

module b17_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P1_MEMORYFETCH_REG_SCAN_IN, 
        DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, 
        DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, 
        DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, 
        DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, 
        DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, 
        DATAI_0_, HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_,
         DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_,
         DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_,
         DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_,
         DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_,
         DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_,
         HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN,
         P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN,
         P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN,
         P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN,
         P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN,
         P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN,
         P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN,
         P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN,
         P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN,
         P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN,
         P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN,
         P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN,
         P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN,
         P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN,
         P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN,
         P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN,
         P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN,
         P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN,
         P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN,
         P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN,
         P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN,
         P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN,
         P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN,
         P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN,
         P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN,
         P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN,
         P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN,
         P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN,
         P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN,
         P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN,
         P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN,
         P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN,
         P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN,
         P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN,
         P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN,
         P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN,
         P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN,
         P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN,
         P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN,
         P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN,
         P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN,
         P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN,
         P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN,
         P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN,
         P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN,
         P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN,
         P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN,
         P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN,
         P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN,
         P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN,
         P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910,
         n11911, n11912, n11913, n11914, n11915, n11916, n11917, n11918,
         n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
         n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934,
         n11935, n11936, n11937, n11938, n11939, n11940, n11941, n11942,
         n11943, n11944, n11945, n11946, n11947, n11948, n11949, n11950,
         n11951, n11952, n11953, n11954, n11955, n11956, n11957, n11958,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974,
         n11975, n11976, n11977, n11978, n11979, n11980, n11981, n11982,
         n11983, n11984, n11985, n11986, n11987, n11988, n11989, n11990,
         n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
         n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006,
         n12007, n12008, n12009, n12010, n12011, n12012, n12013, n12014,
         n12015, n12016, n12017, n12018, n12019, n12020, n12021, n12022,
         n12023, n12024, n12025, n12026, n12027, n12028, n12029, n12030,
         n12031, n12032, n12033, n12034, n12035, n12036, n12037, n12038,
         n12039, n12040, n12041, n12042, n12043, n12044, n12045, n12046,
         n12047, n12048, n12049, n12050, n12051, n12052, n12053, n12054,
         n12055, n12056, n12057, n12058, n12059, n12060, n12061, n12062,
         n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
         n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078,
         n12079, n12080, n12081, n12082, n12083, n12084, n12085, n12086,
         n12087, n12088, n12089, n12090, n12091, n12092, n12093, n12094,
         n12095, n12096, n12097, n12098, n12099, n12100, n12101, n12102,
         n12103, n12104, n12105, n12106, n12107, n12108, n12109, n12110,
         n12111, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
         n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12126,
         n12127, n12128, n12129, n12130, n12131, n12132, n12133, n12134,
         n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142,
         n12143, n12144, n12145, n12146, n12147, n12148, n12149, n12150,
         n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
         n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166,
         n12167, n12168, n12169, n12170, n12171, n12172, n12173, n12174,
         n12175, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12185, n12186, n12187, n12188, n12189, n12190,
         n12191, n12192, n12193, n12194, n12195, n12196, n12197, n12198,
         n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
         n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214,
         n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
         n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230,
         n12231, n12232, n12233, n12234, n12235, n12236, n12237, n12238,
         n12239, n12240, n12241, n12242, n12243, n12244, n12245, n12246,
         n12247, n12248, n12249, n12250, n12251, n12252, n12253, n12254,
         n12255, n12256, n12257, n12258, n12259, n12260, n12261, n12262,
         n12263, n12264, n12265, n12266, n12267, n12268, n12269, n12270,
         n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
         n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286,
         n12287, n12288, n12289, n12290, n12291, n12292, n12293, n12294,
         n12295, n12296, n12297, n12298, n12299, n12300, n12301, n12302,
         n12303, n12304, n12305, n12306, n12307, n12308, n12309, n12310,
         n12311, n12312, n12313, n12314, n12315, n12316, n12317, n12318,
         n12319, n12320, n12321, n12322, n12323, n12324, n12325, n12326,
         n12327, n12328, n12329, n12330, n12331, n12332, n12333, n12334,
         n12335, n12336, n12337, n12338, n12339, n12340, n12341, n12342,
         n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
         n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358,
         n12359, n12360, n12361, n12362, n12363, n12364, n12365, n12366,
         n12367, n12368, n12369, n12370, n12371, n12372, n12373, n12374,
         n12375, n12376, n12377, n12378, n12379, n12380, n12381, n12382,
         n12383, n12384, n12385, n12386, n12387, n12388, n12389, n12390,
         n12391, n12392, n12393, n12394, n12395, n12396, n12397, n12398,
         n12399, n12400, n12401, n12402, n12403, n12404, n12405, n12406,
         n12407, n12408, n12409, n12410, n12411, n12412, n12413, n12414,
         n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
         n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430,
         n12431, n12432, n12433, n12434, n12435, n12436, n12437, n12438,
         n12439, n12440, n12441, n12442, n12443, n12444, n12445, n12446,
         n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
         n12455, n12456, n12457, n12458, n12459, n12460, n12461, n12462,
         n12463, n12464, n12465, n12466, n12467, n12468, n12469, n12470,
         n12471, n12472, n12473, n12474, n12475, n12476, n12477, n12478,
         n12479, n12480, n12481, n12482, n12483, n12484, n12485, n12486,
         n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
         n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502,
         n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510,
         n12511, n12512, n12513, n12514, n12515, n12516, n12517, n12518,
         n12519, n12520, n12521, n12522, n12523, n12524, n12525, n12526,
         n12527, n12528, n12529, n12530, n12531, n12532, n12533, n12534,
         n12535, n12536, n12537, n12538, n12539, n12540, n12541, n12542,
         n12543, n12544, n12545, n12546, n12547, n12548, n12549, n12550,
         n12551, n12552, n12553, n12554, n12555, n12556, n12557, n12558,
         n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
         n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574,
         n12575, n12576, n12577, n12578, n12579, n12580, n12581, n12582,
         n12583, n12584, n12585, n12586, n12587, n12588, n12589, n12590,
         n12591, n12592, n12593, n12594, n12595, n12596, n12597, n12598,
         n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
         n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614,
         n12615, n12616, n12617, n12618, n12619, n12620, n12621, n12622,
         n12623, n12624, n12625, n12626, n12627, n12628, n12629, n12630,
         n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
         n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646,
         n12647, n12648, n12649, n12650, n12651, n12652, n12653, n12654,
         n12655, n12656, n12657, n12658, n12659, n12660, n12661, n12662,
         n12663, n12664, n12665, n12666, n12667, n12668, n12669, n12670,
         n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
         n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686,
         n12687, n12688, n12689, n12690, n12691, n12692, n12693, n12694,
         n12695, n12696, n12697, n12698, n12699, n12700, n12701, n12702,
         n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
         n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718,
         n12719, n12720, n12721, n12722, n12723, n12724, n12725, n12726,
         n12727, n12728, n12729, n12730, n12731, n12732, n12733, n12734,
         n12735, n12736, n12737, n12738, n12739, n12740, n12741, n12742,
         n12743, n12744, n12745, n12746, n12747, n12748, n12749, n12750,
         n12751, n12752, n12753, n12754, n12755, n12756, n12757, n12758,
         n12759, n12760, n12761, n12762, n12763, n12764, n12765, n12766,
         n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
         n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782,
         n12783, n12784, n12785, n12786, n12787, n12788, n12789, n12790,
         n12791, n12792, n12793, n12794, n12795, n12796, n12797, n12798,
         n12799, n12800, n12801, n12802, n12803, n12804, n12805, n12806,
         n12807, n12808, n12809, n12810, n12811, n12812, n12813, n12814,
         n12815, n12816, n12817, n12818, n12819, n12820, n12821, n12822,
         n12823, n12824, n12825, n12826, n12827, n12828, n12829, n12830,
         n12831, n12832, n12833, n12834, n12835, n12836, n12837, n12838,
         n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
         n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854,
         n12855, n12856, n12857, n12858, n12859, n12860, n12861, n12862,
         n12863, n12864, n12865, n12866, n12867, n12868, n12869, n12870,
         n12871, n12872, n12873, n12874, n12875, n12876, n12877, n12878,
         n12879, n12880, n12881, n12882, n12883, n12884, n12885, n12886,
         n12887, n12888, n12889, n12890, n12891, n12892, n12893, n12894,
         n12895, n12896, n12897, n12898, n12899, n12900, n12901, n12902,
         n12903, n12904, n12905, n12906, n12907, n12908, n12909, n12910,
         n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
         n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926,
         n12927, n12928, n12929, n12930, n12931, n12932, n12933, n12934,
         n12935, n12936, n12937, n12938, n12939, n12940, n12941, n12942,
         n12943, n12944, n12945, n12946, n12947, n12948, n12949, n12950,
         n12951, n12952, n12953, n12954, n12955, n12956, n12957, n12958,
         n12959, n12960, n12961, n12962, n12963, n12964, n12965, n12966,
         n12967, n12968, n12969, n12970, n12971, n12972, n12973, n12974,
         n12975, n12976, n12977, n12978, n12979, n12980, n12981, n12982,
         n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
         n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998,
         n12999, n13000, n13001, n13002, n13003, n13004, n13005, n13006,
         n13007, n13008, n13009, n13010, n13011, n13012, n13013, n13014,
         n13015, n13016, n13017, n13018, n13019, n13020, n13021, n13022,
         n13023, n13024, n13025, n13026, n13027, n13028, n13029, n13030,
         n13031, n13032, n13033, n13034, n13035, n13036, n13037, n13038,
         n13039, n13040, n13041, n13042, n13043, n13044, n13045, n13046,
         n13047, n13048, n13049, n13050, n13051, n13052, n13053, n13054,
         n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
         n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070,
         n13071, n13072, n13073, n13074, n13075, n13076, n13077, n13078,
         n13079, n13080, n13081, n13082, n13083, n13084, n13085, n13086,
         n13087, n13088, n13089, n13090, n13091, n13092, n13093, n13094,
         n13095, n13096, n13097, n13098, n13099, n13100, n13101, n13102,
         n13103, n13104, n13105, n13106, n13107, n13108, n13109, n13110,
         n13111, n13112, n13113, n13114, n13115, n13116, n13117, n13118,
         n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
         n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
         n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142,
         n13143, n13144, n13145, n13146, n13147, n13148, n13149, n13150,
         n13151, n13152, n13153, n13154, n13155, n13156, n13157, n13158,
         n13159, n13160, n13161, n13162, n13163, n13164, n13165, n13166,
         n13167, n13168, n13169, n13170, n13171, n13172, n13173, n13174,
         n13175, n13176, n13177, n13178, n13179, n13180, n13181, n13182,
         n13183, n13184, n13185, n13186, n13187, n13188, n13189, n13190,
         n13191, n13192, n13193, n13194, n13195, n13196, n13197, n13198,
         n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
         n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214,
         n13215, n13216, n13217, n13218, n13219, n13220, n13221, n13222,
         n13223, n13224, n13225, n13226, n13227, n13228, n13229, n13230,
         n13231, n13232, n13233, n13234, n13235, n13236, n13237, n13238,
         n13239, n13240, n13241, n13242, n13243, n13244, n13245, n13246,
         n13247, n13248, n13249, n13250, n13251, n13252, n13253, n13254,
         n13255, n13256, n13257, n13258, n13259, n13260, n13261, n13262,
         n13263, n13264, n13265, n13266, n13267, n13268, n13269, n13270,
         n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
         n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286,
         n13287, n13288, n13289, n13290, n13291, n13292, n13293, n13294,
         n13295, n13296, n13297, n13298, n13299, n13300, n13301, n13302,
         n13303, n13304, n13305, n13306, n13307, n13308, n13309, n13310,
         n13311, n13312, n13313, n13314, n13315, n13316, n13317, n13318,
         n13319, n13320, n13321, n13322, n13323, n13324, n13325, n13326,
         n13327, n13328, n13329, n13330, n13331, n13332, n13333, n13334,
         n13335, n13336, n13337, n13338, n13339, n13340, n13341, n13342,
         n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
         n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358,
         n13359, n13360, n13361, n13362, n13363, n13364, n13365, n13366,
         n13367, n13368, n13369, n13370, n13371, n13372, n13373, n13374,
         n13375, n13376, n13377, n13378, n13379, n13380, n13381, n13382,
         n13383, n13384, n13385, n13386, n13387, n13388, n13389, n13390,
         n13391, n13392, n13393, n13394, n13395, n13396, n13397, n13398,
         n13399, n13400, n13401, n13402, n13403, n13404, n13405, n13406,
         n13407, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
         n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422,
         n13423, n13424, n13425, n13426, n13427, n13428, n13429, n13430,
         n13431, n13432, n13433, n13434, n13435, n13436, n13437, n13438,
         n13439, n13440, n13441, n13442, n13443, n13444, n13445, n13446,
         n13447, n13448, n13449, n13450, n13451, n13452, n13453, n13454,
         n13455, n13456, n13457, n13458, n13459, n13460, n13461, n13462,
         n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
         n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478,
         n13479, n13480, n13481, n13482, n13483, n13484, n13485, n13486,
         n13487, n13488, n13489, n13490, n13491, n13492, n13493, n13494,
         n13495, n13496, n13497, n13498, n13499, n13500, n13501, n13502,
         n13503, n13504, n13505, n13506, n13507, n13508, n13509, n13510,
         n13511, n13512, n13513, n13514, n13515, n13516, n13517, n13518,
         n13519, n13520, n13521, n13522, n13523, n13524, n13525, n13526,
         n13527, n13528, n13529, n13530, n13531, n13532, n13533, n13534,
         n13535, n13536, n13537, n13538, n13539, n13540, n13541, n13542,
         n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
         n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558,
         n13559, n13560, n13561, n13562, n13563, n13564, n13565, n13566,
         n13567, n13568, n13569, n13570, n13571, n13572, n13573, n13574,
         n13575, n13576, n13577, n13578, n13579, n13580, n13581, n13582,
         n13583, n13584, n13585, n13586, n13587, n13588, n13589, n13590,
         n13591, n13592, n13593, n13594, n13595, n13596, n13597, n13598,
         n13599, n13600, n13601, n13602, n13603, n13604, n13605, n13606,
         n13607, n13608, n13609, n13610, n13611, n13612, n13613, n13614,
         n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
         n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630,
         n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
         n13639, n13640, n13641, n13642, n13643, n13644, n13645, n13646,
         n13647, n13648, n13649, n13650, n13651, n13652, n13653, n13654,
         n13655, n13656, n13657, n13658, n13659, n13660, n13661, n13662,
         n13663, n13664, n13665, n13666, n13667, n13668, n13669, n13670,
         n13671, n13672, n13673, n13674, n13675, n13676, n13677, n13678,
         n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
         n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
         n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702,
         n13703, n13704, n13705, n13706, n13707, n13708, n13709, n13710,
         n13711, n13712, n13713, n13714, n13715, n13716, n13717, n13718,
         n13719, n13720, n13721, n13722, n13723, n13724, n13725, n13726,
         n13727, n13728, n13729, n13730, n13731, n13732, n13733, n13734,
         n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742,
         n13743, n13744, n13745, n13746, n13747, n13748, n13749, n13750,
         n13751, n13752, n13753, n13754, n13755, n13756, n13757, n13758,
         n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
         n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774,
         n13775, n13776, n13777, n13778, n13779, n13780, n13781, n13782,
         n13783, n13784, n13785, n13786, n13787, n13788, n13789, n13790,
         n13791, n13792, n13793, n13794, n13795, n13796, n13797, n13798,
         n13799, n13800, n13801, n13802, n13803, n13804, n13805, n13806,
         n13807, n13808, n13809, n13810, n13811, n13812, n13813, n13814,
         n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822,
         n13823, n13824, n13825, n13826, n13827, n13828, n13829, n13830,
         n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
         n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846,
         n13847, n13848, n13849, n13850, n13851, n13852, n13853, n13854,
         n13855, n13856, n13857, n13858, n13859, n13860, n13861, n13862,
         n13863, n13864, n13865, n13866, n13867, n13868, n13869, n13870,
         n13871, n13872, n13873, n13874, n13875, n13876, n13877, n13878,
         n13879, n13880, n13881, n13882, n13883, n13884, n13885, n13886,
         n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894,
         n13895, n13896, n13897, n13898, n13899, n13900, n13901, n13902,
         n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
         n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918,
         n13919, n13920, n13921, n13922, n13923, n13924, n13925, n13926,
         n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
         n13935, n13936, n13937, n13938, n13939, n13940, n13941, n13942,
         n13943, n13944, n13945, n13946, n13947, n13948, n13949, n13950,
         n13951, n13952, n13953, n13954, n13955, n13956, n13957, n13958,
         n13959, n13960, n13961, n13962, n13963, n13964, n13965, n13966,
         n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974,
         n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
         n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990,
         n13991, n13992, n13993, n13994, n13995, n13996, n13997, n13998,
         n13999, n14000, n14001, n14002, n14003, n14004, n14005, n14006,
         n14007, n14008, n14009, n14010, n14011, n14012, n14013, n14014,
         n14015, n14016, n14017, n14018, n14019, n14020, n14021, n14022,
         n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030,
         n14031, n14032, n14033, n14034, n14035, n14036, n14037, n14038,
         n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046,
         n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
         n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062,
         n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
         n14071, n14072, n14073, n14074, n14075, n14076, n14077, n14078,
         n14079, n14080, n14081, n14082, n14083, n14084, n14085, n14086,
         n14087, n14088, n14089, n14090, n14091, n14092, n14093, n14094,
         n14095, n14096, n14097, n14098, n14099, n14100, n14101, n14102,
         n14103, n14104, n14105, n14106, n14107, n14108, n14109, n14110,
         n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118,
         n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126,
         n14127, n14128, n14129, n14130, n14131, n14132, n14133, n14134,
         n14135, n14136, n14137, n14138, n14139, n14140, n14141, n14142,
         n14143, n14144, n14145, n14146, n14147, n14148, n14149, n14150,
         n14151, n14152, n14153, n14154, n14155, n14156, n14157, n14158,
         n14159, n14160, n14161, n14162, n14163, n14164, n14165, n14166,
         n14167, n14168, n14169, n14170, n14171, n14172, n14173, n14174,
         n14175, n14176, n14177, n14178, n14179, n14180, n14181, n14182,
         n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190,
         n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198,
         n14199, n14200, n14201, n14202, n14203, n14204, n14205, n14206,
         n14207, n14208, n14209, n14210, n14211, n14212, n14213, n14214,
         n14215, n14216, n14217, n14218, n14219, n14220, n14221, n14222,
         n14223, n14224, n14225, n14226, n14227, n14228, n14229, n14230,
         n14231, n14232, n14233, n14234, n14235, n14236, n14237, n14238,
         n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
         n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
         n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262,
         n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270,
         n14271, n14272, n14273, n14274, n14275, n14276, n14277, n14278,
         n14279, n14280, n14281, n14282, n14283, n14284, n14285, n14286,
         n14287, n14288, n14289, n14290, n14291, n14292, n14293, n14294,
         n14295, n14296, n14297, n14298, n14299, n14300, n14301, n14302,
         n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14310,
         n14311, n14312, n14313, n14314, n14315, n14316, n14317, n14318,
         n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
         n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334,
         n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342,
         n14343, n14344, n14345, n14346, n14347, n14348, n14349, n14350,
         n14351, n14352, n14353, n14354, n14355, n14356, n14357, n14358,
         n14359, n14360, n14361, n14362, n14363, n14364, n14365, n14366,
         n14367, n14368, n14369, n14370, n14371, n14372, n14373, n14374,
         n14375, n14376, n14377, n14378, n14379, n14380, n14381, n14382,
         n14383, n14384, n14385, n14386, n14387, n14388, n14389, n14390,
         n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
         n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406,
         n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414,
         n14415, n14416, n14417, n14418, n14419, n14420, n14421, n14422,
         n14423, n14424, n14425, n14426, n14427, n14428, n14429, n14430,
         n14431, n14432, n14433, n14434, n14435, n14436, n14437, n14438,
         n14439, n14440, n14441, n14442, n14443, n14444, n14445, n14446,
         n14447, n14448, n14449, n14450, n14451, n14452, n14453, n14454,
         n14455, n14456, n14457, n14458, n14459, n14460, n14461, n14462,
         n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
         n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478,
         n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486,
         n14487, n14488, n14489, n14490, n14491, n14492, n14493, n14494,
         n14495, n14496, n14497, n14498, n14499, n14500, n14501, n14502,
         n14503, n14504, n14505, n14506, n14507, n14508, n14509, n14510,
         n14511, n14512, n14513, n14514, n14515, n14516, n14517, n14518,
         n14519, n14520, n14521, n14522, n14523, n14524, n14525, n14526,
         n14527, n14528, n14529, n14530, n14531, n14532, n14533, n14534,
         n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
         n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550,
         n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558,
         n14559, n14560, n14561, n14562, n14563, n14564, n14565, n14566,
         n14567, n14568, n14569, n14570, n14571, n14572, n14573, n14574,
         n14575, n14576, n14577, n14578, n14579, n14580, n14581, n14582,
         n14583, n14584, n14585, n14586, n14587, n14588, n14589, n14590,
         n14591, n14592, n14593, n14594, n14595, n14596, n14597, n14598,
         n14599, n14600, n14601, n14602, n14603, n14604, n14605, n14606,
         n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
         n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622,
         n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630,
         n14631, n14632, n14633, n14634, n14635, n14636, n14637, n14638,
         n14639, n14640, n14641, n14642, n14643, n14644, n14645, n14646,
         n14647, n14648, n14649, n14650, n14651, n14652, n14653, n14654,
         n14655, n14656, n14657, n14658, n14659, n14660, n14661, n14662,
         n14663, n14664, n14665, n14666, n14667, n14668, n14669, n14670,
         n14671, n14672, n14673, n14674, n14675, n14676, n14677, n14678,
         n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
         n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694,
         n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702,
         n14703, n14704, n14705, n14706, n14707, n14708, n14709, n14710,
         n14711, n14712, n14713, n14714, n14715, n14716, n14717, n14718,
         n14719, n14720, n14721, n14722, n14723, n14724, n14725, n14726,
         n14727, n14728, n14729, n14730, n14731, n14732, n14733, n14734,
         n14735, n14736, n14737, n14738, n14739, n14740, n14741, n14742,
         n14743, n14744, n14745, n14746, n14747, n14748, n14749, n14750,
         n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
         n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766,
         n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
         n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782,
         n14783, n14784, n14785, n14786, n14787, n14788, n14789, n14790,
         n14791, n14792, n14793, n14794, n14795, n14796, n14797, n14798,
         n14799, n14800, n14801, n14802, n14803, n14804, n14805, n14806,
         n14807, n14808, n14809, n14810, n14811, n14812, n14813, n14814,
         n14815, n14816, n14817, n14818, n14819, n14820, n14821, n14822,
         n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830,
         n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838,
         n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846,
         n14847, n14848, n14849, n14850, n14851, n14852, n14853, n14854,
         n14855, n14856, n14857, n14858, n14859, n14860, n14861, n14862,
         n14863, n14864, n14865, n14866, n14867, n14868, n14869, n14870,
         n14871, n14872, n14873, n14874, n14875, n14876, n14877, n14878,
         n14879, n14880, n14881, n14882, n14883, n14884, n14885, n14886,
         n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
         n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902,
         n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910,
         n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918,
         n14919, n14920, n14921, n14922, n14923, n14924, n14925, n14926,
         n14927, n14928, n14929, n14930, n14931, n14932, n14933, n14934,
         n14935, n14936, n14937, n14938, n14939, n14940, n14941, n14942,
         n14943, n14944, n14945, n14946, n14947, n14948, n14949, n14950,
         n14951, n14952, n14953, n14954, n14955, n14956, n14957, n14958,
         n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
         n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974,
         n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982,
         n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990,
         n14991, n14992, n14993, n14994, n14995, n14996, n14997, n14998,
         n14999, n15000, n15001, n15002, n15003, n15004, n15005, n15006,
         n15007, n15008, n15009, n15010, n15011, n15012, n15013, n15014,
         n15015, n15016, n15017, n15018, n15019, n15020, n15021, n15022,
         n15023, n15024, n15025, n15026, n15027, n15028, n15029, n15030,
         n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
         n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046,
         n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054,
         n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062,
         n15063, n15064, n15065, n15066, n15067, n15068, n15069, n15070,
         n15071, n15072, n15073, n15074, n15075, n15076, n15077, n15078,
         n15079, n15080, n15081, n15082, n15083, n15084, n15085, n15086,
         n15087, n15088, n15089, n15090, n15091, n15092, n15093, n15094,
         n15095, n15096, n15097, n15098, n15099, n15100, n15101, n15102,
         n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
         n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118,
         n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126,
         n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134,
         n15135, n15136, n15137, n15138, n15139, n15140, n15141, n15142,
         n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150,
         n15151, n15152, n15153, n15154, n15155, n15156, n15157, n15158,
         n15159, n15160, n15161, n15162, n15163, n15164, n15165, n15166,
         n15167, n15168, n15169, n15170, n15171, n15172, n15173, n15174,
         n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
         n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190,
         n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198,
         n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206,
         n15207, n15208, n15209, n15210, n15211, n15212, n15213, n15214,
         n15215, n15216, n15217, n15218, n15219, n15220, n15221, n15222,
         n15223, n15224, n15225, n15226, n15227, n15228, n15229, n15230,
         n15231, n15232, n15233, n15234, n15235, n15236, n15237, n15238,
         n15239, n15240, n15241, n15242, n15243, n15244, n15245, n15246,
         n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
         n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262,
         n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270,
         n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278,
         n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286,
         n15287, n15288, n15289, n15290, n15291, n15292, n15293, n15294,
         n15295, n15296, n15297, n15298, n15299, n15300, n15301, n15302,
         n15303, n15304, n15305, n15306, n15307, n15308, n15309, n15310,
         n15311, n15312, n15313, n15314, n15315, n15316, n15317, n15318,
         n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
         n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334,
         n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342,
         n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350,
         n15351, n15352, n15353, n15354, n15355, n15356, n15357, n15358,
         n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
         n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374,
         n15375, n15376, n15377, n15378, n15379, n15380, n15381, n15382,
         n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390,
         n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
         n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406,
         n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414,
         n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422,
         n15423, n15424, n15425, n15426, n15427, n15428, n15429, n15430,
         n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
         n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446,
         n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454,
         n15455, n15456, n15457, n15458, n15459, n15460, n15461, n15462,
         n15463, n15464, n15465, n15466, n15467, n15468, n15469, n15470,
         n15471, n15472, n15473, n15474, n15475, n15476, n15477, n15478,
         n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486,
         n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494,
         n15495, n15496, n15497, n15498, n15499, n15500, n15501, n15502,
         n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
         n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518,
         n15519, n15520, n15521, n15522, n15523, n15524, n15525, n15526,
         n15527, n15528, n15529, n15530, n15531, n15532, n15533, n15534,
         n15535, n15536, n15537, n15538, n15539, n15540, n15541, n15542,
         n15543, n15544, n15545, n15546, n15547, n15548, n15549, n15550,
         n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558,
         n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566,
         n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
         n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
         n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590,
         n15591, n15592, n15593, n15594, n15595, n15596, n15597, n15598,
         n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606,
         n15607, n15608, n15609, n15610, n15611, n15612, n15613, n15614,
         n15615, n15616, n15617, n15618, n15619, n15620, n15621, n15622,
         n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630,
         n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638,
         n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
         n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654,
         n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662,
         n15663, n15664, n15665, n15666, n15667, n15668, n15669, n15670,
         n15671, n15672, n15673, n15674, n15675, n15676, n15677, n15678,
         n15679, n15680, n15681, n15682, n15683, n15684, n15685, n15686,
         n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694,
         n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702,
         n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710,
         n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718,
         n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726,
         n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15734,
         n15735, n15736, n15737, n15738, n15739, n15740, n15741, n15742,
         n15743, n15744, n15745, n15746, n15747, n15748, n15749, n15750,
         n15751, n15752, n15753, n15754, n15755, n15756, n15757, n15758,
         n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766,
         n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774,
         n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782,
         n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790,
         n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798,
         n15799, n15800, n15801, n15802, n15803, n15804, n15805, n15806,
         n15807, n15808, n15809, n15810, n15811, n15812, n15813, n15814,
         n15815, n15816, n15817, n15818, n15819, n15820, n15821, n15822,
         n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830,
         n15831, n15832, n15833, n15834, n15835, n15836, n15837, n15838,
         n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846,
         n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854,
         n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
         n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870,
         n15871, n15872, n15873, n15874, n15875, n15876, n15877, n15878,
         n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886,
         n15887, n15888, n15889, n15890, n15891, n15892, n15893, n15894,
         n15895, n15896, n15897, n15898, n15899, n15900, n15901, n15902,
         n15903, n15904, n15905, n15906, n15907, n15908, n15909, n15910,
         n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918,
         n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926,
         n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
         n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942,
         n15943, n15944, n15945, n15946, n15947, n15948, n15949, n15950,
         n15951, n15952, n15953, n15954, n15955, n15956, n15957, n15958,
         n15959, n15960, n15961, n15962, n15963, n15964, n15965, n15966,
         n15967, n15968, n15969, n15970, n15971, n15972, n15973, n15974,
         n15975, n15976, n15977, n15978, n15979, n15980, n15981, n15982,
         n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990,
         n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998,
         n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006,
         n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014,
         n16015, n16016, n16017, n16018, n16019, n16020, n16021, n16022,
         n16023, n16024, n16025, n16026, n16027, n16028, n16029, n16030,
         n16031, n16032, n16033, n16034, n16035, n16036, n16037, n16038,
         n16039, n16040, n16041, n16042, n16043, n16044, n16045, n16046,
         n16047, n16048, n16049, n16050, n16051, n16052, n16053, n16054,
         n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062,
         n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070,
         n16071, n16072, n16073, n16074, n16075, n16076, n16077, n16078,
         n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086,
         n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094,
         n16095, n16096, n16097, n16098, n16099, n16100, n16101, n16102,
         n16103, n16104, n16105, n16106, n16107, n16108, n16109, n16110,
         n16111, n16112, n16113, n16114, n16115, n16116, n16117, n16118,
         n16119, n16120, n16121, n16122, n16123, n16124, n16125, n16126,
         n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134,
         n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142,
         n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150,
         n16151, n16152, n16153, n16154, n16155, n16156, n16157, n16158,
         n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
         n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174,
         n16175, n16176, n16177, n16178, n16179, n16180, n16181, n16182,
         n16183, n16184, n16185, n16186, n16187, n16188, n16189, n16190,
         n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198,
         n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206,
         n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214,
         n16215, n16216, n16217, n16218, n16219, n16220, n16221, n16222,
         n16223, n16224, n16225, n16226, n16227, n16228, n16229, n16230,
         n16231, n16232, n16233, n16234, n16235, n16236, n16237, n16238,
         n16239, n16240, n16241, n16242, n16243, n16244, n16245, n16246,
         n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254,
         n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262,
         n16263, n16264, n16265, n16266, n16267, n16268, n16269, n16270,
         n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278,
         n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286,
         n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294,
         n16295, n16296, n16297, n16298, n16299, n16300, n16301, n16302,
         n16303, n16304, n16305, n16306, n16307, n16308, n16309, n16310,
         n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318,
         n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326,
         n16327, n16328, n16329, n16330, n16331, n16332, n16333, n16334,
         n16335, n16336, n16337, n16338, n16339, n16340, n16341, n16342,
         n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350,
         n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358,
         n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366,
         n16367, n16368, n16369, n16370, n16371, n16372, n16373, n16374,
         n16375, n16376, n16377, n16378, n16379, n16380, n16381, n16382,
         n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
         n16391, n16392, n16393, n16394, n16395, n16396, n16397, n16398,
         n16399, n16400, n16401, n16402, n16403, n16404, n16405, n16406,
         n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414,
         n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422,
         n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430,
         n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438,
         n16439, n16440, n16441, n16442, n16443, n16444, n16445, n16446,
         n16447, n16448, n16449, n16450, n16451, n16452, n16453, n16454,
         n16455, n16456, n16457, n16458, n16459, n16460, n16461, n16462,
         n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470,
         n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
         n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486,
         n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494,
         n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502,
         n16503, n16504, n16505, n16506, n16507, n16508, n16509, n16510,
         n16511, n16512, n16513, n16514, n16515, n16516, n16517, n16518,
         n16519, n16520, n16521, n16522, n16523, n16524, n16525, n16526,
         n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534,
         n16535, n16536, n16537, n16538, n16539, n16540, n16541, n16542,
         n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550,
         n16551, n16552, n16553, n16554, n16555, n16556, n16557, n16558,
         n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566,
         n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574,
         n16575, n16576, n16577, n16578, n16579, n16580, n16581, n16582,
         n16583, n16584, n16585, n16586, n16587, n16588, n16589, n16590,
         n16591, n16592, n16593, n16594, n16595, n16596, n16597, n16598,
         n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
         n16607, n16608, n16609, n16610, n16611, n16612, n16613, n16614,
         n16615, n16616, n16617, n16618, n16619, n16620, n16621, n16622,
         n16623, n16624, n16625, n16626, n16627, n16628, n16629, n16630,
         n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638,
         n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646,
         n16647, n16648, n16649, n16650, n16651, n16652, n16653, n16654,
         n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662,
         n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670,
         n16671, n16672, n16673, n16674, n16675, n16676, n16677, n16678,
         n16679, n16680, n16681, n16682, n16683, n16684, n16685, n16686,
         n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694,
         n16695, n16696, n16697, n16698, n16699, n16700, n16701, n16702,
         n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710,
         n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718,
         n16719, n16720, n16721, n16722, n16723, n16724, n16725, n16726,
         n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734,
         n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742,
         n16743, n16744, n16745, n16746, n16747, n16748, n16749, n16750,
         n16751, n16752, n16753, n16754, n16755, n16756, n16757, n16758,
         n16759, n16760, n16761, n16762, n16763, n16764, n16765, n16766,
         n16767, n16768, n16769, n16770, n16771, n16772, n16773, n16774,
         n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782,
         n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790,
         n16791, n16792, n16793, n16794, n16795, n16796, n16797, n16798,
         n16799, n16800, n16801, n16802, n16803, n16804, n16805, n16806,
         n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814,
         n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822,
         n16823, n16824, n16825, n16826, n16827, n16828, n16829, n16830,
         n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838,
         n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846,
         n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854,
         n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862,
         n16863, n16864, n16865, n16866, n16867, n16868, n16869, n16870,
         n16871, n16872, n16873, n16874, n16875, n16876, n16877, n16878,
         n16879, n16880, n16881, n16882, n16883, n16884, n16885, n16886,
         n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894,
         n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16902,
         n16903, n16904, n16905, n16906, n16907, n16908, n16909, n16910,
         n16911, n16912, n16913, n16914, n16915, n16916, n16917, n16918,
         n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926,
         n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934,
         n16935, n16936, n16937, n16938, n16939, n16940, n16941, n16942,
         n16943, n16944, n16945, n16946, n16947, n16948, n16949, n16950,
         n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958,
         n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966,
         n16967, n16968, n16969, n16970, n16971, n16972, n16973, n16974,
         n16975, n16976, n16977, n16978, n16979, n16980, n16981, n16982,
         n16983, n16984, n16985, n16986, n16987, n16988, n16989, n16990,
         n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998,
         n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006,
         n17007, n17008, n17009, n17010, n17011, n17012, n17013, n17014,
         n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022,
         n17023, n17024, n17025, n17026, n17027, n17028, n17029, n17030,
         n17031, n17032, n17033, n17034, n17035, n17036, n17037, n17038,
         n17039, n17040, n17041, n17042, n17043, n17044, n17045, n17046,
         n17047, n17048, n17049, n17050, n17051, n17052, n17053, n17054,
         n17055, n17056, n17057, n17058, n17059, n17060, n17061, n17062,
         n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070,
         n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078,
         n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086,
         n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094,
         n17095, n17096, n17097, n17098, n17099, n17100, n17101, n17102,
         n17103, n17104, n17105, n17106, n17107, n17108, n17109, n17110,
         n17111, n17112, n17113, n17114, n17115, n17116, n17117, n17118,
         n17119, n17120, n17121, n17122, n17123, n17124, n17125, n17126,
         n17127, n17128, n17129, n17130, n17131, n17132, n17133, n17134,
         n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142,
         n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150,
         n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158,
         n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166,
         n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174,
         n17175, n17176, n17177, n17178, n17179, n17180, n17181, n17182,
         n17183, n17184, n17185, n17186, n17187, n17188, n17189, n17190,
         n17191, n17192, n17193, n17194, n17195, n17196, n17197, n17198,
         n17199, n17200, n17201, n17202, n17203, n17204, n17205, n17206,
         n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214,
         n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222,
         n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230,
         n17231, n17232, n17233, n17234, n17235, n17236, n17237, n17238,
         n17239, n17240, n17241, n17242, n17243, n17244, n17245, n17246,
         n17247, n17248, n17249, n17250, n17251, n17252, n17253, n17254,
         n17255, n17256, n17257, n17258, n17259, n17260, n17261, n17262,
         n17263, n17264, n17265, n17266, n17267, n17268, n17269, n17270,
         n17271, n17272, n17273, n17274, n17275, n17276, n17277, n17278,
         n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286,
         n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294,
         n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302,
         n17303, n17304, n17305, n17306, n17307, n17308, n17309, n17310,
         n17311, n17312, n17313, n17314, n17315, n17316, n17317, n17318,
         n17319, n17320, n17321, n17322, n17323, n17324, n17325, n17326,
         n17327, n17328, n17329, n17330, n17331, n17332, n17333, n17334,
         n17335, n17336, n17337, n17338, n17339, n17340, n17341, n17342,
         n17343, n17344, n17345, n17346, n17347, n17348, n17349, n17350,
         n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358,
         n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
         n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374,
         n17375, n17376, n17377, n17378, n17379, n17380, n17381, n17382,
         n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390,
         n17391, n17392, n17393, n17394, n17395, n17396, n17397, n17398,
         n17399, n17400, n17401, n17402, n17403, n17404, n17405, n17406,
         n17407, n17408, n17409, n17410, n17411, n17412, n17413, n17414,
         n17415, n17416, n17417, n17418, n17419, n17420, n17421, n17422,
         n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430,
         n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438,
         n17439, n17440, n17441, n17442, n17443, n17444, n17445, n17446,
         n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454,
         n17455, n17456, n17457, n17458, n17459, n17460, n17461, n17462,
         n17463, n17464, n17465, n17466, n17467, n17468, n17469, n17470,
         n17471, n17472, n17473, n17474, n17475, n17476, n17477, n17478,
         n17479, n17480, n17481, n17482, n17483, n17484, n17485, n17486,
         n17487, n17488, n17489, n17490, n17491, n17492, n17493, n17494,
         n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502,
         n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510,
         n17511, n17512, n17513, n17514, n17515, n17516, n17517, n17518,
         n17519, n17520, n17521, n17522, n17523, n17524, n17525, n17526,
         n17527, n17528, n17529, n17530, n17531, n17532, n17533, n17534,
         n17535, n17536, n17537, n17538, n17539, n17540, n17541, n17542,
         n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550,
         n17551, n17552, n17553, n17554, n17555, n17556, n17557, n17558,
         n17559, n17560, n17561, n17562, n17563, n17564, n17565, n17566,
         n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574,
         n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582,
         n17583, n17584, n17585, n17586, n17587, n17588, n17589, n17590,
         n17591, n17592, n17593, n17594, n17595, n17596, n17597, n17598,
         n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17606,
         n17607, n17608, n17609, n17610, n17611, n17612, n17613, n17614,
         n17615, n17616, n17617, n17618, n17619, n17620, n17621, n17622,
         n17623, n17624, n17625, n17626, n17627, n17628, n17629, n17630,
         n17631, n17632, n17633, n17634, n17635, n17636, n17637, n17638,
         n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646,
         n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654,
         n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17662,
         n17663, n17664, n17665, n17666, n17667, n17668, n17669, n17670,
         n17671, n17672, n17673, n17674, n17675, n17676, n17677, n17678,
         n17679, n17680, n17681, n17682, n17683, n17684, n17685, n17686,
         n17687, n17688, n17689, n17690, n17691, n17692, n17693, n17694,
         n17695, n17696, n17697, n17698, n17699, n17700, n17701, n17702,
         n17703, n17704, n17705, n17706, n17707, n17708, n17709, n17710,
         n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718,
         n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782,
         n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
         n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
         n17799, n17800, n17801, n17802, n17803, n17804, n17805, n17806,
         n17807, n17808, n17809, n17810, n17811, n17812, n17813, n17814,
         n17815, n17816, n17817, n17818, n17819, n17820, n17821, n17822,
         n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
         n17831, n17832, n17833, n17834, n17835, n17836, n17837, n17838,
         n17839, n17840, n17841, n17842, n17843, n17844, n17845, n17846,
         n17847, n17848, n17849, n17850, n17851, n17852, n17853, n17854,
         n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862,
         n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870,
         n17871, n17872, n17873, n17874, n17875, n17876, n17877, n17878,
         n17879, n17880, n17881, n17882, n17883, n17884, n17885, n17886,
         n17887, n17888, n17889, n17890, n17891, n17892, n17893, n17894,
         n17895, n17896, n17897, n17898, n17899, n17900, n17901, n17902,
         n17903, n17904, n17905, n17906, n17907, n17908, n17909, n17910,
         n17911, n17912, n17913, n17914, n17915, n17916, n17917, n17918,
         n17919, n17920, n17921, n17922, n17923, n17924, n17925, n17926,
         n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934,
         n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942,
         n17943, n17944, n17945, n17946, n17947, n17948, n17949, n17950,
         n17951, n17952, n17953, n17954, n17955, n17956, n17957, n17958,
         n17959, n17960, n17961, n17962, n17963, n17964, n17965, n17966,
         n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17974,
         n17975, n17976, n17977, n17978, n17979, n17980, n17981, n17982,
         n17983, n17984, n17985, n17986, n17987, n17988, n17989, n17990,
         n17991, n17992, n17993, n17994, n17995, n17996, n17997, n17998,
         n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006,
         n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014,
         n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022,
         n18023, n18024, n18025, n18026, n18027, n18028, n18029, n18030,
         n18031, n18032, n18033, n18034, n18035, n18036, n18037, n18038,
         n18039, n18040, n18041, n18042, n18043, n18044, n18045, n18046,
         n18047, n18048, n18049, n18050, n18051, n18052, n18053, n18054,
         n18055, n18056, n18057, n18058, n18059, n18060, n18061, n18062,
         n18063, n18064, n18065, n18066, n18067, n18068, n18069, n18070,
         n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078,
         n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086,
         n18087, n18088, n18089, n18090, n18091, n18092, n18093, n18094,
         n18095, n18096, n18097, n18098, n18099, n18100, n18101, n18102,
         n18103, n18104, n18105, n18106, n18107, n18108, n18109, n18110,
         n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
         n18119, n18120, n18121, n18122, n18123, n18124, n18125, n18126,
         n18127, n18128, n18129, n18130, n18131, n18132, n18133, n18134,
         n18135, n18136, n18137, n18138, n18139, n18140, n18141, n18142,
         n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150,
         n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158,
         n18159, n18160, n18161, n18162, n18163, n18164, n18165, n18166,
         n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
         n18175, n18176, n18177, n18178, n18179, n18180, n18181, n18182,
         n18183, n18184, n18185, n18186, n18187, n18188, n18189, n18190,
         n18191, n18192, n18193, n18194, n18195, n18196, n18197, n18198,
         n18199, n18200, n18201, n18202, n18203, n18204, n18205, n18206,
         n18207, n18208, n18209, n18210, n18211, n18212, n18213, n18214,
         n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222,
         n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
         n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238,
         n18239, n18240, n18241, n18242, n18243, n18244, n18245, n18246,
         n18247, n18248, n18249, n18250, n18251, n18252, n18253, n18254,
         n18255, n18256, n18257, n18258, n18259, n18260, n18261, n18262,
         n18263, n18264, n18265, n18266, n18267, n18268, n18269, n18270,
         n18271, n18272, n18273, n18274, n18275, n18276, n18277, n18278,
         n18279, n18280, n18281, n18282, n18283, n18284, n18285, n18286,
         n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294,
         n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302,
         n18303, n18304, n18305, n18306, n18307, n18308, n18309, n18310,
         n18311, n18312, n18313, n18314, n18315, n18316, n18317, n18318,
         n18319, n18320, n18321, n18322, n18323, n18324, n18325, n18326,
         n18327, n18328, n18329, n18330, n18331, n18332, n18333, n18334,
         n18335, n18336, n18337, n18338, n18339, n18340, n18341, n18342,
         n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
         n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358,
         n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366,
         n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374,
         n18375, n18376, n18377, n18378, n18379, n18380, n18381, n18382,
         n18383, n18384, n18385, n18386, n18387, n18388, n18389, n18390,
         n18391, n18392, n18393, n18394, n18395, n18396, n18397, n18398,
         n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
         n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414,
         n18415, n18416, n18417, n18418, n18419, n18420, n18421, n18422,
         n18423, n18424, n18425, n18426, n18427, n18428, n18429, n18430,
         n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438,
         n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446,
         n18447, n18448, n18449, n18450, n18451, n18452, n18453, n18454,
         n18455, n18456, n18457, n18458, n18459, n18460, n18461, n18462,
         n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470,
         n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478,
         n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486,
         n18487, n18488, n18489, n18490, n18491, n18492, n18493, n18494,
         n18495, n18496, n18497, n18498, n18499, n18500, n18501, n18502,
         n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510,
         n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518,
         n18519, n18520, n18521, n18522, n18523, n18524, n18525, n18526,
         n18527, n18528, n18529, n18530, n18531, n18532, n18533, n18534,
         n18535, n18536, n18537, n18538, n18539, n18540, n18541, n18542,
         n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550,
         n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558,
         n18559, n18560, n18561, n18562, n18563, n18564, n18565, n18566,
         n18567, n18568, n18569, n18570, n18571, n18572, n18573, n18574,
         n18575, n18576, n18577, n18578, n18579, n18580, n18581, n18582,
         n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
         n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598,
         n18599, n18600, n18601, n18602, n18603, n18604, n18605, n18606,
         n18607, n18608, n18609, n18610, n18611, n18612, n18613, n18614,
         n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622,
         n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630,
         n18631, n18632, n18633, n18634, n18635, n18636, n18637, n18638,
         n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
         n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654,
         n18655, n18656, n18657, n18658, n18659, n18660, n18661, n18662,
         n18663, n18664, n18665, n18666, n18667, n18668, n18669, n18670,
         n18671, n18672, n18673, n18674, n18675, n18676, n18677, n18678,
         n18679, n18680, n18681, n18682, n18683, n18684, n18685, n18686,
         n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694,
         n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702,
         n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710,
         n18711, n18712, n18713, n18714, n18715, n18716, n18717, n18718,
         n18719, n18720, n18721, n18722, n18723, n18724, n18725, n18726,
         n18727, n18728, n18729, n18730, n18731, n18732, n18733, n18734,
         n18735, n18736, n18737, n18738, n18739, n18740, n18741, n18742,
         n18743, n18744, n18745, n18746, n18747, n18748, n18749, n18750,
         n18751, n18752, n18753, n18754, n18755, n18756, n18757, n18758,
         n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766,
         n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774,
         n18775, n18776, n18777, n18778, n18779, n18780, n18781, n18782,
         n18783, n18784, n18785, n18786, n18787, n18788, n18789, n18790,
         n18791, n18792, n18793, n18794, n18795, n18796, n18797, n18798,
         n18799, n18800, n18801, n18802, n18803, n18804, n18805, n18806,
         n18807, n18808, n18809, n18810, n18811, n18812, n18813, n18814,
         n18815, n18816, n18817, n18818, n18819, n18820, n18821, n18822,
         n18823, n18824, n18825, n18826, n18827, n18828, n18829, n18830,
         n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838,
         n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846,
         n18847, n18848, n18849, n18850, n18851, n18852, n18853, n18854,
         n18855, n18856, n18857, n18858, n18859, n18860, n18861, n18862,
         n18863, n18864, n18865, n18866, n18867, n18868, n18869, n18870,
         n18871, n18872, n18873, n18874, n18875, n18876, n18877, n18878,
         n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
         n18887, n18888, n18889, n18890, n18891, n18892, n18893, n18894,
         n18895, n18896, n18897, n18898, n18899, n18900, n18901, n18902,
         n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910,
         n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918,
         n18919, n18920, n18921, n18922, n18923, n18924, n18925, n18926,
         n18927, n18928, n18929, n18930, n18931, n18932, n18933, n18934,
         n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942,
         n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950,
         n18951, n18952, n18953, n18954, n18955, n18956, n18957, n18958,
         n18959, n18960, n18961, n18962, n18963, n18964, n18965, n18966,
         n18967, n18968, n18969, n18970, n18971, n18972, n18973, n18974,
         n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982,
         n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990,
         n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
         n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006,
         n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014,
         n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022,
         n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030,
         n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038,
         n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046,
         n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
         n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062,
         n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070,
         n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078,
         n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086,
         n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094,
         n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
         n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110,
         n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118,
         n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
         n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134,
         n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142,
         n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150,
         n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158,
         n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166,
         n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
         n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182,
         n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190,
         n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198,
         n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206,
         n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214,
         n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222,
         n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230,
         n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238,
         n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
         n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254,
         n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262,
         n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
         n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278,
         n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286,
         n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294,
         n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302,
         n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310,
         n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
         n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326,
         n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334,
         n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342,
         n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350,
         n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358,
         n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366,
         n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374,
         n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382,
         n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
         n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398,
         n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406,
         n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
         n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422,
         n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430,
         n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438,
         n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446,
         n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454,
         n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
         n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470,
         n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478,
         n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486,
         n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494,
         n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502,
         n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510,
         n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518,
         n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526,
         n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
         n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542,
         n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550,
         n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
         n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566,
         n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574,
         n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582,
         n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590,
         n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598,
         n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
         n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614,
         n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622,
         n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
         n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638,
         n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
         n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
         n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
         n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
         n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710,
         n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
         n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726,
         n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734,
         n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
         n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
         n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758,
         n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766,
         n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
         n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
         n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
         n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
         n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806,
         n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
         n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
         n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830,
         n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838,
         n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
         n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
         n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
         n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870,
         n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
         n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
         n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902,
         n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
         n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
         n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926,
         n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934,
         n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
         n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
         n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
         n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
         n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
         n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982,
         n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
         n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014,
         n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
         n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
         n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
         n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
         n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
         n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142,
         n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
         n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158,
         n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
         n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
         n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
         n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190,
         n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198,
         n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
         n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
         n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
         n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
         n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
         n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246,
         n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
         n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262,
         n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270,
         n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
         n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
         n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
         n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342,
         n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
         n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
         n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
         n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
         n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
         n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
         n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
         n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
         n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
         n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
         n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
         n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
         n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574,
         n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
         n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590,
         n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
         n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
         n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718,
         n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
         n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734,
         n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742,
         n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
         n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
         n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766,
         n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774,
         n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
         n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790,
         n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
         n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806,
         n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814,
         n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822,
         n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
         n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838,
         n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846,
         n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854,
         n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862,
         n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
         n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878,
         n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886,
         n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894,
         n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
         n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910,
         n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918,
         n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
         n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934,
         n20935, n20936, n20937, n20938, n20939, n20940, n20941, n20942,
         n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950,
         n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958,
         n20959, n20960, n20961, n20962, n20963, n20964, n20965, n20966,
         n20967, n20968, n20969, n20970, n20971, n20972, n20973, n20974,
         n20975, n20976, n20977, n20978, n20979, n20980, n20981, n20982,
         n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990,
         n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998,
         n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006,
         n21007, n21008, n21009, n21010, n21011, n21012, n21013, n21014,
         n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022,
         n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030,
         n21031, n21032, n21033, n21034, n21035, n21036, n21037, n21038,
         n21039, n21040, n21041, n21042, n21043, n21044, n21045, n21046,
         n21047, n21048, n21049, n21050, n21051, n21052, n21053, n21054,
         n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062,
         n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070,
         n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078,
         n21079, n21080, n21081, n21082, n21083, n21084, n21085, n21086,
         n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094,
         n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102,
         n21103, n21104, n21105, n21106, n21107, n21108, n21109, n21110,
         n21111, n21112, n21113, n21114, n21115, n21116, n21117, n21118,
         n21119, n21120, n21121, n21122, n21123, n21124, n21125, n21126,
         n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134,
         n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142,
         n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150,
         n21151, n21152, n21153, n21154, n21155, n21156, n21157, n21158,
         n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166,
         n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174,
         n21175, n21176, n21177, n21178, n21179, n21180, n21181, n21182,
         n21183, n21184, n21185, n21186, n21187, n21188, n21189, n21190,
         n21191, n21192, n21193, n21194, n21195, n21196, n21197, n21198,
         n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206,
         n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214,
         n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222,
         n21223, n21224, n21225, n21226, n21227, n21228, n21229, n21230,
         n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238,
         n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246,
         n21247, n21248, n21249, n21250, n21251, n21252, n21253, n21254,
         n21255, n21256, n21257, n21258, n21259, n21260, n21261, n21262,
         n21263, n21264, n21265, n21266, n21267, n21268, n21269, n21270,
         n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278,
         n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286,
         n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294,
         n21295, n21296, n21297, n21298, n21299, n21300, n21301, n21302,
         n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310,
         n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318,
         n21319, n21320, n21321, n21322, n21323, n21324, n21325, n21326,
         n21327, n21328, n21329, n21330, n21331, n21332, n21333, n21334,
         n21335, n21336, n21337, n21338, n21339, n21340, n21341, n21342,
         n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350,
         n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358,
         n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366,
         n21367, n21368, n21369, n21370, n21371, n21372, n21373, n21374,
         n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382,
         n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390,
         n21391, n21392, n21393, n21394, n21395, n21396, n21397, n21398,
         n21399, n21400, n21401, n21402, n21403, n21404, n21405, n21406,
         n21407, n21408, n21409, n21410, n21411, n21412, n21413, n21414,
         n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422,
         n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430,
         n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438,
         n21439, n21440, n21441, n21442, n21443, n21444, n21445, n21446,
         n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454,
         n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462,
         n21463, n21464, n21465, n21466, n21467, n21468, n21469, n21470,
         n21471, n21472, n21473, n21474, n21475, n21476, n21477, n21478,
         n21479, n21480, n21481, n21482, n21483, n21484, n21485, n21486,
         n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494,
         n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502,
         n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510,
         n21511, n21512, n21513, n21514, n21515, n21516, n21517, n21518,
         n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526,
         n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534,
         n21535, n21536, n21537, n21538, n21539, n21540, n21541, n21542,
         n21543, n21544, n21545, n21546, n21547, n21548, n21549, n21550,
         n21551, n21552, n21553, n21554, n21555, n21556, n21557, n21558,
         n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566,
         n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574,
         n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582,
         n21583, n21584, n21585, n21586, n21587, n21588, n21589, n21590,
         n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598,
         n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21606,
         n21607, n21608, n21609, n21610, n21611, n21612, n21613, n21614,
         n21615, n21616, n21617, n21618, n21619, n21620, n21621, n21622,
         n21623, n21624, n21625, n21626, n21627, n21628, n21629, n21630,
         n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638,
         n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646,
         n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21654,
         n21655, n21656, n21657, n21658, n21659, n21660, n21661, n21662,
         n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21670,
         n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678,
         n21679, n21680, n21681, n21682, n21683, n21684, n21685, n21686,
         n21687, n21688, n21689, n21690, n21691, n21692, n21693, n21694,
         n21695, n21696, n21697, n21698, n21699, n21700, n21701, n21702,
         n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710,
         n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718,
         n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726,
         n21727, n21728, n21729, n21730, n21731, n21732, n21733, n21734,
         n21735, n21736, n21737, n21738, n21739, n21740, n21741, n21742,
         n21743, n21744, n21745, n21746, n21747, n21748, n21749, n21750,
         n21751, n21752, n21753, n21754, n21755, n21756, n21757, n21758,
         n21759, n21760, n21761, n21762, n21763, n21764, n21765, n21766,
         n21767, n21768, n21769, n21770, n21771, n21772, n21773, n21774,
         n21775, n21776, n21777, n21778, n21779, n21780, n21781, n21782,
         n21783, n21784, n21785, n21786, n21787, n21788, n21789, n21790,
         n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21798,
         n21799, n21800, n21801, n21802, n21803, n21804, n21805, n21806,
         n21807, n21808, n21809, n21810, n21811, n21812, n21813, n21814,
         n21815, n21816, n21817, n21818, n21819, n21820, n21821, n21822,
         n21823, n21824, n21825, n21826, n21827, n21828, n21829, n21830,
         n21831, n21832, n21833, n21834, n21835, n21836, n21837, n21838,
         n21839, n21840, n21841, n21842, n21843, n21844, n21845, n21846,
         n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854,
         n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862,
         n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870,
         n21871, n21872, n21873, n21874, n21875, n21876, n21877, n21878,
         n21879, n21880, n21881, n21882, n21883, n21884, n21885, n21886,
         n21887, n21888, n21889, n21890, n21891, n21892, n21893, n21894,
         n21895, n21896, n21897, n21898, n21899, n21900, n21901, n21902,
         n21903, n21904, n21905, n21906, n21907, n21908, n21909, n21910,
         n21911, n21912, n21913, n21914, n21915, n21916, n21917, n21918,
         n21919, n21920, n21921, n21922, n21923, n21924, n21925, n21926,
         n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934,
         n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942,
         n21943, n21944, n21945, n21946, n21947, n21948, n21949, n21950,
         n21951, n21952, n21953, n21954, n21955, n21956, n21957, n21958,
         n21959, n21960, n21961, n21962, n21963, n21964, n21965, n21966,
         n21967, n21968, n21969, n21970, n21971, n21972, n21973, n21974,
         n21975, n21976, n21977, n21978, n21979, n21980, n21981, n21982,
         n21983, n21984, n21985, n21986, n21987, n21988, n21989, n21990,
         n21991, n21992, n21993, n21994, n21995, n21996, n21997, n21998,
         n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006,
         n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014,
         n22015, n22016, n22017, n22018, n22019, n22020, n22021, n22022,
         n22023, n22024, n22025, n22026, n22027, n22028, n22029, n22030,
         n22031, n22032, n22033, n22034, n22035, n22036, n22037, n22038,
         n22039, n22040, n22041, n22042, n22043, n22044, n22045, n22046,
         n22047, n22048, n22049, n22050, n22051, n22052, n22053, n22054,
         n22055, n22056, n22057, n22058, n22059, n22060, n22061, n22062,
         n22063, n22064, n22065, n22066, n22067, n22068, n22069, n22070,
         n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078,
         n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086,
         n22087, n22088, n22089, n22090, n22091, n22092, n22093, n22094,
         n22095, n22096, n22097, n22098, n22099, n22100, n22101, n22102,
         n22103, n22104, n22105, n22106, n22107, n22108, n22109, n22110,
         n22111, n22112, n22113, n22114, n22115, n22116, n22117, n22118,
         n22119, n22120, n22121, n22122, n22123, n22124, n22125, n22126,
         n22127, n22128, n22129, n22130, n22131, n22132, n22133, n22134,
         n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142,
         n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150,
         n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158,
         n22159, n22160, n22161, n22162, n22163, n22164, n22165, n22166,
         n22167, n22168, n22169, n22170, n22171, n22172, n22173, n22174,
         n22175, n22176, n22177, n22178, n22179, n22180, n22181, n22182,
         n22183, n22184, n22185, n22186, n22187, n22188, n22189, n22190,
         n22191, n22192, n22193, n22194, n22195, n22196, n22197, n22198,
         n22199, n22200, n22201, n22202, n22203, n22204, n22205, n22206,
         n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214,
         n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222,
         n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230,
         n22231, n22232, n22233, n22234, n22235, n22236, n22237, n22238,
         n22239, n22240, n22241, n22242, n22243, n22244, n22245, n22246,
         n22247, n22248, n22249, n22250, n22251, n22252, n22253, n22254,
         n22255, n22256, n22257, n22258, n22259, n22260, n22261, n22262,
         n22263, n22264, n22265, n22266, n22267, n22268, n22269, n22270,
         n22271, n22272, n22273, n22274, n22275, n22276, n22277, n22278,
         n22279, n22280, n22281, n22282, n22283, n22284, n22285, n22286,
         n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294,
         n22295, n22296, n22297, n22298, n22299, n22300, n22301, n22302,
         n22303, n22304, n22305, n22306, n22307, n22308, n22309, n22310,
         n22311, n22312, n22313;

  AND2_X1 U11065 ( .A1(n12238), .A2(n16208), .ZN(n18526) );
  AOI21_X1 U11066 ( .B1(n12240), .B2(n12238), .A(n12239), .ZN(n18541) );
  NAND2_X1 U11067 ( .A1(n13757), .A2(n15956), .ZN(n15904) );
  AND4_X1 U11068 ( .A1(n11811), .A2(n11810), .A3(n11809), .A4(n11808), .ZN(
        n11820) );
  OR2_X1 U11069 ( .A1(n11782), .A2(n11781), .ZN(n19245) );
  INV_X1 U11070 ( .A(n11774), .ZN(n19621) );
  OAI21_X1 U11071 ( .B1(n12725), .B2(n12724), .A(n14793), .ZN(n14715) );
  INV_X1 U11072 ( .A(n17655), .ZN(n17502) );
  CLKBUF_X1 U11073 ( .A(n17361), .Z(n17535) );
  CLKBUF_X2 U11074 ( .A(n17356), .Z(n13463) );
  CLKBUF_X3 U11075 ( .A(n13456), .Z(n17689) );
  INV_X1 U11076 ( .A(n14019), .ZN(n20734) );
  CLKBUF_X1 U11077 ( .A(n11740), .Z(n13828) );
  BUF_X2 U11078 ( .A(n13934), .Z(n17554) );
  CLKBUF_X1 U11079 ( .A(n13468), .Z(n17721) );
  CLKBUF_X1 U11080 ( .A(n13440), .Z(n17656) );
  CLKBUF_X1 U11081 ( .A(n17510), .Z(n17714) );
  INV_X1 U11082 ( .A(n13479), .ZN(n17546) );
  NAND2_X1 U11083 ( .A1(n11698), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11740) );
  CLKBUF_X2 U11085 ( .A(n12737), .Z(n12679) );
  CLKBUF_X2 U11086 ( .A(n12653), .Z(n13285) );
  AND2_X1 U11087 ( .A1(n15280), .A2(n14198), .ZN(n14222) );
  MUX2_X1 U11088 ( .A(n12626), .B(n12629), .S(n14719), .Z(n12630) );
  AND2_X2 U11089 ( .A1(n11633), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11460) );
  BUF_X2 U11090 ( .A(n11651), .Z(n14370) );
  NAND2_X1 U11091 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n20777) );
  BUF_X1 U11092 ( .A(n11682), .Z(n12286) );
  INV_X1 U11093 ( .A(n11661), .ZN(n11685) );
  INV_X1 U11094 ( .A(n11643), .ZN(n11684) );
  AND4_X1 U11095 ( .A1(n11649), .A2(n11648), .A3(n11647), .A4(n11646), .ZN(
        n11650) );
  AND2_X1 U11096 ( .A1(n14900), .A2(n12520), .ZN(n12690) );
  AND2_X2 U11097 ( .A1(n12519), .A2(n14895), .ZN(n13260) );
  AND2_X1 U11098 ( .A1(n12519), .A2(n14749), .ZN(n12659) );
  INV_X1 U11100 ( .A(n14367), .ZN(n14200) );
  AND2_X2 U11101 ( .A1(n15322), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15319) );
  NOR2_X2 U11102 ( .A1(n11680), .A2(n19685), .ZN(n19604) );
  NAND2_X1 U11103 ( .A1(n12001), .A2(n11346), .ZN(n10958) );
  AND2_X1 U11104 ( .A1(n11882), .A2(n11881), .ZN(n10959) );
  AND2_X1 U11105 ( .A1(n11882), .A2(n11881), .ZN(n10960) );
  INV_X1 U11106 ( .A(n15175), .ZN(n10961) );
  OAI211_X1 U11107 ( .C1(n14452), .C2(n14561), .A(n11702), .B(n11701), .ZN(
        n10962) );
  OAI21_X2 U11108 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n16368), .A(
        n16394), .ZN(n12001) );
  NOR2_X1 U11109 ( .A1(n11696), .A2(n11695), .ZN(n12244) );
  OR2_X1 U11110 ( .A1(n11740), .A2(n11869), .ZN(n11702) );
  NAND2_X2 U11111 ( .A1(n15674), .A2(n15675), .ZN(n15664) );
  AND2_X1 U11113 ( .A1(n11245), .A2(n11680), .ZN(n11699) );
  NOR2_X1 U11114 ( .A1(n13325), .A2(n13324), .ZN(n13339) );
  INV_X2 U11115 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11454) );
  AND2_X2 U11116 ( .A1(n14895), .A2(n14730), .ZN(n12774) );
  AND2_X1 U11117 ( .A1(n14900), .A2(n14895), .ZN(n12653) );
  AOI21_X1 U11118 ( .B1(n11295), .B2(n11292), .A(n11034), .ZN(n11291) );
  AND2_X1 U11119 ( .A1(n14198), .A2(n11414), .ZN(n14225) );
  OR2_X1 U11120 ( .A1(n11941), .A2(n11942), .ZN(n11944) );
  NAND2_X1 U11121 ( .A1(n14388), .A2(n11313), .ZN(n12420) );
  INV_X1 U11122 ( .A(n15124), .ZN(n14719) );
  NAND3_X1 U11123 ( .A1(n12626), .A2(n13357), .A3(n12572), .ZN(n14846) );
  AND2_X1 U11124 ( .A1(n16174), .A2(n15124), .ZN(n14800) );
  INV_X1 U11125 ( .A(n19400), .ZN(n13849) );
  INV_X1 U11126 ( .A(n13395), .ZN(n17683) );
  INV_X1 U11127 ( .A(n20951), .ZN(n21171) );
  INV_X2 U11128 ( .A(n19975), .ZN(n20009) );
  NOR2_X2 U11129 ( .A1(n11959), .A2(n11958), .ZN(n11960) );
  NAND2_X1 U11130 ( .A1(n11684), .A2(n11661), .ZN(n12056) );
  XNOR2_X1 U11132 ( .A(n14449), .B(n14448), .ZN(n15604) );
  OAI221_X1 U11133 ( .B1(n14020), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n18134), .C2(n14019), .A(n14018), .ZN(n18117) );
  OR2_X1 U11134 ( .A1(n15664), .A2(n11265), .ZN(n10987) );
  AND2_X1 U11135 ( .A1(n14489), .A2(n11048), .ZN(n15500) );
  NOR2_X1 U11136 ( .A1(n20688), .A2(n20689), .ZN(n20687) );
  INV_X1 U11137 ( .A(n18055), .ZN(n18038) );
  INV_X1 U11140 ( .A(n10977), .ZN(n18136) );
  OR2_X2 U11141 ( .A1(n13402), .A2(n20777), .ZN(n11009) );
  NAND2_X2 U11142 ( .A1(n11414), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11419) );
  OR2_X1 U11143 ( .A1(n16264), .A2(n16265), .ZN(n10963) );
  NAND2_X2 U11144 ( .A1(n11175), .A2(n11168), .ZN(n11172) );
  NOR2_X2 U11145 ( .A1(n10963), .A2(n15514), .ZN(n15515) );
  OAI22_X2 U11146 ( .A1(n11823), .A2(n19557), .B1(n19245), .B2(n11806), .ZN(
        n11807) );
  NOR2_X1 U11147 ( .A1(n14850), .A2(n13663), .ZN(n12627) );
  OR2_X2 U11148 ( .A1(n12526), .A2(n12525), .ZN(n14850) );
  OR2_X2 U11149 ( .A1(n17756), .A2(n17785), .ZN(n17761) );
  AND2_X2 U11150 ( .A1(n11350), .A2(n11805), .ZN(n11859) );
  NOR4_X2 U11151 ( .A1(n16052), .A2(n16051), .A3(n16050), .A4(n16049), .ZN(
        n16053) );
  NAND2_X2 U11152 ( .A1(n11650), .A2(n11613), .ZN(n11659) );
  NAND2_X1 U11153 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20748), .ZN(
        n13402) );
  NOR2_X2 U11154 ( .A1(n18837), .A2(n20625), .ZN(n20746) );
  INV_X1 U11155 ( .A(n17698), .ZN(n10964) );
  INV_X4 U11156 ( .A(n11005), .ZN(n17698) );
  BUF_X4 U11157 ( .A(n17356), .Z(n17713) );
  NAND2_X1 U11158 ( .A1(n13713), .A2(n13734), .ZN(n10965) );
  NAND2_X1 U11159 ( .A1(n13713), .A2(n13734), .ZN(n13735) );
  INV_X1 U11160 ( .A(n13735), .ZN(n19975) );
  NOR2_X2 U11161 ( .A1(n13799), .A2(n11149), .ZN(n13803) );
  NOR2_X2 U11162 ( .A1(n13419), .A2(n13418), .ZN(n18878) );
  INV_X2 U11163 ( .A(n11691), .ZN(n11700) );
  NOR2_X2 U11164 ( .A1(n13474), .A2(n13473), .ZN(n18961) );
  NOR2_X2 U11165 ( .A1(n10987), .A2(n15623), .ZN(n15622) );
  NOR2_X1 U11166 ( .A1(n19990), .A2(n13743), .ZN(n16000) );
  NOR2_X1 U11167 ( .A1(n21496), .A2(n21494), .ZN(n21510) );
  NOR4_X2 U11168 ( .A1(n20622), .A2(n20621), .A3(n20719), .A4(n20620), .ZN(
        n20721) );
  INV_X1 U11169 ( .A(n15074), .ZN(n11771) );
  INV_X1 U11171 ( .A(n21051), .ZN(n21140) );
  NAND2_X1 U11172 ( .A1(n20760), .A2(n20831), .ZN(n20750) );
  INV_X1 U11173 ( .A(n11719), .ZN(n11741) );
  AND2_X1 U11174 ( .A1(n12263), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11719) );
  AND2_X1 U11175 ( .A1(n12059), .A2(n12246), .ZN(n12275) );
  INV_X4 U11176 ( .A(n12420), .ZN(n12280) );
  NOR2_X1 U11177 ( .A1(n18837), .A2(n13476), .ZN(n13968) );
  NAND2_X1 U11178 ( .A1(n12669), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13314) );
  NAND2_X1 U11180 ( .A1(n13606), .A2(n10979), .ZN(n14684) );
  NAND2_X1 U11181 ( .A1(n19057), .A2(n20661), .ZN(n13494) );
  INV_X1 U11182 ( .A(n13620), .ZN(n13617) );
  OR2_X1 U11183 ( .A1(n13543), .A2(n13534), .ZN(n13620) );
  INV_X2 U11187 ( .A(n12623), .ZN(n16174) );
  INV_X1 U11188 ( .A(n22148), .ZN(n12639) );
  NAND2_X1 U11189 ( .A1(n11015), .A2(n12535), .ZN(n13663) );
  AND2_X1 U11190 ( .A1(n11025), .A2(n12544), .ZN(n12621) );
  BUF_X2 U11191 ( .A(n12659), .Z(n13280) );
  CLKBUF_X2 U11192 ( .A(n11397), .Z(n14373) );
  CLKBUF_X2 U11193 ( .A(n12658), .Z(n13278) );
  CLKBUF_X2 U11194 ( .A(n13982), .Z(n17720) );
  CLKBUF_X2 U11195 ( .A(n13982), .Z(n17585) );
  INV_X4 U11196 ( .A(n11009), .ZN(n17719) );
  BUF_X4 U11198 ( .A(n13897), .Z(n10966) );
  CLKBUF_X2 U11199 ( .A(n19868), .Z(n21257) );
  AND2_X2 U11200 ( .A1(n11413), .A2(n11454), .ZN(n11651) );
  NOR2_X1 U11201 ( .A1(n16543), .A2(n11075), .ZN(n18576) );
  NOR2_X1 U11202 ( .A1(n16554), .A2(n16553), .ZN(n16552) );
  CLKBUF_X1 U11203 ( .A(n16514), .Z(n10972) );
  AND2_X1 U11204 ( .A1(n11082), .A2(n17247), .ZN(n16554) );
  NAND2_X1 U11205 ( .A1(n11209), .A2(n16798), .ZN(n16567) );
  INV_X1 U11206 ( .A(n16796), .ZN(n11209) );
  OR2_X1 U11207 ( .A1(n15586), .A2(n19957), .ZN(n11377) );
  XNOR2_X1 U11208 ( .A(n15622), .B(n13304), .ZN(n13660) );
  AND2_X1 U11209 ( .A1(n11101), .A2(n11100), .ZN(n16591) );
  AND2_X1 U11210 ( .A1(n14460), .A2(n13843), .ZN(n14430) );
  NOR2_X1 U11211 ( .A1(n16290), .A2(n13835), .ZN(n13839) );
  NOR2_X1 U11212 ( .A1(n16250), .A2(n16244), .ZN(n16237) );
  NAND2_X1 U11213 ( .A1(n15361), .A2(n12090), .ZN(n12098) );
  NAND2_X1 U11214 ( .A1(n11905), .A2(n18290), .ZN(n11906) );
  NAND2_X1 U11215 ( .A1(n11853), .A2(n11852), .ZN(n11334) );
  AND2_X1 U11216 ( .A1(n11251), .A2(n11255), .ZN(n15431) );
  NOR2_X1 U11217 ( .A1(n15086), .A2(n11252), .ZN(n11251) );
  OR2_X1 U11218 ( .A1(n15990), .A2(n15989), .ZN(n15999) );
  OR2_X1 U11219 ( .A1(n16014), .A2(n16013), .ZN(n19990) );
  AND2_X1 U11220 ( .A1(n11901), .A2(n11900), .ZN(n12097) );
  AND2_X1 U11221 ( .A1(n11851), .A2(n11850), .ZN(n11854) );
  INV_X1 U11222 ( .A(n18129), .ZN(n18122) );
  AND2_X1 U11223 ( .A1(n15689), .A2(n11226), .ZN(n15640) );
  NAND2_X1 U11224 ( .A1(n17978), .A2(n17977), .ZN(n18129) );
  NAND2_X1 U11225 ( .A1(n14761), .A2(n14088), .ZN(n14916) );
  AND2_X1 U11226 ( .A1(n11784), .A2(n11785), .ZN(n11351) );
  OAI22_X1 U11227 ( .A1(n19530), .A2(n11842), .B1(n11840), .B2(n11815), .ZN(
        n11816) );
  OR2_X1 U11228 ( .A1(n14929), .A2(n14964), .ZN(n14991) );
  CLKBUF_X1 U11229 ( .A(n11826), .Z(n19215) );
  NAND2_X1 U11230 ( .A1(n12795), .A2(n11259), .ZN(n13713) );
  OAI21_X1 U11231 ( .B1(n21769), .B2(n12978), .A(n12855), .ZN(n14976) );
  AOI21_X1 U11232 ( .B1(n11830), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A(
        n19621), .ZN(n11778) );
  INV_X1 U11233 ( .A(n12872), .ZN(n12795) );
  NAND2_X1 U11234 ( .A1(n11277), .A2(n16154), .ZN(n12857) );
  AND2_X1 U11235 ( .A1(n12844), .A2(n12843), .ZN(n14835) );
  NAND2_X1 U11236 ( .A1(n11768), .A2(n18258), .ZN(n11782) );
  NAND2_X1 U11237 ( .A1(n10989), .A2(n11755), .ZN(n19268) );
  AND2_X2 U11238 ( .A1(n14055), .A2(n11762), .ZN(n11834) );
  NAND2_X1 U11239 ( .A1(n11277), .A2(n11276), .ZN(n12872) );
  NOR2_X1 U11240 ( .A1(n10980), .A2(n21836), .ZN(n21782) );
  AOI22_X1 U11241 ( .A1(n21185), .A2(n21183), .B1(n21189), .B2(n17748), .ZN(
        n21196) );
  AND2_X1 U11242 ( .A1(n14921), .A2(n14920), .ZN(n14918) );
  INV_X1 U11243 ( .A(n11767), .ZN(n11776) );
  NOR2_X1 U11244 ( .A1(n11944), .A2(n11176), .ZN(n11584) );
  AND2_X1 U11245 ( .A1(n16154), .A2(n12856), .ZN(n11276) );
  CLKBUF_X1 U11246 ( .A(n15598), .Z(n15880) );
  CLKBUF_X1 U11247 ( .A(n13371), .Z(n15878) );
  AND2_X1 U11248 ( .A1(n12816), .A2(n12814), .ZN(n12749) );
  NAND2_X1 U11249 ( .A1(n12769), .A2(n12768), .ZN(n16154) );
  NAND2_X1 U11250 ( .A1(n20559), .A2(n21051), .ZN(n21190) );
  NOR2_X1 U11251 ( .A1(n21825), .A2(n21675), .ZN(n21935) );
  NAND2_X1 U11252 ( .A1(n11751), .A2(n11754), .ZN(n15074) );
  NAND2_X2 U11253 ( .A1(n15886), .A2(n14949), .ZN(n15890) );
  XNOR2_X1 U11254 ( .A(n14793), .B(n15115), .ZN(n21771) );
  NOR2_X2 U11255 ( .A1(n19351), .A2(n19683), .ZN(n19352) );
  NOR2_X2 U11256 ( .A1(n19183), .A2(n19683), .ZN(n15206) );
  NOR2_X2 U11257 ( .A1(n19398), .A2(n19683), .ZN(n19399) );
  NAND2_X1 U11258 ( .A1(n12725), .A2(n12724), .ZN(n14793) );
  XNOR2_X1 U11259 ( .A(n12126), .B(n12127), .ZN(n12125) );
  NOR2_X1 U11260 ( .A1(n15049), .A2(n15375), .ZN(n15484) );
  NAND2_X1 U11261 ( .A1(n11714), .A2(n11713), .ZN(n11160) );
  INV_X2 U11262 ( .A(n20332), .ZN(n10967) );
  OAI211_X1 U11263 ( .C1(n14452), .C2(n15292), .A(n11743), .B(n11742), .ZN(
        n12126) );
  OR2_X1 U11264 ( .A1(n13828), .A2(n15289), .ZN(n11743) );
  XNOR2_X1 U11265 ( .A(n13998), .B(n11300), .ZN(n18080) );
  NAND2_X1 U11266 ( .A1(n12302), .A2(n12301), .ZN(n11326) );
  BUF_X2 U11267 ( .A(n13828), .Z(n10978) );
  INV_X2 U11268 ( .A(n15031), .ZN(n18562) );
  CLKBUF_X1 U11269 ( .A(n15031), .Z(n18361) );
  NAND2_X1 U11270 ( .A1(n12634), .A2(n12707), .ZN(n12829) );
  NOR2_X1 U11271 ( .A1(n14808), .A2(n12297), .ZN(n12304) );
  OAI211_X1 U11272 ( .C1(n11740), .C2(n11712), .A(n11711), .B(n11710), .ZN(
        n11715) );
  INV_X4 U11273 ( .A(n11741), .ZN(n14450) );
  NOR2_X1 U11274 ( .A1(n11867), .A2(n11868), .ZN(n11862) );
  NAND2_X1 U11275 ( .A1(n11709), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n11711) );
  AND2_X1 U11276 ( .A1(n14650), .A2(n14651), .ZN(n14653) );
  NOR2_X1 U11277 ( .A1(n12276), .A2(n11675), .ZN(n11727) );
  OAI21_X1 U11278 ( .B1(n13889), .B2(n11094), .A(n11091), .ZN(n13493) );
  NAND2_X1 U11279 ( .A1(n11674), .A2(n11673), .ZN(n12276) );
  NOR2_X2 U11280 ( .A1(n13972), .A2(n20593), .ZN(n18010) );
  AOI21_X1 U11281 ( .B1(n15577), .B2(n14705), .A(n12638), .ZN(n12631) );
  AND3_X1 U11282 ( .A1(n11700), .A2(n11699), .A3(n12253), .ZN(n12263) );
  NAND2_X1 U11283 ( .A1(n11670), .A2(n10991), .ZN(n12052) );
  AND2_X1 U11284 ( .A1(n12248), .A2(n12250), .ZN(n11732) );
  AND2_X1 U11285 ( .A1(n12286), .A2(n12056), .ZN(n12248) );
  INV_X2 U11286 ( .A(n12479), .ZN(n12488) );
  OR2_X1 U11287 ( .A1(n12622), .A2(n14703), .ZN(n14705) );
  AND2_X1 U11288 ( .A1(n10991), .A2(n11114), .ZN(n12059) );
  NAND2_X1 U11289 ( .A1(n12056), .A2(n11686), .ZN(n11689) );
  NAND2_X1 U11290 ( .A1(n11693), .A2(n11644), .ZN(n11663) );
  AND2_X1 U11291 ( .A1(n12246), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n18240) );
  OR2_X1 U11292 ( .A1(n13620), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n11376) );
  OR2_X1 U11293 ( .A1(n14725), .A2(n14844), .ZN(n14872) );
  BUF_X2 U11294 ( .A(n11685), .Z(n19400) );
  OR2_X2 U11295 ( .A1(n11572), .A2(n11571), .ZN(n14446) );
  INV_X1 U11296 ( .A(n11686), .ZN(n11245) );
  OR2_X1 U11297 ( .A1(n14717), .A2(n13543), .ZN(n14866) );
  OR2_X1 U11298 ( .A1(n12618), .A2(n12619), .ZN(n15577) );
  NAND2_X1 U11299 ( .A1(n15162), .A2(n15124), .ZN(n13606) );
  NOR2_X1 U11300 ( .A1(n12286), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12287) );
  NAND2_X1 U11301 ( .A1(n11628), .A2(n11627), .ZN(n11668) );
  NAND2_X1 U11302 ( .A1(n11247), .A2(n11246), .ZN(n11686) );
  INV_X1 U11303 ( .A(n11662), .ZN(n12057) );
  OR3_X2 U11304 ( .A1(n11190), .A2(n13991), .A3(n11191), .ZN(n20739) );
  NOR2_X1 U11305 ( .A1(n14871), .A2(n15596), .ZN(n13357) );
  INV_X2 U11306 ( .A(U212), .ZN(n10968) );
  NAND2_X1 U11307 ( .A1(n15596), .A2(n12621), .ZN(n14717) );
  NAND2_X2 U11308 ( .A1(U214), .A2(n20027), .ZN(n20088) );
  OR2_X1 U11309 ( .A1(n12702), .A2(n12701), .ZN(n13675) );
  OR2_X1 U11310 ( .A1(n12685), .A2(n12684), .ZN(n13737) );
  OR2_X2 U11311 ( .A1(n12554), .A2(n12553), .ZN(n15596) );
  NAND2_X1 U11312 ( .A1(n20021), .A2(n15121), .ZN(n22152) );
  AND2_X1 U11313 ( .A1(n11653), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11655) );
  AND4_X1 U11314 ( .A1(n12584), .A2(n12583), .A3(n12582), .A4(n12581), .ZN(
        n12590) );
  AND4_X1 U11315 ( .A1(n12596), .A2(n12595), .A3(n12594), .A4(n12593), .ZN(
        n12612) );
  AND4_X1 U11316 ( .A1(n12576), .A2(n12575), .A3(n12574), .A4(n12573), .ZN(
        n12592) );
  AND4_X1 U11317 ( .A1(n12608), .A2(n12607), .A3(n12606), .A4(n12605), .ZN(
        n12609) );
  AND4_X1 U11318 ( .A1(n12558), .A2(n12557), .A3(n12556), .A4(n12555), .ZN(
        n12563) );
  BUF_X2 U11319 ( .A(n11788), .Z(n14230) );
  AND4_X1 U11320 ( .A1(n12539), .A2(n12538), .A3(n12537), .A4(n12536), .ZN(
        n11025) );
  AND4_X1 U11321 ( .A1(n12543), .A2(n12542), .A3(n12541), .A4(n12540), .ZN(
        n12544) );
  AND4_X1 U11322 ( .A1(n12600), .A2(n12599), .A3(n12598), .A4(n12597), .ZN(
        n12611) );
  AND4_X1 U11323 ( .A1(n12534), .A2(n12533), .A3(n12532), .A4(n12531), .ZN(
        n12535) );
  AND4_X1 U11324 ( .A1(n12588), .A2(n12587), .A3(n12586), .A4(n12585), .ZN(
        n12589) );
  AND4_X1 U11325 ( .A1(n12604), .A2(n12603), .A3(n12602), .A4(n12601), .ZN(
        n12610) );
  AND4_X1 U11326 ( .A1(n12580), .A2(n12579), .A3(n12578), .A4(n12577), .ZN(
        n12591) );
  INV_X2 U11327 ( .A(n19050), .ZN(U215) );
  INV_X2 U11328 ( .A(n13395), .ZN(n20181) );
  AND2_X2 U11329 ( .A1(n11652), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14215) );
  NAND2_X2 U11330 ( .A1(n17340), .A2(n21640), .ZN(n17339) );
  NAND2_X2 U11331 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n17340), .ZN(n17337) );
  CLKBUF_X2 U11332 ( .A(n13986), .Z(n17590) );
  BUF_X2 U11333 ( .A(n11397), .Z(n11633) );
  INV_X2 U11334 ( .A(n19800), .ZN(n19853) );
  BUF_X4 U11335 ( .A(n11396), .Z(n10974) );
  BUF_X2 U11336 ( .A(n11396), .Z(n10975) );
  BUF_X2 U11337 ( .A(n12690), .Z(n12673) );
  OR2_X1 U11338 ( .A1(n20777), .A2(n13400), .ZN(n11005) );
  NOR2_X1 U11339 ( .A1(n20775), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n20769) );
  NAND2_X1 U11340 ( .A1(n20748), .A2(n20759), .ZN(n20146) );
  AND2_X2 U11341 ( .A1(n12512), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12519) );
  INV_X2 U11342 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n20748) );
  NAND2_X1 U11343 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16881) );
  AND2_X1 U11344 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11413) );
  NAND2_X1 U11345 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n20775) );
  AND2_X2 U11346 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n14895) );
  NOR2_X2 U11347 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12520) );
  NAND2_X1 U11348 ( .A1(n11907), .A2(n11079), .ZN(n11078) );
  NAND2_X1 U11349 ( .A1(n11752), .A2(n11349), .ZN(n11159) );
  NOR2_X1 U11350 ( .A1(n14443), .A2(n14441), .ZN(n14416) );
  NAND2_X1 U11351 ( .A1(n14443), .A2(n14442), .ZN(n11120) );
  XNOR2_X1 U11352 ( .A(n11906), .B(n16834), .ZN(n16860) );
  XNOR2_X2 U11353 ( .A(n11745), .B(n11744), .ZN(n14066) );
  OAI21_X2 U11354 ( .B1(n11035), .B2(n12632), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12648) );
  NAND3_X2 U11355 ( .A1(n12617), .A2(n13349), .A3(n14872), .ZN(n11035) );
  NAND2_X1 U11356 ( .A1(n11159), .A2(n11160), .ZN(n10970) );
  OAI21_X1 U11357 ( .B1(n16567), .B2(n16446), .A(n16445), .ZN(n10973) );
  NAND2_X2 U11358 ( .A1(n11616), .A2(n11615), .ZN(n11643) );
  OAI21_X1 U11359 ( .B1(n16567), .B2(n16446), .A(n16445), .ZN(n16516) );
  NAND2_X1 U11361 ( .A1(n11906), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11907) );
  NAND2_X1 U11362 ( .A1(n11159), .A2(n11160), .ZN(n11745) );
  OAI21_X1 U11363 ( .B1(n16567), .B2(n16523), .A(n16522), .ZN(n11082) );
  NAND2_X2 U11364 ( .A1(n13523), .A2(n16174), .ZN(n13349) );
  OAI21_X2 U11365 ( .B1(n11860), .B2(n11859), .A(n12086), .ZN(n15290) );
  NAND2_X1 U11366 ( .A1(n11162), .A2(n11161), .ZN(n11339) );
  XNOR2_X1 U11367 ( .A(n12100), .B(n12097), .ZN(n12092) );
  NOR2_X2 U11368 ( .A1(n16229), .A2(n16224), .ZN(n16216) );
  OAI211_X1 U11369 ( .C1(n14452), .C2(n14561), .A(n11702), .B(n11701), .ZN(
        n11703) );
  NAND2_X1 U11370 ( .A1(n15124), .A2(n12623), .ZN(n13534) );
  AND4_X2 U11371 ( .A1(n12637), .A2(n11280), .A3(n11279), .A4(n11278), .ZN(
        n12635) );
  NAND2_X2 U11372 ( .A1(n11336), .A2(n11017), .ZN(n11842) );
  NOR2_X2 U11373 ( .A1(n15613), .A2(n22310), .ZN(n14804) );
  NAND2_X2 U11374 ( .A1(n13347), .A2(n13346), .ZN(n15613) );
  AND2_X2 U11375 ( .A1(n12635), .A2(n12616), .ZN(n13523) );
  AOI21_X1 U11376 ( .B1(n12129), .B2(n11080), .A(n12128), .ZN(n14921) );
  NAND2_X2 U11377 ( .A1(n12717), .A2(n21783), .ZN(n14906) );
  XNOR2_X2 U11378 ( .A(n13691), .B(n14959), .ZN(n14956) );
  INV_X2 U11379 ( .A(n13547), .ZN(n10979) );
  XNOR2_X2 U11380 ( .A(n13684), .B(n13683), .ZN(n14937) );
  NAND2_X1 U11381 ( .A1(n10989), .A2(n11017), .ZN(n19310) );
  AND2_X2 U11382 ( .A1(n11767), .A2(n18258), .ZN(n10989) );
  AOI211_X2 U11383 ( .C1(n18605), .C2(n17258), .A(n16485), .B(n16484), .ZN(
        n16486) );
  OAI21_X4 U11384 ( .B1(n13731), .B2(n11293), .A(n11291), .ZN(n19974) );
  NAND2_X2 U11385 ( .A1(n15402), .A2(n15401), .ZN(n13731) );
  AND2_X1 U11386 ( .A1(n14895), .A2(n14730), .ZN(n10981) );
  AND2_X2 U11387 ( .A1(n14895), .A2(n14730), .ZN(n10982) );
  AND2_X1 U11388 ( .A1(n12518), .A2(n12519), .ZN(n10983) );
  AND2_X2 U11389 ( .A1(n12518), .A2(n12519), .ZN(n10984) );
  NAND2_X1 U11391 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18060), .ZN(
        n14036) );
  INV_X1 U11392 ( .A(n14409), .ZN(n11343) );
  XNOR2_X1 U11393 ( .A(n15181), .B(n14081), .ZN(n14764) );
  AOI21_X1 U11394 ( .B1(n15074), .B2(n14062), .A(n14077), .ZN(n14765) );
  INV_X1 U11395 ( .A(n12810), .ZN(n11258) );
  NAND2_X1 U11396 ( .A1(n12618), .A2(n13663), .ZN(n12637) );
  NAND2_X1 U11397 ( .A1(n12631), .A2(n12630), .ZN(n12632) );
  NAND2_X1 U11398 ( .A1(n21771), .A2(n16946), .ZN(n12769) );
  INV_X1 U11399 ( .A(n13314), .ZN(n13341) );
  NAND2_X1 U11400 ( .A1(n14871), .A2(n15124), .ZN(n12726) );
  AND2_X1 U11401 ( .A1(n11411), .A2(n11454), .ZN(n11397) );
  AND2_X1 U11402 ( .A1(n11121), .A2(n15478), .ZN(n12099) );
  INV_X1 U11403 ( .A(n12097), .ZN(n12101) );
  AOI22_X1 U11404 ( .A1(n11813), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11812), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11819) );
  AOI21_X1 U11405 ( .B1(n20734), .B2(n20739), .A(n20616), .ZN(n14015) );
  NAND2_X1 U11406 ( .A1(n13880), .A2(n18796), .ZN(n11092) );
  INV_X1 U11407 ( .A(n15367), .ZN(n11253) );
  INV_X1 U11408 ( .A(n13302), .ZN(n13522) );
  INV_X1 U11409 ( .A(n13272), .ZN(n13302) );
  INV_X1 U11410 ( .A(n13232), .ZN(n13296) );
  NOR2_X1 U11411 ( .A1(n11227), .A2(n15638), .ZN(n11226) );
  INV_X1 U11412 ( .A(n11228), .ZN(n11227) );
  NAND2_X1 U11413 ( .A1(n12726), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13345) );
  OR2_X1 U11414 ( .A1(n15200), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n11365) );
  NOR2_X1 U11415 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14198) );
  NOR2_X1 U11416 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n12050), .ZN(
        n12385) );
  AND2_X1 U11417 ( .A1(n18535), .A2(n14446), .ZN(n11587) );
  INV_X1 U11418 ( .A(n18372), .ZN(n11316) );
  NAND2_X1 U11419 ( .A1(n11220), .A2(n15222), .ZN(n11219) );
  INV_X1 U11420 ( .A(n11221), .ZN(n11220) );
  CLKBUF_X1 U11421 ( .A(n12092), .Z(n12093) );
  OAI21_X1 U11422 ( .B1(n21193), .B2(n13965), .A(n21222), .ZN(n16900) );
  NOR2_X1 U11423 ( .A1(n13400), .A2(n13393), .ZN(n13986) );
  NOR2_X1 U11424 ( .A1(n13402), .A2(n13403), .ZN(n13440) );
  OR2_X1 U11425 ( .A1(n20597), .A2(n13973), .ZN(n13972) );
  NAND2_X1 U11426 ( .A1(n18091), .A2(n13996), .ZN(n13998) );
  AND2_X1 U11427 ( .A1(n12166), .A2(n12165), .ZN(n15269) );
  NAND2_X1 U11428 ( .A1(n13839), .A2(n13840), .ZN(n14460) );
  NAND2_X1 U11429 ( .A1(n12001), .A2(n11346), .ZN(n11344) );
  NOR2_X1 U11430 ( .A1(n11347), .A2(n11019), .ZN(n11346) );
  INV_X1 U11431 ( .A(n12000), .ZN(n11347) );
  AND2_X1 U11432 ( .A1(n16545), .A2(n16544), .ZN(n11075) );
  AND2_X1 U11433 ( .A1(n12077), .A2(n18683), .ZN(n12279) );
  AOI21_X1 U11434 ( .B1(n14765), .B2(n14764), .A(n14083), .ZN(n14768) );
  OR2_X1 U11435 ( .A1(n19447), .A2(n18260), .ZN(n19195) );
  AOI21_X1 U11436 ( .B1(n20562), .B2(n20561), .A(n20560), .ZN(n20565) );
  AOI21_X1 U11437 ( .B1(n14037), .B2(n14036), .A(n14035), .ZN(n18051) );
  AND2_X1 U11438 ( .A1(n18641), .A2(n14498), .ZN(n18248) );
  AND2_X1 U11439 ( .A1(n18645), .A2(n18683), .ZN(n18686) );
  AND2_X1 U11440 ( .A1(n16216), .A2(n11234), .ZN(n14456) );
  AND2_X1 U11441 ( .A1(n11017), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11335) );
  AND2_X1 U11442 ( .A1(n12620), .A2(n14948), .ZN(n13650) );
  INV_X1 U11443 ( .A(n13345), .ZN(n13333) );
  NOR2_X1 U11444 ( .A1(n12877), .A2(n11260), .ZN(n11259) );
  INV_X1 U11445 ( .A(n12871), .ZN(n11260) );
  BUF_X1 U11446 ( .A(n13260), .Z(n13279) );
  OR2_X1 U11447 ( .A1(n13315), .A2(n15093), .ZN(n13334) );
  NAND2_X1 U11448 ( .A1(n11666), .A2(n19686), .ZN(n11733) );
  NAND2_X1 U11449 ( .A1(n11428), .A2(n11427), .ZN(n11438) );
  NAND2_X1 U11450 ( .A1(n11603), .A2(n11602), .ZN(n11662) );
  INV_X1 U11451 ( .A(n11685), .ZN(n11081) );
  INV_X1 U11452 ( .A(n20776), .ZN(n13401) );
  NAND2_X1 U11453 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n20764), .ZN(
        n13393) );
  NAND2_X1 U11454 ( .A1(n14717), .A2(n14850), .ZN(n11279) );
  NAND2_X1 U11455 ( .A1(n12619), .A2(n14844), .ZN(n11280) );
  NAND2_X1 U11456 ( .A1(n12615), .A2(n15151), .ZN(n11278) );
  NAND2_X1 U11457 ( .A1(n15649), .A2(n11268), .ZN(n11267) );
  INV_X1 U11458 ( .A(n15665), .ZN(n11268) );
  AND2_X1 U11459 ( .A1(n11271), .A2(n11270), .ZN(n11269) );
  INV_X1 U11460 ( .A(n15691), .ZN(n11270) );
  NOR2_X1 U11461 ( .A1(n15710), .A2(n11274), .ZN(n11273) );
  INV_X1 U11462 ( .A(n15726), .ZN(n11274) );
  NAND2_X1 U11463 ( .A1(n16159), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13299) );
  INV_X1 U11464 ( .A(n15261), .ZN(n11255) );
  INV_X1 U11465 ( .A(n11298), .ZN(n11292) );
  INV_X1 U11466 ( .A(n13534), .ZN(n14687) );
  INV_X1 U11467 ( .A(n12726), .ZN(n12669) );
  XNOR2_X1 U11468 ( .A(n13666), .B(n12747), .ZN(n12826) );
  AOI21_X1 U11469 ( .B1(n12836), .B2(n12835), .A(n12713), .ZN(n12825) );
  NAND2_X1 U11470 ( .A1(n12723), .A2(n12722), .ZN(n12724) );
  INV_X1 U11471 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21794) );
  AOI21_X1 U11472 ( .B1(n21253), .B2(n21583), .A(n21597), .ZN(n15122) );
  NAND2_X1 U11473 ( .A1(n11457), .A2(n11456), .ZN(n12035) );
  NAND2_X1 U11474 ( .A1(n11804), .A2(n11700), .ZN(n11457) );
  NOR2_X1 U11475 ( .A1(n11182), .A2(n11982), .ZN(n11180) );
  NAND2_X1 U11476 ( .A1(n11584), .A2(n11378), .ZN(n11959) );
  OR3_X1 U11477 ( .A1(n11177), .A2(n11938), .A3(n11059), .ZN(n11176) );
  INV_X1 U11478 ( .A(n11374), .ZN(n11177) );
  INV_X1 U11479 ( .A(n11928), .ZN(n11578) );
  NOR2_X1 U11480 ( .A1(n11185), .A2(n11060), .ZN(n11184) );
  INV_X1 U11481 ( .A(n11186), .ZN(n11185) );
  INV_X1 U11482 ( .A(n14320), .ZN(n14298) );
  OR2_X2 U11483 ( .A1(n16881), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14367) );
  NAND2_X1 U11484 ( .A1(n14648), .A2(n11774), .ZN(n14320) );
  AND2_X1 U11485 ( .A1(n11330), .A2(n11329), .ZN(n11328) );
  INV_X1 U11486 ( .A(n16670), .ZN(n11329) );
  AND2_X1 U11487 ( .A1(n16692), .A2(n15551), .ZN(n11330) );
  INV_X1 U11488 ( .A(n16840), .ZN(n11322) );
  NOR2_X1 U11489 ( .A1(n11552), .A2(n11551), .ZN(n12323) );
  AND2_X1 U11490 ( .A1(n11690), .A2(n11699), .ZN(n12254) );
  INV_X1 U11491 ( .A(n16257), .ZN(n11225) );
  INV_X1 U11492 ( .A(n15498), .ZN(n11212) );
  OR2_X1 U11493 ( .A1(n11152), .A2(n11151), .ZN(n11150) );
  NAND2_X1 U11494 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11152) );
  NOR2_X1 U11495 ( .A1(n17223), .A2(n16593), .ZN(n11144) );
  NAND2_X1 U11496 ( .A1(n18523), .A2(n14446), .ZN(n11999) );
  NAND2_X1 U11497 ( .A1(n11174), .A2(n16366), .ZN(n11173) );
  INV_X1 U11498 ( .A(n16401), .ZN(n11174) );
  OR2_X1 U11499 ( .A1(n16419), .A2(n11163), .ZN(n11165) );
  NAND2_X1 U11500 ( .A1(n11170), .A2(n11164), .ZN(n11163) );
  INV_X1 U11501 ( .A(n16421), .ZN(n11164) );
  INV_X1 U11502 ( .A(n18467), .ZN(n11986) );
  NAND2_X1 U11503 ( .A1(n16430), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11978) );
  NAND2_X1 U11504 ( .A1(n16439), .A2(n11932), .ZN(n11162) );
  AND2_X1 U11505 ( .A1(n11957), .A2(n11340), .ZN(n11161) );
  OR2_X1 U11506 ( .A1(n16454), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11340) );
  NAND2_X1 U11507 ( .A1(n11222), .A2(n15060), .ZN(n11221) );
  INV_X1 U11508 ( .A(n14992), .ZN(n11222) );
  OR2_X1 U11509 ( .A1(n12100), .A2(n12101), .ZN(n12104) );
  NAND2_X1 U11510 ( .A1(n12098), .A2(n11104), .ZN(n11103) );
  NAND2_X1 U11511 ( .A1(n12091), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11104) );
  INV_X1 U11512 ( .A(n12099), .ZN(n11105) );
  NAND2_X1 U11513 ( .A1(n12096), .A2(n11108), .ZN(n16862) );
  OAI21_X1 U11514 ( .B1(n12099), .B2(n12098), .A(n12095), .ZN(n11108) );
  NAND2_X1 U11515 ( .A1(n11107), .A2(n11106), .ZN(n16861) );
  NAND2_X1 U11516 ( .A1(n12095), .A2(n15478), .ZN(n11106) );
  OAI21_X1 U11517 ( .B1(n15290), .B2(n15291), .A(n12085), .ZN(n12088) );
  NAND2_X1 U11518 ( .A1(n11748), .A2(n11747), .ZN(n11752) );
  OAI211_X1 U11519 ( .C1(n11741), .C2(n14696), .A(n18656), .B(n11726), .ZN(
        n11730) );
  AND2_X1 U11520 ( .A1(n11671), .A2(n11680), .ZN(n11672) );
  AND2_X1 U11521 ( .A1(n14298), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14072) );
  AOI21_X1 U11522 ( .B1(n15047), .B2(n14062), .A(n14061), .ZN(n14064) );
  OR2_X1 U11523 ( .A1(n14320), .A2(n19557), .ZN(n14063) );
  OR2_X1 U11524 ( .A1(n14064), .A2(n14063), .ZN(n14087) );
  NAND2_X1 U11525 ( .A1(n11638), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11247) );
  NAND2_X1 U11526 ( .A1(n11639), .A2(n11613), .ZN(n11246) );
  OR2_X1 U11527 ( .A1(n12024), .A2(n12023), .ZN(n12026) );
  NOR2_X1 U11528 ( .A1(n13401), .A2(n20146), .ZN(n13392) );
  NOR2_X1 U11529 ( .A1(n13379), .A2(n11133), .ZN(n11132) );
  NOR2_X1 U11530 ( .A1(n11135), .A2(n13378), .ZN(n11134) );
  INV_X1 U11531 ( .A(n11137), .ZN(n11135) );
  OR2_X1 U11532 ( .A1(n18044), .A2(n18010), .ZN(n17775) );
  NAND2_X1 U11533 ( .A1(n18072), .A2(n14001), .ZN(n17773) );
  NOR2_X1 U11534 ( .A1(n18082), .A2(n14027), .ZN(n14029) );
  AND2_X1 U11535 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14026), .ZN(
        n14027) );
  NAND2_X1 U11536 ( .A1(n11200), .A2(n11033), .ZN(n11199) );
  NOR2_X1 U11537 ( .A1(n20748), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13868) );
  AOI21_X1 U11538 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n21214), .A(
        n13507), .ZN(n13874) );
  NAND2_X1 U11539 ( .A1(n20763), .A2(n13882), .ZN(n11094) );
  INV_X1 U11540 ( .A(n13968), .ZN(n11093) );
  INV_X1 U11541 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21204) );
  INV_X1 U11542 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n21214) );
  INV_X1 U11543 ( .A(n21552), .ZN(n21495) );
  INV_X1 U11544 ( .A(n15095), .ZN(n15092) );
  NAND2_X1 U11545 ( .A1(n14685), .A2(n14687), .ZN(n11248) );
  NAND2_X1 U11546 ( .A1(n13128), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13158) );
  AND2_X1 U11547 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n13094), .ZN(
        n13095) );
  AND3_X1 U11548 ( .A1(n12901), .A2(n12900), .A3(n12899), .ZN(n15367) );
  AOI21_X1 U11549 ( .B1(n13694), .B2(n14820), .A(n12868), .ZN(n14998) );
  NAND2_X1 U11550 ( .A1(n13761), .A2(n13760), .ZN(n13771) );
  INV_X1 U11551 ( .A(n13777), .ZN(n13761) );
  NAND2_X1 U11552 ( .A1(n15689), .A2(n11063), .ZN(n15629) );
  INV_X1 U11553 ( .A(n15906), .ZN(n11311) );
  NOR2_X1 U11554 ( .A1(n13740), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11296) );
  NAND2_X1 U11555 ( .A1(n13731), .A2(n11298), .ZN(n11297) );
  AND2_X1 U11556 ( .A1(n21769), .A2(n14911), .ZN(n21809) );
  AND2_X1 U11557 ( .A1(n21819), .A2(n10980), .ZN(n21851) );
  INV_X1 U11558 ( .A(n22145), .ZN(n21825) );
  NOR2_X1 U11559 ( .A1(n21863), .A2(n21825), .ZN(n21942) );
  AND2_X1 U11560 ( .A1(n10980), .A2(n21836), .ZN(n21791) );
  INV_X1 U11561 ( .A(n21921), .ZN(n21914) );
  AOI21_X1 U11562 ( .B1(n21915), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n21825), 
        .ZN(n21923) );
  AND2_X1 U11563 ( .A1(n10980), .A2(n21850), .ZN(n21808) );
  OR2_X1 U11564 ( .A1(n13355), .A2(n13345), .ZN(n13346) );
  OAI21_X1 U11565 ( .B1(n13355), .B2(n13344), .A(n13343), .ZN(n13347) );
  OAI21_X1 U11566 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n12860), .A(n13342), 
        .ZN(n13343) );
  NAND2_X1 U11567 ( .A1(n11995), .A2(n11993), .ZN(n11990) );
  AND2_X1 U11568 ( .A1(n11960), .A2(n11178), .ZN(n11995) );
  NOR2_X1 U11569 ( .A1(n11179), .A2(n11064), .ZN(n11178) );
  INV_X1 U11570 ( .A(n11180), .ZN(n11179) );
  CLKBUF_X1 U11571 ( .A(n12054), .Z(n12055) );
  NAND2_X1 U11572 ( .A1(n11218), .A2(n11217), .ZN(n11216) );
  INV_X1 U11573 ( .A(n15269), .ZN(n11217) );
  INV_X1 U11574 ( .A(n11219), .ZN(n11218) );
  AND2_X1 U11575 ( .A1(n14298), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14915) );
  INV_X1 U11576 ( .A(n11238), .ZN(n11236) );
  NAND2_X1 U11577 ( .A1(n16377), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16378) );
  XNOR2_X1 U11578 ( .A(n16453), .B(n11210), .ZN(n16471) );
  INV_X1 U11579 ( .A(n16454), .ZN(n11210) );
  AOI21_X1 U11580 ( .B1(n16591), .B2(n12109), .A(n11366), .ZN(n16819) );
  AND2_X1 U11581 ( .A1(n16592), .A2(n16820), .ZN(n12109) );
  OR2_X1 U11582 ( .A1(n18304), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16586) );
  AND2_X1 U11583 ( .A1(n12141), .A2(n12140), .ZN(n14931) );
  NOR2_X1 U11584 ( .A1(n16764), .A2(n12265), .ZN(n16833) );
  INV_X1 U11585 ( .A(n16880), .ZN(n11359) );
  AND2_X1 U11586 ( .A1(n15041), .A2(n11771), .ZN(n11211) );
  OAI21_X2 U11587 ( .B1(n18668), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n15191), 
        .ZN(n19312) );
  INV_X1 U11588 ( .A(n19312), .ZN(n19683) );
  NAND2_X1 U11589 ( .A1(n16913), .A2(n11096), .ZN(n13513) );
  INV_X1 U11590 ( .A(n18796), .ZN(n20625) );
  NAND3_X1 U11591 ( .A1(n13386), .A2(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17857) );
  NAND2_X1 U11592 ( .A1(n17975), .A2(n17923), .ZN(n17840) );
  NAND2_X1 U11593 ( .A1(n11282), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11289) );
  AND2_X1 U11594 ( .A1(n18010), .A2(n21135), .ZN(n11288) );
  NAND2_X1 U11595 ( .A1(n13999), .A2(n14000), .ZN(n18073) );
  XNOR2_X1 U11596 ( .A(n14029), .B(n14030), .ZN(n18068) );
  OR2_X1 U11597 ( .A1(n18068), .A2(n20884), .ZN(n11189) );
  OR2_X1 U11598 ( .A1(n18108), .A2(n18107), .ZN(n11200) );
  AOI22_X1 U11599 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13487) );
  AOI22_X1 U11600 ( .A1(n17689), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17585), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13488) );
  AOI211_X1 U11601 ( .C1(n17465), .C2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A(
        n13485), .B(n13484), .ZN(n13486) );
  NAND2_X1 U11602 ( .A1(n13370), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n15599)
         );
  NOR2_X2 U11603 ( .A1(n15124), .A2(n12623), .ZN(n15093) );
  INV_X2 U11604 ( .A(n15886), .ZN(n15887) );
  INV_X1 U11605 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21915) );
  INV_X1 U11606 ( .A(n21836), .ZN(n21850) );
  XNOR2_X1 U11607 ( .A(n14460), .B(n14459), .ZN(n16279) );
  OAI21_X1 U11608 ( .B1(n15604), .B2(n18447), .A(n13864), .ZN(n13865) );
  INV_X1 U11609 ( .A(n18538), .ZN(n18557) );
  AND2_X1 U11610 ( .A1(n18248), .A2(n13834), .ZN(n18560) );
  NOR2_X1 U11611 ( .A1(n19233), .A2(n18536), .ZN(n18537) );
  AND2_X1 U11612 ( .A1(n17222), .A2(n14553), .ZN(n17216) );
  INV_X1 U11613 ( .A(n17228), .ZN(n17258) );
  OR2_X1 U11614 ( .A1(n18686), .A2(n14419), .ZN(n17222) );
  INV_X1 U11615 ( .A(n17257), .ZN(n17227) );
  XNOR2_X1 U11616 ( .A(n11119), .B(n11022), .ZN(n14475) );
  NAND2_X1 U11617 ( .A1(n11120), .A2(n11029), .ZN(n11119) );
  OAI21_X1 U11618 ( .B1(n14473), .B2(n16853), .A(n14466), .ZN(n11117) );
  NAND2_X1 U11619 ( .A1(n11110), .A2(n11109), .ZN(n11113) );
  NOR2_X1 U11620 ( .A1(n11111), .A2(n11070), .ZN(n11109) );
  NAND2_X1 U11621 ( .A1(n10958), .A2(n11345), .ZN(n14410) );
  XNOR2_X1 U11622 ( .A(n16471), .B(n12202), .ZN(n16690) );
  CLKBUF_X1 U11623 ( .A(n16462), .Z(n16469) );
  OAI21_X1 U11624 ( .B1(n18576), .B2(n18575), .A(n11073), .ZN(n11072) );
  INV_X1 U11625 ( .A(n11074), .ZN(n11073) );
  OAI21_X1 U11626 ( .B1(n18579), .B2(n18609), .A(n18578), .ZN(n11074) );
  NAND2_X1 U11627 ( .A1(n11314), .A2(n11317), .ZN(n18371) );
  INV_X1 U11628 ( .A(n18575), .ZN(n18604) );
  INV_X1 U11629 ( .A(n18603), .ZN(n16853) );
  NAND2_X1 U11630 ( .A1(n12279), .A2(n18628), .ZN(n18575) );
  INV_X1 U11631 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19263) );
  NOR2_X1 U11632 ( .A1(n15181), .A2(n11055), .ZN(n18260) );
  INV_X1 U11633 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19233) );
  INV_X1 U11634 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19221) );
  XNOR2_X1 U11635 ( .A(n14765), .B(n14764), .ZN(n19447) );
  XNOR2_X1 U11636 ( .A(n14770), .B(n14769), .ZN(n19559) );
  XNOR2_X1 U11637 ( .A(n11142), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n20332) );
  NOR2_X1 U11638 ( .A1(n13391), .A2(n20538), .ZN(n11142) );
  NOR2_X1 U11639 ( .A1(n20722), .A2(n20565), .ZN(n20690) );
  INV_X1 U11640 ( .A(n20707), .ZN(n20708) );
  INV_X1 U11641 ( .A(n20661), .ZN(n20722) );
  NAND2_X1 U11642 ( .A1(n20729), .A2(P3_EAX_REG_8__SCAN_IN), .ZN(n20728) );
  OR2_X1 U11643 ( .A1(n18051), .A2(n11067), .ZN(n11195) );
  NOR2_X1 U11644 ( .A1(n21041), .A2(n21080), .ZN(n11208) );
  OR2_X1 U11645 ( .A1(n21100), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11207) );
  INV_X1 U11646 ( .A(n21024), .ZN(n11206) );
  NAND2_X1 U11647 ( .A1(n17754), .A2(n20870), .ZN(n21144) );
  NOR2_X1 U11648 ( .A1(n21080), .A2(n21190), .ZN(n20870) );
  AND4_X1 U11649 ( .A1(n11891), .A2(n11890), .A3(n11889), .A4(n11888), .ZN(
        n11897) );
  AND4_X1 U11650 ( .A1(n11839), .A2(n11838), .A3(n11837), .A4(n11836), .ZN(
        n11847) );
  AND2_X1 U11651 ( .A1(n12635), .A2(n12628), .ZN(n12629) );
  NAND2_X1 U11652 ( .A1(n11476), .A2(n11475), .ZN(n11520) );
  XNOR2_X1 U11653 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n11519) );
  OAI211_X1 U11654 ( .C1(n11823), .C2(n19669), .A(n11338), .B(n11337), .ZN(
        n11783) );
  NAND2_X1 U11655 ( .A1(n11336), .A2(n11335), .ZN(n11337) );
  AND2_X1 U11656 ( .A1(n11597), .A2(n11613), .ZN(n11601) );
  OR2_X1 U11657 ( .A1(n13503), .A2(n13504), .ZN(n13499) );
  OR2_X1 U11658 ( .A1(n12805), .A2(n12804), .ZN(n13723) );
  OR2_X1 U11659 ( .A1(n12780), .A2(n12779), .ZN(n13703) );
  INV_X1 U11660 ( .A(n13737), .ZN(n12808) );
  NAND2_X1 U11661 ( .A1(n12829), .A2(n12827), .ZN(n12651) );
  XNOR2_X1 U11662 ( .A(n12649), .B(n11379), .ZN(n15116) );
  NOR2_X1 U11663 ( .A1(n11927), .A2(n11915), .ZN(n11186) );
  CLKBUF_X1 U11664 ( .A(n14200), .Z(n14351) );
  NOR2_X1 U11665 ( .A1(n11910), .A2(n11908), .ZN(n11573) );
  NOR2_X1 U11666 ( .A1(n10992), .A2(n11169), .ZN(n11168) );
  NOR2_X1 U11667 ( .A1(n11925), .A2(n11923), .ZN(n11921) );
  CLKBUF_X1 U11668 ( .A(n12057), .Z(n12252) );
  NAND2_X1 U11669 ( .A1(n11669), .A2(n11640), .ZN(n12250) );
  NOR2_X1 U11670 ( .A1(n11668), .A2(n11661), .ZN(n11640) );
  NAND2_X1 U11671 ( .A1(n11356), .A2(n11331), .ZN(n12063) );
  INV_X1 U11672 ( .A(n11782), .ZN(n11336) );
  AOI22_X1 U11673 ( .A1(n11645), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11633), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11637) );
  AOI22_X1 U11674 ( .A1(n15319), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14200), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11629) );
  AOI22_X1 U11675 ( .A1(n15319), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14200), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11604) );
  AOI21_X1 U11676 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n21204), .A(
        n13498), .ZN(n13504) );
  AND2_X1 U11677 ( .A1(n13868), .A2(n13872), .ZN(n13498) );
  NAND2_X1 U11678 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20795), .ZN(
        n13403) );
  NAND2_X1 U11679 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20759), .ZN(
        n13400) );
  NOR2_X1 U11680 ( .A1(n11275), .A2(n11272), .ZN(n11271) );
  INV_X1 U11681 ( .A(n15697), .ZN(n11275) );
  INV_X1 U11682 ( .A(n11273), .ZN(n11272) );
  NOR2_X1 U11683 ( .A1(n13063), .A2(n11262), .ZN(n11261) );
  INV_X1 U11684 ( .A(n11263), .ZN(n11262) );
  INV_X1 U11685 ( .A(n13299), .ZN(n13269) );
  AND2_X1 U11686 ( .A1(n15540), .A2(n15768), .ZN(n11263) );
  OAI211_X1 U11687 ( .C1(n12795), .C2(n11258), .A(n11257), .B(n11256), .ZN(
        n13721) );
  OR2_X1 U11688 ( .A1(n11259), .A2(n11258), .ZN(n11257) );
  AND2_X1 U11689 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n12811), .ZN(
        n12848) );
  NOR2_X1 U11690 ( .A1(n13615), .A2(n11229), .ZN(n11228) );
  INV_X1 U11691 ( .A(n15676), .ZN(n11229) );
  NOR2_X1 U11692 ( .A1(n15762), .A2(n15746), .ZN(n11244) );
  NOR2_X1 U11693 ( .A1(n15828), .A2(n11242), .ZN(n11241) );
  INV_X1 U11694 ( .A(n15771), .ZN(n11242) );
  INV_X1 U11695 ( .A(n13606), .ZN(n13616) );
  INV_X1 U11696 ( .A(n13700), .ZN(n11285) );
  OR2_X1 U11697 ( .A1(n12767), .A2(n12766), .ZN(n13688) );
  NAND2_X1 U11698 ( .A1(n12625), .A2(n12624), .ZN(n12638) );
  AND2_X1 U11699 ( .A1(n14866), .A2(n15096), .ZN(n12624) );
  NAND2_X1 U11700 ( .A1(n14871), .A2(n14948), .ZN(n12619) );
  NAND2_X1 U11701 ( .A1(n13341), .A2(n13720), .ZN(n13344) );
  OAI21_X1 U11702 ( .B1(n13341), .B2(n13350), .A(n13340), .ZN(n13342) );
  AND3_X1 U11703 ( .A1(n11331), .A2(n11684), .A3(n11685), .ZN(n11114) );
  AND2_X1 U11704 ( .A1(n11691), .A2(n12015), .ZN(n12037) );
  NOR2_X1 U11705 ( .A1(n16298), .A2(n16299), .ZN(n11320) );
  OR2_X1 U11706 ( .A1(n11990), .A2(n11988), .ZN(n11590) );
  NAND2_X1 U11707 ( .A1(n11578), .A2(n11577), .ZN(n11930) );
  NOR2_X1 U11708 ( .A1(n13849), .A2(n11575), .ZN(n11923) );
  NAND2_X1 U11709 ( .A1(n11573), .A2(n11188), .ZN(n11925) );
  INV_X1 U11710 ( .A(n11912), .ZN(n11188) );
  NOR2_X1 U11711 ( .A1(n11856), .A2(n11857), .ZN(n11903) );
  NAND2_X1 U11712 ( .A1(n19400), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n11458) );
  NAND2_X1 U11713 ( .A1(n13849), .A2(n12035), .ZN(n11459) );
  NOR2_X1 U11714 ( .A1(n15419), .A2(n11214), .ZN(n11213) );
  INV_X1 U11715 ( .A(n15408), .ZN(n11214) );
  NOR2_X2 U11716 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11414) );
  CLKBUF_X1 U11717 ( .A(n14373), .Z(n14364) );
  CLKBUF_X1 U11718 ( .A(n15319), .Z(n14372) );
  NOR2_X1 U11719 ( .A1(n16232), .A2(n14282), .ZN(n14303) );
  AND2_X1 U11720 ( .A1(n14280), .A2(n14281), .ZN(n14282) );
  INV_X1 U11721 ( .A(n16251), .ZN(n11361) );
  NAND2_X1 U11722 ( .A1(n16207), .A2(n16217), .ZN(n11238) );
  NOR2_X1 U11723 ( .A1(n18512), .A2(n11154), .ZN(n11153) );
  INV_X1 U11724 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n11154) );
  NOR2_X1 U11725 ( .A1(n16461), .A2(n11148), .ZN(n11147) );
  NAND2_X1 U11726 ( .A1(n11426), .A2(n11425), .ZN(n12298) );
  INV_X1 U11727 ( .A(n11573), .ZN(n11911) );
  NOR2_X1 U11728 ( .A1(n14461), .A2(n16381), .ZN(n11352) );
  NOR2_X1 U11729 ( .A1(n11238), .A2(n12240), .ZN(n11237) );
  NAND2_X1 U11730 ( .A1(n11320), .A2(n11319), .ZN(n16290) );
  INV_X1 U11731 ( .A(n16292), .ZN(n11319) );
  INV_X1 U11732 ( .A(n11168), .ZN(n11167) );
  NOR2_X1 U11733 ( .A1(n18510), .A2(n14411), .ZN(n16368) );
  INV_X1 U11734 ( .A(n11332), .ZN(n11171) );
  OR2_X1 U11735 ( .A1(n11333), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11332) );
  AND2_X1 U11736 ( .A1(n16477), .A2(n16491), .ZN(n16450) );
  AND2_X1 U11737 ( .A1(n16722), .A2(n12271), .ZN(n11353) );
  AND2_X1 U11738 ( .A1(n12174), .A2(n12173), .ZN(n14488) );
  XNOR2_X1 U11739 ( .A(n12104), .B(n14411), .ZN(n12106) );
  NAND2_X1 U11740 ( .A1(n11739), .A2(n11738), .ZN(n11080) );
  AND2_X1 U11741 ( .A1(n11862), .A2(n11861), .ZN(n11872) );
  NAND2_X1 U11742 ( .A1(n11083), .A2(n11822), .ZN(n11860) );
  NAND2_X1 U11743 ( .A1(n11084), .A2(n11774), .ZN(n11083) );
  NAND2_X1 U11744 ( .A1(n11860), .A2(n11859), .ZN(n12086) );
  AOI21_X1 U11745 ( .B1(n12241), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n11707), 
        .ZN(n11708) );
  INV_X1 U11746 ( .A(n12237), .ZN(n11709) );
  NAND2_X1 U11747 ( .A1(n11803), .A2(n11802), .ZN(n12285) );
  OR2_X1 U11748 ( .A1(n14320), .A2(n19669), .ZN(n14081) );
  NAND2_X1 U11749 ( .A1(n11081), .A2(n10971), .ZN(n11660) );
  OAI22_X1 U11750 ( .A1(n11438), .A2(n11437), .B1(n11436), .B2(n11435), .ZN(
        n11682) );
  NAND2_X1 U11751 ( .A1(n11432), .A2(n11431), .ZN(n11436) );
  AND2_X1 U11752 ( .A1(n11669), .A2(n11081), .ZN(n11670) );
  NAND2_X1 U11753 ( .A1(n20661), .A2(n13475), .ZN(n13970) );
  INV_X1 U11754 ( .A(n18878), .ZN(n17346) );
  NOR2_X1 U11755 ( .A1(n13403), .A2(n13400), .ZN(n13982) );
  INV_X1 U11756 ( .A(n13392), .ZN(n13479) );
  NAND2_X1 U11757 ( .A1(n20750), .A2(n13497), .ZN(n20562) );
  NOR2_X1 U11758 ( .A1(n17857), .A2(n17860), .ZN(n17872) );
  NOR2_X1 U11759 ( .A1(n13979), .A2(n14016), .ZN(n13980) );
  AOI211_X1 U11760 ( .C1(n17922), .C2(n14041), .A(n14011), .B(n17876), .ZN(
        n14012) );
  NAND2_X1 U11761 ( .A1(n18043), .A2(n14004), .ZN(n11283) );
  NAND2_X1 U11762 ( .A1(n11189), .A2(n11027), .ZN(n14033) );
  NOR2_X1 U11763 ( .A1(n20746), .A2(n11095), .ZN(n13889) );
  NOR2_X1 U11764 ( .A1(n11096), .A2(n13476), .ZN(n11095) );
  OR2_X1 U11765 ( .A1(n16900), .A2(n11097), .ZN(n20749) );
  OR2_X1 U11766 ( .A1(n20103), .A2(n13491), .ZN(n11097) );
  AND2_X1 U11767 ( .A1(n13490), .A2(n19007), .ZN(n13491) );
  NOR2_X1 U11768 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n20776) );
  NOR2_X1 U11769 ( .A1(n20789), .A2(n20748), .ZN(n17510) );
  NOR2_X1 U11770 ( .A1(n20749), .A2(n20779), .ZN(n20760) );
  INV_X1 U11771 ( .A(n21190), .ZN(n17748) );
  INV_X1 U11772 ( .A(n21459), .ZN(n21483) );
  NAND2_X1 U11773 ( .A1(n15759), .A2(n15760), .ZN(n15762) );
  AND2_X1 U11774 ( .A1(n13549), .A2(n13548), .ZN(n14960) );
  XNOR2_X1 U11775 ( .A(n13541), .B(n14685), .ZN(n21415) );
  AND2_X1 U11776 ( .A1(n14828), .A2(n15617), .ZN(n19857) );
  OR2_X1 U11777 ( .A1(n13236), .A2(n15918), .ZN(n13238) );
  OR2_X1 U11778 ( .A1(n13238), .A2(n13237), .ZN(n13275) );
  INV_X1 U11779 ( .A(n11266), .ZN(n11264) );
  AND2_X1 U11780 ( .A1(n13197), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13198) );
  NAND2_X1 U11781 ( .A1(n13198), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13236) );
  NAND2_X1 U11782 ( .A1(n13160), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n13196) );
  NOR2_X1 U11783 ( .A1(n13127), .A2(n15966), .ZN(n13128) );
  NAND2_X1 U11784 ( .A1(n13753), .A2(n13735), .ZN(n15955) );
  NAND2_X1 U11785 ( .A1(n13755), .A2(n19975), .ZN(n15956) );
  OR2_X1 U11786 ( .A1(n15959), .A2(n13302), .ZN(n13132) );
  AND2_X1 U11787 ( .A1(n13112), .A2(n13111), .ZN(n15726) );
  AND2_X1 U11788 ( .A1(n13097), .A2(n13096), .ZN(n15743) );
  CLKBUF_X1 U11789 ( .A(n15724), .Z(n15725) );
  NOR2_X1 U11790 ( .A1(n13059), .A2(n21545), .ZN(n13026) );
  NAND2_X1 U11791 ( .A1(n13026), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13093) );
  NOR2_X1 U11792 ( .A1(n13025), .A2(n16004), .ZN(n13060) );
  NAND2_X1 U11793 ( .A1(n12995), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n13025) );
  NAND2_X1 U11794 ( .A1(n15787), .A2(n11263), .ZN(n15834) );
  NOR2_X1 U11795 ( .A1(n12981), .A2(n15794), .ZN(n12995) );
  OR2_X1 U11796 ( .A1(n13735), .A2(n21274), .ZN(n19992) );
  AND2_X1 U11797 ( .A1(n15787), .A2(n15540), .ZN(n15769) );
  AND2_X1 U11798 ( .A1(n13735), .A2(n21315), .ZN(n16013) );
  NOR2_X1 U11799 ( .A1(n12933), .A2(n21502), .ZN(n12934) );
  NAND2_X1 U11800 ( .A1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n12934), .ZN(
        n12972) );
  NOR2_X1 U11801 ( .A1(n12903), .A2(n12902), .ZN(n12917) );
  INV_X1 U11802 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12902) );
  CLKBUF_X1 U11803 ( .A(n15431), .Z(n15432) );
  AND2_X1 U11804 ( .A1(n11254), .A2(n11253), .ZN(n11250) );
  NAND2_X1 U11805 ( .A1(n12880), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12903) );
  CLKBUF_X1 U11806 ( .A(n15086), .Z(n15262) );
  NOR2_X1 U11807 ( .A1(n12879), .A2(n21455), .ZN(n12880) );
  AND2_X1 U11808 ( .A1(n12848), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12873) );
  NAND2_X1 U11809 ( .A1(n12870), .A2(n12869), .ZN(n15079) );
  INV_X1 U11810 ( .A(n14998), .ZN(n12869) );
  NAND2_X1 U11811 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12849) );
  OAI21_X1 U11812 ( .B1(n14911), .B2(n12978), .A(n12823), .ZN(n12824) );
  OR2_X1 U11813 ( .A1(n12842), .A2(n14821), .ZN(n12843) );
  INV_X1 U11814 ( .A(n12978), .ZN(n14820) );
  NAND2_X1 U11815 ( .A1(n20009), .A2(n11310), .ZN(n11309) );
  NAND2_X1 U11816 ( .A1(n15689), .A2(n11228), .ZN(n15658) );
  NAND2_X1 U11817 ( .A1(n13759), .A2(n11308), .ZN(n15917) );
  NOR2_X1 U11818 ( .A1(n15727), .A2(n15711), .ZN(n15712) );
  NAND2_X1 U11819 ( .A1(n11244), .A2(n11243), .ZN(n15727) );
  INV_X1 U11820 ( .A(n15729), .ZN(n11243) );
  INV_X1 U11821 ( .A(n11244), .ZN(n15748) );
  AND2_X1 U11822 ( .A1(n15542), .A2(n11239), .ZN(n15823) );
  NOR2_X1 U11823 ( .A1(n11240), .A2(n15822), .ZN(n11239) );
  INV_X1 U11824 ( .A(n11241), .ZN(n11240) );
  OR2_X1 U11825 ( .A1(n13735), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n20007) );
  NAND2_X1 U11826 ( .A1(n15542), .A2(n11241), .ZN(n15831) );
  NAND2_X1 U11827 ( .A1(n15542), .A2(n15771), .ZN(n15829) );
  NOR2_X1 U11828 ( .A1(n15792), .A2(n15791), .ZN(n15790) );
  OR2_X1 U11829 ( .A1(n15535), .A2(n15534), .ZN(n15792) );
  INV_X1 U11830 ( .A(n11295), .ZN(n11293) );
  NOR2_X1 U11831 ( .A1(n15491), .A2(n15490), .ZN(n15524) );
  OR2_X1 U11832 ( .A1(n15446), .A2(n15445), .ZN(n15491) );
  OR2_X1 U11833 ( .A1(n15399), .A2(n15398), .ZN(n15446) );
  AND2_X1 U11834 ( .A1(n15088), .A2(n15089), .ZN(n15276) );
  NAND2_X1 U11835 ( .A1(n15276), .A2(n15275), .ZN(n15399) );
  NOR2_X1 U11836 ( .A1(n15083), .A2(n15082), .ZN(n15088) );
  NAND2_X1 U11837 ( .A1(n14836), .A2(n14960), .ZN(n14985) );
  AND2_X1 U11838 ( .A1(n13552), .A2(n13551), .ZN(n14984) );
  OR2_X1 U11839 ( .A1(n14985), .A2(n14984), .ZN(n15083) );
  AND2_X1 U11840 ( .A1(n14944), .A2(n21401), .ZN(n16031) );
  INV_X1 U11841 ( .A(n21332), .ZN(n16041) );
  NAND2_X1 U11842 ( .A1(n12826), .A2(n12825), .ZN(n12815) );
  OAI21_X1 U11843 ( .B1(n14715), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n12746), 
        .ZN(n12816) );
  INV_X1 U11844 ( .A(n12745), .ZN(n12746) );
  INV_X1 U11846 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14746) );
  OR2_X1 U11847 ( .A1(n10980), .A2(n21850), .ZN(n21893) );
  INV_X1 U11848 ( .A(n15596), .ZN(n15156) );
  NAND2_X1 U11849 ( .A1(n21593), .A2(n15123), .ZN(n16175) );
  OR2_X1 U11850 ( .A1(n14911), .A2(n15112), .ZN(n21921) );
  OR2_X1 U11851 ( .A1(n15613), .A2(n14859), .ZN(n16965) );
  INV_X1 U11852 ( .A(n18630), .ZN(n18640) );
  AND2_X1 U11853 ( .A1(n11997), .A2(n11998), .ZN(n13848) );
  NOR2_X1 U11854 ( .A1(n11590), .A2(n11589), .ZN(n11997) );
  INV_X1 U11855 ( .A(n11320), .ZN(n16301) );
  AND2_X1 U11856 ( .A1(n11328), .A2(n16330), .ZN(n11327) );
  INV_X1 U11857 ( .A(n11584), .ZN(n11934) );
  NOR3_X1 U11858 ( .A1(n11944), .A2(n11177), .A3(n11938), .ZN(n11936) );
  OR2_X1 U11859 ( .A1(n11150), .A2(n18394), .ZN(n11149) );
  AND2_X1 U11860 ( .A1(n11578), .A2(n11184), .ZN(n11946) );
  MUX2_X1 U11861 ( .A(n12292), .B(n11471), .S(n11685), .Z(n11868) );
  AND2_X1 U11862 ( .A1(n11237), .A2(n11235), .ZN(n11234) );
  INV_X1 U11863 ( .A(n14448), .ZN(n11235) );
  AND2_X1 U11864 ( .A1(n12220), .A2(n12219), .ZN(n16244) );
  AND2_X1 U11865 ( .A1(n12196), .A2(n12195), .ZN(n16265) );
  AND2_X1 U11866 ( .A1(n12189), .A2(n12188), .ZN(n15498) );
  NAND2_X1 U11867 ( .A1(n14489), .A2(n11213), .ZN(n15499) );
  NAND2_X1 U11868 ( .A1(n14489), .A2(n15408), .ZN(n15420) );
  OR2_X1 U11870 ( .A1(n11419), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14219) );
  OR2_X1 U11871 ( .A1(n14339), .A2(n14338), .ZN(n16212) );
  AND2_X1 U11872 ( .A1(n16314), .A2(n16315), .ZN(n16309) );
  AND2_X1 U11873 ( .A1(n16691), .A2(n11328), .ZN(n16668) );
  NAND2_X1 U11874 ( .A1(n16691), .A2(n11330), .ZN(n16669) );
  AND2_X1 U11875 ( .A1(n15505), .A2(n14167), .ZN(n15559) );
  AND2_X1 U11876 ( .A1(n14138), .A2(n10997), .ZN(n11362) );
  AND2_X1 U11877 ( .A1(n10990), .A2(n16807), .ZN(n11321) );
  AND3_X1 U11878 ( .A1(n12384), .A2(n12383), .A3(n12382), .ZN(n16792) );
  NAND2_X1 U11879 ( .A1(n12326), .A2(n12325), .ZN(n16870) );
  AND2_X1 U11880 ( .A1(n14624), .A2(n21645), .ZN(n17294) );
  INV_X1 U11881 ( .A(n14398), .ZN(n15196) );
  NAND2_X1 U11882 ( .A1(n13815), .A2(n11153), .ZN(n13821) );
  NAND2_X1 U11883 ( .A1(n15515), .A2(n11058), .ZN(n16255) );
  AND2_X1 U11884 ( .A1(n11058), .A2(n11224), .ZN(n11223) );
  INV_X1 U11885 ( .A(n16248), .ZN(n11224) );
  CLKBUF_X1 U11886 ( .A(n16408), .Z(n16463) );
  INV_X1 U11887 ( .A(n13790), .ZN(n13785) );
  AND2_X1 U11888 ( .A1(n12154), .A2(n12153), .ZN(n14992) );
  NOR2_X1 U11889 ( .A1(n14991), .A2(n14992), .ZN(n15061) );
  NOR2_X1 U11890 ( .A1(n11146), .A2(n17223), .ZN(n11143) );
  NAND2_X1 U11891 ( .A1(n11112), .A2(n16610), .ZN(n11111) );
  INV_X1 U11892 ( .A(n12115), .ZN(n11112) );
  OR2_X1 U11893 ( .A1(n11348), .A2(n11019), .ZN(n11345) );
  NOR2_X1 U11894 ( .A1(n11588), .A2(n12505), .ZN(n14441) );
  INV_X1 U11895 ( .A(n11999), .ZN(n16369) );
  AND2_X1 U11896 ( .A1(n12232), .A2(n12231), .ZN(n16224) );
  AND2_X1 U11897 ( .A1(n12003), .A2(n16637), .ZN(n16400) );
  AND2_X1 U11898 ( .A1(n12004), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16401) );
  AND2_X1 U11899 ( .A1(n11031), .A2(n11342), .ZN(n11341) );
  NAND2_X1 U11900 ( .A1(n16454), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11342) );
  NOR2_X1 U11901 ( .A1(n18436), .A2(n14411), .ZN(n16454) );
  NOR2_X1 U11902 ( .A1(n10996), .A2(n16749), .ZN(n11315) );
  AND2_X1 U11903 ( .A1(n12476), .A2(n12475), .ZN(n16741) );
  NAND2_X1 U11904 ( .A1(n16516), .A2(n16515), .ZN(n16514) );
  NOR2_X1 U11905 ( .A1(n11318), .A2(n18359), .ZN(n11317) );
  INV_X1 U11906 ( .A(n14486), .ZN(n11318) );
  AND2_X1 U11907 ( .A1(n16579), .A2(n18568), .ZN(n16541) );
  NOR2_X1 U11908 ( .A1(n16777), .A2(n18359), .ZN(n18358) );
  NAND2_X1 U11909 ( .A1(n16439), .A2(n16440), .ZN(n16441) );
  AND2_X1 U11910 ( .A1(n12110), .A2(n12105), .ZN(n16820) );
  AND2_X1 U11911 ( .A1(n12149), .A2(n12148), .ZN(n14964) );
  NAND2_X1 U11912 ( .A1(n11102), .A2(n16834), .ZN(n11100) );
  INV_X1 U11913 ( .A(n14931), .ZN(n12142) );
  CLKBUF_X1 U11914 ( .A(n15287), .Z(n15288) );
  NOR2_X1 U11915 ( .A1(n11729), .A2(n11730), .ZN(n11086) );
  AND2_X1 U11916 ( .A1(n12286), .A2(n19233), .ZN(n11313) );
  NOR2_X1 U11917 ( .A1(n14806), .A2(n14807), .ZN(n14808) );
  NAND2_X1 U11918 ( .A1(n12305), .A2(n11325), .ZN(n11324) );
  INV_X1 U11919 ( .A(n14661), .ZN(n11325) );
  INV_X1 U11920 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15176) );
  CLKBUF_X1 U11921 ( .A(n11412), .Z(n15280) );
  NOR2_X1 U11922 ( .A1(n11389), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11411) );
  INV_X1 U11923 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11389) );
  AND2_X1 U11924 ( .A1(n14084), .A2(n14074), .ZN(n14770) );
  AND2_X1 U11925 ( .A1(n14087), .A2(n14065), .ZN(n14760) );
  OR2_X1 U11926 ( .A1(n19447), .A2(n15383), .ZN(n19307) );
  NAND2_X1 U11927 ( .A1(n19312), .A2(n19292), .ZN(n19332) );
  NAND2_X1 U11928 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19312), .ZN(n19685) );
  NAND2_X1 U11929 ( .A1(n19447), .A2(n15383), .ZN(n19290) );
  NAND2_X1 U11930 ( .A1(n19330), .A2(n19559), .ZN(n19198) );
  NAND2_X1 U11931 ( .A1(n12031), .A2(n12030), .ZN(n18626) );
  INV_X1 U11932 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n17266) );
  NOR2_X1 U11933 ( .A1(n16900), .A2(n20562), .ZN(n21187) );
  NAND2_X1 U11934 ( .A1(n20433), .A2(n10967), .ZN(n20443) );
  NAND2_X1 U11935 ( .A1(n20443), .A2(n20444), .ZN(n20442) );
  AND2_X1 U11936 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n11052), .ZN(
        n11137) );
  NOR2_X1 U11937 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n20241), .ZN(n20251) );
  NOR2_X1 U11938 ( .A1(n21223), .A2(n13513), .ZN(n20440) );
  INV_X1 U11939 ( .A(n20769), .ZN(n20155) );
  NAND4_X1 U11940 ( .A1(n21176), .A2(n20099), .A3(n21229), .A4(n21241), .ZN(
        n20548) );
  NOR2_X1 U11941 ( .A1(n20662), .A2(n11089), .ZN(n11088) );
  NAND3_X1 U11942 ( .A1(n13451), .A2(n13450), .A3(n13449), .ZN(n20624) );
  AND4_X1 U11943 ( .A1(n10993), .A2(n13447), .A3(n13446), .A4(n13444), .ZN(
        n13449) );
  OR2_X1 U11944 ( .A1(n20728), .A2(n20576), .ZN(n20622) );
  NOR2_X1 U11945 ( .A1(n13933), .A2(n13932), .ZN(n13978) );
  NOR2_X1 U11946 ( .A1(n20104), .A2(n16912), .ZN(n18192) );
  NAND2_X1 U11947 ( .A1(n17937), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13391) );
  NOR2_X1 U11948 ( .A1(n17962), .A2(n20523), .ZN(n17937) );
  NOR2_X1 U11949 ( .A1(n17893), .A2(n20495), .ZN(n17899) );
  INV_X1 U11950 ( .A(n17895), .ZN(n17893) );
  NOR2_X1 U11951 ( .A1(n17857), .A2(n11139), .ZN(n17895) );
  NAND2_X1 U11952 ( .A1(n11380), .A2(n11140), .ZN(n11139) );
  NOR2_X1 U11953 ( .A1(n17860), .A2(n20485), .ZN(n11140) );
  AND2_X1 U11954 ( .A1(n11131), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11130) );
  AND2_X1 U11955 ( .A1(n11132), .A2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11131) );
  NAND2_X1 U11956 ( .A1(n17974), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17750) );
  NOR2_X1 U11957 ( .A1(n17795), .A2(n20313), .ZN(n17990) );
  NOR2_X1 U11958 ( .A1(n18046), .A2(n20235), .ZN(n18047) );
  NOR2_X1 U11959 ( .A1(n21196), .A2(n21244), .ZN(n17749) );
  OR2_X1 U11960 ( .A1(n21068), .A2(n11201), .ZN(n21023) );
  NAND2_X1 U11961 ( .A1(n21039), .A2(n11202), .ZN(n11201) );
  INV_X1 U11962 ( .A(n11203), .ZN(n11202) );
  AOI21_X1 U11963 ( .B1(n21032), .B2(n21067), .A(n11304), .ZN(n11303) );
  INV_X1 U11964 ( .A(n14048), .ZN(n11304) );
  NOR2_X1 U11965 ( .A1(n17950), .A2(n21011), .ZN(n21030) );
  OAI21_X1 U11966 ( .B1(n14047), .B2(n20593), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11306) );
  NAND2_X1 U11967 ( .A1(n17906), .A2(n17748), .ZN(n14047) );
  NAND2_X1 U11968 ( .A1(n14041), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11203) );
  NAND2_X1 U11969 ( .A1(n11008), .A2(n18010), .ZN(n17915) );
  NOR2_X1 U11970 ( .A1(n17881), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17880) );
  AND2_X1 U11971 ( .A1(n11289), .A2(n21121), .ZN(n11287) );
  INV_X1 U11972 ( .A(n18010), .ZN(n17923) );
  INV_X1 U11973 ( .A(n11283), .ZN(n18012) );
  AND2_X1 U11974 ( .A1(n11198), .A2(n11197), .ZN(n20907) );
  NAND2_X1 U11975 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17775), .ZN(
        n20906) );
  OR2_X1 U11976 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17775), .ZN(
        n18030) );
  NAND2_X1 U11977 ( .A1(n18058), .A2(n14003), .ZN(n18044) );
  NAND2_X1 U11978 ( .A1(n18044), .A2(n18045), .ZN(n18043) );
  OR2_X1 U11979 ( .A1(n18051), .A2(n21172), .ZN(n11198) );
  XNOR2_X1 U11980 ( .A(n17773), .B(n11290), .ZN(n18059) );
  INV_X1 U11981 ( .A(n14002), .ZN(n11290) );
  OR2_X1 U11982 ( .A1(n14033), .A2(n14034), .ZN(n18060) );
  NAND2_X1 U11983 ( .A1(n18073), .A2(n18074), .ZN(n18072) );
  NOR2_X1 U11984 ( .A1(n14025), .A2(n18098), .ZN(n18084) );
  INV_X1 U11985 ( .A(n11199), .ZN(n14023) );
  NOR2_X1 U11986 ( .A1(n18084), .A2(n18083), .ZN(n18082) );
  INV_X1 U11987 ( .A(n13997), .ZN(n11300) );
  NAND2_X1 U11988 ( .A1(n18103), .A2(n13995), .ZN(n18092) );
  NAND2_X1 U11989 ( .A1(n18092), .A2(n18093), .ZN(n18091) );
  XNOR2_X1 U11990 ( .A(n11199), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18100) );
  NOR2_X1 U11991 ( .A1(n18100), .A2(n18099), .ZN(n18098) );
  INV_X1 U11992 ( .A(n20749), .ZN(n13971) );
  OAI21_X1 U11993 ( .B1(n13508), .B2(n13873), .A(n13874), .ZN(n21192) );
  NOR2_X1 U11994 ( .A1(n20093), .A2(n16899), .ZN(n21184) );
  INV_X1 U11995 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n20764) );
  INV_X1 U11996 ( .A(n21184), .ZN(n21119) );
  INV_X1 U11997 ( .A(n20624), .ZN(n18837) );
  NOR2_X2 U11998 ( .A1(n13462), .A2(n13461), .ZN(n18796) );
  NAND2_X1 U11999 ( .A1(n20095), .A2(n18717), .ZN(n19054) );
  INV_X1 U12000 ( .A(n15196), .ZN(n15195) );
  AOI21_X1 U12001 ( .B1(n15633), .B2(n15634), .A(n15632), .ZN(n11232) );
  OR2_X1 U12002 ( .A1(n21411), .A2(n13532), .ZN(n21571) );
  INV_X1 U12003 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n21455) );
  INV_X1 U12004 ( .A(n21571), .ZN(n21541) );
  OR2_X1 U12005 ( .A1(n21411), .A2(n21483), .ZN(n21552) );
  OR2_X1 U12006 ( .A1(n21411), .A2(n21902), .ZN(n21566) );
  NAND3_X1 U12007 ( .A1(n13639), .A2(n13638), .A3(n13637), .ZN(n21559) );
  NAND3_X1 U12008 ( .A1(n13638), .A2(n13636), .A3(n16941), .ZN(n21562) );
  INV_X1 U12009 ( .A(n21565), .ZN(n21535) );
  INV_X1 U12010 ( .A(n21566), .ZN(n21536) );
  AND2_X1 U12011 ( .A1(n13541), .A2(n11248), .ZN(n14838) );
  AND2_X2 U12012 ( .A1(n14690), .A2(n15620), .ZN(n19946) );
  INV_X1 U12013 ( .A(n15595), .ZN(n15877) );
  NOR2_X1 U12014 ( .A1(n15887), .A2(n14949), .ZN(n15888) );
  AND2_X1 U12015 ( .A1(n13359), .A2(n15620), .ZN(n15886) );
  OR2_X1 U12016 ( .A1(n14712), .A2(n13358), .ZN(n13359) );
  OR2_X1 U12017 ( .A1(n21729), .A2(n16174), .ZN(n21761) );
  NAND2_X1 U12018 ( .A1(n10987), .A2(n13781), .ZN(n15586) );
  OR2_X1 U12019 ( .A1(n13780), .A2(n13779), .ZN(n13781) );
  NAND2_X1 U12020 ( .A1(n13701), .A2(n13700), .ZN(n11286) );
  AND2_X1 U12021 ( .A1(n13649), .A2(n21876), .ZN(n20021) );
  XNOR2_X1 U12022 ( .A(n15631), .B(n15630), .ZN(n15802) );
  NAND2_X1 U12023 ( .A1(n13759), .A2(n13758), .ZN(n15924) );
  NAND2_X1 U12024 ( .A1(n11297), .A2(n11294), .ZN(n15457) );
  INV_X1 U12025 ( .A(n11296), .ZN(n11294) );
  AND2_X1 U12026 ( .A1(n14874), .A2(n14873), .ZN(n21394) );
  NAND2_X1 U12027 ( .A1(n14874), .A2(n15609), .ZN(n21332) );
  NAND2_X1 U12028 ( .A1(n14874), .A2(n16162), .ZN(n21402) );
  INV_X1 U12029 ( .A(n21394), .ZN(n21409) );
  AND2_X1 U12030 ( .A1(n14874), .A2(n14863), .ZN(n21406) );
  INV_X1 U12031 ( .A(n16976), .ZN(n21587) );
  INV_X1 U12032 ( .A(n21815), .ZN(n22227) );
  OAI21_X1 U12033 ( .B1(n21826), .B2(n22231), .A(n21942), .ZN(n22234) );
  OAI21_X1 U12034 ( .B1(n22258), .B2(n21867), .A(n21886), .ZN(n22261) );
  AOI21_X1 U12035 ( .B1(n21899), .B2(n21908), .A(n21898), .ZN(n22288) );
  INV_X1 U12036 ( .A(n21880), .ZN(n21934) );
  AND2_X1 U12037 ( .A1(n22145), .A2(n15858), .ZN(n22299) );
  OAI211_X1 U12038 ( .C1(n22296), .C2(n21943), .A(n21942), .B(n21941), .ZN(
        n22302) );
  INV_X1 U12039 ( .A(n21980), .ZN(n21983) );
  INV_X1 U12040 ( .A(n22019), .ZN(n22022) );
  INV_X1 U12041 ( .A(n22057), .ZN(n22060) );
  AND2_X1 U12042 ( .A1(n22145), .A2(n15867), .ZN(n22101) );
  AND2_X1 U12043 ( .A1(n22145), .A2(n22144), .ZN(n22200) );
  INV_X1 U12044 ( .A(n22179), .ZN(n22198) );
  OR2_X1 U12045 ( .A1(n16943), .A2(n16946), .ZN(n22310) );
  NOR2_X1 U12046 ( .A1(n15613), .A2(n21902), .ZN(n21597) );
  INV_X1 U12047 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16973) );
  XNOR2_X1 U12048 ( .A(n11997), .B(n11187), .ZN(n18523) );
  INV_X1 U12049 ( .A(n11998), .ZN(n11187) );
  XNOR2_X1 U12050 ( .A(n11990), .B(n11989), .ZN(n18499) );
  NAND2_X1 U12051 ( .A1(n11960), .A2(n11181), .ZN(n11983) );
  NAND2_X1 U12052 ( .A1(n11960), .A2(n11933), .ZN(n11977) );
  AND2_X1 U12053 ( .A1(n18248), .A2(n13852), .ZN(n18534) );
  OR2_X1 U12054 ( .A1(n15031), .A2(n11036), .ZN(n18384) );
  NAND2_X1 U12055 ( .A1(n18376), .A2(n18375), .ZN(n18374) );
  AND2_X1 U12056 ( .A1(n18248), .A2(n13846), .ZN(n18539) );
  INV_X1 U12057 ( .A(n18551), .ZN(n18536) );
  CLKBUF_X1 U12058 ( .A(n18537), .Z(n18524) );
  INV_X1 U12059 ( .A(n18560), .ZN(n18447) );
  AND2_X1 U12060 ( .A1(n15272), .A2(n15271), .ZN(n18352) );
  AND2_X1 U12061 ( .A1(n15058), .A2(n10997), .ZN(n15265) );
  INV_X1 U12062 ( .A(n14993), .ZN(n15058) );
  NAND2_X1 U12063 ( .A1(n15058), .A2(n11385), .ZN(n15224) );
  AND2_X1 U12064 ( .A1(n14916), .A2(n10999), .ZN(n14995) );
  INV_X1 U12065 ( .A(n16278), .ZN(n16252) );
  INV_X1 U12066 ( .A(n19559), .ZN(n19452) );
  INV_X1 U12067 ( .A(n18260), .ZN(n15383) );
  AND2_X1 U12068 ( .A1(n14647), .A2(n15195), .ZN(n19674) );
  AND2_X1 U12069 ( .A1(n14647), .A2(n15196), .ZN(n19673) );
  INV_X1 U12070 ( .A(n16352), .ZN(n19672) );
  AND2_X1 U12071 ( .A1(n19676), .A2(n19677), .ZN(n19349) );
  INV_X1 U12072 ( .A(n19612), .ZN(n19676) );
  AND2_X1 U12073 ( .A1(n19508), .A2(n14387), .ZN(n19612) );
  INV_X1 U12074 ( .A(n19508), .ZN(n19670) );
  NOR2_X1 U12075 ( .A1(n17294), .A2(n17321), .ZN(n17307) );
  CLKBUF_X1 U12077 ( .A(n17313), .Z(n17321) );
  NAND2_X1 U12078 ( .A1(n14507), .A2(n19621), .ZN(n14622) );
  INV_X1 U12079 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16581) );
  INV_X1 U12080 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16593) );
  INV_X1 U12081 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17223) );
  AND2_X1 U12082 ( .A1(n17222), .A2(n14420), .ZN(n17257) );
  INV_X1 U12083 ( .A(n17222), .ZN(n17245) );
  NAND2_X1 U12084 ( .A1(n11175), .A2(n16420), .ZN(n16412) );
  OR3_X1 U12085 ( .A1(n18597), .A2(n16679), .A3(n16704), .ZN(n16667) );
  AND2_X1 U12086 ( .A1(n16764), .A2(n16830), .ZN(n16774) );
  INV_X1 U12087 ( .A(n16774), .ZN(n16727) );
  XNOR2_X1 U12088 ( .A(n16439), .B(n16825), .ZN(n17237) );
  NAND2_X1 U12089 ( .A1(n15473), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15472) );
  XNOR2_X1 U12090 ( .A(n12098), .B(n12091), .ZN(n15473) );
  INV_X1 U12091 ( .A(n18382), .ZN(n18583) );
  AND2_X1 U12092 ( .A1(n16867), .A2(n16826), .ZN(n16764) );
  NAND2_X1 U12093 ( .A1(n11756), .A2(n11753), .ZN(n11754) );
  INV_X1 U12094 ( .A(n11159), .ZN(n11158) );
  NAND2_X1 U12095 ( .A1(n11326), .A2(n12305), .ZN(n14662) );
  INV_X1 U12096 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18619) );
  NAND2_X1 U12097 ( .A1(n14080), .A2(n14079), .ZN(n15181) );
  OR2_X1 U12098 ( .A1(n18258), .A2(n18652), .ZN(n14080) );
  NAND2_X1 U12099 ( .A1(n15047), .A2(n11359), .ZN(n16895) );
  INV_X1 U12100 ( .A(n19310), .ZN(n19316) );
  OAI21_X1 U12101 ( .B1(n19287), .B2(n19284), .A(n19283), .ZN(n19762) );
  NAND2_X1 U12102 ( .A1(n15198), .A2(n15197), .ZN(n19650) );
  NAND2_X1 U12103 ( .A1(n19273), .A2(n19272), .ZN(n19748) );
  NOR2_X1 U12104 ( .A1(n19256), .A2(n19290), .ZN(n19645) );
  NOR2_X1 U12105 ( .A1(n19276), .A2(n19256), .ZN(n19742) );
  NOR2_X2 U12106 ( .A1(n19220), .A2(n19307), .ZN(n19727) );
  INV_X1 U12107 ( .A(n19597), .ZN(n19607) );
  INV_X1 U12108 ( .A(n19428), .ZN(n19436) );
  INV_X1 U12109 ( .A(n19786), .ZN(n19790) );
  INV_X1 U12110 ( .A(n19545), .ZN(n19554) );
  INV_X1 U12111 ( .A(n19469), .ZN(n19696) );
  OAI21_X1 U12112 ( .B1(n15391), .B2(n15390), .A(n15389), .ZN(n19695) );
  INV_X1 U12113 ( .A(n19771), .ZN(n19793) );
  INV_X1 U12114 ( .A(n19603), .ZN(n19605) );
  INV_X1 U12115 ( .A(n19699), .ZN(n19566) );
  INV_X1 U12116 ( .A(n19433), .ZN(n19435) );
  INV_X1 U12117 ( .A(n19381), .ZN(n19389) );
  OR2_X1 U12118 ( .A1(n19198), .A2(n19290), .ZN(n19699) );
  INV_X1 U12119 ( .A(n19569), .ZN(n19789) );
  NAND2_X1 U12120 ( .A1(n18626), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18668) );
  NAND2_X1 U12121 ( .A1(n21221), .A2(n21188), .ZN(n20104) );
  INV_X1 U12122 ( .A(n16913), .ZN(n20099) );
  INV_X1 U12123 ( .A(n17749), .ZN(n21247) );
  INV_X1 U12124 ( .A(n20544), .ZN(n11123) );
  NAND2_X1 U12125 ( .A1(n20535), .A2(n10967), .ZN(n11126) );
  NAND2_X1 U12126 ( .A1(n11127), .A2(n10967), .ZN(n20530) );
  NOR2_X1 U12127 ( .A1(n11129), .A2(n17913), .ZN(n11128) );
  INV_X1 U12128 ( .A(n20516), .ZN(n11129) );
  NAND2_X1 U12129 ( .A1(n20499), .A2(n10967), .ZN(n20515) );
  NAND2_X1 U12130 ( .A1(n20515), .A2(n20516), .ZN(n20514) );
  NAND2_X1 U12131 ( .A1(n20500), .A2(n20501), .ZN(n20499) );
  NAND2_X1 U12132 ( .A1(n20415), .A2(n10967), .ZN(n20434) );
  NAND2_X1 U12133 ( .A1(n20434), .A2(n20435), .ZN(n20433) );
  NAND2_X1 U12134 ( .A1(n20408), .A2(n10967), .ZN(n20416) );
  NAND2_X1 U12135 ( .A1(n20416), .A2(n20417), .ZN(n20415) );
  INV_X1 U12136 ( .A(n20440), .ZN(n20549) );
  INV_X1 U12137 ( .A(n20546), .ZN(n20508) );
  NAND2_X1 U12138 ( .A1(n11136), .A2(n11137), .ZN(n20265) );
  INV_X1 U12139 ( .A(n20450), .ZN(n20537) );
  NOR2_X2 U12140 ( .A1(n21232), .A2(n20552), .ZN(n20450) );
  INV_X1 U12141 ( .A(n20548), .ZN(n20552) );
  NAND2_X1 U12142 ( .A1(n20697), .A2(n11004), .ZN(n20688) );
  NOR2_X1 U12143 ( .A1(n20702), .A2(n20661), .ZN(n20697) );
  NAND2_X1 U12144 ( .A1(n20697), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n20696) );
  NOR2_X1 U12145 ( .A1(n20710), .A2(n11098), .ZN(n20703) );
  NAND2_X1 U12146 ( .A1(n20703), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n20702) );
  INV_X1 U12147 ( .A(n20642), .ZN(n20631) );
  NOR2_X1 U12148 ( .A1(n20647), .A2(n20652), .ZN(n20646) );
  OR3_X1 U12149 ( .A1(n20661), .A2(n20710), .A3(n20623), .ZN(n20652) );
  NOR2_X1 U12150 ( .A1(n20716), .A2(n20726), .ZN(n20711) );
  NAND2_X1 U12151 ( .A1(n20711), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n20710) );
  NOR2_X1 U12152 ( .A1(n20735), .A2(n11099), .ZN(n20729) );
  NAND2_X1 U12153 ( .A1(n11003), .A2(n11068), .ZN(n11099) );
  NOR2_X1 U12154 ( .A1(n13913), .A2(n13912), .ZN(n20607) );
  AND2_X1 U12155 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n20606), .ZN(n20609) );
  NAND2_X1 U12156 ( .A1(n20746), .A2(n20590), .ZN(n20732) );
  OR4_X1 U12157 ( .A1(n20744), .A2(n20591), .A3(n20618), .A4(n20743), .ZN(
        n20615) );
  NAND2_X1 U12158 ( .A1(n20745), .A2(P3_EAX_REG_1__SCAN_IN), .ZN(n20735) );
  INV_X1 U12159 ( .A(n20690), .ZN(n20736) );
  INV_X1 U12160 ( .A(n13983), .ZN(n11190) );
  NOR2_X1 U12161 ( .A1(n20565), .A2(n20744), .ZN(n20745) );
  INV_X1 U12162 ( .A(n20732), .ZN(n20740) );
  INV_X1 U12163 ( .A(n20610), .ZN(n20741) );
  CLKBUF_X1 U12164 ( .A(n18203), .Z(n18211) );
  NOR2_X1 U12165 ( .A1(n20143), .A2(n20137), .ZN(n20140) );
  INV_X1 U12166 ( .A(n20139), .ZN(n20143) );
  NOR2_X1 U12168 ( .A1(n21068), .A2(n17888), .ZN(n17870) );
  NAND2_X1 U12169 ( .A1(n17974), .A2(n11131), .ZN(n17847) );
  NOR2_X1 U12170 ( .A1(n17778), .A2(n17788), .ZN(n17974) );
  NAND2_X1 U12171 ( .A1(n20593), .A2(n18081), .ZN(n17865) );
  NOR2_X1 U12172 ( .A1(n20938), .A2(n17994), .ZN(n20959) );
  INV_X1 U12173 ( .A(n17865), .ZN(n18052) );
  NOR2_X1 U12174 ( .A1(n18085), .A2(n20206), .ZN(n18070) );
  NAND2_X1 U12175 ( .A1(n18097), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18085) );
  INV_X1 U12176 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20206) );
  AND2_X1 U12177 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18097) );
  INV_X1 U12178 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n18110) );
  INV_X1 U12179 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20157) );
  NAND2_X1 U12180 ( .A1(n11305), .A2(n11301), .ZN(n14049) );
  INV_X1 U12181 ( .A(n11302), .ZN(n11301) );
  NAND2_X1 U12182 ( .A1(n11306), .A2(n17964), .ZN(n11305) );
  OAI21_X1 U12183 ( .B1(n21030), .B2(n21056), .A(n11303), .ZN(n11302) );
  AOI21_X1 U12184 ( .B1(n11196), .B2(n11067), .A(n20938), .ZN(n11193) );
  NAND2_X1 U12185 ( .A1(n21119), .A2(n21175), .ZN(n21147) );
  INV_X1 U12186 ( .A(n11189), .ZN(n18067) );
  INV_X1 U12187 ( .A(n11200), .ZN(n18106) );
  INV_X2 U12188 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n20759) );
  AOI211_X1 U12189 ( .C1(n21221), .C2(n21199), .A(n18718), .B(n16904), .ZN(
        n20796) );
  INV_X1 U12190 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18793) );
  CLKBUF_X2 U12191 ( .A(n21233), .Z(n20098) );
  OR2_X1 U12192 ( .A1(n21658), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18235) );
  INV_X1 U12193 ( .A(n15599), .ZN(n15121) );
  BUF_X1 U12194 ( .A(n18712), .Z(n19050) );
  NAND2_X1 U12195 ( .A1(n11233), .A2(n11230), .ZN(P1_U2810) );
  OR2_X1 U12196 ( .A1(n21562), .A2(n15802), .ZN(n11233) );
  INV_X1 U12197 ( .A(n11231), .ZN(n11230) );
  OAI21_X1 U12198 ( .B1(n15845), .B2(n21571), .A(n11232), .ZN(n11231) );
  AOI211_X1 U12199 ( .C1(n18560), .C2(n16196), .A(n18559), .B(n18558), .ZN(
        n18566) );
  OAI21_X1 U12200 ( .B1(n16209), .B2(P2_EBX_REG_3__SCAN_IN), .A(n11360), .ZN(
        n14763) );
  NAND2_X1 U12201 ( .A1(n16209), .A2(n14055), .ZN(n11360) );
  NAND2_X1 U12202 ( .A1(n11157), .A2(n17256), .ZN(n11156) );
  INV_X1 U12203 ( .A(n16607), .ZN(n11157) );
  OAI21_X1 U12204 ( .B1(n17227), .B2(n14055), .A(n15296), .ZN(n15297) );
  NAND2_X1 U12205 ( .A1(n11007), .A2(n16864), .ZN(n11115) );
  NOR2_X1 U12206 ( .A1(n14464), .A2(n11117), .ZN(n11116) );
  NAND2_X1 U12207 ( .A1(n14475), .A2(n18604), .ZN(n11118) );
  OAI21_X1 U12208 ( .B1(n12509), .B2(n18609), .A(n12508), .ZN(n12510) );
  NAND2_X1 U12209 ( .A1(n16690), .A2(n18604), .ZN(n16710) );
  INV_X1 U12210 ( .A(n11072), .ZN(n18580) );
  OAI21_X1 U12211 ( .B1(n11124), .B2(n21229), .A(n11122), .ZN(P3_U2641) );
  XNOR2_X1 U12212 ( .A(n11126), .B(n11125), .ZN(n11124) );
  NOR4_X1 U12213 ( .A1(n11014), .A2(n20541), .A3(n20540), .A4(n11123), .ZN(
        n11122) );
  INV_X1 U12214 ( .A(n20536), .ZN(n11125) );
  AOI21_X1 U12215 ( .B1(n20670), .B2(P3_EAX_REG_31__SCAN_IN), .A(n20669), .ZN(
        n20671) );
  OAI22_X1 U12216 ( .A1(n20676), .A2(n20690), .B1(P3_EAX_REG_30__SCAN_IN), 
        .B2(n20743), .ZN(n20670) );
  AOI21_X1 U12217 ( .B1(n11205), .B2(n11204), .A(n21025), .ZN(n21035) );
  NOR2_X1 U12218 ( .A1(n21167), .A2(n21033), .ZN(n11204) );
  AND2_X2 U12219 ( .A1(n20769), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13934) );
  OR2_X1 U12220 ( .A1(n15664), .A2(n11267), .ZN(n15635) );
  AND2_X2 U12221 ( .A1(n12520), .A2(n14730), .ZN(n12761) );
  NAND4_X1 U12222 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A4(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n13793) );
  NAND2_X1 U12223 ( .A1(n13789), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13799) );
  NAND2_X1 U12224 ( .A1(n11143), .A2(n11145), .ZN(n13791) );
  AND2_X1 U12225 ( .A1(n10995), .A2(n11385), .ZN(n10985) );
  AND4_X1 U12226 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_21__SCAN_IN), .A4(P3_EAX_REG_19__SCAN_IN), .ZN(n10986)
         );
  NOR2_X1 U12227 ( .A1(n13402), .A2(n13401), .ZN(n13468) );
  NOR2_X1 U12228 ( .A1(n13402), .A2(n13393), .ZN(n17361) );
  INV_X1 U12229 ( .A(n19057), .ZN(n11096) );
  INV_X1 U12230 ( .A(n15086), .ZN(n11254) );
  AND2_X1 U12231 ( .A1(n15724), .A2(n11273), .ZN(n10988) );
  AND2_X1 U12232 ( .A1(n15151), .A2(n13663), .ZN(n12626) );
  NAND2_X1 U12233 ( .A1(n11578), .A2(n11044), .ZN(n11941) );
  AND2_X1 U12234 ( .A1(n11322), .A2(n16847), .ZN(n10990) );
  AND3_X1 U12235 ( .A1(n11686), .A2(n11680), .A3(n11668), .ZN(n10991) );
  AND2_X1 U12236 ( .A1(n11333), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10992) );
  AND3_X1 U12237 ( .A1(n13443), .A2(n13445), .A3(n11041), .ZN(n10993) );
  INV_X1 U12238 ( .A(n11249), .ZN(n15368) );
  INV_X1 U12239 ( .A(n13793), .ZN(n11145) );
  NOR2_X1 U12240 ( .A1(n13788), .A2(n16569), .ZN(n13789) );
  AND3_X1 U12241 ( .A1(n11144), .A2(n11145), .A3(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n13792) );
  AND2_X1 U12242 ( .A1(n14915), .A2(n11375), .ZN(n10994) );
  OR2_X1 U12243 ( .A1(n12381), .A2(n12380), .ZN(n10995) );
  NAND2_X1 U12244 ( .A1(n11317), .A2(n11316), .ZN(n10996) );
  INV_X1 U12245 ( .A(n12057), .ZN(n11331) );
  NOR2_X1 U12246 ( .A1(n13799), .A2(n11152), .ZN(n13801) );
  AND2_X1 U12247 ( .A1(n10985), .A2(n15267), .ZN(n10997) );
  NAND2_X1 U12248 ( .A1(n15505), .A2(n11056), .ZN(n15548) );
  AND2_X1 U12249 ( .A1(n11153), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10998) );
  AND2_X1 U12250 ( .A1(n10994), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10999) );
  AND2_X1 U12251 ( .A1(n13808), .A2(n11147), .ZN(n11000) );
  AND2_X1 U12252 ( .A1(n13806), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13808) );
  AND2_X1 U12253 ( .A1(n14259), .A2(n19621), .ZN(n11001) );
  AND2_X1 U12254 ( .A1(n11056), .A2(n11361), .ZN(n11002) );
  NOR2_X1 U12255 ( .A1(n13819), .A2(n16360), .ZN(n13823) );
  NAND2_X1 U12256 ( .A1(n13815), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13817) );
  AND4_X1 U12257 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(P3_EAX_REG_7__SCAN_IN), 
        .A3(P3_EAX_REG_4__SCAN_IN), .A4(P3_EAX_REG_6__SCAN_IN), .ZN(n11003) );
  AND2_X1 U12258 ( .A1(n11088), .A2(P3_EAX_REG_26__SCAN_IN), .ZN(n11004) );
  INV_X2 U12259 ( .A(n17343), .ZN(n17340) );
  NAND2_X1 U12260 ( .A1(n16555), .A2(n11353), .ZN(n16468) );
  OR2_X1 U12261 ( .A1(n16408), .A2(n12115), .ZN(n11006) );
  XOR2_X1 U12262 ( .A(n11113), .B(n14468), .Z(n11007) );
  INV_X1 U12263 ( .A(n20559), .ZN(n19007) );
  NAND3_X2 U12264 ( .A1(n13488), .A2(n13487), .A3(n13486), .ZN(n20559) );
  AND2_X1 U12265 ( .A1(n11281), .A2(n14051), .ZN(n11008) );
  AND2_X1 U12266 ( .A1(n11172), .A2(n11332), .ZN(n11010) );
  INV_X1 U12267 ( .A(n18961), .ZN(n13476) );
  NAND2_X1 U12268 ( .A1(n15724), .A2(n15726), .ZN(n15709) );
  NOR2_X1 U12269 ( .A1(n16240), .A2(n16239), .ZN(n14280) );
  INV_X1 U12270 ( .A(n11121), .ZN(n12091) );
  NAND2_X1 U12271 ( .A1(n11334), .A2(n12100), .ZN(n11121) );
  NOR2_X1 U12272 ( .A1(n13793), .A2(n17223), .ZN(n13794) );
  NOR2_X1 U12273 ( .A1(n13799), .A2(n16558), .ZN(n13800) );
  AND2_X1 U12274 ( .A1(n11578), .A2(n11186), .ZN(n11011) );
  AND2_X1 U12275 ( .A1(n11960), .A2(n11180), .ZN(n11012) );
  AND2_X1 U12276 ( .A1(n20697), .A2(n11088), .ZN(n11013) );
  NOR2_X1 U12277 ( .A1(n20545), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n11014) );
  AND4_X1 U12278 ( .A1(n12530), .A2(n12529), .A3(n12528), .A4(n12527), .ZN(
        n11015) );
  NAND2_X1 U12279 ( .A1(n15955), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n13757) );
  NAND2_X1 U12280 ( .A1(n10989), .A2(n11211), .ZN(n11825) );
  AND2_X1 U12281 ( .A1(n11160), .A2(n11349), .ZN(n11746) );
  AND2_X1 U12282 ( .A1(n15787), .A2(n11261), .ZN(n11016) );
  INV_X1 U12283 ( .A(n11282), .ZN(n14007) );
  AND2_X1 U12284 ( .A1(n15329), .A2(n15074), .ZN(n11017) );
  OR2_X1 U12285 ( .A1(n11944), .A2(n11938), .ZN(n11018) );
  OR2_X1 U12286 ( .A1(n12005), .A2(n16401), .ZN(n11019) );
  AND2_X1 U12287 ( .A1(n15712), .A2(n15698), .ZN(n11020) );
  NOR2_X1 U12288 ( .A1(n14008), .A2(n11288), .ZN(n11021) );
  INV_X1 U12289 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11146) );
  NAND2_X1 U12290 ( .A1(n15689), .A2(n15676), .ZN(n15654) );
  XOR2_X1 U12291 ( .A(n14447), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .Z(
        n11022) );
  AND4_X1 U12292 ( .A1(n12571), .A2(n12570), .A3(n12569), .A4(n12568), .ZN(
        n11023) );
  NAND2_X1 U12293 ( .A1(n11158), .A2(n11160), .ZN(n11751) );
  NOR3_X1 U12294 ( .A1(n14051), .A2(n21144), .A3(n17908), .ZN(n11024) );
  XNOR2_X1 U12295 ( .A(n11960), .B(n11183), .ZN(n11962) );
  OR2_X2 U12296 ( .A1(n11782), .A2(n11772), .ZN(n11840) );
  AND2_X1 U12297 ( .A1(n14339), .A2(n14338), .ZN(n11026) );
  INV_X1 U12298 ( .A(n14066), .ZN(n15329) );
  NAND2_X1 U12299 ( .A1(n12623), .A2(n13663), .ZN(n13543) );
  INV_X1 U12300 ( .A(n13543), .ZN(n13547) );
  OR2_X1 U12301 ( .A1(n14029), .A2(n14030), .ZN(n11027) );
  AND2_X1 U12302 ( .A1(n11165), .A2(n11166), .ZN(n11028) );
  NOR2_X1 U12303 ( .A1(n14441), .A2(n14440), .ZN(n11029) );
  OR2_X1 U12304 ( .A1(n16364), .A2(n18575), .ZN(n11030) );
  NOR2_X1 U12305 ( .A1(n15456), .A2(n11296), .ZN(n11295) );
  AND2_X1 U12306 ( .A1(n16456), .A2(n11974), .ZN(n11031) );
  AND2_X1 U12307 ( .A1(n11812), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11032) );
  NAND2_X1 U12308 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14022), .ZN(
        n11033) );
  INV_X1 U12309 ( .A(n16408), .ZN(n11110) );
  NOR2_X1 U12310 ( .A1(n13735), .A2(n15466), .ZN(n11034) );
  NOR2_X1 U12311 ( .A1(n11996), .A2(n11171), .ZN(n11170) );
  NAND2_X1 U12312 ( .A1(n15724), .A2(n11271), .ZN(n15690) );
  INV_X1 U12313 ( .A(n20763), .ZN(n13967) );
  AND2_X1 U12314 ( .A1(n11155), .A2(n18375), .ZN(n11036) );
  AND2_X1 U12315 ( .A1(n15329), .A2(n11771), .ZN(n11037) );
  AND2_X1 U12316 ( .A1(n11343), .A2(n11345), .ZN(n11038) );
  INV_X1 U12317 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n20795) );
  AND2_X1 U12318 ( .A1(n11017), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11039) );
  AND2_X1 U12319 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11040) );
  OR2_X1 U12320 ( .A1(n11009), .A2(n13448), .ZN(n11041) );
  INV_X1 U12321 ( .A(n19326), .ZN(n19292) );
  NAND2_X1 U12322 ( .A1(n14916), .A2(n14915), .ZN(n14881) );
  AND2_X1 U12323 ( .A1(n15505), .A2(n11002), .ZN(n11042) );
  NAND2_X1 U12324 ( .A1(n13785), .A2(n11373), .ZN(n13788) );
  NAND2_X1 U12325 ( .A1(n15058), .A2(n11362), .ZN(n15504) );
  NAND2_X1 U12326 ( .A1(n15515), .A2(n15562), .ZN(n15561) );
  NAND2_X1 U12327 ( .A1(n11692), .A2(n11691), .ZN(n12251) );
  NAND2_X1 U12328 ( .A1(n15431), .A2(n15434), .ZN(n15433) );
  INV_X1 U12329 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15068) );
  NOR2_X1 U12330 ( .A1(n14487), .A2(n14488), .ZN(n14489) );
  AND2_X1 U12331 ( .A1(n15790), .A2(n15543), .ZN(n15542) );
  NOR2_X1 U12332 ( .A1(n15079), .A2(n15078), .ZN(n15080) );
  NAND2_X1 U12333 ( .A1(n11872), .A2(n11871), .ZN(n11856) );
  OR2_X1 U12334 ( .A1(n16777), .A2(n10996), .ZN(n11043) );
  NAND2_X1 U12335 ( .A1(n11459), .A2(n11458), .ZN(n11867) );
  NAND2_X1 U12336 ( .A1(n11880), .A2(n18279), .ZN(n15474) );
  NOR2_X1 U12337 ( .A1(n16750), .A2(n16741), .ZN(n16347) );
  AND2_X1 U12338 ( .A1(n15823), .A2(n15815), .ZN(n15759) );
  AND2_X1 U12339 ( .A1(n16691), .A2(n16692), .ZN(n15550) );
  NAND2_X1 U12340 ( .A1(n11255), .A2(n11254), .ZN(n15260) );
  INV_X1 U12341 ( .A(n16420), .ZN(n11169) );
  AND2_X2 U12342 ( .A1(n12518), .A2(n14730), .ZN(n12737) );
  NOR2_X1 U12343 ( .A1(n16332), .A2(n16323), .ZN(n16314) );
  NAND2_X1 U12344 ( .A1(n12063), .A2(n11354), .ZN(n12259) );
  NAND2_X1 U12345 ( .A1(n11250), .A2(n11255), .ZN(n11249) );
  AND2_X1 U12346 ( .A1(n11184), .A2(n11945), .ZN(n11044) );
  AND2_X1 U12347 ( .A1(n11384), .A2(n11517), .ZN(n12313) );
  AND2_X1 U12348 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11045) );
  NAND2_X1 U12349 ( .A1(n11253), .A2(n15441), .ZN(n11252) );
  INV_X1 U12350 ( .A(n11182), .ZN(n11181) );
  OR2_X1 U12351 ( .A1(n11975), .A2(n11183), .ZN(n11182) );
  AND3_X1 U12352 ( .A1(n12474), .A2(n12473), .A3(n12472), .ZN(n16749) );
  OR2_X1 U12353 ( .A1(n20009), .A2(n16077), .ZN(n11046) );
  AND2_X1 U12354 ( .A1(n11259), .A2(n11258), .ZN(n11047) );
  AND2_X1 U12355 ( .A1(n11213), .A2(n11212), .ZN(n11048) );
  AND2_X1 U12356 ( .A1(n11261), .A2(n15755), .ZN(n11049) );
  AND2_X1 U12357 ( .A1(n11147), .A2(n11045), .ZN(n11050) );
  AND2_X1 U12358 ( .A1(n11805), .A2(n12314), .ZN(n11051) );
  AND2_X1 U12359 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11052) );
  AND2_X1 U12360 ( .A1(n11021), .A2(n11289), .ZN(n11053) );
  INV_X1 U12361 ( .A(n12287), .ZN(n12479) );
  NAND2_X1 U12362 ( .A1(n12330), .A2(n12329), .ZN(n16848) );
  AND2_X1 U12363 ( .A1(n18686), .A2(n19621), .ZN(n17256) );
  NAND2_X1 U12364 ( .A1(n17974), .A2(n11132), .ZN(n11054) );
  INV_X1 U12365 ( .A(n11933), .ZN(n11183) );
  NAND2_X1 U12366 ( .A1(n14916), .A2(n10994), .ZN(n14933) );
  NAND2_X1 U12367 ( .A1(n16848), .A2(n16847), .ZN(n16838) );
  NAND3_X1 U12368 ( .A1(n11324), .A2(n15048), .A3(n11326), .ZN(n15049) );
  NAND2_X1 U12369 ( .A1(n13808), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13811) );
  AND2_X1 U12370 ( .A1(n11312), .A2(n14648), .ZN(n11055) );
  AND2_X1 U12371 ( .A1(n15549), .A2(n14167), .ZN(n11056) );
  NOR2_X1 U12372 ( .A1(n14991), .A2(n11216), .ZN(n15270) );
  OR2_X1 U12373 ( .A1(n14991), .A2(n11219), .ZN(n11057) );
  AND2_X1 U12374 ( .A1(n11225), .A2(n15562), .ZN(n11058) );
  INV_X1 U12375 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n16946) );
  AND2_X1 U12376 ( .A1(n19400), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n11059) );
  AND2_X1 U12377 ( .A1(n19400), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n11060) );
  NOR2_X1 U12378 ( .A1(n14991), .A2(n11221), .ZN(n15059) );
  NAND2_X1 U12379 ( .A1(n16848), .A2(n10990), .ZN(n11323) );
  AND2_X1 U12380 ( .A1(n17974), .A2(n11130), .ZN(n13386) );
  NOR2_X1 U12381 ( .A1(n13805), .A2(n16497), .ZN(n13806) );
  OR3_X1 U12382 ( .A1(n17857), .A2(n11141), .A3(n17860), .ZN(n11061) );
  INV_X1 U12383 ( .A(n11381), .ZN(n11155) );
  OR2_X1 U12384 ( .A1(n13799), .A2(n11150), .ZN(n11062) );
  AND2_X2 U12385 ( .A1(n14371), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14172) );
  AND2_X1 U12386 ( .A1(n11226), .A2(n15587), .ZN(n11063) );
  AND2_X1 U12387 ( .A1(n19400), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n11064) );
  NAND2_X1 U12388 ( .A1(n15058), .A2(n10985), .ZN(n11363) );
  INV_X1 U12389 ( .A(n11380), .ZN(n11141) );
  AND2_X1 U12390 ( .A1(n11002), .A2(n16243), .ZN(n11065) );
  INV_X1 U12391 ( .A(n11842), .ZN(n19232) );
  AND2_X1 U12392 ( .A1(n11324), .A2(n11326), .ZN(n11066) );
  NAND2_X1 U12393 ( .A1(n20264), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n17795) );
  AND2_X1 U12394 ( .A1(n13808), .A2(n11050), .ZN(n13813) );
  NAND2_X1 U12395 ( .A1(n13815), .A2(n10998), .ZN(n13819) );
  AND2_X1 U12396 ( .A1(n13813), .A2(n13786), .ZN(n13815) );
  AND3_X1 U12397 ( .A1(n13541), .A2(n11248), .A3(n14837), .ZN(n14836) );
  OR2_X1 U12398 ( .A1(n14040), .A2(n21172), .ZN(n11067) );
  AND2_X1 U12399 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .ZN(n11068) );
  NAND2_X1 U12400 ( .A1(n18070), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n18046) );
  INV_X1 U12401 ( .A(n18046), .ZN(n11136) );
  INV_X1 U12402 ( .A(n11138), .ZN(n20264) );
  NAND2_X1 U12403 ( .A1(n11136), .A2(n11134), .ZN(n11138) );
  AND2_X1 U12404 ( .A1(n11353), .A2(n12113), .ZN(n11069) );
  INV_X1 U12405 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11133) );
  INV_X1 U12406 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n11089) );
  INV_X1 U12407 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n11148) );
  INV_X1 U12408 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n11151) );
  INV_X1 U12409 ( .A(n16078), .ZN(n11310) );
  INV_X1 U12410 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n11090) );
  NAND2_X1 U12411 ( .A1(n11352), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11070) );
  NAND3_X2 U12412 ( .A1(n20095), .A2(n21232), .A3(n21235), .ZN(n21176) );
  OAI22_X2 U12413 ( .A1(n20075), .A2(n22152), .B1(n16178), .B2(n22150), .ZN(
        n21985) );
  OAI22_X2 U12414 ( .A1(n20082), .A2(n22152), .B1(n17101), .B2(n22150), .ZN(
        n22096) );
  OAI22_X2 U12415 ( .A1(n22147), .A2(n22152), .B1(n22146), .B2(n22150), .ZN(
        n22193) );
  AOI22_X2 U12416 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19689), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19690), .ZN(n19500) );
  NOR2_X1 U12417 ( .A1(n20098), .A2(n18192), .ZN(n18203) );
  NOR2_X2 U12418 ( .A1(n21206), .A2(n18755), .ZN(n19117) );
  AOI211_X2 U12419 ( .C1(n16910), .C2(n17744), .A(n19006), .B(n16904), .ZN(
        n18145) );
  OAI22_X2 U12420 ( .A1(n20084), .A2(n22152), .B1(n17118), .B2(n22150), .ZN(
        n22140) );
  CLKBUF_X1 U12421 ( .A(n22259), .Z(n11071) );
  NAND2_X1 U12422 ( .A1(n11076), .A2(n11907), .ZN(n16590) );
  NAND2_X1 U12423 ( .A1(n10960), .A2(n16860), .ZN(n11076) );
  OAI211_X2 U12424 ( .C1(n16860), .C2(n11078), .A(n11077), .B(n16586), .ZN(
        n16439) );
  OR2_X2 U12425 ( .A1(n10959), .A2(n11078), .ZN(n11077) );
  INV_X1 U12426 ( .A(n16587), .ZN(n11079) );
  XNOR2_X2 U12427 ( .A(n11080), .B(n12125), .ZN(n11767) );
  AND2_X2 U12428 ( .A1(n11313), .A2(n11081), .ZN(n12471) );
  AND3_X2 U12429 ( .A1(n11860), .A2(n11051), .A3(n11350), .ZN(n11855) );
  NAND4_X1 U12430 ( .A1(n11820), .A2(n11821), .A3(n11818), .A4(n11819), .ZN(
        n11084) );
  NAND3_X1 U12431 ( .A1(n11737), .A2(n11086), .A3(n11085), .ZN(n11747) );
  NAND2_X1 U12432 ( .A1(n11087), .A2(n11725), .ZN(n11748) );
  OR2_X1 U12433 ( .A1(n11736), .A2(n18669), .ZN(n11085) );
  NAND2_X1 U12434 ( .A1(n11357), .A2(n11720), .ZN(n11087) );
  NAND3_X1 U12435 ( .A1(n11093), .A2(n11092), .A3(n13475), .ZN(n11091) );
  NAND3_X1 U12436 ( .A1(n10986), .A2(P3_EAX_REG_20__SCAN_IN), .A3(
        P3_EAX_REG_22__SCAN_IN), .ZN(n11098) );
  NAND3_X1 U12437 ( .A1(n16862), .A2(n16861), .A3(n11102), .ZN(n11101) );
  NAND3_X1 U12438 ( .A1(n11105), .A2(n12093), .A3(n11103), .ZN(n11102) );
  MUX2_X1 U12439 ( .A(n12101), .B(n15478), .S(n11121), .Z(n11107) );
  NOR2_X2 U12440 ( .A1(n16408), .A2(n11111), .ZN(n16377) );
  NAND3_X1 U12441 ( .A1(n11787), .A2(n11351), .A3(n11786), .ZN(n11350) );
  NAND2_X2 U12442 ( .A1(n11404), .A2(n11403), .ZN(n11661) );
  NAND3_X1 U12443 ( .A1(n11118), .A2(n11116), .A3(n11115), .ZN(P2_U3015) );
  NAND2_X1 U12444 ( .A1(n16555), .A2(n11069), .ZN(n16462) );
  INV_X1 U12445 ( .A(n16462), .ZN(n12114) );
  NAND2_X1 U12446 ( .A1(n20500), .A2(n11128), .ZN(n11127) );
  NAND3_X1 U12447 ( .A1(n11144), .A2(n11040), .A3(n11145), .ZN(n13790) );
  NAND2_X1 U12448 ( .A1(n18562), .A2(n11381), .ZN(n18376) );
  NAND2_X1 U12449 ( .A1(n16376), .A2(n11156), .ZN(P2_U2986) );
  NAND2_X2 U12450 ( .A1(n11855), .A2(n11854), .ZN(n12100) );
  OR2_X2 U12451 ( .A1(n16419), .A2(n16421), .ZN(n11175) );
  AOI21_X1 U12452 ( .B1(n11170), .B2(n11167), .A(n11173), .ZN(n11166) );
  AND2_X2 U12453 ( .A1(n11172), .A2(n11170), .ZN(n16394) );
  AND2_X2 U12454 ( .A1(n15200), .A2(n11685), .ZN(n14388) );
  NAND3_X1 U12455 ( .A1(n13984), .A2(n13985), .A3(n11192), .ZN(n11191) );
  AOI22_X1 U12456 ( .A1(n17585), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11192) );
  INV_X1 U12457 ( .A(n20739), .ZN(n18134) );
  NAND2_X1 U12458 ( .A1(n14038), .A2(n20957), .ZN(n11196) );
  INV_X1 U12459 ( .A(n14038), .ZN(n11197) );
  NAND2_X1 U12460 ( .A1(n11194), .A2(n11193), .ZN(n20962) );
  NAND2_X1 U12461 ( .A1(n18051), .A2(n11196), .ZN(n11194) );
  NAND2_X1 U12462 ( .A1(n11195), .A2(n11196), .ZN(n17987) );
  INV_X1 U12463 ( .A(n11198), .ZN(n18050) );
  OR2_X1 U12464 ( .A1(n21068), .A2(n11203), .ZN(n21011) );
  NAND4_X1 U12465 ( .A1(n21044), .A2(n11208), .A3(n11207), .A4(n11206), .ZN(
        n11205) );
  OR2_X2 U12466 ( .A1(n16575), .A2(n16576), .ZN(n16796) );
  NAND2_X1 U12467 ( .A1(n11039), .A2(n10989), .ZN(n11338) );
  AOI21_X2 U12468 ( .B1(n16493), .B2(n16452), .A(n16451), .ZN(n16453) );
  AND2_X2 U12469 ( .A1(n11215), .A2(n12520), .ZN(n12729) );
  AND2_X2 U12470 ( .A1(n12518), .A2(n11215), .ZN(n12658) );
  AND2_X2 U12471 ( .A1(n15576), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11215) );
  NAND4_X4 U12472 ( .A1(n12612), .A2(n12611), .A3(n12609), .A4(n12610), .ZN(
        n12623) );
  NAND2_X1 U12473 ( .A1(n15515), .A2(n11223), .ZN(n16250) );
  NAND2_X1 U12474 ( .A1(n16216), .A2(n11237), .ZN(n14449) );
  AND2_X1 U12475 ( .A1(n16216), .A2(n16217), .ZN(n16206) );
  NAND2_X1 U12476 ( .A1(n16216), .A2(n11236), .ZN(n12238) );
  NAND2_X2 U12477 ( .A1(n11659), .A2(n11658), .ZN(n11680) );
  NAND2_X1 U12478 ( .A1(n12795), .A2(n11047), .ZN(n11256) );
  NAND2_X1 U12479 ( .A1(n12795), .A2(n12871), .ZN(n12878) );
  NOR2_X1 U12481 ( .A1(n15664), .A2(n15665), .ZN(n15648) );
  NOR2_X1 U12482 ( .A1(n15664), .A2(n11264), .ZN(n13779) );
  NAND2_X1 U12483 ( .A1(n13780), .A2(n11266), .ZN(n11265) );
  NOR2_X1 U12484 ( .A1(n11267), .A2(n15636), .ZN(n11266) );
  AND2_X2 U12485 ( .A1(n15724), .A2(n11269), .ZN(n15674) );
  INV_X1 U12486 ( .A(n12846), .ZN(n11277) );
  NOR2_X4 U12487 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14900) );
  NAND2_X2 U12488 ( .A1(n12819), .A2(n12846), .ZN(n14911) );
  INV_X1 U12489 ( .A(n11281), .ZN(n14046) );
  INV_X1 U12490 ( .A(n14051), .ZN(n17945) );
  NAND2_X1 U12491 ( .A1(n14012), .A2(n21015), .ZN(n14051) );
  OR2_X2 U12492 ( .A1(n14012), .A2(n21015), .ZN(n11281) );
  NAND2_X1 U12493 ( .A1(n11283), .A2(n20950), .ZN(n11282) );
  NAND2_X1 U12494 ( .A1(n13701), .A2(n11284), .ZN(n13712) );
  NOR2_X1 U12495 ( .A1(n19956), .A2(n11285), .ZN(n11284) );
  XNOR2_X1 U12496 ( .A(n11286), .B(n19956), .ZN(n21293) );
  NAND2_X1 U12497 ( .A1(n11287), .A2(n11021), .ZN(n17975) );
  NAND2_X1 U12498 ( .A1(n17840), .A2(n14009), .ZN(n17881) );
  NAND2_X1 U12499 ( .A1(n11297), .A2(n11295), .ZN(n19965) );
  NAND2_X1 U12500 ( .A1(n13731), .A2(n13730), .ZN(n15424) );
  NOR2_X1 U12501 ( .A1(n11299), .A2(n15425), .ZN(n11298) );
  INV_X1 U12502 ( .A(n13730), .ZN(n11299) );
  NAND2_X1 U12503 ( .A1(n13758), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11308) );
  NAND2_X1 U12504 ( .A1(n11307), .A2(n11309), .ZN(n13777) );
  NAND3_X1 U12505 ( .A1(n13759), .A2(n11046), .A3(n11308), .ZN(n11307) );
  NAND3_X1 U12506 ( .A1(n13757), .A2(n11311), .A3(n15956), .ZN(n13756) );
  NAND3_X1 U12507 ( .A1(n20795), .A2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n20789) );
  OR2_X1 U12508 ( .A1(n11313), .A2(n14649), .ZN(n11312) );
  INV_X1 U12509 ( .A(n16777), .ZN(n11314) );
  NAND2_X1 U12510 ( .A1(n11314), .A2(n11315), .ZN(n16750) );
  NAND2_X1 U12511 ( .A1(n16848), .A2(n11321), .ZN(n16793) );
  INV_X1 U12512 ( .A(n11323), .ZN(n16839) );
  NAND2_X1 U12513 ( .A1(n16691), .A2(n11327), .ZN(n16332) );
  INV_X1 U12514 ( .A(n16410), .ZN(n11333) );
  NAND3_X1 U12515 ( .A1(n11334), .A2(n14411), .A3(n12100), .ZN(n11880) );
  NAND2_X1 U12516 ( .A1(n10989), .A2(n11037), .ZN(n11823) );
  NAND2_X2 U12517 ( .A1(n11341), .A2(n11339), .ZN(n16430) );
  NAND2_X1 U12518 ( .A1(n11999), .A2(n16365), .ZN(n11348) );
  AND2_X2 U12519 ( .A1(n11344), .A2(n11038), .ZN(n14443) );
  NAND2_X1 U12520 ( .A1(n11716), .A2(n11715), .ZN(n11349) );
  NAND3_X1 U12521 ( .A1(n11664), .A2(n11663), .A3(n11689), .ZN(n11679) );
  NAND4_X1 U12522 ( .A1(n11663), .A2(n11664), .A3(n11689), .A4(n19686), .ZN(
        n12054) );
  AND2_X1 U12523 ( .A1(n16377), .A2(n11352), .ZN(n14467) );
  NAND2_X1 U12524 ( .A1(n16819), .A2(n12110), .ZN(n16555) );
  AND2_X2 U12525 ( .A1(n16579), .A2(n16722), .ZN(n16487) );
  NAND2_X1 U12526 ( .A1(n12098), .A2(n11104), .ZN(n12094) );
  INV_X1 U12527 ( .A(n12056), .ZN(n12288) );
  NAND2_X1 U12528 ( .A1(n12259), .A2(n11686), .ZN(n11642) );
  AND2_X1 U12529 ( .A1(n11355), .A2(n15200), .ZN(n11354) );
  NAND2_X1 U12530 ( .A1(n12056), .A2(n12057), .ZN(n11355) );
  INV_X1 U12531 ( .A(n12065), .ZN(n11356) );
  NAND2_X1 U12532 ( .A1(n11717), .A2(n11718), .ZN(n11357) );
  INV_X1 U12533 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11358) );
  AND3_X2 U12534 ( .A1(n15176), .A2(n11454), .A3(n11358), .ZN(n11396) );
  INV_X1 U12535 ( .A(n14055), .ZN(n15047) );
  AOI21_X1 U12536 ( .B1(n15505), .B2(n11065), .A(n11001), .ZN(n16240) );
  INV_X1 U12537 ( .A(n11363), .ZN(n15268) );
  NAND2_X1 U12538 ( .A1(n14918), .A2(n14883), .ZN(n14882) );
  INV_X1 U12539 ( .A(n15116), .ZN(n12652) );
  NAND2_X1 U12540 ( .A1(n12717), .A2(n12716), .ZN(n12725) );
  AND2_X1 U12541 ( .A1(n19686), .A2(n11682), .ZN(n11690) );
  NAND2_X1 U12542 ( .A1(n12650), .A2(n15116), .ZN(n12717) );
  INV_X1 U12543 ( .A(n12510), .ZN(n12511) );
  NAND2_X1 U12545 ( .A1(n16487), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16759) );
  AND2_X1 U12546 ( .A1(n11760), .A2(n11759), .ZN(n11764) );
  NAND2_X1 U12547 ( .A1(n12652), .A2(n12651), .ZN(n21783) );
  INV_X1 U12548 ( .A(n12651), .ZN(n12650) );
  NAND2_X2 U12549 ( .A1(n13682), .A2(n13681), .ZN(n13684) );
  OR2_X1 U12550 ( .A1(n14760), .A2(n14759), .ZN(n14762) );
  OR2_X1 U12551 ( .A1(n14437), .A2(n18609), .ZN(n14438) );
  NAND2_X2 U12552 ( .A1(n13672), .A2(n13671), .ZN(n13680) );
  NAND2_X1 U12553 ( .A1(n13660), .A2(n13360), .ZN(n13377) );
  AOI211_X2 U12554 ( .C1(n20000), .C2(n15922), .A(n15921), .B(n15920), .ZN(
        n15923) );
  OR2_X2 U12555 ( .A1(n16228), .A2(n16231), .ZN(n16229) );
  NOR2_X2 U12556 ( .A1(n15504), .A2(n15506), .ZN(n15505) );
  AOI22_X1 U12557 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10974), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11427) );
  INV_X1 U12558 ( .A(n14882), .ZN(n12143) );
  NAND2_X1 U12559 ( .A1(n16223), .A2(n16222), .ZN(n16221) );
  AOI211_X2 U12560 ( .C1(n18541), .C2(n18603), .A(n12507), .B(n12506), .ZN(
        n12508) );
  OAI21_X2 U12561 ( .B1(n14911), .B2(n13732), .A(n13665), .ZN(n14938) );
  AND2_X1 U12562 ( .A1(n19946), .A2(n14948), .ZN(n19942) );
  NAND2_X1 U12563 ( .A1(n19946), .A2(n15597), .ZN(n15837) );
  INV_X1 U12564 ( .A(n20020), .ZN(n21578) );
  NOR2_X2 U12565 ( .A1(n16965), .A2(n22310), .ZN(n20020) );
  NAND2_X1 U12566 ( .A1(n14760), .A2(n14759), .ZN(n14761) );
  INV_X1 U12567 ( .A(n18652), .ZN(n14062) );
  AND2_X1 U12568 ( .A1(n14472), .A2(n14471), .ZN(n11364) );
  NOR2_X1 U12569 ( .A1(n12108), .A2(n16818), .ZN(n11366) );
  NOR2_X1 U12570 ( .A1(n16324), .A2(n16314), .ZN(n11367) );
  AND3_X1 U12571 ( .A1(n13512), .A2(n13518), .A3(n13517), .ZN(n11368) );
  AND4_X1 U12572 ( .A1(n16133), .A2(n21373), .A3(n15964), .A4(n21343), .ZN(
        n11369) );
  INV_X1 U12573 ( .A(n12830), .ZN(n13232) );
  NOR2_X1 U12574 ( .A1(n14948), .A2(n21917), .ZN(n12830) );
  INV_X1 U12575 ( .A(n16704), .ZN(n12113) );
  OR4_X1 U12576 ( .A1(n16600), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14462), .A4(n14461), .ZN(n11370) );
  NOR2_X1 U12577 ( .A1(n16352), .A2(n14402), .ZN(n11371) );
  OR2_X1 U12578 ( .A1(n12623), .A2(n13633), .ZN(n11372) );
  OR2_X1 U12579 ( .A1(n18771), .A2(n19054), .ZN(n19005) );
  NOR2_X1 U12580 ( .A1(n13784), .A2(n16581), .ZN(n11373) );
  OR2_X1 U12581 ( .A1(n13849), .A2(n11582), .ZN(n11374) );
  AND2_X1 U12582 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11375) );
  INV_X1 U12583 ( .A(n11699), .ZN(n12064) );
  OR2_X1 U12584 ( .A1(n13849), .A2(n11583), .ZN(n11378) );
  NAND2_X1 U12585 ( .A1(n11035), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11379) );
  AND2_X1 U12586 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n11380) );
  OR2_X1 U12587 ( .A1(n14483), .A2(n16562), .ZN(n11381) );
  CLKBUF_X3 U12588 ( .A(n17510), .Z(n17497) );
  AND2_X1 U12589 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n10976), .ZN(
        n11382) );
  AND2_X1 U12590 ( .A1(n12054), .A2(n11683), .ZN(n11383) );
  INV_X1 U12591 ( .A(n11680), .ZN(n12069) );
  NOR2_X1 U12592 ( .A1(n18135), .A2(n10977), .ZN(n17925) );
  INV_X1 U12593 ( .A(n17925), .ZN(n17977) );
  AND4_X1 U12594 ( .A1(n11507), .A2(n11506), .A3(n11505), .A4(n11504), .ZN(
        n11384) );
  OR2_X1 U12595 ( .A1(n17214), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n18582) );
  INV_X1 U12596 ( .A(n18582), .ZN(n18382) );
  OR2_X1 U12597 ( .A1(n12364), .A2(n12363), .ZN(n11385) );
  INV_X1 U12598 ( .A(n11682), .ZN(n11671) );
  BUF_X4 U12599 ( .A(n13981), .Z(n17503) );
  AND2_X1 U12600 ( .A1(n15821), .A2(n15818), .ZN(n11386) );
  INV_X1 U12601 ( .A(n12275), .ZN(n11706) );
  AND3_X1 U12602 ( .A1(n17246), .A2(n16566), .A3(n16568), .ZN(n16522) );
  INV_X1 U12603 ( .A(n15505), .ZN(n15558) );
  INV_X1 U12604 ( .A(n11746), .ZN(n11756) );
  AND3_X1 U12605 ( .A1(n12561), .A2(n12560), .A3(n12559), .ZN(n11387) );
  AND4_X1 U12606 ( .A1(n12567), .A2(n12566), .A3(n12565), .A4(n12564), .ZN(
        n11388) );
  INV_X1 U12607 ( .A(n14872), .ZN(n14860) );
  NAND2_X1 U12608 ( .A1(n11831), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11759) );
  NAND2_X1 U12609 ( .A1(n11833), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11777) );
  AND2_X1 U12610 ( .A1(n11645), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11390) );
  NAND2_X1 U12611 ( .A1(n12250), .A2(n11245), .ZN(n11641) );
  AOI22_X1 U12612 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10974), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11394) );
  NAND2_X1 U12613 ( .A1(n19247), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11785) );
  AOI21_X1 U12614 ( .B1(n11520), .B2(n11519), .A(n11518), .ZN(n12022) );
  AND4_X1 U12615 ( .A1(n11662), .A2(n12069), .A3(n11661), .A4(n11668), .ZN(
        n11664) );
  INV_X1 U12616 ( .A(n11405), .ZN(n11410) );
  NAND2_X1 U12617 ( .A1(n12308), .A2(n19621), .ZN(n11822) );
  AOI22_X1 U12618 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10974), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11432) );
  OR2_X1 U12619 ( .A1(n12792), .A2(n12791), .ZN(n13706) );
  OR2_X1 U12620 ( .A1(n12665), .A2(n12664), .ZN(n13667) );
  NAND2_X1 U12621 ( .A1(n12666), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12667) );
  OR2_X1 U12622 ( .A1(n11379), .A2(n12715), .ZN(n12716) );
  AOI22_X1 U12623 ( .A1(n12761), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12774), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12540) );
  OAI211_X1 U12624 ( .C1(n13314), .C2(n12687), .A(n12710), .B(n12686), .ZN(
        n12747) );
  NAND2_X1 U12625 ( .A1(n11691), .A2(n11455), .ZN(n11456) );
  INV_X1 U12626 ( .A(n11927), .ZN(n11577) );
  INV_X1 U12627 ( .A(n14060), .ZN(n14061) );
  OR2_X1 U12628 ( .A1(n15818), .A2(n15817), .ZN(n13063) );
  AND2_X1 U12629 ( .A1(n12807), .A2(n12806), .ZN(n12877) );
  INV_X1 U12630 ( .A(n13093), .ZN(n13094) );
  INV_X1 U12631 ( .A(n12972), .ZN(n12973) );
  AND2_X1 U12632 ( .A1(n13571), .A2(n13570), .ZN(n15523) );
  OR2_X1 U12633 ( .A1(n13606), .A2(n14687), .ZN(n13595) );
  INV_X1 U12634 ( .A(n13732), .ZN(n13720) );
  INV_X1 U12635 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n16161) );
  INV_X1 U12636 ( .A(n11553), .ZN(n11902) );
  AND2_X1 U12637 ( .A1(n14087), .A2(n14086), .ZN(n14088) );
  AND2_X2 U12638 ( .A1(n11358), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11412) );
  INV_X1 U12639 ( .A(n11772), .ZN(n11755) );
  NAND2_X1 U12640 ( .A1(n11443), .A2(n11613), .ZN(n11450) );
  INV_X1 U12641 ( .A(n21559), .ZN(n21533) );
  NAND2_X1 U12642 ( .A1(n14687), .A2(n13543), .ZN(n13612) );
  AND2_X1 U12643 ( .A1(n21917), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13303) );
  AND2_X1 U12644 ( .A1(n13159), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13160) );
  NAND2_X1 U12645 ( .A1(n13754), .A2(n11369), .ZN(n13755) );
  NAND2_X1 U12646 ( .A1(n12973), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12981) );
  NAND2_X1 U12647 ( .A1(n12917), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12933) );
  INV_X1 U12648 ( .A(n14975), .ZN(n12870) );
  OR2_X1 U12649 ( .A1(n13735), .A2(n21361), .ZN(n20005) );
  AND2_X1 U12650 ( .A1(n13574), .A2(n13573), .ZN(n15534) );
  NAND2_X1 U12651 ( .A1(n12754), .A2(n12753), .ZN(n15115) );
  AND2_X1 U12652 ( .A1(n12026), .A2(n12025), .ZN(n12046) );
  INV_X1 U12653 ( .A(n16204), .ZN(n14340) );
  AND2_X1 U12654 ( .A1(n14137), .A2(n15338), .ZN(n14138) );
  INV_X1 U12655 ( .A(n12250), .ZN(n12253) );
  OR2_X1 U12656 ( .A1(n16392), .A2(n16400), .ZN(n11996) );
  AND2_X1 U12657 ( .A1(n12481), .A2(n12480), .ZN(n16340) );
  AND3_X1 U12658 ( .A1(n12455), .A2(n12454), .A3(n12453), .ZN(n18372) );
  OR2_X1 U12659 ( .A1(n13882), .A2(n20762), .ZN(n17345) );
  CLKBUF_X3 U12660 ( .A(n17361), .Z(n17722) );
  INV_X1 U12661 ( .A(n20906), .ZN(n21111) );
  CLKBUF_X3 U12662 ( .A(n13986), .Z(n17723) );
  INV_X1 U12663 ( .A(n13869), .ZN(n13873) );
  INV_X1 U12664 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21210) );
  INV_X1 U12665 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n21502) );
  OAI21_X1 U12666 ( .B1(n16972), .B2(n13528), .A(n14657), .ZN(n13623) );
  NAND2_X1 U12667 ( .A1(n14719), .A2(n12623), .ZN(n15096) );
  OR2_X2 U12668 ( .A1(n15433), .A2(n15520), .ZN(n15529) );
  NAND2_X1 U12669 ( .A1(n13095), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13127) );
  OR2_X1 U12670 ( .A1(n15819), .A2(n15835), .ZN(n15817) );
  INV_X1 U12671 ( .A(n16130), .ZN(n21347) );
  AND2_X1 U12672 ( .A1(n14857), .A2(n15620), .ZN(n14874) );
  AND2_X1 U12673 ( .A1(n21821), .A2(n21820), .ZN(n21854) );
  NOR2_X1 U12674 ( .A1(n21839), .A2(n21825), .ZN(n21886) );
  OR2_X1 U12675 ( .A1(n21769), .A2(n15138), .ZN(n21873) );
  NAND2_X1 U12676 ( .A1(n21870), .A2(n21808), .ZN(n21910) );
  INV_X1 U12677 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21933) );
  INV_X1 U12678 ( .A(n21808), .ZN(n15129) );
  OR2_X1 U12679 ( .A1(n12046), .A2(n12045), .ZN(n18630) );
  OAI22_X1 U12680 ( .A1(n14469), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n18669), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n15031) );
  AND3_X1 U12681 ( .A1(n12317), .A2(n12316), .A3(n12315), .ZN(n15375) );
  INV_X1 U12682 ( .A(n18534), .ZN(n18552) );
  AND2_X1 U12683 ( .A1(n12201), .A2(n12200), .ZN(n15514) );
  BUF_X2 U12684 ( .A(n11767), .Z(n14055) );
  INV_X1 U12685 ( .A(n16212), .ZN(n16213) );
  AND2_X1 U12686 ( .A1(n19508), .A2(n14403), .ZN(n14647) );
  INV_X1 U12687 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16569) );
  OR3_X1 U12688 ( .A1(n16667), .A2(n11987), .A3(n16655), .ZN(n16611) );
  BUF_X1 U12689 ( .A(n16555), .Z(n16579) );
  NAND2_X1 U12690 ( .A1(n12103), .A2(n12102), .ZN(n12110) );
  AND2_X1 U12691 ( .A1(n14640), .A2(n14639), .ZN(n18611) );
  NAND2_X1 U12692 ( .A1(n19453), .A2(n19452), .ZN(n19308) );
  NAND2_X1 U12693 ( .A1(n19453), .A2(n19559), .ZN(n19256) );
  NOR2_X1 U12694 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19295) );
  NAND2_X1 U12695 ( .A1(n19330), .A2(n19452), .ZN(n19220) );
  INV_X1 U12696 ( .A(n19295), .ZN(n19326) );
  AOI211_X1 U12697 ( .C1(n17561), .C2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n13436), .B(n13435), .ZN(n13437) );
  INV_X1 U12698 ( .A(n20964), .ZN(n17816) );
  INV_X1 U12699 ( .A(n21067), .ZN(n21110) );
  NOR2_X1 U12700 ( .A1(n14019), .A2(n13978), .ZN(n14016) );
  NOR2_X1 U12701 ( .A1(n13409), .A2(n13408), .ZN(n18919) );
  INV_X1 U12702 ( .A(n21255), .ZN(n14657) );
  OR2_X1 U12703 ( .A1(n14658), .A2(n13527), .ZN(n21255) );
  OAI21_X1 U12704 ( .B1(n16022), .B2(n21562), .A(n13645), .ZN(n13646) );
  NOR2_X1 U12705 ( .A1(n21482), .A2(n21459), .ZN(n15756) );
  INV_X1 U12706 ( .A(n21562), .ZN(n21469) );
  AND2_X1 U12707 ( .A1(n15124), .A2(n15092), .ZN(n13638) );
  NAND2_X1 U12708 ( .A1(n12873), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12879) );
  NOR2_X1 U12709 ( .A1(n13623), .A2(n21390), .ZN(n21411) );
  INV_X1 U12710 ( .A(n15837), .ZN(n19941) );
  AND2_X1 U12711 ( .A1(n13078), .A2(n13077), .ZN(n15755) );
  INV_X1 U12712 ( .A(n22310), .ZN(n15620) );
  NAND2_X1 U12713 ( .A1(n13060), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13059) );
  INV_X1 U12714 ( .A(n19983), .ZN(n20015) );
  AND2_X1 U12715 ( .A1(n19983), .A2(n13657), .ZN(n20000) );
  INV_X1 U12716 ( .A(n21378), .ZN(n21390) );
  NAND2_X1 U12717 ( .A1(n14870), .A2(n21402), .ZN(n21337) );
  INV_X1 U12718 ( .A(n16031), .ZN(n21334) );
  AND2_X1 U12719 ( .A1(n14874), .A2(n14869), .ZN(n21265) );
  INV_X1 U12720 ( .A(n14715), .ZN(n21821) );
  NOR2_X1 U12721 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15582) );
  AND2_X1 U12722 ( .A1(n21809), .A2(n21862), .ZN(n22214) );
  AND2_X1 U12723 ( .A1(n21809), .A2(n21791), .ZN(n22226) );
  AND2_X1 U12724 ( .A1(n21809), .A2(n21808), .ZN(n22233) );
  INV_X1 U12725 ( .A(n22243), .ZN(n22166) );
  AND2_X1 U12726 ( .A1(n21851), .A2(n21836), .ZN(n22253) );
  INV_X1 U12727 ( .A(n22257), .ZN(n22260) );
  INV_X1 U12728 ( .A(n21893), .ZN(n21862) );
  INV_X1 U12729 ( .A(n21873), .ZN(n21870) );
  NOR2_X1 U12730 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15122), .ZN(n22145) );
  INV_X1 U12731 ( .A(n21910), .ZN(n22283) );
  INV_X1 U12732 ( .A(n22295), .ZN(n22301) );
  INV_X1 U12733 ( .A(n22135), .ZN(n22138) );
  NOR2_X2 U12734 ( .A1(n21921), .A2(n15129), .ZN(n22207) );
  AND2_X1 U12735 ( .A1(n18248), .A2(n13859), .ZN(n18538) );
  OR3_X1 U12736 ( .A1(n18248), .A2(n13854), .A3(n13853), .ZN(n18551) );
  INV_X1 U12737 ( .A(n19349), .ZN(n19396) );
  OR2_X1 U12738 ( .A1(n19672), .A2(n14647), .ZN(n19175) );
  INV_X1 U12739 ( .A(n14622), .ZN(n14606) );
  AND2_X1 U12740 ( .A1(n18373), .A2(n11043), .ZN(n19159) );
  INV_X1 U12741 ( .A(n18609), .ZN(n16864) );
  INV_X1 U12742 ( .A(n16871), .ZN(n18601) );
  AND2_X1 U12743 ( .A1(n12279), .A2(n12243), .ZN(n18603) );
  INV_X1 U12744 ( .A(n19453), .ZN(n19330) );
  OAI21_X1 U12745 ( .B1(n15353), .B2(n15352), .A(n15351), .ZN(n19792) );
  NOR2_X1 U12746 ( .A1(n19195), .A2(n19308), .ZN(n19794) );
  INV_X1 U12747 ( .A(n19770), .ZN(n19653) );
  OAI21_X1 U12748 ( .B1(n19287), .B2(n19286), .A(n19285), .ZN(n19761) );
  INV_X1 U12749 ( .A(n19650), .ZN(n19760) );
  NOR2_X1 U12750 ( .A1(n19256), .A2(n19307), .ZN(n19749) );
  OAI21_X1 U12751 ( .B1(n19250), .B2(n19249), .A(n19248), .ZN(n19735) );
  NOR2_X2 U12752 ( .A1(n19220), .A2(n19195), .ZN(n19734) );
  OAI21_X1 U12753 ( .B1(n19238), .B2(n19237), .A(n19236), .ZN(n19721) );
  NOR2_X1 U12754 ( .A1(n19220), .A2(n19290), .ZN(n19720) );
  NOR2_X1 U12755 ( .A1(n19220), .A2(n19276), .ZN(n19630) );
  INV_X1 U12756 ( .A(n19574), .ZN(n19702) );
  INV_X1 U12757 ( .A(n19644), .ZN(n19666) );
  INV_X1 U12758 ( .A(n15392), .ZN(n19328) );
  AND2_X1 U12759 ( .A1(n18655), .A2(n18654), .ZN(n18672) );
  OAI21_X1 U12760 ( .B1(n11054), .B2(n20312), .A(n10967), .ZN(n20398) );
  AND2_X1 U12761 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17696), .ZN(n17711) );
  NOR2_X1 U12762 ( .A1(n13429), .A2(n13428), .ZN(n19057) );
  NOR3_X1 U12763 ( .A1(n21619), .A2(n21192), .A3(n21244), .ZN(n20561) );
  INV_X1 U12764 ( .A(n13497), .ZN(n20103) );
  AOI21_X1 U12765 ( .B1(n20097), .B2(n20095), .A(n17749), .ZN(n18111) );
  NOR2_X1 U12766 ( .A1(n21247), .A2(n19007), .ZN(n18081) );
  NOR2_X1 U12767 ( .A1(n21176), .A2(n20519), .ZN(n14052) );
  INV_X1 U12768 ( .A(n21144), .ZN(n21166) );
  INV_X1 U12769 ( .A(n20888), .ZN(n21012) );
  INV_X1 U12770 ( .A(n21074), .ZN(n21062) );
  AND2_X1 U12771 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n21621), .ZN(n18230) );
  INV_X1 U12772 ( .A(n13646), .ZN(n13647) );
  NOR2_X1 U12773 ( .A1(n21313), .A2(n21509), .ZN(n21529) );
  OR2_X1 U12774 ( .A1(n21411), .A2(n15101), .ZN(n21565) );
  AND2_X1 U12775 ( .A1(n21571), .A2(n15094), .ZN(n21448) );
  INV_X1 U12776 ( .A(n15888), .ZN(n15885) );
  INV_X1 U12777 ( .A(n19857), .ZN(n19877) );
  NAND2_X2 U12778 ( .A1(n14804), .A2(n14803), .ZN(n21766) );
  INV_X1 U12779 ( .A(n20000), .ZN(n20025) );
  OR2_X1 U12780 ( .A1(n20020), .A2(n13655), .ZN(n19983) );
  INV_X1 U12781 ( .A(n20021), .ZN(n19957) );
  INV_X1 U12782 ( .A(n21406), .ZN(n21327) );
  NAND2_X1 U12783 ( .A1(n21809), .A2(n21782), .ZN(n22219) );
  INV_X1 U12784 ( .A(n21807), .ZN(n22230) );
  OR2_X1 U12785 ( .A1(n21831), .A2(n21836), .ZN(n22245) );
  NAND2_X1 U12786 ( .A1(n21851), .A2(n21850), .ZN(n22257) );
  NAND2_X1 U12787 ( .A1(n21870), .A2(n21862), .ZN(n22270) );
  NAND2_X1 U12788 ( .A1(n21870), .A2(n21782), .ZN(n22279) );
  NAND2_X1 U12789 ( .A1(n21870), .A2(n21791), .ZN(n22273) );
  INV_X1 U12790 ( .A(n22101), .ZN(n22093) );
  INV_X1 U12791 ( .A(n22200), .ZN(n22190) );
  NAND2_X1 U12792 ( .A1(n21914), .A2(n21782), .ZN(n22295) );
  NAND2_X1 U12793 ( .A1(n21914), .A2(n21791), .ZN(n22305) );
  INV_X1 U12794 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n18669) );
  INV_X1 U12795 ( .A(n18539), .ZN(n18567) );
  INV_X1 U12796 ( .A(n16267), .ZN(n16209) );
  NAND2_X1 U12797 ( .A1(n14762), .A2(n14761), .ZN(n19453) );
  AND2_X1 U12798 ( .A1(n14407), .A2(n14406), .ZN(n14408) );
  NAND2_X1 U12799 ( .A1(n12288), .A2(n19508), .ZN(n19677) );
  AND2_X1 U12800 ( .A1(n14386), .A2(n18683), .ZN(n19508) );
  INV_X1 U12801 ( .A(n19175), .ZN(n19619) );
  INV_X1 U12802 ( .A(n17294), .ZN(n17323) );
  CLKBUF_X1 U12803 ( .A(n14568), .Z(n14610) );
  INV_X1 U12804 ( .A(n17256), .ZN(n17224) );
  INV_X1 U12805 ( .A(n17216), .ZN(n17261) );
  NAND2_X1 U12806 ( .A1(n12279), .A2(n18624), .ZN(n18609) );
  INV_X1 U12807 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19294) );
  INV_X1 U12808 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19669) );
  AOI21_X1 U12809 ( .B1(n15347), .B2(n15348), .A(n19683), .ZN(n19798) );
  INV_X1 U12810 ( .A(n19794), .ZN(n19785) );
  OAI21_X1 U12811 ( .B1(n19315), .B2(n19332), .A(n19314), .ZN(n19778) );
  NAND2_X1 U12812 ( .A1(n19278), .A2(n19277), .ZN(n19770) );
  INV_X1 U12813 ( .A(n19749), .ZN(n19758) );
  INV_X1 U12814 ( .A(n19645), .ZN(n19752) );
  INV_X1 U12815 ( .A(n19742), .ZN(n19739) );
  AND2_X1 U12816 ( .A1(n15214), .A2(n15213), .ZN(n19732) );
  AOI211_X2 U12817 ( .C1(n19235), .C2(n19237), .A(n19683), .B(n19234), .ZN(
        n19725) );
  INV_X1 U12818 ( .A(n19720), .ZN(n19633) );
  INV_X1 U12819 ( .A(n19630), .ZN(n19718) );
  OR2_X1 U12820 ( .A1(n19198), .A2(n19307), .ZN(n19574) );
  OR2_X1 U12821 ( .A1(n19198), .A2(n19276), .ZN(n19569) );
  INV_X1 U12822 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n21655) );
  NOR2_X1 U12823 ( .A1(n21187), .A2(n20104), .ZN(n16913) );
  NAND2_X1 U12824 ( .A1(n13519), .A2(n11368), .ZN(n13520) );
  INV_X1 U12825 ( .A(n20547), .ZN(n20525) );
  INV_X1 U12826 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20235) );
  INV_X1 U12827 ( .A(n17640), .ZN(n17644) );
  INV_X1 U12828 ( .A(n17754), .ZN(n20593) );
  NOR2_X1 U12829 ( .A1(n13903), .A2(n13902), .ZN(n20597) );
  INV_X1 U12830 ( .A(n18192), .ZN(n18191) );
  NAND2_X1 U12831 ( .A1(n20103), .A2(n20561), .ZN(n20139) );
  NAND2_X1 U12832 ( .A1(n17754), .A2(n18081), .ZN(n18055) );
  NOR2_X1 U12833 ( .A1(n11024), .A2(n14052), .ZN(n14053) );
  NAND2_X1 U12834 ( .A1(n21151), .A2(n20922), .ZN(n21181) );
  INV_X1 U12835 ( .A(n21151), .ZN(n21080) );
  INV_X1 U12836 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19049) );
  INV_X1 U12837 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18876) );
  INV_X1 U12838 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n21232) );
  INV_X1 U12839 ( .A(n18235), .ZN(n21621) );
  OAI211_X1 U12840 ( .C1(n21578), .C2(n16074), .A(n11377), .B(n13783), .ZN(
        P1_U2970) );
  OR2_X1 U12841 ( .A1(n13521), .A2(n13520), .ZN(P3_U2640) );
  OAI21_X1 U12842 ( .B1(n14054), .B2(n21137), .A(n14053), .ZN(P3_U2834) );
  AND2_X4 U12843 ( .A1(n11412), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14371) );
  INV_X4 U12844 ( .A(n11419), .ZN(n11652) );
  AOI22_X1 U12845 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11651), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11393) );
  AND2_X4 U12846 ( .A1(n15321), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11645) );
  AOI21_X1 U12847 ( .B1(n14373), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n11390), .ZN(n11392) );
  INV_X1 U12848 ( .A(n16881), .ZN(n15322) );
  AOI22_X1 U12849 ( .A1(n15319), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n14200), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11391) );
  NAND4_X1 U12850 ( .A1(n11394), .A2(n11393), .A3(n11392), .A4(n11391), .ZN(
        n11395) );
  NAND2_X1 U12851 ( .A1(n11395), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11404) );
  AOI22_X1 U12852 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10975), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U12853 ( .A1(n11633), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11400) );
  AOI22_X1 U12854 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11651), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11399) );
  AOI22_X1 U12855 ( .A1(n15319), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14200), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11398) );
  NAND4_X1 U12856 ( .A1(n11401), .A2(n11400), .A3(n11399), .A4(n11398), .ZN(
        n11402) );
  NAND2_X1 U12857 ( .A1(n11402), .A2(n11613), .ZN(n11403) );
  NAND2_X1 U12858 ( .A1(n19400), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n13847) );
  AND2_X2 U12859 ( .A1(n15319), .A2(n11613), .ZN(n16892) );
  AND2_X2 U12860 ( .A1(n14200), .A2(n11613), .ZN(n14232) );
  AOI22_X1 U12861 ( .A1(n16892), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14232), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11405) );
  AND2_X2 U12862 ( .A1(n14371), .A2(n11613), .ZN(n14231) );
  AND2_X1 U12863 ( .A1(n14370), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11788) );
  AOI22_X1 U12864 ( .A1(n14231), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11408) );
  NAND3_X1 U12865 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12050) );
  NAND2_X1 U12866 ( .A1(n12385), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n11407) );
  AND2_X2 U12867 ( .A1(n11645), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11481) );
  AOI22_X1 U12868 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11481), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11406) );
  NAND3_X1 U12869 ( .A1(n11408), .A2(n11407), .A3(n11406), .ZN(n11409) );
  NOR2_X1 U12870 ( .A1(n11410), .A2(n11409), .ZN(n11426) );
  AND2_X2 U12871 ( .A1(n11411), .A2(n14198), .ZN(n14223) );
  AOI22_X1 U12872 ( .A1(n14223), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n14222), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11418) );
  NAND2_X1 U12873 ( .A1(n14172), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n11417) );
  AND2_X2 U12874 ( .A1(n14198), .A2(n11413), .ZN(n14224) );
  AOI22_X1 U12875 ( .A1(n14224), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14225), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11416) );
  AND2_X2 U12876 ( .A1(n10974), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11480) );
  NAND2_X1 U12877 ( .A1(n11480), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11415) );
  NAND4_X1 U12878 ( .A1(n11418), .A2(n11417), .A3(n11416), .A4(n11415), .ZN(
        n11424) );
  INV_X1 U12879 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11422) );
  NAND2_X1 U12880 ( .A1(n14215), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n11421) );
  AND2_X2 U12881 ( .A1(n15319), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14216) );
  NAND2_X1 U12882 ( .A1(n14216), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11420) );
  OAI211_X1 U12883 ( .C1(n11422), .C2(n14219), .A(n11421), .B(n11420), .ZN(
        n11423) );
  NOR2_X1 U12884 ( .A1(n11424), .A2(n11423), .ZN(n11425) );
  INV_X1 U12885 ( .A(n12298), .ZN(n11804) );
  AOI22_X1 U12887 ( .A1(n15319), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14360), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11428) );
  AOI22_X1 U12888 ( .A1(n14373), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11430) );
  AOI22_X1 U12889 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11651), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11429) );
  NAND3_X1 U12890 ( .A1(n11430), .A2(n11429), .A3(n11613), .ZN(n11437) );
  AOI22_X1 U12891 ( .A1(n11633), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11431) );
  AOI22_X1 U12892 ( .A1(n15319), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n14360), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11434) );
  AOI22_X1 U12893 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11651), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11433) );
  NAND3_X1 U12894 ( .A1(n11434), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n11433), .ZN(n11435) );
  AOI22_X1 U12895 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11396), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11442) );
  AOI22_X1 U12896 ( .A1(n11633), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11441) );
  AOI22_X1 U12897 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11651), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11440) );
  AOI22_X1 U12898 ( .A1(n15319), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n14200), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11439) );
  NAND4_X1 U12899 ( .A1(n11442), .A2(n11441), .A3(n11440), .A4(n11439), .ZN(
        n11443) );
  AOI22_X1 U12900 ( .A1(n15319), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n14200), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11447) );
  AOI22_X1 U12901 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11396), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11446) );
  AOI22_X1 U12902 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11651), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11445) );
  AOI22_X1 U12903 ( .A1(n11633), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11444) );
  NAND4_X1 U12904 ( .A1(n11447), .A2(n11446), .A3(n11445), .A4(n11444), .ZN(
        n11448) );
  NAND2_X1 U12905 ( .A1(n11448), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11449) );
  NAND2_X2 U12906 ( .A1(n11450), .A2(n11449), .ZN(n11681) );
  NAND2_X2 U12907 ( .A1(n11671), .A2(n11681), .ZN(n11691) );
  XNOR2_X1 U12908 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12033) );
  NAND2_X1 U12909 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19263), .ZN(
        n12007) );
  INV_X1 U12910 ( .A(n12007), .ZN(n11451) );
  NAND2_X1 U12911 ( .A1(n12033), .A2(n11451), .ZN(n11453) );
  NAND2_X1 U12912 ( .A1(n19294), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11452) );
  NAND2_X1 U12913 ( .A1(n11453), .A2(n11452), .ZN(n11474) );
  XNOR2_X1 U12914 ( .A(n11454), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11472) );
  XNOR2_X1 U12915 ( .A(n11474), .B(n11472), .ZN(n12042) );
  INV_X1 U12916 ( .A(n12042), .ZN(n11455) );
  AOI22_X1 U12917 ( .A1(n14172), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14215), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11464) );
  AOI22_X1 U12918 ( .A1(n11480), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n16892), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11463) );
  INV_X1 U12919 ( .A(n14219), .ZN(n14184) );
  AOI22_X1 U12920 ( .A1(n14184), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11481), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11462) );
  AOI22_X1 U12921 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14232), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11461) );
  NAND4_X1 U12922 ( .A1(n11464), .A2(n11463), .A3(n11462), .A4(n11461), .ZN(
        n11470) );
  AOI22_X1 U12923 ( .A1(n14223), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n14224), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11468) );
  AOI22_X1 U12924 ( .A1(n14222), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n14225), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11467) );
  AOI22_X1 U12925 ( .A1(n14231), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11466) );
  AOI22_X1 U12926 ( .A1(n14216), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n14233), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11465) );
  NAND4_X1 U12927 ( .A1(n11468), .A2(n11467), .A3(n11466), .A4(n11465), .ZN(
        n11469) );
  NOR2_X1 U12928 ( .A1(n11470), .A2(n11469), .ZN(n12292) );
  OR2_X1 U12929 ( .A1(P2_EBX_REG_0__SCAN_IN), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(
        n11471) );
  INV_X1 U12930 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n11503) );
  INV_X1 U12931 ( .A(n11472), .ZN(n11473) );
  NAND2_X1 U12932 ( .A1(n11474), .A2(n11473), .ZN(n11476) );
  NAND2_X1 U12933 ( .A1(n19221), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11475) );
  XNOR2_X1 U12934 ( .A(n11520), .B(n11519), .ZN(n12015) );
  INV_X1 U12935 ( .A(n14231), .ZN(n11479) );
  INV_X1 U12936 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12396) );
  INV_X1 U12937 ( .A(n11788), .ZN(n11478) );
  INV_X1 U12938 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11477) );
  OAI22_X1 U12939 ( .A1(n11479), .A2(n12396), .B1(n11478), .B2(n11477), .ZN(
        n11485) );
  INV_X1 U12940 ( .A(n11480), .ZN(n14174) );
  INV_X1 U12941 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11483) );
  INV_X1 U12942 ( .A(n11481), .ZN(n11482) );
  INV_X1 U12943 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n19530) );
  OAI22_X1 U12944 ( .A1(n14174), .A2(n11483), .B1(n11482), .B2(n19530), .ZN(
        n11484) );
  NOR2_X1 U12945 ( .A1(n11485), .A2(n11484), .ZN(n11500) );
  AOI22_X1 U12946 ( .A1(n14223), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n14222), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11489) );
  NAND2_X1 U12947 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n11488) );
  NAND2_X1 U12948 ( .A1(n14172), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11487) );
  AOI22_X1 U12949 ( .A1(n14224), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14225), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11486) );
  AND4_X1 U12950 ( .A1(n11489), .A2(n11488), .A3(n11487), .A4(n11486), .ZN(
        n11499) );
  INV_X1 U12951 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11492) );
  NAND2_X1 U12952 ( .A1(n14215), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11491) );
  NAND2_X1 U12953 ( .A1(n16892), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n11490) );
  OAI211_X1 U12954 ( .C1(n11492), .C2(n14219), .A(n11491), .B(n11490), .ZN(
        n11493) );
  INV_X1 U12955 ( .A(n11493), .ZN(n11498) );
  INV_X1 U12956 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19557) );
  INV_X1 U12957 ( .A(n14216), .ZN(n14187) );
  NAND2_X1 U12958 ( .A1(n14232), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n11495) );
  NAND2_X1 U12959 ( .A1(n14233), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n11494) );
  OAI211_X1 U12960 ( .C1(n19557), .C2(n14187), .A(n11495), .B(n11494), .ZN(
        n11496) );
  INV_X1 U12961 ( .A(n11496), .ZN(n11497) );
  NAND4_X1 U12962 ( .A1(n11500), .A2(n11499), .A3(n11498), .A4(n11497), .ZN(
        n12308) );
  NOR2_X1 U12963 ( .A1(n11691), .A2(n12308), .ZN(n11501) );
  NOR2_X1 U12964 ( .A1(n12037), .A2(n11501), .ZN(n11502) );
  MUX2_X1 U12965 ( .A(n11503), .B(n11502), .S(n13849), .Z(n11861) );
  AOI22_X1 U12966 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11481), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11507) );
  AOI22_X1 U12967 ( .A1(n14172), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14230), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11506) );
  AOI22_X1 U12968 ( .A1(n14216), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n14232), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11505) );
  NAND2_X1 U12969 ( .A1(n12385), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11504) );
  AOI22_X1 U12970 ( .A1(n14223), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n14222), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11511) );
  NAND2_X1 U12971 ( .A1(n14231), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11510) );
  AOI22_X1 U12972 ( .A1(n14224), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14225), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11509) );
  NAND2_X1 U12973 ( .A1(n11480), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11508) );
  NAND4_X1 U12974 ( .A1(n11511), .A2(n11510), .A3(n11509), .A4(n11508), .ZN(
        n11516) );
  INV_X1 U12975 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11514) );
  NAND2_X1 U12976 ( .A1(n14215), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11513) );
  NAND2_X1 U12977 ( .A1(n16892), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11512) );
  OAI211_X1 U12978 ( .C1(n11514), .C2(n14219), .A(n11513), .B(n11512), .ZN(
        n11515) );
  NOR2_X1 U12979 ( .A1(n11516), .A2(n11515), .ZN(n11517) );
  NAND2_X1 U12980 ( .A1(n11700), .A2(n12313), .ZN(n11522) );
  NOR2_X1 U12981 ( .A1(n11613), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11518) );
  NOR2_X1 U12982 ( .A1(n18619), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n11521) );
  AND2_X1 U12983 ( .A1(n12022), .A2(n11521), .ZN(n12016) );
  NAND2_X1 U12984 ( .A1(n11691), .A2(n12016), .ZN(n12019) );
  NAND2_X1 U12985 ( .A1(n11522), .A2(n12019), .ZN(n12038) );
  INV_X1 U12986 ( .A(n12038), .ZN(n11524) );
  INV_X1 U12987 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n11523) );
  MUX2_X1 U12988 ( .A(n11524), .B(n11523), .S(n19400), .Z(n11871) );
  AOI22_X1 U12989 ( .A1(n14172), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11480), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11532) );
  INV_X1 U12990 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11527) );
  NAND2_X1 U12991 ( .A1(n14215), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11526) );
  NAND2_X1 U12992 ( .A1(n14216), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11525) );
  OAI211_X1 U12993 ( .C1(n11527), .C2(n14219), .A(n11526), .B(n11525), .ZN(
        n11528) );
  INV_X1 U12994 ( .A(n11528), .ZN(n11531) );
  AOI22_X1 U12995 ( .A1(n14223), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n14222), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11530) );
  AOI22_X1 U12996 ( .A1(n14224), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14225), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11529) );
  NAND4_X1 U12997 ( .A1(n11532), .A2(n11531), .A3(n11530), .A4(n11529), .ZN(
        n11538) );
  AOI22_X1 U12998 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11481), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U12999 ( .A1(n14231), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14230), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11535) );
  AOI22_X1 U13000 ( .A1(n16892), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14232), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11534) );
  NAND2_X1 U13001 ( .A1(n12385), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11533) );
  NAND4_X1 U13002 ( .A1(n11536), .A2(n11535), .A3(n11534), .A4(n11533), .ZN(
        n11537) );
  NOR2_X1 U13003 ( .A1(n11538), .A2(n11537), .ZN(n12318) );
  MUX2_X1 U13004 ( .A(P2_EBX_REG_5__SCAN_IN), .B(n12318), .S(n13849), .Z(
        n11857) );
  AOI22_X1 U13005 ( .A1(n14172), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11480), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11546) );
  INV_X1 U13006 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11541) );
  NAND2_X1 U13007 ( .A1(n14215), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11540) );
  NAND2_X1 U13008 ( .A1(n14216), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11539) );
  OAI211_X1 U13009 ( .C1(n11541), .C2(n14219), .A(n11540), .B(n11539), .ZN(
        n11542) );
  INV_X1 U13010 ( .A(n11542), .ZN(n11545) );
  AOI22_X1 U13011 ( .A1(n14223), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n14222), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11544) );
  AOI22_X1 U13012 ( .A1(n14224), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14225), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11543) );
  NAND4_X1 U13013 ( .A1(n11546), .A2(n11545), .A3(n11544), .A4(n11543), .ZN(
        n11552) );
  AOI22_X1 U13014 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11481), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11550) );
  AOI22_X1 U13015 ( .A1(n14231), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14230), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11549) );
  AOI22_X1 U13016 ( .A1(n16892), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14232), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11548) );
  NAND2_X1 U13017 ( .A1(n12385), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11547) );
  NAND4_X1 U13018 ( .A1(n11550), .A2(n11549), .A3(n11548), .A4(n11547), .ZN(
        n11551) );
  MUX2_X1 U13019 ( .A(P2_EBX_REG_6__SCAN_IN), .B(n12323), .S(n13849), .Z(
        n11553) );
  NAND2_X1 U13020 ( .A1(n11903), .A2(n11902), .ZN(n11910) );
  AOI22_X1 U13021 ( .A1(n14215), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14184), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11566) );
  AOI22_X1 U13022 ( .A1(n14172), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11480), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11565) );
  INV_X1 U13023 ( .A(n14223), .ZN(n11556) );
  INV_X1 U13024 ( .A(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11555) );
  INV_X1 U13025 ( .A(n14222), .ZN(n11554) );
  INV_X1 U13026 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n19322) );
  OAI22_X1 U13027 ( .A1(n11556), .A2(n11555), .B1(n11554), .B2(n19322), .ZN(
        n11562) );
  INV_X1 U13028 ( .A(n14225), .ZN(n11560) );
  INV_X1 U13029 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11559) );
  INV_X1 U13030 ( .A(n14224), .ZN(n11558) );
  INV_X1 U13031 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11557) );
  OAI22_X1 U13032 ( .A1(n11560), .A2(n11559), .B1(n11558), .B2(n11557), .ZN(
        n11561) );
  NOR2_X1 U13033 ( .A1(n11562), .A2(n11561), .ZN(n11564) );
  NAND2_X1 U13034 ( .A1(n14216), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11563) );
  NAND4_X1 U13035 ( .A1(n11566), .A2(n11565), .A3(n11564), .A4(n11563), .ZN(
        n11572) );
  AOI22_X1 U13036 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11481), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U13037 ( .A1(n14231), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14230), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U13038 ( .A1(n16892), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14232), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11568) );
  NAND2_X1 U13039 ( .A1(n12385), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11567) );
  NAND4_X1 U13040 ( .A1(n11570), .A2(n11569), .A3(n11568), .A4(n11567), .ZN(
        n11571) );
  MUX2_X1 U13041 ( .A(n14411), .B(P2_EBX_REG_7__SCAN_IN), .S(n19400), .Z(
        n11908) );
  INV_X1 U13042 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n11574) );
  NOR2_X1 U13043 ( .A1(n13849), .A2(n11574), .ZN(n11912) );
  INV_X1 U13044 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n11575) );
  NAND2_X1 U13045 ( .A1(n19400), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n11919) );
  NAND2_X1 U13046 ( .A1(n11921), .A2(n11919), .ZN(n11928) );
  INV_X1 U13047 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n11576) );
  NOR2_X1 U13048 ( .A1(n13849), .A2(n11576), .ZN(n11927) );
  INV_X1 U13049 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n11579) );
  NOR2_X1 U13050 ( .A1(n13849), .A2(n11579), .ZN(n11915) );
  NAND2_X1 U13051 ( .A1(n19400), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n11945) );
  INV_X1 U13052 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n11580) );
  NOR2_X1 U13053 ( .A1(n13849), .A2(n11580), .ZN(n11942) );
  INV_X1 U13054 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n11581) );
  NOR2_X1 U13055 ( .A1(n13849), .A2(n11581), .ZN(n11938) );
  INV_X1 U13056 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n11582) );
  INV_X1 U13057 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n11583) );
  INV_X1 U13058 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n18438) );
  NOR2_X1 U13059 ( .A1(n13849), .A2(n18438), .ZN(n11958) );
  NAND2_X1 U13060 ( .A1(n19400), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n11933) );
  INV_X1 U13061 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n11585) );
  NOR2_X1 U13062 ( .A1(n13849), .A2(n11585), .ZN(n11975) );
  INV_X1 U13063 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n18469) );
  NOR2_X1 U13064 ( .A1(n13849), .A2(n18469), .ZN(n11982) );
  NAND2_X1 U13065 ( .A1(n19400), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n11993) );
  INV_X1 U13066 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n11586) );
  NOR2_X1 U13067 ( .A1(n13849), .A2(n11586), .ZN(n11988) );
  INV_X1 U13068 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n18513) );
  NOR2_X1 U13069 ( .A1(n13849), .A2(n18513), .ZN(n11589) );
  NAND2_X1 U13070 ( .A1(n19400), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n11998) );
  XOR2_X1 U13071 ( .A(n13847), .B(n13848), .Z(n18535) );
  NOR2_X1 U13072 ( .A1(n11587), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14409) );
  INV_X1 U13073 ( .A(n11587), .ZN(n11588) );
  INV_X1 U13074 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12505) );
  NOR2_X1 U13075 ( .A1(n14409), .A2(n14441), .ZN(n12006) );
  AND2_X1 U13076 ( .A1(n11590), .A2(n11589), .ZN(n11591) );
  OR2_X1 U13077 ( .A1(n11591), .A2(n11997), .ZN(n18510) );
  AOI22_X1 U13078 ( .A1(n15319), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n14360), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11593) );
  AOI22_X1 U13079 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11651), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11592) );
  AND3_X1 U13080 ( .A1(n11593), .A2(n11592), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11596) );
  AOI22_X1 U13081 ( .A1(n14373), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11595) );
  AOI22_X1 U13082 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10974), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11594) );
  NAND3_X1 U13083 ( .A1(n11596), .A2(n11595), .A3(n11594), .ZN(n11603) );
  AOI22_X1 U13084 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11651), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11597) );
  AOI22_X1 U13085 ( .A1(n14373), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U13086 ( .A1(n15319), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n14200), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11599) );
  AOI22_X1 U13087 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10974), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11598) );
  NAND4_X1 U13088 ( .A1(n11601), .A2(n11600), .A3(n11599), .A4(n11598), .ZN(
        n11602) );
  AOI22_X1 U13089 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10974), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11607) );
  AOI22_X1 U13090 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11651), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11606) );
  AOI22_X1 U13091 ( .A1(n11633), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11605) );
  NAND4_X1 U13092 ( .A1(n11607), .A2(n11606), .A3(n11605), .A4(n11604), .ZN(
        n11608) );
  NAND2_X1 U13093 ( .A1(n11608), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11616) );
  AOI22_X1 U13094 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10975), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11612) );
  AOI22_X1 U13095 ( .A1(n15319), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14360), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11611) );
  AOI22_X1 U13096 ( .A1(n11633), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11610) );
  AOI22_X1 U13097 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11651), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11609) );
  NAND4_X1 U13098 ( .A1(n11612), .A2(n11611), .A3(n11610), .A4(n11609), .ZN(
        n11614) );
  NAND2_X1 U13099 ( .A1(n11614), .A2(n11613), .ZN(n11615) );
  XNOR2_X1 U13100 ( .A(n11661), .B(n11643), .ZN(n12065) );
  AOI22_X1 U13101 ( .A1(n14373), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11620) );
  AOI22_X1 U13102 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10975), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11619) );
  AOI22_X1 U13103 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11651), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U13104 ( .A1(n15319), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n14360), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11617) );
  NAND4_X1 U13105 ( .A1(n11620), .A2(n11619), .A3(n11618), .A4(n11617), .ZN(
        n11621) );
  NAND2_X1 U13106 ( .A1(n11621), .A2(n11613), .ZN(n11628) );
  AOI22_X1 U13107 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10975), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11625) );
  AOI22_X1 U13108 ( .A1(n15319), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n14360), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U13109 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11651), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11623) );
  AOI22_X1 U13110 ( .A1(n11633), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11622) );
  NAND4_X1 U13111 ( .A1(n11625), .A2(n11624), .A3(n11623), .A4(n11622), .ZN(
        n11626) );
  NAND2_X1 U13112 ( .A1(n11626), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11627) );
  CLKBUF_X3 U13113 ( .A(n11668), .Z(n15200) );
  AOI22_X1 U13114 ( .A1(n11633), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11632) );
  AOI22_X1 U13115 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10974), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11631) );
  AOI22_X1 U13116 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11651), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11630) );
  NAND4_X1 U13117 ( .A1(n11632), .A2(n11631), .A3(n11630), .A4(n11629), .ZN(
        n11639) );
  AOI22_X1 U13118 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10974), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11636) );
  AOI22_X1 U13119 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11651), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11635) );
  AOI22_X1 U13120 ( .A1(n15319), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n14360), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11634) );
  NAND4_X1 U13121 ( .A1(n11637), .A2(n11636), .A3(n11635), .A4(n11634), .ZN(
        n11638) );
  NAND2_X1 U13122 ( .A1(n11662), .A2(n11643), .ZN(n11644) );
  INV_X1 U13123 ( .A(n11644), .ZN(n11669) );
  NAND2_X1 U13124 ( .A1(n11642), .A2(n11641), .ZN(n11731) );
  NAND2_X1 U13125 ( .A1(n11731), .A2(n11700), .ZN(n11667) );
  NAND2_X1 U13126 ( .A1(n12057), .A2(n11668), .ZN(n11693) );
  AOI22_X1 U13127 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10975), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11649) );
  AOI22_X1 U13128 ( .A1(n14373), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11648) );
  AOI22_X1 U13129 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11651), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11647) );
  AOI22_X1 U13130 ( .A1(n15319), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14200), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U13131 ( .A1(n15319), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n14360), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U13132 ( .A1(n14373), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11656) );
  AOI22_X1 U13133 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11651), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11653) );
  AOI22_X1 U13134 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10974), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11654) );
  NAND4_X1 U13135 ( .A1(n11657), .A2(n11656), .A3(n11655), .A4(n11654), .ZN(
        n11658) );
  NAND4_X1 U13136 ( .A1(n11689), .A2(n11660), .A3(n11663), .A4(n11680), .ZN(
        n11665) );
  NAND2_X1 U13137 ( .A1(n11665), .A2(n11679), .ZN(n12247) );
  NAND2_X1 U13138 ( .A1(n12247), .A2(n11732), .ZN(n11666) );
  INV_X4 U13139 ( .A(n11681), .ZN(n19686) );
  NAND2_X1 U13140 ( .A1(n11667), .A2(n11733), .ZN(n11676) );
  INV_X1 U13141 ( .A(n12059), .ZN(n11674) );
  NAND2_X1 U13142 ( .A1(n12052), .A2(n11672), .ZN(n11673) );
  INV_X1 U13143 ( .A(n18240), .ZN(n11675) );
  AOI21_X2 U13144 ( .B1(n11676), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n11727), 
        .ZN(n11717) );
  AOI21_X1 U13145 ( .B1(n18669), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n11677) );
  OAI21_X1 U13146 ( .B1(n11717), .B2(n11454), .A(n11677), .ZN(n11704) );
  NAND2_X1 U13147 ( .A1(n12059), .A2(n18240), .ZN(n14502) );
  INV_X1 U13148 ( .A(n14502), .ZN(n11678) );
  INV_X2 U13149 ( .A(n12286), .ZN(n11774) );
  NAND2_X2 U13150 ( .A1(n11678), .A2(n11774), .ZN(n12237) );
  BUF_X8 U13151 ( .A(n12237), .Z(n14452) );
  INV_X1 U13152 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n14561) );
  NAND2_X1 U13153 ( .A1(n12275), .A2(n12286), .ZN(n11697) );
  NAND3_X1 U13154 ( .A1(n12254), .A2(n14388), .A3(n10971), .ZN(n11683) );
  NAND3_X1 U13155 ( .A1(n19686), .A2(n11685), .A3(n11684), .ZN(n11687) );
  NAND2_X1 U13156 ( .A1(n11687), .A2(n11245), .ZN(n11688) );
  NAND2_X1 U13157 ( .A1(n11689), .A2(n11688), .ZN(n11696) );
  INV_X1 U13158 ( .A(n11690), .ZN(n11692) );
  INV_X1 U13159 ( .A(n11693), .ZN(n11694) );
  NAND2_X1 U13160 ( .A1(n12251), .A2(n11694), .ZN(n11695) );
  NAND2_X1 U13161 ( .A1(n12244), .A2(n11699), .ZN(n11721) );
  NAND3_X1 U13162 ( .A1(n11697), .A2(n11383), .A3(n11721), .ZN(n11698) );
  INV_X1 U13163 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11869) );
  AOI22_X1 U13164 ( .A1(n11719), .A2(P2_EBX_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11701) );
  OR2_X2 U13165 ( .A1(n11704), .A2(n11703), .ZN(n11738) );
  NAND2_X1 U13166 ( .A1(n11704), .A2(n10962), .ZN(n11705) );
  AND2_X2 U13167 ( .A1(n11738), .A2(n11705), .ZN(n11744) );
  NAND2_X1 U13168 ( .A1(n11383), .A2(n11706), .ZN(n12241) );
  NAND2_X1 U13169 ( .A1(n18669), .A2(n17266), .ZN(n18656) );
  NOR2_X1 U13170 ( .A1(n18656), .A2(n19294), .ZN(n11707) );
  OAI21_X1 U13171 ( .B1(n11717), .B2(n11358), .A(n11708), .ZN(n11716) );
  INV_X1 U13172 ( .A(n11716), .ZN(n11714) );
  INV_X1 U13173 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11712) );
  AOI22_X1 U13174 ( .A1(n11719), .A2(P2_EBX_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11710) );
  INV_X1 U13175 ( .A(n11715), .ZN(n11713) );
  NAND3_X1 U13176 ( .A1(n11699), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n11700), 
        .ZN(n11718) );
  NAND2_X1 U13177 ( .A1(n11741), .A2(n15176), .ZN(n11720) );
  INV_X1 U13179 ( .A(n11722), .ZN(n11724) );
  NOR2_X1 U13180 ( .A1(n18656), .A2(n19263), .ZN(n11723) );
  AOI21_X1 U13181 ( .B1(n11724), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n11723), 
        .ZN(n11725) );
  NAND2_X1 U13182 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11726) );
  INV_X1 U13183 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n17283) );
  INV_X1 U13184 ( .A(n11727), .ZN(n11728) );
  OAI21_X1 U13185 ( .B1(n12237), .B2(n17283), .A(n11728), .ZN(n11729) );
  INV_X1 U13186 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14682) );
  OR2_X2 U13187 ( .A1(n11740), .A2(n14682), .ZN(n11737) );
  INV_X1 U13188 ( .A(n11732), .ZN(n11735) );
  INV_X1 U13189 ( .A(n11733), .ZN(n11734) );
  AOI21_X1 U13190 ( .B1(n11731), .B2(n11735), .A(n11734), .ZN(n11736) );
  NAND2_X1 U13191 ( .A1(n11744), .A2(n10970), .ZN(n11739) );
  INV_X1 U13192 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n15292) );
  INV_X1 U13193 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n15289) );
  AOI22_X1 U13194 ( .A1(n14450), .A2(P2_EBX_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11742) );
  INV_X1 U13195 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19213) );
  OAI22_X1 U13196 ( .A1(n11717), .A2(n11613), .B1(n18656), .B2(n19213), .ZN(
        n12127) );
  XNOR2_X1 U13197 ( .A(n11748), .B(n11747), .ZN(n11749) );
  INV_X1 U13198 ( .A(n18258), .ZN(n11757) );
  AND2_X1 U13199 ( .A1(n11746), .A2(n11757), .ZN(n11750) );
  AND2_X1 U13200 ( .A1(n15329), .A2(n11750), .ZN(n11761) );
  AND2_X2 U13201 ( .A1(n11776), .A2(n11761), .ZN(n11832) );
  BUF_X2 U13202 ( .A(n14066), .Z(n15041) );
  AND2_X1 U13203 ( .A1(n15041), .A2(n11750), .ZN(n11762) );
  AND2_X2 U13204 ( .A1(n11776), .A2(n11762), .ZN(n11835) );
  AOI22_X1 U13205 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n11832), .B1(
        n11835), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11766) );
  INV_X1 U13206 ( .A(n11752), .ZN(n11753) );
  NAND2_X1 U13207 ( .A1(n15041), .A2(n15074), .ZN(n11772) );
  INV_X1 U13208 ( .A(n19268), .ZN(n19264) );
  NAND2_X1 U13209 ( .A1(n19264), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11765) );
  AND2_X1 U13210 ( .A1(n11757), .A2(n11756), .ZN(n11773) );
  AND2_X1 U13211 ( .A1(n15041), .A2(n11773), .ZN(n11758) );
  AND2_X2 U13212 ( .A1(n14055), .A2(n11758), .ZN(n15203) );
  NAND2_X1 U13213 ( .A1(n15203), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11760) );
  AND2_X2 U13214 ( .A1(n11776), .A2(n11758), .ZN(n11831) );
  AND2_X2 U13215 ( .A1(n14055), .A2(n11761), .ZN(n19301) );
  AOI22_X1 U13216 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19301), .B1(
        n11834), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11763) );
  NAND4_X1 U13217 ( .A1(n11766), .A2(n11765), .A3(n11764), .A4(n11763), .ZN(
        n11770) );
  INV_X1 U13218 ( .A(n11767), .ZN(n11768) );
  NOR2_X1 U13219 ( .A1(n11782), .A2(n15074), .ZN(n11769) );
  NAND2_X1 U13220 ( .A1(n11769), .A2(n15041), .ZN(n11826) );
  INV_X1 U13221 ( .A(n11826), .ZN(n11812) );
  NOR2_X1 U13222 ( .A1(n11770), .A2(n11032), .ZN(n11787) );
  INV_X1 U13223 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11779) );
  AND2_X1 U13224 ( .A1(n15329), .A2(n11773), .ZN(n11775) );
  AND2_X2 U13225 ( .A1(n14055), .A2(n11775), .ZN(n11830) );
  AND2_X2 U13226 ( .A1(n11776), .A2(n11775), .ZN(n11833) );
  OAI211_X1 U13227 ( .C1(n11840), .C2(n11779), .A(n11778), .B(n11777), .ZN(
        n11780) );
  AOI21_X1 U13228 ( .B1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n11813), .A(
        n11780), .ZN(n11786) );
  OR2_X1 U13229 ( .A1(n15074), .A2(n15041), .ZN(n11781) );
  INV_X1 U13230 ( .A(n19245), .ZN(n19247) );
  INV_X1 U13231 ( .A(n11783), .ZN(n11784) );
  AOI22_X1 U13232 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11481), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11792) );
  AOI22_X1 U13233 ( .A1(n14231), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11788), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11791) );
  AOI22_X1 U13234 ( .A1(n16892), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14232), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11790) );
  NAND2_X1 U13235 ( .A1(n12385), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11789) );
  AND4_X1 U13236 ( .A1(n11792), .A2(n11791), .A3(n11790), .A4(n11789), .ZN(
        n11803) );
  AOI22_X1 U13237 ( .A1(n14223), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14222), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11796) );
  NAND2_X1 U13238 ( .A1(n14172), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11795) );
  AOI22_X1 U13239 ( .A1(n14224), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14225), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11794) );
  NAND2_X1 U13240 ( .A1(n11480), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11793) );
  NAND4_X1 U13241 ( .A1(n11796), .A2(n11795), .A3(n11794), .A4(n11793), .ZN(
        n11801) );
  INV_X1 U13242 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11799) );
  NAND2_X1 U13243 ( .A1(n14215), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11798) );
  INV_X1 U13244 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n19797) );
  NAND2_X1 U13245 ( .A1(n14216), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11797) );
  OAI211_X1 U13246 ( .C1(n11799), .C2(n14219), .A(n11798), .B(n11797), .ZN(
        n11800) );
  NOR2_X1 U13247 ( .A1(n11801), .A2(n11800), .ZN(n11802) );
  NAND2_X1 U13248 ( .A1(n12285), .A2(n19621), .ZN(n14549) );
  OR2_X1 U13249 ( .A1(n12292), .A2(n14549), .ZN(n12080) );
  NAND2_X1 U13250 ( .A1(n12080), .A2(n11804), .ZN(n11805) );
  INV_X1 U13251 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11806) );
  INV_X1 U13252 ( .A(n11807), .ZN(n11821) );
  AOI22_X1 U13253 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n11830), .B1(
        n11831), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11811) );
  AOI22_X1 U13254 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n15203), .B1(
        n11835), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11810) );
  AOI22_X1 U13255 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19301), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11809) );
  AOI22_X1 U13256 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11834), .B1(
        n11833), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11808) );
  INV_X1 U13257 ( .A(n11825), .ZN(n11813) );
  INV_X1 U13258 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11814) );
  OAI22_X1 U13259 ( .A1(n11814), .A2(n19310), .B1(n19268), .B2(n12396), .ZN(
        n11817) );
  INV_X1 U13260 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11815) );
  NOR2_X1 U13261 ( .A1(n11817), .A2(n11816), .ZN(n11818) );
  INV_X1 U13262 ( .A(n11855), .ZN(n11853) );
  INV_X1 U13263 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n14932) );
  INV_X1 U13264 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n14329) );
  OAI22_X1 U13265 ( .A1(n14932), .A2(n11823), .B1(n19245), .B2(n14329), .ZN(
        n11824) );
  INV_X1 U13266 ( .A(n11824), .ZN(n11849) );
  INV_X1 U13267 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11828) );
  INV_X1 U13268 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11827) );
  OAI22_X1 U13269 ( .A1(n11828), .A2(n11825), .B1(n19215), .B2(n11827), .ZN(
        n11829) );
  INV_X1 U13270 ( .A(n11829), .ZN(n11848) );
  AOI22_X1 U13271 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n11830), .B1(
        n11831), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11839) );
  AOI22_X1 U13272 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n15203), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11838) );
  AOI22_X1 U13273 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19301), .B1(
        n11833), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U13274 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n11834), .B1(
        n11835), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11836) );
  INV_X1 U13275 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14177) );
  INV_X1 U13276 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11841) );
  OAI22_X1 U13277 ( .A1(n14177), .A2(n19310), .B1(n11840), .B2(n11841), .ZN(
        n11845) );
  INV_X1 U13278 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12424) );
  INV_X1 U13279 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11843) );
  OAI22_X1 U13280 ( .A1(n12424), .A2(n19268), .B1(n11842), .B2(n11843), .ZN(
        n11844) );
  NOR2_X1 U13281 ( .A1(n11845), .A2(n11844), .ZN(n11846) );
  NAND4_X1 U13282 ( .A1(n11849), .A2(n11848), .A3(n11847), .A4(n11846), .ZN(
        n11851) );
  NAND2_X1 U13283 ( .A1(n12318), .A2(n19621), .ZN(n11850) );
  INV_X1 U13284 ( .A(n11854), .ZN(n11852) );
  AND2_X1 U13285 ( .A1(n11856), .A2(n11857), .ZN(n11858) );
  OR2_X1 U13286 ( .A1(n11858), .A2(n11903), .ZN(n18279) );
  NAND2_X1 U13287 ( .A1(n15474), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11879) );
  NOR2_X1 U13288 ( .A1(n11862), .A2(n11861), .ZN(n11863) );
  OR2_X1 U13289 ( .A1(n11872), .A2(n11863), .ZN(n15051) );
  OAI21_X1 U13290 ( .B1(n15290), .B2(n14446), .A(n15051), .ZN(n15287) );
  OAI21_X1 U13291 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19263), .A(
        n12007), .ZN(n12048) );
  INV_X1 U13292 ( .A(n12048), .ZN(n12011) );
  MUX2_X1 U13293 ( .A(n12285), .B(n12011), .S(n11691), .Z(n12034) );
  MUX2_X1 U13294 ( .A(n12034), .B(P2_EBX_REG_0__SCAN_IN), .S(n19400), .Z(
        n18255) );
  AND2_X1 U13295 ( .A1(n18255), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n11866) );
  INV_X1 U13296 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n14696) );
  NAND3_X1 U13297 ( .A1(n19400), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n11864) );
  NAND2_X1 U13298 ( .A1(n11868), .A2(n11864), .ZN(n15072) );
  INV_X1 U13299 ( .A(n15072), .ZN(n11865) );
  NOR2_X1 U13300 ( .A1(n11866), .A2(n11865), .ZN(n14614) );
  AND2_X1 U13301 ( .A1(n11866), .A2(n11865), .ZN(n14613) );
  NOR2_X1 U13302 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14613), .ZN(
        n14612) );
  NOR2_X1 U13303 ( .A1(n14614), .A2(n14612), .ZN(n14557) );
  XNOR2_X1 U13304 ( .A(n11867), .B(n11868), .ZN(n15039) );
  XNOR2_X1 U13305 ( .A(n15039), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n14556) );
  NOR2_X1 U13306 ( .A1(n15039), .A2(n11869), .ZN(n11870) );
  AOI21_X1 U13307 ( .B1(n14557), .B2(n14556), .A(n11870), .ZN(n11873) );
  OAI21_X1 U13308 ( .B1(n11872), .B2(n11871), .A(n11856), .ZN(n18267) );
  INV_X1 U13309 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n15479) );
  AND2_X1 U13310 ( .A1(n18267), .A2(n15479), .ZN(n11874) );
  AOI21_X1 U13311 ( .B1(n11873), .B2(n15289), .A(n11874), .ZN(n11878) );
  INV_X1 U13312 ( .A(n11873), .ZN(n15357) );
  INV_X1 U13313 ( .A(n11874), .ZN(n11875) );
  NAND3_X1 U13314 ( .A1(n15357), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n11875), .ZN(n11876) );
  OAI21_X1 U13315 ( .B1(n15479), .B2(n18267), .A(n11876), .ZN(n11877) );
  AOI21_X1 U13316 ( .B1(n15287), .B2(n11878), .A(n11877), .ZN(n15475) );
  NAND2_X1 U13317 ( .A1(n11879), .A2(n15475), .ZN(n11882) );
  INV_X1 U13318 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n15478) );
  NAND3_X1 U13319 ( .A1(n11880), .A2(n15478), .A3(n18279), .ZN(n11881) );
  INV_X1 U13320 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19392) );
  INV_X1 U13321 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11883) );
  OAI22_X1 U13322 ( .A1(n19392), .A2(n11823), .B1(n19215), .B2(n11883), .ZN(
        n11884) );
  INV_X1 U13323 ( .A(n11884), .ZN(n11899) );
  INV_X1 U13324 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11886) );
  INV_X1 U13325 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11885) );
  OAI22_X1 U13326 ( .A1(n11886), .A2(n11825), .B1(n19245), .B2(n11885), .ZN(
        n11887) );
  INV_X1 U13327 ( .A(n11887), .ZN(n11898) );
  AOI22_X1 U13328 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n11830), .B1(
        n11835), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U13329 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19301), .B1(
        n11831), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11890) );
  AOI22_X1 U13330 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n15203), .B1(
        n11833), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11889) );
  AOI22_X1 U13331 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n11834), .B1(
        n11832), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11888) );
  INV_X1 U13332 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14186) );
  INV_X1 U13333 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12445) );
  OAI22_X1 U13334 ( .A1(n14186), .A2(n19310), .B1(n19268), .B2(n12445), .ZN(
        n11895) );
  INV_X1 U13335 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11893) );
  INV_X1 U13336 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11892) );
  OAI22_X1 U13337 ( .A1(n11893), .A2(n11842), .B1(n11840), .B2(n11892), .ZN(
        n11894) );
  NOR2_X1 U13338 ( .A1(n11895), .A2(n11894), .ZN(n11896) );
  NAND4_X1 U13339 ( .A1(n11899), .A2(n11898), .A3(n11897), .A4(n11896), .ZN(
        n11901) );
  NAND2_X1 U13340 ( .A1(n12323), .A2(n19621), .ZN(n11900) );
  NAND2_X1 U13341 ( .A1(n12092), .A2(n14411), .ZN(n11905) );
  OR2_X1 U13342 ( .A1(n11903), .A2(n11902), .ZN(n11904) );
  NAND2_X1 U13343 ( .A1(n11910), .A2(n11904), .ZN(n18290) );
  INV_X1 U13344 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16834) );
  INV_X1 U13345 ( .A(n11908), .ZN(n11909) );
  XNOR2_X1 U13346 ( .A(n11910), .B(n11909), .ZN(n18304) );
  AND2_X1 U13347 ( .A1(n18304), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16587) );
  NAND2_X1 U13348 ( .A1(n11911), .A2(n11912), .ZN(n11913) );
  NAND2_X1 U13349 ( .A1(n11925), .A2(n11913), .ZN(n18313) );
  AND2_X1 U13350 ( .A1(n14446), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12102) );
  INV_X1 U13351 ( .A(n12102), .ZN(n11914) );
  NOR2_X1 U13352 ( .A1(n18313), .A2(n11914), .ZN(n16823) );
  NAND2_X1 U13353 ( .A1(n16823), .A2(n16586), .ZN(n16440) );
  AND2_X1 U13354 ( .A1(n11930), .A2(n11915), .ZN(n11916) );
  OR2_X1 U13355 ( .A1(n11916), .A2(n11011), .ZN(n18356) );
  INV_X1 U13356 ( .A(n18356), .ZN(n11917) );
  NAND2_X1 U13357 ( .A1(n11917), .A2(n14446), .ZN(n11948) );
  INV_X1 U13358 ( .A(n11948), .ZN(n11918) );
  NAND2_X1 U13359 ( .A1(n11918), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17246) );
  INV_X1 U13360 ( .A(n11919), .ZN(n11920) );
  XNOR2_X1 U13361 ( .A(n11921), .B(n11920), .ZN(n18335) );
  AND2_X1 U13362 ( .A1(n14446), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11922) );
  NAND2_X1 U13363 ( .A1(n18335), .A2(n11922), .ZN(n16797) );
  INV_X1 U13364 ( .A(n11923), .ZN(n11924) );
  XNOR2_X1 U13365 ( .A(n11925), .B(n11924), .ZN(n18322) );
  AND2_X1 U13366 ( .A1(n14446), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11926) );
  NAND2_X1 U13367 ( .A1(n18322), .A2(n11926), .ZN(n16795) );
  AND2_X1 U13368 ( .A1(n16797), .A2(n16795), .ZN(n16566) );
  NAND2_X1 U13369 ( .A1(n11928), .A2(n11927), .ZN(n11929) );
  AND2_X1 U13370 ( .A1(n11930), .A2(n11929), .ZN(n18344) );
  AND2_X1 U13371 ( .A1(n14446), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11931) );
  NAND2_X1 U13372 ( .A1(n18344), .A2(n11931), .ZN(n16568) );
  AND2_X1 U13373 ( .A1(n16440), .A2(n16522), .ZN(n11932) );
  AOI21_X1 U13374 ( .B1(n11962), .B2(n14446), .A(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16455) );
  XNOR2_X1 U13375 ( .A(n11934), .B(n11378), .ZN(n11964) );
  NAND2_X1 U13376 ( .A1(n11964), .A2(n14446), .ZN(n11935) );
  INV_X1 U13377 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n18596) );
  NAND2_X1 U13378 ( .A1(n11935), .A2(n18596), .ZN(n16477) );
  XNOR2_X1 U13379 ( .A(n11936), .B(n11059), .ZN(n18415) );
  NAND2_X1 U13380 ( .A1(n18415), .A2(n14446), .ZN(n11937) );
  INV_X1 U13381 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16489) );
  NAND2_X1 U13382 ( .A1(n11937), .A2(n16489), .ZN(n16491) );
  INV_X1 U13383 ( .A(n11938), .ZN(n11939) );
  XNOR2_X1 U13384 ( .A(n11944), .B(n11939), .ZN(n18391) );
  NAND2_X1 U13385 ( .A1(n18391), .A2(n14446), .ZN(n11940) );
  XNOR2_X1 U13386 ( .A(n11940), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16515) );
  NAND2_X1 U13387 ( .A1(n11941), .A2(n11942), .ZN(n11943) );
  NAND2_X1 U13388 ( .A1(n11944), .A2(n11943), .ZN(n18380) );
  NOR2_X1 U13389 ( .A1(n18380), .A2(n14411), .ZN(n11969) );
  OR2_X1 U13390 ( .A1(n11969), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n16531) );
  XNOR2_X1 U13391 ( .A(n11011), .B(n11060), .ZN(n14484) );
  AOI21_X1 U13392 ( .B1(n14484), .B2(n14446), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16526) );
  INV_X1 U13393 ( .A(n16526), .ZN(n16525) );
  OR2_X1 U13394 ( .A1(n11946), .A2(n11945), .ZN(n11947) );
  NAND2_X1 U13395 ( .A1(n11941), .A2(n11947), .ZN(n18369) );
  NOR2_X1 U13396 ( .A1(n18369), .A2(n14411), .ZN(n11970) );
  OR2_X1 U13397 ( .A1(n11970), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16528) );
  INV_X1 U13398 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17253) );
  NAND2_X1 U13399 ( .A1(n11948), .A2(n17253), .ZN(n17247) );
  NAND4_X1 U13400 ( .A1(n16531), .A2(n16525), .A3(n16528), .A4(n17247), .ZN(
        n16443) );
  NAND2_X1 U13401 ( .A1(n18344), .A2(n14446), .ZN(n11950) );
  INV_X1 U13402 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11949) );
  NAND2_X1 U13403 ( .A1(n11950), .A2(n11949), .ZN(n17248) );
  NAND2_X1 U13404 ( .A1(n18335), .A2(n14446), .ZN(n11951) );
  INV_X1 U13405 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16779) );
  NAND2_X1 U13406 ( .A1(n11951), .A2(n16779), .ZN(n16798) );
  NAND2_X1 U13407 ( .A1(n18322), .A2(n14446), .ZN(n11952) );
  INV_X1 U13408 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16813) );
  NAND2_X1 U13409 ( .A1(n11952), .A2(n16813), .ZN(n16442) );
  INV_X1 U13410 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16837) );
  OAI21_X1 U13411 ( .B1(n18313), .B2(n14411), .A(n16837), .ZN(n16822) );
  NAND4_X1 U13412 ( .A1(n17248), .A2(n16798), .A3(n16442), .A4(n16822), .ZN(
        n11953) );
  NOR2_X1 U13413 ( .A1(n16443), .A2(n11953), .ZN(n11955) );
  XNOR2_X1 U13414 ( .A(n11018), .B(n11374), .ZN(n18403) );
  NAND2_X1 U13415 ( .A1(n18403), .A2(n14446), .ZN(n11954) );
  INV_X1 U13416 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16736) );
  NAND2_X1 U13417 ( .A1(n11954), .A2(n16736), .ZN(n16504) );
  NAND4_X1 U13418 ( .A1(n16450), .A2(n16515), .A3(n11955), .A4(n16504), .ZN(
        n11956) );
  OAI21_X1 U13419 ( .B1(n16455), .B2(n11956), .A(n16522), .ZN(n11957) );
  AND2_X1 U13420 ( .A1(n11959), .A2(n11958), .ZN(n11961) );
  OR2_X1 U13421 ( .A1(n11961), .A2(n11960), .ZN(n18436) );
  AND2_X1 U13422 ( .A1(n14446), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11963) );
  NAND2_X1 U13423 ( .A1(n11962), .A2(n11963), .ZN(n16456) );
  AND2_X1 U13424 ( .A1(n14446), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11965) );
  NAND2_X1 U13425 ( .A1(n11964), .A2(n11965), .ZN(n16476) );
  AND2_X1 U13426 ( .A1(n14446), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11966) );
  NAND2_X1 U13427 ( .A1(n18415), .A2(n11966), .ZN(n16495) );
  NAND2_X1 U13428 ( .A1(n16476), .A2(n16495), .ZN(n16449) );
  AND2_X1 U13429 ( .A1(n14446), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n11967) );
  NAND2_X1 U13430 ( .A1(n18403), .A2(n11967), .ZN(n16503) );
  AND2_X1 U13431 ( .A1(n14446), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11968) );
  NAND2_X1 U13432 ( .A1(n14484), .A2(n11968), .ZN(n16524) );
  NAND2_X1 U13433 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n11969), .ZN(
        n16530) );
  NAND2_X1 U13434 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n11970), .ZN(
        n16527) );
  AND2_X1 U13435 ( .A1(n16530), .A2(n16527), .ZN(n11971) );
  AND2_X1 U13436 ( .A1(n16524), .A2(n11971), .ZN(n16444) );
  AND2_X1 U13437 ( .A1(n14446), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11972) );
  NAND2_X1 U13438 ( .A1(n18391), .A2(n11972), .ZN(n16502) );
  NAND3_X1 U13439 ( .A1(n16503), .A2(n16444), .A3(n16502), .ZN(n11973) );
  NOR2_X1 U13440 ( .A1(n16449), .A2(n11973), .ZN(n11974) );
  INV_X1 U13441 ( .A(n11975), .ZN(n11976) );
  XNOR2_X1 U13442 ( .A(n11977), .B(n11976), .ZN(n18458) );
  NAND2_X1 U13443 ( .A1(n18458), .A2(n14446), .ZN(n16431) );
  NAND2_X1 U13444 ( .A1(n11978), .A2(n16431), .ZN(n11981) );
  INV_X1 U13445 ( .A(n16430), .ZN(n11979) );
  NAND2_X1 U13446 ( .A1(n11979), .A2(n16666), .ZN(n11980) );
  NAND2_X1 U13447 ( .A1(n11981), .A2(n11980), .ZN(n16419) );
  AND2_X1 U13448 ( .A1(n11983), .A2(n11982), .ZN(n11984) );
  OR2_X1 U13449 ( .A1(n11984), .A2(n11012), .ZN(n18467) );
  AOI21_X1 U13450 ( .B1(n11986), .B2(n14446), .A(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16421) );
  AND2_X1 U13451 ( .A1(n14446), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11985) );
  NAND2_X1 U13452 ( .A1(n11986), .A2(n11985), .ZN(n16420) );
  XNOR2_X1 U13453 ( .A(n11012), .B(n11064), .ZN(n18479) );
  NAND2_X1 U13454 ( .A1(n18479), .A2(n14446), .ZN(n16410) );
  INV_X1 U13455 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11987) );
  INV_X1 U13456 ( .A(n11988), .ZN(n11989) );
  NAND2_X1 U13457 ( .A1(n18499), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16366) );
  OR2_X1 U13458 ( .A1(n16366), .A2(n14411), .ZN(n12002) );
  NAND2_X1 U13459 ( .A1(n18499), .A2(n14446), .ZN(n11991) );
  INV_X1 U13460 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16621) );
  NAND2_X1 U13461 ( .A1(n11991), .A2(n16621), .ZN(n11992) );
  NAND2_X1 U13462 ( .A1(n12002), .A2(n11992), .ZN(n16392) );
  INV_X1 U13463 ( .A(n11993), .ZN(n11994) );
  XNOR2_X1 U13464 ( .A(n11995), .B(n11994), .ZN(n18489) );
  NAND2_X1 U13465 ( .A1(n18489), .A2(n14446), .ZN(n12003) );
  INV_X1 U13466 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16637) );
  OAI21_X1 U13467 ( .B1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(n16369), .ZN(n12000) );
  INV_X1 U13468 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16365) );
  INV_X1 U13469 ( .A(n12002), .ZN(n12005) );
  INV_X1 U13470 ( .A(n12003), .ZN(n12004) );
  XOR2_X1 U13471 ( .A(n12006), .B(n14410), .Z(n16364) );
  NAND2_X1 U13472 ( .A1(n19621), .A2(n12048), .ZN(n12008) );
  XNOR2_X1 U13473 ( .A(n12033), .B(n12007), .ZN(n12044) );
  NAND2_X1 U13474 ( .A1(n12008), .A2(n12044), .ZN(n12010) );
  NAND2_X1 U13475 ( .A1(n19621), .A2(n12042), .ZN(n12009) );
  NAND2_X1 U13476 ( .A1(n12010), .A2(n12009), .ZN(n12013) );
  NAND2_X1 U13477 ( .A1(n12033), .A2(n12011), .ZN(n12012) );
  AOI22_X1 U13478 ( .A1(n12013), .A2(n19686), .B1(n11700), .B2(n12012), .ZN(
        n12018) );
  NOR2_X1 U13479 ( .A1(n18240), .A2(n19621), .ZN(n12014) );
  MUX2_X1 U13480 ( .A(n12014), .B(n11700), .S(n12042), .Z(n12017) );
  NOR2_X1 U13481 ( .A1(n12016), .A2(n12015), .ZN(n12041) );
  OAI21_X1 U13482 ( .B1(n12018), .B2(n12017), .A(n12041), .ZN(n12021) );
  INV_X1 U13483 ( .A(n12037), .ZN(n12020) );
  NAND3_X1 U13484 ( .A1(n12021), .A2(n12020), .A3(n12019), .ZN(n12028) );
  INV_X1 U13485 ( .A(n12022), .ZN(n12024) );
  AND2_X1 U13486 ( .A1(n18619), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12023) );
  INV_X1 U13487 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n14646) );
  NAND2_X1 U13488 ( .A1(n14646), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n12025) );
  INV_X1 U13489 ( .A(n12046), .ZN(n12027) );
  NAND2_X1 U13490 ( .A1(n12028), .A2(n12027), .ZN(n12029) );
  MUX2_X1 U13491 ( .A(n12029), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18669), .Z(n12031) );
  NAND2_X1 U13492 ( .A1(n18240), .A2(n12046), .ZN(n12030) );
  NAND2_X1 U13493 ( .A1(n18626), .A2(n11774), .ZN(n14636) );
  NAND2_X1 U13494 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n18675) );
  NAND2_X1 U13495 ( .A1(n21655), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n17343) );
  INV_X1 U13496 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n21640) );
  NOR2_X1 U13497 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_0__SCAN_IN), 
        .ZN(n21641) );
  NAND2_X1 U13498 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n21641), .ZN(n17324) );
  NAND2_X1 U13499 ( .A1(n17339), .A2(n17324), .ZN(n21645) );
  NAND2_X1 U13500 ( .A1(n18675), .A2(n21645), .ZN(n18639) );
  INV_X1 U13501 ( .A(n18639), .ZN(n14637) );
  NAND2_X1 U13502 ( .A1(n14637), .A2(n12069), .ZN(n12076) );
  AOI21_X1 U13503 ( .B1(n12031), .B2(n19686), .A(n11331), .ZN(n12032) );
  NAND2_X1 U13504 ( .A1(n14636), .A2(n12032), .ZN(n12075) );
  NAND2_X1 U13505 ( .A1(n12034), .A2(n12033), .ZN(n12036) );
  NAND2_X1 U13506 ( .A1(n12036), .A2(n12035), .ZN(n12040) );
  NOR2_X1 U13507 ( .A1(n12038), .A2(n12037), .ZN(n12039) );
  AOI21_X1 U13508 ( .B1(n12040), .B2(n12039), .A(n12046), .ZN(n18634) );
  AND2_X1 U13509 ( .A1(n19621), .A2(n12246), .ZN(n12118) );
  NAND2_X1 U13510 ( .A1(n18634), .A2(n12118), .ZN(n14418) );
  NAND2_X1 U13511 ( .A1(n12042), .A2(n12041), .ZN(n12047) );
  INV_X1 U13512 ( .A(n12047), .ZN(n12043) );
  AND2_X1 U13513 ( .A1(n12044), .A2(n12043), .ZN(n12045) );
  OAI21_X1 U13514 ( .B1(n12048), .B2(n12047), .A(n18640), .ZN(n12049) );
  INV_X1 U13515 ( .A(n12049), .ZN(n12051) );
  NAND2_X1 U13516 ( .A1(n12050), .A2(n14646), .ZN(n14642) );
  INV_X1 U13517 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n16921) );
  OAI21_X1 U13518 ( .B1(n14172), .B2(n14642), .A(n16921), .ZN(n17263) );
  MUX2_X1 U13519 ( .A(n12051), .B(n17263), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n18627) );
  NAND2_X1 U13520 ( .A1(n11774), .A2(n18627), .ZN(n12053) );
  AOI21_X1 U13521 ( .B1(n14418), .B2(n12053), .A(n12052), .ZN(n12073) );
  NAND2_X1 U13522 ( .A1(n11355), .A2(n11680), .ZN(n12058) );
  NAND2_X1 U13523 ( .A1(n12055), .A2(n12058), .ZN(n12068) );
  NAND3_X1 U13524 ( .A1(n12059), .A2(n18640), .A3(n14637), .ZN(n12062) );
  NAND2_X1 U13525 ( .A1(n12246), .A2(n15200), .ZN(n12060) );
  OAI211_X1 U13526 ( .C1(n11774), .C2(n11693), .A(n11680), .B(n12060), .ZN(
        n12061) );
  AND4_X1 U13527 ( .A1(n12064), .A2(n12063), .A3(n12062), .A4(n12061), .ZN(
        n12067) );
  NAND2_X1 U13528 ( .A1(n12065), .A2(n15200), .ZN(n12066) );
  NAND2_X1 U13529 ( .A1(n12066), .A2(n12118), .ZN(n12260) );
  AND3_X1 U13530 ( .A1(n12068), .A2(n12067), .A3(n12260), .ZN(n14634) );
  MUX2_X1 U13531 ( .A(n12069), .B(n12059), .S(n11774), .Z(n12070) );
  NAND3_X1 U13532 ( .A1(n12070), .A2(n18640), .A3(n18675), .ZN(n12071) );
  NAND2_X1 U13533 ( .A1(n14634), .A2(n12071), .ZN(n12072) );
  NOR2_X1 U13534 ( .A1(n12073), .A2(n12072), .ZN(n12074) );
  OAI211_X1 U13535 ( .C1(n14636), .C2(n12076), .A(n12075), .B(n12074), .ZN(
        n12077) );
  AND3_X1 U13536 ( .A1(n17266), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n18683) );
  NOR2_X1 U13537 ( .A1(n12052), .A2(n11691), .ZN(n18628) );
  XNOR2_X1 U13538 ( .A(n12292), .B(n12285), .ZN(n12078) );
  AND2_X1 U13539 ( .A1(n14549), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14551) );
  NAND2_X1 U13540 ( .A1(n12078), .A2(n14551), .ZN(n12079) );
  XOR2_X1 U13541 ( .A(n12078), .B(n14551), .Z(n14616) );
  NAND2_X1 U13542 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14616), .ZN(
        n14615) );
  NAND2_X1 U13543 ( .A1(n12079), .A2(n14615), .ZN(n12082) );
  XNOR2_X1 U13544 ( .A(n11869), .B(n12082), .ZN(n14560) );
  INV_X1 U13545 ( .A(n12080), .ZN(n12081) );
  XNOR2_X1 U13546 ( .A(n12298), .B(n12081), .ZN(n14559) );
  NAND2_X1 U13547 ( .A1(n14560), .A2(n14559), .ZN(n14558) );
  NAND2_X1 U13548 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12082), .ZN(
        n12083) );
  NAND2_X1 U13549 ( .A1(n14558), .A2(n12083), .ZN(n12084) );
  XNOR2_X1 U13550 ( .A(n12084), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n15291) );
  NAND2_X1 U13551 ( .A1(n12084), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12085) );
  XNOR2_X1 U13552 ( .A(n12086), .B(n12313), .ZN(n12087) );
  XNOR2_X1 U13553 ( .A(n12088), .B(n12087), .ZN(n15362) );
  NAND2_X1 U13554 ( .A1(n15362), .A2(n15479), .ZN(n15361) );
  INV_X1 U13555 ( .A(n12087), .ZN(n12089) );
  OR2_X1 U13556 ( .A1(n12089), .A2(n12088), .ZN(n12090) );
  NAND2_X1 U13557 ( .A1(n12094), .A2(n12093), .ZN(n12096) );
  INV_X1 U13558 ( .A(n12093), .ZN(n12095) );
  XNOR2_X1 U13559 ( .A(n12106), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16592) );
  INV_X1 U13560 ( .A(n12104), .ZN(n12103) );
  OAI21_X1 U13561 ( .B1(n12104), .B2(n14411), .A(n16837), .ZN(n12105) );
  INV_X1 U13562 ( .A(n16820), .ZN(n12108) );
  INV_X1 U13563 ( .A(n12106), .ZN(n12107) );
  NAND2_X1 U13564 ( .A1(n12107), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16818) );
  AND3_X1 U13565 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16765) );
  AND2_X1 U13566 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12111) );
  AND2_X1 U13567 ( .A1(n16765), .A2(n12111), .ZN(n18568) );
  NAND3_X1 U13568 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16697) );
  INV_X1 U13569 ( .A(n16697), .ZN(n12112) );
  AND2_X1 U13570 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n12112), .ZN(
        n12271) );
  NAND2_X1 U13571 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16704) );
  INV_X1 U13572 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16679) );
  NAND2_X1 U13573 ( .A1(n12114), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n16408) );
  NAND2_X1 U13574 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16655) );
  OR2_X1 U13575 ( .A1(n11987), .A2(n16655), .ZN(n12115) );
  AND2_X1 U13576 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16610) );
  INV_X1 U13577 ( .A(n16378), .ZN(n12116) );
  AOI21_X1 U13578 ( .B1(n12116), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12117) );
  NAND2_X1 U13579 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14461) );
  NOR2_X1 U13580 ( .A1(n12117), .A2(n14467), .ZN(n16356) );
  INV_X1 U13581 ( .A(n16356), .ZN(n12509) );
  INV_X1 U13582 ( .A(n12118), .ZN(n12119) );
  NOR2_X1 U13583 ( .A1(n12052), .A2(n12119), .ZN(n18624) );
  OR2_X1 U13584 ( .A1(n10978), .A2(n12505), .ZN(n12124) );
  INV_X1 U13585 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n17336) );
  NAND2_X1 U13586 ( .A1(n14450), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12121) );
  NAND2_X1 U13587 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12120) );
  OAI211_X1 U13588 ( .C1(n17336), .C2(n14452), .A(n12121), .B(n12120), .ZN(
        n12122) );
  INV_X1 U13589 ( .A(n12122), .ZN(n12123) );
  AND2_X1 U13590 ( .A1(n12124), .A2(n12123), .ZN(n12240) );
  INV_X1 U13591 ( .A(n12125), .ZN(n12129) );
  NOR2_X1 U13592 ( .A1(n12127), .A2(n12126), .ZN(n12128) );
  INV_X1 U13593 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n12132) );
  OR2_X1 U13594 ( .A1(n10978), .A2(n15479), .ZN(n12131) );
  AOI22_X1 U13595 ( .A1(n14450), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12130) );
  OAI211_X1 U13596 ( .C1(n14452), .C2(n12132), .A(n12131), .B(n12130), .ZN(
        n14920) );
  INV_X1 U13597 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n12135) );
  OR2_X1 U13598 ( .A1(n10978), .A2(n15478), .ZN(n12134) );
  AOI22_X1 U13599 ( .A1(n14450), .A2(P2_EBX_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12133) );
  OAI211_X1 U13600 ( .C1(n14452), .C2(n12135), .A(n12134), .B(n12133), .ZN(
        n14883) );
  OR2_X1 U13601 ( .A1(n10978), .A2(n16834), .ZN(n12141) );
  INV_X1 U13602 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n12138) );
  NAND2_X1 U13603 ( .A1(n14450), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n12137) );
  NAND2_X1 U13604 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n12136) );
  OAI211_X1 U13605 ( .C1(n12138), .C2(n14452), .A(n12137), .B(n12136), .ZN(
        n12139) );
  INV_X1 U13606 ( .A(n12139), .ZN(n12140) );
  NAND2_X1 U13607 ( .A1(n12143), .A2(n12142), .ZN(n14929) );
  INV_X1 U13608 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16850) );
  OR2_X1 U13609 ( .A1(n10978), .A2(n16850), .ZN(n12149) );
  INV_X1 U13610 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n12146) );
  NAND2_X1 U13611 ( .A1(n14450), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n12145) );
  NAND2_X1 U13612 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12144) );
  OAI211_X1 U13613 ( .C1(n12146), .C2(n14452), .A(n12145), .B(n12144), .ZN(
        n12147) );
  INV_X1 U13614 ( .A(n12147), .ZN(n12148) );
  OR2_X1 U13615 ( .A1(n10978), .A2(n16837), .ZN(n12154) );
  INV_X1 U13616 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n12349) );
  NAND2_X1 U13617 ( .A1(n14450), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n12151) );
  NAND2_X1 U13618 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12150) );
  OAI211_X1 U13619 ( .C1(n12349), .C2(n14452), .A(n12151), .B(n12150), .ZN(
        n12152) );
  INV_X1 U13620 ( .A(n12152), .ZN(n12153) );
  INV_X1 U13621 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n12157) );
  OR2_X1 U13622 ( .A1(n10978), .A2(n16813), .ZN(n12156) );
  AOI22_X1 U13623 ( .A1(n14450), .A2(P2_EBX_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12155) );
  OAI211_X1 U13624 ( .C1(n14452), .C2(n12157), .A(n12156), .B(n12155), .ZN(
        n15060) );
  INV_X1 U13625 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n12160) );
  OR2_X1 U13626 ( .A1(n10978), .A2(n16779), .ZN(n12159) );
  AOI22_X1 U13627 ( .A1(n14450), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n12158) );
  OAI211_X1 U13628 ( .C1(n14452), .C2(n12160), .A(n12159), .B(n12158), .ZN(
        n15222) );
  OR2_X1 U13629 ( .A1(n10978), .A2(n11949), .ZN(n12166) );
  INV_X1 U13630 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n12163) );
  NAND2_X1 U13631 ( .A1(n14450), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n12162) );
  NAND2_X1 U13632 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12161) );
  OAI211_X1 U13633 ( .C1(n12163), .C2(n14452), .A(n12162), .B(n12161), .ZN(
        n12164) );
  INV_X1 U13634 ( .A(n12164), .ZN(n12165) );
  INV_X1 U13635 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n12419) );
  OR2_X1 U13636 ( .A1(n10978), .A2(n17253), .ZN(n12168) );
  AOI22_X1 U13637 ( .A1(n14450), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n12167) );
  OAI211_X1 U13638 ( .C1(n14452), .C2(n12419), .A(n12168), .B(n12167), .ZN(
        n15299) );
  NAND2_X1 U13639 ( .A1(n15270), .A2(n15299), .ZN(n14487) );
  INV_X1 U13640 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16767) );
  OR2_X1 U13641 ( .A1(n10978), .A2(n16767), .ZN(n12174) );
  INV_X1 U13642 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n12171) );
  NAND2_X1 U13643 ( .A1(n14450), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n12170) );
  NAND2_X1 U13644 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12169) );
  OAI211_X1 U13645 ( .C1(n12171), .C2(n14452), .A(n12170), .B(n12169), .ZN(
        n12172) );
  INV_X1 U13646 ( .A(n12172), .ZN(n12173) );
  INV_X1 U13647 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18571) );
  OR2_X1 U13648 ( .A1(n10978), .A2(n18571), .ZN(n12180) );
  INV_X1 U13649 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n12177) );
  NAND2_X1 U13650 ( .A1(n14450), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n12176) );
  NAND2_X1 U13651 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12175) );
  OAI211_X1 U13652 ( .C1(n12177), .C2(n14452), .A(n12176), .B(n12175), .ZN(
        n12178) );
  INV_X1 U13653 ( .A(n12178), .ZN(n12179) );
  NAND2_X1 U13654 ( .A1(n12180), .A2(n12179), .ZN(n15408) );
  INV_X1 U13655 ( .A(n10978), .ZN(n14454) );
  INV_X1 U13656 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n16534) );
  NAND2_X1 U13657 ( .A1(n14450), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n12182) );
  NAND2_X1 U13658 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12181) );
  OAI211_X1 U13659 ( .C1(n16534), .C2(n14452), .A(n12182), .B(n12181), .ZN(
        n12183) );
  AOI21_X1 U13660 ( .B1(n14454), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n12183), .ZN(n15419) );
  INV_X1 U13661 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12184) );
  OR2_X1 U13662 ( .A1(n10978), .A2(n12184), .ZN(n12189) );
  INV_X1 U13663 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n16743) );
  NAND2_X1 U13664 ( .A1(n14450), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12186) );
  NAND2_X1 U13665 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12185) );
  OAI211_X1 U13666 ( .C1(n16743), .C2(n14452), .A(n12186), .B(n12185), .ZN(
        n12187) );
  INV_X1 U13667 ( .A(n12187), .ZN(n12188) );
  INV_X1 U13668 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n18405) );
  OR2_X1 U13669 ( .A1(n10978), .A2(n16736), .ZN(n12191) );
  AOI22_X1 U13670 ( .A1(n14450), .A2(P2_EBX_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n12190) );
  OAI211_X1 U13671 ( .C1(n14452), .C2(n18405), .A(n12191), .B(n12190), .ZN(
        n16274) );
  NAND2_X1 U13672 ( .A1(n15500), .A2(n16274), .ZN(n16264) );
  OR2_X1 U13673 ( .A1(n10978), .A2(n16489), .ZN(n12196) );
  INV_X1 U13674 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n18417) );
  NAND2_X1 U13675 ( .A1(n14450), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12193) );
  NAND2_X1 U13676 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n12192) );
  OAI211_X1 U13677 ( .C1(n18417), .C2(n14452), .A(n12193), .B(n12192), .ZN(
        n12194) );
  INV_X1 U13678 ( .A(n12194), .ZN(n12195) );
  OR2_X1 U13679 ( .A1(n10978), .A2(n18596), .ZN(n12201) );
  INV_X1 U13680 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n16483) );
  NAND2_X1 U13681 ( .A1(n14450), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n12198) );
  NAND2_X1 U13682 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n12197) );
  OAI211_X1 U13683 ( .C1(n16483), .C2(n14452), .A(n12198), .B(n12197), .ZN(
        n12199) );
  INV_X1 U13684 ( .A(n12199), .ZN(n12200) );
  INV_X1 U13685 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n18437) );
  INV_X1 U13686 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12202) );
  OR2_X1 U13687 ( .A1(n10978), .A2(n12202), .ZN(n12204) );
  AOI22_X1 U13688 ( .A1(n14450), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n12203) );
  OAI211_X1 U13689 ( .C1(n14452), .C2(n18437), .A(n12204), .B(n12203), .ZN(
        n15562) );
  OR2_X1 U13690 ( .A1(n10978), .A2(n16679), .ZN(n12210) );
  INV_X1 U13691 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n12207) );
  NAND2_X1 U13692 ( .A1(n14450), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12206) );
  NAND2_X1 U13693 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n12205) );
  OAI211_X1 U13694 ( .C1(n12207), .C2(n14452), .A(n12206), .B(n12205), .ZN(
        n12208) );
  INV_X1 U13695 ( .A(n12208), .ZN(n12209) );
  AND2_X1 U13696 ( .A1(n12210), .A2(n12209), .ZN(n16257) );
  INV_X1 U13697 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16666) );
  OR2_X1 U13698 ( .A1(n10978), .A2(n16666), .ZN(n12215) );
  INV_X1 U13699 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n16433) );
  NAND2_X1 U13700 ( .A1(n14450), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12212) );
  NAND2_X1 U13701 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n12211) );
  OAI211_X1 U13702 ( .C1(n16433), .C2(n14452), .A(n12212), .B(n12211), .ZN(
        n12213) );
  INV_X1 U13703 ( .A(n12213), .ZN(n12214) );
  AND2_X1 U13704 ( .A1(n12215), .A2(n12214), .ZN(n16248) );
  INV_X1 U13705 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16659) );
  OR2_X1 U13706 ( .A1(n10978), .A2(n16659), .ZN(n12220) );
  INV_X1 U13707 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n16423) );
  NAND2_X1 U13708 ( .A1(n14450), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n12217) );
  NAND2_X1 U13709 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12216) );
  OAI211_X1 U13710 ( .C1(n16423), .C2(n14452), .A(n12217), .B(n12216), .ZN(
        n12218) );
  INV_X1 U13711 ( .A(n12218), .ZN(n12219) );
  INV_X1 U13712 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n16413) );
  OR2_X1 U13713 ( .A1(n10978), .A2(n11987), .ZN(n12222) );
  AOI22_X1 U13714 ( .A1(n14450), .A2(P2_EBX_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n12221) );
  OAI211_X1 U13715 ( .C1(n12237), .C2(n16413), .A(n12222), .B(n12221), .ZN(
        n16238) );
  NAND2_X1 U13716 ( .A1(n16237), .A2(n16238), .ZN(n16228) );
  OR2_X1 U13717 ( .A1(n10978), .A2(n16637), .ZN(n12227) );
  INV_X1 U13718 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n17334) );
  NAND2_X1 U13719 ( .A1(n14450), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12224) );
  NAND2_X1 U13720 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n12223) );
  OAI211_X1 U13721 ( .C1(n17334), .C2(n14452), .A(n12224), .B(n12223), .ZN(
        n12225) );
  INV_X1 U13722 ( .A(n12225), .ZN(n12226) );
  AND2_X1 U13723 ( .A1(n12227), .A2(n12226), .ZN(n16231) );
  OR2_X1 U13724 ( .A1(n10978), .A2(n16621), .ZN(n12232) );
  INV_X1 U13725 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n17335) );
  NAND2_X1 U13726 ( .A1(n14450), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n12229) );
  NAND2_X1 U13727 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12228) );
  OAI211_X1 U13728 ( .C1(n17335), .C2(n14452), .A(n12229), .B(n12228), .ZN(
        n12230) );
  INV_X1 U13729 ( .A(n12230), .ZN(n12231) );
  INV_X1 U13730 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n18511) );
  INV_X1 U13731 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16381) );
  OR2_X1 U13732 ( .A1(n10978), .A2(n16381), .ZN(n12234) );
  AOI22_X1 U13733 ( .A1(n14450), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n12233) );
  OAI211_X1 U13734 ( .C1(n12237), .C2(n18511), .A(n12234), .B(n12233), .ZN(
        n16217) );
  INV_X1 U13735 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n16372) );
  OR2_X1 U13736 ( .A1(n10978), .A2(n16365), .ZN(n12236) );
  AOI22_X1 U13737 ( .A1(n14450), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n12235) );
  OAI211_X1 U13738 ( .C1(n12237), .C2(n16372), .A(n12236), .B(n12235), .ZN(
        n16207) );
  INV_X1 U13739 ( .A(n14449), .ZN(n12239) );
  NAND2_X1 U13740 ( .A1(n12241), .A2(n19621), .ZN(n12242) );
  NAND2_X1 U13741 ( .A1(n12242), .A2(n11722), .ZN(n12243) );
  INV_X1 U13742 ( .A(n14461), .ZN(n12267) );
  AND3_X1 U13743 ( .A1(n11680), .A2(n19621), .A3(n13849), .ZN(n12245) );
  AND2_X1 U13744 ( .A1(n10961), .A2(n12245), .ZN(n18636) );
  NAND2_X1 U13745 ( .A1(n12279), .A2(n18636), .ZN(n16867) );
  MUX2_X1 U13746 ( .A(n12247), .B(n11680), .S(n12246), .Z(n12258) );
  INV_X1 U13747 ( .A(n12248), .ZN(n12249) );
  NAND3_X1 U13748 ( .A1(n12250), .A2(n11699), .A3(n12249), .ZN(n12256) );
  INV_X1 U13749 ( .A(n12251), .ZN(n14504) );
  OAI21_X1 U13750 ( .B1(n11699), .B2(n12252), .A(n14504), .ZN(n12255) );
  NAND2_X1 U13751 ( .A1(n12254), .A2(n12253), .ZN(n14385) );
  AND3_X1 U13752 ( .A1(n12256), .A2(n12255), .A3(n14385), .ZN(n12257) );
  NAND2_X1 U13753 ( .A1(n12258), .A2(n12257), .ZN(n12262) );
  NAND2_X1 U13754 ( .A1(n12259), .A2(n11774), .ZN(n15174) );
  AOI21_X1 U13755 ( .B1(n15174), .B2(n12260), .A(n11245), .ZN(n12261) );
  NOR2_X1 U13756 ( .A1(n12262), .A2(n12261), .ZN(n16880) );
  INV_X1 U13757 ( .A(n12263), .ZN(n15324) );
  NAND2_X1 U13758 ( .A1(n16880), .A2(n15324), .ZN(n12264) );
  NAND2_X1 U13759 ( .A1(n12279), .A2(n12264), .ZN(n16826) );
  NOR2_X1 U13760 ( .A1(n14682), .A2(n11712), .ZN(n14814) );
  NAND2_X1 U13761 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14814), .ZN(
        n16829) );
  INV_X1 U13762 ( .A(n16829), .ZN(n14668) );
  NOR2_X1 U13763 ( .A1(n18636), .A2(n14668), .ZN(n12265) );
  NOR2_X1 U13764 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n14814), .ZN(
        n15307) );
  NOR2_X1 U13765 ( .A1(n15289), .A2(n15307), .ZN(n15371) );
  AND3_X1 U13766 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n15371), .ZN(n16868) );
  NAND2_X1 U13767 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16868), .ZN(
        n16828) );
  NOR3_X1 U13768 ( .A1(n16837), .A2(n16850), .A3(n16828), .ZN(n12269) );
  NAND2_X1 U13769 ( .A1(n16833), .A2(n12269), .ZN(n18570) );
  NAND2_X1 U13770 ( .A1(n18568), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16694) );
  NOR2_X1 U13771 ( .A1(n18570), .A2(n16694), .ZN(n16757) );
  NAND2_X1 U13772 ( .A1(n16757), .A2(n12271), .ZN(n18597) );
  INV_X1 U13773 ( .A(n16611), .ZN(n16638) );
  AND2_X1 U13774 ( .A1(n16610), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12266) );
  NAND2_X1 U13775 ( .A1(n16638), .A2(n12266), .ZN(n16600) );
  AOI211_X1 U13776 ( .C1(n16365), .C2(n12505), .A(n12267), .B(n16600), .ZN(
        n12507) );
  INV_X1 U13777 ( .A(n12279), .ZN(n12268) );
  NAND2_X1 U13778 ( .A1(n19292), .A2(n17266), .ZN(n17214) );
  NAND2_X1 U13779 ( .A1(n12268), .A2(n18583), .ZN(n16830) );
  OAI21_X1 U13780 ( .B1(n16867), .B2(n12269), .A(n16830), .ZN(n16699) );
  AND2_X1 U13781 ( .A1(n12269), .A2(n14668), .ZN(n16695) );
  NOR2_X1 U13782 ( .A1(n16826), .A2(n16695), .ZN(n12270) );
  OR2_X1 U13783 ( .A1(n16699), .A2(n12270), .ZN(n16724) );
  INV_X1 U13784 ( .A(n16724), .ZN(n16810) );
  NAND2_X1 U13785 ( .A1(n12113), .A2(n12271), .ZN(n12272) );
  NOR2_X1 U13786 ( .A1(n16694), .A2(n12272), .ZN(n16680) );
  NAND3_X1 U13787 ( .A1(n16810), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n16680), .ZN(n12273) );
  NAND2_X1 U13788 ( .A1(n12273), .A2(n16727), .ZN(n16665) );
  INV_X1 U13789 ( .A(n16665), .ZN(n12274) );
  AOI211_X1 U13790 ( .C1(n16655), .C2(n16727), .A(n11987), .B(n12274), .ZN(
        n16642) );
  NAND2_X1 U13791 ( .A1(n16642), .A2(n16610), .ZN(n16612) );
  OAI21_X1 U13792 ( .B1(n16612), .B2(n16381), .A(n16727), .ZN(n16599) );
  OR2_X1 U13793 ( .A1(n18582), .A2(n17336), .ZN(n16358) );
  NAND2_X1 U13794 ( .A1(n11706), .A2(n12055), .ZN(n18641) );
  NAND2_X1 U13795 ( .A1(n18641), .A2(n11774), .ZN(n12277) );
  NAND2_X1 U13796 ( .A1(n10961), .A2(n12276), .ZN(n15317) );
  NAND2_X1 U13797 ( .A1(n12277), .A2(n15317), .ZN(n12278) );
  NAND2_X1 U13798 ( .A1(n12279), .A2(n12278), .ZN(n16871) );
  NAND2_X1 U13799 ( .A1(n12280), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n12284) );
  INV_X1 U13800 ( .A(n15200), .ZN(n14387) );
  NAND2_X1 U13801 ( .A1(n14387), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n12281) );
  OAI211_X1 U13802 ( .C1(n12286), .C2(n14682), .A(n12281), .B(n19233), .ZN(
        n12282) );
  INV_X1 U13803 ( .A(n12282), .ZN(n12283) );
  NAND2_X1 U13804 ( .A1(n12284), .A2(n12283), .ZN(n14650) );
  NAND2_X1 U13805 ( .A1(n12471), .A2(n12285), .ZN(n12290) );
  NAND2_X1 U13806 ( .A1(n12287), .A2(n12288), .ZN(n12299) );
  MUX2_X1 U13807 ( .A(n15200), .B(n19263), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12289) );
  NAND3_X1 U13808 ( .A1(n12290), .A2(n12299), .A3(n12289), .ZN(n14651) );
  INV_X1 U13809 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n17298) );
  INV_X1 U13810 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n17326) );
  OAI222_X1 U13811 ( .A1(n11365), .A2(n17298), .B1(n12479), .B2(n11712), .C1(
        n12420), .C2(n17326), .ZN(n12296) );
  XNOR2_X1 U13812 ( .A(n14653), .B(n12296), .ZN(n14806) );
  INV_X1 U13813 ( .A(n12471), .ZN(n12291) );
  OR2_X1 U13814 ( .A1(n12292), .A2(n12291), .ZN(n12295) );
  NAND2_X1 U13815 ( .A1(n12056), .A2(n15200), .ZN(n12293) );
  MUX2_X1 U13816 ( .A(n12293), .B(n19294), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12294) );
  NAND2_X1 U13817 ( .A1(n12295), .A2(n12294), .ZN(n14807) );
  NOR2_X1 U13818 ( .A1(n14653), .A2(n12296), .ZN(n12297) );
  INV_X1 U13819 ( .A(n12304), .ZN(n12302) );
  NAND2_X1 U13820 ( .A1(n12471), .A2(n12298), .ZN(n12300) );
  OAI211_X1 U13821 ( .C1(n19233), .C2(n19221), .A(n12300), .B(n12299), .ZN(
        n12303) );
  INV_X1 U13822 ( .A(n12303), .ZN(n12301) );
  NAND2_X1 U13823 ( .A1(n12304), .A2(n12303), .ZN(n12305) );
  INV_X2 U13824 ( .A(n11365), .ZN(n13836) );
  AOI22_X1 U13825 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_2__SCAN_IN), .ZN(n12307) );
  NAND2_X1 U13826 ( .A1(n12280), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12306) );
  NAND2_X1 U13827 ( .A1(n12307), .A2(n12306), .ZN(n14661) );
  NAND2_X1 U13828 ( .A1(n12280), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n12312) );
  NAND2_X1 U13829 ( .A1(n12471), .A2(n12308), .ZN(n12311) );
  AOI22_X1 U13830 ( .A1(n13836), .A2(P2_EAX_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12310) );
  NAND2_X1 U13831 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12309) );
  NAND4_X1 U13832 ( .A1(n12312), .A2(n12311), .A3(n12310), .A4(n12309), .ZN(
        n15048) );
  AOI22_X1 U13833 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_4__SCAN_IN), .ZN(n12317) );
  INV_X1 U13834 ( .A(n12313), .ZN(n12314) );
  NAND2_X1 U13835 ( .A1(n12471), .A2(n12314), .ZN(n12316) );
  NAND2_X1 U13836 ( .A1(n12280), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n12315) );
  AOI22_X1 U13837 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_5__SCAN_IN), .ZN(n12322) );
  NAND2_X1 U13838 ( .A1(n12280), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n12321) );
  INV_X1 U13839 ( .A(n12318), .ZN(n12319) );
  NAND2_X1 U13840 ( .A1(n12471), .A2(n12319), .ZN(n12320) );
  NAND3_X1 U13841 ( .A1(n12322), .A2(n12321), .A3(n12320), .ZN(n15483) );
  NAND2_X1 U13842 ( .A1(n15484), .A2(n15483), .ZN(n12326) );
  INV_X1 U13843 ( .A(n12323), .ZN(n12324) );
  NAND2_X1 U13844 ( .A1(n12471), .A2(n12324), .ZN(n12325) );
  AOI22_X1 U13845 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_6__SCAN_IN), .ZN(n12328) );
  NAND2_X1 U13846 ( .A1(n12280), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n12327) );
  NAND2_X1 U13847 ( .A1(n12328), .A2(n12327), .ZN(n16869) );
  NAND2_X1 U13848 ( .A1(n16870), .A2(n16869), .ZN(n12330) );
  NAND2_X1 U13849 ( .A1(n12471), .A2(n14446), .ZN(n12329) );
  AOI22_X1 U13850 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_7__SCAN_IN), .ZN(n12332) );
  NAND2_X1 U13851 ( .A1(n12280), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n12331) );
  NAND2_X1 U13852 ( .A1(n12332), .A2(n12331), .ZN(n16847) );
  AOI22_X1 U13853 ( .A1(n14172), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11480), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12336) );
  AOI22_X1 U13854 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n14230), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12335) );
  AOI22_X1 U13855 ( .A1(n14216), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n14232), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12334) );
  NAND2_X1 U13856 ( .A1(n12385), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12333) );
  AND4_X1 U13857 ( .A1(n12336), .A2(n12335), .A3(n12334), .A4(n12333), .ZN(
        n12347) );
  NAND2_X1 U13858 ( .A1(n14231), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12340) );
  AOI22_X1 U13859 ( .A1(n14222), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n14225), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12339) );
  AOI22_X1 U13860 ( .A1(n14223), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n14224), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12338) );
  NAND2_X1 U13861 ( .A1(n11481), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12337) );
  NAND4_X1 U13862 ( .A1(n12340), .A2(n12339), .A3(n12338), .A4(n12337), .ZN(
        n12345) );
  INV_X1 U13863 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12343) );
  NAND2_X1 U13864 ( .A1(n14215), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12342) );
  NAND2_X1 U13865 ( .A1(n16892), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12341) );
  OAI211_X1 U13866 ( .C1(n12343), .C2(n14219), .A(n12342), .B(n12341), .ZN(
        n12344) );
  NOR2_X1 U13867 ( .A1(n12345), .A2(n12344), .ZN(n12346) );
  NAND2_X1 U13868 ( .A1(n12347), .A2(n12346), .ZN(n14994) );
  AOI22_X1 U13869 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_8__SCAN_IN), .ZN(n12348) );
  OAI21_X1 U13870 ( .B1(n12420), .B2(n12349), .A(n12348), .ZN(n12350) );
  AOI21_X1 U13871 ( .B1(n12471), .B2(n14994), .A(n12350), .ZN(n16840) );
  AOI22_X1 U13872 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n12367) );
  NAND2_X1 U13873 ( .A1(n12280), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n12366) );
  AOI22_X1 U13874 ( .A1(n14172), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11480), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12358) );
  INV_X1 U13875 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12353) );
  NAND2_X1 U13876 ( .A1(n14215), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12352) );
  NAND2_X1 U13877 ( .A1(n14216), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12351) );
  OAI211_X1 U13878 ( .C1(n12353), .C2(n14219), .A(n12352), .B(n12351), .ZN(
        n12354) );
  INV_X1 U13879 ( .A(n12354), .ZN(n12357) );
  AOI22_X1 U13880 ( .A1(n14223), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n14222), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12356) );
  AOI22_X1 U13881 ( .A1(n14224), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14225), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12355) );
  NAND4_X1 U13882 ( .A1(n12358), .A2(n12357), .A3(n12356), .A4(n12355), .ZN(
        n12364) );
  AOI22_X1 U13883 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11481), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12362) );
  AOI22_X1 U13884 ( .A1(n14231), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n14230), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12361) );
  AOI22_X1 U13885 ( .A1(n16892), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14232), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12360) );
  NAND2_X1 U13886 ( .A1(n12385), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12359) );
  NAND4_X1 U13887 ( .A1(n12362), .A2(n12361), .A3(n12360), .A4(n12359), .ZN(
        n12363) );
  NAND2_X1 U13888 ( .A1(n12471), .A2(n11385), .ZN(n12365) );
  NAND3_X1 U13889 ( .A1(n12367), .A2(n12366), .A3(n12365), .ZN(n16807) );
  AOI22_X1 U13890 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_10__SCAN_IN), .ZN(n12384) );
  NAND2_X1 U13891 ( .A1(n12280), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n12383) );
  AOI22_X1 U13892 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11481), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12375) );
  INV_X1 U13893 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12370) );
  NAND2_X1 U13894 ( .A1(n14215), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12369) );
  NAND2_X1 U13895 ( .A1(n16892), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12368) );
  OAI211_X1 U13896 ( .C1(n12370), .C2(n14219), .A(n12369), .B(n12368), .ZN(
        n12371) );
  INV_X1 U13897 ( .A(n12371), .ZN(n12374) );
  AOI22_X1 U13898 ( .A1(n14223), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14222), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12373) );
  AOI22_X1 U13899 ( .A1(n14224), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14225), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12372) );
  NAND4_X1 U13900 ( .A1(n12375), .A2(n12374), .A3(n12373), .A4(n12372), .ZN(
        n12381) );
  AOI22_X1 U13901 ( .A1(n14172), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11480), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12379) );
  AOI22_X1 U13902 ( .A1(n14231), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n14230), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12378) );
  AOI22_X1 U13903 ( .A1(n14216), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14232), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12377) );
  NAND2_X1 U13904 ( .A1(n12385), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12376) );
  NAND4_X1 U13905 ( .A1(n12379), .A2(n12378), .A3(n12377), .A4(n12376), .ZN(
        n12380) );
  NAND2_X1 U13906 ( .A1(n12471), .A2(n10995), .ZN(n12382) );
  NOR2_X2 U13907 ( .A1(n16793), .A2(n16792), .ZN(n16775) );
  AOI22_X1 U13908 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n12403) );
  NAND2_X1 U13909 ( .A1(n12280), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n12402) );
  AOI22_X1 U13910 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11481), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12389) );
  AOI22_X1 U13911 ( .A1(n14231), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n14230), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12388) );
  AOI22_X1 U13912 ( .A1(n16892), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14232), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12387) );
  NAND2_X1 U13913 ( .A1(n12385), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12386) );
  AND4_X1 U13914 ( .A1(n12389), .A2(n12388), .A3(n12387), .A4(n12386), .ZN(
        n12400) );
  AOI22_X1 U13915 ( .A1(n14223), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14222), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12393) );
  NAND2_X1 U13916 ( .A1(n14172), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12392) );
  AOI22_X1 U13917 ( .A1(n14224), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14225), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12391) );
  NAND2_X1 U13918 ( .A1(n11480), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12390) );
  NAND4_X1 U13919 ( .A1(n12393), .A2(n12392), .A3(n12391), .A4(n12390), .ZN(
        n12398) );
  NAND2_X1 U13920 ( .A1(n14215), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12395) );
  NAND2_X1 U13921 ( .A1(n14216), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n12394) );
  OAI211_X1 U13922 ( .C1(n12396), .C2(n14219), .A(n12395), .B(n12394), .ZN(
        n12397) );
  NOR2_X1 U13923 ( .A1(n12398), .A2(n12397), .ZN(n12399) );
  NAND2_X1 U13924 ( .A1(n12400), .A2(n12399), .ZN(n15267) );
  NAND2_X1 U13925 ( .A1(n12471), .A2(n15267), .ZN(n12401) );
  NAND3_X1 U13926 ( .A1(n12403), .A2(n12402), .A3(n12401), .ZN(n16776) );
  NAND2_X1 U13927 ( .A1(n16775), .A2(n16776), .ZN(n16777) );
  INV_X1 U13928 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12406) );
  NAND2_X1 U13929 ( .A1(n14215), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12405) );
  NAND2_X1 U13930 ( .A1(n16892), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12404) );
  OAI211_X1 U13931 ( .C1(n12406), .C2(n14219), .A(n12405), .B(n12404), .ZN(
        n12407) );
  INV_X1 U13932 ( .A(n12407), .ZN(n12411) );
  AOI22_X1 U13933 ( .A1(n14172), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n14230), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12410) );
  AOI22_X1 U13934 ( .A1(n14223), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n14224), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12409) );
  AOI22_X1 U13935 ( .A1(n14222), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n14225), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12408) );
  NAND4_X1 U13936 ( .A1(n12411), .A2(n12410), .A3(n12409), .A4(n12408), .ZN(
        n12417) );
  AOI22_X1 U13937 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14231), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12415) );
  AOI22_X1 U13938 ( .A1(n11480), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11481), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12414) );
  AOI22_X1 U13939 ( .A1(n14216), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n14232), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12413) );
  NAND2_X1 U13940 ( .A1(n14233), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12412) );
  NAND4_X1 U13941 ( .A1(n12415), .A2(n12414), .A3(n12413), .A4(n12412), .ZN(
        n12416) );
  OR2_X1 U13942 ( .A1(n12417), .A2(n12416), .ZN(n15301) );
  AOI22_X1 U13943 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_12__SCAN_IN), .ZN(n12418) );
  OAI21_X1 U13944 ( .B1(n12420), .B2(n12419), .A(n12418), .ZN(n12421) );
  AOI21_X1 U13945 ( .B1(n12471), .B2(n15301), .A(n12421), .ZN(n18359) );
  AOI22_X1 U13946 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_13__SCAN_IN), .ZN(n12438) );
  NAND2_X1 U13947 ( .A1(n12280), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n12437) );
  AOI22_X1 U13948 ( .A1(n14172), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11480), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12429) );
  NAND2_X1 U13949 ( .A1(n14215), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12423) );
  NAND2_X1 U13950 ( .A1(n14216), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n12422) );
  OAI211_X1 U13951 ( .C1(n12424), .C2(n14219), .A(n12423), .B(n12422), .ZN(
        n12425) );
  INV_X1 U13952 ( .A(n12425), .ZN(n12428) );
  AOI22_X1 U13953 ( .A1(n14223), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n14222), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12427) );
  AOI22_X1 U13954 ( .A1(n14224), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14225), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12426) );
  NAND4_X1 U13955 ( .A1(n12429), .A2(n12428), .A3(n12427), .A4(n12426), .ZN(
        n12435) );
  AOI22_X1 U13956 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11481), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12433) );
  AOI22_X1 U13957 ( .A1(n14231), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14230), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12432) );
  AOI22_X1 U13958 ( .A1(n16892), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14232), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12431) );
  NAND2_X1 U13959 ( .A1(n14233), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12430) );
  NAND4_X1 U13960 ( .A1(n12433), .A2(n12432), .A3(n12431), .A4(n12430), .ZN(
        n12434) );
  OR2_X1 U13961 ( .A1(n12435), .A2(n12434), .ZN(n15339) );
  NAND2_X1 U13962 ( .A1(n12471), .A2(n15339), .ZN(n12436) );
  NAND3_X1 U13963 ( .A1(n12438), .A2(n12437), .A3(n12436), .ZN(n14486) );
  AOI22_X1 U13964 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n12455) );
  AOI22_X1 U13965 ( .A1(n14172), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n14231), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12442) );
  AOI22_X1 U13966 ( .A1(n11480), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14230), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12441) );
  AOI22_X1 U13967 ( .A1(n14216), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n16892), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12440) );
  NAND2_X1 U13968 ( .A1(n14233), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12439) );
  NAND4_X1 U13969 ( .A1(n12442), .A2(n12441), .A3(n12440), .A4(n12439), .ZN(
        n12452) );
  AOI22_X1 U13970 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11481), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12450) );
  NAND2_X1 U13971 ( .A1(n14215), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n12444) );
  NAND2_X1 U13972 ( .A1(n14232), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n12443) );
  OAI211_X1 U13973 ( .C1(n12445), .C2(n14219), .A(n12444), .B(n12443), .ZN(
        n12446) );
  INV_X1 U13974 ( .A(n12446), .ZN(n12449) );
  AOI22_X1 U13975 ( .A1(n14223), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14224), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12448) );
  AOI22_X1 U13976 ( .A1(n14222), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n14225), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12447) );
  NAND4_X1 U13977 ( .A1(n12450), .A2(n12449), .A3(n12448), .A4(n12447), .ZN(
        n12451) );
  NOR2_X1 U13978 ( .A1(n12452), .A2(n12451), .ZN(n15410) );
  INV_X1 U13979 ( .A(n15410), .ZN(n15411) );
  NAND2_X1 U13980 ( .A1(n12471), .A2(n15411), .ZN(n12454) );
  NAND2_X1 U13981 ( .A1(n12280), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n12453) );
  AOI22_X1 U13982 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_15__SCAN_IN), .ZN(n12474) );
  NAND2_X1 U13983 ( .A1(n12280), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n12473) );
  AOI22_X1 U13984 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11481), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12459) );
  AOI22_X1 U13985 ( .A1(n14231), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n14230), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12458) );
  AOI22_X1 U13986 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n16892), .B1(
        n14232), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12457) );
  NAND2_X1 U13987 ( .A1(n14233), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12456) );
  AND4_X1 U13988 ( .A1(n12459), .A2(n12458), .A3(n12457), .A4(n12456), .ZN(
        n12470) );
  AOI22_X1 U13989 ( .A1(n14223), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n14222), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12463) );
  NAND2_X1 U13990 ( .A1(n14172), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12462) );
  AOI22_X1 U13991 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n14224), .B1(
        n14225), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12461) );
  NAND2_X1 U13992 ( .A1(n11480), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12460) );
  NAND4_X1 U13993 ( .A1(n12463), .A2(n12462), .A3(n12461), .A4(n12460), .ZN(
        n12468) );
  INV_X1 U13994 ( .A(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12466) );
  NAND2_X1 U13995 ( .A1(n14215), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12465) );
  NAND2_X1 U13996 ( .A1(n14216), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n12464) );
  OAI211_X1 U13997 ( .C1(n12466), .C2(n14219), .A(n12465), .B(n12464), .ZN(
        n12467) );
  NOR2_X1 U13998 ( .A1(n12468), .A2(n12467), .ZN(n12469) );
  NAND2_X1 U13999 ( .A1(n12470), .A2(n12469), .ZN(n15417) );
  NAND2_X1 U14000 ( .A1(n12471), .A2(n15417), .ZN(n12472) );
  AOI22_X1 U14001 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_16__SCAN_IN), .ZN(n12476) );
  NAND2_X1 U14002 ( .A1(n12280), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n12475) );
  AOI22_X1 U14003 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_17__SCAN_IN), .ZN(n12478) );
  NAND2_X1 U14004 ( .A1(n12280), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n12477) );
  NAND2_X1 U14005 ( .A1(n12478), .A2(n12477), .ZN(n16348) );
  NAND2_X1 U14006 ( .A1(n16347), .A2(n16348), .ZN(n16339) );
  AOI22_X1 U14007 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_18__SCAN_IN), .ZN(n12481) );
  NAND2_X1 U14008 ( .A1(n12280), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n12480) );
  NOR2_X2 U14009 ( .A1(n16339), .A2(n16340), .ZN(n15507) );
  AOI22_X1 U14010 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_19__SCAN_IN), .ZN(n12483) );
  NAND2_X1 U14011 ( .A1(n12280), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n12482) );
  NAND2_X1 U14012 ( .A1(n12483), .A2(n12482), .ZN(n15509) );
  AND2_X2 U14013 ( .A1(n15507), .A2(n15509), .ZN(n16691) );
  AOI22_X1 U14014 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n12485) );
  NAND2_X1 U14015 ( .A1(n12280), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n12484) );
  NAND2_X1 U14016 ( .A1(n12485), .A2(n12484), .ZN(n16692) );
  AOI22_X1 U14017 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n12487) );
  NAND2_X1 U14018 ( .A1(n12280), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n12486) );
  NAND2_X1 U14019 ( .A1(n12487), .A2(n12486), .ZN(n15551) );
  AOI222_X1 U14020 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n12280), .B1(n12488), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C1(n13836), .C2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16670) );
  AOI22_X1 U14021 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n12490) );
  NAND2_X1 U14022 ( .A1(n12280), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n12489) );
  NAND2_X1 U14023 ( .A1(n12490), .A2(n12489), .ZN(n16330) );
  AOI22_X1 U14024 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n12492) );
  NAND2_X1 U14025 ( .A1(n12280), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12491) );
  AND2_X1 U14026 ( .A1(n12492), .A2(n12491), .ZN(n16323) );
  AOI22_X1 U14027 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n12494) );
  NAND2_X1 U14028 ( .A1(n12280), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12493) );
  NAND2_X1 U14029 ( .A1(n12494), .A2(n12493), .ZN(n16315) );
  AOI22_X1 U14030 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n12496) );
  NAND2_X1 U14031 ( .A1(n12280), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n12495) );
  NAND2_X1 U14032 ( .A1(n12496), .A2(n12495), .ZN(n16308) );
  NAND2_X1 U14033 ( .A1(n16309), .A2(n16308), .ZN(n16298) );
  AOI22_X1 U14034 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n12498) );
  NAND2_X1 U14035 ( .A1(n12280), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12497) );
  AND2_X1 U14036 ( .A1(n12498), .A2(n12497), .ZN(n16299) );
  AOI22_X1 U14037 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n12500) );
  NAND2_X1 U14038 ( .A1(n12280), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12499) );
  AND2_X1 U14039 ( .A1(n12500), .A2(n12499), .ZN(n16292) );
  AOI22_X1 U14040 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n12502) );
  NAND2_X1 U14041 ( .A1(n12280), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n12501) );
  AND2_X1 U14042 ( .A1(n12502), .A2(n12501), .ZN(n13835) );
  INV_X1 U14043 ( .A(n13835), .ZN(n12503) );
  XNOR2_X1 U14044 ( .A(n16290), .B(n12503), .ZN(n18540) );
  NAND2_X1 U14045 ( .A1(n18601), .A2(n18540), .ZN(n12504) );
  OAI211_X1 U14046 ( .C1(n16599), .C2(n12505), .A(n16358), .B(n12504), .ZN(
        n12506) );
  NAND2_X1 U14047 ( .A1(n11030), .A2(n12511), .ZN(P2_U3017) );
  INV_X1 U14048 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12512) );
  AND2_X2 U14049 ( .A1(n12519), .A2(n12520), .ZN(n12759) );
  INV_X2 U14050 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12513) );
  NOR2_X4 U14051 ( .A1(n12513), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12518) );
  AOI22_X1 U14053 ( .A1(n12759), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12658), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12517) );
  AOI22_X1 U14054 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12729), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12516) );
  AND2_X4 U14055 ( .A1(n12513), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14749) );
  AOI22_X1 U14057 ( .A1(n12736), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12735), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12515) );
  AND2_X4 U14058 ( .A1(n12518), .A2(n12519), .ZN(n12727) );
  AOI22_X1 U14059 ( .A1(n12727), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12696), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12514) );
  NAND4_X1 U14060 ( .A1(n12517), .A2(n12516), .A3(n12515), .A4(n12514), .ZN(
        n12526) );
  AND2_X4 U14061 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14730) );
  AND2_X2 U14062 ( .A1(n14749), .A2(n14730), .ZN(n12760) );
  AND2_X2 U14063 ( .A1(n14749), .A2(n14900), .ZN(n12734) );
  AOI22_X1 U14064 ( .A1(n12760), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12734), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12524) );
  AOI22_X1 U14065 ( .A1(n12737), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12690), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12523) );
  AOI22_X1 U14066 ( .A1(n12659), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12653), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12522) );
  AOI22_X1 U14067 ( .A1(n12761), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12521) );
  NAND4_X1 U14068 ( .A1(n12524), .A2(n12523), .A3(n12522), .A4(n12521), .ZN(
        n12525) );
  AOI22_X1 U14069 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13260), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12530) );
  AOI22_X1 U14070 ( .A1(n12659), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12727), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12529) );
  AOI22_X1 U14071 ( .A1(n12735), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12696), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12528) );
  AOI22_X1 U14072 ( .A1(n12736), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12653), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12527) );
  AOI22_X1 U14073 ( .A1(n12760), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12658), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12534) );
  AOI22_X1 U14074 ( .A1(n12734), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12759), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12533) );
  AOI22_X1 U14075 ( .A1(n12737), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12690), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12532) );
  AOI22_X1 U14076 ( .A1(n12761), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12774), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12531) );
  AOI22_X1 U14077 ( .A1(n12659), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10984), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12539) );
  AOI22_X1 U14078 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12729), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12538) );
  AOI22_X1 U14079 ( .A1(n12735), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12696), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12537) );
  AOI22_X1 U14080 ( .A1(n12736), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12653), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12536) );
  AOI22_X1 U14081 ( .A1(n12760), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12658), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12543) );
  AOI22_X1 U14082 ( .A1(n12734), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12759), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12542) );
  AOI22_X1 U14083 ( .A1(n12737), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12690), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12541) );
  INV_X2 U14084 ( .A(n12621), .ZN(n14871) );
  AOI22_X1 U14085 ( .A1(n12760), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12734), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12548) );
  AOI22_X1 U14086 ( .A1(n12727), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12735), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12547) );
  AOI22_X1 U14087 ( .A1(n12737), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12774), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12546) );
  AOI22_X1 U14088 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12761), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12545) );
  NAND4_X1 U14089 ( .A1(n12548), .A2(n12547), .A3(n12546), .A4(n12545), .ZN(
        n12554) );
  AOI22_X1 U14090 ( .A1(n12759), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12658), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12552) );
  AOI22_X1 U14091 ( .A1(n12659), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12696), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12551) );
  AOI22_X1 U14092 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12690), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12550) );
  AOI22_X1 U14093 ( .A1(n12736), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12653), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12549) );
  NAND4_X1 U14094 ( .A1(n12552), .A2(n12551), .A3(n12550), .A4(n12549), .ZN(
        n12553) );
  AOI22_X1 U14095 ( .A1(n12760), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12658), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12558) );
  AOI22_X1 U14096 ( .A1(n12734), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12759), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12557) );
  AOI22_X1 U14097 ( .A1(n12737), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12690), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12556) );
  AOI22_X1 U14098 ( .A1(n12761), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10981), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12555) );
  AOI22_X1 U14099 ( .A1(n12736), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12653), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12561) );
  AOI22_X1 U14100 ( .A1(n12735), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12696), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12560) );
  AOI22_X1 U14101 ( .A1(n12659), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10983), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12559) );
  AOI22_X1 U14102 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12729), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12562) );
  NAND3_X2 U14103 ( .A1(n12563), .A2(n11387), .A3(n12562), .ZN(n22148) );
  AOI22_X1 U14104 ( .A1(n12760), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12759), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12567) );
  AOI22_X1 U14105 ( .A1(n12659), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12729), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12566) );
  AOI22_X1 U14106 ( .A1(n12735), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12696), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12565) );
  AOI22_X1 U14107 ( .A1(n12736), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12653), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12564) );
  AOI22_X1 U14108 ( .A1(n12734), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12658), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12571) );
  AOI22_X1 U14109 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10984), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12570) );
  AOI22_X1 U14110 ( .A1(n12737), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12690), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12569) );
  AOI22_X1 U14111 ( .A1(n12761), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12774), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12568) );
  NAND2_X2 U14112 ( .A1(n11388), .A2(n11023), .ZN(n14948) );
  AND2_X1 U14113 ( .A1(n12639), .A2(n14948), .ZN(n12572) );
  INV_X1 U14114 ( .A(n14846), .ZN(n14702) );
  NAND2_X1 U14115 ( .A1(n12760), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12576) );
  NAND2_X1 U14116 ( .A1(n12734), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12575) );
  NAND2_X1 U14117 ( .A1(n12759), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12574) );
  NAND2_X1 U14118 ( .A1(n12658), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12573) );
  NAND2_X1 U14119 ( .A1(n12727), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12580) );
  NAND2_X1 U14120 ( .A1(n12659), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12579) );
  NAND2_X1 U14121 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12578) );
  NAND2_X1 U14122 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n12577) );
  NAND2_X1 U14123 ( .A1(n12735), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n12584) );
  NAND2_X1 U14124 ( .A1(n12736), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12583) );
  NAND2_X1 U14125 ( .A1(n12696), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12582) );
  NAND2_X1 U14126 ( .A1(n12653), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n12581) );
  NAND2_X1 U14127 ( .A1(n12737), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12588) );
  NAND2_X1 U14128 ( .A1(n12690), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12587) );
  NAND2_X1 U14129 ( .A1(n12761), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12586) );
  NAND2_X1 U14130 ( .A1(n12774), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12585) );
  NAND4_X4 U14131 ( .A1(n12592), .A2(n12591), .A3(n12590), .A4(n12589), .ZN(
        n15124) );
  NAND2_X1 U14132 ( .A1(n14702), .A2(n15124), .ZN(n14546) );
  INV_X1 U14133 ( .A(n14546), .ZN(n12614) );
  NAND2_X1 U14134 ( .A1(n12760), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n12596) );
  NAND2_X1 U14135 ( .A1(n12734), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12595) );
  NAND2_X1 U14136 ( .A1(n12759), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n12594) );
  NAND2_X1 U14137 ( .A1(n12658), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12593) );
  NAND2_X1 U14138 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12600) );
  NAND2_X1 U14139 ( .A1(n12659), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12599) );
  NAND2_X1 U14140 ( .A1(n12727), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12598) );
  NAND2_X1 U14141 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n12597) );
  NAND2_X1 U14142 ( .A1(n12735), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n12604) );
  NAND2_X1 U14143 ( .A1(n12736), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12603) );
  NAND2_X1 U14144 ( .A1(n12696), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12602) );
  NAND2_X1 U14145 ( .A1(n12653), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n12601) );
  NAND2_X1 U14146 ( .A1(n12737), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12608) );
  NAND2_X1 U14147 ( .A1(n12690), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12607) );
  NAND2_X1 U14148 ( .A1(n12761), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12606) );
  NAND2_X1 U14149 ( .A1(n12774), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12605) );
  INV_X1 U14150 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n12613) );
  XNOR2_X1 U14151 ( .A(n12613), .B(P1_STATE_REG_1__SCAN_IN), .ZN(n13633) );
  NAND2_X1 U14152 ( .A1(n12614), .A2(n11372), .ZN(n12617) );
  NAND2_X1 U14153 ( .A1(n22148), .A2(n14948), .ZN(n14844) );
  AND2_X1 U14154 ( .A1(n22148), .A2(n15596), .ZN(n12615) );
  INV_X2 U14155 ( .A(n14850), .ZN(n15151) );
  NOR2_X1 U14156 ( .A1(n14717), .A2(n15124), .ZN(n12616) );
  NAND3_X1 U14157 ( .A1(n15093), .A2(n12627), .A3(n15156), .ZN(n14725) );
  NAND2_X1 U14158 ( .A1(n15156), .A2(n22148), .ZN(n12620) );
  NAND2_X1 U14159 ( .A1(n13650), .A2(n15245), .ZN(n12622) );
  INV_X1 U14160 ( .A(n12618), .ZN(n14703) );
  NAND2_X1 U14161 ( .A1(n12622), .A2(n14800), .ZN(n12625) );
  INV_X1 U14162 ( .A(n12627), .ZN(n12628) );
  INV_X1 U14163 ( .A(n12648), .ZN(n12718) );
  NAND2_X1 U14164 ( .A1(n12718), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12634) );
  NAND2_X1 U14165 ( .A1(n16973), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16943) );
  INV_X1 U14166 ( .A(n16943), .ZN(n12633) );
  NAND2_X1 U14167 ( .A1(n15582), .A2(n16946), .ZN(n13654) );
  MUX2_X1 U14168 ( .A(n12633), .B(n13654), .S(n21915), .Z(n12707) );
  INV_X1 U14169 ( .A(n12635), .ZN(n12636) );
  OAI21_X1 U14170 ( .B1(n15093), .B2(n12637), .A(n12636), .ZN(n12645) );
  NAND3_X1 U14171 ( .A1(n14705), .A2(n12623), .A3(n15577), .ZN(n12644) );
  INV_X1 U14172 ( .A(n12638), .ZN(n12643) );
  NAND2_X1 U14173 ( .A1(n12627), .A2(n12639), .ZN(n14865) );
  NAND2_X1 U14174 ( .A1(n15582), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12640) );
  AOI21_X1 U14175 ( .B1(n14850), .B2(n15124), .A(n12640), .ZN(n12641) );
  AND2_X1 U14176 ( .A1(n14865), .A2(n12641), .ZN(n12642) );
  NAND4_X1 U14177 ( .A1(n12645), .A2(n12644), .A3(n12643), .A4(n12642), .ZN(
        n12827) );
  XNOR2_X1 U14178 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21903) );
  NAND2_X1 U14179 ( .A1(n16943), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n12714) );
  OAI21_X1 U14180 ( .B1(n13654), .B2(n21903), .A(n12714), .ZN(n12646) );
  INV_X1 U14181 ( .A(n12646), .ZN(n12647) );
  OAI21_X2 U14182 ( .B1(n12648), .B2(n16161), .A(n12647), .ZN(n12649) );
  NAND2_X1 U14183 ( .A1(n14906), .A2(n16946), .ZN(n12668) );
  AOI22_X1 U14184 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12727), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12657) );
  BUF_X1 U14185 ( .A(n12734), .Z(n12688) );
  AOI22_X1 U14186 ( .A1(n12688), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12679), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12656) );
  AOI22_X1 U14187 ( .A1(n12678), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12774), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12655) );
  AOI22_X1 U14188 ( .A1(n12671), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12654) );
  NAND4_X1 U14189 ( .A1(n12657), .A2(n12656), .A3(n12655), .A4(n12654), .ZN(
        n12665) );
  AOI22_X1 U14190 ( .A1(n12689), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12663) );
  AOI22_X1 U14191 ( .A1(n12670), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12728), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12662) );
  BUF_X1 U14192 ( .A(n12759), .Z(n12695) );
  AOI22_X1 U14193 ( .A1(n12695), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12661) );
  AOI22_X1 U14194 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12672), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12660) );
  NAND4_X1 U14195 ( .A1(n12663), .A2(n12662), .A3(n12661), .A4(n12660), .ZN(
        n12664) );
  NAND2_X1 U14196 ( .A1(n15245), .A2(n13667), .ZN(n12666) );
  NAND2_X2 U14197 ( .A1(n12668), .A2(n12667), .ZN(n13666) );
  INV_X1 U14198 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12687) );
  NOR2_X1 U14199 ( .A1(n14871), .A2(n16946), .ZN(n12708) );
  AOI22_X1 U14200 ( .A1(n12688), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12658), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12677) );
  AOI22_X1 U14201 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12727), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12676) );
  BUF_X1 U14203 ( .A(n12735), .Z(n12670) );
  AOI22_X1 U14204 ( .A1(n12736), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12670), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12675) );
  AOI22_X1 U14206 ( .A1(n12673), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12672), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12674) );
  NAND4_X1 U14207 ( .A1(n12677), .A2(n12676), .A3(n12675), .A4(n12674), .ZN(
        n12685) );
  AOI22_X1 U14208 ( .A1(n12689), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12695), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12683) );
  BUF_X1 U14209 ( .A(n12729), .Z(n12678) );
  AOI22_X1 U14210 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12678), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12682) );
  AOI22_X1 U14211 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12774), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12681) );
  AOI22_X1 U14212 ( .A1(n12728), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12680) );
  NAND4_X1 U14213 ( .A1(n12683), .A2(n12682), .A3(n12681), .A4(n12680), .ZN(
        n12684) );
  NAND2_X1 U14214 ( .A1(n12708), .A2(n12808), .ZN(n12710) );
  NAND3_X1 U14215 ( .A1(n14719), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n13667), 
        .ZN(n12686) );
  NAND2_X1 U14216 ( .A1(n13341), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12706) );
  BUF_X1 U14217 ( .A(n12760), .Z(n12689) );
  AOI22_X1 U14218 ( .A1(n12689), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12688), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12694) );
  AOI22_X1 U14219 ( .A1(n12727), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12671), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12693) );
  AOI22_X1 U14220 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12692) );
  AOI22_X1 U14221 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12774), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12691) );
  NAND4_X1 U14222 ( .A1(n12694), .A2(n12693), .A3(n12692), .A4(n12691), .ZN(
        n12702) );
  AOI22_X1 U14223 ( .A1(n12695), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12658), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12700) );
  AOI22_X1 U14224 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12728), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12699) );
  AOI22_X1 U14225 ( .A1(n12678), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12672), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12698) );
  AOI22_X1 U14226 ( .A1(n12670), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12697) );
  NAND4_X1 U14227 ( .A1(n12700), .A2(n12699), .A3(n12698), .A4(n12697), .ZN(
        n12701) );
  NAND2_X1 U14228 ( .A1(n14719), .A2(n13675), .ZN(n12703) );
  OAI211_X1 U14229 ( .C1(n12808), .C2(n14871), .A(P1_STATE2_REG_0__SCAN_IN), 
        .B(n12703), .ZN(n12704) );
  INV_X1 U14230 ( .A(n12704), .ZN(n12705) );
  NAND2_X1 U14231 ( .A1(n12706), .A2(n12705), .ZN(n12836) );
  NAND2_X1 U14232 ( .A1(n12707), .A2(n16946), .ZN(n12712) );
  NAND2_X1 U14233 ( .A1(n12708), .A2(n13737), .ZN(n13733) );
  INV_X1 U14234 ( .A(n13675), .ZN(n12709) );
  MUX2_X1 U14235 ( .A(n12710), .B(n13733), .S(n12709), .Z(n12711) );
  NAND2_X1 U14236 ( .A1(n12712), .A2(n12711), .ZN(n12835) );
  INV_X1 U14237 ( .A(n13733), .ZN(n12713) );
  AND2_X1 U14238 ( .A1(n12714), .A2(n16161), .ZN(n12715) );
  NAND2_X1 U14239 ( .A1(n12718), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12723) );
  INV_X1 U14240 ( .A(n13654), .ZN(n12752) );
  INV_X1 U14241 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21900) );
  NAND2_X1 U14242 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12719) );
  NAND2_X1 U14243 ( .A1(n21900), .A2(n12719), .ZN(n12721) );
  NAND2_X1 U14244 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21932) );
  INV_X1 U14245 ( .A(n21932), .ZN(n12720) );
  NAND2_X1 U14246 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n12720), .ZN(
        n12750) );
  AND2_X1 U14247 ( .A1(n12721), .A2(n12750), .ZN(n21772) );
  AOI22_X1 U14248 ( .A1(n12752), .A2(n21772), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16943), .ZN(n12722) );
  INV_X1 U14249 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12744) );
  AOI22_X1 U14250 ( .A1(n12689), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12733) );
  AOI22_X1 U14251 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n13279), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12732) );
  AOI22_X1 U14252 ( .A1(n12727), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12728), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12731) );
  AOI22_X1 U14253 ( .A1(n12678), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12730) );
  NAND4_X1 U14254 ( .A1(n12733), .A2(n12732), .A3(n12731), .A4(n12730), .ZN(
        n12743) );
  AOI22_X1 U14255 ( .A1(n12688), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12695), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12741) );
  AOI22_X1 U14256 ( .A1(n12670), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12672), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12740) );
  AOI22_X1 U14257 ( .A1(n12671), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12739) );
  AOI22_X1 U14258 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12774), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12738) );
  NAND4_X1 U14259 ( .A1(n12741), .A2(n12740), .A3(n12739), .A4(n12738), .ZN(
        n12742) );
  NOR2_X1 U14260 ( .A1(n12743), .A2(n12742), .ZN(n13662) );
  OAI22_X1 U14261 ( .A1(n13314), .A2(n12744), .B1(n13345), .B2(n13662), .ZN(
        n12745) );
  INV_X1 U14262 ( .A(n12747), .ZN(n12748) );
  NAND2_X1 U14263 ( .A1(n13666), .A2(n12748), .ZN(n12814) );
  NAND2_X2 U14264 ( .A1(n12815), .A2(n12749), .ZN(n12846) );
  NAND2_X1 U14265 ( .A1(n12718), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12754) );
  INV_X1 U14266 ( .A(n12750), .ZN(n15117) );
  NAND2_X1 U14267 ( .A1(n15117), .A2(n21933), .ZN(n21852) );
  NAND2_X1 U14268 ( .A1(n12750), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12751) );
  NAND2_X1 U14269 ( .A1(n21852), .A2(n12751), .ZN(n21904) );
  AOI22_X1 U14270 ( .A1(n12752), .A2(n21904), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n16943), .ZN(n12753) );
  AOI22_X1 U14271 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12678), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12758) );
  AOI22_X1 U14272 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12727), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12757) );
  AOI22_X1 U14273 ( .A1(n12670), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12728), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12756) );
  AOI22_X1 U14274 ( .A1(n12671), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12755) );
  NAND4_X1 U14275 ( .A1(n12758), .A2(n12757), .A3(n12756), .A4(n12755), .ZN(
        n12767) );
  AOI22_X1 U14276 ( .A1(n12688), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12695), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12765) );
  AOI22_X1 U14277 ( .A1(n12689), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12764) );
  AOI22_X1 U14278 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12763) );
  AOI22_X1 U14279 ( .A1(n12672), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12774), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12762) );
  NAND4_X1 U14280 ( .A1(n12765), .A2(n12764), .A3(n12763), .A4(n12762), .ZN(
        n12766) );
  AOI22_X1 U14281 ( .A1(n13341), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13333), .B2(n13688), .ZN(n12768) );
  NAND2_X1 U14282 ( .A1(n13341), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12782) );
  AOI22_X1 U14283 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12695), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12773) );
  AOI22_X1 U14284 ( .A1(n10984), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12670), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12772) );
  AOI22_X1 U14285 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12678), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12771) );
  AOI22_X1 U14286 ( .A1(n12671), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12770) );
  NAND4_X1 U14287 ( .A1(n12773), .A2(n12772), .A3(n12771), .A4(n12770), .ZN(
        n12780) );
  AOI22_X1 U14288 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12688), .B1(
        n12689), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12778) );
  AOI22_X1 U14289 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12728), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12777) );
  AOI22_X1 U14290 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12679), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12776) );
  AOI22_X1 U14291 ( .A1(n12672), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12774), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12775) );
  NAND4_X1 U14292 ( .A1(n12778), .A2(n12777), .A3(n12776), .A4(n12775), .ZN(
        n12779) );
  NAND2_X1 U14293 ( .A1(n13333), .A2(n13703), .ZN(n12781) );
  NAND2_X1 U14294 ( .A1(n12782), .A2(n12781), .ZN(n12856) );
  NAND2_X1 U14295 ( .A1(n13341), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12794) );
  AOI22_X1 U14296 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12678), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12786) );
  AOI22_X1 U14297 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12727), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12785) );
  AOI22_X1 U14298 ( .A1(n12670), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12728), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12784) );
  AOI22_X1 U14299 ( .A1(n12671), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12783) );
  NAND4_X1 U14300 ( .A1(n12786), .A2(n12785), .A3(n12784), .A4(n12783), .ZN(
        n12792) );
  AOI22_X1 U14301 ( .A1(n12688), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12695), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12790) );
  AOI22_X1 U14302 ( .A1(n12689), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12789) );
  AOI22_X1 U14303 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12788) );
  AOI22_X1 U14304 ( .A1(n12672), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12774), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12787) );
  NAND4_X1 U14305 ( .A1(n12790), .A2(n12789), .A3(n12788), .A4(n12787), .ZN(
        n12791) );
  NAND2_X1 U14306 ( .A1(n13333), .A2(n13706), .ZN(n12793) );
  NAND2_X1 U14307 ( .A1(n12794), .A2(n12793), .ZN(n12871) );
  NAND2_X1 U14308 ( .A1(n13341), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12807) );
  AOI22_X1 U14309 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n13279), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12799) );
  AOI22_X1 U14310 ( .A1(n12689), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12798) );
  AOI22_X1 U14311 ( .A1(n12695), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12672), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12797) );
  AOI22_X1 U14312 ( .A1(n12728), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12796) );
  NAND4_X1 U14313 ( .A1(n12799), .A2(n12798), .A3(n12797), .A4(n12796), .ZN(
        n12805) );
  AOI22_X1 U14314 ( .A1(n12671), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12670), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12803) );
  AOI22_X1 U14315 ( .A1(n10984), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12678), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12802) );
  AOI22_X1 U14316 ( .A1(n12688), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12801) );
  AOI22_X1 U14317 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12774), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12800) );
  NAND4_X1 U14318 ( .A1(n12803), .A2(n12802), .A3(n12801), .A4(n12800), .ZN(
        n12804) );
  NAND2_X1 U14319 ( .A1(n13333), .A2(n13723), .ZN(n12806) );
  INV_X1 U14320 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12809) );
  OAI22_X1 U14321 ( .A1(n13314), .A2(n12809), .B1(n13345), .B2(n12808), .ZN(
        n12810) );
  NAND2_X1 U14322 ( .A1(n12639), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12978) );
  INV_X2 U14323 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n21917) );
  INV_X1 U14324 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n15264) );
  NOR2_X1 U14325 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13272) );
  INV_X1 U14326 ( .A(n12849), .ZN(n12811) );
  OAI21_X1 U14327 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n12880), .A(
        n12903), .ZN(n21478) );
  AOI22_X1 U14328 ( .A1(n13522), .A2(n21478), .B1(n13303), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12812) );
  OAI21_X1 U14329 ( .B1(n13232), .B2(n15264), .A(n12812), .ZN(n12813) );
  AOI21_X1 U14330 ( .B1(n13721), .B2(n14820), .A(n12813), .ZN(n15261) );
  NAND2_X1 U14331 ( .A1(n12815), .A2(n12814), .ZN(n12818) );
  INV_X1 U14332 ( .A(n12816), .ZN(n12817) );
  NAND2_X1 U14333 ( .A1(n12818), .A2(n12817), .ZN(n12819) );
  INV_X1 U14334 ( .A(n14844), .ZN(n13373) );
  NAND2_X1 U14335 ( .A1(n13373), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12861) );
  XNOR2_X1 U14336 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n15103) );
  AOI21_X1 U14337 ( .B1(n13272), .B2(n15103), .A(n13303), .ZN(n12821) );
  NAND2_X1 U14338 ( .A1(n13296), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n12820) );
  OAI211_X1 U14339 ( .C1(n12861), .C2(n14731), .A(n12821), .B(n12820), .ZN(
        n12822) );
  INV_X1 U14340 ( .A(n12822), .ZN(n12823) );
  NAND2_X1 U14341 ( .A1(n13303), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12845) );
  NAND2_X1 U14342 ( .A1(n12824), .A2(n12845), .ZN(n14834) );
  XNOR2_X1 U14343 ( .A(n12826), .B(n12825), .ZN(n14819) );
  INV_X1 U14344 ( .A(n12827), .ZN(n12828) );
  XNOR2_X1 U14345 ( .A(n12829), .B(n12828), .ZN(n21581) );
  NAND2_X1 U14346 ( .A1(n21581), .A2(n14820), .ZN(n12834) );
  AOI22_X1 U14347 ( .A1(n12830), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n21917), .ZN(n12832) );
  INV_X1 U14348 ( .A(n12861), .ZN(n12839) );
  NAND2_X1 U14349 ( .A1(n12839), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12831) );
  AND2_X1 U14350 ( .A1(n12832), .A2(n12831), .ZN(n12833) );
  NAND2_X1 U14351 ( .A1(n12834), .A2(n12833), .ZN(n14693) );
  XNOR2_X1 U14352 ( .A(n12836), .B(n12835), .ZN(n21836) );
  AOI21_X1 U14353 ( .B1(n21836), .B2(n12639), .A(n21917), .ZN(n14692) );
  NAND2_X1 U14354 ( .A1(n14693), .A2(n14692), .ZN(n14691) );
  OR2_X1 U14355 ( .A1(n14693), .A2(n13302), .ZN(n12837) );
  NAND2_X1 U14356 ( .A1(n14691), .A2(n12837), .ZN(n14823) );
  AND2_X1 U14357 ( .A1(n14820), .A2(n14823), .ZN(n12838) );
  NAND2_X1 U14358 ( .A1(n14819), .A2(n12838), .ZN(n12844) );
  INV_X1 U14359 ( .A(n14823), .ZN(n12842) );
  AOI22_X1 U14360 ( .A1(n13296), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n21917), .ZN(n12841) );
  NAND2_X1 U14361 ( .A1(n12839), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12840) );
  AND2_X1 U14362 ( .A1(n12841), .A2(n12840), .ZN(n14821) );
  OAI21_X2 U14363 ( .B1(n14834), .B2(n14835), .A(n12845), .ZN(n14977) );
  INV_X1 U14364 ( .A(n16154), .ZN(n15112) );
  NAND2_X1 U14365 ( .A1(n12846), .A2(n15112), .ZN(n12847) );
  NAND2_X1 U14366 ( .A1(n12857), .A2(n12847), .ZN(n21769) );
  INV_X1 U14367 ( .A(n12848), .ZN(n12863) );
  INV_X1 U14368 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12850) );
  NAND2_X1 U14369 ( .A1(n12850), .A2(n12849), .ZN(n12851) );
  NAND2_X1 U14370 ( .A1(n12863), .A2(n12851), .ZN(n15240) );
  AOI22_X1 U14371 ( .A1(n15240), .A2(n13522), .B1(n13303), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12853) );
  NAND2_X1 U14372 ( .A1(n13296), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n12852) );
  OAI211_X1 U14373 ( .C1(n12861), .C2(n14746), .A(n12853), .B(n12852), .ZN(
        n12854) );
  INV_X1 U14374 ( .A(n12854), .ZN(n12855) );
  NAND2_X1 U14375 ( .A1(n14977), .A2(n14976), .ZN(n14975) );
  XNOR2_X1 U14376 ( .A(n12857), .B(n12856), .ZN(n13694) );
  INV_X1 U14377 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12860) );
  NAND2_X1 U14378 ( .A1(n21917), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12859) );
  NAND2_X1 U14379 ( .A1(n13296), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12858) );
  OAI211_X1 U14380 ( .C1(n12861), .C2(n12860), .A(n12859), .B(n12858), .ZN(
        n12862) );
  NAND2_X1 U14381 ( .A1(n12862), .A2(n13302), .ZN(n12867) );
  INV_X1 U14382 ( .A(n12873), .ZN(n12865) );
  INV_X1 U14383 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n21428) );
  NAND2_X1 U14384 ( .A1(n12863), .A2(n21428), .ZN(n12864) );
  NAND2_X1 U14385 ( .A1(n12865), .A2(n12864), .ZN(n21437) );
  NAND2_X1 U14386 ( .A1(n21437), .A2(n13522), .ZN(n12866) );
  NAND2_X1 U14387 ( .A1(n12867), .A2(n12866), .ZN(n12868) );
  XNOR2_X1 U14388 ( .A(n12872), .B(n12871), .ZN(n13702) );
  INV_X1 U14389 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n12875) );
  OAI21_X1 U14390 ( .B1(n12873), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n12879), .ZN(n21452) );
  AOI22_X1 U14391 ( .A1(n21452), .A2(n13522), .B1(n13303), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12874) );
  OAI21_X1 U14392 ( .B1(n13232), .B2(n12875), .A(n12874), .ZN(n12876) );
  AOI21_X1 U14393 ( .B1(n13702), .B2(n14820), .A(n12876), .ZN(n15078) );
  NAND2_X1 U14394 ( .A1(n12878), .A2(n12877), .ZN(n13714) );
  NAND2_X1 U14395 ( .A1(n13714), .A2(n14820), .ZN(n12887) );
  INV_X1 U14396 ( .A(n13303), .ZN(n12884) );
  NAND2_X1 U14397 ( .A1(n12879), .A2(n21455), .ZN(n12882) );
  INV_X1 U14398 ( .A(n12880), .ZN(n12881) );
  NAND2_X1 U14399 ( .A1(n12882), .A2(n12881), .ZN(n21463) );
  NAND2_X1 U14400 ( .A1(n21463), .A2(n13522), .ZN(n12883) );
  OAI21_X1 U14401 ( .B1(n21455), .B2(n12884), .A(n12883), .ZN(n12885) );
  AOI21_X1 U14402 ( .B1(n13296), .B2(P1_EAX_REG_6__SCAN_IN), .A(n12885), .ZN(
        n12886) );
  NAND2_X1 U14403 ( .A1(n12887), .A2(n12886), .ZN(n15087) );
  NAND2_X1 U14404 ( .A1(n15080), .A2(n15087), .ZN(n15086) );
  AOI22_X1 U14405 ( .A1(n12689), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12891) );
  AOI22_X1 U14406 ( .A1(n12688), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12695), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12890) );
  AOI22_X1 U14407 ( .A1(n12671), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12670), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12889) );
  AOI22_X1 U14408 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12728), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12888) );
  NAND4_X1 U14409 ( .A1(n12891), .A2(n12890), .A3(n12889), .A4(n12888), .ZN(
        n12897) );
  AOI22_X1 U14410 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12678), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12895) );
  AOI22_X1 U14411 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12894) );
  AOI22_X1 U14412 ( .A1(n10984), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12893) );
  AOI22_X1 U14413 ( .A1(n12672), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12774), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12892) );
  NAND4_X1 U14414 ( .A1(n12895), .A2(n12894), .A3(n12893), .A4(n12892), .ZN(
        n12896) );
  OAI21_X1 U14415 ( .B1(n12897), .B2(n12896), .A(n14820), .ZN(n12901) );
  INV_X1 U14416 ( .A(n12903), .ZN(n12898) );
  XNOR2_X1 U14417 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n12898), .ZN(
        n21480) );
  AOI22_X1 U14418 ( .A1(n13522), .A2(n21480), .B1(n13303), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12900) );
  NAND2_X1 U14419 ( .A1(n13296), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12899) );
  XOR2_X1 U14420 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n12917), .Z(n15460) );
  AOI22_X1 U14421 ( .A1(n12689), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12688), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12907) );
  AOI22_X1 U14422 ( .A1(n12727), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12678), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12906) );
  AOI22_X1 U14423 ( .A1(n12670), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12728), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12905) );
  AOI22_X1 U14424 ( .A1(n12671), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12904) );
  NAND4_X1 U14425 ( .A1(n12907), .A2(n12906), .A3(n12905), .A4(n12904), .ZN(
        n12913) );
  AOI22_X1 U14426 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n13279), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12911) );
  AOI22_X1 U14427 ( .A1(n12695), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12910) );
  AOI22_X1 U14428 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12909) );
  AOI22_X1 U14429 ( .A1(n12672), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12908) );
  NAND4_X1 U14430 ( .A1(n12911), .A2(n12910), .A3(n12909), .A4(n12908), .ZN(
        n12912) );
  OR2_X1 U14431 ( .A1(n12913), .A2(n12912), .ZN(n12914) );
  AOI22_X1 U14432 ( .A1(n14820), .A2(n12914), .B1(n13303), .B2(
        P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n12916) );
  NAND2_X1 U14433 ( .A1(n13296), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12915) );
  OAI211_X1 U14434 ( .C1(n15460), .C2(n13302), .A(n12916), .B(n12915), .ZN(
        n15441) );
  XNOR2_X1 U14435 ( .A(n12933), .B(n21502), .ZN(n19971) );
  NAND2_X1 U14436 ( .A1(n19971), .A2(n13522), .ZN(n12932) );
  AOI22_X1 U14437 ( .A1(n12689), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12688), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12921) );
  AOI22_X1 U14438 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10984), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12920) );
  AOI22_X1 U14439 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12678), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12919) );
  AOI22_X1 U14440 ( .A1(n12728), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12918) );
  NAND4_X1 U14441 ( .A1(n12921), .A2(n12920), .A3(n12919), .A4(n12918), .ZN(
        n12927) );
  AOI22_X1 U14442 ( .A1(n12695), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12925) );
  AOI22_X1 U14443 ( .A1(n12671), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12670), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12924) );
  AOI22_X1 U14444 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12923) );
  AOI22_X1 U14445 ( .A1(n12672), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12774), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12922) );
  NAND4_X1 U14446 ( .A1(n12925), .A2(n12924), .A3(n12923), .A4(n12922), .ZN(
        n12926) );
  OAI21_X1 U14447 ( .B1(n12927), .B2(n12926), .A(n14820), .ZN(n12930) );
  NAND2_X1 U14448 ( .A1(n13296), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n12929) );
  NAND2_X1 U14449 ( .A1(n13303), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12928) );
  AND3_X1 U14450 ( .A1(n12930), .A2(n12929), .A3(n12928), .ZN(n12931) );
  NAND2_X1 U14451 ( .A1(n12932), .A2(n12931), .ZN(n15434) );
  NAND2_X1 U14452 ( .A1(n13296), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n12936) );
  OAI21_X1 U14453 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12934), .A(
        n12972), .ZN(n21515) );
  AOI22_X1 U14454 ( .A1(n13522), .A2(n21515), .B1(n13303), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12935) );
  AND2_X1 U14455 ( .A1(n12936), .A2(n12935), .ZN(n15520) );
  AOI22_X1 U14456 ( .A1(n12760), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12940) );
  AOI22_X1 U14457 ( .A1(n12695), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n12679), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12939) );
  AOI22_X1 U14458 ( .A1(n10984), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12735), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12938) );
  AOI22_X1 U14459 ( .A1(n12761), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12937) );
  NAND4_X1 U14460 ( .A1(n12940), .A2(n12939), .A3(n12938), .A4(n12937), .ZN(
        n12946) );
  AOI22_X1 U14461 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12678), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12944) );
  AOI22_X1 U14462 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12696), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12943) );
  AOI22_X1 U14463 ( .A1(n12734), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12942) );
  AOI22_X1 U14464 ( .A1(n12736), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12941) );
  NAND4_X1 U14465 ( .A1(n12944), .A2(n12943), .A3(n12942), .A4(n12941), .ZN(
        n12945) );
  OR2_X1 U14466 ( .A1(n12946), .A2(n12945), .ZN(n12947) );
  NAND2_X1 U14467 ( .A1(n14820), .A2(n12947), .ZN(n15530) );
  OR2_X2 U14468 ( .A1(n15433), .A2(n15530), .ZN(n12980) );
  AOI22_X1 U14469 ( .A1(n10984), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12696), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12951) );
  AOI22_X1 U14470 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12688), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12950) );
  AOI22_X1 U14471 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12672), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12949) );
  AOI22_X1 U14472 ( .A1(n12736), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12948) );
  NAND4_X1 U14473 ( .A1(n12951), .A2(n12950), .A3(n12949), .A4(n12948), .ZN(
        n12957) );
  AOI22_X1 U14474 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12760), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12955) );
  AOI22_X1 U14475 ( .A1(n12695), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12737), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12954) );
  AOI22_X1 U14476 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12735), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12953) );
  AOI22_X1 U14477 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12952) );
  NAND4_X1 U14478 ( .A1(n12955), .A2(n12954), .A3(n12953), .A4(n12952), .ZN(
        n12956) );
  OAI21_X1 U14479 ( .B1(n12957), .B2(n12956), .A(n14820), .ZN(n12961) );
  NAND2_X1 U14480 ( .A1(n13296), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n12960) );
  XNOR2_X1 U14481 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12972), .ZN(
        n21525) );
  INV_X1 U14482 ( .A(n21525), .ZN(n12958) );
  AOI22_X1 U14483 ( .A1(n12958), .A2(n13522), .B1(n13303), .B2(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12959) );
  NAND3_X1 U14484 ( .A1(n12961), .A2(n12960), .A3(n12959), .ZN(n15532) );
  AOI22_X1 U14485 ( .A1(n12760), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12737), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12965) );
  AOI22_X1 U14486 ( .A1(n12671), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12735), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12964) );
  AOI22_X1 U14487 ( .A1(n10984), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12729), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12963) );
  AOI22_X1 U14488 ( .A1(n12672), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12962) );
  NAND4_X1 U14489 ( .A1(n12965), .A2(n12964), .A3(n12963), .A4(n12962), .ZN(
        n12971) );
  AOI22_X1 U14490 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13279), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12969) );
  AOI22_X1 U14491 ( .A1(n12695), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12968) );
  AOI22_X1 U14492 ( .A1(n12688), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12967) );
  AOI22_X1 U14493 ( .A1(n12728), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12966) );
  NAND4_X1 U14494 ( .A1(n12969), .A2(n12968), .A3(n12967), .A4(n12966), .ZN(
        n12970) );
  NOR2_X1 U14495 ( .A1(n12971), .A2(n12970), .ZN(n12977) );
  INV_X1 U14496 ( .A(n12981), .ZN(n12974) );
  XNOR2_X1 U14497 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n12974), .ZN(
        n16017) );
  AOI22_X1 U14498 ( .A1(n13522), .A2(n16017), .B1(n13303), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12976) );
  NAND2_X1 U14499 ( .A1(n13296), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12975) );
  OAI211_X1 U14500 ( .C1(n12978), .C2(n12977), .A(n12976), .B(n12975), .ZN(
        n15786) );
  NAND2_X1 U14501 ( .A1(n15532), .A2(n15786), .ZN(n12979) );
  AOI21_X4 U14502 ( .B1(n15529), .B2(n12980), .A(n12979), .ZN(n15787) );
  INV_X1 U14503 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15794) );
  XOR2_X1 U14504 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n12995), .Z(
        n19999) );
  AOI22_X1 U14505 ( .A1(n12688), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12695), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12985) );
  AOI22_X1 U14506 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n13279), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12984) );
  AOI22_X1 U14507 ( .A1(n12727), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12671), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12983) );
  AOI22_X1 U14508 ( .A1(n12689), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12982) );
  NAND4_X1 U14509 ( .A1(n12985), .A2(n12984), .A3(n12983), .A4(n12982), .ZN(
        n12991) );
  AOI22_X1 U14510 ( .A1(n12678), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12728), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12989) );
  AOI22_X1 U14511 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12988) );
  AOI22_X1 U14512 ( .A1(n12670), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12987) );
  AOI22_X1 U14513 ( .A1(n12672), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12986) );
  NAND4_X1 U14514 ( .A1(n12989), .A2(n12988), .A3(n12987), .A4(n12986), .ZN(
        n12990) );
  OR2_X1 U14515 ( .A1(n12991), .A2(n12990), .ZN(n12992) );
  AOI22_X1 U14516 ( .A1(n14820), .A2(n12992), .B1(n13303), .B2(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12994) );
  NAND2_X1 U14517 ( .A1(n13296), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12993) );
  OAI211_X1 U14518 ( .C1(n19999), .C2(n13302), .A(n12994), .B(n12993), .ZN(
        n15540) );
  INV_X1 U14519 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16004) );
  XNOR2_X1 U14520 ( .A(n13025), .B(n16004), .ZN(n16003) );
  NAND2_X1 U14521 ( .A1(n16003), .A2(n13522), .ZN(n13010) );
  AOI22_X1 U14522 ( .A1(n12689), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12695), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12999) );
  AOI22_X1 U14523 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12670), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12998) );
  AOI22_X1 U14524 ( .A1(n12734), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12997) );
  AOI22_X1 U14525 ( .A1(n12671), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12996) );
  NAND4_X1 U14526 ( .A1(n12999), .A2(n12998), .A3(n12997), .A4(n12996), .ZN(
        n13005) );
  AOI22_X1 U14527 ( .A1(n13278), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12679), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13003) );
  AOI22_X1 U14528 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12678), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13002) );
  AOI22_X1 U14529 ( .A1(n10984), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12696), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13001) );
  AOI22_X1 U14530 ( .A1(n12761), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12774), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13000) );
  NAND4_X1 U14531 ( .A1(n13003), .A2(n13002), .A3(n13001), .A4(n13000), .ZN(
        n13004) );
  OAI21_X1 U14532 ( .B1(n13005), .B2(n13004), .A(n14820), .ZN(n13008) );
  NAND2_X1 U14533 ( .A1(n13296), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n13007) );
  NAND2_X1 U14534 ( .A1(n13303), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13006) );
  AND3_X1 U14535 ( .A1(n13008), .A2(n13007), .A3(n13006), .ZN(n13009) );
  NAND2_X1 U14536 ( .A1(n13010), .A2(n13009), .ZN(n15768) );
  INV_X1 U14537 ( .A(n15577), .ZN(n16159) );
  AOI22_X1 U14538 ( .A1(n12760), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13014) );
  AOI22_X1 U14539 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13279), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13013) );
  AOI22_X1 U14540 ( .A1(n12727), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12735), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13012) );
  AOI22_X1 U14541 ( .A1(n12688), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12761), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13011) );
  NAND4_X1 U14542 ( .A1(n13014), .A2(n13013), .A3(n13012), .A4(n13011), .ZN(
        n13020) );
  AOI22_X1 U14543 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12696), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13018) );
  AOI22_X1 U14544 ( .A1(n12759), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13017) );
  AOI22_X1 U14545 ( .A1(n12671), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13016) );
  AOI22_X1 U14546 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13015) );
  NAND4_X1 U14547 ( .A1(n13018), .A2(n13017), .A3(n13016), .A4(n13015), .ZN(
        n13019) );
  NOR2_X1 U14548 ( .A1(n13020), .A2(n13019), .ZN(n13024) );
  NAND2_X1 U14549 ( .A1(n21917), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13021) );
  NAND2_X1 U14550 ( .A1(n13302), .A2(n13021), .ZN(n13022) );
  AOI21_X1 U14551 ( .B1(n13296), .B2(P1_EAX_REG_18__SCAN_IN), .A(n13022), .ZN(
        n13023) );
  OAI21_X1 U14552 ( .B1(n13299), .B2(n13024), .A(n13023), .ZN(n13029) );
  INV_X1 U14553 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n21545) );
  OAI21_X1 U14554 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n13026), .A(
        n13093), .ZN(n21564) );
  INV_X1 U14555 ( .A(n21564), .ZN(n13027) );
  NAND2_X1 U14556 ( .A1(n13027), .A2(n13522), .ZN(n13028) );
  NAND2_X1 U14557 ( .A1(n13029), .A2(n13028), .ZN(n15818) );
  AOI22_X1 U14558 ( .A1(n12688), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12695), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13033) );
  AOI22_X1 U14559 ( .A1(n10984), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12671), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13032) );
  AOI22_X1 U14560 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12678), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13031) );
  AOI22_X1 U14561 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13030) );
  NAND4_X1 U14562 ( .A1(n13033), .A2(n13032), .A3(n13031), .A4(n13030), .ZN(
        n13039) );
  AOI22_X1 U14563 ( .A1(n12689), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13037) );
  AOI22_X1 U14564 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12696), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13036) );
  AOI22_X1 U14565 ( .A1(n12673), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12761), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13035) );
  AOI22_X1 U14566 ( .A1(n12670), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13034) );
  NAND4_X1 U14567 ( .A1(n13037), .A2(n13036), .A3(n13035), .A4(n13034), .ZN(
        n13038) );
  OR2_X1 U14568 ( .A1(n13039), .A2(n13038), .ZN(n13044) );
  INV_X1 U14569 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13042) );
  INV_X1 U14570 ( .A(n13059), .ZN(n13040) );
  XNOR2_X1 U14571 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n13040), .ZN(
        n21546) );
  AOI22_X1 U14572 ( .A1(n13522), .A2(n21546), .B1(n13303), .B2(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n13041) );
  OAI21_X1 U14573 ( .B1(n13232), .B2(n13042), .A(n13041), .ZN(n13043) );
  AOI21_X1 U14574 ( .B1(n13269), .B2(n13044), .A(n13043), .ZN(n15819) );
  AOI22_X1 U14575 ( .A1(n12689), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12688), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13048) );
  AOI22_X1 U14576 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13279), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13047) );
  AOI22_X1 U14577 ( .A1(n12671), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12728), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13046) );
  AOI22_X1 U14578 ( .A1(n12673), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12761), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13045) );
  NAND4_X1 U14579 ( .A1(n13048), .A2(n13047), .A3(n13046), .A4(n13045), .ZN(
        n13054) );
  AOI22_X1 U14580 ( .A1(n12695), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13052) );
  AOI22_X1 U14581 ( .A1(n12727), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12678), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13051) );
  AOI22_X1 U14582 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13050) );
  AOI22_X1 U14583 ( .A1(n12670), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13049) );
  NAND4_X1 U14584 ( .A1(n13052), .A2(n13051), .A3(n13050), .A4(n13049), .ZN(
        n13053) );
  NOR2_X1 U14585 ( .A1(n13054), .A2(n13053), .ZN(n13058) );
  NAND2_X1 U14586 ( .A1(n21917), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n13055) );
  NAND2_X1 U14587 ( .A1(n13302), .A2(n13055), .ZN(n13056) );
  AOI21_X1 U14588 ( .B1(n13296), .B2(P1_EAX_REG_16__SCAN_IN), .A(n13056), .ZN(
        n13057) );
  OAI21_X1 U14589 ( .B1(n13299), .B2(n13058), .A(n13057), .ZN(n13062) );
  OAI21_X1 U14590 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n13060), .A(
        n13059), .ZN(n20014) );
  INV_X1 U14591 ( .A(n20014), .ZN(n21534) );
  NAND2_X1 U14592 ( .A1(n21534), .A2(n13522), .ZN(n13061) );
  NAND2_X1 U14593 ( .A1(n13062), .A2(n13061), .ZN(n15835) );
  AOI22_X1 U14594 ( .A1(n12734), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12759), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13067) );
  AOI22_X1 U14595 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13279), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13066) );
  AOI22_X1 U14596 ( .A1(n12671), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12735), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13065) );
  AOI22_X1 U14597 ( .A1(n12678), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12761), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13064) );
  NAND4_X1 U14598 ( .A1(n13067), .A2(n13066), .A3(n13065), .A4(n13064), .ZN(
        n13073) );
  AOI22_X1 U14599 ( .A1(n12689), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13071) );
  AOI22_X1 U14600 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13070) );
  AOI22_X1 U14601 ( .A1(n12728), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13069) );
  AOI22_X1 U14602 ( .A1(n12727), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13068) );
  NAND4_X1 U14603 ( .A1(n13071), .A2(n13070), .A3(n13069), .A4(n13068), .ZN(
        n13072) );
  NOR2_X1 U14604 ( .A1(n13073), .A2(n13072), .ZN(n13076) );
  INV_X1 U14605 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15982) );
  OAI21_X1 U14606 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15982), .A(n13302), 
        .ZN(n13074) );
  AOI21_X1 U14607 ( .B1(n13296), .B2(P1_EAX_REG_19__SCAN_IN), .A(n13074), .ZN(
        n13075) );
  OAI21_X1 U14608 ( .B1(n13299), .B2(n13076), .A(n13075), .ZN(n13078) );
  XNOR2_X1 U14609 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n13093), .ZN(
        n15986) );
  NAND2_X1 U14610 ( .A1(n13522), .A2(n15986), .ZN(n13077) );
  AOI22_X1 U14611 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12759), .B1(
        n12688), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13082) );
  AOI22_X1 U14612 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n12689), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13081) );
  AOI22_X1 U14613 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13080) );
  AOI22_X1 U14614 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13079) );
  NAND4_X1 U14615 ( .A1(n13082), .A2(n13081), .A3(n13080), .A4(n13079), .ZN(
        n13088) );
  AOI22_X1 U14616 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12736), .B1(
        n12735), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13086) );
  AOI22_X1 U14617 ( .A1(n12727), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12728), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13085) );
  AOI22_X1 U14618 ( .A1(n12737), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13084) );
  AOI22_X1 U14619 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12672), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13083) );
  NAND4_X1 U14620 ( .A1(n13086), .A2(n13085), .A3(n13084), .A4(n13083), .ZN(
        n13087) );
  NOR2_X1 U14621 ( .A1(n13088), .A2(n13087), .ZN(n13092) );
  NAND2_X1 U14622 ( .A1(n21917), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13089) );
  NAND2_X1 U14623 ( .A1(n13302), .A2(n13089), .ZN(n13090) );
  AOI21_X1 U14624 ( .B1(n13296), .B2(P1_EAX_REG_20__SCAN_IN), .A(n13090), .ZN(
        n13091) );
  OAI21_X1 U14625 ( .B1(n13299), .B2(n13092), .A(n13091), .ZN(n13097) );
  OAI21_X1 U14626 ( .B1(n13095), .B2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n13127), .ZN(n15973) );
  OR2_X1 U14627 ( .A1(n15973), .A2(n13302), .ZN(n13096) );
  AND2_X2 U14628 ( .A1(n15740), .A2(n15743), .ZN(n15724) );
  AOI22_X1 U14629 ( .A1(n12760), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12734), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13101) );
  AOI22_X1 U14630 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12727), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13100) );
  AOI22_X1 U14631 ( .A1(n12673), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12672), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13099) );
  AOI22_X1 U14632 ( .A1(n12735), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13098) );
  NAND4_X1 U14633 ( .A1(n13101), .A2(n13100), .A3(n13099), .A4(n13098), .ZN(
        n13107) );
  AOI22_X1 U14634 ( .A1(n12759), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13105) );
  AOI22_X1 U14635 ( .A1(n13279), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12678), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13104) );
  AOI22_X1 U14636 ( .A1(n12736), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12728), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13103) );
  AOI22_X1 U14637 ( .A1(n12737), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12774), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13102) );
  NAND4_X1 U14638 ( .A1(n13105), .A2(n13104), .A3(n13103), .A4(n13102), .ZN(
        n13106) );
  NOR2_X1 U14639 ( .A1(n13107), .A2(n13106), .ZN(n13110) );
  INV_X1 U14640 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15966) );
  OAI21_X1 U14641 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15966), .A(n13302), 
        .ZN(n13108) );
  AOI21_X1 U14642 ( .B1(n13296), .B2(P1_EAX_REG_21__SCAN_IN), .A(n13108), .ZN(
        n13109) );
  OAI21_X1 U14643 ( .B1(n13299), .B2(n13110), .A(n13109), .ZN(n13112) );
  XNOR2_X1 U14644 ( .A(n13127), .B(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15970) );
  NAND2_X1 U14645 ( .A1(n15970), .A2(n13522), .ZN(n13111) );
  AOI22_X1 U14646 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10984), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13116) );
  AOI22_X1 U14647 ( .A1(n12759), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13115) );
  AOI22_X1 U14648 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13114) );
  AOI22_X1 U14649 ( .A1(n12670), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13113) );
  NAND4_X1 U14650 ( .A1(n13116), .A2(n13115), .A3(n13114), .A4(n13113), .ZN(
        n13122) );
  AOI22_X1 U14651 ( .A1(n12689), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12688), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13120) );
  AOI22_X1 U14652 ( .A1(n12736), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12728), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13119) );
  AOI22_X1 U14653 ( .A1(n12737), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12774), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13118) );
  AOI22_X1 U14654 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12761), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13117) );
  NAND4_X1 U14655 ( .A1(n13120), .A2(n13119), .A3(n13118), .A4(n13117), .ZN(
        n13121) );
  NOR2_X1 U14656 ( .A1(n13122), .A2(n13121), .ZN(n13126) );
  INV_X1 U14657 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n21936) );
  OAI21_X1 U14658 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n21936), .A(
        n21917), .ZN(n13123) );
  INV_X1 U14659 ( .A(n13123), .ZN(n13124) );
  AOI21_X1 U14660 ( .B1(n13296), .B2(P1_EAX_REG_22__SCAN_IN), .A(n13124), .ZN(
        n13125) );
  OAI21_X1 U14661 ( .B1(n13299), .B2(n13126), .A(n13125), .ZN(n13133) );
  INV_X1 U14662 ( .A(n13128), .ZN(n13130) );
  INV_X1 U14663 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n13129) );
  NAND2_X1 U14664 ( .A1(n13130), .A2(n13129), .ZN(n13131) );
  NAND2_X1 U14665 ( .A1(n13158), .A2(n13131), .ZN(n15959) );
  NAND2_X1 U14666 ( .A1(n13133), .A2(n13132), .ZN(n15710) );
  AOI22_X1 U14667 ( .A1(n12695), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13137) );
  AOI22_X1 U14668 ( .A1(n12671), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12728), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13136) );
  AOI22_X1 U14669 ( .A1(n12688), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13135) );
  AOI22_X1 U14670 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12774), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13134) );
  NAND4_X1 U14671 ( .A1(n13137), .A2(n13136), .A3(n13135), .A4(n13134), .ZN(
        n13143) );
  AOI22_X1 U14672 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10984), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13141) );
  AOI22_X1 U14673 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12678), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13140) );
  AOI22_X1 U14674 ( .A1(n12689), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12672), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13139) );
  AOI22_X1 U14675 ( .A1(n12670), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13138) );
  NAND4_X1 U14676 ( .A1(n13141), .A2(n13140), .A3(n13139), .A4(n13138), .ZN(
        n13142) );
  NOR2_X1 U14677 ( .A1(n13143), .A2(n13142), .ZN(n13164) );
  AOI22_X1 U14678 ( .A1(n12670), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12728), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n13147) );
  AOI22_X1 U14679 ( .A1(n13278), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13146) );
  AOI22_X1 U14680 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12672), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13145) );
  AOI22_X1 U14681 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n13144) );
  NAND4_X1 U14682 ( .A1(n13147), .A2(n13146), .A3(n13145), .A4(n13144), .ZN(
        n13153) );
  AOI22_X1 U14683 ( .A1(n12689), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12695), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13151) );
  AOI22_X1 U14684 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12727), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13150) );
  AOI22_X1 U14685 ( .A1(n12688), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12678), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13149) );
  AOI22_X1 U14686 ( .A1(n12671), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13148) );
  NAND4_X1 U14687 ( .A1(n13151), .A2(n13150), .A3(n13149), .A4(n13148), .ZN(
        n13152) );
  NOR2_X1 U14688 ( .A1(n13153), .A2(n13152), .ZN(n13165) );
  XOR2_X1 U14689 ( .A(n13164), .B(n13165), .Z(n13154) );
  NAND2_X1 U14690 ( .A1(n13269), .A2(n13154), .ZN(n13157) );
  INV_X1 U14691 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15949) );
  NOR2_X1 U14692 ( .A1(n15949), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13155) );
  AOI211_X1 U14693 ( .C1(n13296), .C2(P1_EAX_REG_23__SCAN_IN), .A(n13522), .B(
        n13155), .ZN(n13156) );
  XNOR2_X1 U14694 ( .A(n13158), .B(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15953) );
  AOI22_X1 U14695 ( .A1(n13157), .A2(n13156), .B1(n13522), .B2(n15953), .ZN(
        n15697) );
  INV_X1 U14696 ( .A(n13158), .ZN(n13159) );
  INV_X1 U14697 ( .A(n13160), .ZN(n13162) );
  INV_X1 U14698 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n13161) );
  NAND2_X1 U14699 ( .A1(n13162), .A2(n13161), .ZN(n13163) );
  NAND2_X1 U14700 ( .A1(n13196), .A2(n13163), .ZN(n15943) );
  NOR2_X1 U14701 ( .A1(n13165), .A2(n13164), .ZN(n13191) );
  AOI22_X1 U14702 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12678), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13169) );
  AOI22_X1 U14703 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10984), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13168) );
  AOI22_X1 U14704 ( .A1(n12670), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12728), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13167) );
  AOI22_X1 U14705 ( .A1(n12736), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13166) );
  NAND4_X1 U14706 ( .A1(n13169), .A2(n13168), .A3(n13167), .A4(n13166), .ZN(
        n13175) );
  AOI22_X1 U14707 ( .A1(n12688), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12695), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13173) );
  AOI22_X1 U14708 ( .A1(n12689), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13172) );
  AOI22_X1 U14709 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13171) );
  AOI22_X1 U14710 ( .A1(n12672), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13170) );
  NAND4_X1 U14711 ( .A1(n13173), .A2(n13172), .A3(n13171), .A4(n13170), .ZN(
        n13174) );
  OR2_X1 U14712 ( .A1(n13175), .A2(n13174), .ZN(n13190) );
  XNOR2_X1 U14713 ( .A(n13191), .B(n13190), .ZN(n13178) );
  AOI21_X1 U14714 ( .B1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n21917), .A(
        n13522), .ZN(n13177) );
  NAND2_X1 U14715 ( .A1(n13296), .A2(P1_EAX_REG_24__SCAN_IN), .ZN(n13176) );
  OAI211_X1 U14716 ( .C1(n13178), .C2(n13299), .A(n13177), .B(n13176), .ZN(
        n13179) );
  OAI21_X1 U14717 ( .B1(n13302), .B2(n15943), .A(n13179), .ZN(n15691) );
  AOI22_X1 U14718 ( .A1(n12688), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13183) );
  AOI22_X1 U14719 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12678), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13182) );
  AOI22_X1 U14720 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13181) );
  AOI22_X1 U14721 ( .A1(n12736), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13180) );
  NAND4_X1 U14722 ( .A1(n13183), .A2(n13182), .A3(n13181), .A4(n13180), .ZN(
        n13189) );
  AOI22_X1 U14723 ( .A1(n12760), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12695), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13187) );
  AOI22_X1 U14724 ( .A1(n12727), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n13279), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13186) );
  AOI22_X1 U14725 ( .A1(n12670), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12696), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13185) );
  AOI22_X1 U14726 ( .A1(n12673), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12672), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13184) );
  NAND4_X1 U14727 ( .A1(n13187), .A2(n13186), .A3(n13185), .A4(n13184), .ZN(
        n13188) );
  NOR2_X1 U14728 ( .A1(n13189), .A2(n13188), .ZN(n13203) );
  NAND2_X1 U14729 ( .A1(n13191), .A2(n13190), .ZN(n13202) );
  XOR2_X1 U14730 ( .A(n13203), .B(n13202), .Z(n13192) );
  NAND2_X1 U14731 ( .A1(n13192), .A2(n13269), .ZN(n13195) );
  INV_X1 U14732 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15930) );
  NOR2_X1 U14733 ( .A1(n15930), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13193) );
  AOI211_X1 U14734 ( .C1(n13296), .C2(P1_EAX_REG_25__SCAN_IN), .A(n13522), .B(
        n13193), .ZN(n13194) );
  XNOR2_X1 U14735 ( .A(n13196), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15932) );
  AOI22_X1 U14736 ( .A1(n13195), .A2(n13194), .B1(n13272), .B2(n15932), .ZN(
        n15675) );
  INV_X1 U14737 ( .A(n13196), .ZN(n13197) );
  INV_X1 U14738 ( .A(n13198), .ZN(n13200) );
  INV_X1 U14739 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n13199) );
  NAND2_X1 U14740 ( .A1(n13200), .A2(n13199), .ZN(n13201) );
  NAND2_X1 U14741 ( .A1(n13236), .A2(n13201), .ZN(n15926) );
  NOR2_X1 U14742 ( .A1(n13203), .A2(n13202), .ZN(n13229) );
  AOI22_X1 U14743 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12678), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13207) );
  AOI22_X1 U14744 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10984), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13206) );
  AOI22_X1 U14745 ( .A1(n12670), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12728), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13205) );
  AOI22_X1 U14746 ( .A1(n12671), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13204) );
  NAND4_X1 U14747 ( .A1(n13207), .A2(n13206), .A3(n13205), .A4(n13204), .ZN(
        n13213) );
  AOI22_X1 U14748 ( .A1(n12734), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12695), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13211) );
  AOI22_X1 U14749 ( .A1(n12760), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13210) );
  AOI22_X1 U14750 ( .A1(n12679), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13209) );
  AOI22_X1 U14751 ( .A1(n12672), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13208) );
  NAND4_X1 U14752 ( .A1(n13211), .A2(n13210), .A3(n13209), .A4(n13208), .ZN(
        n13212) );
  OR2_X1 U14753 ( .A1(n13213), .A2(n13212), .ZN(n13228) );
  XNOR2_X1 U14754 ( .A(n13229), .B(n13228), .ZN(n13216) );
  AOI21_X1 U14755 ( .B1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n21917), .A(
        n13522), .ZN(n13215) );
  NAND2_X1 U14756 ( .A1(n13296), .A2(P1_EAX_REG_26__SCAN_IN), .ZN(n13214) );
  OAI211_X1 U14757 ( .C1(n13216), .C2(n13299), .A(n13215), .B(n13214), .ZN(
        n13217) );
  OAI21_X1 U14758 ( .B1(n13302), .B2(n15926), .A(n13217), .ZN(n15665) );
  XNOR2_X1 U14759 ( .A(n13236), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15922) );
  AOI22_X1 U14760 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12734), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13221) );
  AOI22_X1 U14761 ( .A1(n12729), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12696), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13220) );
  AOI22_X1 U14762 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12679), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13219) );
  AOI22_X1 U14763 ( .A1(n12672), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12774), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13218) );
  NAND4_X1 U14764 ( .A1(n13221), .A2(n13220), .A3(n13219), .A4(n13218), .ZN(
        n13227) );
  AOI22_X1 U14765 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12759), .B1(
        n12760), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13225) );
  AOI22_X1 U14766 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n13280), .B1(
        n13279), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13224) );
  AOI22_X1 U14767 ( .A1(n12727), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12670), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13223) );
  AOI22_X1 U14768 ( .A1(n12671), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13222) );
  NAND4_X1 U14769 ( .A1(n13225), .A2(n13224), .A3(n13223), .A4(n13222), .ZN(
        n13226) );
  NOR2_X1 U14770 ( .A1(n13227), .A2(n13226), .ZN(n13241) );
  NAND2_X1 U14771 ( .A1(n13229), .A2(n13228), .ZN(n13240) );
  XOR2_X1 U14772 ( .A(n13241), .B(n13240), .Z(n13234) );
  INV_X1 U14773 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n13231) );
  NAND2_X1 U14774 ( .A1(n21917), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13230) );
  OAI211_X1 U14775 ( .C1(n13232), .C2(n13231), .A(n13302), .B(n13230), .ZN(
        n13233) );
  AOI21_X1 U14776 ( .B1(n13234), .B2(n13269), .A(n13233), .ZN(n13235) );
  AOI21_X1 U14777 ( .B1(n13272), .B2(n15922), .A(n13235), .ZN(n15649) );
  INV_X1 U14778 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15918) );
  INV_X1 U14779 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13237) );
  NAND2_X1 U14780 ( .A1(n13238), .A2(n13237), .ZN(n13239) );
  NAND2_X1 U14781 ( .A1(n13275), .A2(n13239), .ZN(n15902) );
  NOR2_X1 U14782 ( .A1(n13241), .A2(n13240), .ZN(n13268) );
  AOI22_X1 U14783 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12729), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13245) );
  AOI22_X1 U14784 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12727), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13244) );
  AOI22_X1 U14785 ( .A1(n12670), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12728), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13243) );
  AOI22_X1 U14786 ( .A1(n12671), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13242) );
  NAND4_X1 U14787 ( .A1(n13245), .A2(n13244), .A3(n13243), .A4(n13242), .ZN(
        n13251) );
  AOI22_X1 U14788 ( .A1(n12734), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12695), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13249) );
  AOI22_X1 U14789 ( .A1(n12689), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13248) );
  AOI22_X1 U14790 ( .A1(n12737), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13247) );
  AOI22_X1 U14791 ( .A1(n12672), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13246) );
  NAND4_X1 U14792 ( .A1(n13249), .A2(n13248), .A3(n13247), .A4(n13246), .ZN(
        n13250) );
  OR2_X1 U14793 ( .A1(n13251), .A2(n13250), .ZN(n13267) );
  XNOR2_X1 U14794 ( .A(n13268), .B(n13267), .ZN(n13254) );
  AOI21_X1 U14795 ( .B1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n21917), .A(
        n13522), .ZN(n13253) );
  NAND2_X1 U14796 ( .A1(n13296), .A2(P1_EAX_REG_28__SCAN_IN), .ZN(n13252) );
  OAI211_X1 U14797 ( .C1(n13254), .C2(n13299), .A(n13253), .B(n13252), .ZN(
        n13255) );
  OAI21_X1 U14798 ( .B1(n13302), .B2(n15902), .A(n13255), .ZN(n15636) );
  AOI22_X1 U14799 ( .A1(n12689), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13278), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13259) );
  AOI22_X1 U14800 ( .A1(n12737), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13258) );
  AOI22_X1 U14801 ( .A1(n10984), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13257) );
  AOI22_X1 U14802 ( .A1(n12678), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10982), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13256) );
  NAND4_X1 U14803 ( .A1(n13259), .A2(n13258), .A3(n13257), .A4(n13256), .ZN(
        n13266) );
  AOI22_X1 U14804 ( .A1(n12734), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12759), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13264) );
  AOI22_X1 U14805 ( .A1(n12671), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12735), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13263) );
  AOI22_X1 U14806 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12696), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13262) );
  AOI22_X1 U14807 ( .A1(n13260), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12672), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13261) );
  NAND4_X1 U14808 ( .A1(n13264), .A2(n13263), .A3(n13262), .A4(n13261), .ZN(
        n13265) );
  NOR2_X1 U14809 ( .A1(n13266), .A2(n13265), .ZN(n13293) );
  NAND2_X1 U14810 ( .A1(n13268), .A2(n13267), .ZN(n13292) );
  XOR2_X1 U14811 ( .A(n13293), .B(n13292), .Z(n13270) );
  NAND2_X1 U14812 ( .A1(n13270), .A2(n13269), .ZN(n13274) );
  INV_X1 U14813 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15588) );
  AOI21_X1 U14814 ( .B1(n15588), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n13271) );
  AOI21_X1 U14815 ( .B1(n12830), .B2(P1_EAX_REG_29__SCAN_IN), .A(n13271), .ZN(
        n13273) );
  XNOR2_X1 U14816 ( .A(n13275), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n15591) );
  AOI22_X1 U14817 ( .A1(n13274), .A2(n13273), .B1(n13272), .B2(n15591), .ZN(
        n13780) );
  INV_X1 U14818 ( .A(n13275), .ZN(n13276) );
  NAND2_X1 U14819 ( .A1(n13276), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13529) );
  INV_X1 U14820 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13277) );
  XNOR2_X1 U14821 ( .A(n13529), .B(n13277), .ZN(n15898) );
  AOI22_X1 U14822 ( .A1(n13278), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12737), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13284) );
  AOI22_X1 U14823 ( .A1(n13280), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13279), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13283) );
  AOI22_X1 U14824 ( .A1(n12736), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12728), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13282) );
  AOI22_X1 U14825 ( .A1(n12761), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12774), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n13281) );
  NAND4_X1 U14826 ( .A1(n13284), .A2(n13283), .A3(n13282), .A4(n13281), .ZN(
        n13291) );
  AOI22_X1 U14827 ( .A1(n12689), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12759), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13289) );
  AOI22_X1 U14828 ( .A1(n12727), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12729), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13288) );
  AOI22_X1 U14829 ( .A1(n12688), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12673), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13287) );
  AOI22_X1 U14830 ( .A1(n12670), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n13285), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13286) );
  NAND4_X1 U14831 ( .A1(n13289), .A2(n13288), .A3(n13287), .A4(n13286), .ZN(
        n13290) );
  NOR2_X1 U14832 ( .A1(n13291), .A2(n13290), .ZN(n13295) );
  NOR2_X1 U14833 ( .A1(n13293), .A2(n13292), .ZN(n13294) );
  XOR2_X1 U14834 ( .A(n13295), .B(n13294), .Z(n13300) );
  AOI21_X1 U14835 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n21917), .A(
        n13522), .ZN(n13298) );
  NAND2_X1 U14836 ( .A1(n13296), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n13297) );
  OAI211_X1 U14837 ( .C1(n13300), .C2(n13299), .A(n13298), .B(n13297), .ZN(
        n13301) );
  OAI21_X1 U14838 ( .B1(n13302), .B2(n15898), .A(n13301), .ZN(n15623) );
  AOI22_X1 U14839 ( .A1(n12830), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n13303), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13304) );
  NAND2_X1 U14840 ( .A1(n21915), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13312) );
  INV_X1 U14841 ( .A(n13312), .ZN(n13305) );
  XNOR2_X1 U14842 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13313) );
  AOI22_X1 U14843 ( .A1(n13305), .A2(n13313), .B1(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n21794), .ZN(n13326) );
  XNOR2_X1 U14844 ( .A(n14731), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13327) );
  OAI22_X1 U14845 ( .A1(n13326), .A2(n13327), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n14731), .ZN(n13310) );
  OAI21_X1 U14846 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n21933), .A(
        n13310), .ZN(n13306) );
  OAI21_X1 U14847 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n14746), .A(
        n13306), .ZN(n13308) );
  INV_X1 U14848 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n16977) );
  NAND2_X1 U14849 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n12860), .ZN(
        n13307) );
  OAI221_X1 U14850 ( .B1(n13308), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), 
        .C1(n13308), .C2(n16977), .A(n13307), .ZN(n13355) );
  NAND2_X1 U14851 ( .A1(n15596), .A2(n12623), .ZN(n13732) );
  NOR3_X1 U14852 ( .A1(n13308), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        n16977), .ZN(n13332) );
  XNOR2_X1 U14853 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n13309) );
  XNOR2_X1 U14854 ( .A(n13310), .B(n13309), .ZN(n13330) );
  NOR2_X1 U14855 ( .A1(n13332), .A2(n13330), .ZN(n13350) );
  OAI21_X1 U14856 ( .B1(n21915), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n13312), .ZN(n13316) );
  INV_X1 U14857 ( .A(n13316), .ZN(n13311) );
  NAND2_X1 U14858 ( .A1(n13333), .A2(n13311), .ZN(n13319) );
  XNOR2_X1 U14859 ( .A(n13313), .B(n13312), .ZN(n13353) );
  NAND2_X1 U14860 ( .A1(n15156), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13320) );
  OAI21_X1 U14861 ( .B1(n13314), .B2(n13353), .A(n13320), .ZN(n13321) );
  NOR3_X1 U14862 ( .A1(n13321), .A2(n12623), .A3(n13353), .ZN(n13318) );
  INV_X1 U14863 ( .A(n14717), .ZN(n13653) );
  AND2_X1 U14864 ( .A1(n16174), .A2(n15596), .ZN(n13315) );
  AOI211_X1 U14865 ( .C1(n13653), .C2(n15124), .A(n13316), .B(n13334), .ZN(
        n13317) );
  AOI211_X1 U14866 ( .C1(n13344), .C2(n13319), .A(n13318), .B(n13317), .ZN(
        n13325) );
  INV_X1 U14867 ( .A(n13353), .ZN(n13323) );
  NAND3_X1 U14868 ( .A1(n13345), .A2(n13320), .A3(n12623), .ZN(n13329) );
  AOI21_X1 U14869 ( .B1(n13333), .B2(n12623), .A(n13321), .ZN(n13322) );
  AOI21_X1 U14870 ( .B1(n13323), .B2(n13329), .A(n13322), .ZN(n13324) );
  XOR2_X1 U14871 ( .A(n13327), .B(n13326), .Z(n13351) );
  INV_X1 U14872 ( .A(n13351), .ZN(n13328) );
  AOI21_X1 U14873 ( .B1(n13341), .B2(n13328), .A(n13334), .ZN(n13338) );
  INV_X1 U14874 ( .A(n13329), .ZN(n13331) );
  AOI22_X1 U14875 ( .A1(n13332), .A2(n13331), .B1(n13720), .B2(n13330), .ZN(
        n13337) );
  INV_X1 U14876 ( .A(n13339), .ZN(n13335) );
  OAI211_X1 U14877 ( .C1(n13335), .C2(n13334), .A(n13333), .B(n13351), .ZN(
        n13336) );
  OAI211_X1 U14878 ( .C1(n13339), .C2(n13338), .A(n13337), .B(n13336), .ZN(
        n13340) );
  INV_X1 U14879 ( .A(n12626), .ZN(n13348) );
  NOR2_X1 U14880 ( .A1(n13348), .A2(n15577), .ZN(n14729) );
  NAND2_X1 U14881 ( .A1(n14729), .A2(n15093), .ZN(n14858) );
  NAND2_X1 U14882 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n21622) );
  INV_X1 U14883 ( .A(n21622), .ZN(n21624) );
  AND2_X1 U14884 ( .A1(n13351), .A2(n13350), .ZN(n13352) );
  NAND2_X1 U14885 ( .A1(n13353), .A2(n13352), .ZN(n13354) );
  NAND2_X1 U14886 ( .A1(n13355), .A2(n13354), .ZN(n15608) );
  OR2_X1 U14887 ( .A1(n13349), .A2(n15608), .ZN(n13524) );
  OAI22_X1 U14888 ( .A1(n15613), .A2(n14858), .B1(n21624), .B2(n13524), .ZN(
        n14712) );
  OR2_X1 U14889 ( .A1(n14846), .A2(n10976), .ZN(n14862) );
  INV_X1 U14890 ( .A(n14862), .ZN(n13356) );
  NAND2_X1 U14891 ( .A1(n13356), .A2(n21622), .ZN(n14700) );
  INV_X1 U14892 ( .A(n15093), .ZN(n14724) );
  INV_X1 U14893 ( .A(n14948), .ZN(n15597) );
  NAND4_X1 U14894 ( .A1(n12627), .A2(n13357), .A3(n15597), .A4(n22148), .ZN(
        n14688) );
  OAI22_X1 U14895 ( .A1(n15613), .A2(n14700), .B1(n14724), .B2(n14688), .ZN(
        n13358) );
  AND2_X1 U14896 ( .A1(n15886), .A2(n15597), .ZN(n13360) );
  NOR4_X1 U14897 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13364) );
  NOR4_X1 U14898 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n13363) );
  NOR4_X1 U14899 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13362) );
  NOR4_X1 U14900 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n13361) );
  AND4_X1 U14901 ( .A1(n13364), .A2(n13363), .A3(n13362), .A4(n13361), .ZN(
        n13369) );
  NOR4_X1 U14902 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n13367) );
  NOR4_X1 U14903 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n13366) );
  NOR4_X1 U14904 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13365) );
  INV_X1 U14905 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n19879) );
  AND4_X1 U14906 ( .A1(n13367), .A2(n13366), .A3(n13365), .A4(n19879), .ZN(
        n13368) );
  NAND2_X1 U14907 ( .A1(n13369), .A2(n13368), .ZN(n13370) );
  NOR3_X1 U14908 ( .A1(n15887), .A2(n14844), .A3(n15599), .ZN(n13371) );
  AOI22_X1 U14909 ( .A1(n15878), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P1_EAX_REG_31__SCAN_IN), .B2(n15887), .ZN(n13372) );
  INV_X1 U14910 ( .A(n13372), .ZN(n13375) );
  NAND3_X1 U14911 ( .A1(n15886), .A2(n13373), .A3(n15599), .ZN(n15595) );
  INV_X1 U14912 ( .A(DATAI_31_), .ZN(n15167) );
  NOR2_X1 U14913 ( .A1(n15595), .A2(n15167), .ZN(n13374) );
  NOR2_X1 U14914 ( .A1(n13375), .A2(n13374), .ZN(n13376) );
  NAND2_X1 U14915 ( .A1(n13377), .A2(n13376), .ZN(P1_U2873) );
  INV_X1 U14916 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13378) );
  NAND2_X1 U14917 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n20313) );
  NAND2_X1 U14918 ( .A1(n17990), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17778) );
  INV_X1 U14919 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n20339) );
  INV_X1 U14920 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n20357) );
  NOR2_X1 U14921 ( .A1(n20339), .A2(n20357), .ZN(n20351) );
  INV_X1 U14922 ( .A(n20351), .ZN(n17788) );
  INV_X1 U14923 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n13379) );
  INV_X1 U14924 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17846) );
  INV_X1 U14925 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17860) );
  INV_X1 U14926 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n20485) );
  INV_X1 U14927 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n20495) );
  NAND2_X1 U14928 ( .A1(n17899), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n17962) );
  INV_X1 U14929 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n20523) );
  XNOR2_X1 U14930 ( .A(n13391), .B(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n20536) );
  INV_X1 U14931 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n20095) );
  INV_X1 U14932 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n21098) );
  INV_X1 U14933 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n21612) );
  NAND4_X1 U14934 ( .A1(n20095), .A2(n21098), .A3(n21612), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n21229) );
  INV_X1 U14935 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n17940) );
  INV_X1 U14936 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n20538) );
  AND2_X1 U14937 ( .A1(n17899), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13381) );
  INV_X1 U14938 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20150) );
  NOR2_X1 U14939 ( .A1(n17962), .A2(n20150), .ZN(n17938) );
  INV_X1 U14940 ( .A(n17938), .ZN(n13380) );
  OAI21_X1 U14941 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n13381), .A(
        n13380), .ZN(n20516) );
  NAND2_X1 U14942 ( .A1(n17895), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13382) );
  AOI21_X1 U14943 ( .B1(n20495), .B2(n13382), .A(n13381), .ZN(n17913) );
  INV_X1 U14944 ( .A(n17913), .ZN(n20501) );
  NOR2_X1 U14945 ( .A1(n11061), .A2(n20150), .ZN(n13383) );
  OAI21_X1 U14946 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n13383), .A(
        n13382), .ZN(n20490) );
  INV_X1 U14947 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n20454) );
  NAND2_X1 U14948 ( .A1(n17872), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13385) );
  NOR2_X1 U14949 ( .A1(n20454), .A2(n13385), .ZN(n13384) );
  INV_X1 U14950 ( .A(n13383), .ZN(n17897) );
  OAI21_X1 U14951 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n13384), .A(
        n17897), .ZN(n20477) );
  XNOR2_X1 U14952 ( .A(n20454), .B(n13385), .ZN(n20462) );
  NOR2_X1 U14953 ( .A1(n17857), .A2(n20150), .ZN(n13387) );
  OAI21_X1 U14954 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n13387), .A(
        n13385), .ZN(n20444) );
  INV_X1 U14955 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17821) );
  NAND2_X1 U14956 ( .A1(n13386), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13390) );
  NOR2_X1 U14957 ( .A1(n17821), .A2(n13390), .ZN(n13388) );
  INV_X1 U14958 ( .A(n13387), .ZN(n17859) );
  OAI21_X1 U14959 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n13388), .A(
        n17859), .ZN(n20435) );
  NOR2_X1 U14960 ( .A1(n17847), .A2(n20150), .ZN(n17823) );
  OAI21_X1 U14961 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17823), .A(
        n13390), .ZN(n20410) );
  NOR2_X1 U14962 ( .A1(n11054), .A2(n20150), .ZN(n17751) );
  INV_X1 U14963 ( .A(n17823), .ZN(n13389) );
  OAI21_X1 U14964 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17751), .A(
        n13389), .ZN(n20399) );
  INV_X1 U14965 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n20553) );
  NAND2_X1 U14966 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n20553), .ZN(
        n20312) );
  NAND2_X1 U14967 ( .A1(n20399), .A2(n20398), .ZN(n20397) );
  NAND2_X1 U14968 ( .A1(n10967), .A2(n20397), .ZN(n20409) );
  NAND2_X1 U14969 ( .A1(n20410), .A2(n20409), .ZN(n20408) );
  XOR2_X1 U14970 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n13390), .Z(
        n20417) );
  NAND2_X1 U14971 ( .A1(n10967), .A2(n20442), .ZN(n20461) );
  NAND2_X1 U14972 ( .A1(n20462), .A2(n20461), .ZN(n20460) );
  NAND2_X1 U14973 ( .A1(n10967), .A2(n20460), .ZN(n20476) );
  NAND2_X1 U14974 ( .A1(n20477), .A2(n20476), .ZN(n20475) );
  NAND2_X1 U14975 ( .A1(n10967), .A2(n20475), .ZN(n20489) );
  NAND2_X1 U14976 ( .A1(n20490), .A2(n20489), .ZN(n20488) );
  NAND2_X1 U14977 ( .A1(n20488), .A2(n10967), .ZN(n20500) );
  OAI21_X1 U14978 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n17938), .A(
        n13391), .ZN(n20531) );
  NAND2_X1 U14979 ( .A1(n20530), .A2(n20531), .ZN(n20535) );
  NOR4_X1 U14980 ( .A1(n20536), .A2(n21229), .A3(n20332), .A4(n20535), .ZN(
        n13521) );
  NAND2_X1 U14981 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n21659) );
  AOI22_X1 U14982 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17722), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13399) );
  NOR2_X2 U14983 ( .A1(n20146), .A2(n13393), .ZN(n13456) );
  AOI22_X1 U14984 ( .A1(n17688), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13456), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13398) );
  NOR3_X1 U14985 ( .A1(n20748), .A2(n20759), .A3(n20777), .ZN(n13394) );
  INV_X1 U14986 ( .A(n13394), .ZN(n13395) );
  AOI22_X1 U14987 ( .A1(n20181), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13397) );
  NOR2_X2 U14988 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n20155), .ZN(
        n17356) );
  AOI22_X1 U14989 ( .A1(n13934), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17713), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13396) );
  NAND4_X1 U14990 ( .A1(n13399), .A2(n13398), .A3(n13397), .A4(n13396), .ZN(
        n13409) );
  BUF_X2 U14991 ( .A(n13440), .Z(n17465) );
  AOI22_X1 U14992 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13407) );
  NOR2_X2 U14993 ( .A1(n13401), .A2(n13400), .ZN(n13897) );
  AOI22_X1 U14994 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n13406) );
  OR2_X2 U14995 ( .A1(n20146), .A2(n20777), .ZN(n17655) );
  AOI22_X1 U14996 ( .A1(n17585), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17703), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13405) );
  NOR2_X2 U14997 ( .A1(n13403), .A2(n20146), .ZN(n13981) );
  AOI22_X1 U14998 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n13981), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13404) );
  NAND4_X1 U14999 ( .A1(n13407), .A2(n13406), .A3(n13405), .A4(n13404), .ZN(
        n13408) );
  INV_X1 U15000 ( .A(n18919), .ZN(n13475) );
  AOI22_X1 U15001 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13413) );
  AOI22_X1 U15002 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13412) );
  AOI22_X1 U15003 ( .A1(n13934), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n13463), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13411) );
  AOI22_X1 U15004 ( .A1(n17683), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13410) );
  NAND4_X1 U15005 ( .A1(n13413), .A2(n13412), .A3(n13411), .A4(n13410), .ZN(
        n13419) );
  AOI22_X1 U15006 ( .A1(n17585), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n13981), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13417) );
  AOI22_X1 U15007 ( .A1(n17719), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17689), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13416) );
  AOI22_X1 U15008 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17502), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13415) );
  INV_X2 U15009 ( .A(n13479), .ZN(n17688) );
  AOI22_X1 U15010 ( .A1(n17688), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17535), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13414) );
  NAND4_X1 U15011 ( .A1(n13417), .A2(n13416), .A3(n13415), .A4(n13414), .ZN(
        n13418) );
  CLKBUF_X3 U15012 ( .A(n13468), .Z(n17561) );
  AOI22_X1 U15013 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13423) );
  AOI22_X1 U15014 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17535), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13422) );
  AOI22_X1 U15015 ( .A1(n13934), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n20181), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13421) );
  AOI22_X1 U15016 ( .A1(n17713), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13420) );
  NAND4_X1 U15017 ( .A1(n13423), .A2(n13422), .A3(n13421), .A4(n13420), .ZN(
        n13429) );
  AOI22_X1 U15018 ( .A1(n17688), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13427) );
  AOI22_X1 U15019 ( .A1(n17585), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17502), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n13426) );
  AOI22_X1 U15020 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17689), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13425) );
  AOI22_X1 U15021 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13424) );
  NAND4_X1 U15022 ( .A1(n13427), .A2(n13426), .A3(n13425), .A4(n13424), .ZN(
        n13428) );
  AOI22_X1 U15023 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13439) );
  AOI22_X1 U15024 ( .A1(n17722), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13438) );
  AOI22_X1 U15025 ( .A1(n17689), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13430) );
  OAI21_X1 U15026 ( .B1(n13479), .B2(n18793), .A(n13430), .ZN(n13436) );
  AOI22_X1 U15027 ( .A1(n17719), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17723), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13434) );
  AOI22_X1 U15028 ( .A1(n17703), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13433) );
  AOI22_X1 U15029 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17683), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13432) );
  AOI22_X1 U15030 ( .A1(n17713), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17714), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13431) );
  NAND4_X1 U15031 ( .A1(n13434), .A2(n13433), .A3(n13432), .A4(n13431), .ZN(
        n13435) );
  NAND3_X2 U15032 ( .A1(n13439), .A2(n13438), .A3(n13437), .ZN(n20661) );
  AOI22_X1 U15033 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n13456), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13451) );
  AOI22_X1 U15034 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13450) );
  INV_X1 U15035 ( .A(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13448) );
  AOI22_X1 U15036 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13441) );
  OAI21_X1 U15037 ( .B1(n13479), .B2(n18876), .A(n13441), .ZN(n13442) );
  INV_X1 U15038 ( .A(n13442), .ZN(n13447) );
  AOI22_X1 U15039 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17502), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13446) );
  AOI22_X1 U15040 ( .A1(n17722), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n13981), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13445) );
  AOI22_X1 U15041 ( .A1(n13934), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n13463), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13444) );
  AOI22_X1 U15042 ( .A1(n17683), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13443) );
  AOI22_X1 U15043 ( .A1(n17688), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17585), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13455) );
  AOI22_X1 U15044 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17502), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13454) );
  AOI22_X1 U15045 ( .A1(n17683), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n13463), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13453) );
  AOI22_X1 U15046 ( .A1(n13934), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13452) );
  NAND4_X1 U15047 ( .A1(n13455), .A2(n13454), .A3(n13453), .A4(n13452), .ZN(
        n13462) );
  AOI22_X1 U15048 ( .A1(n17689), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17535), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13460) );
  AOI22_X1 U15049 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17723), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13459) );
  AOI22_X1 U15050 ( .A1(n17719), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13458) );
  AOI22_X1 U15051 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13457) );
  NAND4_X1 U15052 ( .A1(n13460), .A2(n13459), .A3(n13458), .A4(n13457), .ZN(
        n13461) );
  NAND2_X1 U15053 ( .A1(n20624), .A2(n20625), .ZN(n13877) );
  NOR4_X2 U15054 ( .A1(n13475), .A2(n17346), .A3(n13494), .A4(n13877), .ZN(
        n20831) );
  AOI22_X1 U15055 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13981), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13467) );
  AOI22_X1 U15056 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13466) );
  AOI22_X1 U15057 ( .A1(n13934), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n13463), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13465) );
  AOI22_X1 U15058 ( .A1(n17683), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13464) );
  NAND4_X1 U15059 ( .A1(n13467), .A2(n13466), .A3(n13465), .A4(n13464), .ZN(
        n13474) );
  AOI22_X1 U15060 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17689), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13472) );
  AOI22_X1 U15061 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17535), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13471) );
  AOI22_X1 U15062 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13470) );
  AOI22_X1 U15063 ( .A1(n17719), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17502), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n13469) );
  NAND4_X1 U15064 ( .A1(n13472), .A2(n13471), .A3(n13470), .A4(n13469), .ZN(
        n13473) );
  NAND2_X1 U15065 ( .A1(n20831), .A2(n13476), .ZN(n13883) );
  INV_X1 U15066 ( .A(n13883), .ZN(n13477) );
  NAND2_X1 U15067 ( .A1(n17346), .A2(n18796), .ZN(n20763) );
  NAND2_X1 U15068 ( .A1(n18837), .A2(n20625), .ZN(n13882) );
  NOR2_X1 U15069 ( .A1(n13476), .A2(n17346), .ZN(n13880) );
  NOR3_X1 U15070 ( .A1(n20624), .A2(n13970), .A3(n13493), .ZN(n13489) );
  NOR2_X1 U15071 ( .A1(n13477), .A2(n13489), .ZN(n21193) );
  AOI22_X1 U15072 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13478) );
  OAI21_X1 U15073 ( .B1(n13479), .B2(n19049), .A(n13478), .ZN(n13485) );
  AOI22_X1 U15074 ( .A1(n17722), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13483) );
  AOI22_X1 U15075 ( .A1(n17703), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13482) );
  AOI22_X1 U15076 ( .A1(n17713), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13481) );
  AOI22_X1 U15077 ( .A1(n13934), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n20181), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13480) );
  NAND4_X1 U15078 ( .A1(n13483), .A2(n13482), .A3(n13481), .A4(n13480), .ZN(
        n13484) );
  NAND2_X1 U15079 ( .A1(n19057), .A2(n20559), .ZN(n13965) );
  NAND2_X1 U15080 ( .A1(n19007), .A2(n13489), .ZN(n21222) );
  NAND2_X1 U15081 ( .A1(n20559), .A2(n13489), .ZN(n13497) );
  NAND2_X1 U15082 ( .A1(n18961), .A2(n18919), .ZN(n20762) );
  NOR2_X1 U15083 ( .A1(n13494), .A2(n17345), .ZN(n13490) );
  NAND2_X1 U15084 ( .A1(n18961), .A2(n13965), .ZN(n13885) );
  AOI21_X1 U15085 ( .B1(n20661), .B2(n13877), .A(n18878), .ZN(n13492) );
  AOI21_X1 U15086 ( .B1(n13877), .B2(n13885), .A(n13492), .ZN(n13496) );
  NAND2_X1 U15087 ( .A1(n11096), .A2(n19007), .ZN(n13966) );
  NOR2_X1 U15088 ( .A1(n20722), .A2(n20746), .ZN(n20563) );
  NOR2_X1 U15089 ( .A1(n13966), .A2(n20563), .ZN(n13881) );
  AOI211_X1 U15090 ( .C1(n13494), .C2(n18919), .A(n13881), .B(n13493), .ZN(
        n13495) );
  NAND2_X1 U15091 ( .A1(n13496), .A2(n13495), .ZN(n20779) );
  INV_X1 U15092 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n20754) );
  NAND2_X1 U15093 ( .A1(n20754), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n21225) );
  NOR2_X1 U15094 ( .A1(n21098), .A2(n21225), .ZN(n21221) );
  OAI22_X1 U15095 ( .A1(n20759), .A2(n21204), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13872) );
  XNOR2_X1 U15096 ( .A(n13868), .B(n13872), .ZN(n13508) );
  AOI22_X1 U15097 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n21210), .B2(n20764), .ZN(
        n13503) );
  OAI21_X1 U15098 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n20764), .A(
        n13499), .ZN(n13500) );
  OAI22_X1 U15099 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21214), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13500), .ZN(n13505) );
  NOR2_X1 U15100 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21214), .ZN(
        n13501) );
  NAND2_X1 U15101 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13500), .ZN(
        n13506) );
  AOI22_X1 U15102 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13505), .B1(
        n13501), .B2(n13506), .ZN(n13871) );
  OAI21_X1 U15103 ( .B1(n13504), .B2(n13503), .A(n13871), .ZN(n13502) );
  AOI21_X1 U15104 ( .B1(n13504), .B2(n13503), .A(n13502), .ZN(n13869) );
  AOI21_X1 U15105 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n13506), .A(
        n13505), .ZN(n13507) );
  INV_X1 U15106 ( .A(n21192), .ZN(n21188) );
  NAND2_X1 U15107 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n20559), .ZN(n13509) );
  AOI211_X4 U15108 ( .C1(n21659), .C2(n21612), .A(n13513), .B(n13509), .ZN(
        n20546) );
  NOR3_X1 U15109 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_1__SCAN_IN), .ZN(n20176) );
  INV_X1 U15110 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n20175) );
  NAND2_X1 U15111 ( .A1(n20176), .A2(n20175), .ZN(n20183) );
  NOR2_X1 U15112 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n20183), .ZN(n20203) );
  INV_X1 U15113 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n20202) );
  NAND2_X1 U15114 ( .A1(n20203), .A2(n20202), .ZN(n20209) );
  NOR2_X1 U15115 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n20209), .ZN(n20232) );
  INV_X1 U15116 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n20231) );
  NAND2_X1 U15117 ( .A1(n20232), .A2(n20231), .ZN(n20241) );
  INV_X1 U15118 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n20252) );
  NAND2_X1 U15119 ( .A1(n20251), .A2(n20252), .ZN(n20269) );
  NOR2_X1 U15120 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n20269), .ZN(n20284) );
  INV_X1 U15121 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n20283) );
  NAND2_X1 U15122 ( .A1(n20284), .A2(n20283), .ZN(n20289) );
  NOR2_X1 U15123 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n20289), .ZN(n20305) );
  INV_X1 U15124 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n20308) );
  NAND2_X1 U15125 ( .A1(n20305), .A2(n20308), .ZN(n20319) );
  NOR2_X1 U15126 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n20319), .ZN(n20337) );
  INV_X1 U15127 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n20336) );
  NAND2_X1 U15128 ( .A1(n20337), .A2(n20336), .ZN(n20353) );
  NOR2_X1 U15129 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n20353), .ZN(n20372) );
  INV_X1 U15130 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n20378) );
  NAND2_X1 U15131 ( .A1(n20372), .A2(n20378), .ZN(n20379) );
  NOR2_X1 U15132 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n20379), .ZN(n20389) );
  INV_X1 U15133 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n20390) );
  NAND2_X1 U15134 ( .A1(n20389), .A2(n20390), .ZN(n20405) );
  NOR2_X1 U15135 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n20405), .ZN(n20419) );
  INV_X1 U15136 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n20418) );
  NAND2_X1 U15137 ( .A1(n20419), .A2(n20418), .ZN(n20426) );
  NOR2_X1 U15138 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n20426), .ZN(n20445) );
  INV_X1 U15139 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n20448) );
  NAND2_X1 U15140 ( .A1(n20445), .A2(n20448), .ZN(n20453) );
  NOR2_X1 U15141 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n20453), .ZN(n20474) );
  INV_X1 U15142 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n20473) );
  NAND2_X1 U15143 ( .A1(n20474), .A2(n20473), .ZN(n20481) );
  NOR2_X1 U15144 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n20481), .ZN(n20498) );
  INV_X1 U15145 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n20497) );
  NAND2_X1 U15146 ( .A1(n20498), .A2(n20497), .ZN(n20509) );
  NOR2_X1 U15147 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n20509), .ZN(n20521) );
  INV_X1 U15148 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n20524) );
  NAND2_X1 U15149 ( .A1(n20521), .A2(n20524), .ZN(n20522) );
  NOR2_X1 U15150 ( .A1(n20508), .A2(n20522), .ZN(n20543) );
  INV_X1 U15151 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n17495) );
  NAND2_X1 U15152 ( .A1(n20543), .A2(n17495), .ZN(n13519) );
  INV_X1 U15153 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n21658) );
  INV_X1 U15154 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n21618) );
  NAND2_X1 U15155 ( .A1(P3_STATE_REG_2__SCAN_IN), .A2(n21618), .ZN(n21664) );
  AOI21_X1 U15156 ( .B1(n18235), .B2(n21664), .A(n18230), .ZN(n20091) );
  OAI211_X1 U15157 ( .C1(n20559), .C2(n20091), .A(n21659), .B(n21612), .ZN(
        n21223) );
  NAND3_X1 U15158 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n13510) );
  NOR2_X1 U15159 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n21235) );
  NAND2_X1 U15160 ( .A1(n21098), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18770) );
  OR2_X1 U15161 ( .A1(n21225), .A2(n18770), .ZN(n21241) );
  INV_X1 U15162 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n20471) );
  INV_X1 U15163 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18223) );
  INV_X1 U15164 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n20366) );
  INV_X1 U15165 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n20344) );
  INV_X1 U15166 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n20343) );
  INV_X1 U15167 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n20263) );
  INV_X1 U15168 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n20920) );
  INV_X1 U15169 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n20239) );
  INV_X1 U15170 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n20875) );
  INV_X1 U15171 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n20186) );
  NAND3_X1 U15172 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .A3(P3_REIP_REG_1__SCAN_IN), .ZN(n20182) );
  NOR2_X1 U15173 ( .A1(n20186), .A2(n20182), .ZN(n20196) );
  NAND2_X1 U15174 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n20196), .ZN(n20207) );
  NOR2_X1 U15175 ( .A1(n20875), .A2(n20207), .ZN(n20226) );
  NAND2_X1 U15176 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n20226), .ZN(n20240) );
  NOR2_X1 U15177 ( .A1(n20239), .A2(n20240), .ZN(n20257) );
  NAND2_X1 U15178 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n20257), .ZN(n20262) );
  NOR3_X1 U15179 ( .A1(n20263), .A2(n20920), .A3(n20262), .ZN(n20290) );
  NAND2_X1 U15180 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n20290), .ZN(n20342) );
  NOR3_X1 U15181 ( .A1(n20344), .A2(n20343), .A3(n20342), .ZN(n20320) );
  NAND3_X1 U15182 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .A3(n20320), .ZN(n20367) );
  NOR2_X1 U15183 ( .A1(n20366), .A2(n20367), .ZN(n20381) );
  NAND2_X1 U15184 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n20381), .ZN(n20392) );
  NOR2_X1 U15185 ( .A1(n18223), .A2(n20392), .ZN(n20414) );
  AND2_X1 U15186 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n20414), .ZN(n20404) );
  NAND4_X1 U15187 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(P3_REIP_REG_22__SCAN_IN), 
        .A3(P3_REIP_REG_21__SCAN_IN), .A4(n20404), .ZN(n20439) );
  INV_X1 U15188 ( .A(n20439), .ZN(n20458) );
  NAND2_X1 U15189 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n20458), .ZN(n20466) );
  NOR2_X1 U15190 ( .A1(n20471), .A2(n20466), .ZN(n20482) );
  NAND2_X1 U15191 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n20482), .ZN(n13511) );
  NAND2_X1 U15192 ( .A1(n20440), .A2(n13511), .ZN(n20483) );
  NAND2_X1 U15193 ( .A1(n20548), .A2(n20483), .ZN(n20505) );
  AOI21_X1 U15194 ( .B1(n20440), .B2(n13510), .A(n20505), .ZN(n20539) );
  INV_X1 U15195 ( .A(n20539), .ZN(n20527) );
  INV_X1 U15196 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n20519) );
  NOR2_X1 U15197 ( .A1(n20549), .A2(n13511), .ZN(n20507) );
  NAND2_X1 U15198 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n20507), .ZN(n20511) );
  NOR2_X1 U15199 ( .A1(n20519), .A2(n20511), .ZN(n20529) );
  NAND2_X1 U15200 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n20529), .ZN(n13515) );
  NOR2_X1 U15201 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n13515), .ZN(n20541) );
  OAI21_X1 U15202 ( .B1(n20527), .B2(n20541), .A(P3_REIP_REG_31__SCAN_IN), 
        .ZN(n13512) );
  INV_X1 U15203 ( .A(n21223), .ZN(n13514) );
  AOI211_X4 U15204 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n20559), .A(n13514), .B(
        n13513), .ZN(n20547) );
  INV_X1 U15205 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n21037) );
  NOR3_X1 U15206 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n13515), .A3(n21037), 
        .ZN(n13516) );
  AOI21_X1 U15207 ( .B1(n20547), .B2(P3_EBX_REG_31__SCAN_IN), .A(n13516), .ZN(
        n13518) );
  OR2_X1 U15208 ( .A1(n20537), .A2(n17940), .ZN(n13517) );
  NAND2_X1 U15209 ( .A1(n16973), .A2(n21917), .ZN(n21253) );
  INV_X1 U15210 ( .A(n21253), .ZN(n21596) );
  AOI21_X1 U15211 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21596), .A(n16946), 
        .ZN(n16972) );
  AOI21_X1 U15212 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(n13522), .A(
        P1_STATE2_REG_0__SCAN_IN), .ZN(n13528) );
  AND2_X1 U15213 ( .A1(n13523), .A2(n12623), .ZN(n16162) );
  NAND2_X1 U15214 ( .A1(n14804), .A2(n16162), .ZN(n14827) );
  INV_X1 U15215 ( .A(n13524), .ZN(n13525) );
  NAND2_X1 U15216 ( .A1(n13525), .A2(n15620), .ZN(n13526) );
  NAND2_X1 U15217 ( .A1(n14827), .A2(n13526), .ZN(n14658) );
  NAND2_X1 U15218 ( .A1(n14804), .A2(n12614), .ZN(n14802) );
  INV_X1 U15219 ( .A(n14802), .ZN(n13527) );
  OR2_X1 U15220 ( .A1(n13654), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21378) );
  INV_X1 U15221 ( .A(n13529), .ZN(n13530) );
  NAND2_X1 U15222 ( .A1(n13530), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13531) );
  INV_X1 U15223 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13640) );
  XNOR2_X1 U15224 ( .A(n13531), .B(n13640), .ZN(n15100) );
  OR2_X1 U15225 ( .A1(n15100), .A2(n16973), .ZN(n13532) );
  NAND2_X1 U15226 ( .A1(n13660), .A2(n21541), .ZN(n13648) );
  INV_X1 U15227 ( .A(n13663), .ZN(n15162) );
  OAI22_X1 U15228 ( .A1(n14684), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        P1_EBX_REG_30__SCAN_IN), .B2(n10976), .ZN(n15630) );
  INV_X1 U15229 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13533) );
  NAND2_X1 U15230 ( .A1(n13606), .A2(n13533), .ZN(n13536) );
  INV_X1 U15231 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n21412) );
  NAND2_X1 U15232 ( .A1(n14687), .A2(n21412), .ZN(n13535) );
  NAND3_X1 U15233 ( .A1(n13536), .A2(n13535), .A3(n10979), .ZN(n13537) );
  NAND2_X1 U15234 ( .A1(n11376), .A2(n13537), .ZN(n13541) );
  NAND2_X1 U15235 ( .A1(n13606), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13540) );
  INV_X1 U15236 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13538) );
  NAND2_X1 U15237 ( .A1(n10979), .A2(n13538), .ZN(n13539) );
  NAND2_X1 U15238 ( .A1(n13540), .A2(n13539), .ZN(n14685) );
  INV_X1 U15239 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13683) );
  NAND2_X1 U15240 ( .A1(n13606), .A2(n13683), .ZN(n13545) );
  INV_X1 U15241 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13542) );
  NAND2_X1 U15242 ( .A1(n14687), .A2(n13542), .ZN(n13544) );
  NAND3_X1 U15243 ( .A1(n13545), .A2(n13544), .A3(n10979), .ZN(n13546) );
  OAI21_X1 U15244 ( .B1(P1_EBX_REG_2__SCAN_IN), .B2(n13620), .A(n13546), .ZN(
        n14837) );
  MUX2_X1 U15245 ( .A(n13612), .B(n10979), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n13549) );
  OR2_X1 U15246 ( .A1(n14684), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13548) );
  INV_X1 U15247 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n15016) );
  NAND2_X1 U15248 ( .A1(n13617), .A2(n15016), .ZN(n13552) );
  INV_X1 U15249 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13698) );
  NAND2_X1 U15250 ( .A1(n13606), .A2(n13698), .ZN(n13550) );
  OAI211_X1 U15251 ( .C1(n10976), .C2(P1_EBX_REG_4__SCAN_IN), .A(n13550), .B(
        n10979), .ZN(n13551) );
  MUX2_X1 U15252 ( .A(n13612), .B(n10979), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n13553) );
  OAI21_X1 U15253 ( .B1(n14684), .B2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n13553), .ZN(n15082) );
  MUX2_X1 U15254 ( .A(n13617), .B(n13616), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n13554) );
  INV_X1 U15255 ( .A(n13554), .ZN(n13557) );
  NAND2_X1 U15256 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n10976), .ZN(
        n13555) );
  AND2_X1 U15257 ( .A1(n13595), .A2(n13555), .ZN(n13556) );
  NAND2_X1 U15258 ( .A1(n13557), .A2(n13556), .ZN(n15089) );
  OR2_X1 U15259 ( .A1(n14684), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13559) );
  MUX2_X1 U15260 ( .A(n13612), .B(n10979), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n13558) );
  AND2_X1 U15261 ( .A1(n13559), .A2(n13558), .ZN(n15275) );
  MUX2_X1 U15262 ( .A(n13617), .B(n13616), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n13562) );
  NAND2_X1 U15263 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n10976), .ZN(
        n13560) );
  NAND2_X1 U15264 ( .A1(n13595), .A2(n13560), .ZN(n13561) );
  NOR2_X1 U15265 ( .A1(n13562), .A2(n13561), .ZN(n15398) );
  OR2_X1 U15266 ( .A1(n13612), .A2(P1_EBX_REG_9__SCAN_IN), .ZN(n13565) );
  NAND2_X1 U15267 ( .A1(n10979), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13563) );
  OAI211_X1 U15268 ( .C1(n10976), .C2(P1_EBX_REG_9__SCAN_IN), .A(n13606), .B(
        n13563), .ZN(n13564) );
  NAND2_X1 U15269 ( .A1(n13565), .A2(n13564), .ZN(n15445) );
  MUX2_X1 U15270 ( .A(n13617), .B(n13616), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n13568) );
  NAND2_X1 U15271 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n10976), .ZN(
        n13566) );
  NAND2_X1 U15272 ( .A1(n13595), .A2(n13566), .ZN(n13567) );
  NOR2_X1 U15273 ( .A1(n13568), .A2(n13567), .ZN(n15490) );
  OR2_X1 U15274 ( .A1(n13612), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n13571) );
  NAND2_X1 U15275 ( .A1(n10979), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13569) );
  OAI211_X1 U15276 ( .C1(n10976), .C2(P1_EBX_REG_11__SCAN_IN), .A(n13606), .B(
        n13569), .ZN(n13570) );
  NAND2_X1 U15277 ( .A1(n15524), .A2(n15523), .ZN(n15535) );
  INV_X1 U15278 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n21521) );
  NAND2_X1 U15279 ( .A1(n13617), .A2(n21521), .ZN(n13574) );
  INV_X1 U15280 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n21315) );
  NAND2_X1 U15281 ( .A1(n13606), .A2(n21315), .ZN(n13572) );
  OAI211_X1 U15282 ( .C1(n10976), .C2(P1_EBX_REG_12__SCAN_IN), .A(n13572), .B(
        n10979), .ZN(n13573) );
  MUX2_X1 U15283 ( .A(n13612), .B(n10979), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n13576) );
  OR2_X1 U15284 ( .A1(n14684), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n13575) );
  NAND2_X1 U15285 ( .A1(n13576), .A2(n13575), .ZN(n15791) );
  INV_X1 U15286 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n21272) );
  NAND2_X1 U15287 ( .A1(n13606), .A2(n21272), .ZN(n13578) );
  INV_X1 U15288 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n15777) );
  NAND2_X1 U15289 ( .A1(n14687), .A2(n15777), .ZN(n13577) );
  NAND3_X1 U15290 ( .A1(n13578), .A2(n13577), .A3(n10979), .ZN(n13579) );
  OAI21_X1 U15291 ( .B1(P1_EBX_REG_14__SCAN_IN), .B2(n13620), .A(n13579), .ZN(
        n15543) );
  OR2_X1 U15292 ( .A1(n14684), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n13581) );
  MUX2_X1 U15293 ( .A(n13612), .B(n10979), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n13580) );
  AND2_X1 U15294 ( .A1(n13581), .A2(n13580), .ZN(n15771) );
  MUX2_X1 U15295 ( .A(n13617), .B(n13616), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n13584) );
  NAND2_X1 U15296 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n10976), .ZN(
        n13582) );
  NAND2_X1 U15297 ( .A1(n13595), .A2(n13582), .ZN(n13583) );
  NOR2_X1 U15298 ( .A1(n13584), .A2(n13583), .ZN(n15828) );
  OR2_X1 U15299 ( .A1(n13612), .A2(P1_EBX_REG_17__SCAN_IN), .ZN(n13587) );
  NAND2_X1 U15300 ( .A1(n10979), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13585) );
  OAI211_X1 U15301 ( .C1(n10976), .C2(P1_EBX_REG_17__SCAN_IN), .A(n13606), .B(
        n13585), .ZN(n13586) );
  NAND2_X1 U15302 ( .A1(n13587), .A2(n13586), .ZN(n15822) );
  MUX2_X1 U15303 ( .A(n13617), .B(n13616), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n13588) );
  INV_X1 U15304 ( .A(n13588), .ZN(n13591) );
  NAND2_X1 U15305 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n10976), .ZN(
        n13589) );
  AND2_X1 U15306 ( .A1(n13595), .A2(n13589), .ZN(n13590) );
  NAND2_X1 U15307 ( .A1(n13591), .A2(n13590), .ZN(n15815) );
  MUX2_X1 U15308 ( .A(n13612), .B(n10979), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n13593) );
  OR2_X1 U15309 ( .A1(n14684), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13592) );
  AND2_X1 U15310 ( .A1(n13593), .A2(n13592), .ZN(n15760) );
  MUX2_X1 U15311 ( .A(n13617), .B(n13616), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n13597) );
  NAND2_X1 U15312 ( .A1(n10976), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13594) );
  NAND2_X1 U15313 ( .A1(n13595), .A2(n13594), .ZN(n13596) );
  NOR2_X1 U15314 ( .A1(n13597), .A2(n13596), .ZN(n15746) );
  MUX2_X1 U15315 ( .A(n13612), .B(n10979), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n13599) );
  OR2_X1 U15316 ( .A1(n14684), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n13598) );
  NAND2_X1 U15317 ( .A1(n13599), .A2(n13598), .ZN(n15729) );
  MUX2_X1 U15318 ( .A(n13617), .B(n13616), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n13600) );
  NOR2_X1 U15319 ( .A1(n13600), .A2(n11382), .ZN(n15711) );
  MUX2_X1 U15320 ( .A(n13612), .B(n13543), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n13602) );
  OR2_X1 U15321 ( .A1(n14684), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n13601) );
  AND2_X1 U15322 ( .A1(n13602), .A2(n13601), .ZN(n15698) );
  INV_X1 U15323 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16118) );
  NAND2_X1 U15324 ( .A1(n13606), .A2(n16118), .ZN(n13603) );
  OAI211_X1 U15325 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n10976), .A(n13603), .B(
        n10979), .ZN(n13604) );
  OAI21_X1 U15326 ( .B1(P1_EBX_REG_24__SCAN_IN), .B2(n13620), .A(n13604), .ZN(
        n15687) );
  AND2_X2 U15327 ( .A1(n11020), .A2(n15687), .ZN(n15689) );
  OR2_X1 U15328 ( .A1(n13612), .A2(P1_EBX_REG_25__SCAN_IN), .ZN(n13608) );
  NAND2_X1 U15329 ( .A1(n10979), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n13605) );
  OAI211_X1 U15330 ( .C1(P1_EBX_REG_25__SCAN_IN), .C2(n10976), .A(n13606), .B(
        n13605), .ZN(n13607) );
  AND2_X1 U15331 ( .A1(n13608), .A2(n13607), .ZN(n15676) );
  MUX2_X1 U15332 ( .A(n13617), .B(n13616), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n13609) );
  INV_X1 U15333 ( .A(n13609), .ZN(n13611) );
  NAND2_X1 U15334 ( .A1(n10976), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n13610) );
  NAND2_X1 U15335 ( .A1(n13611), .A2(n13610), .ZN(n15655) );
  MUX2_X1 U15336 ( .A(n13612), .B(n10979), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n13614) );
  OR2_X1 U15337 ( .A1(n14684), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n13613) );
  AND2_X1 U15338 ( .A1(n13614), .A2(n13613), .ZN(n15656) );
  NAND2_X1 U15339 ( .A1(n15655), .A2(n15656), .ZN(n13615) );
  MUX2_X1 U15340 ( .A(n13617), .B(n13616), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n13619) );
  AND2_X1 U15341 ( .A1(n10976), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n13618) );
  NOR2_X1 U15342 ( .A1(n13619), .A2(n13618), .ZN(n15638) );
  OAI22_X1 U15343 ( .A1(n14684), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        P1_EBX_REG_29__SCAN_IN), .B2(n10976), .ZN(n15627) );
  OAI22_X1 U15344 ( .A1(n15627), .A2(n13547), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n13620), .ZN(n15587) );
  MUX2_X1 U15345 ( .A(n15630), .B(n13543), .S(n15629), .Z(n13622) );
  OAI22_X1 U15346 ( .A1(n14684), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        P1_EBX_REG_31__SCAN_IN), .B2(n10976), .ZN(n13621) );
  XNOR2_X2 U15347 ( .A(n13622), .B(n13621), .ZN(n16022) );
  NAND2_X1 U15348 ( .A1(n13623), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15095) );
  AND2_X1 U15349 ( .A1(n12623), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13636) );
  NAND2_X1 U15350 ( .A1(n21622), .A2(n21936), .ZN(n16941) );
  NAND2_X1 U15351 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .ZN(n21433) );
  NAND4_X1 U15352 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_4__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n13624)
         );
  NOR2_X1 U15353 ( .A1(n21433), .A2(n13624), .ZN(n21465) );
  NAND2_X1 U15354 ( .A1(n21465), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n21485) );
  INV_X1 U15355 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n21487) );
  NOR2_X1 U15356 ( .A1(n21485), .A2(n21487), .ZN(n15448) );
  NAND3_X1 U15357 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_19__SCAN_IN), .ZN(n13627) );
  NAND4_X1 U15358 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .A3(P1_REIP_REG_13__SCAN_IN), .A4(P1_REIP_REG_10__SCAN_IN), .ZN(n13626) );
  NAND4_X1 U15359 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .A3(P1_REIP_REG_12__SCAN_IN), .A4(P1_REIP_REG_17__SCAN_IN), .ZN(n13625) );
  NOR3_X1 U15360 ( .A1(n13627), .A2(n13626), .A3(n13625), .ZN(n15745) );
  NAND3_X1 U15361 ( .A1(n15448), .A2(n15745), .A3(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n15714) );
  NOR2_X1 U15362 ( .A1(n21411), .A2(n15714), .ZN(n15730) );
  NAND2_X1 U15363 ( .A1(n15730), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15717) );
  NAND3_X1 U15364 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(P1_REIP_REG_23__SCAN_IN), 
        .A3(P1_REIP_REG_25__SCAN_IN), .ZN(n15666) );
  INV_X1 U15365 ( .A(n15666), .ZN(n13628) );
  NAND3_X1 U15366 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .A3(n13628), .ZN(n13629) );
  NOR2_X1 U15367 ( .A1(n15717), .A2(n13629), .ZN(n15650) );
  AND2_X1 U15368 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n13630) );
  NAND2_X1 U15369 ( .A1(n15650), .A2(n13630), .ZN(n15625) );
  NAND2_X1 U15370 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n13631) );
  NOR2_X1 U15371 ( .A1(n15625), .A2(n13631), .ZN(n13641) );
  INV_X1 U15372 ( .A(n13638), .ZN(n13635) );
  INV_X1 U15373 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n13632) );
  NAND2_X1 U15374 ( .A1(n13633), .A2(n13632), .ZN(n21633) );
  NAND2_X1 U15375 ( .A1(n16174), .A2(n21633), .ZN(n14843) );
  INV_X1 U15376 ( .A(n16941), .ZN(n13634) );
  NAND2_X1 U15377 ( .A1(n14843), .A2(n13634), .ZN(n13639) );
  OR2_X2 U15378 ( .A1(n13635), .A2(n13639), .ZN(n21459) );
  NOR2_X1 U15379 ( .A1(n13641), .A2(n21495), .ZN(n15634) );
  INV_X1 U15380 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n15801) );
  INV_X1 U15381 ( .A(n13636), .ZN(n13637) );
  OAI22_X1 U15382 ( .A1(n21566), .A2(n13640), .B1(n15801), .B2(n21559), .ZN(
        n13644) );
  INV_X1 U15383 ( .A(n13641), .ZN(n13642) );
  NOR3_X1 U15384 ( .A1(n13642), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n21459), 
        .ZN(n13643) );
  AOI211_X1 U15385 ( .C1(n15634), .C2(P1_REIP_REG_31__SCAN_IN), .A(n13644), 
        .B(n13643), .ZN(n13645) );
  NAND2_X1 U15386 ( .A1(n13648), .A2(n13647), .ZN(P1_U2809) );
  NAND3_X1 U15387 ( .A1(n16946), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n21589) );
  INV_X1 U15388 ( .A(n21589), .ZN(n13649) );
  NOR2_X1 U15389 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n21876) );
  OR2_X1 U15390 ( .A1(n14717), .A2(n22148), .ZN(n13651) );
  AND2_X1 U15391 ( .A1(n13651), .A2(n13650), .ZN(n14716) );
  NAND2_X1 U15392 ( .A1(n15577), .A2(n14719), .ZN(n13652) );
  AND3_X1 U15393 ( .A1(n14716), .A2(n12626), .A3(n13652), .ZN(n14706) );
  NAND2_X1 U15394 ( .A1(n14706), .A2(n13653), .ZN(n14859) );
  INV_X1 U15395 ( .A(n21876), .ZN(n21919) );
  NAND2_X1 U15396 ( .A1(n21919), .A2(n13654), .ZN(n21256) );
  AND2_X1 U15397 ( .A1(n21256), .A2(n16946), .ZN(n13655) );
  NAND2_X1 U15398 ( .A1(n16946), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n16944) );
  NAND2_X1 U15399 ( .A1(n21936), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13656) );
  AND2_X1 U15400 ( .A1(n16944), .A2(n13656), .ZN(n19952) );
  INV_X1 U15401 ( .A(n19952), .ZN(n13657) );
  INV_X1 U15402 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n17189) );
  NOR2_X1 U15403 ( .A1(n21378), .A2(n17189), .ZN(n16051) );
  AOI21_X1 U15404 ( .B1(n20015), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n16051), .ZN(n13658) );
  OAI21_X1 U15405 ( .B1(n20025), .B2(n15100), .A(n13658), .ZN(n13659) );
  AOI21_X1 U15406 ( .B1(n13660), .B2(n20021), .A(n13659), .ZN(n13774) );
  NAND2_X1 U15407 ( .A1(n13675), .A2(n13667), .ZN(n13661) );
  NAND2_X1 U15408 ( .A1(n13661), .A2(n13662), .ZN(n13687) );
  OAI21_X1 U15409 ( .B1(n13662), .B2(n13661), .A(n13687), .ZN(n13664) );
  AND2_X1 U15410 ( .A1(n14719), .A2(n13663), .ZN(n13673) );
  AOI21_X1 U15411 ( .B1(n13664), .B2(n14800), .A(n13673), .ZN(n13665) );
  NAND2_X1 U15412 ( .A1(n13666), .A2(n13720), .ZN(n13672) );
  INV_X1 U15413 ( .A(n13667), .ZN(n13668) );
  XNOR2_X1 U15414 ( .A(n13668), .B(n13675), .ZN(n13670) );
  NAND2_X1 U15415 ( .A1(n15151), .A2(n15596), .ZN(n13669) );
  AOI21_X1 U15416 ( .B1(n13670), .B2(n14800), .A(n13669), .ZN(n13671) );
  NAND2_X1 U15417 ( .A1(n21850), .A2(n13720), .ZN(n13678) );
  INV_X1 U15418 ( .A(n14800), .ZN(n21250) );
  INV_X1 U15419 ( .A(n13673), .ZN(n13674) );
  OAI21_X1 U15420 ( .B1(n21250), .B2(n13675), .A(n13674), .ZN(n13676) );
  INV_X1 U15421 ( .A(n13676), .ZN(n13677) );
  NAND2_X1 U15422 ( .A1(n13678), .A2(n13677), .ZN(n19947) );
  NAND2_X1 U15423 ( .A1(n19947), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13679) );
  NAND2_X1 U15425 ( .A1(n14842), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13682) );
  INV_X1 U15426 ( .A(n13679), .ZN(n19948) );
  NAND2_X1 U15427 ( .A1(n13680), .A2(n19948), .ZN(n13681) );
  NAND2_X1 U15428 ( .A1(n14938), .A2(n14937), .ZN(n13686) );
  NAND2_X1 U15429 ( .A1(n13684), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13685) );
  NAND2_X2 U15430 ( .A1(n13686), .A2(n13685), .ZN(n13691) );
  INV_X1 U15431 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n14959) );
  OR2_X1 U15432 ( .A1(n21769), .A2(n13732), .ZN(n13690) );
  NAND2_X1 U15433 ( .A1(n13687), .A2(n13688), .ZN(n13705) );
  OAI211_X1 U15434 ( .C1(n13688), .C2(n13687), .A(n13705), .B(n14800), .ZN(
        n13689) );
  NAND2_X1 U15435 ( .A1(n13690), .A2(n13689), .ZN(n14955) );
  NAND2_X1 U15436 ( .A1(n14956), .A2(n14955), .ZN(n13693) );
  NAND2_X1 U15437 ( .A1(n13691), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13692) );
  NAND2_X1 U15438 ( .A1(n13693), .A2(n13692), .ZN(n14982) );
  NAND2_X1 U15439 ( .A1(n13694), .A2(n13720), .ZN(n13697) );
  XNOR2_X1 U15440 ( .A(n13705), .B(n13703), .ZN(n13695) );
  NAND2_X1 U15441 ( .A1(n13695), .A2(n14800), .ZN(n13696) );
  NAND2_X1 U15442 ( .A1(n13697), .A2(n13696), .ZN(n13699) );
  XNOR2_X1 U15443 ( .A(n13699), .B(n13698), .ZN(n14981) );
  NAND2_X1 U15444 ( .A1(n14982), .A2(n14981), .ZN(n13701) );
  NAND2_X1 U15445 ( .A1(n13699), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13700) );
  NAND2_X1 U15446 ( .A1(n13702), .A2(n13720), .ZN(n13709) );
  INV_X1 U15447 ( .A(n13703), .ZN(n13704) );
  NOR2_X1 U15448 ( .A1(n13705), .A2(n13704), .ZN(n13707) );
  NAND2_X1 U15449 ( .A1(n13707), .A2(n13706), .ZN(n13722) );
  OAI211_X1 U15450 ( .C1(n13707), .C2(n13706), .A(n13722), .B(n14800), .ZN(
        n13708) );
  NAND2_X1 U15451 ( .A1(n13709), .A2(n13708), .ZN(n13710) );
  XNOR2_X1 U15452 ( .A(n13710), .B(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n19956) );
  OR2_X1 U15453 ( .A1(n13710), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13711) );
  NAND2_X1 U15454 ( .A1(n13712), .A2(n13711), .ZN(n15253) );
  NAND3_X1 U15455 ( .A1(n13713), .A2(n13720), .A3(n13714), .ZN(n13717) );
  XNOR2_X1 U15456 ( .A(n13722), .B(n13723), .ZN(n13715) );
  NAND2_X1 U15457 ( .A1(n13715), .A2(n14800), .ZN(n13716) );
  NAND2_X1 U15458 ( .A1(n13717), .A2(n13716), .ZN(n13718) );
  XNOR2_X1 U15459 ( .A(n13718), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15252) );
  OR2_X2 U15460 ( .A1(n15253), .A2(n15252), .ZN(n15255) );
  NAND2_X1 U15461 ( .A1(n13718), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13719) );
  NAND2_X2 U15462 ( .A1(n15255), .A2(n13719), .ZN(n15402) );
  NAND2_X1 U15463 ( .A1(n13721), .A2(n13720), .ZN(n13727) );
  INV_X1 U15464 ( .A(n13722), .ZN(n13724) );
  NAND2_X1 U15465 ( .A1(n13724), .A2(n13723), .ZN(n13736) );
  XNOR2_X1 U15466 ( .A(n13736), .B(n13737), .ZN(n13725) );
  NAND2_X1 U15467 ( .A1(n13725), .A2(n14800), .ZN(n13726) );
  NAND2_X1 U15468 ( .A1(n13727), .A2(n13726), .ZN(n13729) );
  INV_X1 U15469 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n13728) );
  XNOR2_X1 U15470 ( .A(n13729), .B(n13728), .ZN(n15401) );
  NAND2_X1 U15471 ( .A1(n13729), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13730) );
  NOR2_X1 U15472 ( .A1(n13733), .A2(n13732), .ZN(n13734) );
  INV_X1 U15473 ( .A(n13736), .ZN(n13738) );
  NAND3_X1 U15474 ( .A1(n13738), .A2(n14800), .A3(n13737), .ZN(n13739) );
  NAND2_X1 U15475 ( .A1(n10965), .A2(n13739), .ZN(n13740) );
  XNOR2_X1 U15476 ( .A(n13740), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15425) );
  INV_X1 U15477 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15466) );
  XNOR2_X1 U15478 ( .A(n13735), .B(n15466), .ZN(n15456) );
  INV_X1 U15479 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21274) );
  NAND2_X1 U15480 ( .A1(n13735), .A2(n21274), .ZN(n13741) );
  NAND2_X1 U15481 ( .A1(n19992), .A2(n13741), .ZN(n16014) );
  NAND3_X1 U15482 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n13742) );
  AND2_X1 U15483 ( .A1(n13735), .A2(n13742), .ZN(n13743) );
  NAND2_X1 U15484 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21353) );
  INV_X1 U15485 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21352) );
  NOR2_X1 U15486 ( .A1(n21353), .A2(n21352), .ZN(n21348) );
  INV_X1 U15487 ( .A(n21348), .ZN(n13744) );
  NAND2_X1 U15488 ( .A1(n20007), .A2(n13744), .ZN(n13745) );
  NAND3_X1 U15489 ( .A1(n19974), .A2(n16000), .A3(n13745), .ZN(n13751) );
  OR2_X1 U15490 ( .A1(n13735), .A2(n21272), .ZN(n13746) );
  NAND2_X1 U15491 ( .A1(n19992), .A2(n13746), .ZN(n15990) );
  NOR2_X1 U15492 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16010) );
  AND2_X1 U15493 ( .A1(n16010), .A2(n21315), .ZN(n13747) );
  NOR2_X1 U15494 ( .A1(n13735), .A2(n13747), .ZN(n15989) );
  NOR2_X1 U15495 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n13748) );
  INV_X1 U15496 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21361) );
  OAI21_X1 U15497 ( .B1(n13748), .B2(n13735), .A(n20005), .ZN(n13749) );
  NOR2_X1 U15498 ( .A1(n15999), .A2(n13749), .ZN(n13750) );
  NAND2_X2 U15499 ( .A1(n13751), .A2(n13750), .ZN(n20018) );
  AND2_X1 U15500 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16134) );
  NAND2_X1 U15501 ( .A1(n16134), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n21381) );
  INV_X1 U15502 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21343) );
  NOR2_X1 U15503 ( .A1(n21381), .A2(n21343), .ZN(n13752) );
  NAND2_X1 U15504 ( .A1(n20018), .A2(n13752), .ZN(n13753) );
  INV_X1 U15505 ( .A(n20018), .ZN(n13754) );
  INV_X1 U15506 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n16133) );
  INV_X1 U15507 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n21373) );
  INV_X1 U15508 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15964) );
  INV_X1 U15509 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16113) );
  INV_X1 U15510 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n16104) );
  NAND3_X1 U15511 ( .A1(n16113), .A2(n16104), .A3(n16118), .ZN(n15906) );
  NAND2_X1 U15512 ( .A1(n13756), .A2(n19975), .ZN(n13759) );
  AND2_X1 U15513 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16105) );
  NAND2_X1 U15514 ( .A1(n16105), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16045) );
  NAND2_X1 U15515 ( .A1(n20009), .A2(n16045), .ZN(n15905) );
  NAND2_X1 U15516 ( .A1(n13757), .A2(n20009), .ZN(n15933) );
  AND2_X1 U15517 ( .A1(n15905), .A2(n15933), .ZN(n13758) );
  INV_X1 U15518 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n16037) );
  NOR2_X1 U15519 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16077) );
  AND2_X1 U15520 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16078) );
  INV_X1 U15521 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13765) );
  AND2_X1 U15522 ( .A1(n20009), .A2(n13765), .ZN(n13775) );
  INV_X1 U15523 ( .A(n13775), .ZN(n13760) );
  INV_X1 U15524 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n16038) );
  XNOR2_X1 U15525 ( .A(n20009), .B(n16038), .ZN(n13763) );
  INV_X1 U15526 ( .A(n13763), .ZN(n13762) );
  INV_X1 U15527 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16048) );
  NAND2_X1 U15528 ( .A1(n20009), .A2(n16048), .ZN(n13766) );
  NAND2_X1 U15529 ( .A1(n13762), .A2(n13766), .ZN(n13770) );
  NOR2_X1 U15530 ( .A1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13764) );
  OAI211_X1 U15531 ( .C1(n13764), .C2(n20009), .A(n13771), .B(n13763), .ZN(
        n13769) );
  OR2_X1 U15532 ( .A1(n20009), .A2(n13765), .ZN(n15894) );
  OAI211_X1 U15533 ( .C1(n20009), .C2(n16048), .A(n15894), .B(n13766), .ZN(
        n13767) );
  NAND2_X1 U15534 ( .A1(n13767), .A2(n16038), .ZN(n13768) );
  OAI211_X1 U15535 ( .C1(n13771), .C2(n13770), .A(n13769), .B(n13768), .ZN(
        n16054) );
  INV_X1 U15536 ( .A(n16054), .ZN(n13772) );
  NAND2_X1 U15537 ( .A1(n13772), .A2(n20020), .ZN(n13773) );
  NAND2_X1 U15538 ( .A1(n13774), .A2(n13773), .ZN(P1_U2968) );
  INV_X1 U15539 ( .A(n15894), .ZN(n13776) );
  NOR2_X1 U15540 ( .A1(n13776), .A2(n13775), .ZN(n13778) );
  XOR2_X1 U15541 ( .A(n13778), .B(n13777), .Z(n16074) );
  NAND2_X1 U15542 ( .A1(n21390), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n16067) );
  OAI21_X1 U15543 ( .B1(n19983), .B2(n15588), .A(n16067), .ZN(n13782) );
  AOI21_X1 U15544 ( .B1(n20000), .B2(n15591), .A(n13782), .ZN(n13783) );
  INV_X1 U15545 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n13784) );
  INV_X1 U15546 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16558) );
  INV_X1 U15547 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18394) );
  NAND2_X1 U15548 ( .A1(n13803), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n13805) );
  INV_X1 U15549 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n16497) );
  INV_X1 U15550 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n16482) );
  INV_X1 U15551 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n16461) );
  AND2_X1 U15552 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n13786) );
  INV_X1 U15553 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n18512) );
  INV_X1 U15554 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n13820) );
  INV_X1 U15555 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16360) );
  NAND2_X1 U15556 ( .A1(n13823), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13787) );
  XNOR2_X1 U15557 ( .A(n13787), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14469) );
  AOI21_X1 U15558 ( .B1(n16569), .B2(n13788), .A(n13789), .ZN(n18350) );
  NOR2_X1 U15559 ( .A1(n16581), .A2(n13790), .ZN(n13798) );
  AOI21_X1 U15560 ( .B1(n16581), .B2(n13790), .A(n13798), .ZN(n18327) );
  AOI21_X1 U15561 ( .B1(n16593), .B2(n13791), .A(n13792), .ZN(n18301) );
  AOI21_X1 U15562 ( .B1(n17223), .B2(n13793), .A(n13794), .ZN(n18284) );
  INV_X1 U15563 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n15293) );
  NAND2_X1 U15564 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13796) );
  NOR2_X1 U15565 ( .A1(n15293), .A2(n13796), .ZN(n13797) );
  AOI21_X1 U15566 ( .B1(n15293), .B2(n13796), .A(n13797), .ZN(n15295) );
  OAI22_X1 U15567 ( .A1(n18669), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n13795) );
  INV_X1 U15568 ( .A(n13795), .ZN(n18253) );
  AOI22_X1 U15569 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n11712), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18669), .ZN(n15067) );
  NOR2_X1 U15570 ( .A1(n18253), .A2(n15067), .ZN(n15066) );
  OAI21_X1 U15571 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n13796), .ZN(n15032) );
  NAND2_X1 U15572 ( .A1(n15066), .A2(n15032), .ZN(n15044) );
  NOR2_X1 U15573 ( .A1(n15295), .A2(n15044), .ZN(n18271) );
  OAI21_X1 U15574 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13797), .A(
        n13793), .ZN(n18270) );
  NAND2_X1 U15575 ( .A1(n18271), .A2(n18270), .ZN(n18282) );
  NOR2_X1 U15576 ( .A1(n18284), .A2(n18282), .ZN(n18293) );
  OAI21_X1 U15577 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13794), .A(
        n13791), .ZN(n18294) );
  NAND2_X1 U15578 ( .A1(n18293), .A2(n18294), .ZN(n18300) );
  NOR2_X1 U15579 ( .A1(n18301), .A2(n18300), .ZN(n18315) );
  OAI21_X1 U15580 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n13792), .A(
        n13790), .ZN(n18316) );
  NAND2_X1 U15581 ( .A1(n18315), .A2(n18316), .ZN(n18325) );
  NOR2_X1 U15582 ( .A1(n18327), .A2(n18325), .ZN(n18332) );
  OAI21_X1 U15583 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n13798), .A(
        n13788), .ZN(n18334) );
  NAND2_X1 U15584 ( .A1(n18332), .A2(n18334), .ZN(n18348) );
  NOR2_X1 U15585 ( .A1(n18350), .A2(n18348), .ZN(n18360) );
  OAI21_X1 U15586 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n13789), .A(
        n13799), .ZN(n18362) );
  NAND2_X1 U15587 ( .A1(n18360), .A2(n18362), .ZN(n14483) );
  AOI21_X1 U15588 ( .B1(n16558), .B2(n13799), .A(n13800), .ZN(n16562) );
  INV_X1 U15589 ( .A(n13801), .ZN(n13802) );
  OAI21_X1 U15590 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n13800), .A(
        n13802), .ZN(n18375) );
  OAI21_X1 U15591 ( .B1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n13801), .A(
        n11062), .ZN(n18385) );
  NAND2_X1 U15592 ( .A1(n18384), .A2(n18385), .ZN(n18383) );
  NAND2_X1 U15593 ( .A1(n18562), .A2(n18383), .ZN(n18398) );
  AOI21_X1 U15594 ( .B1(n18394), .B2(n11062), .A(n13803), .ZN(n13804) );
  INV_X1 U15595 ( .A(n13804), .ZN(n18399) );
  NAND2_X1 U15596 ( .A1(n18398), .A2(n18399), .ZN(n18397) );
  NAND2_X1 U15597 ( .A1(n18562), .A2(n18397), .ZN(n18411) );
  OAI21_X1 U15598 ( .B1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n13803), .A(
        n13805), .ZN(n18412) );
  NAND2_X1 U15599 ( .A1(n18411), .A2(n18412), .ZN(n18410) );
  NAND2_X1 U15600 ( .A1(n18562), .A2(n18410), .ZN(n18423) );
  INV_X1 U15601 ( .A(n13805), .ZN(n13807) );
  INV_X1 U15602 ( .A(n13806), .ZN(n13809) );
  OAI21_X1 U15603 ( .B1(n13807), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n13809), .ZN(n18424) );
  NAND2_X1 U15604 ( .A1(n18423), .A2(n18424), .ZN(n18422) );
  NAND2_X1 U15605 ( .A1(n18562), .A2(n18422), .ZN(n18431) );
  AOI21_X1 U15606 ( .B1(n16482), .B2(n13809), .A(n13808), .ZN(n13810) );
  INV_X1 U15607 ( .A(n13810), .ZN(n18432) );
  NAND2_X1 U15608 ( .A1(n18431), .A2(n18432), .ZN(n18430) );
  NAND2_X1 U15609 ( .A1(n18562), .A2(n18430), .ZN(n18443) );
  OR2_X1 U15610 ( .A1(n13808), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n13812) );
  NAND2_X1 U15611 ( .A1(n13811), .A2(n13812), .ZN(n18444) );
  NAND2_X1 U15612 ( .A1(n18443), .A2(n18444), .ZN(n18442) );
  NAND2_X1 U15613 ( .A1(n18562), .A2(n18442), .ZN(n18452) );
  AOI21_X1 U15614 ( .B1(n16461), .B2(n13811), .A(n11000), .ZN(n16466) );
  INV_X1 U15615 ( .A(n16466), .ZN(n18453) );
  NAND2_X1 U15616 ( .A1(n18452), .A2(n18453), .ZN(n18451) );
  NAND2_X1 U15617 ( .A1(n18562), .A2(n18451), .ZN(n18461) );
  XNOR2_X1 U15618 ( .A(n11000), .B(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n18462) );
  NAND2_X1 U15619 ( .A1(n18461), .A2(n18462), .ZN(n18460) );
  NAND2_X1 U15620 ( .A1(n18562), .A2(n18460), .ZN(n18474) );
  AOI21_X1 U15621 ( .B1(n11000), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n13814) );
  OR2_X1 U15622 ( .A1(n13814), .A2(n13813), .ZN(n18475) );
  NAND2_X1 U15623 ( .A1(n18474), .A2(n18475), .ZN(n18473) );
  NAND2_X1 U15624 ( .A1(n18562), .A2(n18473), .ZN(n18483) );
  XNOR2_X1 U15625 ( .A(n13813), .B(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n18484) );
  NAND2_X1 U15626 ( .A1(n18483), .A2(n18484), .ZN(n18482) );
  NAND2_X1 U15627 ( .A1(n18562), .A2(n18482), .ZN(n18493) );
  AOI21_X1 U15628 ( .B1(n13813), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n13816) );
  OR2_X1 U15629 ( .A1(n13815), .A2(n13816), .ZN(n18494) );
  NAND2_X1 U15630 ( .A1(n18493), .A2(n18494), .ZN(n18492) );
  NAND2_X1 U15631 ( .A1(n18562), .A2(n18492), .ZN(n18504) );
  OAI21_X1 U15632 ( .B1(n13815), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n13817), .ZN(n18505) );
  NAND2_X1 U15633 ( .A1(n18504), .A2(n18505), .ZN(n18503) );
  NAND2_X1 U15634 ( .A1(n18562), .A2(n18503), .ZN(n18518) );
  INV_X1 U15635 ( .A(n13821), .ZN(n13818) );
  AOI21_X1 U15636 ( .B1(n18512), .B2(n13817), .A(n13818), .ZN(n16386) );
  INV_X1 U15637 ( .A(n16386), .ZN(n18519) );
  NAND2_X1 U15638 ( .A1(n18518), .A2(n18519), .ZN(n18517) );
  NAND2_X1 U15639 ( .A1(n18562), .A2(n18517), .ZN(n18528) );
  NAND2_X1 U15640 ( .A1(n13821), .A2(n13820), .ZN(n13822) );
  NAND2_X1 U15641 ( .A1(n13819), .A2(n13822), .ZN(n18529) );
  NAND2_X1 U15642 ( .A1(n18528), .A2(n18529), .ZN(n18527) );
  NAND2_X1 U15643 ( .A1(n18562), .A2(n18527), .ZN(n18543) );
  AOI21_X1 U15644 ( .B1(n16360), .B2(n13819), .A(n13823), .ZN(n16357) );
  INV_X1 U15645 ( .A(n16357), .ZN(n18544) );
  NAND2_X1 U15646 ( .A1(n18543), .A2(n18544), .ZN(n18542) );
  NAND2_X1 U15647 ( .A1(n18562), .A2(n18542), .ZN(n18561) );
  INV_X1 U15648 ( .A(n18561), .ZN(n13825) );
  XNOR2_X1 U15649 ( .A(n13823), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n18563) );
  INV_X1 U15650 ( .A(n18563), .ZN(n13824) );
  NAND2_X1 U15651 ( .A1(n13825), .A2(n13824), .ZN(n13827) );
  NAND2_X1 U15652 ( .A1(n18563), .A2(n18561), .ZN(n13826) );
  OR4_X1 U15653 ( .A1(n17266), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(
        P2_STATE2_REG_2__SCAN_IN), .A4(P2_STATEBS16_REG_SCAN_IN), .ZN(n18663)
         );
  INV_X2 U15654 ( .A(n18663), .ZN(n18564) );
  NAND3_X1 U15655 ( .A1(n13827), .A2(n13826), .A3(n18564), .ZN(n13867) );
  INV_X1 U15656 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14462) );
  OR2_X1 U15657 ( .A1(n10978), .A2(n14462), .ZN(n13833) );
  INV_X1 U15658 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n17338) );
  NAND2_X1 U15659 ( .A1(n14450), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13830) );
  NAND2_X1 U15660 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13829) );
  OAI211_X1 U15661 ( .C1(n17338), .C2(n14452), .A(n13830), .B(n13829), .ZN(
        n13831) );
  INV_X1 U15662 ( .A(n13831), .ZN(n13832) );
  AND2_X1 U15663 ( .A1(n13833), .A2(n13832), .ZN(n14448) );
  INV_X1 U15664 ( .A(n18683), .ZN(n18657) );
  NOR2_X1 U15665 ( .A1(n18630), .A2(n18657), .ZN(n14498) );
  INV_X1 U15666 ( .A(n18675), .ZN(n21639) );
  OR2_X1 U15667 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n21639), .ZN(n13856) );
  NOR2_X1 U15668 ( .A1(n11691), .A2(n13856), .ZN(n13834) );
  AOI22_X1 U15669 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_30__SCAN_IN), .ZN(n13838) );
  NAND2_X1 U15670 ( .A1(n12280), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n13837) );
  NAND2_X1 U15671 ( .A1(n13838), .A2(n13837), .ZN(n13840) );
  INV_X1 U15672 ( .A(n13839), .ZN(n13842) );
  INV_X1 U15673 ( .A(n13840), .ZN(n13841) );
  NAND2_X1 U15674 ( .A1(n13842), .A2(n13841), .ZN(n13843) );
  INV_X1 U15675 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n21607) );
  NAND2_X1 U15676 ( .A1(n19621), .A2(n21607), .ZN(n13844) );
  NOR2_X1 U15677 ( .A1(n18639), .A2(n13844), .ZN(n13845) );
  NAND2_X1 U15678 ( .A1(n12275), .A2(n13845), .ZN(n18654) );
  INV_X1 U15679 ( .A(n18654), .ZN(n13846) );
  NAND2_X1 U15680 ( .A1(n13848), .A2(n13847), .ZN(n14444) );
  INV_X1 U15681 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n13861) );
  NOR2_X1 U15682 ( .A1(n13849), .A2(n13861), .ZN(n13850) );
  XNOR2_X1 U15683 ( .A(n14444), .B(n13850), .ZN(n14412) );
  OAI21_X1 U15684 ( .B1(P2_STATEBS16_REG_SCAN_IN), .B2(n21639), .A(
        P2_EBX_REG_31__SCAN_IN), .ZN(n13851) );
  NOR2_X1 U15685 ( .A1(n11691), .A2(n13851), .ZN(n13852) );
  INV_X1 U15686 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n18247) );
  NAND2_X1 U15687 ( .A1(n18247), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n18676) );
  OR3_X1 U15688 ( .A1(n19233), .A2(n18676), .A3(P2_STATE2_REG_1__SCAN_IN), 
        .ZN(n18674) );
  INV_X1 U15689 ( .A(n18674), .ZN(n13854) );
  NAND2_X1 U15690 ( .A1(n18583), .A2(n18663), .ZN(n13853) );
  OAI22_X1 U15691 ( .A1(n14412), .A2(n18552), .B1(n17338), .B2(n18551), .ZN(
        n13863) );
  OR2_X1 U15692 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n18639), .ZN(n13855) );
  NAND2_X1 U15693 ( .A1(n19621), .A2(n13855), .ZN(n13858) );
  INV_X1 U15694 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n18556) );
  NAND2_X1 U15695 ( .A1(n18556), .A2(n13856), .ZN(n13857) );
  AOI21_X1 U15696 ( .B1(n13858), .B2(n13857), .A(n19686), .ZN(n13859) );
  INV_X1 U15697 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13860) );
  INV_X1 U15698 ( .A(n18537), .ZN(n18554) );
  OAI22_X1 U15699 ( .A1(n18557), .A2(n13861), .B1(n13860), .B2(n18554), .ZN(
        n13862) );
  AOI211_X1 U15700 ( .C1(n14430), .C2(n18539), .A(n13863), .B(n13862), .ZN(
        n13864) );
  INV_X1 U15701 ( .A(n13865), .ZN(n13866) );
  NAND2_X1 U15702 ( .A1(n13867), .A2(n13866), .ZN(P2_U2825) );
  AOI21_X1 U15703 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n20748), .A(
        n13868), .ZN(n13870) );
  AOI21_X1 U15704 ( .B1(n13869), .B2(n13870), .A(n21192), .ZN(n21189) );
  NAND2_X1 U15705 ( .A1(n21189), .A2(n20559), .ZN(n13878) );
  INV_X1 U15706 ( .A(n13870), .ZN(n13876) );
  NAND2_X1 U15707 ( .A1(n13872), .A2(n13871), .ZN(n13875) );
  OAI211_X1 U15708 ( .C1(n13876), .C2(n13875), .A(n13874), .B(n13873), .ZN(
        n17747) );
  OAI22_X1 U15709 ( .A1(n18796), .A2(n13878), .B1(n17747), .B2(n13877), .ZN(
        n13891) );
  XNOR2_X1 U15710 ( .A(n20559), .B(n18961), .ZN(n13879) );
  OAI21_X1 U15711 ( .B1(n13879), .B2(n20091), .A(n21659), .ZN(n21191) );
  NOR3_X1 U15712 ( .A1(n13968), .A2(n21192), .A3(n21191), .ZN(n13890) );
  INV_X1 U15713 ( .A(n13880), .ZN(n13888) );
  INV_X1 U15714 ( .A(n13881), .ZN(n13887) );
  INV_X1 U15715 ( .A(n13970), .ZN(n13969) );
  OAI211_X1 U15716 ( .C1(n20746), .C2(n18878), .A(n13969), .B(n13882), .ZN(
        n13884) );
  OAI21_X1 U15717 ( .B1(n13885), .B2(n13884), .A(n13883), .ZN(n13886) );
  OAI211_X1 U15718 ( .C1(n13889), .C2(n13888), .A(n13887), .B(n13886), .ZN(
        n16902) );
  AOI211_X1 U15719 ( .C1(n18961), .C2(n13891), .A(n13890), .B(n16902), .ZN(
        n13892) );
  INV_X1 U15720 ( .A(n21221), .ZN(n21244) );
  AOI221_X4 U15721 ( .B1(n18878), .B2(n13892), .C1(n17747), .C2(n13892), .A(
        n21244), .ZN(n21151) );
  AOI22_X1 U15722 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17688), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13896) );
  AOI22_X1 U15723 ( .A1(n17585), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17703), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n13895) );
  AOI22_X1 U15724 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17713), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13894) );
  AOI22_X1 U15725 ( .A1(n20181), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17714), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13893) );
  NAND4_X1 U15726 ( .A1(n13896), .A2(n13895), .A3(n13894), .A4(n13893), .ZN(
        n13903) );
  AOI22_X1 U15727 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13901) );
  AOI22_X1 U15728 ( .A1(n17689), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13900) );
  AOI22_X1 U15729 ( .A1(n17722), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13899) );
  AOI22_X1 U15730 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13898) );
  NAND4_X1 U15731 ( .A1(n13901), .A2(n13900), .A3(n13899), .A4(n13898), .ZN(
        n13902) );
  AOI22_X1 U15732 ( .A1(n17585), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13907) );
  AOI22_X1 U15733 ( .A1(n17719), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17722), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13906) );
  AOI22_X1 U15734 ( .A1(n20181), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17713), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13905) );
  AOI22_X1 U15735 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17714), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13904) );
  NAND4_X1 U15736 ( .A1(n13907), .A2(n13906), .A3(n13905), .A4(n13904), .ZN(
        n13913) );
  AOI22_X1 U15737 ( .A1(n17688), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13911) );
  AOI22_X1 U15738 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13910) );
  AOI22_X1 U15739 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13909) );
  AOI22_X1 U15740 ( .A1(n17689), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17703), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n13908) );
  NAND4_X1 U15741 ( .A1(n13911), .A2(n13910), .A3(n13909), .A4(n13908), .ZN(
        n13912) );
  AOI22_X1 U15742 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17720), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n10966), .ZN(n13917) );
  AOI22_X1 U15743 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n13981), .B1(
        n17722), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13916) );
  AOI22_X1 U15744 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n13934), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17713), .ZN(n13915) );
  AOI22_X1 U15745 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20181), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17714), .ZN(n13914) );
  NAND4_X1 U15746 ( .A1(n13917), .A2(n13916), .A3(n13915), .A4(n13914), .ZN(
        n13923) );
  AOI22_X1 U15747 ( .A1(n13440), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17703), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n13921) );
  AOI22_X1 U15748 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17590), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13920) );
  AOI22_X1 U15749 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n17698), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n13456), .ZN(n13919) );
  AOI22_X1 U15750 ( .A1(n13392), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13918) );
  NAND4_X1 U15751 ( .A1(n13921), .A2(n13920), .A3(n13919), .A4(n13918), .ZN(
        n13922) );
  NOR2_X2 U15752 ( .A1(n13923), .A2(n13922), .ZN(n14019) );
  AOI22_X1 U15753 ( .A1(n17585), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n13981), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13927) );
  AOI22_X1 U15754 ( .A1(n13440), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17722), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13926) );
  AOI22_X1 U15755 ( .A1(n20181), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17714), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13925) );
  AOI22_X1 U15756 ( .A1(n13934), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17713), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13924) );
  NAND4_X1 U15757 ( .A1(n13927), .A2(n13926), .A3(n13925), .A4(n13924), .ZN(
        n13933) );
  AOI22_X1 U15758 ( .A1(n13392), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n13456), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13931) );
  AOI22_X1 U15759 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13930) );
  AOI22_X1 U15760 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17703), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13929) );
  AOI22_X1 U15761 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13928) );
  NAND4_X1 U15762 ( .A1(n13931), .A2(n13930), .A3(n13929), .A4(n13928), .ZN(
        n13932) );
  AOI22_X1 U15763 ( .A1(n17688), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13944) );
  AOI22_X1 U15764 ( .A1(n17703), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n13943) );
  INV_X1 U15765 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18958) );
  AOI22_X1 U15766 ( .A1(n17713), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17714), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13935) );
  OAI21_X1 U15767 ( .B1(n13395), .B2(n18958), .A(n13935), .ZN(n13941) );
  AOI22_X1 U15768 ( .A1(n17585), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13939) );
  AOI22_X1 U15769 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17722), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13938) );
  AOI22_X1 U15770 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17689), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13937) );
  AOI22_X1 U15771 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13936) );
  NAND4_X1 U15772 ( .A1(n13939), .A2(n13938), .A3(n13937), .A4(n13936), .ZN(
        n13940) );
  AOI211_X1 U15773 ( .C1(n17554), .C2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n13941), .B(n13940), .ZN(n13942) );
  NAND3_X1 U15774 ( .A1(n13944), .A2(n13943), .A3(n13942), .ZN(n20612) );
  NAND2_X1 U15775 ( .A1(n14016), .A2(n20612), .ZN(n13976) );
  NOR2_X1 U15776 ( .A1(n20607), .A2(n13976), .ZN(n13975) );
  AOI22_X1 U15777 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13954) );
  AOI22_X1 U15778 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17722), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13953) );
  AOI22_X1 U15779 ( .A1(n17713), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17714), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13945) );
  OAI21_X1 U15780 ( .B1(n13395), .B2(n18876), .A(n13945), .ZN(n13951) );
  AOI22_X1 U15781 ( .A1(n17689), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13949) );
  AOI22_X1 U15782 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13948) );
  AOI22_X1 U15783 ( .A1(n17688), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n13947) );
  AOI22_X1 U15784 ( .A1(n17719), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17703), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13946) );
  NAND4_X1 U15785 ( .A1(n13949), .A2(n13948), .A3(n13947), .A4(n13946), .ZN(
        n13950) );
  AOI211_X1 U15786 ( .C1(n17554), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n13951), .B(n13950), .ZN(n13952) );
  NAND3_X1 U15787 ( .A1(n13954), .A2(n13953), .A3(n13952), .ZN(n20601) );
  NAND2_X1 U15788 ( .A1(n13975), .A2(n20601), .ZN(n13973) );
  AOI22_X1 U15789 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17703), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n13964) );
  AOI22_X1 U15790 ( .A1(n17688), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13963) );
  AOI22_X1 U15791 ( .A1(n17713), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17714), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13955) );
  OAI21_X1 U15792 ( .B1(n13395), .B2(n18793), .A(n13955), .ZN(n13961) );
  AOI22_X1 U15793 ( .A1(n17719), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13959) );
  AOI22_X1 U15794 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13958) );
  AOI22_X1 U15795 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17689), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13957) );
  AOI22_X1 U15796 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17722), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13956) );
  NAND4_X1 U15797 ( .A1(n13959), .A2(n13958), .A3(n13957), .A4(n13956), .ZN(
        n13960) );
  AOI211_X1 U15798 ( .C1(n17554), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n13961), .B(n13960), .ZN(n13962) );
  NAND3_X1 U15799 ( .A1(n13964), .A2(n13963), .A3(n13962), .ZN(n17754) );
  NAND2_X1 U15800 ( .A1(n13966), .A2(n13965), .ZN(n20093) );
  NAND3_X1 U15801 ( .A1(n13969), .A2(n13968), .A3(n13967), .ZN(n16899) );
  NAND2_X1 U15802 ( .A1(n13971), .A2(n20750), .ZN(n20903) );
  INV_X4 U15803 ( .A(n20903), .ZN(n21175) );
  NAND2_X1 U15804 ( .A1(n20559), .A2(n13970), .ZN(n20761) );
  NAND2_X1 U15805 ( .A1(n20762), .A2(n20761), .ZN(n20829) );
  AOI21_X2 U15806 ( .B1(n13971), .B2(n20829), .A(n20779), .ZN(n20951) );
  NOR2_X4 U15807 ( .A1(n21147), .A2(n21171), .ZN(n21051) );
  NOR2_X1 U15808 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18010), .ZN(
        n17944) );
  AOI21_X1 U15809 ( .B1(n18010), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n17944), .ZN(n17908) );
  INV_X1 U15810 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21135) );
  NAND2_X1 U15811 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n20916) );
  INV_X1 U15812 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n18009) );
  NOR2_X1 U15813 ( .A1(n20916), .A2(n18009), .ZN(n20923) );
  NAND2_X1 U15814 ( .A1(n20923), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n20937) );
  INV_X1 U15815 ( .A(n20937), .ZN(n20929) );
  NAND2_X1 U15816 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n20929), .ZN(
        n14040) );
  INV_X1 U15817 ( .A(n14040), .ZN(n20957) );
  NAND2_X1 U15818 ( .A1(n20957), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n20953) );
  INV_X1 U15819 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n20958) );
  NOR2_X1 U15820 ( .A1(n20953), .A2(n20958), .ZN(n20950) );
  INV_X1 U15821 ( .A(n20950), .ZN(n21122) );
  NAND2_X1 U15822 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17923), .ZN(
        n14004) );
  INV_X1 U15823 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n21172) );
  AOI22_X1 U15824 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17923), .B1(
        n18010), .B2(n21172), .ZN(n18045) );
  AOI21_X1 U15825 ( .B1(n20593), .B2(n13972), .A(n18010), .ZN(n14002) );
  XOR2_X1 U15826 ( .A(n20597), .B(n13973), .Z(n13974) );
  NAND2_X1 U15827 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n13974), .ZN(
        n14001) );
  XOR2_X1 U15828 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n13974), .Z(
        n18074) );
  XOR2_X1 U15829 ( .A(n20601), .B(n13975), .Z(n13997) );
  XOR2_X1 U15830 ( .A(n20607), .B(n13976), .Z(n13977) );
  NAND2_X1 U15831 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13977), .ZN(
        n13996) );
  XOR2_X1 U15832 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n13977), .Z(
        n18093) );
  INV_X1 U15833 ( .A(n13978), .ZN(n20616) );
  NOR2_X1 U15834 ( .A1(n20734), .A2(n20616), .ZN(n13979) );
  NAND2_X1 U15835 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13980), .ZN(
        n13993) );
  XOR2_X1 U15836 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n13980), .Z(
        n18121) );
  NAND2_X1 U15837 ( .A1(n14019), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13992) );
  XNOR2_X1 U15838 ( .A(n20734), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18126) );
  AOI22_X1 U15839 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13981), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n13985) );
  AOI22_X1 U15840 ( .A1(n17713), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17714), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n13984) );
  AOI22_X1 U15841 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17683), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13983) );
  AOI22_X1 U15842 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17722), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n13990) );
  AOI22_X1 U15843 ( .A1(n17719), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17703), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n13989) );
  AOI22_X1 U15844 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13456), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n13988) );
  AOI22_X1 U15845 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13987) );
  NAND4_X1 U15846 ( .A1(n13990), .A2(n13989), .A3(n13988), .A4(n13987), .ZN(
        n13991) );
  INV_X1 U15847 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20827) );
  NOR2_X1 U15848 ( .A1(n18134), .A2(n20827), .ZN(n18133) );
  NAND2_X1 U15849 ( .A1(n18126), .A2(n18133), .ZN(n18125) );
  NAND2_X1 U15850 ( .A1(n13992), .A2(n18125), .ZN(n18120) );
  NAND2_X1 U15851 ( .A1(n18121), .A2(n18120), .ZN(n18119) );
  NAND2_X1 U15852 ( .A1(n13993), .A2(n18119), .ZN(n13994) );
  NAND2_X1 U15853 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13994), .ZN(
        n13995) );
  INV_X1 U15854 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20865) );
  XNOR2_X1 U15855 ( .A(n20865), .B(n13994), .ZN(n18105) );
  XOR2_X1 U15856 ( .A(n20612), .B(n14016), .Z(n18104) );
  NAND2_X1 U15857 ( .A1(n18105), .A2(n18104), .ZN(n18103) );
  NAND2_X1 U15858 ( .A1(n13997), .A2(n13998), .ZN(n14000) );
  NAND2_X1 U15859 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18080), .ZN(
        n13999) );
  NAND2_X1 U15860 ( .A1(n18059), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n18058) );
  NAND2_X1 U15861 ( .A1(n14002), .A2(n17773), .ZN(n14003) );
  INV_X1 U15862 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18041) );
  INV_X1 U15863 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18028) );
  NAND2_X1 U15864 ( .A1(n18041), .A2(n18028), .ZN(n18025) );
  INV_X1 U15865 ( .A(n18025), .ZN(n18016) );
  NOR4_X1 U15866 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14005) );
  NAND2_X1 U15867 ( .A1(n18016), .A2(n14005), .ZN(n17776) );
  NOR2_X1 U15868 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17776), .ZN(
        n14006) );
  AOI21_X1 U15869 ( .B1(n18012), .B2(n14006), .A(n18010), .ZN(n14008) );
  INV_X1 U15870 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21121) );
  NOR2_X1 U15871 ( .A1(n14008), .A2(n14007), .ZN(n17785) );
  NAND2_X1 U15872 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17756) );
  INV_X1 U15873 ( .A(n17756), .ZN(n21109) );
  NAND2_X1 U15874 ( .A1(n21109), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17764) );
  NAND2_X1 U15875 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n20806) );
  INV_X1 U15876 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n20807) );
  NOR2_X1 U15877 ( .A1(n20806), .A2(n20807), .ZN(n14010) );
  INV_X1 U15878 ( .A(n14010), .ZN(n20972) );
  NOR2_X1 U15879 ( .A1(n17764), .A2(n20972), .ZN(n17817) );
  NAND3_X1 U15880 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17817), .ZN(n17887) );
  NOR2_X1 U15881 ( .A1(n18010), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17842) );
  INV_X1 U15882 ( .A(n17842), .ZN(n17760) );
  NOR4_X1 U15883 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A4(n17760), .ZN(n17820) );
  INV_X1 U15884 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n20974) );
  NAND2_X1 U15885 ( .A1(n17820), .A2(n20974), .ZN(n17855) );
  OAI22_X1 U15886 ( .A1(n17785), .A2(n17887), .B1(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17855), .ZN(n14009) );
  NAND2_X1 U15887 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21079) );
  NAND2_X1 U15888 ( .A1(n17840), .A2(n17761), .ZN(n17759) );
  NAND3_X1 U15889 ( .A1(n14010), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17759), .ZN(n17818) );
  NOR3_X2 U15890 ( .A1(n17880), .A2(n21079), .A3(n17818), .ZN(n17922) );
  NAND2_X1 U15891 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17904) );
  INV_X1 U15892 ( .A(n17904), .ZN(n14041) );
  INV_X1 U15893 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n20998) );
  INV_X1 U15894 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n20986) );
  AOI21_X1 U15895 ( .B1(n20998), .B2(n20986), .A(n18010), .ZN(n14011) );
  NOR2_X1 U15896 ( .A1(n18010), .A2(n17880), .ZN(n17876) );
  INV_X1 U15897 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21015) );
  NAND2_X1 U15898 ( .A1(n17915), .A2(n14051), .ZN(n17907) );
  NAND2_X1 U15899 ( .A1(n17908), .A2(n17907), .ZN(n17906) );
  NOR2_X1 U15900 ( .A1(n21122), .A2(n17764), .ZN(n20798) );
  INV_X1 U15901 ( .A(n14015), .ZN(n14013) );
  NAND2_X1 U15902 ( .A1(n14013), .A2(n20612), .ZN(n14024) );
  NOR2_X1 U15903 ( .A1(n20607), .A2(n14024), .ZN(n14014) );
  NAND2_X1 U15904 ( .A1(n14014), .A2(n20601), .ZN(n14028) );
  NOR2_X1 U15905 ( .A1(n20597), .A2(n14028), .ZN(n14031) );
  NAND2_X1 U15906 ( .A1(n14031), .A2(n17754), .ZN(n14032) );
  XOR2_X1 U15907 ( .A(n20601), .B(n14014), .Z(n14026) );
  XNOR2_X1 U15908 ( .A(n20612), .B(n14015), .ZN(n14022) );
  AOI21_X1 U15909 ( .B1(n14016), .B2(n20739), .A(n14015), .ZN(n14017) );
  INV_X1 U15910 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14039) );
  NOR2_X1 U15911 ( .A1(n14017), .A2(n14039), .ZN(n14021) );
  XOR2_X1 U15912 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n14017), .Z(
        n18118) );
  NOR2_X1 U15913 ( .A1(n14019), .A2(n20827), .ZN(n14020) );
  NAND3_X1 U15914 ( .A1(n18134), .A2(n14019), .A3(n20827), .ZN(n14018) );
  NOR2_X1 U15915 ( .A1(n18118), .A2(n18117), .ZN(n18116) );
  NOR2_X1 U15916 ( .A1(n14021), .A2(n18116), .ZN(n18108) );
  XOR2_X1 U15917 ( .A(n20865), .B(n14022), .Z(n18107) );
  INV_X1 U15918 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20866) );
  NOR2_X1 U15919 ( .A1(n14023), .A2(n20866), .ZN(n14025) );
  XNOR2_X1 U15920 ( .A(n20607), .B(n14024), .ZN(n18099) );
  INV_X1 U15921 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n20873) );
  XOR2_X1 U15922 ( .A(n20873), .B(n14026), .Z(n18083) );
  XNOR2_X1 U15923 ( .A(n20597), .B(n14028), .ZN(n14030) );
  INV_X1 U15924 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n20884) );
  XOR2_X1 U15925 ( .A(n17754), .B(n14031), .Z(n14034) );
  NOR2_X1 U15926 ( .A1(n14032), .A2(n14036), .ZN(n14038) );
  INV_X1 U15927 ( .A(n14032), .ZN(n14037) );
  NAND2_X1 U15928 ( .A1(n14034), .A2(n14033), .ZN(n18061) );
  OAI21_X1 U15929 ( .B1(n14037), .B2(n14036), .A(n18061), .ZN(n14035) );
  NOR2_X4 U15930 ( .A1(n20559), .A2(n21140), .ZN(n21183) );
  INV_X1 U15931 ( .A(n21183), .ZN(n21056) );
  NOR2_X2 U15932 ( .A1(n17754), .A2(n21190), .ZN(n21067) );
  OAI22_X1 U15933 ( .A1(n20907), .A2(n21056), .B1(n21110), .B2(n20906), .ZN(
        n20915) );
  AOI21_X1 U15934 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n21171), .A(
        n20903), .ZN(n20842) );
  INV_X1 U15935 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n20898) );
  NOR2_X1 U15936 ( .A1(n20898), .A2(n21172), .ZN(n20912) );
  NAND3_X1 U15937 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20878) );
  NAND2_X1 U15938 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20844) );
  NOR2_X1 U15939 ( .A1(n20878), .A2(n20844), .ZN(n20863) );
  AND2_X1 U15940 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n20863), .ZN(
        n21174) );
  NAND2_X1 U15941 ( .A1(n20912), .A2(n21174), .ZN(n20904) );
  INV_X1 U15942 ( .A(n20904), .ZN(n21113) );
  NAND2_X1 U15943 ( .A1(n20798), .A2(n21113), .ZN(n14042) );
  INV_X1 U15944 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20832) );
  OAI21_X1 U15945 ( .B1(n20832), .B2(n20827), .A(n14039), .ZN(n20846) );
  INV_X1 U15946 ( .A(n20846), .ZN(n20843) );
  NOR2_X1 U15947 ( .A1(n20843), .A2(n20878), .ZN(n20861) );
  NAND3_X1 U15948 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n20861), .A3(
        n20912), .ZN(n20908) );
  NOR3_X1 U15949 ( .A1(n21122), .A2(n17756), .A3(n20908), .ZN(n21120) );
  NAND2_X1 U15950 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n21120), .ZN(
        n20801) );
  OAI22_X1 U15951 ( .A1(n20842), .A2(n14042), .B1(n21119), .B2(n20801), .ZN(
        n21026) );
  AOI21_X1 U15952 ( .B1(n20798), .B2(n20915), .A(n21026), .ZN(n20973) );
  NOR2_X1 U15953 ( .A1(n20974), .A2(n20972), .ZN(n21029) );
  INV_X1 U15954 ( .A(n21029), .ZN(n14044) );
  NOR2_X1 U15955 ( .A1(n20973), .A2(n14044), .ZN(n21075) );
  INV_X1 U15956 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n21071) );
  INV_X1 U15957 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17888) );
  NOR2_X1 U15958 ( .A1(n21071), .A2(n17888), .ZN(n20999) );
  NAND2_X1 U15959 ( .A1(n14041), .A2(n20999), .ZN(n14043) );
  INV_X1 U15960 ( .A(n14043), .ZN(n21028) );
  NAND2_X1 U15961 ( .A1(n21075), .A2(n21028), .ZN(n21014) );
  OAI22_X1 U15962 ( .A1(n17923), .A2(n14047), .B1(n21014), .B2(n21015), .ZN(
        n14050) );
  INV_X1 U15963 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17905) );
  NOR2_X1 U15964 ( .A1(n17905), .A2(n21015), .ZN(n21027) );
  INV_X1 U15965 ( .A(n21027), .ZN(n17950) );
  INV_X1 U15966 ( .A(n17887), .ZN(n17903) );
  NOR2_X2 U15967 ( .A1(n20958), .A2(n20962), .ZN(n21108) );
  NAND2_X1 U15968 ( .A1(n17903), .A2(n21108), .ZN(n21068) );
  INV_X1 U15969 ( .A(n14042), .ZN(n20799) );
  NAND2_X1 U15970 ( .A1(n20799), .A2(n21029), .ZN(n20983) );
  NOR2_X1 U15971 ( .A1(n14043), .A2(n20983), .ZN(n21021) );
  NAND2_X1 U15972 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n21021), .ZN(
        n14045) );
  NAND2_X1 U15973 ( .A1(n21176), .A2(n21080), .ZN(n21074) );
  OAI21_X1 U15974 ( .B1(n20801), .B2(n14044), .A(n21184), .ZN(n21073) );
  OAI21_X1 U15975 ( .B1(n21028), .B2(n21119), .A(n21073), .ZN(n21008) );
  AOI221_X1 U15976 ( .B1(n20827), .B2(n21171), .C1(n14045), .C2(n21171), .A(
        n21008), .ZN(n21038) );
  OAI21_X1 U15977 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n21119), .A(
        n21038), .ZN(n21024) );
  AOI211_X1 U15978 ( .C1(n20903), .C2(n14045), .A(n21062), .B(n21024), .ZN(
        n14048) );
  INV_X1 U15979 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n20938) );
  NAND2_X1 U15980 ( .A1(n21111), .A2(n20957), .ZN(n17994) );
  NAND2_X1 U15981 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n20959), .ZN(
        n20964) );
  NAND2_X1 U15982 ( .A1(n17903), .A2(n17816), .ZN(n21066) );
  INV_X1 U15983 ( .A(n21066), .ZN(n17866) );
  NAND2_X1 U15984 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17866), .ZN(
        n17875) );
  NOR2_X1 U15985 ( .A1(n17904), .A2(n17875), .ZN(n17952) );
  INV_X1 U15986 ( .A(n17952), .ZN(n21009) );
  NOR2_X1 U15987 ( .A1(n17950), .A2(n21009), .ZN(n17963) );
  INV_X1 U15988 ( .A(n17963), .ZN(n21032) );
  NAND3_X1 U15989 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n18010), .A3(
        n14046), .ZN(n17964) );
  OAI221_X1 U15990 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n21151), 
        .C1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n14050), .A(n14049), .ZN(
        n14054) );
  INV_X1 U15991 ( .A(n21176), .ZN(n21137) );
  NAND2_X1 U15992 ( .A1(n18669), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n18652) );
  NAND2_X1 U15993 ( .A1(n10971), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n14056) );
  NAND2_X1 U15994 ( .A1(n14056), .A2(n19233), .ZN(n14078) );
  NAND2_X1 U15995 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19291) );
  INV_X1 U15996 ( .A(n19291), .ZN(n14057) );
  AND2_X1 U15997 ( .A1(n14057), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14058) );
  NAND2_X1 U15998 ( .A1(n14058), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n15345) );
  INV_X1 U15999 ( .A(n14058), .ZN(n14068) );
  NAND2_X1 U16000 ( .A1(n14068), .A2(n19213), .ZN(n14059) );
  AND3_X1 U16001 ( .A1(n15345), .A2(n19292), .A3(n14059), .ZN(n19205) );
  AOI21_X1 U16002 ( .B1(n14078), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19205), .ZN(n14060) );
  NOR2_X1 U16003 ( .A1(n10971), .A2(n18669), .ZN(n14648) );
  NAND2_X1 U16004 ( .A1(n14064), .A2(n14063), .ZN(n14065) );
  NAND2_X1 U16005 ( .A1(n14066), .A2(n14062), .ZN(n14071) );
  NAND2_X1 U16006 ( .A1(n19291), .A2(n19221), .ZN(n14067) );
  NAND2_X1 U16007 ( .A1(n14068), .A2(n14067), .ZN(n19206) );
  NOR2_X1 U16008 ( .A1(n19206), .A2(n19326), .ZN(n14069) );
  AOI21_X1 U16009 ( .B1(n14078), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n14069), .ZN(n14070) );
  NAND2_X1 U16010 ( .A1(n14071), .A2(n14070), .ZN(n14073) );
  NAND2_X1 U16011 ( .A1(n14073), .A2(n14072), .ZN(n14084) );
  OR2_X1 U16012 ( .A1(n14073), .A2(n14072), .ZN(n14074) );
  NAND2_X1 U16013 ( .A1(n14078), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n14076) );
  NAND2_X1 U16014 ( .A1(n19294), .A2(n19263), .ZN(n14075) );
  AND2_X1 U16015 ( .A1(n14075), .A2(n19291), .ZN(n19270) );
  NAND2_X1 U16016 ( .A1(n19270), .A2(n19292), .ZN(n19318) );
  NAND2_X1 U16017 ( .A1(n14076), .A2(n19318), .ZN(n14077) );
  AOI22_X1 U16018 ( .A1(n14078), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19292), .B2(n19263), .ZN(n14079) );
  INV_X1 U16019 ( .A(n14081), .ZN(n14082) );
  NOR2_X1 U16020 ( .A1(n15181), .A2(n14082), .ZN(n14083) );
  NAND2_X1 U16021 ( .A1(n14770), .A2(n14768), .ZN(n14085) );
  NAND2_X1 U16022 ( .A1(n14085), .A2(n14084), .ZN(n14759) );
  NAND2_X1 U16023 ( .A1(n10971), .A2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n14086) );
  INV_X1 U16024 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15356) );
  NAND2_X1 U16025 ( .A1(n14995), .A2(n14994), .ZN(n14993) );
  AOI22_X1 U16026 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11481), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n14092) );
  AOI22_X1 U16027 ( .A1(n14231), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14230), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14091) );
  AOI22_X1 U16028 ( .A1(n16892), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14232), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n14090) );
  NAND2_X1 U16029 ( .A1(n14233), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n14089) );
  AND4_X1 U16030 ( .A1(n14092), .A2(n14091), .A3(n14090), .A4(n14089), .ZN(
        n14103) );
  AOI22_X1 U16031 ( .A1(n14223), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n14222), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n14096) );
  NAND2_X1 U16032 ( .A1(n14172), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14095) );
  AOI22_X1 U16033 ( .A1(n14224), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14225), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14094) );
  NAND2_X1 U16034 ( .A1(n11480), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n14093) );
  NAND4_X1 U16035 ( .A1(n14096), .A2(n14095), .A3(n14094), .A4(n14093), .ZN(
        n14101) );
  INV_X1 U16036 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14099) );
  NAND2_X1 U16037 ( .A1(n14215), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n14098) );
  NAND2_X1 U16038 ( .A1(n14216), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n14097) );
  OAI211_X1 U16039 ( .C1(n14099), .C2(n14219), .A(n14098), .B(n14097), .ZN(
        n14100) );
  NOR2_X1 U16040 ( .A1(n14101), .A2(n14100), .ZN(n14102) );
  NAND2_X1 U16041 ( .A1(n14103), .A2(n14102), .ZN(n16263) );
  AOI22_X1 U16042 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11481), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n14107) );
  AOI22_X1 U16043 ( .A1(n14231), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14230), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14106) );
  AOI22_X1 U16044 ( .A1(n16892), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n14232), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14105) );
  NAND2_X1 U16045 ( .A1(n14233), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n14104) );
  AND4_X1 U16046 ( .A1(n14107), .A2(n14106), .A3(n14105), .A4(n14104), .ZN(
        n14118) );
  AOI22_X1 U16047 ( .A1(n14223), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14222), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n14111) );
  NAND2_X1 U16048 ( .A1(n14172), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14110) );
  AOI22_X1 U16049 ( .A1(n14224), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14225), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14109) );
  NAND2_X1 U16050 ( .A1(n11480), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n14108) );
  NAND4_X1 U16051 ( .A1(n14111), .A2(n14110), .A3(n14109), .A4(n14108), .ZN(
        n14116) );
  INV_X1 U16052 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14114) );
  NAND2_X1 U16053 ( .A1(n14215), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n14113) );
  NAND2_X1 U16054 ( .A1(n14216), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n14112) );
  OAI211_X1 U16055 ( .C1(n14114), .C2(n14219), .A(n14113), .B(n14112), .ZN(
        n14115) );
  NOR2_X1 U16056 ( .A1(n14116), .A2(n14115), .ZN(n14117) );
  NAND2_X1 U16057 ( .A1(n14118), .A2(n14117), .ZN(n15495) );
  INV_X1 U16058 ( .A(n15495), .ZN(n14120) );
  INV_X1 U16059 ( .A(n15417), .ZN(n14119) );
  OR2_X1 U16060 ( .A1(n14119), .A2(n15410), .ZN(n15415) );
  OR2_X1 U16061 ( .A1(n14120), .A2(n15415), .ZN(n15493) );
  AOI22_X1 U16062 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11481), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n14124) );
  AOI22_X1 U16063 ( .A1(n14231), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14230), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14123) );
  AOI22_X1 U16064 ( .A1(n16892), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n14232), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n14122) );
  NAND2_X1 U16065 ( .A1(n14233), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n14121) );
  AND4_X1 U16066 ( .A1(n14124), .A2(n14123), .A3(n14122), .A4(n14121), .ZN(
        n14135) );
  AOI22_X1 U16067 ( .A1(n14223), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14222), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n14128) );
  NAND2_X1 U16068 ( .A1(n14172), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n14127) );
  AOI22_X1 U16069 ( .A1(n14224), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14225), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14126) );
  NAND2_X1 U16070 ( .A1(n11480), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n14125) );
  NAND4_X1 U16071 ( .A1(n14128), .A2(n14127), .A3(n14126), .A4(n14125), .ZN(
        n14133) );
  INV_X1 U16072 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14131) );
  NAND2_X1 U16073 ( .A1(n14215), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n14130) );
  NAND2_X1 U16074 ( .A1(n14216), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n14129) );
  OAI211_X1 U16075 ( .C1(n14131), .C2(n14219), .A(n14130), .B(n14129), .ZN(
        n14132) );
  NOR2_X1 U16076 ( .A1(n14133), .A2(n14132), .ZN(n14134) );
  NAND2_X1 U16077 ( .A1(n14135), .A2(n14134), .ZN(n16272) );
  INV_X1 U16078 ( .A(n16272), .ZN(n14136) );
  NOR2_X1 U16079 ( .A1(n15493), .A2(n14136), .ZN(n16261) );
  AND2_X1 U16080 ( .A1(n16263), .A2(n16261), .ZN(n14137) );
  AND2_X1 U16081 ( .A1(n15339), .A2(n15301), .ZN(n15338) );
  AOI22_X1 U16082 ( .A1(n14172), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11480), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14146) );
  INV_X1 U16083 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14141) );
  NAND2_X1 U16084 ( .A1(n14215), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n14140) );
  NAND2_X1 U16085 ( .A1(n14216), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n14139) );
  OAI211_X1 U16086 ( .C1(n14141), .C2(n14219), .A(n14140), .B(n14139), .ZN(
        n14142) );
  INV_X1 U16087 ( .A(n14142), .ZN(n14145) );
  AOI22_X1 U16088 ( .A1(n14223), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n14222), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n14144) );
  AOI22_X1 U16089 ( .A1(n14224), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14225), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14143) );
  NAND4_X1 U16090 ( .A1(n14146), .A2(n14145), .A3(n14144), .A4(n14143), .ZN(
        n14152) );
  AOI22_X1 U16091 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11481), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n14150) );
  AOI22_X1 U16092 ( .A1(n14231), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14230), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14149) );
  AOI22_X1 U16093 ( .A1(n16892), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14232), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14148) );
  NAND2_X1 U16094 ( .A1(n14233), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n14147) );
  NAND4_X1 U16095 ( .A1(n14150), .A2(n14149), .A3(n14148), .A4(n14147), .ZN(
        n14151) );
  NOR2_X1 U16096 ( .A1(n14152), .A2(n14151), .ZN(n15506) );
  AOI22_X1 U16097 ( .A1(n14172), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11480), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14160) );
  INV_X1 U16098 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14155) );
  NAND2_X1 U16099 ( .A1(n14215), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n14154) );
  NAND2_X1 U16100 ( .A1(n14216), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n14153) );
  OAI211_X1 U16101 ( .C1(n14155), .C2(n14219), .A(n14154), .B(n14153), .ZN(
        n14156) );
  INV_X1 U16102 ( .A(n14156), .ZN(n14159) );
  AOI22_X1 U16103 ( .A1(n14223), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14222), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n14158) );
  AOI22_X1 U16104 ( .A1(n14224), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14225), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14157) );
  NAND4_X1 U16105 ( .A1(n14160), .A2(n14159), .A3(n14158), .A4(n14157), .ZN(
        n14166) );
  AOI22_X1 U16106 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11481), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14164) );
  AOI22_X1 U16107 ( .A1(n14231), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14230), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14163) );
  AOI22_X1 U16108 ( .A1(n16892), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n14232), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14162) );
  NAND2_X1 U16109 ( .A1(n14233), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n14161) );
  NAND4_X1 U16110 ( .A1(n14164), .A2(n14163), .A3(n14162), .A4(n14161), .ZN(
        n14165) );
  NOR2_X1 U16111 ( .A1(n14166), .A2(n14165), .ZN(n15557) );
  INV_X1 U16112 ( .A(n15557), .ZN(n14167) );
  AOI22_X1 U16113 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11481), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14171) );
  AOI22_X1 U16114 ( .A1(n14231), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n14230), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14170) );
  AOI22_X1 U16115 ( .A1(n16892), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14232), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14169) );
  NAND2_X1 U16116 ( .A1(n14233), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n14168) );
  NAND4_X1 U16117 ( .A1(n14171), .A2(n14170), .A3(n14169), .A4(n14168), .ZN(
        n14183) );
  INV_X1 U16118 ( .A(n14172), .ZN(n14175) );
  INV_X1 U16119 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14173) );
  OAI22_X1 U16120 ( .A1(n14175), .A2(n14932), .B1(n14174), .B2(n14173), .ZN(
        n14182) );
  AOI22_X1 U16121 ( .A1(n14184), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n14215), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14176) );
  OAI21_X1 U16122 ( .B1(n14187), .B2(n14177), .A(n14176), .ZN(n14181) );
  AOI22_X1 U16123 ( .A1(n14223), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14222), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n14179) );
  AOI22_X1 U16124 ( .A1(n14224), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14225), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14178) );
  NAND2_X1 U16125 ( .A1(n14179), .A2(n14178), .ZN(n14180) );
  OR4_X1 U16126 ( .A1(n14183), .A2(n14182), .A3(n14181), .A4(n14180), .ZN(
        n15549) );
  AOI22_X1 U16127 ( .A1(n14184), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14215), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14185) );
  OAI21_X1 U16128 ( .B1(n14187), .B2(n14186), .A(n14185), .ZN(n14197) );
  AOI22_X1 U16129 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11481), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n14191) );
  AOI22_X1 U16130 ( .A1(n14231), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n14230), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n14190) );
  AOI22_X1 U16131 ( .A1(n16892), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14232), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n14189) );
  NAND2_X1 U16132 ( .A1(n14233), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n14188) );
  NAND4_X1 U16133 ( .A1(n14191), .A2(n14190), .A3(n14189), .A4(n14188), .ZN(
        n14196) );
  AOI22_X1 U16134 ( .A1(n14172), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11480), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14194) );
  AOI22_X1 U16135 ( .A1(n14223), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14222), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n14193) );
  AOI22_X1 U16136 ( .A1(n14224), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14225), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14192) );
  NAND3_X1 U16137 ( .A1(n14194), .A2(n14193), .A3(n14192), .ZN(n14195) );
  NOR3_X1 U16138 ( .A1(n14197), .A2(n14196), .A3(n14195), .ZN(n16251) );
  AOI22_X1 U16139 ( .A1(n10974), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14206) );
  AND2_X1 U16140 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n14199) );
  OR2_X1 U16141 ( .A1(n14199), .A2(n14198), .ZN(n14369) );
  INV_X1 U16142 ( .A(n14369), .ZN(n14346) );
  NAND2_X1 U16143 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n14202) );
  NAND2_X1 U16144 ( .A1(n14351), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n14201) );
  AND3_X1 U16145 ( .A1(n14346), .A2(n14202), .A3(n14201), .ZN(n14205) );
  AOI22_X1 U16146 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n14370), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14204) );
  AOI22_X1 U16147 ( .A1(n14364), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n14372), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14203) );
  NAND4_X1 U16148 ( .A1(n14206), .A2(n14205), .A3(n14204), .A4(n14203), .ZN(
        n14214) );
  AOI22_X1 U16149 ( .A1(n10975), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14212) );
  AOI22_X1 U16150 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n14370), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n14211) );
  NAND2_X1 U16151 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n14208) );
  NAND2_X1 U16152 ( .A1(n14351), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n14207) );
  AND3_X1 U16153 ( .A1(n14208), .A2(n14369), .A3(n14207), .ZN(n14210) );
  AOI22_X1 U16154 ( .A1(n14364), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14372), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n14209) );
  NAND4_X1 U16155 ( .A1(n14212), .A2(n14211), .A3(n14210), .A4(n14209), .ZN(
        n14213) );
  NAND2_X1 U16156 ( .A1(n14214), .A2(n14213), .ZN(n14241) );
  AOI22_X1 U16157 ( .A1(n14172), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11480), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14229) );
  INV_X1 U16158 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14220) );
  NAND2_X1 U16159 ( .A1(n14215), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n14218) );
  NAND2_X1 U16160 ( .A1(n14216), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n14217) );
  OAI211_X1 U16161 ( .C1(n14220), .C2(n14219), .A(n14218), .B(n14217), .ZN(
        n14221) );
  INV_X1 U16162 ( .A(n14221), .ZN(n14228) );
  AOI22_X1 U16163 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n14223), .B1(
        n14222), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14227) );
  AOI22_X1 U16164 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n14225), .B1(
        n14224), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n14226) );
  NAND4_X1 U16165 ( .A1(n14229), .A2(n14228), .A3(n14227), .A4(n14226), .ZN(
        n14239) );
  AOI22_X1 U16166 ( .A1(n11460), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11481), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14237) );
  AOI22_X1 U16167 ( .A1(n14231), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n14230), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14236) );
  AOI22_X1 U16168 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n14232), .B1(
        n16892), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14235) );
  NAND2_X1 U16169 ( .A1(n14233), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n14234) );
  NAND4_X1 U16170 ( .A1(n14237), .A2(n14236), .A3(n14235), .A4(n14234), .ZN(
        n14238) );
  NOR2_X1 U16171 ( .A1(n14239), .A2(n14238), .ZN(n14240) );
  XOR2_X1 U16172 ( .A(n14241), .B(n14240), .Z(n16243) );
  INV_X1 U16173 ( .A(n14240), .ZN(n14243) );
  INV_X1 U16174 ( .A(n14241), .ZN(n14242) );
  AND2_X1 U16175 ( .A1(n14243), .A2(n14242), .ZN(n14259) );
  AOI22_X1 U16176 ( .A1(n10974), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n14249) );
  NAND2_X1 U16177 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n14245) );
  NAND2_X1 U16178 ( .A1(n14351), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n14244) );
  AND3_X1 U16179 ( .A1(n14346), .A2(n14245), .A3(n14244), .ZN(n14248) );
  AOI22_X1 U16180 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14370), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14247) );
  AOI22_X1 U16181 ( .A1(n14364), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n14372), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n14246) );
  NAND4_X1 U16182 ( .A1(n14249), .A2(n14248), .A3(n14247), .A4(n14246), .ZN(
        n14257) );
  AOI22_X1 U16183 ( .A1(n10975), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n14255) );
  AOI22_X1 U16184 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n14370), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n14254) );
  NAND2_X1 U16185 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n14251) );
  NAND2_X1 U16186 ( .A1(n14351), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n14250) );
  AND3_X1 U16187 ( .A1(n14251), .A2(n14369), .A3(n14250), .ZN(n14253) );
  AOI22_X1 U16188 ( .A1(n14364), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n14372), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n14252) );
  NAND4_X1 U16189 ( .A1(n14255), .A2(n14254), .A3(n14253), .A4(n14252), .ZN(
        n14256) );
  NAND2_X1 U16190 ( .A1(n14257), .A2(n14256), .ZN(n14260) );
  INV_X1 U16191 ( .A(n14260), .ZN(n14258) );
  NAND2_X1 U16192 ( .A1(n14259), .A2(n14258), .ZN(n14277) );
  INV_X1 U16193 ( .A(n14259), .ZN(n14261) );
  OAI21_X1 U16194 ( .B1(n14320), .B2(n14261), .A(n14260), .ZN(n14262) );
  OAI21_X1 U16195 ( .B1(n19621), .B2(n14277), .A(n14262), .ZN(n16239) );
  AOI22_X1 U16196 ( .A1(n10974), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14268) );
  NAND2_X1 U16197 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n14264) );
  NAND2_X1 U16198 ( .A1(n14351), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n14263) );
  AND3_X1 U16199 ( .A1(n14346), .A2(n14264), .A3(n14263), .ZN(n14267) );
  AOI22_X1 U16200 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14370), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14266) );
  AOI22_X1 U16201 ( .A1(n14364), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n14372), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n14265) );
  NAND4_X1 U16202 ( .A1(n14268), .A2(n14267), .A3(n14266), .A4(n14265), .ZN(
        n14276) );
  AOI22_X1 U16203 ( .A1(n10975), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14274) );
  AOI22_X1 U16204 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n14370), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n14273) );
  NAND2_X1 U16205 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n14270) );
  NAND2_X1 U16206 ( .A1(n14351), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n14269) );
  AND3_X1 U16207 ( .A1(n14270), .A2(n14369), .A3(n14269), .ZN(n14272) );
  AOI22_X1 U16208 ( .A1(n14364), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n14372), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n14271) );
  NAND4_X1 U16209 ( .A1(n14274), .A2(n14273), .A3(n14272), .A4(n14271), .ZN(
        n14275) );
  NAND2_X1 U16210 ( .A1(n14276), .A2(n14275), .ZN(n14278) );
  NOR2_X1 U16211 ( .A1(n14277), .A2(n14278), .ZN(n14319) );
  AOI211_X1 U16212 ( .C1(n14278), .C2(n14277), .A(n14320), .B(n14319), .ZN(
        n14281) );
  XNOR2_X1 U16213 ( .A(n14280), .B(n14281), .ZN(n16234) );
  INV_X1 U16214 ( .A(n14278), .ZN(n14279) );
  NAND2_X1 U16215 ( .A1(n19621), .A2(n14279), .ZN(n16233) );
  NOR2_X1 U16216 ( .A1(n16234), .A2(n16233), .ZN(n16232) );
  INV_X1 U16217 ( .A(n14319), .ZN(n14297) );
  AOI22_X1 U16218 ( .A1(n10974), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14288) );
  NAND2_X1 U16219 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n14284) );
  NAND2_X1 U16220 ( .A1(n14351), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n14283) );
  AND3_X1 U16221 ( .A1(n14346), .A2(n14284), .A3(n14283), .ZN(n14287) );
  AOI22_X1 U16222 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n14370), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14286) );
  AOI22_X1 U16223 ( .A1(n14364), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n14372), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14285) );
  NAND4_X1 U16224 ( .A1(n14288), .A2(n14287), .A3(n14286), .A4(n14285), .ZN(
        n14296) );
  AOI22_X1 U16225 ( .A1(n10975), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n14294) );
  AOI22_X1 U16226 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n14370), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n14293) );
  NAND2_X1 U16227 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n14290) );
  NAND2_X1 U16228 ( .A1(n14351), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n14289) );
  AND3_X1 U16229 ( .A1(n14290), .A2(n14369), .A3(n14289), .ZN(n14292) );
  AOI22_X1 U16230 ( .A1(n14364), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n14372), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n14291) );
  NAND4_X1 U16231 ( .A1(n14294), .A2(n14293), .A3(n14292), .A4(n14291), .ZN(
        n14295) );
  AND2_X1 U16232 ( .A1(n14296), .A2(n14295), .ZN(n14318) );
  XNOR2_X1 U16233 ( .A(n14297), .B(n14318), .ZN(n14299) );
  NAND2_X1 U16234 ( .A1(n14299), .A2(n14298), .ZN(n14302) );
  INV_X1 U16235 ( .A(n14302), .ZN(n14300) );
  XNOR2_X1 U16236 ( .A(n14303), .B(n14300), .ZN(n16223) );
  INV_X1 U16237 ( .A(n14318), .ZN(n14301) );
  NOR2_X1 U16238 ( .A1(n11774), .A2(n14301), .ZN(n16222) );
  OAI21_X1 U16239 ( .B1(n14303), .B2(n14302), .A(n16221), .ZN(n14339) );
  AOI22_X1 U16240 ( .A1(n10974), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14309) );
  NAND2_X1 U16241 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n14305) );
  NAND2_X1 U16242 ( .A1(n14351), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n14304) );
  AND3_X1 U16243 ( .A1(n14346), .A2(n14305), .A3(n14304), .ZN(n14308) );
  AOI22_X1 U16244 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n14370), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n14307) );
  AOI22_X1 U16245 ( .A1(n14373), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n14372), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n14306) );
  NAND4_X1 U16246 ( .A1(n14309), .A2(n14308), .A3(n14307), .A4(n14306), .ZN(
        n14317) );
  AOI22_X1 U16247 ( .A1(n10975), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n14315) );
  AOI22_X1 U16248 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n14370), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n14314) );
  NAND2_X1 U16249 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n14311) );
  NAND2_X1 U16250 ( .A1(n14351), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n14310) );
  AND3_X1 U16251 ( .A1(n14311), .A2(n14369), .A3(n14310), .ZN(n14313) );
  AOI22_X1 U16252 ( .A1(n14364), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14372), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14312) );
  NAND4_X1 U16253 ( .A1(n14315), .A2(n14314), .A3(n14313), .A4(n14312), .ZN(
        n14316) );
  NAND2_X1 U16254 ( .A1(n14317), .A2(n14316), .ZN(n14322) );
  NAND2_X1 U16255 ( .A1(n14319), .A2(n14318), .ZN(n14321) );
  NOR2_X1 U16256 ( .A1(n14321), .A2(n14322), .ZN(n16203) );
  AOI211_X1 U16257 ( .C1(n14322), .C2(n14321), .A(n14320), .B(n16203), .ZN(
        n14338) );
  INV_X1 U16258 ( .A(n14322), .ZN(n14323) );
  NAND2_X1 U16259 ( .A1(n19621), .A2(n14323), .ZN(n16215) );
  INV_X1 U16260 ( .A(n16215), .ZN(n14341) );
  AOI22_X1 U16261 ( .A1(n14364), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n14372), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n14326) );
  NAND2_X1 U16262 ( .A1(n14351), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n14325) );
  NAND2_X1 U16263 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n14324) );
  NAND4_X1 U16264 ( .A1(n14326), .A2(n14369), .A3(n14325), .A4(n14324), .ZN(
        n14337) );
  AOI22_X1 U16265 ( .A1(n10974), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n14328) );
  AOI22_X1 U16266 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n14370), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n14327) );
  NAND2_X1 U16267 ( .A1(n14328), .A2(n14327), .ZN(n14336) );
  NOR2_X1 U16268 ( .A1(n11419), .A2(n14329), .ZN(n14330) );
  AOI211_X1 U16269 ( .C1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .C2(n14351), .A(
        n14369), .B(n14330), .ZN(n14334) );
  AOI22_X1 U16270 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n14370), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14333) );
  AOI22_X1 U16271 ( .A1(n10975), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14332) );
  AOI22_X1 U16272 ( .A1(n14364), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n14372), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14331) );
  NAND4_X1 U16273 ( .A1(n14334), .A2(n14333), .A3(n14332), .A4(n14331), .ZN(
        n14335) );
  OAI21_X1 U16274 ( .B1(n14337), .B2(n14336), .A(n14335), .ZN(n16204) );
  OAI211_X1 U16275 ( .C1(n11026), .C2(n14341), .A(n14340), .B(n16212), .ZN(
        n14342) );
  INV_X1 U16276 ( .A(n14342), .ZN(n16200) );
  INV_X1 U16277 ( .A(n16203), .ZN(n14343) );
  NOR3_X1 U16278 ( .A1(n14343), .A2(n19621), .A3(n16204), .ZN(n16197) );
  AOI22_X1 U16279 ( .A1(n10974), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n14350) );
  NAND2_X1 U16280 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n14345) );
  NAND2_X1 U16281 ( .A1(n14351), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n14344) );
  AND3_X1 U16282 ( .A1(n14346), .A2(n14345), .A3(n14344), .ZN(n14349) );
  AOI22_X1 U16283 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14370), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n14348) );
  AOI22_X1 U16284 ( .A1(n14364), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n14372), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n14347) );
  NAND4_X1 U16285 ( .A1(n14350), .A2(n14349), .A3(n14348), .A4(n14347), .ZN(
        n14359) );
  AOI22_X1 U16286 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n14357) );
  NAND2_X1 U16287 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n14353) );
  NAND2_X1 U16288 ( .A1(n14351), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n14352) );
  AND3_X1 U16289 ( .A1(n14353), .A2(n14369), .A3(n14352), .ZN(n14356) );
  AOI22_X1 U16290 ( .A1(n14364), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14370), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n14355) );
  AOI22_X1 U16291 ( .A1(n10975), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14372), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n14354) );
  NAND4_X1 U16292 ( .A1(n14357), .A2(n14356), .A3(n14355), .A4(n14354), .ZN(
        n14358) );
  AND2_X1 U16293 ( .A1(n14359), .A2(n14358), .ZN(n16198) );
  OAI21_X1 U16294 ( .B1(n16200), .B2(n16197), .A(n16198), .ZN(n14382) );
  AOI22_X1 U16295 ( .A1(n11645), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14372), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14363) );
  NAND2_X1 U16296 ( .A1(n11652), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n14362) );
  NAND2_X1 U16297 ( .A1(n14360), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n14361) );
  NAND4_X1 U16298 ( .A1(n14363), .A2(n14362), .A3(n14361), .A4(n14369), .ZN(
        n14380) );
  AOI22_X1 U16299 ( .A1(n14364), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10974), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14366) );
  AOI22_X1 U16300 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n14370), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14365) );
  NAND2_X1 U16301 ( .A1(n14366), .A2(n14365), .ZN(n14379) );
  INV_X1 U16302 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n19241) );
  NOR2_X1 U16303 ( .A1(n14367), .A2(n19241), .ZN(n14368) );
  AOI211_X1 U16304 ( .C1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .C2(n11652), .A(
        n14369), .B(n14368), .ZN(n14377) );
  AOI22_X1 U16305 ( .A1(n14371), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14370), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14376) );
  AOI22_X1 U16306 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n11645), .B1(
        n10975), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14375) );
  AOI22_X1 U16307 ( .A1(n14373), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n14372), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n14374) );
  NAND4_X1 U16308 ( .A1(n14377), .A2(n14376), .A3(n14375), .A4(n14374), .ZN(
        n14378) );
  OAI21_X1 U16309 ( .B1(n14380), .B2(n14379), .A(n14378), .ZN(n14381) );
  XNOR2_X1 U16310 ( .A(n14382), .B(n14381), .ZN(n15607) );
  NAND2_X1 U16311 ( .A1(n12251), .A2(n18675), .ZN(n18638) );
  NOR2_X1 U16312 ( .A1(n18638), .A2(n18630), .ZN(n14383) );
  AND2_X1 U16313 ( .A1(n18641), .A2(n14383), .ZN(n14384) );
  AOI21_X1 U16314 ( .B1(n18626), .B2(n18636), .A(n14384), .ZN(n14635) );
  NAND2_X1 U16315 ( .A1(n14635), .A2(n14385), .ZN(n14386) );
  AOI22_X1 U16316 ( .A1(n14430), .A2(n19612), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n19670), .ZN(n14407) );
  NAND2_X1 U16317 ( .A1(n19508), .A2(n14388), .ZN(n16352) );
  NOR4_X1 U16318 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_12__SCAN_IN), .A4(
        P2_ADDRESS_REG_11__SCAN_IN), .ZN(n14392) );
  NOR4_X1 U16319 ( .A1(P2_ADDRESS_REG_18__SCAN_IN), .A2(
        P2_ADDRESS_REG_17__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n14391) );
  NOR4_X1 U16320 ( .A1(P2_ADDRESS_REG_6__SCAN_IN), .A2(
        P2_ADDRESS_REG_5__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n14390) );
  NOR4_X1 U16321 ( .A1(P2_ADDRESS_REG_10__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n14389) );
  NAND4_X1 U16322 ( .A1(n14392), .A2(n14391), .A3(n14390), .A4(n14389), .ZN(
        n14397) );
  NOR4_X1 U16323 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_1__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n14395) );
  NOR4_X1 U16324 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_20__SCAN_IN), .A4(
        P2_ADDRESS_REG_19__SCAN_IN), .ZN(n14394) );
  NOR4_X1 U16325 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n14393) );
  INV_X1 U16326 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n17327) );
  NAND4_X1 U16327 ( .A1(n14395), .A2(n14394), .A3(n14393), .A4(n17327), .ZN(
        n14396) );
  OAI21_X1 U16328 ( .B1(n14397), .B2(n14396), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n14398) );
  NAND2_X1 U16329 ( .A1(n15195), .A2(BUF2_REG_14__SCAN_IN), .ZN(n14401) );
  INV_X1 U16330 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n14399) );
  OR2_X1 U16331 ( .A1(n15195), .A2(n14399), .ZN(n14400) );
  NAND2_X1 U16332 ( .A1(n14401), .A2(n14400), .ZN(n19158) );
  INV_X1 U16333 ( .A(n19158), .ZN(n14402) );
  AND2_X1 U16334 ( .A1(n10971), .A2(n15200), .ZN(n14403) );
  AOI22_X1 U16335 ( .A1(n19673), .A2(BUF1_REG_30__SCAN_IN), .B1(n19674), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n14404) );
  INV_X1 U16336 ( .A(n14404), .ZN(n14405) );
  NOR2_X1 U16337 ( .A1(n11371), .A2(n14405), .ZN(n14406) );
  OAI21_X1 U16338 ( .B1(n15607), .B2(n19677), .A(n14408), .ZN(P2_U2889) );
  NOR3_X1 U16339 ( .A1(n14412), .A2(n14411), .A3(n14462), .ZN(n14440) );
  OR2_X1 U16340 ( .A1(n14412), .A2(n14411), .ZN(n14413) );
  NAND2_X1 U16341 ( .A1(n14413), .A2(n14462), .ZN(n14442) );
  INV_X1 U16342 ( .A(n14442), .ZN(n14414) );
  NOR2_X1 U16343 ( .A1(n14440), .A2(n14414), .ZN(n14415) );
  XNOR2_X1 U16344 ( .A(n14416), .B(n14415), .ZN(n14436) );
  NAND2_X1 U16345 ( .A1(n11700), .A2(n18627), .ZN(n14417) );
  AOI21_X1 U16346 ( .B1(n14418), .B2(n14417), .A(n12052), .ZN(n18645) );
  NAND2_X1 U16347 ( .A1(n18686), .A2(n11774), .ZN(n17228) );
  NAND2_X1 U16348 ( .A1(n14436), .A2(n17258), .ZN(n14428) );
  XNOR2_X1 U16349 ( .A(n14467), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14437) );
  NAND2_X1 U16350 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_2__SCAN_IN), .ZN(n15190) );
  INV_X1 U16351 ( .A(n15190), .ZN(n17262) );
  NOR2_X1 U16352 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n17262), .ZN(n18250) );
  AND2_X1 U16353 ( .A1(n18250), .A2(n18669), .ZN(n14419) );
  AND2_X1 U16354 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n14420) );
  NOR2_X1 U16355 ( .A1(n18583), .A2(n17338), .ZN(n14429) );
  NAND2_X1 U16356 ( .A1(n21607), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n14421) );
  NAND2_X1 U16357 ( .A1(n18652), .A2(n14421), .ZN(n14553) );
  NOR2_X1 U16358 ( .A1(n18563), .A2(n17261), .ZN(n14422) );
  AOI211_X1 U16359 ( .C1(n17245), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14429), .B(n14422), .ZN(n14423) );
  OAI21_X1 U16360 ( .B1(n15604), .B2(n17227), .A(n14423), .ZN(n14424) );
  INV_X1 U16361 ( .A(n14424), .ZN(n14425) );
  OAI21_X1 U16362 ( .B1(n14437), .B2(n17224), .A(n14425), .ZN(n14426) );
  INV_X1 U16363 ( .A(n14426), .ZN(n14427) );
  NAND2_X1 U16364 ( .A1(n14428), .A2(n14427), .ZN(P2_U2984) );
  AOI21_X1 U16365 ( .B1(n14430), .B2(n18601), .A(n14429), .ZN(n14434) );
  OAI21_X1 U16366 ( .B1(n14461), .B2(n14462), .A(n16727), .ZN(n14431) );
  NAND2_X1 U16367 ( .A1(n16599), .A2(n14431), .ZN(n14465) );
  OAI21_X1 U16368 ( .B1(n16600), .B2(n14461), .A(n14462), .ZN(n14432) );
  NAND2_X1 U16369 ( .A1(n14465), .A2(n14432), .ZN(n14433) );
  OAI211_X1 U16370 ( .C1(n15604), .C2(n16853), .A(n14434), .B(n14433), .ZN(
        n14435) );
  AOI21_X1 U16371 ( .B1(n14436), .B2(n18604), .A(n14435), .ZN(n14439) );
  NAND2_X1 U16372 ( .A1(n14439), .A2(n14438), .ZN(P2_U3016) );
  NOR2_X1 U16373 ( .A1(n14444), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n14445) );
  MUX2_X1 U16374 ( .A(n11911), .B(n14445), .S(n19400), .Z(n18549) );
  NAND2_X1 U16375 ( .A1(n18549), .A2(n14446), .ZN(n14447) );
  INV_X1 U16376 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n18550) );
  AOI22_X1 U16377 ( .A1(n14450), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n14451) );
  OAI21_X1 U16378 ( .B1(n14452), .B2(n18550), .A(n14451), .ZN(n14453) );
  AOI21_X1 U16379 ( .B1(n14454), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n14453), .ZN(n14455) );
  XNOR2_X1 U16380 ( .A(n14456), .B(n14455), .ZN(n16196) );
  INV_X1 U16381 ( .A(n16196), .ZN(n14473) );
  AOI22_X1 U16382 ( .A1(n12488), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n13836), .B2(P2_EAX_REG_31__SCAN_IN), .ZN(n14458) );
  NAND2_X1 U16383 ( .A1(n12280), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14457) );
  AND2_X1 U16384 ( .A1(n14458), .A2(n14457), .ZN(n14459) );
  NOR2_X1 U16385 ( .A1(n18583), .A2(n18550), .ZN(n14470) );
  INV_X1 U16386 ( .A(n14470), .ZN(n14463) );
  OAI211_X1 U16387 ( .C1(n16871), .C2(n16279), .A(n14463), .B(n11370), .ZN(
        n14464) );
  NAND2_X1 U16388 ( .A1(n14465), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14466) );
  INV_X1 U16389 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14468) );
  NAND2_X1 U16390 ( .A1(n14469), .A2(n17216), .ZN(n14472) );
  AOI21_X1 U16391 ( .B1(n17245), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14470), .ZN(n14471) );
  OAI21_X1 U16392 ( .B1(n14473), .B2(n17227), .A(n11364), .ZN(n14474) );
  AOI21_X1 U16393 ( .B1(n14475), .B2(n17258), .A(n14474), .ZN(n14477) );
  NAND2_X1 U16394 ( .A1(n11007), .A2(n17256), .ZN(n14476) );
  NAND2_X1 U16395 ( .A1(n14477), .A2(n14476), .ZN(P2_U2983) );
  INV_X1 U16396 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20090) );
  NOR3_X1 U16397 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n20090), .ZN(n14479) );
  NOR4_X1 U16398 ( .A1(P1_ADS_N_REG_SCAN_IN), .A2(P1_D_C_N_REG_SCAN_IN), .A3(
        P1_BE_N_REG_1__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n14478) );
  NAND4_X1 U16399 ( .A1(n15121), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n14479), .A4(
        n14478), .ZN(U214) );
  NOR2_X1 U16400 ( .A1(P2_BE_N_REG_3__SCAN_IN), .A2(P2_BE_N_REG_2__SCAN_IN), 
        .ZN(n14481) );
  NOR4_X1 U16401 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n14480) );
  NAND4_X1 U16402 ( .A1(n14481), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n14480), .ZN(n14482) );
  OR2_X1 U16403 ( .A1(n15195), .A2(n14482), .ZN(n20027) );
  INV_X2 U16404 ( .A(U214), .ZN(n20078) );
  OR2_X1 U16405 ( .A1(n20027), .A2(n20078), .ZN(U212) );
  NOR2_X1 U16406 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n14482), .ZN(n18712)
         );
  AOI211_X1 U16407 ( .C1(n16562), .C2(n14483), .A(n18663), .B(n18376), .ZN(
        n14495) );
  INV_X1 U16408 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n15343) );
  OAI22_X1 U16409 ( .A1(n18557), .A2(n15343), .B1(n16558), .B2(n18554), .ZN(
        n14494) );
  NOR2_X1 U16410 ( .A1(n18663), .A2(n18562), .ZN(n15069) );
  AOI22_X1 U16411 ( .A1(n14484), .A2(n18534), .B1(n16562), .B2(n15069), .ZN(
        n14485) );
  OAI211_X1 U16412 ( .C1(n12171), .C2(n18551), .A(n14485), .B(n18582), .ZN(
        n14493) );
  XNOR2_X1 U16413 ( .A(n14486), .B(n18358), .ZN(n19164) );
  NAND2_X1 U16414 ( .A1(n14488), .A2(n14487), .ZN(n14491) );
  INV_X1 U16415 ( .A(n14489), .ZN(n14490) );
  NAND2_X1 U16416 ( .A1(n14491), .A2(n14490), .ZN(n16559) );
  OAI22_X1 U16417 ( .A1(n18567), .A2(n19164), .B1(n18447), .B2(n16559), .ZN(
        n14492) );
  OR4_X1 U16418 ( .A1(n14495), .A2(n14494), .A3(n14493), .A4(n14492), .ZN(
        P2_U2842) );
  NAND2_X1 U16419 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n17743) );
  NOR2_X1 U16420 ( .A1(n20095), .A2(n17743), .ZN(n16910) );
  INV_X1 U16421 ( .A(n20777), .ZN(n14496) );
  AOI21_X1 U16422 ( .B1(n14496), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16905) );
  NAND2_X1 U16423 ( .A1(n16905), .A2(n10964), .ZN(n17744) );
  INV_X1 U16424 ( .A(n21235), .ZN(n20094) );
  NOR2_X1 U16425 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n21232), .ZN(
        n21234) );
  AOI21_X1 U16426 ( .B1(n20094), .B2(n17743), .A(n21234), .ZN(n14497) );
  INV_X1 U16427 ( .A(n14497), .ZN(n18717) );
  INV_X1 U16428 ( .A(n19054), .ZN(n19006) );
  INV_X1 U16429 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n21248) );
  INV_X1 U16430 ( .A(n16910), .ZN(n21230) );
  NOR2_X1 U16431 ( .A1(n21248), .A2(n21230), .ZN(n16904) );
  AND2_X1 U16432 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18145), .ZN(
        P3_U2867) );
  INV_X1 U16433 ( .A(n14498), .ZN(n14499) );
  OR2_X1 U16434 ( .A1(n12055), .A2(n14499), .ZN(n15077) );
  INV_X1 U16435 ( .A(n15077), .ZN(n18269) );
  INV_X1 U16436 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n14503) );
  NAND2_X1 U16437 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n17266), .ZN(n18653) );
  INV_X1 U16438 ( .A(n18653), .ZN(n14500) );
  NAND2_X1 U16439 ( .A1(n18640), .A2(n14500), .ZN(n14501) );
  OR2_X1 U16440 ( .A1(n14502), .A2(n14501), .ZN(n14506) );
  OAI211_X1 U16441 ( .C1(n18269), .C2(n14503), .A(n17214), .B(n14506), .ZN(
        P2_U2814) );
  NOR2_X1 U16442 ( .A1(n18248), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n14505)
         );
  AOI22_X1 U16443 ( .A1(n14505), .A2(n17214), .B1(n14504), .B2(n18248), .ZN(
        P2_U3612) );
  INV_X1 U16444 ( .A(n14506), .ZN(n14507) );
  OAI21_X1 U16445 ( .B1(n14506), .B2(n21639), .A(n14622), .ZN(n14568) );
  INV_X1 U16446 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n14508) );
  NAND3_X1 U16447 ( .A1(n14507), .A2(n11774), .A3(n18675), .ZN(n14591) );
  AOI22_X1 U16448 ( .A1(n15196), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n15195), .ZN(n19155) );
  INV_X1 U16449 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19156) );
  OAI222_X1 U16450 ( .A1(n14568), .A2(n14508), .B1(n14591), .B2(n19155), .C1(
        n14622), .C2(n19156), .ZN(P2_U2982) );
  INV_X1 U16451 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n14510) );
  AOI22_X1 U16452 ( .A1(n15196), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n15195), .ZN(n19517) );
  NOR2_X1 U16453 ( .A1(n14591), .A2(n19517), .ZN(n14603) );
  AOI21_X1 U16454 ( .B1(n14606), .B2(P2_EAX_REG_3__SCAN_IN), .A(n14603), .ZN(
        n14509) );
  OAI21_X1 U16455 ( .B1(n14568), .B2(n14510), .A(n14509), .ZN(P2_U2970) );
  INV_X1 U16456 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n14512) );
  AOI22_X1 U16457 ( .A1(n15196), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n15195), .ZN(n19398) );
  NOR2_X1 U16458 ( .A1(n14591), .A2(n19398), .ZN(n14573) );
  AOI21_X1 U16459 ( .B1(n14606), .B2(P2_EAX_REG_5__SCAN_IN), .A(n14573), .ZN(
        n14511) );
  OAI21_X1 U16460 ( .B1(n14568), .B2(n14512), .A(n14511), .ZN(P2_U2972) );
  INV_X1 U16461 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n14515) );
  INV_X1 U16462 ( .A(n14591), .ZN(n14540) );
  AOI22_X1 U16463 ( .A1(n15196), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n15195), .ZN(n19162) );
  INV_X1 U16464 ( .A(n19162), .ZN(n14513) );
  NAND2_X1 U16465 ( .A1(n14540), .A2(n14513), .ZN(n14526) );
  NAND2_X1 U16466 ( .A1(n14606), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n14514) );
  OAI211_X1 U16467 ( .C1(n14568), .C2(n14515), .A(n14526), .B(n14514), .ZN(
        P2_U2980) );
  INV_X1 U16468 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n14518) );
  AOI22_X1 U16469 ( .A1(n15196), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n15195), .ZN(n19620) );
  INV_X1 U16470 ( .A(n19620), .ZN(n14516) );
  NAND2_X1 U16471 ( .A1(n14540), .A2(n14516), .ZN(n14535) );
  NAND2_X1 U16472 ( .A1(n14606), .A2(P2_EAX_REG_1__SCAN_IN), .ZN(n14517) );
  OAI211_X1 U16473 ( .C1(n14568), .C2(n14518), .A(n14535), .B(n14517), .ZN(
        P2_U2968) );
  INV_X1 U16474 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n14791) );
  INV_X1 U16475 ( .A(n14568), .ZN(n14542) );
  NAND2_X1 U16476 ( .A1(n14542), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n14519) );
  NAND2_X1 U16477 ( .A1(n14540), .A2(n19158), .ZN(n14543) );
  OAI211_X1 U16478 ( .C1(n14791), .C2(n14622), .A(n14519), .B(n14543), .ZN(
        P2_U2966) );
  INV_X1 U16479 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19179) );
  NAND2_X1 U16480 ( .A1(n14542), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n14522) );
  NAND2_X1 U16481 ( .A1(n15195), .A2(BUF2_REG_9__SCAN_IN), .ZN(n14521) );
  INV_X1 U16482 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n20046) );
  OR2_X1 U16483 ( .A1(n15195), .A2(n20046), .ZN(n14520) );
  NAND2_X1 U16484 ( .A1(n14521), .A2(n14520), .ZN(n19176) );
  NAND2_X1 U16485 ( .A1(n14540), .A2(n19176), .ZN(n14528) );
  OAI211_X1 U16486 ( .C1(n19179), .C2(n14622), .A(n14522), .B(n14528), .ZN(
        P2_U2976) );
  INV_X1 U16487 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n14774) );
  NAND2_X1 U16488 ( .A1(n14542), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n14525) );
  NAND2_X1 U16489 ( .A1(n15195), .A2(BUF2_REG_10__SCAN_IN), .ZN(n14524) );
  INV_X1 U16490 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n20048) );
  OR2_X1 U16491 ( .A1(n15195), .A2(n20048), .ZN(n14523) );
  NAND2_X1 U16492 ( .A1(n14524), .A2(n14523), .ZN(n19172) );
  NAND2_X1 U16493 ( .A1(n14540), .A2(n19172), .ZN(n14530) );
  OAI211_X1 U16494 ( .C1(n14774), .C2(n14622), .A(n14525), .B(n14530), .ZN(
        P2_U2962) );
  INV_X1 U16495 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14780) );
  NAND2_X1 U16496 ( .A1(n14542), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n14527) );
  OAI211_X1 U16497 ( .C1(n14622), .C2(n14780), .A(n14527), .B(n14526), .ZN(
        P2_U2965) );
  INV_X1 U16498 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n14630) );
  NAND2_X1 U16499 ( .A1(n14542), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n14529) );
  OAI211_X1 U16500 ( .C1(n14622), .C2(n14630), .A(n14529), .B(n14528), .ZN(
        P2_U2961) );
  INV_X1 U16501 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n17315) );
  NAND2_X1 U16502 ( .A1(n14542), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n14531) );
  OAI211_X1 U16503 ( .C1(n17315), .C2(n14622), .A(n14531), .B(n14530), .ZN(
        P2_U2977) );
  INV_X1 U16504 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19168) );
  NAND2_X1 U16505 ( .A1(n14542), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n14534) );
  NAND2_X1 U16506 ( .A1(n15195), .A2(BUF2_REG_12__SCAN_IN), .ZN(n14533) );
  INV_X1 U16507 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n20052) );
  OR2_X1 U16508 ( .A1(n15195), .A2(n20052), .ZN(n14532) );
  NAND2_X1 U16509 ( .A1(n14533), .A2(n14532), .ZN(n19165) );
  NAND2_X1 U16510 ( .A1(n14540), .A2(n19165), .ZN(n14537) );
  OAI211_X1 U16511 ( .C1(n19168), .C2(n14622), .A(n14534), .B(n14537), .ZN(
        P2_U2979) );
  INV_X1 U16512 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14788) );
  NAND2_X1 U16513 ( .A1(n14542), .A2(P2_UWORD_REG_1__SCAN_IN), .ZN(n14536) );
  OAI211_X1 U16514 ( .C1(n14622), .C2(n14788), .A(n14536), .B(n14535), .ZN(
        P2_U2953) );
  INV_X1 U16515 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n14776) );
  NAND2_X1 U16516 ( .A1(n14542), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n14538) );
  OAI211_X1 U16517 ( .C1(n14776), .C2(n14622), .A(n14538), .B(n14537), .ZN(
        P2_U2964) );
  INV_X1 U16518 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14782) );
  NAND2_X1 U16519 ( .A1(n14542), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n14541) );
  AOI22_X1 U16520 ( .A1(n15196), .A2(BUF1_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n15195), .ZN(n19169) );
  INV_X1 U16521 ( .A(n19169), .ZN(n14539) );
  NAND2_X1 U16522 ( .A1(n14540), .A2(n14539), .ZN(n14608) );
  OAI211_X1 U16523 ( .C1(n14622), .C2(n14782), .A(n14541), .B(n14608), .ZN(
        P2_U2963) );
  INV_X1 U16524 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19161) );
  NAND2_X1 U16525 ( .A1(n14542), .A2(P2_LWORD_REG_14__SCAN_IN), .ZN(n14544) );
  OAI211_X1 U16526 ( .C1(n19161), .C2(n14622), .A(n14544), .B(n14543), .ZN(
        P2_U2981) );
  INV_X1 U16527 ( .A(n15608), .ZN(n14545) );
  NAND2_X1 U16528 ( .A1(n14545), .A2(n13523), .ZN(n22311) );
  AOI22_X1 U16529 ( .A1(n15613), .A2(n14724), .B1(n14546), .B2(n22311), .ZN(
        n15619) );
  INV_X1 U16530 ( .A(P1_CODEFETCH_REG_SCAN_IN), .ZN(n17168) );
  AOI21_X1 U16531 ( .B1(n15619), .B2(n15620), .A(n17168), .ZN(n14548) );
  INV_X1 U16532 ( .A(n15582), .ZN(n16171) );
  NOR3_X1 U16533 ( .A1(n16171), .A2(P1_STATE2_REG_2__SCAN_IN), .A3(n16946), 
        .ZN(n14547) );
  OR2_X1 U16534 ( .A1(n14548), .A2(n14547), .ZN(P1_U2803) );
  NOR2_X1 U16535 ( .A1(n14549), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14550) );
  NOR2_X1 U16536 ( .A1(n14551), .A2(n14550), .ZN(n14677) );
  XNOR2_X1 U16537 ( .A(n18255), .B(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14676) );
  OR2_X1 U16538 ( .A1(n18583), .A2(n17283), .ZN(n14678) );
  OAI21_X1 U16539 ( .B1(n17228), .B2(n14676), .A(n14678), .ZN(n14552) );
  AOI21_X1 U16540 ( .B1(n17256), .B2(n14677), .A(n14552), .ZN(n14555) );
  OAI21_X1 U16541 ( .B1(n17245), .B2(n14553), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14554) );
  OAI211_X1 U16542 ( .C1(n18258), .C2(n17227), .A(n14555), .B(n14554), .ZN(
        P2_U3014) );
  XNOR2_X1 U16543 ( .A(n14557), .B(n14556), .ZN(n14672) );
  INV_X1 U16544 ( .A(n14672), .ZN(n14566) );
  OAI21_X1 U16545 ( .B1(n14560), .B2(n14559), .A(n14558), .ZN(n14666) );
  INV_X1 U16546 ( .A(n15032), .ZN(n14563) );
  INV_X1 U16547 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n15035) );
  OR2_X1 U16548 ( .A1(n18582), .A2(n14561), .ZN(n14664) );
  OAI21_X1 U16549 ( .B1(n17222), .B2(n15035), .A(n14664), .ZN(n14562) );
  AOI21_X1 U16550 ( .B1(n17216), .B2(n14563), .A(n14562), .ZN(n14564) );
  OAI21_X1 U16551 ( .B1(n14666), .B2(n17224), .A(n14564), .ZN(n14565) );
  AOI21_X1 U16552 ( .B1(n14566), .B2(n17258), .A(n14565), .ZN(n14567) );
  OAI21_X1 U16553 ( .B1(n15329), .B2(n17227), .A(n14567), .ZN(P2_U3012) );
  INV_X1 U16554 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n14570) );
  INV_X1 U16555 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n20040) );
  INV_X1 U16556 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n20600) );
  AOI22_X1 U16557 ( .A1(n15196), .A2(n20040), .B1(n20600), .B2(n15195), .ZN(
        n19342) );
  INV_X1 U16558 ( .A(n19342), .ZN(n19351) );
  NOR2_X1 U16559 ( .A1(n14591), .A2(n19351), .ZN(n14578) );
  AOI21_X1 U16560 ( .B1(n14606), .B2(P2_EAX_REG_6__SCAN_IN), .A(n14578), .ZN(
        n14569) );
  OAI21_X1 U16561 ( .B1(n14610), .B2(n14570), .A(n14569), .ZN(P2_U2973) );
  INV_X1 U16562 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n14572) );
  AOI22_X1 U16563 ( .A1(n15196), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n15195), .ZN(n19183) );
  NOR2_X1 U16564 ( .A1(n14591), .A2(n19183), .ZN(n14581) );
  AOI21_X1 U16565 ( .B1(n14606), .B2(P2_EAX_REG_23__SCAN_IN), .A(n14581), .ZN(
        n14571) );
  OAI21_X1 U16566 ( .B1(n14610), .B2(n14572), .A(n14571), .ZN(P2_U2959) );
  INV_X1 U16567 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n14575) );
  AOI21_X1 U16568 ( .B1(n14606), .B2(P2_EAX_REG_21__SCAN_IN), .A(n14573), .ZN(
        n14574) );
  OAI21_X1 U16569 ( .B1(n14610), .B2(n14575), .A(n14574), .ZN(P2_U2957) );
  INV_X1 U16570 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n14577) );
  OAI22_X1 U16571 ( .A1(n15195), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n15196), .ZN(n19684) );
  NOR2_X1 U16572 ( .A1(n14591), .A2(n19684), .ZN(n14597) );
  AOI21_X1 U16573 ( .B1(n14606), .B2(P2_EAX_REG_0__SCAN_IN), .A(n14597), .ZN(
        n14576) );
  OAI21_X1 U16574 ( .B1(n14610), .B2(n14577), .A(n14576), .ZN(P2_U2967) );
  INV_X1 U16575 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n14580) );
  AOI21_X1 U16576 ( .B1(n14606), .B2(P2_EAX_REG_22__SCAN_IN), .A(n14578), .ZN(
        n14579) );
  OAI21_X1 U16577 ( .B1(n14610), .B2(n14580), .A(n14579), .ZN(P2_U2958) );
  INV_X1 U16578 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n14583) );
  AOI21_X1 U16579 ( .B1(n14606), .B2(P2_EAX_REG_7__SCAN_IN), .A(n14581), .ZN(
        n14582) );
  OAI21_X1 U16580 ( .B1(n14610), .B2(n14583), .A(n14582), .ZN(P2_U2974) );
  INV_X1 U16581 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n14585) );
  AOI22_X1 U16582 ( .A1(n15196), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n15195), .ZN(n19565) );
  NOR2_X1 U16583 ( .A1(n14591), .A2(n19565), .ZN(n14588) );
  AOI21_X1 U16584 ( .B1(n14606), .B2(P2_EAX_REG_18__SCAN_IN), .A(n14588), .ZN(
        n14584) );
  OAI21_X1 U16585 ( .B1(n14610), .B2(n14585), .A(n14584), .ZN(P2_U2954) );
  INV_X1 U16586 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n14587) );
  INV_X1 U16587 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n20036) );
  INV_X1 U16588 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n20611) );
  AOI22_X1 U16589 ( .A1(n15196), .A2(n20036), .B1(n20611), .B2(n15195), .ZN(
        n19439) );
  INV_X1 U16590 ( .A(n19439), .ZN(n19461) );
  NOR2_X1 U16591 ( .A1(n14591), .A2(n19461), .ZN(n14600) );
  AOI21_X1 U16592 ( .B1(n14606), .B2(P2_EAX_REG_20__SCAN_IN), .A(n14600), .ZN(
        n14586) );
  OAI21_X1 U16593 ( .B1(n14610), .B2(n14587), .A(n14586), .ZN(P2_U2956) );
  INV_X1 U16594 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n14590) );
  AOI21_X1 U16595 ( .B1(P2_EAX_REG_2__SCAN_IN), .B2(n14606), .A(n14588), .ZN(
        n14589) );
  OAI21_X1 U16596 ( .B1(n14610), .B2(n14590), .A(n14589), .ZN(P2_U2969) );
  INV_X1 U16597 ( .A(P2_UWORD_REG_8__SCAN_IN), .ZN(n14593) );
  AOI22_X1 U16598 ( .A1(n15196), .A2(BUF1_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n15195), .ZN(n19182) );
  NOR2_X1 U16599 ( .A1(n14591), .A2(n19182), .ZN(n14594) );
  AOI21_X1 U16600 ( .B1(n14606), .B2(P2_EAX_REG_24__SCAN_IN), .A(n14594), .ZN(
        n14592) );
  OAI21_X1 U16601 ( .B1(n14610), .B2(n14593), .A(n14592), .ZN(P2_U2960) );
  INV_X1 U16602 ( .A(P2_LWORD_REG_8__SCAN_IN), .ZN(n14596) );
  AOI21_X1 U16603 ( .B1(n14606), .B2(P2_EAX_REG_8__SCAN_IN), .A(n14594), .ZN(
        n14595) );
  OAI21_X1 U16604 ( .B1(n14610), .B2(n14596), .A(n14595), .ZN(P2_U2975) );
  INV_X1 U16605 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n14599) );
  AOI21_X1 U16606 ( .B1(n14606), .B2(P2_EAX_REG_16__SCAN_IN), .A(n14597), .ZN(
        n14598) );
  OAI21_X1 U16607 ( .B1(n14610), .B2(n14599), .A(n14598), .ZN(P2_U2952) );
  INV_X1 U16608 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n14602) );
  AOI21_X1 U16609 ( .B1(n14606), .B2(P2_EAX_REG_4__SCAN_IN), .A(n14600), .ZN(
        n14601) );
  OAI21_X1 U16610 ( .B1(n14610), .B2(n14602), .A(n14601), .ZN(P2_U2971) );
  INV_X1 U16611 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n14605) );
  AOI21_X1 U16612 ( .B1(n14606), .B2(P2_EAX_REG_19__SCAN_IN), .A(n14603), .ZN(
        n14604) );
  OAI21_X1 U16613 ( .B1(n14610), .B2(n14605), .A(n14604), .ZN(P2_U2955) );
  INV_X1 U16614 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n14609) );
  NAND2_X1 U16615 ( .A1(n14606), .A2(P2_EAX_REG_11__SCAN_IN), .ZN(n14607) );
  OAI211_X1 U16616 ( .C1(n14610), .C2(n14609), .A(n14608), .B(n14607), .ZN(
        P2_U2978) );
  INV_X1 U16617 ( .A(n14614), .ZN(n14611) );
  AOI222_X1 U16618 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14614), .B1(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n14613), .C1(n14612), .C2(
        n14611), .ZN(n14818) );
  OAI21_X1 U16619 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n14616), .A(
        n14615), .ZN(n14617) );
  INV_X1 U16620 ( .A(n14617), .ZN(n14811) );
  NAND2_X1 U16621 ( .A1(n17256), .A2(n14811), .ZN(n14618) );
  NAND2_X1 U16622 ( .A1(n18382), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n14812) );
  OAI211_X1 U16623 ( .C1(n15068), .C2(n17222), .A(n14618), .B(n14812), .ZN(
        n14620) );
  NOR2_X1 U16624 ( .A1(n17261), .A2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14619) );
  AOI211_X1 U16625 ( .C1(n17257), .C2(n15074), .A(n14620), .B(n14619), .ZN(
        n14621) );
  OAI21_X1 U16626 ( .B1(n14818), .B2(n17228), .A(n14621), .ZN(P2_U3013) );
  INV_X1 U16627 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14626) );
  OR2_X1 U16628 ( .A1(n12055), .A2(n18657), .ZN(n14623) );
  OAI21_X1 U16629 ( .B1(n14636), .B2(n14623), .A(n14622), .ZN(n14624) );
  NAND2_X1 U16630 ( .A1(n17294), .A2(n18240), .ZN(n14790) );
  NOR2_X1 U16631 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15190), .ZN(n17313) );
  AOI22_X1 U16632 ( .A1(n17321), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n17307), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n14625) );
  OAI21_X1 U16633 ( .B1(n14626), .B2(n14790), .A(n14625), .ZN(P2_U2929) );
  INV_X1 U16634 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n14628) );
  AOI22_X1 U16635 ( .A1(n17321), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n17307), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n14627) );
  OAI21_X1 U16636 ( .B1(n14628), .B2(n14790), .A(n14627), .ZN(P2_U2930) );
  AOI22_X1 U16637 ( .A1(n17321), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n17307), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n14629) );
  OAI21_X1 U16638 ( .B1(n14630), .B2(n14790), .A(n14629), .ZN(P2_U2926) );
  INV_X1 U16639 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n16333) );
  AOI22_X1 U16640 ( .A1(n17321), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n17307), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n14631) );
  OAI21_X1 U16641 ( .B1(n16333), .B2(n14790), .A(n14631), .ZN(P2_U2928) );
  INV_X1 U16642 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n14633) );
  AOI22_X1 U16643 ( .A1(n17321), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n17307), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n14632) );
  OAI21_X1 U16644 ( .B1(n14633), .B2(n14790), .A(n14632), .ZN(P2_U2927) );
  NOR2_X1 U16645 ( .A1(n18669), .A2(n15190), .ZN(n18665) );
  INV_X1 U16646 ( .A(n18626), .ZN(n18637) );
  INV_X1 U16647 ( .A(n15317), .ZN(n18625) );
  NAND2_X1 U16648 ( .A1(n18637), .A2(n18625), .ZN(n14694) );
  AND3_X1 U16649 ( .A1(n14635), .A2(n14694), .A3(n14634), .ZN(n14640) );
  INV_X1 U16650 ( .A(n14636), .ZN(n14638) );
  INV_X1 U16651 ( .A(n12055), .ZN(n14643) );
  NAND3_X1 U16652 ( .A1(n14638), .A2(n14643), .A3(n14637), .ZN(n14639) );
  OAI22_X1 U16653 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19233), .B1(n18611), 
        .B2(n18657), .ZN(n14641) );
  AOI21_X1 U16654 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n18665), .A(n14641), .ZN(
        n16897) );
  INV_X1 U16655 ( .A(n16897), .ZN(n14645) );
  NOR2_X1 U16656 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15334) );
  INV_X1 U16657 ( .A(n15334), .ZN(n18658) );
  NAND2_X1 U16658 ( .A1(n14643), .A2(n14642), .ZN(n18642) );
  OR4_X1 U16659 ( .A1(n16897), .A2(n18658), .A3(n11774), .A4(n18642), .ZN(
        n14644) );
  OAI21_X1 U16660 ( .B1(n14646), .B2(n14645), .A(n14644), .ZN(P2_U3595) );
  NOR2_X1 U16661 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n14649) );
  NOR2_X1 U16662 ( .A1(n14651), .A2(n14650), .ZN(n14652) );
  OR2_X1 U16663 ( .A1(n14653), .A2(n14652), .ZN(n14675) );
  INV_X1 U16664 ( .A(n14675), .ZN(n18254) );
  NOR2_X1 U16665 ( .A1(n15383), .A2(n14675), .ZN(n19614) );
  INV_X1 U16666 ( .A(n19614), .ZN(n14654) );
  INV_X1 U16667 ( .A(n19677), .ZN(n19561) );
  OAI211_X1 U16668 ( .C1(n18260), .C2(n18254), .A(n14654), .B(n19561), .ZN(
        n14656) );
  AOI22_X1 U16669 ( .A1(n19612), .A2(n18254), .B1(n19670), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n14655) );
  OAI211_X1 U16670 ( .C1(n19619), .C2(n19684), .A(n14656), .B(n14655), .ZN(
        P2_U2919) );
  NAND2_X1 U16671 ( .A1(n21925), .A2(n16973), .ZN(n15449) );
  AND2_X1 U16672 ( .A1(n14802), .A2(n15449), .ZN(n22312) );
  INV_X1 U16673 ( .A(n22312), .ZN(n14659) );
  OAI33_X1 U16674 ( .A1(n14659), .A2(P1_READREQUEST_REG_SCAN_IN), .A3(n14658), 
        .B1(n13547), .B2(n15093), .B3(n14657), .ZN(n14660) );
  INV_X1 U16675 ( .A(n14660), .ZN(P1_U3487) );
  XNOR2_X1 U16676 ( .A(n14662), .B(n14661), .ZN(n19558) );
  INV_X1 U16677 ( .A(n16867), .ZN(n15308) );
  INV_X1 U16678 ( .A(n15307), .ZN(n15304) );
  NAND2_X1 U16679 ( .A1(n16829), .A2(n15304), .ZN(n14663) );
  NAND2_X1 U16680 ( .A1(n15308), .A2(n14663), .ZN(n14665) );
  OAI211_X1 U16681 ( .C1(n14666), .C2(n18609), .A(n14665), .B(n14664), .ZN(
        n14667) );
  INV_X1 U16682 ( .A(n14667), .ZN(n14671) );
  NOR2_X1 U16683 ( .A1(n16826), .A2(n14668), .ZN(n15305) );
  OAI21_X1 U16684 ( .B1(n16826), .B2(n14814), .A(n16830), .ZN(n14669) );
  AOI22_X1 U16685 ( .A1(n15305), .A2(n14814), .B1(n14669), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14670) );
  OAI211_X1 U16686 ( .C1(n14672), .C2(n18575), .A(n14671), .B(n14670), .ZN(
        n14673) );
  AOI21_X1 U16687 ( .B1(n18601), .B2(n19558), .A(n14673), .ZN(n14674) );
  OAI21_X1 U16688 ( .B1(n15329), .B2(n16853), .A(n14674), .ZN(P2_U3044) );
  INV_X1 U16689 ( .A(n16764), .ZN(n16696) );
  OAI22_X1 U16690 ( .A1(n14676), .A2(n18575), .B1(n16871), .B2(n14675), .ZN(
        n14681) );
  NAND2_X1 U16691 ( .A1(n16864), .A2(n14677), .ZN(n14679) );
  OAI211_X1 U16692 ( .C1(n16830), .C2(n14682), .A(n14679), .B(n14678), .ZN(
        n14680) );
  AOI211_X1 U16693 ( .C1(n14682), .C2(n16696), .A(n14681), .B(n14680), .ZN(
        n14683) );
  OAI21_X1 U16694 ( .B1(n18258), .B2(n16853), .A(n14683), .ZN(P2_U3046) );
  OR2_X1 U16695 ( .A1(n14684), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14686) );
  NAND2_X1 U16696 ( .A1(n14686), .A2(n14685), .ZN(n21410) );
  AND2_X1 U16697 ( .A1(n14729), .A2(n14687), .ZN(n15609) );
  NAND2_X1 U16698 ( .A1(n15613), .A2(n15609), .ZN(n14710) );
  OR2_X1 U16699 ( .A1(n14688), .A2(n10976), .ZN(n14689) );
  NAND2_X1 U16700 ( .A1(n14710), .A2(n14689), .ZN(n14690) );
  OAI21_X1 U16701 ( .B1(n14693), .B2(n14692), .A(n14691), .ZN(n19955) );
  INV_X2 U16702 ( .A(n19942), .ZN(n15842) );
  OAI222_X1 U16703 ( .A1(n21410), .A2(n15837), .B1(n13538), .B2(n19946), .C1(
        n19955), .C2(n15842), .ZN(P1_U2872) );
  NAND2_X1 U16704 ( .A1(n14694), .A2(n15324), .ZN(n14695) );
  NAND2_X2 U16705 ( .A1(n14695), .A2(n18683), .ZN(n16267) );
  NAND2_X1 U16706 ( .A1(n16209), .A2(n15200), .ZN(n16278) );
  MUX2_X1 U16707 ( .A(n18258), .B(n14696), .S(n16267), .Z(n14697) );
  OAI21_X1 U16708 ( .B1(n15383), .B2(n16278), .A(n14697), .ZN(P2_U2887) );
  INV_X1 U16709 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n14699) );
  AOI22_X1 U16710 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n17320), .B1(n17321), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n14698) );
  OAI21_X1 U16711 ( .B1(n14699), .B2(n14790), .A(n14698), .ZN(P2_U2935) );
  INV_X1 U16712 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n21902) );
  NOR2_X1 U16713 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21902), .ZN(n21593) );
  OAI21_X1 U16714 ( .B1(n21624), .B2(n21633), .A(n14700), .ZN(n14701) );
  OAI21_X1 U16715 ( .B1(n16162), .B2(n14702), .A(n14701), .ZN(n14711) );
  AOI21_X1 U16716 ( .B1(n14703), .B2(n12623), .A(n14719), .ZN(n14704) );
  NAND2_X1 U16717 ( .A1(n14705), .A2(n14704), .ZN(n14722) );
  AND2_X1 U16718 ( .A1(n14706), .A2(n14722), .ZN(n14707) );
  NOR2_X1 U16719 ( .A1(n14707), .A2(n13523), .ZN(n14853) );
  NOR2_X1 U16720 ( .A1(n15096), .A2(n14850), .ZN(n14708) );
  NOR2_X1 U16721 ( .A1(n14853), .A2(n14708), .ZN(n14709) );
  OAI211_X1 U16722 ( .C1(n15613), .C2(n14711), .A(n14710), .B(n14709), .ZN(
        n14713) );
  OR2_X1 U16723 ( .A1(n14713), .A2(n14712), .ZN(n16947) );
  NOR2_X1 U16724 ( .A1(n16946), .A2(n16973), .ZN(n21588) );
  AND2_X1 U16725 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21588), .ZN(n21592) );
  AOI22_X1 U16726 ( .A1(n16947), .A2(n15620), .B1(P1_FLUSH_REG_SCAN_IN), .B2(
        n21592), .ZN(n14714) );
  INV_X1 U16727 ( .A(n14714), .ZN(n14792) );
  NOR2_X1 U16728 ( .A1(n21593), .A2(n14792), .ZN(n16172) );
  NAND2_X1 U16729 ( .A1(n14716), .A2(n12628), .ZN(n14721) );
  INV_X1 U16730 ( .A(n15096), .ZN(n14728) );
  NAND2_X1 U16731 ( .A1(n14728), .A2(n14717), .ZN(n14718) );
  OAI21_X1 U16732 ( .B1(n12626), .B2(n14719), .A(n14718), .ZN(n14720) );
  AOI21_X1 U16733 ( .B1(n14721), .B2(n12623), .A(n14720), .ZN(n14723) );
  OAI211_X1 U16734 ( .C1(n12635), .C2(n14724), .A(n14723), .B(n14722), .ZN(
        n14868) );
  NAND3_X1 U16735 ( .A1(n14846), .A2(n14725), .A3(n14866), .ZN(n14726) );
  NOR2_X1 U16736 ( .A1(n14868), .A2(n14726), .ZN(n14727) );
  NAND2_X1 U16737 ( .A1(n14727), .A2(n13349), .ZN(n15579) );
  INV_X1 U16738 ( .A(n15579), .ZN(n16164) );
  XNOR2_X1 U16739 ( .A(n16161), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14734) );
  NOR2_X1 U16740 ( .A1(n14728), .A2(n14800), .ZN(n15618) );
  NAND2_X1 U16741 ( .A1(n14729), .A2(n15618), .ZN(n14743) );
  INV_X1 U16742 ( .A(n14743), .ZN(n14733) );
  XNOR2_X1 U16743 ( .A(n14730), .B(n14731), .ZN(n14737) );
  INV_X1 U16744 ( .A(n14737), .ZN(n14732) );
  AOI22_X1 U16745 ( .A1(n16162), .A2(n14734), .B1(n14733), .B2(n14732), .ZN(
        n14736) );
  NAND3_X1 U16746 ( .A1(n16164), .A2(n12627), .A3(n14737), .ZN(n14735) );
  OAI211_X1 U16747 ( .C1(n14715), .C2(n16164), .A(n14736), .B(n14735), .ZN(
        n14889) );
  OAI22_X1 U16748 ( .A1(n13533), .A2(n16038), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n16165) );
  INV_X1 U16749 ( .A(n16165), .ZN(n14738) );
  INV_X1 U16750 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21400) );
  NOR2_X1 U16751 ( .A1(n16973), .A2(n21400), .ZN(n16166) );
  AOI222_X1 U16752 ( .A1(n14889), .A2(n15582), .B1(n14738), .B2(n16166), .C1(
        n21597), .C2(n14737), .ZN(n14740) );
  NAND2_X1 U16753 ( .A1(n16172), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14739) );
  OAI21_X1 U16754 ( .B1(n16172), .B2(n14740), .A(n14739), .ZN(P1_U3472) );
  INV_X1 U16755 ( .A(n21771), .ZN(n15239) );
  AOI21_X1 U16756 ( .B1(n14730), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n14746), .ZN(n14741) );
  NOR2_X1 U16757 ( .A1(n12737), .A2(n14741), .ZN(n14755) );
  NOR3_X1 U16758 ( .A1(n15579), .A2(n14755), .A3(n12628), .ZN(n14753) );
  INV_X1 U16759 ( .A(n16162), .ZN(n15581) );
  NAND2_X1 U16760 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14745) );
  INV_X1 U16761 ( .A(n14745), .ZN(n14742) );
  NOR2_X1 U16762 ( .A1(n15581), .A2(n14742), .ZN(n14748) );
  NOR2_X1 U16763 ( .A1(n14730), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n14744) );
  OAI22_X1 U16764 ( .A1(n15581), .A2(n14745), .B1(n14744), .B2(n14743), .ZN(
        n14747) );
  MUX2_X1 U16765 ( .A(n14748), .B(n14747), .S(n14746), .Z(n14752) );
  INV_X1 U16766 ( .A(n14749), .ZN(n14750) );
  NOR2_X1 U16767 ( .A1(n14730), .A2(n14750), .ZN(n14751) );
  NOR3_X1 U16768 ( .A1(n14753), .A2(n14752), .A3(n14751), .ZN(n14754) );
  OAI21_X1 U16769 ( .B1(n15239), .B2(n16164), .A(n14754), .ZN(n14888) );
  INV_X1 U16770 ( .A(n14755), .ZN(n14756) );
  AOI22_X1 U16771 ( .A1(n14888), .A2(n15582), .B1(n21597), .B2(n14756), .ZN(
        n14758) );
  NAND2_X1 U16772 ( .A1(n16172), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n14757) );
  OAI21_X1 U16773 ( .B1(n16172), .B2(n14758), .A(n14757), .ZN(P1_U3469) );
  OAI21_X1 U16774 ( .B1(n19453), .B2(n16278), .A(n14763), .ZN(P2_U2884) );
  INV_X1 U16775 ( .A(n19447), .ZN(n19448) );
  NOR2_X1 U16776 ( .A1(n11771), .A2(n16267), .ZN(n14766) );
  AOI21_X1 U16777 ( .B1(P2_EBX_REG_1__SCAN_IN), .B2(n16267), .A(n14766), .ZN(
        n14767) );
  OAI21_X1 U16778 ( .B1(n19448), .B2(n16278), .A(n14767), .ZN(P2_U2886) );
  INV_X1 U16779 ( .A(n14768), .ZN(n14769) );
  INV_X1 U16780 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n14771) );
  MUX2_X1 U16781 ( .A(n14771), .B(n15329), .S(n16209), .Z(n14772) );
  OAI21_X1 U16782 ( .B1(n19452), .B2(n16278), .A(n14772), .ZN(P2_U2885) );
  AOI22_X1 U16783 ( .A1(n17321), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n17320), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n14773) );
  OAI21_X1 U16784 ( .B1(n14774), .B2(n14790), .A(n14773), .ZN(P2_U2925) );
  AOI22_X1 U16785 ( .A1(n17321), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n17320), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n14775) );
  OAI21_X1 U16786 ( .B1(n14776), .B2(n14790), .A(n14775), .ZN(P2_U2923) );
  INV_X1 U16787 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n14778) );
  AOI22_X1 U16788 ( .A1(n17321), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n17320), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n14777) );
  OAI21_X1 U16789 ( .B1(n14778), .B2(n14790), .A(n14777), .ZN(P2_U2931) );
  AOI22_X1 U16790 ( .A1(n17321), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n17320), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n14779) );
  OAI21_X1 U16791 ( .B1(n14780), .B2(n14790), .A(n14779), .ZN(P2_U2922) );
  AOI22_X1 U16792 ( .A1(n17321), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n17320), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n14781) );
  OAI21_X1 U16793 ( .B1(n14782), .B2(n14790), .A(n14781), .ZN(P2_U2924) );
  INV_X1 U16794 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n14784) );
  AOI22_X1 U16795 ( .A1(n17313), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n17320), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n14783) );
  OAI21_X1 U16796 ( .B1(n14784), .B2(n14790), .A(n14783), .ZN(P2_U2933) );
  INV_X1 U16797 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n14786) );
  AOI22_X1 U16798 ( .A1(n17313), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n17320), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n14785) );
  OAI21_X1 U16799 ( .B1(n14786), .B2(n14790), .A(n14785), .ZN(P2_U2932) );
  AOI22_X1 U16800 ( .A1(n17313), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n17320), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n14787) );
  OAI21_X1 U16801 ( .B1(n14788), .B2(n14790), .A(n14787), .ZN(P2_U2934) );
  AOI22_X1 U16802 ( .A1(n17313), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n17320), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n14789) );
  OAI21_X1 U16803 ( .B1(n14791), .B2(n14790), .A(n14789), .ZN(P2_U2921) );
  INV_X1 U16804 ( .A(n16172), .ZN(n15585) );
  NAND2_X1 U16805 ( .A1(n15582), .A2(n14792), .ZN(n14796) );
  INV_X1 U16806 ( .A(n15115), .ZN(n21820) );
  OR2_X1 U16807 ( .A1(n14793), .A2(n21820), .ZN(n14794) );
  XNOR2_X1 U16808 ( .A(n14794), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n21424) );
  INV_X1 U16809 ( .A(n13349), .ZN(n14795) );
  NAND2_X1 U16810 ( .A1(n21424), .A2(n14795), .ZN(n14890) );
  OAI22_X1 U16811 ( .A1(n15585), .A2(n12860), .B1(n14796), .B2(n14890), .ZN(
        P1_U3468) );
  INV_X1 U16812 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n14797) );
  OR2_X1 U16813 ( .A1(n15599), .A2(n14797), .ZN(n14799) );
  NAND2_X1 U16814 ( .A1(n15599), .A2(DATAI_15_), .ZN(n14798) );
  AND2_X1 U16815 ( .A1(n14799), .A2(n14798), .ZN(n15884) );
  NOR2_X1 U16816 ( .A1(n14800), .A2(n21622), .ZN(n14801) );
  OR2_X2 U16817 ( .A1(n14802), .A2(n14801), .ZN(n21729) );
  OR2_X1 U16818 ( .A1(n14846), .A2(n21250), .ZN(n16940) );
  INV_X1 U16819 ( .A(n16940), .ZN(n14803) );
  INV_X1 U16820 ( .A(n21766), .ZN(n21692) );
  AOI22_X1 U16821 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n21729), .B1(n21692), 
        .B2(P1_EAX_REG_15__SCAN_IN), .ZN(n14805) );
  OAI21_X1 U16822 ( .B1(n15884), .B2(n21761), .A(n14805), .ZN(P1_U2967) );
  NAND2_X1 U16823 ( .A1(n14807), .A2(n14806), .ZN(n14810) );
  INV_X1 U16824 ( .A(n14808), .ZN(n14809) );
  AND2_X1 U16825 ( .A1(n14810), .A2(n14809), .ZN(n19449) );
  INV_X1 U16826 ( .A(n16830), .ZN(n15306) );
  AOI22_X1 U16827 ( .A1(n15306), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n16864), .B2(n14811), .ZN(n14813) );
  OAI211_X1 U16828 ( .C1(n19449), .C2(n16871), .A(n14813), .B(n14812), .ZN(
        n14816) );
  AOI211_X1 U16829 ( .C1(n11712), .C2(n14682), .A(n14814), .B(n16764), .ZN(
        n14815) );
  AOI211_X1 U16830 ( .C1(n18603), .C2(n15074), .A(n14816), .B(n14815), .ZN(
        n14817) );
  OAI21_X1 U16831 ( .B1(n14818), .B2(n18575), .A(n14817), .ZN(P2_U3045) );
  NAND2_X1 U16832 ( .A1(n10980), .A2(n14820), .ZN(n14822) );
  NAND2_X1 U16833 ( .A1(n14822), .A2(n14821), .ZN(n14824) );
  OAI21_X1 U16834 ( .B1(n14824), .B2(n14823), .A(n14835), .ZN(n21419) );
  XNOR2_X1 U16835 ( .A(n21415), .B(n10976), .ZN(n14875) );
  INV_X1 U16836 ( .A(n14875), .ZN(n14825) );
  INV_X1 U16837 ( .A(n19946), .ZN(n15840) );
  AOI22_X1 U16838 ( .A1(n19941), .A2(n14825), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n15840), .ZN(n14826) );
  OAI21_X1 U16839 ( .B1(n21419), .B2(n15842), .A(n14826), .ZN(P1_U2871) );
  INV_X1 U16840 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n21714) );
  NAND2_X1 U16841 ( .A1(n21766), .A2(n14827), .ZN(n14828) );
  INV_X1 U16842 ( .A(n21633), .ZN(n15617) );
  NAND2_X1 U16843 ( .A1(n19857), .A2(n15124), .ZN(n15030) );
  NAND2_X1 U16844 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n21583) );
  NOR2_X1 U16845 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n21583), .ZN(n19868) );
  NOR2_X4 U16846 ( .A1(n19857), .A2(n21257), .ZN(n19865) );
  AOI22_X1 U16847 ( .A1(n19868), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n14829) );
  OAI21_X1 U16848 ( .B1(n21714), .B2(n15030), .A(n14829), .ZN(P1_U2913) );
  INV_X1 U16849 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n21708) );
  AOI22_X1 U16850 ( .A1(n21257), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n14830) );
  OAI21_X1 U16851 ( .B1(n21708), .B2(n15030), .A(n14830), .ZN(P1_U2914) );
  INV_X1 U16852 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n21727) );
  AOI22_X1 U16853 ( .A1(n21257), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n14831) );
  OAI21_X1 U16854 ( .B1(n21727), .B2(n15030), .A(n14831), .ZN(P1_U2911) );
  INV_X1 U16855 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n21735) );
  AOI22_X1 U16856 ( .A1(n21257), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n14832) );
  OAI21_X1 U16857 ( .B1(n21735), .B2(n15030), .A(n14832), .ZN(P1_U2910) );
  INV_X1 U16858 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n21720) );
  AOI22_X1 U16859 ( .A1(n21257), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n14833) );
  OAI21_X1 U16860 ( .B1(n21720), .B2(n15030), .A(n14833), .ZN(P1_U2912) );
  XNOR2_X1 U16861 ( .A(n14834), .B(n14835), .ZN(n15107) );
  NOR2_X1 U16862 ( .A1(n14838), .A2(n14837), .ZN(n14839) );
  OR2_X1 U16863 ( .A1(n14836), .A2(n14839), .ZN(n15099) );
  INV_X1 U16864 ( .A(n15099), .ZN(n14840) );
  AOI22_X1 U16865 ( .A1(n19941), .A2(n14840), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n15840), .ZN(n14841) );
  OAI21_X1 U16866 ( .B1(n15107), .B2(n15842), .A(n14841), .ZN(P1_U2870) );
  XNOR2_X1 U16867 ( .A(n14842), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14924) );
  INV_X1 U16868 ( .A(n15613), .ZN(n15610) );
  NAND2_X1 U16869 ( .A1(n14843), .A2(n21622), .ZN(n14845) );
  OAI211_X1 U16870 ( .C1(n14846), .C2(n14845), .A(n15124), .B(n14844), .ZN(
        n14847) );
  NAND2_X1 U16871 ( .A1(n15610), .A2(n14847), .ZN(n14852) );
  NAND2_X1 U16872 ( .A1(n12623), .A2(n21633), .ZN(n14848) );
  NAND2_X1 U16873 ( .A1(n14848), .A2(n21622), .ZN(n14849) );
  OR2_X1 U16874 ( .A1(n15608), .A2(n14849), .ZN(n14851) );
  MUX2_X1 U16875 ( .A(n14852), .B(n14851), .S(n14850), .Z(n14856) );
  NOR2_X1 U16876 ( .A1(n15577), .A2(n16174), .ZN(n14854) );
  AOI21_X1 U16877 ( .B1(n15613), .B2(n14854), .A(n14853), .ZN(n14855) );
  NAND2_X1 U16878 ( .A1(n14856), .A2(n14855), .ZN(n14857) );
  AND2_X1 U16879 ( .A1(n14859), .A2(n14858), .ZN(n15611) );
  NAND2_X1 U16880 ( .A1(n14860), .A2(n14871), .ZN(n14861) );
  NAND4_X1 U16881 ( .A1(n13349), .A2(n15611), .A3(n14862), .A4(n14861), .ZN(
        n14863) );
  INV_X1 U16882 ( .A(n14874), .ZN(n14864) );
  NAND2_X1 U16883 ( .A1(n14864), .A2(n21378), .ZN(n21401) );
  OAI21_X1 U16884 ( .B1(n14866), .B2(n15124), .A(n14865), .ZN(n14867) );
  OR2_X1 U16885 ( .A1(n14868), .A2(n14867), .ZN(n14869) );
  OAI21_X1 U16886 ( .B1(n16041), .B2(n21265), .A(n21400), .ZN(n21407) );
  AOI21_X1 U16887 ( .B1(n21401), .B2(n21407), .A(n13533), .ZN(n14879) );
  INV_X1 U16888 ( .A(n21265), .ZN(n14870) );
  OR2_X1 U16889 ( .A1(n21337), .A2(n16041), .ZN(n16130) );
  NAND2_X1 U16890 ( .A1(n21402), .A2(n21400), .ZN(n14939) );
  AND3_X1 U16891 ( .A1(n16130), .A2(n13533), .A3(n14939), .ZN(n14878) );
  INV_X1 U16892 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n21418) );
  NOR2_X1 U16893 ( .A1(n21378), .A2(n21418), .ZN(n14877) );
  OAI21_X1 U16894 ( .B1(n14872), .B2(n14871), .A(n16940), .ZN(n14873) );
  NOR2_X1 U16895 ( .A1(n21409), .A2(n14875), .ZN(n14876) );
  NOR4_X1 U16896 ( .A1(n14879), .A2(n14878), .A3(n14877), .A4(n14876), .ZN(
        n14880) );
  OAI21_X1 U16897 ( .B1(n14924), .B2(n21327), .A(n14880), .ZN(P1_U3030) );
  XOR2_X1 U16898 ( .A(n14881), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n14887)
         );
  OR2_X1 U16899 ( .A1(n14918), .A2(n14883), .ZN(n14884) );
  AND2_X1 U16900 ( .A1(n14882), .A2(n14884), .ZN(n18286) );
  INV_X1 U16901 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n18278) );
  NOR2_X1 U16902 ( .A1(n16209), .A2(n18278), .ZN(n14885) );
  AOI21_X1 U16903 ( .B1(n18286), .B2(n16209), .A(n14885), .ZN(n14886) );
  OAI21_X1 U16904 ( .B1(n14887), .B2(n16278), .A(n14886), .ZN(P2_U2882) );
  MUX2_X1 U16905 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n14888), .S(
        n16947), .Z(n16962) );
  MUX2_X1 U16906 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14889), .S(
        n16947), .Z(n16957) );
  NAND3_X1 U16907 ( .A1(n16962), .A2(n16973), .A3(n16957), .ZN(n14898) );
  NAND2_X1 U16908 ( .A1(n16947), .A2(n14890), .ZN(n14891) );
  OAI211_X1 U16909 ( .C1(n16947), .C2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n14891), .B(n16973), .ZN(n14893) );
  NOR2_X1 U16910 ( .A1(n16973), .A2(P1_FLUSH_REG_SCAN_IN), .ZN(n14894) );
  NAND2_X1 U16911 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n14894), .ZN(
        n14892) );
  NAND2_X1 U16912 ( .A1(n14893), .A2(n14892), .ZN(n14899) );
  AND2_X1 U16913 ( .A1(n14895), .A2(n14894), .ZN(n14896) );
  NOR2_X1 U16914 ( .A1(n14899), .A2(n14896), .ZN(n14897) );
  NAND2_X1 U16915 ( .A1(n14898), .A2(n14897), .ZN(n16968) );
  INV_X1 U16916 ( .A(n14899), .ZN(n14901) );
  NAND2_X1 U16917 ( .A1(n14901), .A2(n14900), .ZN(n14902) );
  NAND2_X1 U16918 ( .A1(n16968), .A2(n14902), .ZN(n21582) );
  INV_X1 U16919 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n14903) );
  NAND2_X1 U16920 ( .A1(n21582), .A2(n14903), .ZN(n14904) );
  NAND2_X1 U16921 ( .A1(n14904), .A2(n21592), .ZN(n14905) );
  NAND2_X1 U16922 ( .A1(n14905), .A2(n21825), .ZN(n16976) );
  INV_X1 U16923 ( .A(n14906), .ZN(n21938) );
  NAND2_X1 U16924 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21902), .ZN(n21580) );
  INV_X1 U16925 ( .A(n10980), .ZN(n21818) );
  NAND2_X1 U16926 ( .A1(n10980), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n21802) );
  INV_X1 U16927 ( .A(n21919), .ZN(n21925) );
  NAND2_X1 U16928 ( .A1(n21802), .A2(n21925), .ZN(n14910) );
  AOI21_X1 U16929 ( .B1(n21936), .B2(n21818), .A(n14910), .ZN(n14907) );
  AOI21_X1 U16930 ( .B1(n21938), .B2(n21580), .A(n14907), .ZN(n14909) );
  NAND2_X1 U16931 ( .A1(n21587), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n14908) );
  OAI21_X1 U16932 ( .B1(n21587), .B2(n14909), .A(n14908), .ZN(P1_U3477) );
  INV_X1 U16933 ( .A(n14910), .ZN(n15114) );
  NOR2_X1 U16934 ( .A1(n21802), .A2(n21919), .ZN(n15139) );
  MUX2_X1 U16935 ( .A(n15114), .B(n15139), .S(n14911), .Z(n14912) );
  AOI21_X1 U16936 ( .B1(n21580), .B2(n21821), .A(n14912), .ZN(n14914) );
  NAND2_X1 U16937 ( .A1(n21587), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14913) );
  OAI21_X1 U16938 ( .B1(n21587), .B2(n14914), .A(n14913), .ZN(P1_U3476) );
  OR2_X1 U16939 ( .A1(n14916), .A2(n14915), .ZN(n14917) );
  AND2_X1 U16940 ( .A1(n14881), .A2(n14917), .ZN(n19393) );
  INV_X1 U16941 ( .A(n19393), .ZN(n19455) );
  INV_X1 U16942 ( .A(n14918), .ZN(n14919) );
  OAI21_X1 U16943 ( .B1(n14921), .B2(n14920), .A(n14919), .ZN(n18277) );
  NOR2_X1 U16944 ( .A1(n18277), .A2(n16267), .ZN(n14922) );
  AOI21_X1 U16945 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n16267), .A(n14922), .ZN(
        n14923) );
  OAI21_X1 U16946 ( .B1(n19455), .B2(n16278), .A(n14923), .ZN(P2_U2883) );
  INV_X1 U16947 ( .A(n14924), .ZN(n14927) );
  AOI22_X1 U16948 ( .A1(n20015), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n21390), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n14925) );
  OAI21_X1 U16949 ( .B1(n20025), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n14925), .ZN(n14926) );
  AOI21_X1 U16950 ( .B1(n20020), .B2(n14927), .A(n14926), .ZN(n14928) );
  OAI21_X1 U16951 ( .B1(n19957), .B2(n21419), .A(n14928), .ZN(P1_U2998) );
  INV_X1 U16952 ( .A(n14929), .ZN(n14930) );
  AOI21_X1 U16953 ( .B1(n14931), .B2(n14882), .A(n14930), .ZN(n18297) );
  INV_X1 U16954 ( .A(n18297), .ZN(n17226) );
  NOR2_X1 U16955 ( .A1(n14881), .A2(n14932), .ZN(n14934) );
  OAI211_X1 U16956 ( .C1(n14934), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n16252), .B(n14933), .ZN(n14936) );
  NAND2_X1 U16957 ( .A1(n16267), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n14935) );
  OAI211_X1 U16958 ( .C1(n17226), .C2(n16267), .A(n14936), .B(n14935), .ZN(
        P2_U2881) );
  XNOR2_X1 U16959 ( .A(n14938), .B(n14937), .ZN(n14974) );
  AOI21_X1 U16960 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n15403) );
  INV_X1 U16961 ( .A(n15403), .ZN(n14958) );
  OAI22_X1 U16962 ( .A1(n21332), .A2(n14958), .B1(n21409), .B2(n15099), .ZN(
        n14941) );
  AND2_X1 U16963 ( .A1(n21390), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n14969) );
  NAND2_X1 U16964 ( .A1(n21337), .A2(n14939), .ZN(n16116) );
  NOR3_X1 U16965 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13533), .A3(
        n16116), .ZN(n14940) );
  NOR3_X1 U16966 ( .A1(n14941), .A2(n14969), .A3(n14940), .ZN(n14947) );
  INV_X1 U16967 ( .A(n21337), .ZN(n14943) );
  NAND2_X1 U16968 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14942) );
  OAI22_X1 U16969 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n14943), .B1(
        n14942), .B2(n21332), .ZN(n14945) );
  NAND2_X1 U16970 ( .A1(n21265), .A2(n21400), .ZN(n14944) );
  OAI21_X1 U16971 ( .B1(n14945), .B2(n21334), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n14946) );
  OAI211_X1 U16972 ( .C1(n14974), .C2(n21327), .A(n14947), .B(n14946), .ZN(
        P1_U3029) );
  NAND2_X1 U16973 ( .A1(n12618), .A2(n14948), .ZN(n14949) );
  INV_X1 U16974 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n21680) );
  INV_X1 U16975 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n14950) );
  OR2_X1 U16976 ( .A1(n15599), .A2(n14950), .ZN(n14952) );
  NAND2_X1 U16977 ( .A1(n15599), .A2(DATAI_0_), .ZN(n14951) );
  AND2_X1 U16978 ( .A1(n14952), .A2(n14951), .ZN(n21675) );
  OAI222_X1 U16979 ( .A1(n15890), .A2(n19955), .B1(n15886), .B2(n21680), .C1(
        n15885), .C2(n21675), .ZN(P1_U2904) );
  INV_X1 U16980 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n21691) );
  INV_X1 U16981 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n20032) );
  NOR2_X1 U16982 ( .A1(n15121), .A2(DATAI_2_), .ZN(n14953) );
  AOI21_X1 U16983 ( .B1(n15121), .B2(n20032), .A(n14953), .ZN(n15872) );
  INV_X1 U16984 ( .A(n15872), .ZN(n21686) );
  OAI222_X1 U16985 ( .A1(n15107), .A2(n15890), .B1(n15886), .B2(n21691), .C1(
        n15885), .C2(n21686), .ZN(P1_U2902) );
  INV_X1 U16986 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n21685) );
  INV_X1 U16987 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n20030) );
  NOR2_X1 U16988 ( .A1(n15121), .A2(DATAI_1_), .ZN(n14954) );
  AOI21_X1 U16989 ( .B1(n15121), .B2(n20030), .A(n14954), .ZN(n16177) );
  INV_X1 U16990 ( .A(n16177), .ZN(n21681) );
  OAI222_X1 U16991 ( .A1(n21419), .A2(n15890), .B1(n15886), .B2(n21685), .C1(
        n15885), .C2(n21681), .ZN(P1_U2903) );
  XNOR2_X1 U16992 ( .A(n14956), .B(n14955), .ZN(n15008) );
  NAND2_X1 U16993 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n21283) );
  AOI21_X1 U16994 ( .B1(n21283), .B2(n21337), .A(n21334), .ZN(n14957) );
  OAI21_X1 U16995 ( .B1(n21332), .B2(n14958), .A(n14957), .ZN(n14988) );
  NOR2_X1 U16996 ( .A1(n21283), .A2(n16116), .ZN(n21285) );
  AOI21_X1 U16997 ( .B1(n16041), .B2(n14958), .A(n21285), .ZN(n21295) );
  INV_X1 U16998 ( .A(n21295), .ZN(n14983) );
  AOI22_X1 U16999 ( .A1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n14988), .B1(
        n14983), .B2(n14959), .ZN(n14963) );
  OAI21_X1 U17000 ( .B1(n14836), .B2(n14960), .A(n14985), .ZN(n14980) );
  INV_X1 U17001 ( .A(n14980), .ZN(n15236) );
  INV_X1 U17002 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n14961) );
  NOR2_X1 U17003 ( .A1(n21378), .A2(n14961), .ZN(n15003) );
  AOI21_X1 U17004 ( .B1(n21394), .B2(n15236), .A(n15003), .ZN(n14962) );
  OAI211_X1 U17005 ( .C1(n21327), .C2(n15008), .A(n14963), .B(n14962), .ZN(
        P1_U3028) );
  XOR2_X1 U17006 ( .A(n14933), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .Z(n14968)
         );
  NAND2_X1 U17007 ( .A1(n14929), .A2(n14964), .ZN(n14965) );
  NAND2_X1 U17008 ( .A1(n14991), .A2(n14965), .ZN(n18303) );
  INV_X1 U17009 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n14966) );
  MUX2_X1 U17010 ( .A(n18303), .B(n14966), .S(n16267), .Z(n14967) );
  OAI21_X1 U17011 ( .B1(n14968), .B2(n16278), .A(n14967), .ZN(P2_U2880) );
  INV_X1 U17012 ( .A(n15107), .ZN(n14972) );
  AOI21_X1 U17013 ( .B1(n20015), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n14969), .ZN(n14970) );
  OAI21_X1 U17014 ( .B1(n20025), .B2(n15103), .A(n14970), .ZN(n14971) );
  AOI21_X1 U17015 ( .B1(n14972), .B2(n20021), .A(n14971), .ZN(n14973) );
  OAI21_X1 U17016 ( .B1(n21578), .B2(n14974), .A(n14973), .ZN(P1_U2997) );
  OAI21_X1 U17017 ( .B1(n14977), .B2(n14976), .A(n14975), .ZN(n15244) );
  INV_X1 U17018 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n19862) );
  INV_X1 U17019 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n20034) );
  NOR2_X1 U17020 ( .A1(n15121), .A2(DATAI_3_), .ZN(n14978) );
  AOI21_X1 U17021 ( .B1(n15121), .B2(n20034), .A(n14978), .ZN(n17209) );
  INV_X1 U17022 ( .A(n17209), .ZN(n14979) );
  OAI222_X1 U17023 ( .A1(n15244), .A2(n15890), .B1(n15886), .B2(n19862), .C1(
        n15885), .C2(n14979), .ZN(P1_U2901) );
  INV_X1 U17024 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n15234) );
  OAI222_X1 U17025 ( .A1(n15244), .A2(n15842), .B1(n15234), .B2(n19946), .C1(
        n14980), .C2(n15837), .ZN(P1_U2869) );
  XNOR2_X1 U17026 ( .A(n14982), .B(n14981), .ZN(n15015) );
  NAND2_X1 U17027 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n21284) );
  OAI211_X1 U17028 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n14983), .B(n21284), .ZN(n14990) );
  AND2_X1 U17029 ( .A1(n21390), .A2(P1_REIP_REG_4__SCAN_IN), .ZN(n15009) );
  NAND2_X1 U17030 ( .A1(n14985), .A2(n14984), .ZN(n14986) );
  NAND2_X1 U17031 ( .A1(n15083), .A2(n14986), .ZN(n21427) );
  NOR2_X1 U17032 ( .A1(n21409), .A2(n21427), .ZN(n14987) );
  AOI211_X1 U17033 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n14988), .A(
        n15009), .B(n14987), .ZN(n14989) );
  OAI211_X1 U17034 ( .C1(n15015), .C2(n21327), .A(n14990), .B(n14989), .ZN(
        P1_U3027) );
  AOI21_X1 U17035 ( .B1(n14992), .B2(n14991), .A(n15061), .ZN(n17236) );
  INV_X1 U17036 ( .A(n17236), .ZN(n18321) );
  OAI211_X1 U17037 ( .C1(n14995), .C2(n14994), .A(n14993), .B(n16252), .ZN(
        n14997) );
  NAND2_X1 U17038 ( .A1(n16267), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n14996) );
  OAI211_X1 U17039 ( .C1(n18321), .C2(n16267), .A(n14997), .B(n14996), .ZN(
        P2_U2879) );
  NAND2_X1 U17040 ( .A1(n14975), .A2(n14998), .ZN(n14999) );
  AND2_X1 U17041 ( .A1(n15079), .A2(n14999), .ZN(n21432) );
  INV_X1 U17042 ( .A(n21432), .ZN(n15002) );
  INV_X1 U17043 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n21700) );
  OR2_X1 U17044 ( .A1(n15599), .A2(n20036), .ZN(n15001) );
  NAND2_X1 U17045 ( .A1(n15599), .A2(DATAI_4_), .ZN(n15000) );
  NAND2_X1 U17046 ( .A1(n15001), .A2(n15000), .ZN(n15867) );
  INV_X1 U17047 ( .A(n15867), .ZN(n21695) );
  OAI222_X1 U17048 ( .A1(n15890), .A2(n15002), .B1(n15886), .B2(n21700), .C1(
        n15885), .C2(n21695), .ZN(P1_U2900) );
  INV_X1 U17049 ( .A(n15244), .ZN(n15006) );
  AOI21_X1 U17050 ( .B1(n20015), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n15003), .ZN(n15004) );
  OAI21_X1 U17051 ( .B1(n20025), .B2(n15240), .A(n15004), .ZN(n15005) );
  AOI21_X1 U17052 ( .B1(n15006), .B2(n20021), .A(n15005), .ZN(n15007) );
  OAI21_X1 U17053 ( .B1(n15008), .B2(n21578), .A(n15007), .ZN(P1_U2996) );
  INV_X1 U17054 ( .A(n21437), .ZN(n15012) );
  INV_X1 U17055 ( .A(n15009), .ZN(n15010) );
  OAI21_X1 U17056 ( .B1(n19983), .B2(n21428), .A(n15010), .ZN(n15011) );
  AOI21_X1 U17057 ( .B1(n15012), .B2(n20000), .A(n15011), .ZN(n15014) );
  NAND2_X1 U17058 ( .A1(n21432), .A2(n20021), .ZN(n15013) );
  OAI211_X1 U17059 ( .C1(n15015), .C2(n21578), .A(n15014), .B(n15013), .ZN(
        P1_U2995) );
  OAI22_X1 U17060 ( .A1(n15837), .A2(n21427), .B1(n15016), .B2(n19946), .ZN(
        n15017) );
  AOI21_X1 U17061 ( .B1(n21432), .B2(n19942), .A(n15017), .ZN(n15018) );
  INV_X1 U17062 ( .A(n15018), .ZN(P1_U2868) );
  INV_X1 U17063 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n21677) );
  AOI22_X1 U17064 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n19865), .B1(n19868), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n15019) );
  OAI21_X1 U17065 ( .B1(n21677), .B2(n15030), .A(n15019), .ZN(P1_U2920) );
  INV_X1 U17066 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n15021) );
  AOI22_X1 U17067 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n19868), .B1(n19865), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n15020) );
  OAI21_X1 U17068 ( .B1(n15021), .B2(n15030), .A(n15020), .ZN(P1_U2917) );
  AOI22_X1 U17069 ( .A1(n19868), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n15022) );
  OAI21_X1 U17070 ( .B1(n13042), .B2(n15030), .A(n15022), .ZN(P1_U2919) );
  AOI22_X1 U17071 ( .A1(n21257), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n15023) );
  OAI21_X1 U17072 ( .B1(n13231), .B2(n15030), .A(n15023), .ZN(P1_U2909) );
  INV_X1 U17073 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n21688) );
  AOI22_X1 U17074 ( .A1(n21257), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n15024) );
  OAI21_X1 U17075 ( .B1(n21688), .B2(n15030), .A(n15024), .ZN(P1_U2918) );
  INV_X1 U17076 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n21748) );
  AOI22_X1 U17077 ( .A1(n21257), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n15025) );
  OAI21_X1 U17078 ( .B1(n21748), .B2(n15030), .A(n15025), .ZN(P1_U2908) );
  INV_X1 U17079 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n21703) );
  AOI22_X1 U17080 ( .A1(n21257), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n15026) );
  OAI21_X1 U17081 ( .B1(n21703), .B2(n15030), .A(n15026), .ZN(P1_U2915) );
  INV_X1 U17082 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n21697) );
  AOI22_X1 U17083 ( .A1(n21257), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n15027) );
  OAI21_X1 U17084 ( .B1(n21697), .B2(n15030), .A(n15027), .ZN(P1_U2916) );
  INV_X1 U17085 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n21763) );
  AOI22_X1 U17086 ( .A1(n21257), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n15028) );
  OAI21_X1 U17087 ( .B1(n21763), .B2(n15030), .A(n15028), .ZN(P1_U2906) );
  INV_X1 U17088 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n21755) );
  AOI22_X1 U17089 ( .A1(n21257), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n15029) );
  OAI21_X1 U17090 ( .B1(n21755), .B2(n15030), .A(n15029), .ZN(P1_U2907) );
  NOR2_X1 U17091 ( .A1(n18361), .A2(n15066), .ZN(n15033) );
  XNOR2_X1 U17092 ( .A(n15033), .B(n15032), .ZN(n15034) );
  NAND2_X1 U17093 ( .A1(n15034), .A2(n18564), .ZN(n15043) );
  NAND2_X1 U17094 ( .A1(n19558), .A2(n18539), .ZN(n15038) );
  OAI22_X1 U17095 ( .A1(n15035), .A2(n18554), .B1(n14561), .B2(n18551), .ZN(
        n15036) );
  AOI21_X1 U17096 ( .B1(n18538), .B2(P2_EBX_REG_2__SCAN_IN), .A(n15036), .ZN(
        n15037) );
  OAI211_X1 U17097 ( .C1(n18552), .C2(n15039), .A(n15038), .B(n15037), .ZN(
        n15040) );
  AOI21_X1 U17098 ( .B1(n15041), .B2(n18560), .A(n15040), .ZN(n15042) );
  OAI211_X1 U17099 ( .C1(n15077), .C2(n19452), .A(n15043), .B(n15042), .ZN(
        P2_U2853) );
  NAND2_X1 U17100 ( .A1(n18562), .A2(n15044), .ZN(n15045) );
  XNOR2_X1 U17101 ( .A(n15295), .B(n15045), .ZN(n15046) );
  NAND2_X1 U17102 ( .A1(n15046), .A2(n18564), .ZN(n15057) );
  OR2_X1 U17103 ( .A1(n11066), .A2(n15048), .ZN(n15050) );
  NAND2_X1 U17104 ( .A1(n15050), .A2(n15049), .ZN(n19509) );
  OAI22_X1 U17105 ( .A1(n15051), .A2(n18552), .B1(n18567), .B2(n19509), .ZN(
        n15053) );
  NOR2_X1 U17106 ( .A1(n18557), .A2(n11503), .ZN(n15052) );
  AOI211_X1 U17107 ( .C1(n18524), .C2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n15053), .B(n15052), .ZN(n15054) );
  OAI21_X1 U17108 ( .B1(n15292), .B2(n18551), .A(n15054), .ZN(n15055) );
  AOI21_X1 U17109 ( .B1(n15047), .B2(n18560), .A(n15055), .ZN(n15056) );
  OAI211_X1 U17110 ( .C1(n15077), .C2(n19453), .A(n15057), .B(n15056), .ZN(
        P2_U2852) );
  OAI211_X1 U17111 ( .C1(n15058), .C2(n11385), .A(n16252), .B(n15224), .ZN(
        n15065) );
  NOR2_X1 U17112 ( .A1(n15061), .A2(n15060), .ZN(n15062) );
  OR2_X1 U17113 ( .A1(n15059), .A2(n15062), .ZN(n18331) );
  INV_X1 U17114 ( .A(n18331), .ZN(n15063) );
  NAND2_X1 U17115 ( .A1(n15063), .A2(n16209), .ZN(n15064) );
  OAI211_X1 U17116 ( .C1(n16209), .C2(n11575), .A(n15065), .B(n15064), .ZN(
        P2_U2878) );
  AOI211_X1 U17117 ( .C1(n18253), .C2(n15067), .A(n18361), .B(n15066), .ZN(
        n15283) );
  AOI22_X1 U17118 ( .A1(n15283), .A2(n18564), .B1(n15069), .B2(n15068), .ZN(
        n15076) );
  INV_X1 U17119 ( .A(n19449), .ZN(n19611) );
  AOI22_X1 U17120 ( .A1(n18536), .A2(P2_REIP_REG_1__SCAN_IN), .B1(n18539), 
        .B2(n19611), .ZN(n15071) );
  AOI22_X1 U17121 ( .A1(n18538), .A2(P2_EBX_REG_1__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18524), .ZN(n15070) );
  OAI211_X1 U17122 ( .C1(n18552), .C2(n15072), .A(n15071), .B(n15070), .ZN(
        n15073) );
  AOI21_X1 U17123 ( .B1(n15074), .B2(n18560), .A(n15073), .ZN(n15075) );
  OAI211_X1 U17124 ( .C1(n19448), .C2(n15077), .A(n15076), .B(n15075), .ZN(
        P2_U2854) );
  AND2_X1 U17125 ( .A1(n15079), .A2(n15078), .ZN(n15081) );
  OR2_X1 U17126 ( .A1(n15081), .A2(n15080), .ZN(n21449) );
  AND2_X1 U17127 ( .A1(n15083), .A2(n15082), .ZN(n15084) );
  NOR2_X1 U17128 ( .A1(n15088), .A2(n15084), .ZN(n21438) );
  AOI22_X1 U17129 ( .A1(n19941), .A2(n21438), .B1(P1_EBX_REG_5__SCAN_IN), .B2(
        n15840), .ZN(n15085) );
  OAI21_X1 U17130 ( .B1(n21449), .B2(n15842), .A(n15085), .ZN(P1_U2867) );
  OAI21_X1 U17131 ( .B1(n15080), .B2(n15087), .A(n15262), .ZN(n15256) );
  XOR2_X1 U17132 ( .A(n15089), .B(n15088), .Z(n21453) );
  AOI22_X1 U17133 ( .A1(n19941), .A2(n21453), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n15840), .ZN(n15090) );
  OAI21_X1 U17134 ( .B1(n15256), .B2(n15842), .A(n15090), .ZN(P1_U2866) );
  INV_X1 U17135 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n20038) );
  NOR2_X1 U17136 ( .A1(n15121), .A2(DATAI_5_), .ZN(n15091) );
  AOI21_X1 U17137 ( .B1(n15121), .B2(n20038), .A(n15091), .ZN(n15864) );
  INV_X1 U17138 ( .A(n15864), .ZN(n21701) );
  OAI222_X1 U17139 ( .A1(n21449), .A2(n15890), .B1(n15886), .B2(n12875), .C1(
        n15885), .C2(n21701), .ZN(P1_U2899) );
  NAND2_X1 U17140 ( .A1(n15093), .A2(n15092), .ZN(n15094) );
  NOR2_X1 U17141 ( .A1(n21459), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n21413) );
  OR2_X1 U17142 ( .A1(n21411), .A2(n21413), .ZN(n15230) );
  NOR2_X1 U17143 ( .A1(n15096), .A2(n15095), .ZN(n21423) );
  NAND2_X1 U17144 ( .A1(n21821), .A2(n21423), .ZN(n15098) );
  NOR2_X1 U17145 ( .A1(n21459), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n15231) );
  AOI22_X1 U17146 ( .A1(n15231), .A2(P1_REIP_REG_1__SCAN_IN), .B1(n21533), 
        .B2(P1_EBX_REG_2__SCAN_IN), .ZN(n15097) );
  OAI211_X1 U17147 ( .C1(n15099), .C2(n21562), .A(n15098), .B(n15097), .ZN(
        n15105) );
  NAND2_X1 U17148 ( .A1(n15100), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15101) );
  INV_X1 U17149 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n15102) );
  OAI22_X1 U17150 ( .A1(n15103), .A2(n21565), .B1(n21566), .B2(n15102), .ZN(
        n15104) );
  AOI211_X1 U17151 ( .C1(P1_REIP_REG_2__SCAN_IN), .C2(n15230), .A(n15105), .B(
        n15104), .ZN(n15106) );
  OAI21_X1 U17152 ( .B1(n21448), .B2(n15107), .A(n15106), .ZN(P1_U2838) );
  OAI22_X1 U17153 ( .A1(n21410), .A2(n21562), .B1(n21559), .B2(n13538), .ZN(
        n15109) );
  INV_X1 U17154 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n19950) );
  NOR2_X1 U17155 ( .A1(n21495), .A2(n19950), .ZN(n15108) );
  AOI211_X1 U17156 ( .C1(n21423), .C2(n21581), .A(n15109), .B(n15108), .ZN(
        n15111) );
  OAI21_X1 U17157 ( .B1(n21536), .B2(n21535), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n15110) );
  OAI211_X1 U17158 ( .C1(n21448), .C2(n19955), .A(n15111), .B(n15110), .ZN(
        P1_U2840) );
  OR2_X1 U17159 ( .A1(n21933), .A2(n21932), .ZN(n15125) );
  NOR2_X1 U17160 ( .A1(n21914), .A2(n21919), .ZN(n15113) );
  AOI211_X1 U17161 ( .C1(n15125), .C2(n21919), .A(n15114), .B(n15113), .ZN(
        n15120) );
  NAND2_X1 U17162 ( .A1(n21821), .A2(n15115), .ZN(n21931) );
  AND2_X1 U17163 ( .A1(n15116), .A2(n21581), .ZN(n21853) );
  INV_X1 U17164 ( .A(n21853), .ZN(n15118) );
  NAND2_X1 U17165 ( .A1(n15117), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n16176) );
  OAI21_X1 U17166 ( .B1(n21931), .B2(n15118), .A(n16176), .ZN(n15119) );
  AND2_X1 U17167 ( .A1(n15119), .A2(n21876), .ZN(n15128) );
  OAI21_X1 U17168 ( .B1(n15120), .B2(n15128), .A(n21923), .ZN(n22202) );
  INV_X1 U17169 ( .A(n22202), .ZN(n15135) );
  INV_X1 U17170 ( .A(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15134) );
  INV_X1 U17171 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n20073) );
  INV_X1 U17172 ( .A(DATAI_24_), .ZN(n17105) );
  NAND2_X1 U17173 ( .A1(n20021), .A2(n15599), .ZN(n22150) );
  OAI22_X2 U17174 ( .A1(n20073), .A2(n22152), .B1(n17105), .B2(n22150), .ZN(
        n21944) );
  INV_X1 U17175 ( .A(n22305), .ZN(n16191) );
  INV_X1 U17176 ( .A(n15122), .ZN(n15123) );
  INV_X1 U17177 ( .A(n16175), .ZN(n22149) );
  NAND2_X1 U17178 ( .A1(n22149), .A2(n15124), .ZN(n21880) );
  INV_X1 U17179 ( .A(n15125), .ZN(n15126) );
  AND2_X1 U17180 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n15126), .ZN(n15127) );
  OR2_X1 U17181 ( .A1(n15128), .A2(n15127), .ZN(n22199) );
  NAND2_X1 U17182 ( .A1(n21935), .A2(n22199), .ZN(n15131) );
  INV_X1 U17183 ( .A(DATAI_16_), .ZN(n17125) );
  INV_X1 U17184 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n20058) );
  OAI22_X1 U17185 ( .A1(n17125), .A2(n22150), .B1(n20058), .B2(n22152), .ZN(
        n21901) );
  NAND2_X1 U17186 ( .A1(n22207), .A2(n21901), .ZN(n15130) );
  OAI211_X1 U17187 ( .C1(n16176), .C2(n21880), .A(n15131), .B(n15130), .ZN(
        n15132) );
  AOI21_X1 U17188 ( .B1(n21944), .B2(n16191), .A(n15132), .ZN(n15133) );
  OAI21_X1 U17189 ( .B1(n15135), .B2(n15134), .A(n15133), .ZN(P1_U3153) );
  INV_X1 U17190 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n21711) );
  OR2_X1 U17191 ( .A1(n15599), .A2(n20040), .ZN(n15137) );
  NAND2_X1 U17192 ( .A1(n15599), .A2(DATAI_6_), .ZN(n15136) );
  NAND2_X1 U17193 ( .A1(n15137), .A2(n15136), .ZN(n22144) );
  INV_X1 U17194 ( .A(n22144), .ZN(n21706) );
  OAI222_X1 U17195 ( .A1(n15256), .A2(n15890), .B1(n21711), .B2(n15886), .C1(
        n15885), .C2(n21706), .ZN(P1_U2898) );
  INV_X1 U17196 ( .A(n14911), .ZN(n15138) );
  AND2_X1 U17197 ( .A1(n21870), .A2(n15139), .ZN(n15140) );
  NOR3_X1 U17198 ( .A1(n21933), .A2(n21794), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21879) );
  OAI21_X1 U17199 ( .B1(n15140), .B2(n21879), .A(n21923), .ZN(n22185) );
  INV_X1 U17200 ( .A(n22185), .ZN(n15251) );
  INV_X1 U17201 ( .A(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n15150) );
  INV_X1 U17202 ( .A(n22273), .ZN(n15248) );
  INV_X1 U17203 ( .A(n21901), .ZN(n21947) );
  AND2_X1 U17204 ( .A1(n21771), .A2(n14715), .ZN(n21884) );
  NAND2_X1 U17205 ( .A1(n21884), .A2(n21853), .ZN(n15143) );
  INV_X1 U17206 ( .A(n21879), .ZN(n15141) );
  NOR2_X1 U17207 ( .A1(n21915), .A2(n15141), .ZN(n22183) );
  INV_X1 U17208 ( .A(n22183), .ZN(n15142) );
  NAND2_X1 U17209 ( .A1(n15143), .A2(n15142), .ZN(n15144) );
  NAND2_X1 U17210 ( .A1(n15144), .A2(n21925), .ZN(n15146) );
  NAND2_X1 U17211 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21879), .ZN(n15145) );
  NAND2_X1 U17212 ( .A1(n15146), .A2(n15145), .ZN(n22184) );
  AOI22_X1 U17213 ( .A1(n21935), .A2(n22184), .B1(n21934), .B2(n22183), .ZN(
        n15147) );
  OAI21_X1 U17214 ( .B1(n21910), .B2(n21947), .A(n15147), .ZN(n15148) );
  AOI21_X1 U17215 ( .B1(n21944), .B2(n15248), .A(n15148), .ZN(n15149) );
  OAI21_X1 U17216 ( .B1(n15251), .B2(n15150), .A(n15149), .ZN(P1_U3121) );
  INV_X1 U17217 ( .A(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15155) );
  INV_X1 U17218 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n20077) );
  INV_X1 U17219 ( .A(DATAI_26_), .ZN(n17107) );
  OAI22_X2 U17220 ( .A1(n20077), .A2(n22152), .B1(n17107), .B2(n22150), .ZN(
        n22024) );
  INV_X1 U17221 ( .A(DATAI_18_), .ZN(n16994) );
  INV_X1 U17222 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n20062) );
  OAI22_X1 U17223 ( .A1(n16994), .A2(n22150), .B1(n20062), .B2(n22152), .ZN(
        n22016) );
  INV_X1 U17224 ( .A(n22016), .ZN(n22027) );
  NOR2_X2 U17225 ( .A1(n16175), .A2(n15151), .ZN(n22023) );
  NAND2_X1 U17226 ( .A1(n22145), .A2(n15872), .ZN(n22019) );
  AOI22_X1 U17227 ( .A1(n22023), .A2(n22183), .B1(n22022), .B2(n22184), .ZN(
        n15152) );
  OAI21_X1 U17228 ( .B1(n21910), .B2(n22027), .A(n15152), .ZN(n15153) );
  AOI21_X1 U17229 ( .B1(n22024), .B2(n15248), .A(n15153), .ZN(n15154) );
  OAI21_X1 U17230 ( .B1(n15251), .B2(n15155), .A(n15154), .ZN(P1_U3123) );
  INV_X1 U17231 ( .A(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15160) );
  INV_X1 U17232 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n20084) );
  INV_X1 U17233 ( .A(DATAI_29_), .ZN(n17118) );
  INV_X1 U17234 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n20068) );
  INV_X1 U17235 ( .A(DATAI_21_), .ZN(n16999) );
  OAI22_X1 U17236 ( .A1(n20068), .A2(n22152), .B1(n16999), .B2(n22150), .ZN(
        n22132) );
  INV_X1 U17237 ( .A(n22132), .ZN(n22143) );
  NOR2_X2 U17238 ( .A1(n16175), .A2(n15156), .ZN(n22139) );
  NAND2_X1 U17239 ( .A1(n22145), .A2(n15864), .ZN(n22135) );
  AOI22_X1 U17240 ( .A1(n22139), .A2(n22183), .B1(n22138), .B2(n22184), .ZN(
        n15157) );
  OAI21_X1 U17241 ( .B1(n21910), .B2(n22143), .A(n15157), .ZN(n15158) );
  AOI21_X1 U17242 ( .B1(n22140), .B2(n15248), .A(n15158), .ZN(n15159) );
  OAI21_X1 U17243 ( .B1(n15251), .B2(n15160), .A(n15159), .ZN(P1_U3126) );
  INV_X1 U17244 ( .A(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15166) );
  INV_X1 U17245 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n20080) );
  INV_X1 U17246 ( .A(DATAI_27_), .ZN(n17104) );
  OAI22_X2 U17247 ( .A1(n20080), .A2(n22152), .B1(n17104), .B2(n22150), .ZN(
        n22062) );
  INV_X1 U17248 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n20064) );
  INV_X1 U17249 ( .A(DATAI_19_), .ZN(n15161) );
  OAI22_X1 U17250 ( .A1(n20064), .A2(n22152), .B1(n15161), .B2(n22150), .ZN(
        n22054) );
  INV_X1 U17251 ( .A(n22054), .ZN(n22065) );
  NOR2_X2 U17252 ( .A1(n16175), .A2(n15162), .ZN(n22061) );
  NAND2_X1 U17253 ( .A1(n22145), .A2(n17209), .ZN(n22057) );
  AOI22_X1 U17254 ( .A1(n22061), .A2(n22183), .B1(n22060), .B2(n22184), .ZN(
        n15163) );
  OAI21_X1 U17255 ( .B1(n21910), .B2(n22065), .A(n15163), .ZN(n15164) );
  AOI21_X1 U17256 ( .B1(n22062), .B2(n15248), .A(n15164), .ZN(n15165) );
  OAI21_X1 U17257 ( .B1(n15251), .B2(n15166), .A(n15165), .ZN(P1_U3124) );
  INV_X1 U17258 ( .A(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15173) );
  INV_X1 U17259 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n20087) );
  OAI22_X1 U17260 ( .A1(n15167), .A2(n22150), .B1(n20087), .B2(n22152), .ZN(
        n22300) );
  INV_X1 U17261 ( .A(DATAI_23_), .ZN(n17108) );
  INV_X1 U17262 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n20071) );
  OAI22_X1 U17263 ( .A1(n17108), .A2(n22150), .B1(n20071), .B2(n22152), .ZN(
        n22282) );
  INV_X1 U17264 ( .A(n22282), .ZN(n22306) );
  INV_X1 U17265 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n20042) );
  OR2_X1 U17266 ( .A1(n15599), .A2(n20042), .ZN(n15169) );
  NAND2_X1 U17267 ( .A1(n15599), .A2(DATAI_7_), .ZN(n15168) );
  NAND2_X1 U17268 ( .A1(n15169), .A2(n15168), .ZN(n15858) );
  NOR2_X2 U17269 ( .A1(n16175), .A2(n15597), .ZN(n22297) );
  AOI22_X1 U17270 ( .A1(n22299), .A2(n22184), .B1(n22297), .B2(n22183), .ZN(
        n15170) );
  OAI21_X1 U17271 ( .B1(n21910), .B2(n22306), .A(n15170), .ZN(n15171) );
  AOI21_X1 U17272 ( .B1(n22300), .B2(n15248), .A(n15171), .ZN(n15172) );
  OAI21_X1 U17273 ( .B1(n15251), .B2(n15173), .A(n15172), .ZN(P1_U3128) );
  OR2_X1 U17274 ( .A1(n18258), .A2(n16880), .ZN(n15180) );
  INV_X1 U17275 ( .A(n12241), .ZN(n15178) );
  INV_X1 U17276 ( .A(n12244), .ZN(n15175) );
  NAND2_X1 U17277 ( .A1(n15175), .A2(n15174), .ZN(n15279) );
  INV_X1 U17278 ( .A(n15279), .ZN(n15177) );
  MUX2_X1 U17279 ( .A(n15178), .B(n15177), .S(n15176), .Z(n15179) );
  NAND2_X1 U17280 ( .A1(n15180), .A2(n15179), .ZN(n18613) );
  INV_X1 U17281 ( .A(n15181), .ZN(n15182) );
  INV_X1 U17282 ( .A(n18668), .ZN(n15333) );
  AOI22_X1 U17283 ( .A1(n18361), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n18253), .B2(n18562), .ZN(n15284) );
  AOI222_X1 U17284 ( .A1(n18613), .A2(n15334), .B1(n15182), .B2(n15333), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n15284), .ZN(n15184) );
  NAND2_X1 U17285 ( .A1(n16897), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15183) );
  OAI21_X1 U17286 ( .B1(n15184), .B2(n16897), .A(n15183), .ZN(P2_U3601) );
  INV_X1 U17287 ( .A(n22300), .ZN(n22280) );
  NAND2_X1 U17288 ( .A1(n22202), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n15188) );
  INV_X1 U17289 ( .A(n22299), .ZN(n22287) );
  INV_X1 U17290 ( .A(n22199), .ZN(n15185) );
  INV_X1 U17291 ( .A(n22297), .ZN(n22272) );
  OAI22_X1 U17292 ( .A1(n22287), .A2(n15185), .B1(n16176), .B2(n22272), .ZN(
        n15186) );
  AOI21_X1 U17293 ( .B1(n22207), .B2(n22282), .A(n15186), .ZN(n15187) );
  OAI211_X1 U17294 ( .C1(n22305), .C2(n22280), .A(n15188), .B(n15187), .ZN(
        P1_U3160) );
  OR2_X1 U17295 ( .A1(n19447), .A2(n21607), .ZN(n19197) );
  OAI21_X1 U17296 ( .B1(n19256), .B2(n19197), .A(n19295), .ZN(n15205) );
  NAND2_X1 U17297 ( .A1(n19213), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19266) );
  INV_X1 U17298 ( .A(n19266), .ZN(n19269) );
  NAND2_X1 U17299 ( .A1(n19269), .A2(n19294), .ZN(n19279) );
  INV_X1 U17300 ( .A(n19279), .ZN(n15189) );
  OR2_X1 U17301 ( .A1(n15205), .A2(n15189), .ZN(n15194) );
  NAND2_X1 U17302 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n18669), .ZN(n18246) );
  NAND2_X1 U17303 ( .A1(n18652), .A2(n18246), .ZN(n18667) );
  NAND2_X1 U17304 ( .A1(n15190), .A2(n18667), .ZN(n15191) );
  NAND2_X1 U17305 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19294), .ZN(
        n19324) );
  NOR2_X1 U17306 ( .A1(n19324), .A2(n19266), .ZN(n19753) );
  INV_X1 U17307 ( .A(n19753), .ZN(n15201) );
  NOR2_X1 U17308 ( .A1(n15191), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19331) );
  NAND2_X1 U17309 ( .A1(n15203), .A2(n19331), .ZN(n15192) );
  OAI211_X1 U17310 ( .C1(n19683), .C2(n15201), .A(n15192), .B(n19332), .ZN(
        n15193) );
  NAND2_X1 U17311 ( .A1(n15194), .A2(n15193), .ZN(n19755) );
  INV_X1 U17312 ( .A(n19755), .ZN(n19376) );
  INV_X1 U17313 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15209) );
  NOR3_X4 U17314 ( .A1(n21607), .A2(n15195), .A3(n19332), .ZN(n19690) );
  NOR3_X4 U17315 ( .A1(n15196), .A2(n21607), .A3(n19332), .ZN(n19689) );
  AOI22_X1 U17316 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19690), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19689), .ZN(n19341) );
  INV_X1 U17317 ( .A(n19341), .ZN(n19319) );
  INV_X1 U17318 ( .A(n19256), .ZN(n15198) );
  INV_X1 U17319 ( .A(n19195), .ZN(n15197) );
  INV_X1 U17320 ( .A(n19690), .ZN(n19464) );
  INV_X1 U17321 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n20706) );
  INV_X1 U17322 ( .A(n19689), .ZN(n19462) );
  OAI22_X2 U17323 ( .A1(n20071), .A2(n19464), .B1(n20706), .B2(n19462), .ZN(
        n19338) );
  INV_X1 U17324 ( .A(n19338), .ZN(n15394) );
  INV_X1 U17325 ( .A(n19685), .ZN(n15199) );
  NAND2_X1 U17326 ( .A1(n15200), .A2(n15199), .ZN(n15392) );
  OAI22_X1 U17327 ( .A1(n15394), .A2(n19758), .B1(n15392), .B2(n15201), .ZN(
        n15202) );
  AOI21_X1 U17328 ( .B1(n19319), .B2(n19760), .A(n15202), .ZN(n15208) );
  OAI21_X1 U17329 ( .B1(n15203), .B2(n19753), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15204) );
  OAI21_X1 U17330 ( .B1(n15205), .B2(n19279), .A(n15204), .ZN(n19754) );
  NAND2_X1 U17331 ( .A1(n19754), .A2(n15206), .ZN(n15207) );
  OAI211_X1 U17332 ( .C1(n19376), .C2(n15209), .A(n15208), .B(n15207), .ZN(
        P2_U3095) );
  OR2_X1 U17333 ( .A1(n19559), .A2(n19197), .ZN(n19329) );
  OAI21_X1 U17334 ( .B1(n19453), .B2(n19329), .A(n19295), .ZN(n15218) );
  NAND3_X1 U17335 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19294), .A3(
        n19221), .ZN(n19242) );
  INV_X1 U17336 ( .A(n19242), .ZN(n15210) );
  OR2_X1 U17337 ( .A1(n15218), .A2(n15210), .ZN(n15214) );
  NAND2_X1 U17338 ( .A1(n11833), .A2(n19331), .ZN(n15212) );
  NOR2_X1 U17339 ( .A1(n19263), .A2(n19242), .ZN(n19726) );
  OAI21_X1 U17340 ( .B1(n19295), .B2(n19726), .A(n19312), .ZN(n15211) );
  NAND2_X1 U17341 ( .A1(n15212), .A2(n15211), .ZN(n15213) );
  INV_X1 U17342 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15221) );
  INV_X1 U17343 ( .A(n19727), .ZN(n19229) );
  INV_X1 U17344 ( .A(n19726), .ZN(n15215) );
  OAI22_X1 U17345 ( .A1(n15394), .A2(n19229), .B1(n15392), .B2(n15215), .ZN(
        n15216) );
  AOI21_X1 U17346 ( .B1(n19319), .B2(n19734), .A(n15216), .ZN(n15220) );
  OAI21_X1 U17347 ( .B1(n11833), .B2(n19726), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15217) );
  OAI21_X1 U17348 ( .B1(n15218), .B2(n19242), .A(n15217), .ZN(n19728) );
  NAND2_X1 U17349 ( .A1(n19728), .A2(n15206), .ZN(n15219) );
  OAI211_X1 U17350 ( .C1(n19732), .C2(n15221), .A(n15220), .B(n15219), .ZN(
        P2_U3127) );
  OR2_X1 U17351 ( .A1(n15059), .A2(n15222), .ZN(n15223) );
  AND2_X1 U17352 ( .A1(n15223), .A2(n11057), .ZN(n18341) );
  INV_X1 U17353 ( .A(n18341), .ZN(n15228) );
  INV_X1 U17354 ( .A(n15224), .ZN(n15225) );
  OAI211_X1 U17355 ( .C1(n15225), .C2(n10995), .A(n11363), .B(n16252), .ZN(
        n15227) );
  NAND2_X1 U17356 ( .A1(n16267), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n15226) );
  OAI211_X1 U17357 ( .C1(n15228), .C2(n16267), .A(n15227), .B(n15226), .ZN(
        P2_U2877) );
  INV_X1 U17358 ( .A(n21423), .ZN(n15238) );
  INV_X1 U17359 ( .A(n21433), .ZN(n15229) );
  NAND3_X1 U17360 ( .A1(n21483), .A2(n14961), .A3(n15229), .ZN(n15233) );
  OAI21_X1 U17361 ( .B1(n15231), .B2(n15230), .A(P1_REIP_REG_3__SCAN_IN), .ZN(
        n15232) );
  OAI211_X1 U17362 ( .C1(n15234), .C2(n21559), .A(n15233), .B(n15232), .ZN(
        n15235) );
  AOI21_X1 U17363 ( .B1(n15236), .B2(n21469), .A(n15235), .ZN(n15237) );
  OAI21_X1 U17364 ( .B1(n15239), .B2(n15238), .A(n15237), .ZN(n15242) );
  NOR2_X1 U17365 ( .A1(n21565), .A2(n15240), .ZN(n15241) );
  AOI211_X1 U17366 ( .C1(n21536), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n15242), .B(n15241), .ZN(n15243) );
  OAI21_X1 U17367 ( .B1(n21448), .B2(n15244), .A(n15243), .ZN(P1_U2837) );
  INV_X1 U17368 ( .A(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15250) );
  INV_X1 U17369 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n20082) );
  INV_X1 U17370 ( .A(DATAI_28_), .ZN(n17101) );
  INV_X1 U17371 ( .A(DATAI_20_), .ZN(n17120) );
  INV_X1 U17372 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n20066) );
  OAI22_X1 U17373 ( .A1(n17120), .A2(n22150), .B1(n20066), .B2(n22152), .ZN(
        n22102) );
  INV_X1 U17374 ( .A(n22102), .ZN(n22099) );
  NOR2_X2 U17375 ( .A1(n16175), .A2(n15245), .ZN(n22100) );
  AOI22_X1 U17376 ( .A1(n22101), .A2(n22184), .B1(n22183), .B2(n22100), .ZN(
        n15246) );
  OAI21_X1 U17377 ( .B1(n21910), .B2(n22099), .A(n15246), .ZN(n15247) );
  AOI21_X1 U17378 ( .B1(n22096), .B2(n15248), .A(n15247), .ZN(n15249) );
  OAI21_X1 U17379 ( .B1(n15251), .B2(n15250), .A(n15249), .ZN(P1_U3125) );
  NAND2_X1 U17380 ( .A1(n15253), .A2(n15252), .ZN(n15254) );
  NAND2_X1 U17381 ( .A1(n15255), .A2(n15254), .ZN(n21287) );
  INV_X1 U17382 ( .A(n15256), .ZN(n21457) );
  INV_X1 U17383 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n19886) );
  NOR2_X1 U17384 ( .A1(n21378), .A2(n19886), .ZN(n21289) );
  AOI21_X1 U17385 ( .B1(n20015), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n21289), .ZN(n15257) );
  OAI21_X1 U17386 ( .B1(n20025), .B2(n21463), .A(n15257), .ZN(n15258) );
  AOI21_X1 U17387 ( .B1(n21457), .B2(n20021), .A(n15258), .ZN(n15259) );
  OAI21_X1 U17388 ( .B1(n21287), .B2(n21578), .A(n15259), .ZN(P1_U2993) );
  NAND2_X1 U17389 ( .A1(n15262), .A2(n15261), .ZN(n15263) );
  AND2_X1 U17390 ( .A1(n15260), .A2(n15263), .ZN(n21475) );
  INV_X1 U17391 ( .A(n21475), .ZN(n15278) );
  INV_X1 U17392 ( .A(n15858), .ZN(n21712) );
  OAI222_X1 U17393 ( .A1(n15278), .A2(n15890), .B1(n15264), .B2(n15886), .C1(
        n15885), .C2(n21712), .ZN(P1_U2897) );
  INV_X1 U17394 ( .A(n15265), .ZN(n15266) );
  OAI211_X1 U17395 ( .C1(n15268), .C2(n15267), .A(n15266), .B(n16252), .ZN(
        n15274) );
  NAND2_X1 U17396 ( .A1(n15269), .A2(n11057), .ZN(n15272) );
  INV_X1 U17397 ( .A(n15270), .ZN(n15271) );
  NAND2_X1 U17398 ( .A1(n16209), .A2(n18352), .ZN(n15273) );
  OAI211_X1 U17399 ( .C1(n16209), .C2(n11576), .A(n15274), .B(n15273), .ZN(
        P2_U2876) );
  OR2_X1 U17400 ( .A1(n15276), .A2(n15275), .ZN(n15277) );
  NAND2_X1 U17401 ( .A1(n15399), .A2(n15277), .ZN(n21464) );
  INV_X1 U17402 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n21467) );
  OAI222_X1 U17403 ( .A1(n21464), .A2(n15837), .B1(n21467), .B2(n19946), .C1(
        n15278), .C2(n15842), .ZN(P1_U2865) );
  OAI21_X1 U17404 ( .B1(n11411), .B2(n15280), .A(n15279), .ZN(n15282) );
  NAND2_X1 U17405 ( .A1(n12241), .A2(n11358), .ZN(n15281) );
  OAI211_X1 U17406 ( .C1(n11771), .C2(n16880), .A(n15282), .B(n15281), .ZN(
        n18617) );
  AOI21_X1 U17407 ( .B1(n18361), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n15283), .ZN(n15330) );
  NOR2_X1 U17408 ( .A1(n15284), .A2(n17266), .ZN(n15331) );
  AOI222_X1 U17409 ( .A1(n18617), .A2(n15334), .B1(n15330), .B2(n15331), .C1(
        n19447), .C2(n15333), .ZN(n15286) );
  NAND2_X1 U17410 ( .A1(n16897), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n15285) );
  OAI21_X1 U17411 ( .B1(n15286), .B2(n16897), .A(n15285), .ZN(P2_U3600) );
  XNOR2_X1 U17412 ( .A(n15288), .B(n15289), .ZN(n15358) );
  XNOR2_X1 U17413 ( .A(n15358), .B(n15357), .ZN(n15316) );
  XOR2_X1 U17414 ( .A(n15290), .B(n15291), .Z(n15313) );
  OAI22_X1 U17415 ( .A1(n17222), .A2(n15293), .B1(n15292), .B2(n18582), .ZN(
        n15294) );
  AOI21_X1 U17416 ( .B1(n17216), .B2(n15295), .A(n15294), .ZN(n15296) );
  AOI21_X1 U17417 ( .B1(n15313), .B2(n17256), .A(n15297), .ZN(n15298) );
  OAI21_X1 U17418 ( .B1(n15316), .B2(n17228), .A(n15298), .ZN(P2_U3011) );
  OR2_X1 U17419 ( .A1(n15299), .A2(n15270), .ZN(n15300) );
  NAND2_X1 U17420 ( .A1(n15300), .A2(n14487), .ZN(n18367) );
  NAND2_X1 U17421 ( .A1(n15265), .A2(n15301), .ZN(n15337) );
  OAI211_X1 U17422 ( .C1(n15265), .C2(n15301), .A(n15337), .B(n16252), .ZN(
        n15303) );
  NAND2_X1 U17423 ( .A1(n16267), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n15302) );
  OAI211_X1 U17424 ( .C1(n18367), .C2(n16267), .A(n15303), .B(n15302), .ZN(
        P2_U2875) );
  AND2_X1 U17425 ( .A1(n16833), .A2(n15304), .ZN(n15310) );
  AOI211_X1 U17426 ( .C1(n15308), .C2(n15307), .A(n15306), .B(n15305), .ZN(
        n15372) );
  INV_X1 U17427 ( .A(n15372), .ZN(n15309) );
  MUX2_X1 U17428 ( .A(n15310), .B(n15309), .S(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n15312) );
  OAI22_X1 U17429 ( .A1(n19509), .A2(n16871), .B1(n15292), .B2(n18583), .ZN(
        n15311) );
  AOI211_X1 U17430 ( .C1(n18603), .C2(n15047), .A(n15312), .B(n15311), .ZN(
        n15315) );
  NAND2_X1 U17431 ( .A1(n15313), .A2(n16864), .ZN(n15314) );
  OAI211_X1 U17432 ( .C1(n15316), .C2(n18575), .A(n15315), .B(n15314), .ZN(
        P2_U3043) );
  INV_X1 U17433 ( .A(n18636), .ZN(n15318) );
  NAND2_X1 U17434 ( .A1(n15318), .A2(n15317), .ZN(n16887) );
  INV_X1 U17435 ( .A(n15319), .ZN(n16882) );
  INV_X1 U17436 ( .A(n11413), .ZN(n15320) );
  NAND2_X1 U17437 ( .A1(n15320), .A2(n11454), .ZN(n16886) );
  NAND2_X1 U17438 ( .A1(n16882), .A2(n16886), .ZN(n15325) );
  NOR2_X1 U17439 ( .A1(n15321), .A2(n15322), .ZN(n15323) );
  AOI22_X1 U17440 ( .A1(n16887), .A2(n15325), .B1(n12241), .B2(n15323), .ZN(
        n15328) );
  NAND2_X1 U17441 ( .A1(n11722), .A2(n15324), .ZN(n16883) );
  INV_X1 U17442 ( .A(n15325), .ZN(n15326) );
  NAND2_X1 U17443 ( .A1(n16883), .A2(n15326), .ZN(n15327) );
  OAI211_X1 U17444 ( .C1(n15329), .C2(n16880), .A(n15328), .B(n15327), .ZN(
        n18610) );
  INV_X1 U17445 ( .A(n15330), .ZN(n15332) );
  AOI222_X1 U17446 ( .A1(n18610), .A2(n15334), .B1(n15333), .B2(n19559), .C1(
        n15332), .C2(n15331), .ZN(n15336) );
  NAND2_X1 U17447 ( .A1(n16897), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15335) );
  OAI21_X1 U17448 ( .B1(n15336), .B2(n16897), .A(n15335), .ZN(P2_U3599) );
  INV_X1 U17449 ( .A(n15337), .ZN(n15340) );
  NAND2_X1 U17450 ( .A1(n15265), .A2(n15338), .ZN(n15494) );
  OAI211_X1 U17451 ( .C1(n15340), .C2(n15339), .A(n16252), .B(n15494), .ZN(
        n15342) );
  INV_X1 U17452 ( .A(n16559), .ZN(n16770) );
  NAND2_X1 U17453 ( .A1(n16209), .A2(n16770), .ZN(n15341) );
  OAI211_X1 U17454 ( .C1(n16209), .C2(n15343), .A(n15342), .B(n15341), .ZN(
        P2_U2874) );
  NAND2_X1 U17455 ( .A1(n19447), .A2(n18260), .ZN(n19276) );
  OAI21_X1 U17456 ( .B1(n19789), .B2(n19794), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n15344) );
  NAND2_X1 U17457 ( .A1(n15344), .A2(n19292), .ZN(n15353) );
  INV_X1 U17458 ( .A(n15345), .ZN(n19687) );
  INV_X1 U17459 ( .A(n19331), .ZN(n19297) );
  OAI21_X1 U17460 ( .B1(n11823), .B2(n19297), .A(n19332), .ZN(n15346) );
  OAI21_X1 U17461 ( .B1(n15353), .B2(n19687), .A(n15346), .ZN(n15347) );
  NAND2_X1 U17462 ( .A1(n19221), .A2(n19213), .ZN(n19323) );
  NOR2_X1 U17463 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19323), .ZN(
        n19336) );
  INV_X1 U17464 ( .A(n19336), .ZN(n19327) );
  NOR2_X1 U17465 ( .A1(n19327), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19788) );
  INV_X1 U17466 ( .A(n19788), .ZN(n15348) );
  OAI22_X1 U17467 ( .A1(n15394), .A2(n19785), .B1(n15392), .B2(n15348), .ZN(
        n15349) );
  AOI21_X1 U17468 ( .B1(n19789), .B2(n19319), .A(n15349), .ZN(n15355) );
  NOR2_X1 U17469 ( .A1(n19687), .A2(n19788), .ZN(n15352) );
  INV_X1 U17470 ( .A(n11823), .ZN(n15350) );
  OAI21_X1 U17471 ( .B1(n15350), .B2(n19788), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15351) );
  NAND2_X1 U17472 ( .A1(n19792), .A2(n15206), .ZN(n15354) );
  OAI211_X1 U17473 ( .C1(n19798), .C2(n15356), .A(n15355), .B(n15354), .ZN(
        P2_U3055) );
  AOI22_X1 U17474 ( .A1(n15358), .A2(n15357), .B1(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n15288), .ZN(n15360) );
  XNOR2_X1 U17475 ( .A(n18267), .B(n15479), .ZN(n15359) );
  XNOR2_X1 U17476 ( .A(n15360), .B(n15359), .ZN(n15382) );
  OAI21_X1 U17477 ( .B1(n15362), .B2(n15479), .A(n15361), .ZN(n15380) );
  OAI22_X1 U17478 ( .A1(n12132), .A2(n18582), .B1(n17261), .B2(n18270), .ZN(
        n15363) );
  AOI21_X1 U17479 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17245), .A(
        n15363), .ZN(n15364) );
  OAI21_X1 U17480 ( .B1(n17227), .B2(n18277), .A(n15364), .ZN(n15365) );
  AOI21_X1 U17481 ( .B1(n15380), .B2(n17256), .A(n15365), .ZN(n15366) );
  OAI21_X1 U17482 ( .B1(n15382), .B2(n17228), .A(n15366), .ZN(P2_U3010) );
  AND2_X1 U17483 ( .A1(n15260), .A2(n15367), .ZN(n15369) );
  OR2_X1 U17484 ( .A1(n15369), .A2(n15368), .ZN(n21488) );
  MUX2_X1 U17485 ( .A(BUF1_REG_8__SCAN_IN), .B(DATAI_8_), .S(n15599), .Z(
        n21717) );
  AOI22_X1 U17486 ( .A1(n15888), .A2(n21717), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n15887), .ZN(n15370) );
  OAI21_X1 U17487 ( .B1(n21488), .B2(n15890), .A(n15370), .ZN(P1_U2896) );
  NAND2_X1 U17488 ( .A1(n15371), .A2(n16833), .ZN(n15477) );
  OAI21_X1 U17489 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n16764), .A(
        n15372), .ZN(n15482) );
  INV_X1 U17490 ( .A(n15482), .ZN(n15374) );
  NAND2_X1 U17491 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n18382), .ZN(n15373) );
  OAI221_X1 U17492 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n15477), .C1(
        n15479), .C2(n15374), .A(n15373), .ZN(n15379) );
  NAND2_X1 U17493 ( .A1(n15375), .A2(n15049), .ZN(n15377) );
  INV_X1 U17494 ( .A(n15484), .ZN(n15376) );
  NAND2_X1 U17495 ( .A1(n15377), .A2(n15376), .ZN(n19454) );
  OAI22_X1 U17496 ( .A1(n18277), .A2(n16853), .B1(n16871), .B2(n19454), .ZN(
        n15378) );
  AOI211_X1 U17497 ( .C1(n15380), .C2(n16864), .A(n15379), .B(n15378), .ZN(
        n15381) );
  OAI21_X1 U17498 ( .B1(n15382), .B2(n18575), .A(n15381), .ZN(P2_U3042) );
  INV_X1 U17499 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n15397) );
  NAND3_X1 U17500 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19187) );
  INV_X1 U17501 ( .A(n19187), .ZN(n19191) );
  NAND2_X1 U17502 ( .A1(n19191), .A2(n19263), .ZN(n15387) );
  OAI21_X1 U17503 ( .B1(n19702), .B2(n19566), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n15384) );
  NAND2_X1 U17504 ( .A1(n15384), .A2(n19292), .ZN(n15391) );
  NAND3_X1 U17505 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19294), .ZN(n19209) );
  NOR2_X1 U17506 ( .A1(n19263), .A2(n19209), .ZN(n19700) );
  OAI21_X1 U17507 ( .B1(n11840), .B2(n19297), .A(n19332), .ZN(n15385) );
  OAI21_X1 U17508 ( .B1(n15391), .B2(n19700), .A(n15385), .ZN(n15386) );
  OAI21_X1 U17509 ( .B1(n19683), .B2(n15387), .A(n15386), .ZN(n19469) );
  INV_X1 U17510 ( .A(n19700), .ZN(n19199) );
  AND2_X1 U17511 ( .A1(n15387), .A2(n19199), .ZN(n15390) );
  INV_X1 U17512 ( .A(n11840), .ZN(n15388) );
  INV_X1 U17513 ( .A(n15387), .ZN(n19694) );
  OAI21_X1 U17514 ( .B1(n15388), .B2(n19694), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15389) );
  AOI22_X1 U17515 ( .A1(n19319), .A2(n19702), .B1(n19328), .B2(n19694), .ZN(
        n15393) );
  OAI21_X1 U17516 ( .B1(n15394), .B2(n19699), .A(n15393), .ZN(n15395) );
  AOI21_X1 U17517 ( .B1(n19695), .B2(n15206), .A(n15395), .ZN(n15396) );
  OAI21_X1 U17518 ( .B1(n15397), .B2(n19469), .A(n15396), .ZN(P2_U3167) );
  NAND2_X1 U17519 ( .A1(n15399), .A2(n15398), .ZN(n15400) );
  NAND2_X1 U17520 ( .A1(n15446), .A2(n15400), .ZN(n21493) );
  INV_X1 U17521 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n21479) );
  OAI222_X1 U17522 ( .A1(n21493), .A2(n15837), .B1(n21479), .B2(n19946), .C1(
        n21488), .C2(n15842), .ZN(P1_U2864) );
  XOR2_X1 U17523 ( .A(n15402), .B(n15401), .Z(n19962) );
  INV_X1 U17524 ( .A(n19962), .ZN(n15407) );
  INV_X1 U17525 ( .A(n21284), .ZN(n21294) );
  NAND2_X1 U17526 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n21294), .ZN(
        n15464) );
  NOR2_X1 U17527 ( .A1(n15403), .A2(n15464), .ZN(n16025) );
  INV_X1 U17528 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n21292) );
  AOI211_X1 U17529 ( .C1(n21283), .C2(n21337), .A(n21292), .B(n21334), .ZN(
        n15404) );
  AOI22_X1 U17530 ( .A1(n16025), .A2(n15404), .B1(n21347), .B2(n16031), .ZN(
        n15428) );
  NOR2_X1 U17531 ( .A1(n21295), .A2(n15464), .ZN(n21316) );
  INV_X1 U17532 ( .A(n21316), .ZN(n21286) );
  NOR2_X1 U17533 ( .A1(n21292), .A2(n21286), .ZN(n15426) );
  NAND2_X1 U17534 ( .A1(n21390), .A2(P1_REIP_REG_7__SCAN_IN), .ZN(n19963) );
  OAI21_X1 U17535 ( .B1(n21409), .B2(n21464), .A(n19963), .ZN(n15405) );
  AOI221_X1 U17536 ( .B1(n15428), .B2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(
        n15426), .C2(n13728), .A(n15405), .ZN(n15406) );
  OAI21_X1 U17537 ( .B1(n15407), .B2(n21327), .A(n15406), .ZN(P1_U3024) );
  OR2_X1 U17538 ( .A1(n15408), .A2(n14489), .ZN(n15409) );
  AND2_X1 U17539 ( .A1(n15409), .A2(n15420), .ZN(n18577) );
  INV_X1 U17540 ( .A(n18577), .ZN(n16547) );
  INV_X1 U17541 ( .A(n15494), .ZN(n16262) );
  OR2_X1 U17542 ( .A1(n15494), .A2(n15410), .ZN(n15414) );
  OAI211_X1 U17543 ( .C1(n16262), .C2(n15411), .A(n16252), .B(n15414), .ZN(
        n15413) );
  NAND2_X1 U17544 ( .A1(n16267), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n15412) );
  OAI211_X1 U17545 ( .C1(n16547), .C2(n16267), .A(n15413), .B(n15412), .ZN(
        P2_U2873) );
  INV_X1 U17546 ( .A(n15414), .ZN(n15418) );
  NOR2_X1 U17547 ( .A1(n15494), .A2(n15415), .ZN(n15496) );
  INV_X1 U17548 ( .A(n15496), .ZN(n15416) );
  OAI211_X1 U17549 ( .C1(n15418), .C2(n15417), .A(n15416), .B(n16252), .ZN(
        n15423) );
  NAND2_X1 U17550 ( .A1(n15420), .A2(n15419), .ZN(n15421) );
  AND2_X1 U17551 ( .A1(n15499), .A2(n15421), .ZN(n18389) );
  NAND2_X1 U17552 ( .A1(n16209), .A2(n18389), .ZN(n15422) );
  OAI211_X1 U17553 ( .C1(n16209), .C2(n11580), .A(n15423), .B(n15422), .ZN(
        P2_U2872) );
  XOR2_X1 U17554 ( .A(n15425), .B(n15424), .Z(n15440) );
  NAND2_X1 U17555 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15463) );
  OAI211_X1 U17556 ( .C1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n15426), .B(n15463), .ZN(n15430) );
  OAI22_X1 U17557 ( .A1(n21378), .A2(n21487), .B1(n21409), .B2(n21493), .ZN(
        n15427) );
  AOI21_X1 U17558 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n15428), .A(
        n15427), .ZN(n15429) );
  OAI211_X1 U17559 ( .C1(n15440), .C2(n21327), .A(n15430), .B(n15429), .ZN(
        P1_U3023) );
  OAI21_X1 U17560 ( .B1(n15432), .B2(n15434), .A(n15433), .ZN(n19970) );
  MUX2_X1 U17561 ( .A(BUF1_REG_10__SCAN_IN), .B(DATAI_10_), .S(n15599), .Z(
        n21732) );
  AOI22_X1 U17562 ( .A1(n15888), .A2(n21732), .B1(P1_EAX_REG_10__SCAN_IN), 
        .B2(n15887), .ZN(n15435) );
  OAI21_X1 U17563 ( .B1(n19970), .B2(n15890), .A(n15435), .ZN(P1_U2894) );
  INV_X1 U17564 ( .A(n21488), .ZN(n15438) );
  AOI22_X1 U17565 ( .A1(n20015), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n21390), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n15436) );
  OAI21_X1 U17566 ( .B1(n20025), .B2(n21480), .A(n15436), .ZN(n15437) );
  AOI21_X1 U17567 ( .B1(n15438), .B2(n20021), .A(n15437), .ZN(n15439) );
  OAI21_X1 U17568 ( .B1(n15440), .B2(n21578), .A(n15439), .ZN(P1_U2991) );
  INV_X1 U17569 ( .A(n15441), .ZN(n15442) );
  AOI21_X1 U17570 ( .B1(n15442), .B2(n11249), .A(n15432), .ZN(n19943) );
  INV_X1 U17571 ( .A(n19943), .ZN(n15455) );
  MUX2_X1 U17572 ( .A(BUF1_REG_9__SCAN_IN), .B(DATAI_9_), .S(n15599), .Z(
        n21724) );
  AOI22_X1 U17573 ( .A1(n15888), .A2(n21724), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n15887), .ZN(n15443) );
  OAI21_X1 U17574 ( .B1(n15455), .B2(n15890), .A(n15443), .ZN(P1_U2895) );
  INV_X1 U17575 ( .A(n15491), .ZN(n15444) );
  AOI21_X1 U17576 ( .B1(n15446), .B2(n15445), .A(n15444), .ZN(n19940) );
  INV_X1 U17577 ( .A(n19940), .ZN(n15447) );
  INV_X1 U17578 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n19945) );
  OAI22_X1 U17579 ( .A1(n15447), .A2(n21562), .B1(n19945), .B2(n21559), .ZN(
        n15453) );
  INV_X1 U17580 ( .A(n15448), .ZN(n21482) );
  OAI21_X1 U17581 ( .B1(n21411), .B2(n21482), .A(n21552), .ZN(n21486) );
  INV_X1 U17582 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n15451) );
  AOI22_X1 U17583 ( .A1(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n21536), .B1(
        n15756), .B2(n15451), .ZN(n15450) );
  OR2_X1 U17584 ( .A1(n21411), .A2(n15449), .ZN(n21560) );
  OAI211_X1 U17585 ( .C1(n21486), .C2(n15451), .A(n15450), .B(n21560), .ZN(
        n15452) );
  AOI211_X1 U17586 ( .C1(n15460), .C2(n21535), .A(n15453), .B(n15452), .ZN(
        n15454) );
  OAI21_X1 U17587 ( .B1(n15455), .B2(n21571), .A(n15454), .ZN(P1_U2831) );
  NAND2_X1 U17588 ( .A1(n15457), .A2(n15456), .ZN(n15458) );
  NAND2_X1 U17589 ( .A1(n19965), .A2(n15458), .ZN(n15471) );
  NOR2_X1 U17590 ( .A1(n21378), .A2(n15451), .ZN(n15468) );
  AND2_X1 U17591 ( .A1(n20015), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15459) );
  AOI211_X1 U17592 ( .C1(n20000), .C2(n15460), .A(n15468), .B(n15459), .ZN(
        n15462) );
  NAND2_X1 U17593 ( .A1(n19943), .A2(n20021), .ZN(n15461) );
  OAI211_X1 U17594 ( .C1(n15471), .C2(n21578), .A(n15462), .B(n15461), .ZN(
        P1_U2990) );
  NOR2_X1 U17595 ( .A1(n21292), .A2(n15463), .ZN(n16024) );
  NOR2_X1 U17596 ( .A1(n15464), .A2(n21283), .ZN(n16028) );
  INV_X1 U17597 ( .A(n16028), .ZN(n15465) );
  OAI21_X1 U17598 ( .B1(n16025), .B2(n21332), .A(n16031), .ZN(n21282) );
  AOI21_X1 U17599 ( .B1(n15465), .B2(n21337), .A(n21282), .ZN(n21312) );
  OAI21_X1 U17600 ( .B1(n16024), .B2(n21347), .A(n21312), .ZN(n21308) );
  NAND2_X1 U17601 ( .A1(n16024), .A2(n21316), .ZN(n21305) );
  INV_X1 U17602 ( .A(n21305), .ZN(n15467) );
  AOI22_X1 U17603 ( .A1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n21308), .B1(
        n15467), .B2(n15466), .ZN(n15470) );
  AOI21_X1 U17604 ( .B1(n21394), .B2(n19940), .A(n15468), .ZN(n15469) );
  OAI211_X1 U17605 ( .C1(n15471), .C2(n21327), .A(n15470), .B(n15469), .ZN(
        P1_U3022) );
  OAI21_X1 U17606 ( .B1(n15473), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n15472), .ZN(n17218) );
  XNOR2_X1 U17607 ( .A(n15475), .B(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15476) );
  XNOR2_X1 U17608 ( .A(n15474), .B(n15476), .ZN(n17217) );
  AOI221_X1 U17609 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C1(n15479), .C2(n15478), .A(
        n15477), .ZN(n15481) );
  NOR2_X1 U17610 ( .A1(n12135), .A2(n18583), .ZN(n15480) );
  AOI211_X1 U17611 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n15482), .A(
        n15481), .B(n15480), .ZN(n15487) );
  XNOR2_X1 U17612 ( .A(n15484), .B(n15483), .ZN(n19394) );
  NOR2_X1 U17613 ( .A1(n16871), .A2(n19394), .ZN(n15485) );
  AOI21_X1 U17614 ( .B1(n18286), .B2(n18603), .A(n15485), .ZN(n15486) );
  OAI211_X1 U17615 ( .C1(n17217), .C2(n18575), .A(n15487), .B(n15486), .ZN(
        n15488) );
  INV_X1 U17616 ( .A(n15488), .ZN(n15489) );
  OAI21_X1 U17617 ( .B1(n17218), .B2(n18609), .A(n15489), .ZN(P2_U3041) );
  AND2_X1 U17618 ( .A1(n15491), .A2(n15490), .ZN(n15492) );
  OR2_X1 U17619 ( .A1(n15492), .A2(n15524), .ZN(n21499) );
  INV_X1 U17620 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n21498) );
  OAI222_X1 U17621 ( .A1(n21499), .A2(n15837), .B1(n21498), .B2(n19946), .C1(
        n19970), .C2(n15842), .ZN(P1_U2862) );
  NOR2_X1 U17622 ( .A1(n15494), .A2(n15493), .ZN(n16273) );
  NOR2_X1 U17623 ( .A1(n15496), .A2(n15495), .ZN(n15497) );
  OR2_X1 U17624 ( .A1(n16273), .A2(n15497), .ZN(n19678) );
  AND2_X1 U17625 ( .A1(n15499), .A2(n15498), .ZN(n15501) );
  OR2_X1 U17626 ( .A1(n15501), .A2(n15500), .ZN(n18402) );
  NOR2_X1 U17627 ( .A1(n18402), .A2(n16267), .ZN(n15502) );
  AOI21_X1 U17628 ( .B1(P2_EBX_REG_16__SCAN_IN), .B2(n16267), .A(n15502), .ZN(
        n15503) );
  OAI21_X1 U17629 ( .B1(n19678), .B2(n16278), .A(n15503), .ZN(P2_U2871) );
  AOI21_X1 U17630 ( .B1(n15506), .B2(n15504), .A(n15505), .ZN(n15517) );
  AOI22_X1 U17631 ( .A1(n19673), .A2(BUF1_REG_19__SCAN_IN), .B1(n19674), .B2(
        BUF2_REG_19__SCAN_IN), .ZN(n15511) );
  INV_X1 U17632 ( .A(n15507), .ZN(n15508) );
  XNOR2_X1 U17633 ( .A(n15509), .B(n15508), .ZN(n18600) );
  AOI22_X1 U17634 ( .A1(n19612), .A2(n18600), .B1(n19670), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n15510) );
  OAI211_X1 U17635 ( .C1(n19517), .C2(n16352), .A(n15511), .B(n15510), .ZN(
        n15512) );
  AOI21_X1 U17636 ( .B1(n15517), .B2(n19561), .A(n15512), .ZN(n15513) );
  INV_X1 U17637 ( .A(n15513), .ZN(P2_U2900) );
  AND2_X1 U17638 ( .A1(n10963), .A2(n15514), .ZN(n15516) );
  OR2_X1 U17639 ( .A1(n15516), .A2(n15515), .ZN(n18429) );
  NAND2_X1 U17640 ( .A1(n15517), .A2(n16252), .ZN(n15519) );
  NAND2_X1 U17641 ( .A1(n16267), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n15518) );
  OAI211_X1 U17642 ( .C1(n18429), .C2(n16267), .A(n15519), .B(n15518), .ZN(
        P2_U2868) );
  NAND2_X1 U17643 ( .A1(n15433), .A2(n15520), .ZN(n15521) );
  NAND2_X1 U17644 ( .A1(n15529), .A2(n15521), .ZN(n15531) );
  INV_X1 U17645 ( .A(n15530), .ZN(n15522) );
  XNOR2_X1 U17646 ( .A(n15531), .B(n15522), .ZN(n19980) );
  INV_X1 U17647 ( .A(n19980), .ZN(n21514) );
  OR2_X1 U17648 ( .A1(n15524), .A2(n15523), .ZN(n15525) );
  NAND2_X1 U17649 ( .A1(n15535), .A2(n15525), .ZN(n21512) );
  INV_X1 U17650 ( .A(n21512), .ZN(n15526) );
  AOI22_X1 U17651 ( .A1(n19941), .A2(n15526), .B1(P1_EBX_REG_11__SCAN_IN), 
        .B2(n15840), .ZN(n15527) );
  OAI21_X1 U17652 ( .B1(n21514), .B2(n15842), .A(n15527), .ZN(P1_U2861) );
  MUX2_X1 U17653 ( .A(BUF1_REG_11__SCAN_IN), .B(DATAI_11_), .S(n15599), .Z(
        n21739) );
  AOI22_X1 U17654 ( .A1(n15888), .A2(n21739), .B1(P1_EAX_REG_11__SCAN_IN), 
        .B2(n15887), .ZN(n15528) );
  OAI21_X1 U17655 ( .B1(n21514), .B2(n15890), .A(n15528), .ZN(P1_U2893) );
  OAI21_X1 U17656 ( .B1(n15531), .B2(n15530), .A(n15529), .ZN(n15533) );
  NAND2_X1 U17657 ( .A1(n15533), .A2(n15532), .ZN(n15789) );
  OAI21_X1 U17658 ( .B1(n15533), .B2(n15532), .A(n15789), .ZN(n19987) );
  NAND2_X1 U17659 ( .A1(n15535), .A2(n15534), .ZN(n15536) );
  NAND2_X1 U17660 ( .A1(n15792), .A2(n15536), .ZN(n21522) );
  INV_X1 U17661 ( .A(n21522), .ZN(n15537) );
  AOI22_X1 U17662 ( .A1(n15537), .A2(n19941), .B1(P1_EBX_REG_12__SCAN_IN), 
        .B2(n15840), .ZN(n15538) );
  OAI21_X1 U17663 ( .B1(n19987), .B2(n15842), .A(n15538), .ZN(P1_U2860) );
  MUX2_X1 U17664 ( .A(BUF1_REG_12__SCAN_IN), .B(DATAI_12_), .S(n15599), .Z(
        n21745) );
  AOI22_X1 U17665 ( .A1(n15888), .A2(n21745), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n15887), .ZN(n15539) );
  OAI21_X1 U17666 ( .B1(n19987), .B2(n15890), .A(n15539), .ZN(P1_U2892) );
  NOR2_X1 U17667 ( .A1(n15787), .A2(n15540), .ZN(n15541) );
  OR2_X1 U17668 ( .A1(n15769), .A2(n15541), .ZN(n19998) );
  NOR2_X1 U17669 ( .A1(n15790), .A2(n15543), .ZN(n15544) );
  OR2_X1 U17670 ( .A1(n15542), .A2(n15544), .ZN(n21281) );
  OAI22_X1 U17671 ( .A1(n21281), .A2(n15837), .B1(n15777), .B2(n19946), .ZN(
        n15545) );
  INV_X1 U17672 ( .A(n15545), .ZN(n15546) );
  OAI21_X1 U17673 ( .B1(n19998), .B2(n15842), .A(n15546), .ZN(P1_U2858) );
  MUX2_X1 U17674 ( .A(BUF1_REG_14__SCAN_IN), .B(DATAI_14_), .S(n15599), .Z(
        n21759) );
  AOI22_X1 U17675 ( .A1(n15888), .A2(n21759), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n15887), .ZN(n15547) );
  OAI21_X1 U17676 ( .B1(n19998), .B2(n15890), .A(n15547), .ZN(P1_U2890) );
  OAI21_X1 U17677 ( .B1(n15559), .B2(n15549), .A(n15548), .ZN(n16260) );
  AOI22_X1 U17678 ( .A1(n19673), .A2(BUF1_REG_21__SCAN_IN), .B1(n19674), .B2(
        BUF2_REG_21__SCAN_IN), .ZN(n15554) );
  OR2_X1 U17679 ( .A1(n15550), .A2(n15551), .ZN(n15552) );
  AND2_X1 U17680 ( .A1(n15552), .A2(n16669), .ZN(n18449) );
  AOI22_X1 U17681 ( .A1(n19612), .A2(n18449), .B1(n19670), .B2(
        P2_EAX_REG_21__SCAN_IN), .ZN(n15553) );
  OAI211_X1 U17682 ( .C1(n19398), .C2(n16352), .A(n15554), .B(n15553), .ZN(
        n15555) );
  INV_X1 U17683 ( .A(n15555), .ZN(n15556) );
  OAI21_X1 U17684 ( .B1(n16260), .B2(n19677), .A(n15556), .ZN(P2_U2898) );
  AND2_X1 U17685 ( .A1(n15558), .A2(n15557), .ZN(n15560) );
  OR2_X1 U17686 ( .A1(n15560), .A2(n15559), .ZN(n19441) );
  OR2_X1 U17687 ( .A1(n15515), .A2(n15562), .ZN(n15563) );
  NAND2_X1 U17688 ( .A1(n15561), .A2(n15563), .ZN(n18448) );
  NOR2_X1 U17689 ( .A1(n18448), .A2(n16267), .ZN(n15564) );
  AOI21_X1 U17690 ( .B1(P2_EBX_REG_20__SCAN_IN), .B2(n16267), .A(n15564), .ZN(
        n15565) );
  OAI21_X1 U17691 ( .B1(n19441), .B2(n16278), .A(n15565), .ZN(P2_U2867) );
  INV_X1 U17692 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21201) );
  INV_X1 U17693 ( .A(n17743), .ZN(n15572) );
  NOR2_X1 U17694 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n15572), .ZN(n20097) );
  NOR2_X1 U17695 ( .A1(n20754), .A2(n21612), .ZN(n18001) );
  INV_X1 U17696 ( .A(n18001), .ZN(n18096) );
  NAND2_X1 U17697 ( .A1(n20097), .A2(n18096), .ZN(n15566) );
  OAI21_X1 U17698 ( .B1(n21201), .B2(n21232), .A(n15566), .ZN(n18142) );
  INV_X1 U17699 ( .A(n18142), .ZN(n15567) );
  NOR2_X1 U17700 ( .A1(n18145), .A2(n15567), .ZN(n15569) );
  NAND3_X1 U17701 ( .A1(n21098), .A2(n21232), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18771) );
  INV_X1 U17702 ( .A(n18771), .ZN(n15570) );
  NOR2_X1 U17703 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21232), .ZN(
        n18715) );
  OR3_X1 U17704 ( .A1(n15570), .A2(n18715), .A3(n18145), .ZN(n15568) );
  MUX2_X1 U17705 ( .A(n15569), .B(n15568), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  AOI21_X1 U17706 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18142), .A(
        n15570), .ZN(n15571) );
  NOR2_X1 U17707 ( .A1(n18145), .A2(n15571), .ZN(n15575) );
  NAND2_X1 U17708 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18714) );
  OAI21_X1 U17709 ( .B1(n15572), .B2(n18001), .A(n21232), .ZN(n15573) );
  AOI211_X1 U17710 ( .C1(n18714), .C2(n15573), .A(n18145), .B(n18715), .ZN(
        n18143) );
  INV_X1 U17711 ( .A(n18143), .ZN(n15574) );
  MUX2_X1 U17712 ( .A(n15575), .B(n15574), .S(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .Z(P3_U2865) );
  NOR2_X1 U17713 ( .A1(n15577), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15578) );
  AOI21_X1 U17714 ( .B1(n21581), .B2(n15579), .A(n15578), .ZN(n16953) );
  AOI22_X1 U17715 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n21400), .B1(n15576), 
        .B2(n21597), .ZN(n15580) );
  OAI21_X1 U17716 ( .B1(n16953), .B2(n16171), .A(n15580), .ZN(n15583) );
  NOR2_X1 U17717 ( .A1(n15581), .A2(n15576), .ZN(n16951) );
  AOI22_X1 U17718 ( .A1(n15585), .A2(n15583), .B1(n15582), .B2(n16951), .ZN(
        n15584) );
  OAI21_X1 U17719 ( .B1(n15576), .B2(n15585), .A(n15584), .ZN(P1_U3474) );
  OAI21_X1 U17720 ( .B1(n15640), .B2(n15587), .A(n15629), .ZN(n15602) );
  INV_X1 U17721 ( .A(n15602), .ZN(n16071) );
  INV_X1 U17722 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n15624) );
  NAND2_X1 U17723 ( .A1(n15625), .A2(n21552), .ZN(n15642) );
  INV_X1 U17724 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n15603) );
  OAI22_X1 U17725 ( .A1(n21566), .A2(n15588), .B1(n21559), .B2(n15603), .ZN(
        n15590) );
  NOR3_X1 U17726 ( .A1(n15625), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n21459), 
        .ZN(n15589) );
  AOI211_X1 U17727 ( .C1(n21535), .C2(n15591), .A(n15590), .B(n15589), .ZN(
        n15592) );
  OAI21_X1 U17728 ( .B1(n15624), .B2(n15642), .A(n15592), .ZN(n15593) );
  AOI21_X1 U17729 ( .B1(n16071), .B2(n21469), .A(n15593), .ZN(n15594) );
  OAI21_X1 U17730 ( .B1(n15586), .B2(n21571), .A(n15594), .ZN(P1_U2811) );
  AOI22_X1 U17731 ( .A1(n15877), .A2(DATAI_29_), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n15887), .ZN(n15601) );
  NOR3_X1 U17732 ( .A1(n15887), .A2(n15597), .A3(n15596), .ZN(n15598) );
  MUX2_X1 U17733 ( .A(BUF1_REG_13__SCAN_IN), .B(DATAI_13_), .S(n15599), .Z(
        n21752) );
  AOI22_X1 U17734 ( .A1(n15880), .A2(n21752), .B1(BUF1_REG_29__SCAN_IN), .B2(
        n15878), .ZN(n15600) );
  OAI211_X1 U17735 ( .C1(n15586), .C2(n15890), .A(n15601), .B(n15600), .ZN(
        P1_U2875) );
  OAI222_X1 U17736 ( .A1(n15842), .A2(n15586), .B1(n15603), .B2(n19946), .C1(
        n15602), .C2(n15837), .ZN(P1_U2843) );
  NOR2_X1 U17737 ( .A1(n15604), .A2(n16267), .ZN(n15605) );
  AOI21_X1 U17738 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n16267), .A(n15605), .ZN(
        n15606) );
  OAI21_X1 U17739 ( .B1(n15607), .B2(n16278), .A(n15606), .ZN(P2_U2857) );
  AOI22_X1 U17740 ( .A1(n15613), .A2(n12614), .B1(n13523), .B2(n15608), .ZN(
        n15616) );
  NAND2_X1 U17741 ( .A1(n15610), .A2(n15609), .ZN(n15615) );
  INV_X1 U17742 ( .A(n15611), .ZN(n15612) );
  NAND2_X1 U17743 ( .A1(n15613), .A2(n15612), .ZN(n15614) );
  AND3_X1 U17744 ( .A1(n15616), .A2(n15615), .A3(n15614), .ZN(n16966) );
  INV_X1 U17745 ( .A(n16966), .ZN(n15621) );
  NOR2_X1 U17746 ( .A1(n15618), .A2(n15617), .ZN(n21252) );
  OAI21_X1 U17747 ( .B1(n21624), .B2(n21252), .A(n15619), .ZN(n16964) );
  AND2_X1 U17748 ( .A1(n16964), .A2(n15620), .ZN(n21579) );
  MUX2_X1 U17749 ( .A(P1_MORE_REG_SCAN_IN), .B(n15621), .S(n21579), .Z(
        P1_U3484) );
  AOI21_X1 U17750 ( .B1(n15623), .B2(n10987), .A(n15622), .ZN(n15900) );
  INV_X1 U17751 ( .A(n15900), .ZN(n15845) );
  INV_X1 U17752 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n17089) );
  OAI21_X1 U17753 ( .B1(n15625), .B2(n15624), .A(n17089), .ZN(n15633) );
  AOI22_X1 U17754 ( .A1(n21536), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B1(
        n21533), .B2(P1_EBX_REG_30__SCAN_IN), .ZN(n15626) );
  OAI21_X1 U17755 ( .B1(n15898), .B2(n21565), .A(n15626), .ZN(n15632) );
  INV_X1 U17756 ( .A(n15627), .ZN(n15628) );
  AOI22_X1 U17757 ( .A1(n15629), .A2(n13547), .B1(n15628), .B2(n15640), .ZN(
        n15631) );
  AOI21_X1 U17758 ( .B1(n15636), .B2(n15635), .A(n13779), .ZN(n15637) );
  INV_X1 U17759 ( .A(n15637), .ZN(n15915) );
  AND2_X1 U17760 ( .A1(n15658), .A2(n15638), .ZN(n15639) );
  NOR2_X1 U17761 ( .A1(n15640), .A2(n15639), .ZN(n16075) );
  INV_X1 U17762 ( .A(n15717), .ZN(n15678) );
  INV_X1 U17763 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n17081) );
  NOR2_X1 U17764 ( .A1(n21459), .A2(n17081), .ZN(n15641) );
  NAND2_X1 U17765 ( .A1(n15678), .A2(n15641), .ZN(n15700) );
  INV_X1 U17766 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n16981) );
  NOR3_X1 U17767 ( .A1(n15700), .A2(n15666), .A3(n16981), .ZN(n15662) );
  AOI21_X1 U17768 ( .B1(n15662), .B2(P1_REIP_REG_27__SCAN_IN), .A(
        P1_REIP_REG_28__SCAN_IN), .ZN(n15643) );
  NOR2_X1 U17769 ( .A1(n15643), .A2(n15642), .ZN(n15646) );
  AOI22_X1 U17770 ( .A1(n21536), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .B1(
        n21533), .B2(P1_EBX_REG_28__SCAN_IN), .ZN(n15644) );
  OAI21_X1 U17771 ( .B1(n15902), .B2(n21565), .A(n15644), .ZN(n15645) );
  AOI211_X1 U17772 ( .C1(n16075), .C2(n21469), .A(n15646), .B(n15645), .ZN(
        n15647) );
  OAI21_X1 U17773 ( .B1(n15915), .B2(n21571), .A(n15647), .ZN(P1_U2812) );
  OAI21_X2 U17774 ( .B1(n15648), .B2(n15649), .A(n15635), .ZN(n15919) );
  INV_X1 U17775 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n17194) );
  INV_X1 U17776 ( .A(n15922), .ZN(n15653) );
  NOR2_X1 U17777 ( .A1(n21495), .A2(n15650), .ZN(n15672) );
  NAND2_X1 U17778 ( .A1(n15672), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n15652) );
  AOI22_X1 U17779 ( .A1(n21536), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B1(
        n21533), .B2(P1_EBX_REG_27__SCAN_IN), .ZN(n15651) );
  OAI211_X1 U17780 ( .C1(n21565), .C2(n15653), .A(n15652), .B(n15651), .ZN(
        n15661) );
  INV_X1 U17781 ( .A(n15655), .ZN(n15668) );
  INV_X1 U17782 ( .A(n15656), .ZN(n15657) );
  OAI21_X1 U17783 ( .B1(n15654), .B2(n15668), .A(n15657), .ZN(n15659) );
  NAND2_X1 U17784 ( .A1(n15659), .A2(n15658), .ZN(n16086) );
  NOR2_X1 U17785 ( .A1(n16086), .A2(n21562), .ZN(n15660) );
  AOI211_X1 U17786 ( .C1(n15662), .C2(n17194), .A(n15661), .B(n15660), .ZN(
        n15663) );
  OAI21_X1 U17787 ( .B1(n15919), .B2(n21571), .A(n15663), .ZN(P1_U2813) );
  AOI21_X1 U17788 ( .B1(n15665), .B2(n15664), .A(n15648), .ZN(n15928) );
  INV_X1 U17789 ( .A(n15928), .ZN(n15852) );
  OAI21_X1 U17790 ( .B1(n15700), .B2(n15666), .A(n16981), .ZN(n15671) );
  AOI22_X1 U17791 ( .A1(n21536), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n21533), .B2(P1_EBX_REG_26__SCAN_IN), .ZN(n15667) );
  OAI21_X1 U17792 ( .B1(n15926), .B2(n21565), .A(n15667), .ZN(n15670) );
  XNOR2_X1 U17793 ( .A(n15654), .B(n15668), .ZN(n16096) );
  NOR2_X1 U17794 ( .A1(n16096), .A2(n21562), .ZN(n15669) );
  AOI211_X1 U17795 ( .C1(n15672), .C2(n15671), .A(n15670), .B(n15669), .ZN(
        n15673) );
  OAI21_X1 U17796 ( .B1(n15852), .B2(n21571), .A(n15673), .ZN(P1_U2814) );
  OAI21_X1 U17797 ( .B1(n15674), .B2(n15675), .A(n15664), .ZN(n15938) );
  OR2_X1 U17798 ( .A1(n15689), .A2(n15676), .ZN(n15677) );
  NAND2_X1 U17799 ( .A1(n15654), .A2(n15677), .ZN(n16108) );
  INV_X1 U17800 ( .A(n16108), .ZN(n15685) );
  INV_X1 U17801 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n16983) );
  NAND3_X1 U17802 ( .A1(n15678), .A2(P1_REIP_REG_22__SCAN_IN), .A3(
        P1_REIP_REG_23__SCAN_IN), .ZN(n15679) );
  AND2_X1 U17803 ( .A1(n15679), .A2(n21552), .ZN(n15702) );
  AOI21_X1 U17804 ( .B1(n21483), .B2(n16983), .A(n15702), .ZN(n15683) );
  INV_X1 U17805 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n17085) );
  INV_X1 U17806 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n15807) );
  OAI22_X1 U17807 ( .A1(n21566), .A2(n15930), .B1(n21559), .B2(n15807), .ZN(
        n15681) );
  INV_X1 U17808 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n17086) );
  NOR4_X1 U17809 ( .A1(n15700), .A2(P1_REIP_REG_25__SCAN_IN), .A3(n16983), 
        .A4(n17086), .ZN(n15680) );
  AOI211_X1 U17810 ( .C1(n21535), .C2(n15932), .A(n15681), .B(n15680), .ZN(
        n15682) );
  OAI21_X1 U17811 ( .B1(n15683), .B2(n17085), .A(n15682), .ZN(n15684) );
  AOI21_X1 U17812 ( .B1(n15685), .B2(n21469), .A(n15684), .ZN(n15686) );
  OAI21_X1 U17813 ( .B1(n15938), .B2(n21571), .A(n15686), .ZN(P1_U2815) );
  NOR2_X1 U17814 ( .A1(n11020), .A2(n15687), .ZN(n15688) );
  OR2_X1 U17815 ( .A1(n15689), .A2(n15688), .ZN(n16122) );
  AOI21_X1 U17816 ( .B1(n15691), .B2(n15690), .A(n15674), .ZN(n15945) );
  NAND2_X1 U17817 ( .A1(n15945), .A2(n21541), .ZN(n15696) );
  NOR3_X1 U17818 ( .A1(n15700), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n17086), 
        .ZN(n15694) );
  AOI22_X1 U17819 ( .A1(n21536), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n21533), .B2(P1_EBX_REG_24__SCAN_IN), .ZN(n15692) );
  OAI21_X1 U17820 ( .B1(n15943), .B2(n21565), .A(n15692), .ZN(n15693) );
  AOI211_X1 U17821 ( .C1(n15702), .C2(P1_REIP_REG_24__SCAN_IN), .A(n15694), 
        .B(n15693), .ZN(n15695) );
  OAI211_X1 U17822 ( .C1(n16122), .C2(n21562), .A(n15696), .B(n15695), .ZN(
        P1_U2816) );
  OAI21_X1 U17823 ( .B1(n10988), .B2(n15697), .A(n15690), .ZN(n15950) );
  NOR2_X1 U17824 ( .A1(n15712), .A2(n15698), .ZN(n15699) );
  OR2_X1 U17825 ( .A1(n11020), .A2(n15699), .ZN(n15809) );
  INV_X1 U17826 ( .A(n15809), .ZN(n21393) );
  INV_X1 U17827 ( .A(n15953), .ZN(n15706) );
  NAND2_X1 U17828 ( .A1(n15700), .A2(n17086), .ZN(n15701) );
  NAND2_X1 U17829 ( .A1(n15702), .A2(n15701), .ZN(n15705) );
  INV_X1 U17830 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n15810) );
  OAI22_X1 U17831 ( .A1(n21566), .A2(n15949), .B1(n21559), .B2(n15810), .ZN(
        n15703) );
  INV_X1 U17832 ( .A(n15703), .ZN(n15704) );
  OAI211_X1 U17833 ( .C1(n21565), .C2(n15706), .A(n15705), .B(n15704), .ZN(
        n15707) );
  AOI21_X1 U17834 ( .B1(n21393), .B2(n21469), .A(n15707), .ZN(n15708) );
  OAI21_X1 U17835 ( .B1(n15950), .B2(n21571), .A(n15708), .ZN(P1_U2817) );
  AOI21_X1 U17836 ( .B1(n15710), .B2(n15709), .A(n10988), .ZN(n15961) );
  AND2_X1 U17837 ( .A1(n15727), .A2(n15711), .ZN(n15713) );
  OR2_X1 U17838 ( .A1(n15713), .A2(n15712), .ZN(n21389) );
  INV_X1 U17839 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15811) );
  INV_X1 U17840 ( .A(n15714), .ZN(n15732) );
  NAND3_X1 U17841 ( .A1(n15732), .A2(P1_REIP_REG_21__SCAN_IN), .A3(n17081), 
        .ZN(n15715) );
  OAI22_X1 U17842 ( .A1(n21559), .A2(n15811), .B1(n21459), .B2(n15715), .ZN(
        n15716) );
  AOI21_X1 U17843 ( .B1(n21536), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15716), .ZN(n15721) );
  NAND3_X1 U17844 ( .A1(n21552), .A2(n15717), .A3(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n15718) );
  OAI21_X1 U17845 ( .B1(n21565), .B2(n15959), .A(n15718), .ZN(n15719) );
  INV_X1 U17846 ( .A(n15719), .ZN(n15720) );
  OAI211_X1 U17847 ( .C1(n21389), .C2(n21562), .A(n15721), .B(n15720), .ZN(
        n15722) );
  AOI21_X1 U17848 ( .B1(n15961), .B2(n21541), .A(n15722), .ZN(n15723) );
  INV_X1 U17849 ( .A(n15723), .ZN(P1_U2818) );
  OAI21_X1 U17850 ( .B1(n15725), .B2(n15726), .A(n15709), .ZN(n15967) );
  INV_X1 U17851 ( .A(n15727), .ZN(n15728) );
  AOI21_X1 U17852 ( .B1(n15729), .B2(n15748), .A(n15728), .ZN(n16136) );
  NOR2_X1 U17853 ( .A1(n15730), .A2(n21495), .ZN(n15744) );
  AOI22_X1 U17854 ( .A1(n15970), .A2(n21535), .B1(P1_REIP_REG_21__SCAN_IN), 
        .B2(n15744), .ZN(n15737) );
  INV_X1 U17855 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15734) );
  INV_X1 U17856 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n15731) );
  NAND2_X1 U17857 ( .A1(n15732), .A2(n15731), .ZN(n15733) );
  OAI22_X1 U17858 ( .A1(n21559), .A2(n15734), .B1(n21459), .B2(n15733), .ZN(
        n15735) );
  INV_X1 U17859 ( .A(n15735), .ZN(n15736) );
  OAI211_X1 U17860 ( .C1(n15966), .C2(n21566), .A(n15737), .B(n15736), .ZN(
        n15738) );
  AOI21_X1 U17861 ( .B1(n16136), .B2(n21469), .A(n15738), .ZN(n15739) );
  OAI21_X1 U17862 ( .B1(n15967), .B2(n21571), .A(n15739), .ZN(P1_U2819) );
  INV_X1 U17864 ( .A(n15725), .ZN(n15742) );
  OAI21_X1 U17865 ( .B1(n15743), .B2(n15741), .A(n15742), .ZN(n15979) );
  OAI221_X1 U17866 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(n15745), .C1(
        P1_REIP_REG_20__SCAN_IN), .C2(n15756), .A(n15744), .ZN(n15753) );
  NAND2_X1 U17867 ( .A1(n15762), .A2(n15746), .ZN(n15747) );
  NAND2_X1 U17868 ( .A1(n15748), .A2(n15747), .ZN(n16143) );
  OAI22_X1 U17869 ( .A1(n16143), .A2(n21562), .B1(n15973), .B2(n21565), .ZN(
        n15751) );
  INV_X1 U17870 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15749) );
  INV_X1 U17871 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15813) );
  OAI22_X1 U17872 ( .A1(n21566), .A2(n15749), .B1(n21559), .B2(n15813), .ZN(
        n15750) );
  NOR2_X1 U17873 ( .A1(n15751), .A2(n15750), .ZN(n15752) );
  OAI211_X1 U17874 ( .C1(n15979), .C2(n21571), .A(n15753), .B(n15752), .ZN(
        P1_U2820) );
  INV_X1 U17875 ( .A(n15741), .ZN(n15754) );
  OAI21_X1 U17876 ( .B1(n15755), .B2(n11016), .A(n15754), .ZN(n15983) );
  INV_X1 U17877 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n21359) );
  INV_X1 U17878 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n19894) );
  INV_X1 U17879 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n21313) );
  INV_X1 U17880 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n21496) );
  NAND2_X1 U17881 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n15756), .ZN(n21494) );
  NAND2_X1 U17882 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n21510), .ZN(n21509) );
  NAND2_X1 U17883 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n21529), .ZN(n15785) );
  NOR2_X1 U17884 ( .A1(n19894), .A2(n15785), .ZN(n15770) );
  NAND2_X1 U17885 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n15770), .ZN(n21530) );
  NOR2_X1 U17886 ( .A1(n21359), .A2(n21530), .ZN(n21554) );
  NAND2_X1 U17887 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n21554), .ZN(n21577) );
  INV_X1 U17888 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n21576) );
  NOR2_X1 U17889 ( .A1(n21577), .A2(n21576), .ZN(n15758) );
  AOI21_X1 U17890 ( .B1(n15758), .B2(P1_REIP_REG_19__SCAN_IN), .A(n21495), 
        .ZN(n15757) );
  OAI21_X1 U17891 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(n15758), .A(n15757), 
        .ZN(n15767) );
  OR2_X1 U17892 ( .A1(n15759), .A2(n15760), .ZN(n15761) );
  NAND2_X1 U17893 ( .A1(n15762), .A2(n15761), .ZN(n21370) );
  INV_X1 U17894 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n15814) );
  OAI22_X1 U17895 ( .A1(n21370), .A2(n21562), .B1(n21559), .B2(n15814), .ZN(
        n15763) );
  INV_X1 U17896 ( .A(n15763), .ZN(n15764) );
  OAI211_X1 U17897 ( .C1(n21566), .C2(n15982), .A(n15764), .B(n21560), .ZN(
        n15765) );
  AOI21_X1 U17898 ( .B1(n21535), .B2(n15986), .A(n15765), .ZN(n15766) );
  OAI211_X1 U17899 ( .C1(n15983), .C2(n21571), .A(n15767), .B(n15766), .ZN(
        P1_U2821) );
  OAI21_X1 U17900 ( .B1(n15769), .B2(n15768), .A(n15834), .ZN(n16009) );
  NOR2_X1 U17901 ( .A1(n21495), .A2(n15770), .ZN(n15783) );
  INV_X1 U17902 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n21338) );
  AOI22_X1 U17903 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n15783), .B1(n15770), 
        .B2(n21338), .ZN(n15776) );
  OAI21_X1 U17904 ( .B1(n15542), .B2(n15771), .A(n15829), .ZN(n15839) );
  INV_X1 U17905 ( .A(n15839), .ZN(n21330) );
  INV_X1 U17906 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n15838) );
  OAI22_X1 U17907 ( .A1(n21565), .A2(n16003), .B1(n15838), .B2(n21559), .ZN(
        n15772) );
  INV_X1 U17908 ( .A(n15772), .ZN(n15773) );
  OAI211_X1 U17909 ( .C1(n21566), .C2(n16004), .A(n15773), .B(n21560), .ZN(
        n15774) );
  AOI21_X1 U17910 ( .B1(n21330), .B2(n21469), .A(n15774), .ZN(n15775) );
  OAI211_X1 U17911 ( .C1(n16009), .C2(n21571), .A(n15776), .B(n15775), .ZN(
        P1_U2825) );
  NAND2_X1 U17912 ( .A1(n19894), .A2(n15785), .ZN(n15782) );
  AOI22_X1 U17913 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n21536), .B1(
        n21535), .B2(n19999), .ZN(n15780) );
  INV_X1 U17914 ( .A(n21560), .ZN(n21532) );
  OAI22_X1 U17915 ( .A1(n21281), .A2(n21562), .B1(n15777), .B2(n21559), .ZN(
        n15778) );
  NOR2_X1 U17916 ( .A1(n21532), .A2(n15778), .ZN(n15779) );
  NAND2_X1 U17917 ( .A1(n15780), .A2(n15779), .ZN(n15781) );
  AOI21_X1 U17918 ( .B1(n15783), .B2(n15782), .A(n15781), .ZN(n15784) );
  OAI21_X1 U17919 ( .B1(n19998), .B2(n21571), .A(n15784), .ZN(P1_U2826) );
  AOI21_X1 U17920 ( .B1(P1_REIP_REG_13__SCAN_IN), .B2(n21552), .A(n21529), 
        .ZN(n15800) );
  INV_X1 U17921 ( .A(n15785), .ZN(n15799) );
  INV_X1 U17922 ( .A(n15786), .ZN(n15788) );
  AOI21_X1 U17923 ( .B1(n15789), .B2(n15788), .A(n15787), .ZN(n16019) );
  NAND2_X1 U17924 ( .A1(n16019), .A2(n21541), .ZN(n15798) );
  INV_X1 U17925 ( .A(n16017), .ZN(n15796) );
  AOI21_X1 U17926 ( .B1(n15792), .B2(n15791), .A(n15790), .ZN(n21261) );
  AOI22_X1 U17927 ( .A1(n21469), .A2(n21261), .B1(n21533), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n15793) );
  OAI211_X1 U17928 ( .C1(n21566), .C2(n15794), .A(n15793), .B(n21560), .ZN(
        n15795) );
  AOI21_X1 U17929 ( .B1(n21535), .B2(n15796), .A(n15795), .ZN(n15797) );
  OAI211_X1 U17930 ( .C1(n15800), .C2(n15799), .A(n15798), .B(n15797), .ZN(
        P1_U2827) );
  OAI22_X1 U17931 ( .A1(n16022), .A2(n15837), .B1(n19946), .B2(n15801), .ZN(
        P1_U2841) );
  INV_X1 U17932 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n15803) );
  OAI222_X1 U17933 ( .A1(n15845), .A2(n15842), .B1(n15803), .B2(n19946), .C1(
        n15837), .C2(n15802), .ZN(P1_U2842) );
  AOI22_X1 U17934 ( .A1(n16075), .A2(n19941), .B1(P1_EBX_REG_28__SCAN_IN), 
        .B2(n15840), .ZN(n15804) );
  OAI21_X1 U17935 ( .B1(n15915), .B2(n15842), .A(n15804), .ZN(P1_U2844) );
  INV_X1 U17936 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n15805) );
  OAI222_X1 U17937 ( .A1(n15842), .A2(n15919), .B1(n15805), .B2(n19946), .C1(
        n16086), .C2(n15837), .ZN(P1_U2845) );
  INV_X1 U17938 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n15806) );
  OAI222_X1 U17939 ( .A1(n15852), .A2(n15842), .B1(n15806), .B2(n19946), .C1(
        n15837), .C2(n16096), .ZN(P1_U2846) );
  OAI222_X1 U17940 ( .A1(n15938), .A2(n15842), .B1(n15807), .B2(n19946), .C1(
        n16108), .C2(n15837), .ZN(P1_U2847) );
  INV_X1 U17941 ( .A(n15945), .ZN(n15857) );
  INV_X1 U17942 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n15808) );
  OAI222_X1 U17943 ( .A1(n15842), .A2(n15857), .B1(n15808), .B2(n19946), .C1(
        n16122), .C2(n15837), .ZN(P1_U2848) );
  OAI222_X1 U17944 ( .A1(n15950), .A2(n15842), .B1(n15810), .B2(n19946), .C1(
        n15809), .C2(n15837), .ZN(P1_U2849) );
  INV_X1 U17945 ( .A(n15961), .ZN(n15863) );
  OAI222_X1 U17946 ( .A1(n21389), .A2(n15837), .B1(n15811), .B2(n19946), .C1(
        n15863), .C2(n15842), .ZN(P1_U2850) );
  AOI22_X1 U17947 ( .A1(n16136), .A2(n19941), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n15840), .ZN(n15812) );
  OAI21_X1 U17948 ( .B1(n15967), .B2(n15842), .A(n15812), .ZN(P1_U2851) );
  OAI222_X1 U17949 ( .A1(n15979), .A2(n15842), .B1(n15813), .B2(n19946), .C1(
        n16143), .C2(n15837), .ZN(P1_U2852) );
  OAI222_X1 U17950 ( .A1(n15983), .A2(n15842), .B1(n15814), .B2(n19946), .C1(
        n21370), .C2(n15837), .ZN(P1_U2853) );
  NOR2_X1 U17951 ( .A1(n15823), .A2(n15815), .ZN(n15816) );
  OR2_X1 U17952 ( .A1(n15759), .A2(n15816), .ZN(n21563) );
  INV_X1 U17953 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n21558) );
  OR2_X1 U17954 ( .A1(n15834), .A2(n15817), .ZN(n15821) );
  OR2_X1 U17955 ( .A1(n11386), .A2(n11016), .ZN(n21572) );
  OAI222_X1 U17956 ( .A1(n21563), .A2(n15837), .B1(n21558), .B2(n19946), .C1(
        n21572), .C2(n15842), .ZN(P1_U2854) );
  OR2_X1 U17957 ( .A1(n15834), .A2(n15835), .ZN(n15832) );
  NAND2_X1 U17958 ( .A1(n15832), .A2(n15819), .ZN(n15820) );
  NAND2_X1 U17959 ( .A1(n15821), .A2(n15820), .ZN(n21550) );
  AND2_X1 U17960 ( .A1(n15831), .A2(n15822), .ZN(n15824) );
  OR2_X1 U17961 ( .A1(n15824), .A2(n15823), .ZN(n21557) );
  INV_X1 U17962 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n15825) );
  OAI22_X1 U17963 ( .A1(n21557), .A2(n15837), .B1(n15825), .B2(n19946), .ZN(
        n15826) );
  INV_X1 U17964 ( .A(n15826), .ZN(n15827) );
  OAI21_X1 U17965 ( .B1(n21550), .B2(n15842), .A(n15827), .ZN(P1_U2855) );
  NAND2_X1 U17966 ( .A1(n15829), .A2(n15828), .ZN(n15830) );
  NAND2_X1 U17967 ( .A1(n15831), .A2(n15830), .ZN(n21544) );
  INV_X1 U17968 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n15836) );
  INV_X1 U17969 ( .A(n15832), .ZN(n15833) );
  AOI21_X1 U17970 ( .B1(n15835), .B2(n15834), .A(n15833), .ZN(n21542) );
  INV_X1 U17971 ( .A(n21542), .ZN(n15883) );
  OAI222_X1 U17972 ( .A1(n21544), .A2(n15837), .B1(n15836), .B2(n19946), .C1(
        n15883), .C2(n15842), .ZN(P1_U2856) );
  OAI222_X1 U17973 ( .A1(n15839), .A2(n15837), .B1(n15838), .B2(n19946), .C1(
        n16009), .C2(n15842), .ZN(P1_U2857) );
  INV_X1 U17974 ( .A(n16019), .ZN(n15891) );
  AOI22_X1 U17975 ( .A1(n21261), .A2(n19941), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n15840), .ZN(n15841) );
  OAI21_X1 U17976 ( .B1(n15891), .B2(n15842), .A(n15841), .ZN(P1_U2859) );
  AOI22_X1 U17977 ( .A1(n15877), .A2(DATAI_30_), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n15887), .ZN(n15844) );
  AOI22_X1 U17978 ( .A1(n15880), .A2(n21759), .B1(BUF1_REG_30__SCAN_IN), .B2(
        n15878), .ZN(n15843) );
  OAI211_X1 U17979 ( .C1(n15845), .C2(n15890), .A(n15844), .B(n15843), .ZN(
        P1_U2874) );
  AOI22_X1 U17980 ( .A1(n15877), .A2(DATAI_28_), .B1(P1_EAX_REG_28__SCAN_IN), 
        .B2(n15887), .ZN(n15847) );
  AOI22_X1 U17981 ( .A1(n15880), .A2(n21745), .B1(BUF1_REG_28__SCAN_IN), .B2(
        n15878), .ZN(n15846) );
  OAI211_X1 U17982 ( .C1(n15915), .C2(n15890), .A(n15847), .B(n15846), .ZN(
        P1_U2876) );
  AOI22_X1 U17983 ( .A1(n15877), .A2(DATAI_27_), .B1(P1_EAX_REG_27__SCAN_IN), 
        .B2(n15887), .ZN(n15849) );
  AOI22_X1 U17984 ( .A1(n15880), .A2(n21739), .B1(BUF1_REG_27__SCAN_IN), .B2(
        n15878), .ZN(n15848) );
  OAI211_X1 U17985 ( .C1(n15919), .C2(n15890), .A(n15849), .B(n15848), .ZN(
        P1_U2877) );
  AOI22_X1 U17986 ( .A1(n15877), .A2(DATAI_26_), .B1(P1_EAX_REG_26__SCAN_IN), 
        .B2(n15887), .ZN(n15851) );
  AOI22_X1 U17987 ( .A1(n15880), .A2(n21732), .B1(BUF1_REG_26__SCAN_IN), .B2(
        n15878), .ZN(n15850) );
  OAI211_X1 U17988 ( .C1(n15852), .C2(n15890), .A(n15851), .B(n15850), .ZN(
        P1_U2878) );
  AOI22_X1 U17989 ( .A1(n15877), .A2(DATAI_25_), .B1(P1_EAX_REG_25__SCAN_IN), 
        .B2(n15887), .ZN(n15854) );
  AOI22_X1 U17990 ( .A1(n15880), .A2(n21724), .B1(n15878), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n15853) );
  OAI211_X1 U17991 ( .C1(n15938), .C2(n15890), .A(n15854), .B(n15853), .ZN(
        P1_U2879) );
  AOI22_X1 U17992 ( .A1(n15877), .A2(DATAI_24_), .B1(P1_EAX_REG_24__SCAN_IN), 
        .B2(n15887), .ZN(n15856) );
  AOI22_X1 U17993 ( .A1(n15880), .A2(n21717), .B1(n15878), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n15855) );
  OAI211_X1 U17994 ( .C1(n15857), .C2(n15890), .A(n15856), .B(n15855), .ZN(
        P1_U2880) );
  AOI22_X1 U17995 ( .A1(n15877), .A2(DATAI_23_), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n15887), .ZN(n15860) );
  AOI22_X1 U17996 ( .A1(n15880), .A2(n15858), .B1(n15878), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n15859) );
  OAI211_X1 U17997 ( .C1(n15950), .C2(n15890), .A(n15860), .B(n15859), .ZN(
        P1_U2881) );
  AOI22_X1 U17998 ( .A1(n15877), .A2(DATAI_22_), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n15887), .ZN(n15862) );
  AOI22_X1 U17999 ( .A1(n15880), .A2(n22144), .B1(n15878), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n15861) );
  OAI211_X1 U18000 ( .C1(n15863), .C2(n15890), .A(n15862), .B(n15861), .ZN(
        P1_U2882) );
  AOI22_X1 U18001 ( .A1(n15877), .A2(DATAI_21_), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n15887), .ZN(n15866) );
  AOI22_X1 U18002 ( .A1(n15880), .A2(n15864), .B1(n15878), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n15865) );
  OAI211_X1 U18003 ( .C1(n15967), .C2(n15890), .A(n15866), .B(n15865), .ZN(
        P1_U2883) );
  AOI22_X1 U18004 ( .A1(n15877), .A2(DATAI_20_), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n15887), .ZN(n15869) );
  AOI22_X1 U18005 ( .A1(n15880), .A2(n15867), .B1(n15878), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n15868) );
  OAI211_X1 U18006 ( .C1(n15979), .C2(n15890), .A(n15869), .B(n15868), .ZN(
        P1_U2884) );
  AOI22_X1 U18007 ( .A1(n15877), .A2(DATAI_19_), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n15887), .ZN(n15871) );
  AOI22_X1 U18008 ( .A1(n15880), .A2(n17209), .B1(n15878), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n15870) );
  OAI211_X1 U18009 ( .C1(n15983), .C2(n15890), .A(n15871), .B(n15870), .ZN(
        P1_U2885) );
  AOI22_X1 U18010 ( .A1(n15877), .A2(DATAI_18_), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n15887), .ZN(n15874) );
  AOI22_X1 U18011 ( .A1(n15880), .A2(n15872), .B1(n15878), .B2(
        BUF1_REG_18__SCAN_IN), .ZN(n15873) );
  OAI211_X1 U18012 ( .C1(n21572), .C2(n15890), .A(n15874), .B(n15873), .ZN(
        P1_U2886) );
  AOI22_X1 U18013 ( .A1(n15877), .A2(DATAI_17_), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n15887), .ZN(n15876) );
  AOI22_X1 U18014 ( .A1(n15880), .A2(n16177), .B1(n15878), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n15875) );
  OAI211_X1 U18015 ( .C1(n21550), .C2(n15890), .A(n15876), .B(n15875), .ZN(
        P1_U2887) );
  AOI22_X1 U18016 ( .A1(n15877), .A2(DATAI_16_), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n15887), .ZN(n15882) );
  INV_X1 U18017 ( .A(n21675), .ZN(n15879) );
  AOI22_X1 U18018 ( .A1(n15880), .A2(n15879), .B1(n15878), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n15881) );
  OAI211_X1 U18019 ( .C1(n15883), .C2(n15890), .A(n15882), .B(n15881), .ZN(
        P1_U2888) );
  INV_X1 U18020 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n19878) );
  OAI222_X1 U18021 ( .A1(n16009), .A2(n15890), .B1(n15886), .B2(n19878), .C1(
        n15885), .C2(n15884), .ZN(P1_U2889) );
  AOI22_X1 U18022 ( .A1(n15888), .A2(n21752), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n15887), .ZN(n15889) );
  OAI21_X1 U18023 ( .B1(n15891), .B2(n15890), .A(n15889), .ZN(P1_U2891) );
  INV_X1 U18024 ( .A(n16077), .ZN(n15892) );
  NOR2_X1 U18025 ( .A1(n20009), .A2(n15892), .ZN(n15893) );
  AND2_X1 U18026 ( .A1(n16078), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16046) );
  MUX2_X1 U18027 ( .A(n15893), .B(n16046), .S(n15917), .Z(n15895) );
  NAND2_X1 U18028 ( .A1(n15895), .A2(n15894), .ZN(n15896) );
  XNOR2_X1 U18029 ( .A(n15896), .B(n16048), .ZN(n16066) );
  NOR2_X1 U18030 ( .A1(n21378), .A2(n17089), .ZN(n16058) );
  AOI21_X1 U18031 ( .B1(n20015), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n16058), .ZN(n15897) );
  OAI21_X1 U18032 ( .B1(n20025), .B2(n15898), .A(n15897), .ZN(n15899) );
  AOI21_X1 U18033 ( .B1(n15900), .B2(n20021), .A(n15899), .ZN(n15901) );
  OAI21_X1 U18034 ( .B1(n16066), .B2(n21578), .A(n15901), .ZN(P1_U2969) );
  INV_X1 U18035 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n17192) );
  NOR2_X1 U18036 ( .A1(n21378), .A2(n17192), .ZN(n16080) );
  NOR2_X1 U18037 ( .A1(n20025), .A2(n15902), .ZN(n15903) );
  AOI211_X1 U18038 ( .C1(n20015), .C2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16080), .B(n15903), .ZN(n15914) );
  NAND3_X1 U18039 ( .A1(n15904), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n15905), .ZN(n15908) );
  OR3_X1 U18040 ( .A1(n15904), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n15906), .ZN(n15907) );
  NAND2_X1 U18041 ( .A1(n15908), .A2(n15907), .ZN(n15911) );
  INV_X1 U18042 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15909) );
  MUX2_X1 U18043 ( .A(n15909), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n20009), .Z(n15910) );
  NAND2_X1 U18044 ( .A1(n15911), .A2(n15910), .ZN(n15912) );
  XNOR2_X1 U18045 ( .A(n15912), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16076) );
  NAND2_X1 U18046 ( .A1(n16076), .A2(n20020), .ZN(n15913) );
  OAI211_X1 U18047 ( .C1(n15915), .C2(n19957), .A(n15914), .B(n15913), .ZN(
        P1_U2971) );
  XNOR2_X1 U18048 ( .A(n20009), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15916) );
  XNOR2_X1 U18049 ( .A(n15917), .B(n15916), .ZN(n16091) );
  NAND2_X1 U18050 ( .A1(n21390), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n16084) );
  OAI21_X1 U18051 ( .B1(n19983), .B2(n15918), .A(n16084), .ZN(n15921) );
  NOR2_X1 U18052 ( .A1(n15919), .A2(n19957), .ZN(n15920) );
  OAI21_X1 U18053 ( .B1(n16091), .B2(n21578), .A(n15923), .ZN(P1_U2972) );
  XOR2_X1 U18054 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n15924), .Z(
        n16100) );
  NOR2_X1 U18055 ( .A1(n21378), .A2(n16981), .ZN(n16095) );
  AOI21_X1 U18056 ( .B1(n20015), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16095), .ZN(n15925) );
  OAI21_X1 U18057 ( .B1(n20025), .B2(n15926), .A(n15925), .ZN(n15927) );
  AOI21_X1 U18058 ( .B1(n15928), .B2(n20021), .A(n15927), .ZN(n15929) );
  OAI21_X1 U18059 ( .B1(n21578), .B2(n16100), .A(n15929), .ZN(P1_U2973) );
  NOR2_X1 U18060 ( .A1(n21378), .A2(n17085), .ZN(n16102) );
  NOR2_X1 U18061 ( .A1(n19983), .A2(n15930), .ZN(n15931) );
  AOI211_X1 U18062 ( .C1(n20000), .C2(n15932), .A(n16102), .B(n15931), .ZN(
        n15937) );
  NOR2_X1 U18063 ( .A1(n15904), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15934) );
  NAND2_X1 U18064 ( .A1(n19975), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15947) );
  OAI211_X1 U18065 ( .C1(n15934), .C2(n16105), .A(n15947), .B(n15933), .ZN(
        n15935) );
  XNOR2_X1 U18066 ( .A(n15935), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n16101) );
  NAND2_X1 U18067 ( .A1(n16101), .A2(n20020), .ZN(n15936) );
  OAI211_X1 U18068 ( .C1(n15938), .C2(n19957), .A(n15937), .B(n15936), .ZN(
        P1_U2974) );
  OR2_X1 U18069 ( .A1(n15904), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15940) );
  NAND2_X1 U18070 ( .A1(n15904), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15939) );
  MUX2_X1 U18071 ( .A(n15940), .B(n15939), .S(n20009), .Z(n15941) );
  XNOR2_X1 U18072 ( .A(n15941), .B(n16118), .ZN(n16126) );
  NOR2_X1 U18073 ( .A1(n21378), .A2(n16983), .ZN(n16117) );
  AOI21_X1 U18074 ( .B1(n20015), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16117), .ZN(n15942) );
  OAI21_X1 U18075 ( .B1(n20025), .B2(n15943), .A(n15942), .ZN(n15944) );
  AOI21_X1 U18076 ( .B1(n15945), .B2(n20021), .A(n15944), .ZN(n15946) );
  OAI21_X1 U18077 ( .B1(n21578), .B2(n16126), .A(n15946), .ZN(P1_U2975) );
  OAI21_X1 U18078 ( .B1(n19975), .B2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15947), .ZN(n15948) );
  XOR2_X1 U18079 ( .A(n15948), .B(n15904), .Z(n21392) );
  OAI22_X1 U18080 ( .A1(n19983), .A2(n15949), .B1(n21378), .B2(n17086), .ZN(
        n15952) );
  NOR2_X1 U18081 ( .A1(n15950), .A2(n19957), .ZN(n15951) );
  AOI211_X1 U18082 ( .C1(n20000), .C2(n15953), .A(n15952), .B(n15951), .ZN(
        n15954) );
  OAI21_X1 U18083 ( .B1(n21392), .B2(n21578), .A(n15954), .ZN(P1_U2976) );
  NAND2_X1 U18084 ( .A1(n15956), .A2(n15955), .ZN(n15957) );
  XOR2_X1 U18085 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n15957), .Z(
        n21380) );
  NOR2_X1 U18086 ( .A1(n21378), .A2(n17081), .ZN(n21383) );
  AOI21_X1 U18087 ( .B1(n20015), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n21383), .ZN(n15958) );
  OAI21_X1 U18088 ( .B1(n20025), .B2(n15959), .A(n15958), .ZN(n15960) );
  AOI21_X1 U18089 ( .B1(n15961), .B2(n20021), .A(n15960), .ZN(n15962) );
  OAI21_X1 U18090 ( .B1(n21578), .B2(n21380), .A(n15962), .ZN(P1_U2977) );
  XNOR2_X1 U18091 ( .A(n20009), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n20017) );
  NAND2_X1 U18092 ( .A1(n20018), .A2(n20017), .ZN(n20016) );
  OAI21_X1 U18093 ( .B1(n21343), .B2(n20009), .A(n20016), .ZN(n15981) );
  AOI22_X1 U18094 ( .A1(n15981), .A2(n21373), .B1(n20009), .B2(n20016), .ZN(
        n15975) );
  NAND2_X1 U18095 ( .A1(n15964), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15963) );
  OAI211_X1 U18096 ( .C1(n15964), .C2(n20009), .A(n15975), .B(n15963), .ZN(
        n15965) );
  XNOR2_X1 U18097 ( .A(n15965), .B(n16133), .ZN(n16141) );
  NAND2_X1 U18098 ( .A1(n21390), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n16137) );
  OAI21_X1 U18099 ( .B1(n19983), .B2(n15966), .A(n16137), .ZN(n15969) );
  NOR2_X1 U18100 ( .A1(n15967), .A2(n19957), .ZN(n15968) );
  AOI211_X1 U18101 ( .C1(n20000), .C2(n15970), .A(n15969), .B(n15968), .ZN(
        n15971) );
  OAI21_X1 U18102 ( .B1(n21578), .B2(n16141), .A(n15971), .ZN(P1_U2978) );
  INV_X1 U18103 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n15972) );
  NOR2_X1 U18104 ( .A1(n21378), .A2(n15972), .ZN(n16145) );
  NOR2_X1 U18105 ( .A1(n20025), .A2(n15973), .ZN(n15974) );
  AOI211_X1 U18106 ( .C1(n20015), .C2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16145), .B(n15974), .ZN(n15978) );
  OAI21_X1 U18107 ( .B1(n20009), .B2(n21373), .A(n15975), .ZN(n15976) );
  XNOR2_X1 U18108 ( .A(n15976), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n16142) );
  NAND2_X1 U18109 ( .A1(n16142), .A2(n20020), .ZN(n15977) );
  OAI211_X1 U18110 ( .C1(n15979), .C2(n19957), .A(n15978), .B(n15977), .ZN(
        P1_U2979) );
  XNOR2_X1 U18111 ( .A(n20009), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15980) );
  XNOR2_X1 U18112 ( .A(n15981), .B(n15980), .ZN(n21369) );
  OAI22_X1 U18113 ( .A1(n19983), .A2(n15982), .B1(n21378), .B2(n21379), .ZN(
        n15985) );
  NOR2_X1 U18114 ( .A1(n15983), .A2(n19957), .ZN(n15984) );
  AOI211_X1 U18115 ( .C1(n20000), .C2(n15986), .A(n15985), .B(n15984), .ZN(
        n15987) );
  OAI21_X1 U18116 ( .B1(n21369), .B2(n21578), .A(n15987), .ZN(P1_U2980) );
  INV_X1 U18117 ( .A(n21353), .ZN(n15988) );
  NAND2_X1 U18118 ( .A1(n20009), .A2(n15988), .ZN(n15992) );
  OR2_X1 U18119 ( .A1(n19974), .A2(n15989), .ZN(n19995) );
  INV_X1 U18120 ( .A(n20005), .ZN(n16001) );
  AOI211_X1 U18121 ( .C1(n19995), .C2(n16000), .A(n16001), .B(n15990), .ZN(
        n15991) );
  MUX2_X1 U18122 ( .A(n15992), .B(n20007), .S(n15991), .Z(n15993) );
  XNOR2_X1 U18123 ( .A(n15993), .B(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n21356) );
  NAND2_X1 U18124 ( .A1(n21356), .A2(n20020), .ZN(n15998) );
  INV_X1 U18125 ( .A(n21546), .ZN(n15996) );
  INV_X1 U18126 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n15994) );
  OAI22_X1 U18127 ( .A1(n19983), .A2(n21545), .B1(n21378), .B2(n15994), .ZN(
        n15995) );
  AOI21_X1 U18128 ( .B1(n20000), .B2(n15996), .A(n15995), .ZN(n15997) );
  OAI211_X1 U18129 ( .C1(n19957), .C2(n21550), .A(n15998), .B(n15997), .ZN(
        P1_U2982) );
  AOI21_X1 U18130 ( .B1(n19974), .B2(n16000), .A(n15999), .ZN(n20006) );
  NOR2_X1 U18131 ( .A1(n19975), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n20004) );
  NOR2_X1 U18132 ( .A1(n20004), .A2(n16001), .ZN(n16002) );
  XNOR2_X1 U18133 ( .A(n20006), .B(n16002), .ZN(n21329) );
  NAND2_X1 U18134 ( .A1(n21329), .A2(n20020), .ZN(n16008) );
  INV_X1 U18135 ( .A(n16003), .ZN(n16006) );
  OAI22_X1 U18136 ( .A1(n19983), .A2(n16004), .B1(n21378), .B2(n21338), .ZN(
        n16005) );
  AOI21_X1 U18137 ( .B1(n20000), .B2(n16006), .A(n16005), .ZN(n16007) );
  OAI211_X1 U18138 ( .C1(n19957), .C2(n16009), .A(n16008), .B(n16007), .ZN(
        P1_U2984) );
  INV_X1 U18139 ( .A(n19974), .ZN(n16011) );
  AOI21_X1 U18140 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n19975), .ZN(n19991) );
  OAI22_X1 U18141 ( .A1(n16011), .A2(n19991), .B1(n16010), .B2(n20009), .ZN(
        n19986) );
  INV_X1 U18142 ( .A(n16013), .ZN(n16012) );
  OAI21_X1 U18143 ( .B1(n20009), .B2(n21315), .A(n16012), .ZN(n19985) );
  NOR2_X1 U18144 ( .A1(n19986), .A2(n19985), .ZN(n19984) );
  NOR2_X1 U18145 ( .A1(n19984), .A2(n16013), .ZN(n16015) );
  XNOR2_X1 U18146 ( .A(n16015), .B(n16014), .ZN(n21262) );
  INV_X1 U18147 ( .A(n21262), .ZN(n16021) );
  AOI22_X1 U18148 ( .A1(n20015), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n21390), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n16016) );
  OAI21_X1 U18149 ( .B1(n20025), .B2(n16017), .A(n16016), .ZN(n16018) );
  AOI21_X1 U18150 ( .B1(n16019), .B2(n20021), .A(n16018), .ZN(n16020) );
  OAI21_X1 U18151 ( .B1(n16021), .B2(n21578), .A(n16020), .ZN(P1_U2986) );
  NOR2_X1 U18152 ( .A1(n16022), .A2(n21409), .ZN(n16052) );
  INV_X1 U18153 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16023) );
  NOR2_X1 U18154 ( .A1(n21381), .A2(n16023), .ZN(n16114) );
  INV_X1 U18155 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n21324) );
  NAND3_X1 U18156 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n16024), .ZN(n21311) );
  NOR3_X1 U18157 ( .A1(n21315), .A2(n21324), .A3(n21311), .ZN(n16029) );
  NAND2_X1 U18158 ( .A1(n16029), .A2(n16025), .ZN(n16040) );
  NOR2_X1 U18159 ( .A1(n21274), .A2(n21272), .ZN(n21344) );
  AND2_X1 U18160 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n21344), .ZN(
        n16026) );
  AND2_X1 U18161 ( .A1(n21348), .A2(n16026), .ZN(n16043) );
  INV_X1 U18162 ( .A(n16043), .ZN(n16027) );
  NOR2_X1 U18163 ( .A1(n16040), .A2(n16027), .ZN(n16127) );
  NAND3_X1 U18164 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n16114), .A3(
        n16127), .ZN(n16033) );
  NAND2_X1 U18165 ( .A1(n16029), .A2(n16028), .ZN(n21264) );
  INV_X1 U18166 ( .A(n21264), .ZN(n21331) );
  NAND2_X1 U18167 ( .A1(n21331), .A2(n16043), .ZN(n16030) );
  NAND2_X1 U18168 ( .A1(n21337), .A2(n16030), .ZN(n16032) );
  NAND2_X1 U18169 ( .A1(n16032), .A2(n16031), .ZN(n16129) );
  AOI21_X1 U18170 ( .B1(n16041), .B2(n16033), .A(n16129), .ZN(n16035) );
  INV_X1 U18171 ( .A(n16114), .ZN(n16044) );
  NAND2_X1 U18172 ( .A1(n21337), .A2(n16044), .ZN(n16034) );
  NAND2_X1 U18173 ( .A1(n16035), .A2(n16034), .ZN(n21391) );
  AND2_X1 U18174 ( .A1(n16130), .A2(n16045), .ZN(n16036) );
  OR2_X1 U18175 ( .A1(n21391), .A2(n16036), .ZN(n16110) );
  NOR2_X1 U18176 ( .A1(n16110), .A2(n16037), .ZN(n16056) );
  NOR3_X1 U18177 ( .A1(n21337), .A2(n16129), .A3(n16041), .ZN(n16055) );
  NOR2_X1 U18178 ( .A1(n16056), .A2(n16055), .ZN(n16089) );
  NOR2_X1 U18179 ( .A1(n16089), .A2(n16048), .ZN(n16062) );
  NOR2_X1 U18180 ( .A1(n21347), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16057) );
  NOR2_X1 U18181 ( .A1(n16057), .A2(n11310), .ZN(n16039) );
  AOI211_X1 U18182 ( .C1(n16062), .C2(n16039), .A(n16055), .B(n16038), .ZN(
        n16050) );
  OR2_X1 U18183 ( .A1(n16116), .A2(n21264), .ZN(n16042) );
  INV_X1 U18184 ( .A(n16040), .ZN(n21333) );
  NAND2_X1 U18185 ( .A1(n16041), .A2(n21333), .ZN(n16147) );
  NAND2_X1 U18186 ( .A1(n16042), .A2(n16147), .ZN(n21342) );
  NAND2_X1 U18187 ( .A1(n21342), .A2(n16043), .ZN(n21399) );
  OR2_X1 U18188 ( .A1(n21399), .A2(n16044), .ZN(n16103) );
  NOR2_X1 U18189 ( .A1(n16103), .A2(n16045), .ZN(n16092) );
  NAND2_X1 U18190 ( .A1(n16092), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16085) );
  INV_X1 U18191 ( .A(n16046), .ZN(n16047) );
  OR2_X1 U18192 ( .A1(n16085), .A2(n16047), .ZN(n16061) );
  NOR3_X1 U18193 ( .A1(n16061), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n16048), .ZN(n16049) );
  OAI21_X1 U18194 ( .B1(n16054), .B2(n21327), .A(n16053), .ZN(P1_U3000) );
  INV_X1 U18195 ( .A(n15802), .ZN(n16064) );
  AOI21_X1 U18196 ( .B1(n16056), .B2(n16078), .A(n16055), .ZN(n16070) );
  OAI21_X1 U18197 ( .B1(n16070), .B2(n16057), .A(
        P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16060) );
  INV_X1 U18198 ( .A(n16058), .ZN(n16059) );
  OAI211_X1 U18199 ( .C1(n16062), .C2(n16061), .A(n16060), .B(n16059), .ZN(
        n16063) );
  AOI21_X1 U18200 ( .B1(n16064), .B2(n21394), .A(n16063), .ZN(n16065) );
  OAI21_X1 U18201 ( .B1(n16066), .B2(n21327), .A(n16065), .ZN(P1_U3001) );
  INV_X1 U18202 ( .A(n16067), .ZN(n16069) );
  NOR3_X1 U18203 ( .A1(n16085), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11310), .ZN(n16068) );
  AOI211_X1 U18204 ( .C1(n16070), .C2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n16069), .B(n16068), .ZN(n16073) );
  NAND2_X1 U18205 ( .A1(n16071), .A2(n21394), .ZN(n16072) );
  OAI211_X1 U18206 ( .C1(n16074), .C2(n21327), .A(n16073), .B(n16072), .ZN(
        P1_U3002) );
  INV_X1 U18207 ( .A(n16075), .ZN(n16083) );
  NAND2_X1 U18208 ( .A1(n16076), .A2(n21406), .ZN(n16082) );
  NOR3_X1 U18209 ( .A1(n16085), .A2(n16078), .A3(n16077), .ZN(n16079) );
  AOI211_X1 U18210 ( .C1(n16089), .C2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n16080), .B(n16079), .ZN(n16081) );
  OAI211_X1 U18211 ( .C1(n21409), .C2(n16083), .A(n16082), .B(n16081), .ZN(
        P1_U3003) );
  OAI21_X1 U18212 ( .B1(n16085), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16084), .ZN(n16088) );
  NOR2_X1 U18213 ( .A1(n16086), .A2(n21409), .ZN(n16087) );
  AOI211_X1 U18214 ( .C1(n16089), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16088), .B(n16087), .ZN(n16090) );
  OAI21_X1 U18215 ( .B1(n16091), .B2(n21327), .A(n16090), .ZN(P1_U3004) );
  INV_X1 U18216 ( .A(n16092), .ZN(n16093) );
  NOR2_X1 U18217 ( .A1(n16093), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n16094) );
  AOI211_X1 U18218 ( .C1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n16110), .A(
        n16095), .B(n16094), .ZN(n16099) );
  INV_X1 U18219 ( .A(n16096), .ZN(n16097) );
  NAND2_X1 U18220 ( .A1(n16097), .A2(n21394), .ZN(n16098) );
  OAI211_X1 U18221 ( .C1(n16100), .C2(n21327), .A(n16099), .B(n16098), .ZN(
        P1_U3005) );
  INV_X1 U18222 ( .A(n16101), .ZN(n16112) );
  INV_X1 U18223 ( .A(n16102), .ZN(n16107) );
  INV_X1 U18224 ( .A(n16103), .ZN(n16119) );
  NAND3_X1 U18225 ( .A1(n16119), .A2(n16105), .A3(n16104), .ZN(n16106) );
  OAI211_X1 U18226 ( .C1(n16108), .C2(n21409), .A(n16107), .B(n16106), .ZN(
        n16109) );
  AOI21_X1 U18227 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n16110), .A(
        n16109), .ZN(n16111) );
  OAI21_X1 U18228 ( .B1(n16112), .B2(n21327), .A(n16111), .ZN(P1_U3006) );
  NAND2_X1 U18229 ( .A1(n16114), .A2(n16113), .ZN(n21398) );
  INV_X1 U18230 ( .A(n21391), .ZN(n16115) );
  OAI21_X1 U18231 ( .B1(n16116), .B2(n21398), .A(n16115), .ZN(n16124) );
  INV_X1 U18232 ( .A(n16117), .ZN(n16121) );
  NAND3_X1 U18233 ( .A1(n16119), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n16118), .ZN(n16120) );
  OAI211_X1 U18234 ( .C1(n16122), .C2(n21409), .A(n16121), .B(n16120), .ZN(
        n16123) );
  AOI21_X1 U18235 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n16124), .A(
        n16123), .ZN(n16125) );
  OAI21_X1 U18236 ( .B1(n16126), .B2(n21327), .A(n16125), .ZN(P1_U3007) );
  NOR2_X1 U18237 ( .A1(n21332), .A2(n16127), .ZN(n16128) );
  OR2_X1 U18238 ( .A1(n16129), .A2(n16128), .ZN(n21375) );
  INV_X1 U18239 ( .A(n16134), .ZN(n16131) );
  OAI22_X1 U18240 ( .A1(n21375), .A2(n16131), .B1(n16130), .B2(n21334), .ZN(
        n16132) );
  INV_X1 U18241 ( .A(n16132), .ZN(n21386) );
  NAND2_X1 U18242 ( .A1(n16134), .A2(n16133), .ZN(n16135) );
  NOR2_X1 U18243 ( .A1(n21399), .A2(n16135), .ZN(n21385) );
  INV_X1 U18244 ( .A(n16136), .ZN(n16138) );
  OAI21_X1 U18245 ( .B1(n16138), .B2(n21409), .A(n16137), .ZN(n16139) );
  AOI211_X1 U18246 ( .C1(n21386), .C2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n21385), .B(n16139), .ZN(n16140) );
  OAI21_X1 U18247 ( .B1(n16141), .B2(n21327), .A(n16140), .ZN(P1_U3010) );
  INV_X1 U18248 ( .A(n16142), .ZN(n16153) );
  INV_X1 U18249 ( .A(n16143), .ZN(n16146) );
  NOR3_X1 U18250 ( .A1(n21399), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n21373), .ZN(n16144) );
  AOI211_X1 U18251 ( .C1(n21394), .C2(n16146), .A(n16145), .B(n16144), .ZN(
        n16152) );
  NAND2_X1 U18252 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21265), .ZN(
        n16148) );
  OAI21_X1 U18253 ( .B1(n21264), .B2(n16148), .A(n16147), .ZN(n21271) );
  INV_X1 U18254 ( .A(n21271), .ZN(n16149) );
  AOI21_X1 U18255 ( .B1(n16149), .B2(n21402), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16150) );
  OAI21_X1 U18256 ( .B1(n16150), .B2(n21375), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n16151) );
  OAI211_X1 U18257 ( .C1(n16153), .C2(n21327), .A(n16152), .B(n16151), .ZN(
        P1_U3011) );
  NOR2_X1 U18258 ( .A1(n14911), .A2(n16154), .ZN(n21819) );
  NAND2_X1 U18259 ( .A1(n21851), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n21857) );
  INV_X1 U18260 ( .A(n21769), .ZN(n16155) );
  OAI211_X1 U18261 ( .C1(n14911), .C2(n21802), .A(n16155), .B(n21925), .ZN(
        n16157) );
  NAND2_X1 U18262 ( .A1(n21771), .A2(n21580), .ZN(n16156) );
  OAI211_X1 U18263 ( .C1(n21857), .C2(n21919), .A(n16157), .B(n16156), .ZN(
        n16158) );
  MUX2_X1 U18264 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n16158), .S(
        n16976), .Z(P1_U3475) );
  NOR2_X1 U18265 ( .A1(n14900), .A2(n14730), .ZN(n16160) );
  AOI22_X1 U18266 ( .A1(n16162), .A2(n16161), .B1(n16160), .B2(n16159), .ZN(
        n16163) );
  OAI21_X1 U18267 ( .B1(n14906), .B2(n16164), .A(n16163), .ZN(n16950) );
  INV_X1 U18268 ( .A(n16950), .ZN(n16948) );
  NAND2_X1 U18269 ( .A1(n16166), .A2(n16165), .ZN(n16170) );
  INV_X1 U18270 ( .A(n14900), .ZN(n16168) );
  INV_X1 U18271 ( .A(n14730), .ZN(n16167) );
  NAND3_X1 U18272 ( .A1(n16168), .A2(n21597), .A3(n16167), .ZN(n16169) );
  OAI211_X1 U18273 ( .C1(n16948), .C2(n16171), .A(n16170), .B(n16169), .ZN(
        n16173) );
  MUX2_X1 U18274 ( .A(n16173), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n16172), .Z(P1_U3473) );
  NAND2_X1 U18275 ( .A1(n22202), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n16182) );
  NOR2_X2 U18276 ( .A1(n16175), .A2(n16174), .ZN(n21984) );
  INV_X1 U18277 ( .A(n16176), .ZN(n22197) );
  NAND2_X1 U18278 ( .A1(n22145), .A2(n16177), .ZN(n21980) );
  AOI22_X1 U18279 ( .A1(n21984), .A2(n22197), .B1(n22199), .B2(n21983), .ZN(
        n16181) );
  INV_X1 U18280 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20075) );
  INV_X1 U18281 ( .A(DATAI_25_), .ZN(n16178) );
  NAND2_X1 U18282 ( .A1(n16191), .A2(n21985), .ZN(n16180) );
  INV_X1 U18283 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n20060) );
  INV_X1 U18284 ( .A(DATAI_17_), .ZN(n16993) );
  OAI22_X1 U18285 ( .A1(n20060), .A2(n22152), .B1(n16993), .B2(n22150), .ZN(
        n21977) );
  NAND2_X1 U18286 ( .A1(n22207), .A2(n21977), .ZN(n16179) );
  NAND4_X1 U18287 ( .A1(n16182), .A2(n16181), .A3(n16180), .A4(n16179), .ZN(
        P1_U3154) );
  NAND2_X1 U18288 ( .A1(n22202), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n16186) );
  AOI22_X1 U18289 ( .A1(n22023), .A2(n22197), .B1(n22199), .B2(n22022), .ZN(
        n16185) );
  NAND2_X1 U18290 ( .A1(n16191), .A2(n22024), .ZN(n16184) );
  NAND2_X1 U18291 ( .A1(n22207), .A2(n22016), .ZN(n16183) );
  NAND4_X1 U18292 ( .A1(n16186), .A2(n16185), .A3(n16184), .A4(n16183), .ZN(
        P1_U3155) );
  NAND2_X1 U18293 ( .A1(n22202), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n16190) );
  AOI22_X1 U18294 ( .A1(n22061), .A2(n22197), .B1(n22199), .B2(n22060), .ZN(
        n16189) );
  NAND2_X1 U18295 ( .A1(n16191), .A2(n22062), .ZN(n16188) );
  NAND2_X1 U18296 ( .A1(n22207), .A2(n22054), .ZN(n16187) );
  NAND4_X1 U18297 ( .A1(n16190), .A2(n16189), .A3(n16188), .A4(n16187), .ZN(
        P1_U3156) );
  NAND2_X1 U18298 ( .A1(n22202), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n16195) );
  AOI22_X1 U18299 ( .A1(n22139), .A2(n22197), .B1(n22199), .B2(n22138), .ZN(
        n16194) );
  NAND2_X1 U18300 ( .A1(n16191), .A2(n22140), .ZN(n16193) );
  NAND2_X1 U18301 ( .A1(n22207), .A2(n22132), .ZN(n16192) );
  NAND4_X1 U18302 ( .A1(n16195), .A2(n16194), .A3(n16193), .A4(n16192), .ZN(
        P1_U3158) );
  MUX2_X1 U18303 ( .A(P2_EBX_REG_31__SCAN_IN), .B(n16196), .S(n16209), .Z(
        P2_U2856) );
  XOR2_X1 U18304 ( .A(n16198), .B(n16197), .Z(n16199) );
  XNOR2_X1 U18305 ( .A(n16200), .B(n16199), .ZN(n16289) );
  NAND2_X1 U18306 ( .A1(n16267), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n16202) );
  NAND2_X1 U18307 ( .A1(n18541), .A2(n16209), .ZN(n16201) );
  OAI211_X1 U18308 ( .C1(n16289), .C2(n16278), .A(n16202), .B(n16201), .ZN(
        P2_U2858) );
  NOR2_X1 U18309 ( .A1(n11026), .A2(n16203), .ZN(n16205) );
  XNOR2_X1 U18310 ( .A(n16205), .B(n16204), .ZN(n16297) );
  NAND2_X1 U18311 ( .A1(n16267), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n16211) );
  OR2_X1 U18312 ( .A1(n16206), .A2(n16207), .ZN(n16208) );
  NAND2_X1 U18313 ( .A1(n18526), .A2(n16209), .ZN(n16210) );
  OAI211_X1 U18314 ( .C1(n16297), .C2(n16278), .A(n16211), .B(n16210), .ZN(
        P2_U2859) );
  NOR2_X1 U18315 ( .A1(n16213), .A2(n11026), .ZN(n16214) );
  XOR2_X1 U18316 ( .A(n16215), .B(n16214), .Z(n16307) );
  NOR2_X1 U18317 ( .A1(n16216), .A2(n16217), .ZN(n16218) );
  OR2_X1 U18318 ( .A1(n16206), .A2(n16218), .ZN(n16609) );
  NOR2_X1 U18319 ( .A1(n16609), .A2(n16267), .ZN(n16219) );
  AOI21_X1 U18320 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n16267), .A(n16219), .ZN(
        n16220) );
  OAI21_X1 U18321 ( .B1(n16307), .B2(n16278), .A(n16220), .ZN(P2_U2860) );
  OAI21_X1 U18322 ( .B1(n16223), .B2(n16222), .A(n16221), .ZN(n16313) );
  AND2_X1 U18323 ( .A1(n16229), .A2(n16224), .ZN(n16225) );
  OR2_X1 U18324 ( .A1(n16225), .A2(n16216), .ZN(n18500) );
  NOR2_X1 U18325 ( .A1(n18500), .A2(n16267), .ZN(n16226) );
  AOI21_X1 U18326 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n16267), .A(n16226), .ZN(
        n16227) );
  OAI21_X1 U18327 ( .B1(n16313), .B2(n16278), .A(n16227), .ZN(P2_U2861) );
  INV_X1 U18328 ( .A(n16229), .ZN(n16230) );
  AOI21_X1 U18329 ( .B1(n16231), .B2(n16228), .A(n16230), .ZN(n18490) );
  INV_X1 U18330 ( .A(n18490), .ZN(n16634) );
  AOI21_X1 U18331 ( .B1(n16234), .B2(n16233), .A(n16232), .ZN(n16321) );
  NAND2_X1 U18332 ( .A1(n16321), .A2(n16252), .ZN(n16236) );
  NAND2_X1 U18333 ( .A1(n16267), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n16235) );
  OAI211_X1 U18334 ( .C1(n16634), .C2(n16267), .A(n16236), .B(n16235), .ZN(
        P2_U2862) );
  OAI21_X1 U18335 ( .B1(n16237), .B2(n16238), .A(n16228), .ZN(n18480) );
  AOI21_X1 U18336 ( .B1(n16240), .B2(n16239), .A(n14280), .ZN(n16328) );
  NAND2_X1 U18337 ( .A1(n16328), .A2(n16252), .ZN(n16242) );
  NAND2_X1 U18338 ( .A1(n16267), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n16241) );
  OAI211_X1 U18339 ( .C1(n18480), .C2(n16267), .A(n16242), .B(n16241), .ZN(
        P2_U2863) );
  XNOR2_X1 U18340 ( .A(n11042), .B(n16243), .ZN(n16338) );
  AND2_X1 U18341 ( .A1(n16250), .A2(n16244), .ZN(n16245) );
  OR2_X1 U18342 ( .A1(n16245), .A2(n16237), .ZN(n16652) );
  NOR2_X1 U18343 ( .A1(n16652), .A2(n16267), .ZN(n16246) );
  AOI21_X1 U18344 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n16267), .A(n16246), .ZN(
        n16247) );
  OAI21_X1 U18345 ( .B1(n16338), .B2(n16278), .A(n16247), .ZN(P2_U2864) );
  NAND2_X1 U18346 ( .A1(n16255), .A2(n16248), .ZN(n16249) );
  AND2_X1 U18347 ( .A1(n16250), .A2(n16249), .ZN(n18459) );
  INV_X1 U18348 ( .A(n18459), .ZN(n16672) );
  AOI21_X1 U18349 ( .B1(n16251), .B2(n15548), .A(n11042), .ZN(n19344) );
  NAND2_X1 U18350 ( .A1(n19344), .A2(n16252), .ZN(n16254) );
  NAND2_X1 U18351 ( .A1(n16267), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n16253) );
  OAI211_X1 U18352 ( .C1(n16672), .C2(n16267), .A(n16254), .B(n16253), .ZN(
        P2_U2865) );
  INV_X1 U18353 ( .A(n16255), .ZN(n16256) );
  AOI21_X1 U18354 ( .B1(n16257), .B2(n15561), .A(n16256), .ZN(n18450) );
  INV_X1 U18355 ( .A(n18450), .ZN(n16683) );
  NOR2_X1 U18356 ( .A1(n16683), .A2(n16267), .ZN(n16258) );
  AOI21_X1 U18357 ( .B1(P2_EBX_REG_21__SCAN_IN), .B2(n16267), .A(n16258), .ZN(
        n16259) );
  OAI21_X1 U18358 ( .B1(n16260), .B2(n16278), .A(n16259), .ZN(P2_U2866) );
  AND2_X1 U18359 ( .A1(n16262), .A2(n16261), .ZN(n16270) );
  OAI21_X1 U18360 ( .B1(n16270), .B2(n16263), .A(n15504), .ZN(n16346) );
  NAND2_X1 U18361 ( .A1(n16267), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n16269) );
  NAND2_X1 U18362 ( .A1(n16264), .A2(n16265), .ZN(n16266) );
  NAND2_X1 U18363 ( .A1(n10963), .A2(n16266), .ZN(n18418) );
  OR2_X1 U18364 ( .A1(n18418), .A2(n16267), .ZN(n16268) );
  OAI211_X1 U18365 ( .C1(n16346), .C2(n16278), .A(n16269), .B(n16268), .ZN(
        P2_U2869) );
  INV_X1 U18366 ( .A(n16270), .ZN(n16271) );
  OAI21_X1 U18367 ( .B1(n16273), .B2(n16272), .A(n16271), .ZN(n16355) );
  OR2_X1 U18368 ( .A1(n15500), .A2(n16274), .ZN(n16275) );
  NAND2_X1 U18369 ( .A1(n16264), .A2(n16275), .ZN(n18406) );
  NOR2_X1 U18370 ( .A1(n18406), .A2(n16267), .ZN(n16276) );
  AOI21_X1 U18371 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n16267), .A(n16276), .ZN(
        n16277) );
  OAI21_X1 U18372 ( .B1(n16355), .B2(n16278), .A(n16277), .ZN(P2_U2870) );
  INV_X1 U18373 ( .A(n19674), .ZN(n16284) );
  INV_X1 U18374 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n16283) );
  INV_X1 U18375 ( .A(n16279), .ZN(n16280) );
  AOI22_X1 U18376 ( .A1(n16280), .A2(n19612), .B1(P2_EAX_REG_31__SCAN_IN), 
        .B2(n19670), .ZN(n16282) );
  NAND2_X1 U18377 ( .A1(n19673), .A2(BUF1_REG_31__SCAN_IN), .ZN(n16281) );
  OAI211_X1 U18378 ( .C1(n16284), .C2(n16283), .A(n16282), .B(n16281), .ZN(
        P2_U2888) );
  AOI22_X1 U18379 ( .A1(n19673), .A2(BUF1_REG_29__SCAN_IN), .B1(n19674), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n16286) );
  AOI22_X1 U18380 ( .A1(n19612), .A2(n18540), .B1(n19670), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n16285) );
  OAI211_X1 U18381 ( .C1(n19162), .C2(n16352), .A(n16286), .B(n16285), .ZN(
        n16287) );
  INV_X1 U18382 ( .A(n16287), .ZN(n16288) );
  OAI21_X1 U18383 ( .B1(n16289), .B2(n19677), .A(n16288), .ZN(P2_U2890) );
  INV_X1 U18384 ( .A(n16290), .ZN(n16291) );
  AOI21_X1 U18385 ( .B1(n16292), .B2(n16301), .A(n16291), .ZN(n18525) );
  INV_X1 U18386 ( .A(n18525), .ZN(n16293) );
  OAI22_X1 U18387 ( .A1(n16293), .A2(n19676), .B1(n19508), .B2(n14776), .ZN(
        n16294) );
  AOI21_X1 U18388 ( .B1(n19672), .B2(n19165), .A(n16294), .ZN(n16296) );
  AOI22_X1 U18389 ( .A1(n19673), .A2(BUF1_REG_28__SCAN_IN), .B1(n19674), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n16295) );
  OAI211_X1 U18390 ( .C1(n16297), .C2(n19677), .A(n16296), .B(n16295), .ZN(
        P2_U2891) );
  AOI22_X1 U18391 ( .A1(n19673), .A2(BUF1_REG_27__SCAN_IN), .B1(n19674), .B2(
        BUF2_REG_27__SCAN_IN), .ZN(n16304) );
  NAND2_X1 U18392 ( .A1(n16298), .A2(n16299), .ZN(n16300) );
  NAND2_X1 U18393 ( .A1(n16301), .A2(n16300), .ZN(n18522) );
  INV_X1 U18394 ( .A(n18522), .ZN(n16302) );
  AOI22_X1 U18395 ( .A1(n19612), .A2(n16302), .B1(n19670), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n16303) );
  OAI211_X1 U18396 ( .C1(n19169), .C2(n16352), .A(n16304), .B(n16303), .ZN(
        n16305) );
  INV_X1 U18397 ( .A(n16305), .ZN(n16306) );
  OAI21_X1 U18398 ( .B1(n16307), .B2(n19677), .A(n16306), .ZN(P2_U2892) );
  OAI21_X1 U18399 ( .B1(n16309), .B2(n16308), .A(n16298), .ZN(n16620) );
  OAI22_X1 U18400 ( .A1(n19676), .A2(n16620), .B1(n19508), .B2(n14774), .ZN(
        n16310) );
  AOI21_X1 U18401 ( .B1(n19672), .B2(n19172), .A(n16310), .ZN(n16312) );
  AOI22_X1 U18402 ( .A1(n19673), .A2(BUF1_REG_26__SCAN_IN), .B1(n19674), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n16311) );
  OAI211_X1 U18403 ( .C1(n16313), .C2(n19677), .A(n16312), .B(n16311), .ZN(
        P2_U2893) );
  INV_X1 U18404 ( .A(n19176), .ZN(n16319) );
  AOI22_X1 U18405 ( .A1(n19673), .A2(BUF1_REG_25__SCAN_IN), .B1(n19674), .B2(
        BUF2_REG_25__SCAN_IN), .ZN(n16318) );
  INV_X1 U18406 ( .A(n16315), .ZN(n16316) );
  XNOR2_X1 U18407 ( .A(n16314), .B(n16316), .ZN(n18491) );
  AOI22_X1 U18408 ( .A1(n19612), .A2(n18491), .B1(n19670), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n16317) );
  OAI211_X1 U18409 ( .C1(n16319), .C2(n16352), .A(n16318), .B(n16317), .ZN(
        n16320) );
  AOI21_X1 U18410 ( .B1(n16321), .B2(n19561), .A(n16320), .ZN(n16322) );
  INV_X1 U18411 ( .A(n16322), .ZN(P2_U2894) );
  AOI22_X1 U18412 ( .A1(n19673), .A2(BUF1_REG_24__SCAN_IN), .B1(n19674), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n16326) );
  AND2_X1 U18413 ( .A1(n16332), .A2(n16323), .ZN(n16324) );
  AOI22_X1 U18414 ( .A1(n19612), .A2(n11367), .B1(n19670), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n16325) );
  OAI211_X1 U18415 ( .C1(n19182), .C2(n16352), .A(n16326), .B(n16325), .ZN(
        n16327) );
  AOI21_X1 U18416 ( .B1(n16328), .B2(n19561), .A(n16327), .ZN(n16329) );
  INV_X1 U18417 ( .A(n16329), .ZN(P2_U2895) );
  INV_X1 U18418 ( .A(n19183), .ZN(n16335) );
  OR2_X1 U18419 ( .A1(n16330), .A2(n16668), .ZN(n16331) );
  NAND2_X1 U18420 ( .A1(n16332), .A2(n16331), .ZN(n18478) );
  OAI22_X1 U18421 ( .A1(n19676), .A2(n18478), .B1(n16333), .B2(n19508), .ZN(
        n16334) );
  AOI21_X1 U18422 ( .B1(n19672), .B2(n16335), .A(n16334), .ZN(n16337) );
  AOI22_X1 U18423 ( .A1(n19673), .A2(BUF1_REG_23__SCAN_IN), .B1(n19674), .B2(
        BUF2_REG_23__SCAN_IN), .ZN(n16336) );
  OAI211_X1 U18424 ( .C1(n16338), .C2(n19677), .A(n16337), .B(n16336), .ZN(
        P2_U2896) );
  AOI22_X1 U18425 ( .A1(n19673), .A2(BUF1_REG_18__SCAN_IN), .B1(n19674), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n16343) );
  XNOR2_X1 U18426 ( .A(n16339), .B(n16340), .ZN(n18419) );
  INV_X1 U18427 ( .A(n18419), .ZN(n16341) );
  AOI22_X1 U18428 ( .A1(n19612), .A2(n16341), .B1(n19670), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16342) );
  OAI211_X1 U18429 ( .C1(n19565), .C2(n16352), .A(n16343), .B(n16342), .ZN(
        n16344) );
  INV_X1 U18430 ( .A(n16344), .ZN(n16345) );
  OAI21_X1 U18431 ( .B1(n16346), .B2(n19677), .A(n16345), .ZN(P2_U2901) );
  AOI22_X1 U18432 ( .A1(n19673), .A2(BUF1_REG_17__SCAN_IN), .B1(n19674), .B2(
        BUF2_REG_17__SCAN_IN), .ZN(n16351) );
  OR2_X1 U18433 ( .A1(n16347), .A2(n16348), .ZN(n16349) );
  NAND2_X1 U18434 ( .A1(n16339), .A2(n16349), .ZN(n18407) );
  INV_X1 U18435 ( .A(n18407), .ZN(n16729) );
  AOI22_X1 U18436 ( .A1(n19612), .A2(n16729), .B1(n19670), .B2(
        P2_EAX_REG_17__SCAN_IN), .ZN(n16350) );
  OAI211_X1 U18437 ( .C1(n19620), .C2(n16352), .A(n16351), .B(n16350), .ZN(
        n16353) );
  INV_X1 U18438 ( .A(n16353), .ZN(n16354) );
  OAI21_X1 U18439 ( .B1(n16355), .B2(n19677), .A(n16354), .ZN(P2_U2902) );
  NAND2_X1 U18440 ( .A1(n16356), .A2(n17256), .ZN(n16363) );
  NAND2_X1 U18441 ( .A1(n16357), .A2(n17216), .ZN(n16359) );
  OAI211_X1 U18442 ( .C1(n17222), .C2(n16360), .A(n16359), .B(n16358), .ZN(
        n16361) );
  AOI21_X1 U18443 ( .B1(n18541), .B2(n17257), .A(n16361), .ZN(n16362) );
  OAI211_X1 U18444 ( .C1(n16364), .C2(n17228), .A(n16363), .B(n16362), .ZN(
        P2_U2985) );
  XNOR2_X1 U18445 ( .A(n16378), .B(n16365), .ZN(n16607) );
  INV_X1 U18446 ( .A(n16368), .ZN(n16367) );
  NOR2_X1 U18447 ( .A1(n11028), .A2(n16367), .ZN(n16380) );
  NOR2_X1 U18448 ( .A1(n16380), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16379) );
  NOR2_X1 U18449 ( .A1(n16394), .A2(n16368), .ZN(n16382) );
  NOR2_X1 U18450 ( .A1(n16379), .A2(n16382), .ZN(n16371) );
  XNOR2_X1 U18451 ( .A(n16369), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16370) );
  XNOR2_X1 U18452 ( .A(n16371), .B(n16370), .ZN(n16605) );
  NAND2_X1 U18453 ( .A1(n18526), .A2(n17257), .ZN(n16374) );
  NOR2_X1 U18454 ( .A1(n18583), .A2(n16372), .ZN(n16598) );
  AOI21_X1 U18455 ( .B1(n17245), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n16598), .ZN(n16373) );
  OAI211_X1 U18456 ( .C1(n17261), .C2(n18529), .A(n16374), .B(n16373), .ZN(
        n16375) );
  AOI21_X1 U18457 ( .B1(n16605), .B2(n17258), .A(n16375), .ZN(n16376) );
  OAI21_X1 U18458 ( .B1(n16377), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n16378), .ZN(n16619) );
  INV_X1 U18459 ( .A(n16379), .ZN(n16384) );
  OAI21_X1 U18460 ( .B1(n16380), .B2(n16382), .A(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n16383) );
  AOI22_X1 U18461 ( .A1(n16384), .A2(n16383), .B1(n16382), .B2(n16381), .ZN(
        n16608) );
  NAND2_X1 U18462 ( .A1(n18382), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n16613) );
  OAI21_X1 U18463 ( .B1(n17222), .B2(n18512), .A(n16613), .ZN(n16385) );
  AOI21_X1 U18464 ( .B1(n16386), .B2(n17216), .A(n16385), .ZN(n16387) );
  OAI21_X1 U18465 ( .B1(n17227), .B2(n16609), .A(n16387), .ZN(n16388) );
  AOI21_X1 U18466 ( .B1(n16608), .B2(n17258), .A(n16388), .ZN(n16389) );
  OAI21_X1 U18467 ( .B1(n17224), .B2(n16619), .A(n16389), .ZN(P2_U2987) );
  NOR2_X1 U18468 ( .A1(n11006), .A2(n16637), .ZN(n16403) );
  INV_X1 U18469 ( .A(n16377), .ZN(n16390) );
  OAI21_X1 U18470 ( .B1(n16403), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n16390), .ZN(n16630) );
  INV_X1 U18471 ( .A(n16400), .ZN(n16391) );
  OAI21_X1 U18472 ( .B1(n11010), .B2(n16401), .A(n16391), .ZN(n16393) );
  MUX2_X1 U18473 ( .A(n16401), .B(n16393), .S(n16392), .Z(n16395) );
  NOR2_X1 U18474 ( .A1(n16395), .A2(n16394), .ZN(n16628) );
  NOR2_X1 U18475 ( .A1(n18582), .A2(n17335), .ZN(n16623) );
  NOR2_X1 U18476 ( .A1(n18505), .A2(n17261), .ZN(n16396) );
  AOI211_X1 U18477 ( .C1(n17245), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n16623), .B(n16396), .ZN(n16397) );
  OAI21_X1 U18478 ( .B1(n17227), .B2(n18500), .A(n16397), .ZN(n16398) );
  AOI21_X1 U18479 ( .B1(n16628), .B2(n17258), .A(n16398), .ZN(n16399) );
  OAI21_X1 U18480 ( .B1(n16630), .B2(n17224), .A(n16399), .ZN(P2_U2988) );
  NOR2_X1 U18481 ( .A1(n16401), .A2(n16400), .ZN(n16402) );
  XNOR2_X1 U18482 ( .A(n11010), .B(n16402), .ZN(n16641) );
  AOI21_X1 U18483 ( .B1(n16637), .B2(n11006), .A(n16403), .ZN(n16631) );
  NAND2_X1 U18484 ( .A1(n16631), .A2(n17256), .ZN(n16407) );
  NOR2_X1 U18485 ( .A1(n18583), .A2(n17334), .ZN(n16632) );
  AOI21_X1 U18486 ( .B1(n17245), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16632), .ZN(n16404) );
  OAI21_X1 U18487 ( .B1(n18494), .B2(n17261), .A(n16404), .ZN(n16405) );
  AOI21_X1 U18488 ( .B1(n18490), .B2(n17257), .A(n16405), .ZN(n16406) );
  OAI211_X1 U18489 ( .C1(n17228), .C2(n16641), .A(n16407), .B(n16406), .ZN(
        P2_U2989) );
  OR2_X1 U18490 ( .A1(n16463), .A2(n16655), .ZN(n16418) );
  INV_X1 U18491 ( .A(n16418), .ZN(n16409) );
  OAI21_X1 U18492 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n16409), .A(
        n11006), .ZN(n16651) );
  XOR2_X1 U18493 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n16410), .Z(
        n16411) );
  XNOR2_X1 U18494 ( .A(n16412), .B(n16411), .ZN(n16649) );
  NOR2_X1 U18495 ( .A1(n18582), .A2(n16413), .ZN(n16645) );
  NOR2_X1 U18496 ( .A1(n18480), .A2(n17227), .ZN(n16414) );
  AOI211_X1 U18497 ( .C1(n17245), .C2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n16645), .B(n16414), .ZN(n16415) );
  OAI21_X1 U18498 ( .B1(n17261), .B2(n18484), .A(n16415), .ZN(n16416) );
  AOI21_X1 U18499 ( .B1(n16649), .B2(n17258), .A(n16416), .ZN(n16417) );
  OAI21_X1 U18500 ( .B1(n16651), .B2(n17224), .A(n16417), .ZN(P2_U2990) );
  NOR2_X1 U18501 ( .A1(n16463), .A2(n16666), .ZN(n16428) );
  OAI21_X1 U18502 ( .B1(n16428), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n16418), .ZN(n16663) );
  NOR2_X1 U18503 ( .A1(n16421), .A2(n11169), .ZN(n16422) );
  XNOR2_X1 U18504 ( .A(n16419), .B(n16422), .ZN(n16661) );
  NOR2_X1 U18505 ( .A1(n18582), .A2(n16423), .ZN(n16654) );
  NOR2_X1 U18506 ( .A1(n16652), .A2(n17227), .ZN(n16424) );
  AOI211_X1 U18507 ( .C1(n17245), .C2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16654), .B(n16424), .ZN(n16425) );
  OAI21_X1 U18508 ( .B1(n17261), .B2(n18475), .A(n16425), .ZN(n16426) );
  AOI21_X1 U18509 ( .B1(n16661), .B2(n17258), .A(n16426), .ZN(n16427) );
  OAI21_X1 U18510 ( .B1(n16663), .B2(n17224), .A(n16427), .ZN(P2_U2991) );
  INV_X1 U18511 ( .A(n16428), .ZN(n16429) );
  OAI21_X1 U18512 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n11110), .A(
        n16429), .ZN(n16677) );
  XOR2_X1 U18513 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n16431), .Z(
        n16432) );
  XNOR2_X1 U18514 ( .A(n16430), .B(n16432), .ZN(n16675) );
  INV_X1 U18515 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16434) );
  OAI22_X1 U18516 ( .A1(n17222), .A2(n16434), .B1(n16433), .B2(n18583), .ZN(
        n16435) );
  AOI21_X1 U18517 ( .B1(n18459), .B2(n17257), .A(n16435), .ZN(n16436) );
  OAI21_X1 U18518 ( .B1(n18462), .B2(n17261), .A(n16436), .ZN(n16437) );
  AOI21_X1 U18519 ( .B1(n16675), .B2(n17258), .A(n16437), .ZN(n16438) );
  OAI21_X1 U18520 ( .B1(n16677), .B2(n17224), .A(n16438), .ZN(P2_U2992) );
  NAND2_X1 U18521 ( .A1(n16441), .A2(n16822), .ZN(n16575) );
  INV_X1 U18522 ( .A(n16442), .ZN(n16576) );
  INV_X1 U18523 ( .A(n17248), .ZN(n16523) );
  OR2_X1 U18524 ( .A1(n16443), .A2(n16523), .ZN(n16446) );
  AND2_X1 U18525 ( .A1(n16522), .A2(n16444), .ZN(n16445) );
  AND2_X1 U18526 ( .A1(n16503), .A2(n16502), .ZN(n16447) );
  NAND2_X1 U18527 ( .A1(n16514), .A2(n16447), .ZN(n16448) );
  NAND2_X1 U18528 ( .A1(n16448), .A2(n16504), .ZN(n16493) );
  INV_X1 U18529 ( .A(n16449), .ZN(n16452) );
  INV_X1 U18530 ( .A(n16450), .ZN(n16451) );
  AOI22_X1 U18531 ( .A1(n16471), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n16454), .B2(n16453), .ZN(n16459) );
  INV_X1 U18532 ( .A(n16455), .ZN(n16457) );
  NAND2_X1 U18533 ( .A1(n16457), .A2(n16456), .ZN(n16458) );
  XNOR2_X1 U18534 ( .A(n16459), .B(n16458), .ZN(n16689) );
  NAND2_X1 U18535 ( .A1(n18450), .A2(n17257), .ZN(n16460) );
  NAND2_X1 U18536 ( .A1(n18382), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n16682) );
  OAI211_X1 U18537 ( .C1(n17222), .C2(n16461), .A(n16460), .B(n16682), .ZN(
        n16465) );
  OAI21_X1 U18538 ( .B1(n12114), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n16463), .ZN(n16678) );
  NOR2_X1 U18539 ( .A1(n16678), .A2(n17224), .ZN(n16464) );
  AOI211_X1 U18540 ( .C1(n17216), .C2(n16466), .A(n16465), .B(n16464), .ZN(
        n16467) );
  OAI21_X1 U18541 ( .B1(n16689), .B2(n17228), .A(n16467), .ZN(P2_U2993) );
  NOR2_X1 U18542 ( .A1(n16468), .A2(n18596), .ZN(n16470) );
  OAI21_X1 U18543 ( .B1(n16470), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n16469), .ZN(n16711) );
  NAND2_X1 U18544 ( .A1(n16690), .A2(n17258), .ZN(n16475) );
  INV_X1 U18545 ( .A(n18448), .ZN(n16708) );
  OAI22_X1 U18546 ( .A1(n17222), .A2(n11148), .B1(n18437), .B2(n18583), .ZN(
        n16473) );
  NOR2_X1 U18547 ( .A1(n18444), .A2(n17261), .ZN(n16472) );
  AOI211_X1 U18548 ( .C1(n17257), .C2(n16708), .A(n16473), .B(n16472), .ZN(
        n16474) );
  OAI211_X1 U18549 ( .C1(n17224), .C2(n16711), .A(n16475), .B(n16474), .ZN(
        P2_U2994) );
  XNOR2_X1 U18550 ( .A(n16468), .B(n18596), .ZN(n18608) );
  NAND2_X1 U18551 ( .A1(n16477), .A2(n16476), .ZN(n16481) );
  INV_X1 U18552 ( .A(n16491), .ZN(n16478) );
  NOR2_X1 U18553 ( .A1(n16493), .A2(n16478), .ZN(n16496) );
  INV_X1 U18554 ( .A(n16495), .ZN(n16479) );
  NOR2_X1 U18555 ( .A1(n16496), .A2(n16479), .ZN(n16480) );
  XOR2_X1 U18556 ( .A(n16481), .B(n16480), .Z(n18605) );
  OAI22_X1 U18557 ( .A1(n16482), .A2(n17222), .B1(n17261), .B2(n18432), .ZN(
        n16485) );
  OAI22_X1 U18558 ( .A1(n18429), .A2(n17227), .B1(n16483), .B2(n18583), .ZN(
        n16484) );
  OAI21_X1 U18559 ( .B1(n17224), .B2(n18608), .A(n16486), .ZN(P2_U2995) );
  INV_X1 U18560 ( .A(n16759), .ZN(n16488) );
  NAND2_X1 U18561 ( .A1(n16488), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16725) );
  OAI21_X1 U18562 ( .B1(n16725), .B2(n16736), .A(n16489), .ZN(n16490) );
  NAND2_X1 U18563 ( .A1(n16490), .A2(n16468), .ZN(n16721) );
  NAND2_X1 U18564 ( .A1(n16491), .A2(n16495), .ZN(n16492) );
  AND2_X1 U18565 ( .A1(n16493), .A2(n16492), .ZN(n16494) );
  AOI21_X1 U18566 ( .B1(n16496), .B2(n16495), .A(n16494), .ZN(n16719) );
  INV_X1 U18567 ( .A(n18418), .ZN(n16714) );
  NOR2_X1 U18568 ( .A1(n18582), .A2(n18417), .ZN(n16713) );
  NOR2_X1 U18569 ( .A1(n17222), .A2(n16497), .ZN(n16498) );
  AOI211_X1 U18570 ( .C1(n16714), .C2(n17257), .A(n16713), .B(n16498), .ZN(
        n16499) );
  OAI21_X1 U18571 ( .B1(n17261), .B2(n18424), .A(n16499), .ZN(n16500) );
  AOI21_X1 U18572 ( .B1(n16719), .B2(n17258), .A(n16500), .ZN(n16501) );
  OAI21_X1 U18573 ( .B1(n16721), .B2(n17224), .A(n16501), .ZN(P2_U2996) );
  XNOR2_X1 U18574 ( .A(n16725), .B(n16736), .ZN(n16513) );
  NAND2_X1 U18575 ( .A1(n10972), .A2(n16502), .ZN(n16506) );
  NAND2_X1 U18576 ( .A1(n16504), .A2(n16503), .ZN(n16505) );
  XNOR2_X1 U18577 ( .A(n16506), .B(n16505), .ZN(n16732) );
  INV_X1 U18578 ( .A(n18412), .ZN(n16509) );
  NOR2_X1 U18579 ( .A1(n18582), .A2(n18405), .ZN(n16728) );
  INV_X1 U18580 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16507) );
  NOR2_X1 U18581 ( .A1(n17222), .A2(n16507), .ZN(n16508) );
  AOI211_X1 U18582 ( .C1(n17216), .C2(n16509), .A(n16728), .B(n16508), .ZN(
        n16510) );
  OAI21_X1 U18583 ( .B1(n17227), .B2(n18406), .A(n16510), .ZN(n16511) );
  AOI21_X1 U18584 ( .B1(n16732), .B2(n17258), .A(n16511), .ZN(n16512) );
  OAI21_X1 U18585 ( .B1(n16513), .B2(n17224), .A(n16512), .ZN(P2_U2997) );
  OAI21_X1 U18586 ( .B1(n10973), .B2(n16515), .A(n10972), .ZN(n16748) );
  XNOR2_X1 U18587 ( .A(n16759), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16517) );
  NAND2_X1 U18588 ( .A1(n16517), .A2(n17256), .ZN(n16521) );
  INV_X1 U18589 ( .A(n18402), .ZN(n16745) );
  OAI22_X1 U18590 ( .A1(n17222), .A2(n18394), .B1(n16743), .B2(n18582), .ZN(
        n16519) );
  NOR2_X1 U18591 ( .A1(n18399), .A2(n17261), .ZN(n16518) );
  AOI211_X1 U18592 ( .C1(n17257), .C2(n16745), .A(n16519), .B(n16518), .ZN(
        n16520) );
  OAI211_X1 U18593 ( .C1(n17228), .C2(n16748), .A(n16521), .B(n16520), .ZN(
        P2_U2998) );
  INV_X1 U18594 ( .A(n16528), .ZN(n16529) );
  NAND2_X1 U18595 ( .A1(n16525), .A2(n16524), .ZN(n16553) );
  NOR2_X1 U18596 ( .A1(n16526), .A2(n16552), .ZN(n16545) );
  NAND2_X1 U18597 ( .A1(n16528), .A2(n16527), .ZN(n16544) );
  NOR2_X1 U18598 ( .A1(n16545), .A2(n16544), .ZN(n16543) );
  NOR2_X1 U18599 ( .A1(n16529), .A2(n16543), .ZN(n16533) );
  NAND2_X1 U18600 ( .A1(n16531), .A2(n16530), .ZN(n16532) );
  XOR2_X1 U18601 ( .A(n16533), .B(n16532), .Z(n16762) );
  OAI22_X1 U18602 ( .A1(n11151), .A2(n17222), .B1(n17261), .B2(n18385), .ZN(
        n16537) );
  INV_X1 U18603 ( .A(n18389), .ZN(n16535) );
  OAI22_X1 U18604 ( .A1(n16535), .A2(n17227), .B1(n16534), .B2(n18583), .ZN(
        n16536) );
  NOR2_X1 U18605 ( .A1(n16537), .A2(n16536), .ZN(n16540) );
  INV_X1 U18606 ( .A(n16487), .ZN(n16538) );
  INV_X1 U18607 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n16756) );
  NAND2_X1 U18608 ( .A1(n16538), .A2(n16756), .ZN(n16758) );
  NAND3_X1 U18609 ( .A1(n16759), .A2(n17256), .A3(n16758), .ZN(n16539) );
  OAI211_X1 U18610 ( .C1(n16762), .C2(n17228), .A(n16540), .B(n16539), .ZN(
        P2_U2999) );
  NOR2_X1 U18611 ( .A1(n16541), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n16542) );
  OR2_X1 U18612 ( .A1(n16487), .A2(n16542), .ZN(n18579) );
  INV_X1 U18613 ( .A(n18576), .ZN(n16550) );
  OAI22_X1 U18614 ( .A1(n12177), .A2(n18582), .B1(n17261), .B2(n18375), .ZN(
        n16549) );
  INV_X1 U18615 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n16546) );
  OAI22_X1 U18616 ( .A1(n17227), .A2(n16547), .B1(n16546), .B2(n17222), .ZN(
        n16548) );
  AOI211_X1 U18617 ( .C1(n16550), .C2(n17258), .A(n16549), .B(n16548), .ZN(
        n16551) );
  OAI21_X1 U18618 ( .B1(n17224), .B2(n18579), .A(n16551), .ZN(P2_U3000) );
  AOI21_X1 U18619 ( .B1(n16554), .B2(n16553), .A(n16552), .ZN(n16773) );
  NAND2_X1 U18620 ( .A1(n16579), .A2(n16765), .ZN(n17254) );
  INV_X1 U18621 ( .A(n17254), .ZN(n16556) );
  AOI21_X1 U18622 ( .B1(n16556), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16557) );
  NOR2_X1 U18623 ( .A1(n16557), .A2(n16541), .ZN(n16763) );
  NAND2_X1 U18624 ( .A1(n16763), .A2(n17256), .ZN(n16564) );
  OAI22_X1 U18625 ( .A1(n16558), .A2(n17222), .B1(n12171), .B2(n18582), .ZN(
        n16561) );
  NOR2_X1 U18626 ( .A1(n17227), .A2(n16559), .ZN(n16560) );
  AOI211_X1 U18627 ( .C1(n17216), .C2(n16562), .A(n16561), .B(n16560), .ZN(
        n16563) );
  OAI211_X1 U18628 ( .C1(n16773), .C2(n17228), .A(n16564), .B(n16563), .ZN(
        P2_U3001) );
  NAND2_X1 U18629 ( .A1(n16579), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16805) );
  OAI21_X1 U18630 ( .B1(n16805), .B2(n16779), .A(n11949), .ZN(n16565) );
  NAND2_X1 U18631 ( .A1(n16565), .A2(n17254), .ZN(n16788) );
  NAND2_X1 U18632 ( .A1(n16567), .A2(n16566), .ZN(n17250) );
  NAND2_X1 U18633 ( .A1(n17248), .A2(n16568), .ZN(n17249) );
  XNOR2_X1 U18634 ( .A(n17250), .B(n17249), .ZN(n16786) );
  OAI22_X1 U18635 ( .A1(n16569), .A2(n17222), .B1(n12163), .B2(n18582), .ZN(
        n16573) );
  INV_X1 U18636 ( .A(n18352), .ZN(n16571) );
  INV_X1 U18637 ( .A(n18350), .ZN(n16570) );
  OAI22_X1 U18638 ( .A1(n17227), .A2(n16571), .B1(n17261), .B2(n16570), .ZN(
        n16572) );
  AOI211_X1 U18639 ( .C1(n16786), .C2(n17258), .A(n16573), .B(n16572), .ZN(
        n16574) );
  OAI21_X1 U18640 ( .B1(n16788), .B2(n17224), .A(n16574), .ZN(P2_U3003) );
  INV_X1 U18641 ( .A(n16795), .ZN(n16578) );
  OAI21_X1 U18642 ( .B1(n16576), .B2(n16578), .A(n16575), .ZN(n16577) );
  OAI21_X1 U18643 ( .B1(n16796), .B2(n16578), .A(n16577), .ZN(n16817) );
  INV_X1 U18644 ( .A(n16579), .ZN(n16580) );
  NAND2_X1 U18645 ( .A1(n16580), .A2(n16813), .ZN(n16806) );
  NAND3_X1 U18646 ( .A1(n16806), .A2(n17256), .A3(n16805), .ZN(n16585) );
  OAI22_X1 U18647 ( .A1(n16581), .A2(n17222), .B1(n12157), .B2(n18582), .ZN(
        n16583) );
  NOR2_X1 U18648 ( .A1(n18331), .A2(n17227), .ZN(n16582) );
  AOI211_X1 U18649 ( .C1(n17216), .C2(n18327), .A(n16583), .B(n16582), .ZN(
        n16584) );
  OAI211_X1 U18650 ( .C1(n17228), .C2(n16817), .A(n16585), .B(n16584), .ZN(
        P2_U3005) );
  INV_X1 U18651 ( .A(n16586), .ZN(n16588) );
  NOR2_X1 U18652 ( .A1(n16588), .A2(n16587), .ZN(n16589) );
  XNOR2_X1 U18653 ( .A(n16590), .B(n16589), .ZN(n16859) );
  OR2_X1 U18654 ( .A1(n16591), .A2(n16592), .ZN(n16846) );
  NAND2_X1 U18655 ( .A1(n16591), .A2(n16592), .ZN(n16845) );
  NAND3_X1 U18656 ( .A1(n16846), .A2(n16845), .A3(n17256), .ZN(n16597) );
  OAI22_X1 U18657 ( .A1(n16593), .A2(n17222), .B1(n12146), .B2(n18582), .ZN(
        n16595) );
  NOR2_X1 U18658 ( .A1(n18303), .A2(n17227), .ZN(n16594) );
  AOI211_X1 U18659 ( .C1(n17216), .C2(n18301), .A(n16595), .B(n16594), .ZN(
        n16596) );
  OAI211_X1 U18660 ( .C1(n16859), .C2(n17228), .A(n16597), .B(n16596), .ZN(
        P2_U3007) );
  INV_X1 U18661 ( .A(n18526), .ZN(n16603) );
  AOI21_X1 U18662 ( .B1(n18525), .B2(n18601), .A(n16598), .ZN(n16602) );
  MUX2_X1 U18663 ( .A(n16600), .B(n16599), .S(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .Z(n16601) );
  OAI211_X1 U18664 ( .C1(n16603), .C2(n16853), .A(n16602), .B(n16601), .ZN(
        n16604) );
  AOI21_X1 U18665 ( .B1(n16605), .B2(n18604), .A(n16604), .ZN(n16606) );
  OAI21_X1 U18666 ( .B1(n18609), .B2(n16607), .A(n16606), .ZN(P2_U3018) );
  NAND2_X1 U18667 ( .A1(n16608), .A2(n18604), .ZN(n16618) );
  INV_X1 U18668 ( .A(n16609), .ZN(n18516) );
  INV_X1 U18669 ( .A(n16610), .ZN(n16624) );
  NOR3_X1 U18670 ( .A1(n16611), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n16624), .ZN(n16616) );
  NAND3_X1 U18671 ( .A1(n16612), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n16727), .ZN(n16614) );
  OAI211_X1 U18672 ( .C1(n16871), .C2(n18522), .A(n16614), .B(n16613), .ZN(
        n16615) );
  AOI211_X1 U18673 ( .C1(n18516), .C2(n18603), .A(n16616), .B(n16615), .ZN(
        n16617) );
  OAI211_X1 U18674 ( .C1(n16619), .C2(n18609), .A(n16618), .B(n16617), .ZN(
        P2_U3019) );
  INV_X1 U18675 ( .A(n16620), .ZN(n18501) );
  NOR3_X1 U18676 ( .A1(n16642), .A2(n16774), .A3(n16621), .ZN(n16622) );
  AOI211_X1 U18677 ( .C1(n18601), .C2(n18501), .A(n16623), .B(n16622), .ZN(
        n16626) );
  OAI211_X1 U18678 ( .C1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(n16638), .B(n16624), .ZN(
        n16625) );
  OAI211_X1 U18679 ( .C1(n18500), .C2(n16853), .A(n16626), .B(n16625), .ZN(
        n16627) );
  AOI21_X1 U18680 ( .B1(n16628), .B2(n18604), .A(n16627), .ZN(n16629) );
  OAI21_X1 U18681 ( .B1(n16630), .B2(n18609), .A(n16629), .ZN(P2_U3020) );
  NAND2_X1 U18682 ( .A1(n16631), .A2(n16864), .ZN(n16640) );
  NOR3_X1 U18683 ( .A1(n16642), .A2(n16774), .A3(n16637), .ZN(n16636) );
  AOI21_X1 U18684 ( .B1(n18601), .B2(n18491), .A(n16632), .ZN(n16633) );
  OAI21_X1 U18685 ( .B1(n16634), .B2(n16853), .A(n16633), .ZN(n16635) );
  AOI211_X1 U18686 ( .C1(n16638), .C2(n16637), .A(n16636), .B(n16635), .ZN(
        n16639) );
  OAI211_X1 U18687 ( .C1(n16641), .C2(n18575), .A(n16640), .B(n16639), .ZN(
        P2_U3021) );
  NOR2_X1 U18688 ( .A1(n16667), .A2(n16655), .ZN(n16644) );
  INV_X1 U18689 ( .A(n16642), .ZN(n16643) );
  OAI21_X1 U18690 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n16644), .A(
        n16643), .ZN(n16647) );
  AOI21_X1 U18691 ( .B1(n18601), .B2(n11367), .A(n16645), .ZN(n16646) );
  OAI211_X1 U18692 ( .C1(n18480), .C2(n16853), .A(n16647), .B(n16646), .ZN(
        n16648) );
  AOI21_X1 U18693 ( .B1(n16649), .B2(n18604), .A(n16648), .ZN(n16650) );
  OAI21_X1 U18694 ( .B1(n16651), .B2(n18609), .A(n16650), .ZN(P2_U3022) );
  INV_X1 U18695 ( .A(n16652), .ZN(n18472) );
  NOR2_X1 U18696 ( .A1(n16871), .A2(n18478), .ZN(n16653) );
  AOI211_X1 U18697 ( .C1(n18472), .C2(n18603), .A(n16654), .B(n16653), .ZN(
        n16658) );
  INV_X1 U18698 ( .A(n16667), .ZN(n16656) );
  OAI211_X1 U18699 ( .C1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n16656), .B(n16655), .ZN(
        n16657) );
  OAI211_X1 U18700 ( .C1(n16665), .C2(n16659), .A(n16658), .B(n16657), .ZN(
        n16660) );
  AOI21_X1 U18701 ( .B1(n16661), .B2(n18604), .A(n16660), .ZN(n16662) );
  OAI21_X1 U18702 ( .B1(n16663), .B2(n18609), .A(n16662), .ZN(P2_U3023) );
  NAND2_X1 U18703 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n18382), .ZN(n16664) );
  OAI221_X1 U18704 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n16667), 
        .C1(n16666), .C2(n16665), .A(n16664), .ZN(n16674) );
  AOI21_X1 U18705 ( .B1(n16670), .B2(n16669), .A(n16668), .ZN(n19343) );
  INV_X1 U18706 ( .A(n19343), .ZN(n16671) );
  OAI22_X1 U18707 ( .A1(n16672), .A2(n16853), .B1(n16871), .B2(n16671), .ZN(
        n16673) );
  AOI211_X1 U18708 ( .C1(n16675), .C2(n18604), .A(n16674), .B(n16673), .ZN(
        n16676) );
  OAI21_X1 U18709 ( .B1(n16677), .B2(n18609), .A(n16676), .ZN(P2_U3024) );
  NOR2_X1 U18710 ( .A1(n16678), .A2(n18609), .ZN(n16687) );
  NOR3_X1 U18711 ( .A1(n18597), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n16704), .ZN(n16686) );
  AOI211_X1 U18712 ( .C1(n16810), .C2(n16680), .A(n16679), .B(n16774), .ZN(
        n16685) );
  NAND2_X1 U18713 ( .A1(n18601), .A2(n18449), .ZN(n16681) );
  OAI211_X1 U18714 ( .C1(n16683), .C2(n16853), .A(n16682), .B(n16681), .ZN(
        n16684) );
  NOR4_X1 U18715 ( .A1(n16687), .A2(n16686), .A3(n16685), .A4(n16684), .ZN(
        n16688) );
  OAI21_X1 U18716 ( .B1(n16689), .B2(n18575), .A(n16688), .ZN(P2_U3025) );
  NOR2_X1 U18717 ( .A1(n16692), .A2(n16691), .ZN(n16693) );
  OR2_X1 U18718 ( .A1(n15550), .A2(n16693), .ZN(n19440) );
  INV_X1 U18719 ( .A(n16757), .ZN(n16733) );
  NOR3_X1 U18720 ( .A1(n16733), .A2(n16697), .A3(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n16718) );
  INV_X1 U18721 ( .A(n16694), .ZN(n16722) );
  AOI21_X1 U18722 ( .B1(n16722), .B2(n16695), .A(n16826), .ZN(n16698) );
  OAI21_X1 U18723 ( .B1(n16698), .B2(n16697), .A(n16696), .ZN(n16701) );
  INV_X1 U18724 ( .A(n16699), .ZN(n16700) );
  OAI211_X1 U18725 ( .C1(n16722), .C2(n16867), .A(n16701), .B(n16700), .ZN(
        n16712) );
  NOR2_X1 U18726 ( .A1(n16718), .A2(n16712), .ZN(n18595) );
  INV_X1 U18727 ( .A(n18595), .ZN(n16702) );
  AOI22_X1 U18728 ( .A1(n18382), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n16702), .ZN(n16703) );
  OAI21_X1 U18729 ( .B1(n16871), .B2(n19440), .A(n16703), .ZN(n16707) );
  OAI21_X1 U18730 ( .B1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(n16704), .ZN(n16705) );
  NOR2_X1 U18731 ( .A1(n18597), .A2(n16705), .ZN(n16706) );
  AOI211_X1 U18732 ( .C1(n16708), .C2(n18603), .A(n16707), .B(n16706), .ZN(
        n16709) );
  OAI211_X1 U18733 ( .C1(n16711), .C2(n18609), .A(n16710), .B(n16709), .ZN(
        P2_U3026) );
  NAND2_X1 U18734 ( .A1(n16712), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n16716) );
  AOI21_X1 U18735 ( .B1(n16714), .B2(n18603), .A(n16713), .ZN(n16715) );
  OAI211_X1 U18736 ( .C1(n18419), .C2(n16871), .A(n16716), .B(n16715), .ZN(
        n16717) );
  AOI211_X1 U18737 ( .C1(n16719), .C2(n18604), .A(n16718), .B(n16717), .ZN(
        n16720) );
  OAI21_X1 U18738 ( .B1(n16721), .B2(n18609), .A(n16720), .ZN(P2_U3028) );
  OAI22_X1 U18739 ( .A1(n16764), .A2(n16722), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n16826), .ZN(n16723) );
  NOR2_X1 U18740 ( .A1(n16724), .A2(n16723), .ZN(n16754) );
  NAND2_X1 U18741 ( .A1(n16754), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n16739) );
  INV_X1 U18742 ( .A(n16725), .ZN(n16726) );
  AOI21_X1 U18743 ( .B1(n18609), .B2(n16867), .A(n16726), .ZN(n16740) );
  AOI21_X1 U18744 ( .B1(n16727), .B2(n16739), .A(n16740), .ZN(n16737) );
  AOI21_X1 U18745 ( .B1(n18601), .B2(n16729), .A(n16728), .ZN(n16730) );
  OAI21_X1 U18746 ( .B1(n18406), .B2(n16853), .A(n16730), .ZN(n16731) );
  AOI21_X1 U18747 ( .B1(n16732), .B2(n18604), .A(n16731), .ZN(n16735) );
  OAI22_X1 U18748 ( .A1(n16759), .A2(n18609), .B1(n16756), .B2(n16733), .ZN(
        n16738) );
  NAND3_X1 U18749 ( .A1(n16738), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n16736), .ZN(n16734) );
  OAI211_X1 U18750 ( .C1(n16737), .C2(n16736), .A(n16735), .B(n16734), .ZN(
        P2_U3029) );
  OAI22_X1 U18751 ( .A1(n16740), .A2(n16739), .B1(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n16738), .ZN(n16747) );
  AND2_X1 U18752 ( .A1(n16750), .A2(n16741), .ZN(n16742) );
  OR2_X1 U18753 ( .A1(n16347), .A2(n16742), .ZN(n19675) );
  OAI22_X1 U18754 ( .A1(n16871), .A2(n19675), .B1(n16743), .B2(n18583), .ZN(
        n16744) );
  AOI21_X1 U18755 ( .B1(n18603), .B2(n16745), .A(n16744), .ZN(n16746) );
  OAI211_X1 U18756 ( .C1(n16748), .C2(n18575), .A(n16747), .B(n16746), .ZN(
        P2_U3030) );
  NAND2_X1 U18757 ( .A1(n16749), .A2(n11043), .ZN(n16751) );
  NAND2_X1 U18758 ( .A1(n16751), .A2(n16750), .ZN(n19157) );
  OAI22_X1 U18759 ( .A1(n16871), .A2(n19157), .B1(n16534), .B2(n18582), .ZN(
        n16752) );
  AOI21_X1 U18760 ( .B1(n18603), .B2(n18389), .A(n16752), .ZN(n16753) );
  OAI21_X1 U18761 ( .B1(n16754), .B2(n16756), .A(n16753), .ZN(n16755) );
  AOI21_X1 U18762 ( .B1(n16757), .B2(n16756), .A(n16755), .ZN(n16761) );
  NAND3_X1 U18763 ( .A1(n16759), .A2(n16864), .A3(n16758), .ZN(n16760) );
  OAI211_X1 U18764 ( .C1(n16762), .C2(n18575), .A(n16761), .B(n16760), .ZN(
        P2_U3031) );
  NAND2_X1 U18765 ( .A1(n16763), .A2(n16864), .ZN(n16772) );
  OAI22_X1 U18766 ( .A1(n16871), .A2(n19164), .B1(n12171), .B2(n18583), .ZN(
        n16769) );
  NOR4_X1 U18767 ( .A1(n11949), .A2(n16779), .A3(n16813), .A4(n18570), .ZN(
        n18584) );
  OAI21_X1 U18768 ( .B1(n16765), .B2(n16764), .A(n16810), .ZN(n16766) );
  AOI21_X1 U18769 ( .B1(n18584), .B2(n17253), .A(n16766), .ZN(n18585) );
  NAND2_X1 U18770 ( .A1(n18584), .A2(n16767), .ZN(n18572) );
  OAI22_X1 U18771 ( .A1(n18585), .A2(n16767), .B1(n17253), .B2(n18572), .ZN(
        n16768) );
  AOI211_X1 U18772 ( .C1(n16770), .C2(n18603), .A(n16769), .B(n16768), .ZN(
        n16771) );
  OAI211_X1 U18773 ( .C1(n16773), .C2(n18575), .A(n16772), .B(n16771), .ZN(
        P2_U3033) );
  AOI21_X1 U18774 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16810), .A(
        n16774), .ZN(n16791) );
  NOR3_X1 U18775 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n16813), .A3(
        n18570), .ZN(n16790) );
  OAI21_X1 U18776 ( .B1(n16791), .B2(n16790), .A(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16784) );
  OR2_X1 U18777 ( .A1(n16776), .A2(n16775), .ZN(n16778) );
  NAND2_X1 U18778 ( .A1(n16778), .A2(n16777), .ZN(n19171) );
  NOR3_X1 U18779 ( .A1(n16779), .A2(n16813), .A3(n18570), .ZN(n16780) );
  AOI22_X1 U18780 ( .A1(n18382), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n11949), 
        .B2(n16780), .ZN(n16781) );
  OAI21_X1 U18781 ( .B1(n16871), .B2(n19171), .A(n16781), .ZN(n16782) );
  AOI21_X1 U18782 ( .B1(n18603), .B2(n18352), .A(n16782), .ZN(n16783) );
  NAND2_X1 U18783 ( .A1(n16784), .A2(n16783), .ZN(n16785) );
  AOI21_X1 U18784 ( .B1(n16786), .B2(n18604), .A(n16785), .ZN(n16787) );
  OAI21_X1 U18785 ( .B1(n16788), .B2(n18609), .A(n16787), .ZN(P2_U3035) );
  XNOR2_X1 U18786 ( .A(n16805), .B(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17241) );
  NAND2_X1 U18787 ( .A1(n17241), .A2(n16864), .ZN(n16804) );
  NOR2_X1 U18788 ( .A1(n12160), .A2(n18583), .ZN(n16789) );
  AOI211_X1 U18789 ( .C1(n16791), .C2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n16790), .B(n16789), .ZN(n16803) );
  XNOR2_X1 U18790 ( .A(n16793), .B(n16792), .ZN(n19174) );
  NOR2_X1 U18791 ( .A1(n16871), .A2(n19174), .ZN(n16794) );
  AOI21_X1 U18792 ( .B1(n18341), .B2(n18603), .A(n16794), .ZN(n16802) );
  NAND2_X1 U18793 ( .A1(n16796), .A2(n16795), .ZN(n16800) );
  NAND2_X1 U18794 ( .A1(n16798), .A2(n16797), .ZN(n16799) );
  XNOR2_X1 U18795 ( .A(n16800), .B(n16799), .ZN(n17242) );
  NAND2_X1 U18796 ( .A1(n17242), .A2(n18604), .ZN(n16801) );
  NAND4_X1 U18797 ( .A1(n16804), .A2(n16803), .A3(n16802), .A4(n16801), .ZN(
        P2_U3036) );
  NAND3_X1 U18798 ( .A1(n16806), .A2(n16864), .A3(n16805), .ZN(n16816) );
  INV_X1 U18799 ( .A(n18570), .ZN(n16814) );
  NAND2_X1 U18800 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n18382), .ZN(n16809) );
  XNOR2_X1 U18801 ( .A(n16807), .B(n11323), .ZN(n19177) );
  NAND2_X1 U18802 ( .A1(n18601), .A2(n19177), .ZN(n16808) );
  OAI211_X1 U18803 ( .C1(n16810), .C2(n16813), .A(n16809), .B(n16808), .ZN(
        n16812) );
  NOR2_X1 U18804 ( .A1(n18331), .A2(n16853), .ZN(n16811) );
  AOI211_X1 U18805 ( .C1(n16814), .C2(n16813), .A(n16812), .B(n16811), .ZN(
        n16815) );
  OAI211_X1 U18806 ( .C1(n16817), .C2(n18575), .A(n16816), .B(n16815), .ZN(
        P2_U3037) );
  NAND2_X1 U18807 ( .A1(n16845), .A2(n16818), .ZN(n16821) );
  OAI21_X1 U18808 ( .B1(n16821), .B2(n16820), .A(n16819), .ZN(n17235) );
  INV_X1 U18809 ( .A(n16822), .ZN(n16824) );
  NOR2_X1 U18810 ( .A1(n16824), .A2(n16823), .ZN(n16825) );
  INV_X1 U18811 ( .A(n16828), .ZN(n16832) );
  INV_X1 U18812 ( .A(n16826), .ZN(n16827) );
  OAI21_X1 U18813 ( .B1(n16829), .B2(n16828), .A(n16827), .ZN(n16831) );
  AND2_X1 U18814 ( .A1(n16831), .A2(n16830), .ZN(n16866) );
  OAI21_X1 U18815 ( .B1(n16832), .B2(n16867), .A(n16866), .ZN(n16856) );
  NAND2_X1 U18816 ( .A1(n16833), .A2(n16868), .ZN(n16876) );
  NOR2_X1 U18817 ( .A1(n16834), .A2(n16876), .ZN(n16851) );
  NAND2_X1 U18818 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16835) );
  AOI22_X1 U18819 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n16856), .B1(
        n16851), .B2(n16835), .ZN(n16836) );
  AOI21_X1 U18820 ( .B1(n16837), .B2(n16850), .A(n16836), .ZN(n16843) );
  AOI21_X1 U18821 ( .B1(n16840), .B2(n16838), .A(n16839), .ZN(n19180) );
  AOI22_X1 U18822 ( .A1(n18601), .A2(n19180), .B1(n18382), .B2(
        P2_REIP_REG_8__SCAN_IN), .ZN(n16841) );
  OAI21_X1 U18823 ( .B1(n18321), .B2(n16853), .A(n16841), .ZN(n16842) );
  AOI211_X1 U18824 ( .C1(n17237), .C2(n18604), .A(n16843), .B(n16842), .ZN(
        n16844) );
  OAI21_X1 U18825 ( .B1(n17235), .B2(n18609), .A(n16844), .ZN(P2_U3038) );
  NAND3_X1 U18826 ( .A1(n16846), .A2(n16845), .A3(n16864), .ZN(n16858) );
  OR2_X1 U18827 ( .A1(n16848), .A2(n16847), .ZN(n16849) );
  NAND2_X1 U18828 ( .A1(n16849), .A2(n16838), .ZN(n19185) );
  AOI22_X1 U18829 ( .A1(n18382), .A2(P2_REIP_REG_7__SCAN_IN), .B1(n16851), 
        .B2(n16850), .ZN(n16852) );
  OAI21_X1 U18830 ( .B1(n16871), .B2(n19185), .A(n16852), .ZN(n16855) );
  NOR2_X1 U18831 ( .A1(n18303), .A2(n16853), .ZN(n16854) );
  AOI211_X1 U18832 ( .C1(n16856), .C2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n16855), .B(n16854), .ZN(n16857) );
  OAI211_X1 U18833 ( .C1(n16859), .C2(n18575), .A(n16858), .B(n16857), .ZN(
        P2_U3039) );
  XNOR2_X1 U18834 ( .A(n16860), .B(n10960), .ZN(n17229) );
  NAND2_X1 U18835 ( .A1(n16862), .A2(n16861), .ZN(n16863) );
  NOR2_X1 U18836 ( .A1(n16863), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17225) );
  INV_X1 U18837 ( .A(n17225), .ZN(n16865) );
  NAND2_X1 U18838 ( .A1(n16863), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17231) );
  NAND3_X1 U18839 ( .A1(n16865), .A2(n16864), .A3(n17231), .ZN(n16879) );
  OAI21_X1 U18840 ( .B1(n16868), .B2(n16867), .A(n16866), .ZN(n16874) );
  NOR2_X1 U18841 ( .A1(n12138), .A2(n18583), .ZN(n16873) );
  XNOR2_X1 U18842 ( .A(n16870), .B(n16869), .ZN(n19350) );
  NOR2_X1 U18843 ( .A1(n16871), .A2(n19350), .ZN(n16872) );
  AOI211_X1 U18844 ( .C1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n16874), .A(
        n16873), .B(n16872), .ZN(n16875) );
  OAI21_X1 U18845 ( .B1(n16876), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n16875), .ZN(n16877) );
  AOI21_X1 U18846 ( .B1(n18297), .B2(n18603), .A(n16877), .ZN(n16878) );
  OAI211_X1 U18847 ( .C1(n17229), .C2(n18575), .A(n16879), .B(n16878), .ZN(
        P2_U3040) );
  NAND2_X1 U18848 ( .A1(n12241), .A2(n16881), .ZN(n16885) );
  NAND2_X1 U18849 ( .A1(n16883), .A2(n16882), .ZN(n16884) );
  NAND3_X1 U18850 ( .A1(n16885), .A2(n16886), .A3(n16884), .ZN(n16891) );
  NAND2_X1 U18851 ( .A1(n16887), .A2(n16886), .ZN(n16889) );
  NAND2_X1 U18852 ( .A1(n12241), .A2(n15322), .ZN(n16888) );
  NAND2_X1 U18853 ( .A1(n16889), .A2(n16888), .ZN(n16890) );
  MUX2_X1 U18854 ( .A(n16891), .B(n16890), .S(n11613), .Z(n16893) );
  NOR2_X1 U18855 ( .A1(n16893), .A2(n16892), .ZN(n16894) );
  NAND2_X1 U18856 ( .A1(n16895), .A2(n16894), .ZN(n18612) );
  INV_X1 U18857 ( .A(n18612), .ZN(n16896) );
  OAI22_X1 U18858 ( .A1(n19453), .A2(n18668), .B1(n16896), .B2(n18658), .ZN(
        n16898) );
  MUX2_X1 U18859 ( .A(n16898), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n16897), .Z(P2_U3596) );
  NOR2_X1 U18860 ( .A1(n17747), .A2(n16899), .ZN(n17348) );
  INV_X1 U18861 ( .A(n20562), .ZN(n16901) );
  NAND2_X1 U18862 ( .A1(n20091), .A2(n16900), .ZN(n16912) );
  INV_X1 U18863 ( .A(n21659), .ZN(n21619) );
  AOI211_X1 U18864 ( .C1(n16901), .C2(n16912), .A(n21619), .B(n21192), .ZN(
        n16903) );
  NOR3_X1 U18865 ( .A1(n17348), .A2(n16903), .A3(n16902), .ZN(n21208) );
  INV_X1 U18866 ( .A(n21208), .ZN(n21199) );
  NOR2_X1 U18867 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n21232), .ZN(n18718) );
  INV_X1 U18868 ( .A(n20796), .ZN(n20793) );
  INV_X1 U18869 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n21197) );
  NOR2_X1 U18870 ( .A1(n16905), .A2(n20750), .ZN(n21220) );
  NOR2_X1 U18871 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n20791) );
  NAND3_X1 U18872 ( .A1(n20793), .A2(n21220), .A3(n20791), .ZN(n16906) );
  OAI21_X1 U18873 ( .B1(n20793), .B2(n21197), .A(n16906), .ZN(P3_U3284) );
  INV_X1 U18874 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n16907) );
  OAI21_X1 U18875 ( .B1(P3_STATE_REG_2__SCAN_IN), .B2(n21658), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n18214) );
  NAND2_X1 U18876 ( .A1(n18235), .A2(n18214), .ZN(n16909) );
  INV_X1 U18877 ( .A(n16909), .ZN(n21615) );
  INV_X1 U18878 ( .A(n21615), .ZN(n16908) );
  INV_X1 U18879 ( .A(BS16), .ZN(n17157) );
  INV_X1 U18880 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n21666) );
  NAND2_X1 U18881 ( .A1(n21666), .A2(n21658), .ZN(n21617) );
  AOI21_X1 U18882 ( .B1(n17157), .B2(n21617), .A(n16908), .ZN(n21611) );
  AOI21_X1 U18883 ( .B1(n16907), .B2(n16908), .A(n21611), .ZN(P3_U3280) );
  AND2_X1 U18884 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n16908), .ZN(P3_U3028) );
  AND2_X1 U18885 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n16908), .ZN(P3_U3027) );
  AND2_X1 U18886 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n16908), .ZN(P3_U3026) );
  AND2_X1 U18887 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n16908), .ZN(P3_U3025) );
  AND2_X1 U18888 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n16908), .ZN(P3_U3024) );
  AND2_X1 U18889 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n16908), .ZN(P3_U3023) );
  AND2_X1 U18890 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n16908), .ZN(P3_U3022) );
  AND2_X1 U18891 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n16908), .ZN(P3_U3021) );
  AND2_X1 U18892 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n16908), .ZN(
        P3_U3020) );
  AND2_X1 U18893 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n16908), .ZN(
        P3_U3019) );
  AND2_X1 U18894 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n16908), .ZN(
        P3_U3018) );
  AND2_X1 U18895 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n16908), .ZN(
        P3_U3017) );
  AND2_X1 U18896 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n16908), .ZN(
        P3_U3016) );
  AND2_X1 U18897 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n16909), .ZN(
        P3_U3015) );
  AND2_X1 U18898 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n16909), .ZN(
        P3_U3014) );
  AND2_X1 U18899 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n16909), .ZN(
        P3_U3013) );
  AND2_X1 U18900 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n16909), .ZN(
        P3_U3012) );
  AND2_X1 U18901 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n16909), .ZN(
        P3_U3011) );
  AND2_X1 U18902 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n16909), .ZN(
        P3_U3010) );
  AND2_X1 U18903 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n16909), .ZN(
        P3_U3009) );
  AND2_X1 U18904 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n16909), .ZN(
        P3_U3008) );
  AND2_X1 U18905 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n16909), .ZN(
        P3_U3007) );
  AND2_X1 U18906 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n16909), .ZN(
        P3_U3006) );
  AND2_X1 U18907 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n16909), .ZN(
        P3_U3005) );
  AND2_X1 U18908 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n16909), .ZN(
        P3_U3004) );
  AND2_X1 U18909 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n16909), .ZN(
        P3_U3003) );
  AND2_X1 U18910 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n16909), .ZN(
        P3_U3002) );
  AND2_X1 U18911 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n16908), .ZN(
        P3_U3001) );
  AND2_X1 U18912 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n16908), .ZN(
        P3_U3000) );
  AND2_X1 U18913 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n16909), .ZN(
        P3_U2999) );
  AOI21_X1 U18914 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n16911)
         );
  NOR4_X1 U18915 ( .A1(n20754), .A2(n20095), .A3(n21659), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n21182) );
  AOI211_X1 U18916 ( .C1(n18096), .C2(n16911), .A(n16910), .B(n21182), .ZN(
        P3_U2998) );
  NAND2_X1 U18917 ( .A1(n20095), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18135) );
  NOR2_X1 U18918 ( .A1(n20754), .A2(n18135), .ZN(n21233) );
  AND2_X1 U18919 ( .A1(n18203), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  AOI21_X1 U18920 ( .B1(n21235), .B2(n21232), .A(n16913), .ZN(n16914) );
  INV_X1 U18921 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18168) );
  AOI22_X1 U18922 ( .A1(n16914), .A2(n18168), .B1(n16913), .B2(n20093), .ZN(
        P3_U3298) );
  INV_X1 U18923 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18167) );
  NOR2_X1 U18924 ( .A1(n11096), .A2(n20099), .ZN(n20550) );
  AOI21_X1 U18925 ( .B1(n16914), .B2(n18167), .A(n20550), .ZN(P3_U3299) );
  INV_X1 U18926 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n16915) );
  NOR2_X1 U18927 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n16915), .ZN(n21647) );
  AOI21_X1 U18928 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n21647), .A(n21641), 
        .ZN(n16917) );
  INV_X1 U18929 ( .A(n16917), .ZN(n21610) );
  INV_X1 U18930 ( .A(n21610), .ZN(n16918) );
  INV_X1 U18931 ( .A(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n16932) );
  NAND2_X1 U18932 ( .A1(n21640), .A2(n16915), .ZN(n16916) );
  AOI21_X1 U18933 ( .B1(n17157), .B2(n16916), .A(n16918), .ZN(n21606) );
  AOI21_X1 U18934 ( .B1(n16918), .B2(n16932), .A(n21606), .ZN(P2_U3591) );
  AND2_X1 U18935 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n16918), .ZN(P2_U3208) );
  AND2_X1 U18936 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n16918), .ZN(P2_U3207) );
  AND2_X1 U18937 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n16918), .ZN(P2_U3206) );
  AND2_X1 U18938 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n16918), .ZN(P2_U3205) );
  AND2_X1 U18939 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n16918), .ZN(P2_U3204) );
  AND2_X1 U18940 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n16918), .ZN(P2_U3203) );
  AND2_X1 U18941 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n16918), .ZN(P2_U3202) );
  AND2_X1 U18942 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n16918), .ZN(P2_U3201) );
  AND2_X1 U18943 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n16918), .ZN(
        P2_U3200) );
  AND2_X1 U18944 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n16918), .ZN(
        P2_U3199) );
  AND2_X1 U18945 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n16918), .ZN(
        P2_U3198) );
  AND2_X1 U18946 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n16918), .ZN(
        P2_U3197) );
  AND2_X1 U18947 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n16918), .ZN(
        P2_U3196) );
  AND2_X1 U18948 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n16918), .ZN(
        P2_U3195) );
  AND2_X1 U18949 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n16917), .ZN(
        P2_U3194) );
  AND2_X1 U18950 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n16917), .ZN(
        P2_U3193) );
  AND2_X1 U18951 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n16917), .ZN(
        P2_U3192) );
  AND2_X1 U18952 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n16917), .ZN(
        P2_U3191) );
  AND2_X1 U18953 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n16917), .ZN(
        P2_U3190) );
  AND2_X1 U18954 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n16917), .ZN(
        P2_U3189) );
  AND2_X1 U18955 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n16917), .ZN(
        P2_U3188) );
  AND2_X1 U18956 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n16917), .ZN(
        P2_U3187) );
  AND2_X1 U18957 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n16917), .ZN(
        P2_U3186) );
  AND2_X1 U18958 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n16917), .ZN(
        P2_U3185) );
  AND2_X1 U18959 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n16917), .ZN(
        P2_U3184) );
  AND2_X1 U18960 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n16917), .ZN(
        P2_U3183) );
  AND2_X1 U18961 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n16918), .ZN(
        P2_U3182) );
  AND2_X1 U18962 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n16918), .ZN(
        P2_U3181) );
  AND2_X1 U18963 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n16918), .ZN(
        P2_U3180) );
  AND2_X1 U18964 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n16918), .ZN(
        P2_U3179) );
  OAI221_X1 U18965 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(
        P2_STATEBS16_REG_SCAN_IN), .C1(n18669), .C2(n18675), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n16919) );
  AOI21_X1 U18966 ( .B1(n16919), .B2(n18247), .A(n18665), .ZN(P2_U3178) );
  INV_X1 U18967 ( .A(n18665), .ZN(n16920) );
  OAI221_X1 U18968 ( .B1(n16921), .B2(n16920), .C1(n18627), .C2(n16920), .A(
        n19683), .ZN(n17279) );
  NOR2_X1 U18969 ( .A1(n18619), .A2(n17279), .ZN(P2_U3047) );
  AND2_X1 U18970 ( .A1(n17307), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  NOR4_X1 U18971 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_12__SCAN_IN), .A3(P2_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16925) );
  NOR4_X1 U18972 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16924) );
  NOR4_X1 U18973 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16923) );
  NOR4_X1 U18974 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16922) );
  NAND4_X1 U18975 ( .A1(n16925), .A2(n16924), .A3(n16923), .A4(n16922), .ZN(
        n16931) );
  NOR4_X1 U18976 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_28__SCAN_IN), .A3(P2_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_26__SCAN_IN), .ZN(n16929) );
  AOI211_X1 U18977 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_31__SCAN_IN), .B(
        P2_DATAWIDTH_REG_30__SCAN_IN), .ZN(n16928) );
  NOR4_X1 U18978 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16927) );
  NOR4_X1 U18979 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_24__SCAN_IN), .A3(P2_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n16926) );
  NAND4_X1 U18980 ( .A1(n16929), .A2(n16928), .A3(n16927), .A4(n16926), .ZN(
        n16930) );
  NOR2_X1 U18981 ( .A1(n16931), .A2(n16930), .ZN(n17290) );
  INV_X1 U18982 ( .A(n17290), .ZN(n17288) );
  NOR2_X1 U18983 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n17288), .ZN(n17282) );
  INV_X1 U18984 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21609) );
  NAND3_X1 U18985 ( .A1(n17283), .A2(n21609), .A3(n16932), .ZN(n17287) );
  INV_X1 U18986 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16933) );
  AOI22_X1 U18987 ( .A1(n17282), .A2(n17287), .B1(n17288), .B2(n16933), .ZN(
        P2_U2821) );
  INV_X1 U18988 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n16934) );
  AOI22_X1 U18989 ( .A1(n17282), .A2(n17283), .B1(n17288), .B2(n16934), .ZN(
        P2_U2820) );
  INV_X1 U18990 ( .A(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(n16937) );
  INV_X1 U18991 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n16935) );
  NOR2_X1 U18992 ( .A1(n16935), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n21631) );
  NAND2_X1 U18993 ( .A1(n13632), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n22308) );
  OAI21_X1 U18994 ( .B1(n21631), .B2(n13632), .A(n22308), .ZN(n16938) );
  NOR2_X1 U18995 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n21625) );
  INV_X1 U18996 ( .A(n16938), .ZN(n21605) );
  OAI21_X1 U18997 ( .B1(BS16), .B2(n21625), .A(n21605), .ZN(n21603) );
  INV_X1 U18998 ( .A(n21603), .ZN(n16936) );
  AOI21_X1 U18999 ( .B1(n16937), .B2(n16938), .A(n16936), .ZN(P1_U3464) );
  AND2_X1 U19000 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n16938), .ZN(P1_U3193) );
  AND2_X1 U19001 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n16938), .ZN(P1_U3192) );
  AND2_X1 U19002 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n16938), .ZN(P1_U3191) );
  AND2_X1 U19003 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n16938), .ZN(P1_U3190) );
  AND2_X1 U19004 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n16938), .ZN(P1_U3189) );
  AND2_X1 U19005 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n16938), .ZN(P1_U3188) );
  AND2_X1 U19006 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n16938), .ZN(P1_U3187) );
  AND2_X1 U19007 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n16938), .ZN(P1_U3186) );
  AND2_X1 U19008 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n16938), .ZN(
        P1_U3185) );
  INV_X1 U19009 ( .A(n21605), .ZN(n16939) );
  AND2_X1 U19010 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n16939), .ZN(
        P1_U3184) );
  AND2_X1 U19011 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n16939), .ZN(
        P1_U3183) );
  AND2_X1 U19012 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n16939), .ZN(
        P1_U3182) );
  AND2_X1 U19013 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n16939), .ZN(
        P1_U3181) );
  AND2_X1 U19014 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n16939), .ZN(
        P1_U3180) );
  AND2_X1 U19015 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n16939), .ZN(
        P1_U3179) );
  AND2_X1 U19016 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n16939), .ZN(
        P1_U3178) );
  AND2_X1 U19017 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n16939), .ZN(
        P1_U3177) );
  AND2_X1 U19018 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n16939), .ZN(
        P1_U3176) );
  AND2_X1 U19019 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n16939), .ZN(
        P1_U3175) );
  AND2_X1 U19020 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n16939), .ZN(
        P1_U3174) );
  AND2_X1 U19021 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n16939), .ZN(
        P1_U3173) );
  AND2_X1 U19022 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n16939), .ZN(
        P1_U3172) );
  AND2_X1 U19023 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n16939), .ZN(
        P1_U3171) );
  AND2_X1 U19024 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n16939), .ZN(
        P1_U3170) );
  AND2_X1 U19025 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n16939), .ZN(
        P1_U3169) );
  AND2_X1 U19026 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n16939), .ZN(
        P1_U3168) );
  AND2_X1 U19027 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n16939), .ZN(
        P1_U3167) );
  AND2_X1 U19028 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n16939), .ZN(
        P1_U3166) );
  AND2_X1 U19029 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n16939), .ZN(
        P1_U3165) );
  AND2_X1 U19030 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n16939), .ZN(
        P1_U3164) );
  NOR2_X1 U19031 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21622), .ZN(n16945) );
  NOR3_X1 U19032 ( .A1(n16941), .A2(n21633), .A3(n16940), .ZN(n16942) );
  AOI221_X1 U19033 ( .B1(n16944), .B2(n16943), .C1(n21622), .C2(n16943), .A(
        n16942), .ZN(n16971) );
  AOI21_X1 U19034 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n16945), .A(n16971), 
        .ZN(n16975) );
  OAI221_X1 U19035 ( .B1(n16973), .B2(n16946), .C1(n16973), .C2(n21936), .A(
        n21583), .ZN(n16974) );
  INV_X1 U19036 ( .A(n16947), .ZN(n16949) );
  OAI21_X1 U19037 ( .B1(n16949), .B2(n16948), .A(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n16956) );
  NAND2_X1 U19038 ( .A1(n16950), .A2(n21794), .ZN(n16954) );
  INV_X1 U19039 ( .A(n16951), .ZN(n16952) );
  NAND4_X1 U19040 ( .A1(n16954), .A2(n16953), .A3(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A4(n16952), .ZN(n16955) );
  NAND2_X1 U19041 ( .A1(n16956), .A2(n16955), .ZN(n16959) );
  INV_X1 U19042 ( .A(n16957), .ZN(n16958) );
  AOI222_X1 U19043 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n16959), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16958), .C1(n16959), 
        .C2(n16958), .ZN(n16961) );
  AND2_X1 U19044 ( .A1(n16962), .A2(n21933), .ZN(n16960) );
  OAI221_X1 U19045 ( .B1(n16962), .B2(n21933), .C1(n16961), .C2(n16960), .A(
        n16977), .ZN(n16963) );
  INV_X1 U19046 ( .A(n16963), .ZN(n16970) );
  INV_X1 U19047 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n17057) );
  AOI21_X1 U19048 ( .B1(n14903), .B2(n17057), .A(n16964), .ZN(n16969) );
  NAND2_X1 U19049 ( .A1(n16966), .A2(n16965), .ZN(n16967) );
  NOR4_X1 U19050 ( .A1(n16970), .A2(n16969), .A3(n16968), .A4(n16967), .ZN(
        n21602) );
  OAI221_X1 U19051 ( .B1(P1_STATE2_REG_1__SCAN_IN), .B2(
        P1_STATE2_REG_0__SCAN_IN), .C1(P1_STATE2_REG_1__SCAN_IN), .C2(n21602), 
        .A(n16971), .ZN(n21591) );
  OAI211_X1 U19052 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n21622), .A(n16972), 
        .B(n21591), .ZN(n21599) );
  AOI22_X1 U19053 ( .A1(n16975), .A2(n16974), .B1(n16973), .B2(n21599), .ZN(
        P1_U3162) );
  NOR2_X1 U19054 ( .A1(n16977), .A2(n16976), .ZN(P1_U3032) );
  AND2_X1 U19055 ( .A1(n19865), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR2_X1 U19056 ( .A1(n21631), .A2(n13632), .ZN(n16978) );
  INV_X1 U19057 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n17164) );
  INV_X1 U19058 ( .A(n22308), .ZN(n22307) );
  AOI21_X1 U19059 ( .B1(n16978), .B2(n17164), .A(n22307), .ZN(P1_U2802) );
  OAI22_X1 U19060 ( .A1(n17081), .A2(keyinput_125), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(keyinput_126), .ZN(n16979) );
  AOI221_X1 U19061 ( .B1(n17081), .B2(keyinput_125), .C1(keyinput_126), .C2(
        P1_REIP_REG_21__SCAN_IN), .A(n16979), .ZN(n17208) );
  OAI22_X1 U19062 ( .A1(n17086), .A2(keyinput_124), .B1(n16981), .B2(
        keyinput_121), .ZN(n16980) );
  AOI221_X1 U19063 ( .B1(n17086), .B2(keyinput_124), .C1(keyinput_121), .C2(
        n16981), .A(n16980), .ZN(n17079) );
  OAI22_X1 U19064 ( .A1(n16983), .A2(keyinput_123), .B1(
        P1_REIP_REG_25__SCAN_IN), .B2(keyinput_122), .ZN(n16982) );
  AOI221_X1 U19065 ( .B1(n16983), .B2(keyinput_123), .C1(keyinput_122), .C2(
        P1_REIP_REG_25__SCAN_IN), .A(n16982), .ZN(n17078) );
  INV_X1 U19066 ( .A(keyinput_120), .ZN(n17076) );
  INV_X1 U19067 ( .A(keyinput_119), .ZN(n17074) );
  INV_X1 U19068 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17184) );
  INV_X1 U19069 ( .A(keyinput_115), .ZN(n17068) );
  INV_X1 U19070 ( .A(keyinput_114), .ZN(n17066) );
  INV_X1 U19071 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n19931) );
  INV_X1 U19072 ( .A(keyinput_113), .ZN(n17064) );
  INV_X1 U19073 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19935) );
  INV_X1 U19074 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n19938) );
  INV_X1 U19075 ( .A(keyinput_112), .ZN(n17062) );
  INV_X1 U19076 ( .A(keyinput_104), .ZN(n17050) );
  INV_X1 U19077 ( .A(keyinput_103), .ZN(n17048) );
  INV_X1 U19078 ( .A(P1_READREQUEST_REG_SCAN_IN), .ZN(n17162) );
  INV_X1 U19079 ( .A(READY1), .ZN(n17092) );
  OAI22_X1 U19080 ( .A1(n17092), .A2(keyinput_100), .B1(READY2), .B2(
        keyinput_101), .ZN(n16984) );
  AOI221_X1 U19081 ( .B1(n17092), .B2(keyinput_100), .C1(keyinput_101), .C2(
        READY2), .A(n16984), .ZN(n17045) );
  INV_X1 U19082 ( .A(keyinput_99), .ZN(n17043) );
  INV_X1 U19083 ( .A(HOLD), .ZN(n21665) );
  INV_X1 U19084 ( .A(keyinput_95), .ZN(n17037) );
  INV_X1 U19085 ( .A(DATAI_1_), .ZN(n17149) );
  INV_X1 U19086 ( .A(DATAI_3_), .ZN(n16986) );
  AOI22_X1 U19087 ( .A1(DATAI_4_), .A2(keyinput_92), .B1(n16986), .B2(
        keyinput_93), .ZN(n16985) );
  OAI221_X1 U19088 ( .B1(DATAI_4_), .B2(keyinput_92), .C1(n16986), .C2(
        keyinput_93), .A(n16985), .ZN(n17034) );
  INV_X1 U19089 ( .A(DATAI_5_), .ZN(n17142) );
  INV_X1 U19090 ( .A(keyinput_91), .ZN(n17032) );
  INV_X1 U19091 ( .A(keyinput_90), .ZN(n17030) );
  INV_X1 U19092 ( .A(DATAI_6_), .ZN(n17139) );
  INV_X1 U19093 ( .A(DATAI_7_), .ZN(n17096) );
  INV_X1 U19094 ( .A(DATAI_10_), .ZN(n17023) );
  INV_X1 U19095 ( .A(DATAI_11_), .ZN(n16989) );
  INV_X1 U19096 ( .A(DATAI_13_), .ZN(n16988) );
  AOI22_X1 U19097 ( .A1(n16989), .A2(keyinput_85), .B1(n16988), .B2(
        keyinput_83), .ZN(n16987) );
  OAI221_X1 U19098 ( .B1(n16989), .B2(keyinput_85), .C1(n16988), .C2(
        keyinput_83), .A(n16987), .ZN(n17021) );
  INV_X1 U19099 ( .A(DATAI_12_), .ZN(n17019) );
  INV_X1 U19100 ( .A(DATAI_15_), .ZN(n16991) );
  OAI22_X1 U19101 ( .A1(n16991), .A2(keyinput_81), .B1(keyinput_82), .B2(
        DATAI_14_), .ZN(n16990) );
  AOI221_X1 U19102 ( .B1(n16991), .B2(keyinput_81), .C1(DATAI_14_), .C2(
        keyinput_82), .A(n16990), .ZN(n17017) );
  AOI22_X1 U19103 ( .A1(n16994), .A2(keyinput_78), .B1(keyinput_79), .B2(
        n16993), .ZN(n16992) );
  OAI221_X1 U19104 ( .B1(n16994), .B2(keyinput_78), .C1(n16993), .C2(
        keyinput_79), .A(n16992), .ZN(n17015) );
  AOI22_X1 U19105 ( .A1(DATAI_22_), .A2(keyinput_74), .B1(DATAI_23_), .B2(
        keyinput_73), .ZN(n16995) );
  OAI221_X1 U19106 ( .B1(DATAI_22_), .B2(keyinput_74), .C1(DATAI_23_), .C2(
        keyinput_73), .A(n16995), .ZN(n17003) );
  AOI22_X1 U19107 ( .A1(DATAI_24_), .A2(keyinput_72), .B1(DATAI_25_), .B2(
        keyinput_71), .ZN(n16996) );
  OAI221_X1 U19108 ( .B1(DATAI_24_), .B2(keyinput_72), .C1(DATAI_25_), .C2(
        keyinput_71), .A(n16996), .ZN(n17002) );
  AOI22_X1 U19109 ( .A1(n17101), .A2(keyinput_68), .B1(keyinput_70), .B2(
        n17107), .ZN(n16997) );
  OAI221_X1 U19110 ( .B1(n17101), .B2(keyinput_68), .C1(n17107), .C2(
        keyinput_70), .A(n16997), .ZN(n17001) );
  AOI22_X1 U19111 ( .A1(n16999), .A2(keyinput_75), .B1(n17104), .B2(
        keyinput_69), .ZN(n16998) );
  OAI221_X1 U19112 ( .B1(n16999), .B2(keyinput_75), .C1(n17104), .C2(
        keyinput_69), .A(n16998), .ZN(n17000) );
  NOR4_X1 U19113 ( .A1(n17003), .A2(n17002), .A3(n17001), .A4(n17000), .ZN(
        n17012) );
  INV_X1 U19114 ( .A(keyinput_67), .ZN(n17008) );
  INV_X1 U19115 ( .A(keyinput_66), .ZN(n17006) );
  INV_X1 U19116 ( .A(DATAI_30_), .ZN(n22146) );
  AOI22_X1 U19117 ( .A1(P1_MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_64), .B1(
        DATAI_31_), .B2(keyinput_65), .ZN(n17004) );
  OAI221_X1 U19118 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_64), .C1(
        DATAI_31_), .C2(keyinput_65), .A(n17004), .ZN(n17005) );
  OAI221_X1 U19119 ( .B1(DATAI_30_), .B2(n17006), .C1(n22146), .C2(keyinput_66), .A(n17005), .ZN(n17007) );
  OAI221_X1 U19120 ( .B1(DATAI_29_), .B2(keyinput_67), .C1(n17118), .C2(n17008), .A(n17007), .ZN(n17011) );
  AOI22_X1 U19121 ( .A1(DATAI_19_), .A2(keyinput_77), .B1(n17120), .B2(
        keyinput_76), .ZN(n17009) );
  OAI221_X1 U19122 ( .B1(DATAI_19_), .B2(keyinput_77), .C1(n17120), .C2(
        keyinput_76), .A(n17009), .ZN(n17010) );
  AOI21_X1 U19123 ( .B1(n17012), .B2(n17011), .A(n17010), .ZN(n17014) );
  NAND2_X1 U19124 ( .A1(n17125), .A2(keyinput_80), .ZN(n17013) );
  OAI221_X1 U19125 ( .B1(n17015), .B2(n17014), .C1(n17125), .C2(keyinput_80), 
        .A(n17013), .ZN(n17016) );
  AOI22_X1 U19126 ( .A1(n17017), .A2(n17016), .B1(keyinput_84), .B2(n17019), 
        .ZN(n17018) );
  OAI21_X1 U19127 ( .B1(keyinput_84), .B2(n17019), .A(n17018), .ZN(n17020) );
  OAI22_X1 U19128 ( .A1(keyinput_86), .A2(n17023), .B1(n17021), .B2(n17020), 
        .ZN(n17022) );
  AOI21_X1 U19129 ( .B1(keyinput_86), .B2(n17023), .A(n17022), .ZN(n17028) );
  INV_X1 U19130 ( .A(DATAI_9_), .ZN(n17025) );
  OAI22_X1 U19131 ( .A1(n17025), .A2(keyinput_87), .B1(keyinput_88), .B2(
        DATAI_8_), .ZN(n17024) );
  AOI221_X1 U19132 ( .B1(n17025), .B2(keyinput_87), .C1(DATAI_8_), .C2(
        keyinput_88), .A(n17024), .ZN(n17026) );
  OAI21_X1 U19133 ( .B1(keyinput_89), .B2(n17096), .A(n17026), .ZN(n17027) );
  AOI211_X1 U19134 ( .C1(keyinput_89), .C2(n17096), .A(n17028), .B(n17027), 
        .ZN(n17029) );
  AOI221_X1 U19135 ( .B1(DATAI_6_), .B2(n17030), .C1(n17139), .C2(keyinput_90), 
        .A(n17029), .ZN(n17031) );
  AOI221_X1 U19136 ( .B1(DATAI_5_), .B2(keyinput_91), .C1(n17142), .C2(n17032), 
        .A(n17031), .ZN(n17033) );
  OAI22_X1 U19137 ( .A1(n17034), .A2(n17033), .B1(keyinput_94), .B2(DATAI_2_), 
        .ZN(n17035) );
  AOI21_X1 U19138 ( .B1(keyinput_94), .B2(DATAI_2_), .A(n17035), .ZN(n17036)
         );
  AOI221_X1 U19139 ( .B1(DATAI_1_), .B2(n17037), .C1(n17149), .C2(keyinput_95), 
        .A(n17036), .ZN(n17040) );
  INV_X1 U19140 ( .A(DATAI_0_), .ZN(n17152) );
  INV_X1 U19141 ( .A(NA), .ZN(n21667) );
  AOI22_X1 U19142 ( .A1(n17152), .A2(keyinput_96), .B1(keyinput_98), .B2(
        n21667), .ZN(n17038) );
  OAI221_X1 U19143 ( .B1(n17152), .B2(keyinput_96), .C1(n21667), .C2(
        keyinput_98), .A(n17038), .ZN(n17039) );
  AOI211_X1 U19144 ( .C1(n21665), .C2(keyinput_97), .A(n17040), .B(n17039), 
        .ZN(n17041) );
  OAI21_X1 U19145 ( .B1(n21665), .B2(keyinput_97), .A(n17041), .ZN(n17042) );
  OAI221_X1 U19146 ( .B1(BS16), .B2(keyinput_99), .C1(n17157), .C2(n17043), 
        .A(n17042), .ZN(n17044) );
  OAI211_X1 U19147 ( .C1(n17162), .C2(keyinput_102), .A(n17045), .B(n17044), 
        .ZN(n17046) );
  AOI21_X1 U19148 ( .B1(n17162), .B2(keyinput_102), .A(n17046), .ZN(n17047) );
  AOI221_X1 U19149 ( .B1(P1_ADS_N_REG_SCAN_IN), .B2(keyinput_103), .C1(n17164), 
        .C2(n17048), .A(n17047), .ZN(n17049) );
  AOI221_X1 U19150 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_104), .C1(
        n17168), .C2(n17050), .A(n17049), .ZN(n17052) );
  XOR2_X1 U19151 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(keyinput_105), .Z(n17051) );
  OAI22_X1 U19152 ( .A1(n17052), .A2(n17051), .B1(P1_D_C_N_REG_SCAN_IN), .B2(
        keyinput_106), .ZN(n17055) );
  OAI22_X1 U19153 ( .A1(n21936), .A2(keyinput_108), .B1(keyinput_107), .B2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n17053) );
  AOI221_X1 U19154 ( .B1(n21936), .B2(keyinput_108), .C1(
        P1_REQUESTPENDING_REG_SCAN_IN), .C2(keyinput_107), .A(n17053), .ZN(
        n17054) );
  OAI221_X1 U19155 ( .B1(n17055), .B2(keyinput_106), .C1(n17055), .C2(
        P1_D_C_N_REG_SCAN_IN), .A(n17054), .ZN(n17060) );
  OAI22_X1 U19156 ( .A1(n17057), .A2(keyinput_109), .B1(P1_FLUSH_REG_SCAN_IN), 
        .B2(keyinput_110), .ZN(n17056) );
  AOI221_X1 U19157 ( .B1(n17057), .B2(keyinput_109), .C1(keyinput_110), .C2(
        P1_FLUSH_REG_SCAN_IN), .A(n17056), .ZN(n17059) );
  NOR2_X1 U19158 ( .A1(P1_W_R_N_REG_SCAN_IN), .A2(keyinput_111), .ZN(n17058)
         );
  AOI221_X1 U19159 ( .B1(n17060), .B2(n17059), .C1(keyinput_111), .C2(
        P1_W_R_N_REG_SCAN_IN), .A(n17058), .ZN(n17061) );
  AOI221_X1 U19160 ( .B1(P1_BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_112), 
        .C1(n19938), .C2(n17062), .A(n17061), .ZN(n17063) );
  AOI221_X1 U19161 ( .B1(P1_BYTEENABLE_REG_1__SCAN_IN), .B2(n17064), .C1(
        n19935), .C2(keyinput_113), .A(n17063), .ZN(n17065) );
  AOI221_X1 U19162 ( .B1(P1_BYTEENABLE_REG_2__SCAN_IN), .B2(n17066), .C1(
        n19931), .C2(keyinput_114), .A(n17065), .ZN(n17067) );
  AOI221_X1 U19163 ( .B1(P1_BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput_115), 
        .C1(n17184), .C2(n17068), .A(n17067), .ZN(n17071) );
  AOI22_X1 U19164 ( .A1(P1_REIP_REG_31__SCAN_IN), .A2(keyinput_116), .B1(
        n17089), .B2(keyinput_117), .ZN(n17069) );
  OAI221_X1 U19165 ( .B1(P1_REIP_REG_31__SCAN_IN), .B2(keyinput_116), .C1(
        n17089), .C2(keyinput_117), .A(n17069), .ZN(n17070) );
  AOI211_X1 U19166 ( .C1(P1_REIP_REG_29__SCAN_IN), .C2(keyinput_118), .A(
        n17071), .B(n17070), .ZN(n17072) );
  OAI21_X1 U19167 ( .B1(P1_REIP_REG_29__SCAN_IN), .B2(keyinput_118), .A(n17072), .ZN(n17073) );
  OAI221_X1 U19168 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(keyinput_119), .C1(
        n17192), .C2(n17074), .A(n17073), .ZN(n17075) );
  OAI221_X1 U19169 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n17076), .C1(n17194), 
        .C2(keyinput_120), .A(n17075), .ZN(n17077) );
  NAND3_X1 U19170 ( .A1(n17079), .A2(n17078), .A3(n17077), .ZN(n17207) );
  OAI22_X1 U19171 ( .A1(n17081), .A2(keyinput_61), .B1(P1_REIP_REG_21__SCAN_IN), .B2(keyinput_62), .ZN(n17080) );
  AOI221_X1 U19172 ( .B1(n17081), .B2(keyinput_61), .C1(keyinput_62), .C2(
        P1_REIP_REG_21__SCAN_IN), .A(n17080), .ZN(n17201) );
  AOI22_X1 U19173 ( .A1(P1_REIP_REG_26__SCAN_IN), .A2(keyinput_57), .B1(
        P1_REIP_REG_24__SCAN_IN), .B2(keyinput_59), .ZN(n17082) );
  OAI221_X1 U19174 ( .B1(P1_REIP_REG_26__SCAN_IN), .B2(keyinput_57), .C1(
        P1_REIP_REG_24__SCAN_IN), .C2(keyinput_59), .A(n17082), .ZN(n17083) );
  INV_X1 U19175 ( .A(n17083), .ZN(n17199) );
  AOI22_X1 U19176 ( .A1(n17086), .A2(keyinput_60), .B1(keyinput_58), .B2(
        n17085), .ZN(n17084) );
  OAI221_X1 U19177 ( .B1(n17086), .B2(keyinput_60), .C1(n17085), .C2(
        keyinput_58), .A(n17084), .ZN(n17087) );
  INV_X1 U19178 ( .A(n17087), .ZN(n17198) );
  INV_X1 U19179 ( .A(keyinput_56), .ZN(n17195) );
  INV_X1 U19180 ( .A(keyinput_55), .ZN(n17191) );
  OAI22_X1 U19181 ( .A1(n17089), .A2(keyinput_53), .B1(P1_REIP_REG_29__SCAN_IN), .B2(keyinput_54), .ZN(n17088) );
  AOI221_X1 U19182 ( .B1(n17089), .B2(keyinput_53), .C1(keyinput_54), .C2(
        P1_REIP_REG_29__SCAN_IN), .A(n17088), .ZN(n17187) );
  INV_X1 U19183 ( .A(keyinput_51), .ZN(n17185) );
  INV_X1 U19184 ( .A(keyinput_50), .ZN(n17182) );
  INV_X1 U19185 ( .A(keyinput_49), .ZN(n17180) );
  INV_X1 U19186 ( .A(keyinput_48), .ZN(n17178) );
  OAI22_X1 U19187 ( .A1(n14903), .A2(keyinput_46), .B1(P1_MORE_REG_SCAN_IN), 
        .B2(keyinput_45), .ZN(n17090) );
  AOI221_X1 U19188 ( .B1(n14903), .B2(keyinput_46), .C1(keyinput_45), .C2(
        P1_MORE_REG_SCAN_IN), .A(n17090), .ZN(n17175) );
  INV_X1 U19189 ( .A(keyinput_40), .ZN(n17167) );
  INV_X1 U19190 ( .A(keyinput_39), .ZN(n17165) );
  OAI22_X1 U19191 ( .A1(n17092), .A2(keyinput_36), .B1(keyinput_37), .B2(
        READY2), .ZN(n17091) );
  AOI221_X1 U19192 ( .B1(n17092), .B2(keyinput_36), .C1(READY2), .C2(
        keyinput_37), .A(n17091), .ZN(n17160) );
  INV_X1 U19193 ( .A(keyinput_35), .ZN(n17158) );
  INV_X1 U19194 ( .A(keyinput_31), .ZN(n17150) );
  INV_X1 U19195 ( .A(DATAI_2_), .ZN(n17147) );
  INV_X1 U19196 ( .A(DATAI_4_), .ZN(n17094) );
  AOI22_X1 U19197 ( .A1(DATAI_3_), .A2(keyinput_29), .B1(n17094), .B2(
        keyinput_28), .ZN(n17093) );
  OAI221_X1 U19198 ( .B1(DATAI_3_), .B2(keyinput_29), .C1(n17094), .C2(
        keyinput_28), .A(n17093), .ZN(n17145) );
  INV_X1 U19199 ( .A(keyinput_27), .ZN(n17143) );
  INV_X1 U19200 ( .A(keyinput_26), .ZN(n17140) );
  INV_X1 U19201 ( .A(DATAI_8_), .ZN(n17097) );
  OAI22_X1 U19202 ( .A1(n17097), .A2(keyinput_24), .B1(n17096), .B2(
        keyinput_25), .ZN(n17095) );
  AOI221_X1 U19203 ( .B1(n17097), .B2(keyinput_24), .C1(keyinput_25), .C2(
        n17096), .A(n17095), .ZN(n17136) );
  OAI22_X1 U19204 ( .A1(DATAI_14_), .A2(keyinput_18), .B1(DATAI_15_), .B2(
        keyinput_17), .ZN(n17098) );
  AOI221_X1 U19205 ( .B1(DATAI_14_), .B2(keyinput_18), .C1(keyinput_17), .C2(
        DATAI_15_), .A(n17098), .ZN(n17129) );
  AOI22_X1 U19206 ( .A1(DATAI_17_), .A2(keyinput_15), .B1(DATAI_18_), .B2(
        keyinput_14), .ZN(n17099) );
  OAI221_X1 U19207 ( .B1(DATAI_17_), .B2(keyinput_15), .C1(DATAI_18_), .C2(
        keyinput_14), .A(n17099), .ZN(n17127) );
  AOI22_X1 U19208 ( .A1(DATAI_21_), .A2(keyinput_11), .B1(n17101), .B2(
        keyinput_4), .ZN(n17100) );
  OAI221_X1 U19209 ( .B1(DATAI_21_), .B2(keyinput_11), .C1(n17101), .C2(
        keyinput_4), .A(n17100), .ZN(n17112) );
  AOI22_X1 U19210 ( .A1(DATAI_22_), .A2(keyinput_10), .B1(DATAI_25_), .B2(
        keyinput_7), .ZN(n17102) );
  OAI221_X1 U19211 ( .B1(DATAI_22_), .B2(keyinput_10), .C1(DATAI_25_), .C2(
        keyinput_7), .A(n17102), .ZN(n17111) );
  AOI22_X1 U19212 ( .A1(n17105), .A2(keyinput_8), .B1(n17104), .B2(keyinput_5), 
        .ZN(n17103) );
  OAI221_X1 U19213 ( .B1(n17105), .B2(keyinput_8), .C1(n17104), .C2(keyinput_5), .A(n17103), .ZN(n17110) );
  AOI22_X1 U19214 ( .A1(n17108), .A2(keyinput_9), .B1(n17107), .B2(keyinput_6), 
        .ZN(n17106) );
  OAI221_X1 U19215 ( .B1(n17108), .B2(keyinput_9), .C1(n17107), .C2(keyinput_6), .A(n17106), .ZN(n17109) );
  NOR4_X1 U19216 ( .A1(n17112), .A2(n17111), .A3(n17110), .A4(n17109), .ZN(
        n17123) );
  INV_X1 U19217 ( .A(keyinput_3), .ZN(n17117) );
  INV_X1 U19218 ( .A(keyinput_2), .ZN(n17115) );
  AOI22_X1 U19219 ( .A1(P1_MEMORYFETCH_REG_SCAN_IN), .A2(keyinput_0), .B1(
        DATAI_31_), .B2(keyinput_1), .ZN(n17113) );
  OAI221_X1 U19220 ( .B1(P1_MEMORYFETCH_REG_SCAN_IN), .B2(keyinput_0), .C1(
        DATAI_31_), .C2(keyinput_1), .A(n17113), .ZN(n17114) );
  OAI221_X1 U19221 ( .B1(DATAI_30_), .B2(n17115), .C1(n22146), .C2(keyinput_2), 
        .A(n17114), .ZN(n17116) );
  OAI221_X1 U19222 ( .B1(DATAI_29_), .B2(keyinput_3), .C1(n17118), .C2(n17117), 
        .A(n17116), .ZN(n17122) );
  AOI22_X1 U19223 ( .A1(DATAI_19_), .A2(keyinput_13), .B1(n17120), .B2(
        keyinput_12), .ZN(n17119) );
  OAI221_X1 U19224 ( .B1(DATAI_19_), .B2(keyinput_13), .C1(n17120), .C2(
        keyinput_12), .A(n17119), .ZN(n17121) );
  AOI21_X1 U19225 ( .B1(n17123), .B2(n17122), .A(n17121), .ZN(n17126) );
  NAND2_X1 U19226 ( .A1(n17125), .A2(keyinput_16), .ZN(n17124) );
  OAI221_X1 U19227 ( .B1(n17127), .B2(n17126), .C1(n17125), .C2(keyinput_16), 
        .A(n17124), .ZN(n17128) );
  AOI22_X1 U19228 ( .A1(n17129), .A2(n17128), .B1(DATAI_13_), .B2(keyinput_19), 
        .ZN(n17130) );
  OAI21_X1 U19229 ( .B1(DATAI_13_), .B2(keyinput_19), .A(n17130), .ZN(n17134)
         );
  AOI22_X1 U19230 ( .A1(DATAI_11_), .A2(keyinput_21), .B1(DATAI_12_), .B2(
        keyinput_20), .ZN(n17131) );
  OAI221_X1 U19231 ( .B1(DATAI_11_), .B2(keyinput_21), .C1(DATAI_12_), .C2(
        keyinput_20), .A(n17131), .ZN(n17133) );
  NAND2_X1 U19232 ( .A1(DATAI_10_), .A2(keyinput_22), .ZN(n17132) );
  OAI221_X1 U19233 ( .B1(n17134), .B2(n17133), .C1(DATAI_10_), .C2(keyinput_22), .A(n17132), .ZN(n17135) );
  OAI211_X1 U19234 ( .C1(DATAI_9_), .C2(keyinput_23), .A(n17136), .B(n17135), 
        .ZN(n17137) );
  AOI21_X1 U19235 ( .B1(DATAI_9_), .B2(keyinput_23), .A(n17137), .ZN(n17138)
         );
  AOI221_X1 U19236 ( .B1(DATAI_6_), .B2(n17140), .C1(n17139), .C2(keyinput_26), 
        .A(n17138), .ZN(n17141) );
  AOI221_X1 U19237 ( .B1(DATAI_5_), .B2(n17143), .C1(n17142), .C2(keyinput_27), 
        .A(n17141), .ZN(n17144) );
  OAI22_X1 U19238 ( .A1(keyinput_30), .A2(n17147), .B1(n17145), .B2(n17144), 
        .ZN(n17146) );
  AOI21_X1 U19239 ( .B1(keyinput_30), .B2(n17147), .A(n17146), .ZN(n17148) );
  AOI221_X1 U19240 ( .B1(DATAI_1_), .B2(n17150), .C1(n17149), .C2(keyinput_31), 
        .A(n17148), .ZN(n17154) );
  AOI22_X1 U19241 ( .A1(HOLD), .A2(keyinput_33), .B1(n17152), .B2(keyinput_32), 
        .ZN(n17151) );
  OAI221_X1 U19242 ( .B1(HOLD), .B2(keyinput_33), .C1(n17152), .C2(keyinput_32), .A(n17151), .ZN(n17153) );
  AOI211_X1 U19243 ( .C1(n21667), .C2(keyinput_34), .A(n17154), .B(n17153), 
        .ZN(n17155) );
  OAI21_X1 U19244 ( .B1(n21667), .B2(keyinput_34), .A(n17155), .ZN(n17156) );
  OAI221_X1 U19245 ( .B1(BS16), .B2(n17158), .C1(n17157), .C2(keyinput_35), 
        .A(n17156), .ZN(n17159) );
  OAI211_X1 U19246 ( .C1(n17162), .C2(keyinput_38), .A(n17160), .B(n17159), 
        .ZN(n17161) );
  AOI21_X1 U19247 ( .B1(n17162), .B2(keyinput_38), .A(n17161), .ZN(n17163) );
  AOI221_X1 U19248 ( .B1(P1_ADS_N_REG_SCAN_IN), .B2(n17165), .C1(n17164), .C2(
        keyinput_39), .A(n17163), .ZN(n17166) );
  AOI221_X1 U19249 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput_40), .C1(
        n17168), .C2(n17167), .A(n17166), .ZN(n17170) );
  XOR2_X1 U19250 ( .A(P1_M_IO_N_REG_SCAN_IN), .B(keyinput_41), .Z(n17169) );
  OAI22_X1 U19251 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(keyinput_42), .B1(n17170), 
        .B2(n17169), .ZN(n17173) );
  OAI22_X1 U19252 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(keyinput_44), .B1(
        P1_REQUESTPENDING_REG_SCAN_IN), .B2(keyinput_43), .ZN(n17171) );
  AOI221_X1 U19253 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(keyinput_44), .C1(
        keyinput_43), .C2(P1_REQUESTPENDING_REG_SCAN_IN), .A(n17171), .ZN(
        n17172) );
  OAI221_X1 U19254 ( .B1(n17173), .B2(keyinput_42), .C1(n17173), .C2(
        P1_D_C_N_REG_SCAN_IN), .A(n17172), .ZN(n17174) );
  AOI22_X1 U19255 ( .A1(n17175), .A2(n17174), .B1(keyinput_47), .B2(
        P1_W_R_N_REG_SCAN_IN), .ZN(n17176) );
  OAI21_X1 U19256 ( .B1(keyinput_47), .B2(P1_W_R_N_REG_SCAN_IN), .A(n17176), 
        .ZN(n17177) );
  OAI221_X1 U19257 ( .B1(P1_BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput_48), .C1(
        n19938), .C2(n17178), .A(n17177), .ZN(n17179) );
  OAI221_X1 U19258 ( .B1(P1_BYTEENABLE_REG_1__SCAN_IN), .B2(n17180), .C1(
        n19935), .C2(keyinput_49), .A(n17179), .ZN(n17181) );
  OAI221_X1 U19259 ( .B1(P1_BYTEENABLE_REG_2__SCAN_IN), .B2(keyinput_50), .C1(
        n19931), .C2(n17182), .A(n17181), .ZN(n17183) );
  OAI221_X1 U19260 ( .B1(P1_BYTEENABLE_REG_3__SCAN_IN), .B2(n17185), .C1(
        n17184), .C2(keyinput_51), .A(n17183), .ZN(n17186) );
  OAI211_X1 U19261 ( .C1(n17189), .C2(keyinput_52), .A(n17187), .B(n17186), 
        .ZN(n17188) );
  AOI21_X1 U19262 ( .B1(n17189), .B2(keyinput_52), .A(n17188), .ZN(n17190) );
  AOI221_X1 U19263 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(keyinput_55), .C1(
        n17192), .C2(n17191), .A(n17190), .ZN(n17193) );
  AOI221_X1 U19264 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n17195), .C1(n17194), 
        .C2(keyinput_56), .A(n17193), .ZN(n17196) );
  INV_X1 U19265 ( .A(n17196), .ZN(n17197) );
  NAND3_X1 U19266 ( .A1(n17199), .A2(n17198), .A3(n17197), .ZN(n17200) );
  NAND2_X1 U19267 ( .A1(n17201), .A2(n17200), .ZN(n17203) );
  AOI21_X1 U19268 ( .B1(keyinput_63), .B2(n17203), .A(keyinput_127), .ZN(
        n17205) );
  INV_X1 U19269 ( .A(keyinput_63), .ZN(n17202) );
  AOI21_X1 U19270 ( .B1(n17203), .B2(n17202), .A(n15972), .ZN(n17204) );
  AOI22_X1 U19271 ( .A1(n15972), .A2(n17205), .B1(keyinput_127), .B2(n17204), 
        .ZN(n17206) );
  AOI21_X1 U19272 ( .B1(n17208), .B2(n17207), .A(n17206), .ZN(n17213) );
  INV_X1 U19273 ( .A(n21761), .ZN(n17210) );
  NAND2_X1 U19274 ( .A1(n17210), .A2(n17209), .ZN(n21693) );
  AOI22_X1 U19275 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n21729), .B1(n21692), 
        .B2(P1_EAX_REG_19__SCAN_IN), .ZN(n17211) );
  NAND2_X1 U19276 ( .A1(n21693), .A2(n17211), .ZN(n17212) );
  XOR2_X1 U19277 ( .A(n17213), .B(n17212), .Z(P1_U2940) );
  INV_X1 U19278 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n17215) );
  OAI22_X1 U19279 ( .A1(n18248), .A2(n17215), .B1(n18669), .B2(n17214), .ZN(
        P2_U2816) );
  AOI22_X1 U19280 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n18382), .B1(n17216), 
        .B2(n18284), .ZN(n17221) );
  OAI22_X1 U19281 ( .A1(n17218), .A2(n17224), .B1(n17228), .B2(n17217), .ZN(
        n17219) );
  AOI21_X1 U19282 ( .B1(n17257), .B2(n18286), .A(n17219), .ZN(n17220) );
  OAI211_X1 U19283 ( .C1(n17223), .C2(n17222), .A(n17221), .B(n17220), .ZN(
        P2_U3009) );
  AOI22_X1 U19284 ( .A1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17245), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n18382), .ZN(n17234) );
  NOR2_X1 U19285 ( .A1(n17225), .A2(n17224), .ZN(n17232) );
  OAI22_X1 U19286 ( .A1(n17229), .A2(n17228), .B1(n17227), .B2(n17226), .ZN(
        n17230) );
  AOI21_X1 U19287 ( .B1(n17232), .B2(n17231), .A(n17230), .ZN(n17233) );
  OAI211_X1 U19288 ( .C1(n17261), .C2(n18294), .A(n17234), .B(n17233), .ZN(
        P2_U3008) );
  AOI22_X1 U19289 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n17245), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n18382), .ZN(n17240) );
  INV_X1 U19290 ( .A(n17235), .ZN(n17238) );
  AOI222_X1 U19291 ( .A1(n17238), .A2(n17256), .B1(n17258), .B2(n17237), .C1(
        n17257), .C2(n17236), .ZN(n17239) );
  OAI211_X1 U19292 ( .C1(n17261), .C2(n18316), .A(n17240), .B(n17239), .ZN(
        P2_U3006) );
  AOI22_X1 U19293 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17245), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n18382), .ZN(n17244) );
  AOI222_X1 U19294 ( .A1(n17242), .A2(n17258), .B1(n17257), .B2(n18341), .C1(
        n17256), .C2(n17241), .ZN(n17243) );
  OAI211_X1 U19295 ( .C1(n17261), .C2(n18334), .A(n17244), .B(n17243), .ZN(
        P2_U3004) );
  AOI22_X1 U19296 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17245), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n18382), .ZN(n17260) );
  NAND2_X1 U19297 ( .A1(n17247), .A2(n17246), .ZN(n17252) );
  OAI21_X1 U19298 ( .B1(n17250), .B2(n17249), .A(n17248), .ZN(n17251) );
  XOR2_X1 U19299 ( .A(n17252), .B(n17251), .Z(n18590) );
  INV_X1 U19300 ( .A(n18367), .ZN(n18589) );
  XNOR2_X1 U19301 ( .A(n17254), .B(n17253), .ZN(n18593) );
  INV_X1 U19302 ( .A(n18593), .ZN(n17255) );
  AOI222_X1 U19303 ( .A1(n18590), .A2(n17258), .B1(n17257), .B2(n18589), .C1(
        n17256), .C2(n17255), .ZN(n17259) );
  OAI211_X1 U19304 ( .C1(n17261), .C2(n18362), .A(n17260), .B(n17259), .ZN(
        P2_U3002) );
  INV_X1 U19305 ( .A(n17279), .ZN(n17281) );
  NOR2_X1 U19306 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19233), .ZN(
        n17264) );
  AND2_X1 U19307 ( .A1(n17263), .A2(n17262), .ZN(n18671) );
  AOI211_X1 U19308 ( .C1(n18260), .C2(n18250), .A(n17264), .B(n18671), .ZN(
        n17265) );
  AOI22_X1 U19309 ( .A1(n17281), .A2(n19263), .B1(n17265), .B2(n17279), .ZN(
        P2_U3605) );
  NAND2_X1 U19310 ( .A1(n19447), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19255) );
  OR2_X1 U19311 ( .A1(n19559), .A2(n19255), .ZN(n19293) );
  OR2_X1 U19312 ( .A1(n19255), .A2(n17266), .ZN(n17267) );
  AND2_X1 U19313 ( .A1(n17267), .A2(n18250), .ZN(n17276) );
  NAND2_X1 U19314 ( .A1(n19559), .A2(n17276), .ZN(n17269) );
  NAND2_X1 U19315 ( .A1(n19558), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n17268) );
  OAI211_X1 U19316 ( .C1(n19293), .C2(n19326), .A(n17269), .B(n17268), .ZN(
        n17270) );
  INV_X1 U19317 ( .A(n17270), .ZN(n17271) );
  AOI22_X1 U19318 ( .A1(n17281), .A2(n19221), .B1(n17271), .B2(n17279), .ZN(
        P2_U3603) );
  NOR2_X1 U19319 ( .A1(n19326), .A2(n21607), .ZN(n17277) );
  OR2_X1 U19320 ( .A1(n19447), .A2(n17277), .ZN(n17273) );
  NOR2_X1 U19321 ( .A1(n19449), .A2(n19233), .ZN(n17272) );
  AOI21_X1 U19322 ( .B1(n17276), .B2(n17273), .A(n17272), .ZN(n17274) );
  AOI22_X1 U19323 ( .A1(n17281), .A2(n19294), .B1(n17274), .B2(n17279), .ZN(
        P2_U3604) );
  OAI21_X1 U19324 ( .B1(n19256), .B2(n19448), .A(n19220), .ZN(n17278) );
  INV_X1 U19325 ( .A(n19509), .ZN(n17275) );
  AOI222_X1 U19326 ( .A1(n17278), .A2(n17277), .B1(n19330), .B2(n17276), .C1(
        P2_STATE2_REG_3__SCAN_IN), .C2(n17275), .ZN(n17280) );
  AOI22_X1 U19327 ( .A1(n17281), .A2(n19213), .B1(n17280), .B2(n17279), .ZN(
        P2_U3602) );
  NAND2_X1 U19328 ( .A1(n17282), .A2(n21609), .ZN(n17286) );
  OAI21_X1 U19329 ( .B1(n17326), .B2(n17283), .A(n17290), .ZN(n17284) );
  OAI21_X1 U19330 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n17290), .A(n17284), 
        .ZN(n17285) );
  OAI221_X1 U19331 ( .B1(n17286), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n17286), .C2(P2_REIP_REG_0__SCAN_IN), .A(n17285), .ZN(P2_U2822) );
  INV_X1 U19332 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n17289) );
  OAI221_X1 U19333 ( .B1(n17290), .B2(n17289), .C1(n17288), .C2(n17287), .A(
        n17286), .ZN(P2_U2823) );
  OAI22_X1 U19334 ( .A1(n17343), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n17340), .ZN(n17291) );
  INV_X1 U19335 ( .A(n17291), .ZN(P2_U3611) );
  INV_X1 U19336 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n17292) );
  AOI22_X1 U19337 ( .A1(n17340), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n17292), 
        .B2(n17343), .ZN(P2_U3608) );
  AOI21_X1 U19338 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n21610), .ZN(n17293) );
  INV_X1 U19339 ( .A(n17293), .ZN(P2_U2815) );
  INV_X1 U19340 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n17296) );
  AOI22_X1 U19341 ( .A1(n17321), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n17320), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n17295) );
  OAI21_X1 U19342 ( .B1(n17296), .B2(n17323), .A(n17295), .ZN(P2_U2951) );
  AOI22_X1 U19343 ( .A1(n17321), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n17320), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n17297) );
  OAI21_X1 U19344 ( .B1(n17298), .B2(n17323), .A(n17297), .ZN(P2_U2950) );
  INV_X1 U19345 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n17300) );
  AOI22_X1 U19346 ( .A1(n17321), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n17307), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n17299) );
  OAI21_X1 U19347 ( .B1(n17300), .B2(n17323), .A(n17299), .ZN(P2_U2949) );
  INV_X1 U19348 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n17302) );
  AOI22_X1 U19349 ( .A1(n17313), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n17307), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n17301) );
  OAI21_X1 U19350 ( .B1(n17302), .B2(n17323), .A(n17301), .ZN(P2_U2948) );
  INV_X1 U19351 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n17304) );
  AOI22_X1 U19352 ( .A1(n17321), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n17307), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n17303) );
  OAI21_X1 U19353 ( .B1(n17304), .B2(n17323), .A(n17303), .ZN(P2_U2947) );
  INV_X1 U19354 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n17306) );
  AOI22_X1 U19355 ( .A1(n17313), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n17307), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n17305) );
  OAI21_X1 U19356 ( .B1(n17306), .B2(n17323), .A(n17305), .ZN(P2_U2946) );
  INV_X1 U19357 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19348) );
  AOI22_X1 U19358 ( .A1(n17313), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n17307), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n17308) );
  OAI21_X1 U19359 ( .B1(n19348), .B2(n17323), .A(n17308), .ZN(P2_U2945) );
  INV_X1 U19360 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19184) );
  AOI22_X1 U19361 ( .A1(n17313), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n17320), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n17309) );
  OAI21_X1 U19362 ( .B1(n19184), .B2(n17323), .A(n17309), .ZN(P2_U2944) );
  INV_X1 U19363 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n17311) );
  AOI22_X1 U19364 ( .A1(n17313), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n17320), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n17310) );
  OAI21_X1 U19365 ( .B1(n17311), .B2(n17323), .A(n17310), .ZN(P2_U2943) );
  AOI22_X1 U19366 ( .A1(n17321), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n17320), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n17312) );
  OAI21_X1 U19367 ( .B1(n19179), .B2(n17323), .A(n17312), .ZN(P2_U2942) );
  AOI22_X1 U19368 ( .A1(n17313), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n17320), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n17314) );
  OAI21_X1 U19369 ( .B1(n17315), .B2(n17323), .A(n17314), .ZN(P2_U2941) );
  INV_X1 U19370 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19170) );
  AOI22_X1 U19371 ( .A1(n17321), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n17320), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n17316) );
  OAI21_X1 U19372 ( .B1(n19170), .B2(n17323), .A(n17316), .ZN(P2_U2940) );
  AOI22_X1 U19373 ( .A1(n17321), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n17320), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n17317) );
  OAI21_X1 U19374 ( .B1(n19168), .B2(n17323), .A(n17317), .ZN(P2_U2939) );
  INV_X1 U19375 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19163) );
  AOI22_X1 U19376 ( .A1(n17321), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n17320), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n17318) );
  OAI21_X1 U19377 ( .B1(n19163), .B2(n17323), .A(n17318), .ZN(P2_U2938) );
  AOI22_X1 U19378 ( .A1(n17321), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n17320), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n17319) );
  OAI21_X1 U19379 ( .B1(n19161), .B2(n17323), .A(n17319), .ZN(P2_U2937) );
  AOI22_X1 U19380 ( .A1(n17321), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n17320), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n17322) );
  OAI21_X1 U19381 ( .B1(n19156), .B2(n17323), .A(n17322), .ZN(P2_U2936) );
  AOI21_X1 U19382 ( .B1(n21655), .B2(n17324), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n17325) );
  AOI21_X1 U19383 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n17340), .A(n17325), 
        .ZN(P2_U2817) );
  OAI222_X1 U19384 ( .A1(n17339), .A2(n14561), .B1(n17327), .B2(n17340), .C1(
        n17326), .C2(n17337), .ZN(P2_U3212) );
  INV_X1 U19385 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n17328) );
  OAI222_X1 U19386 ( .A1(n17339), .A2(n15292), .B1(n17328), .B2(n17340), .C1(
        n14561), .C2(n17337), .ZN(P2_U3213) );
  INV_X1 U19387 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n17329) );
  OAI222_X1 U19388 ( .A1(n17339), .A2(n12132), .B1(n17329), .B2(n17340), .C1(
        n15292), .C2(n17337), .ZN(P2_U3214) );
  INV_X1 U19389 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n17330) );
  OAI222_X1 U19390 ( .A1(n17339), .A2(n12135), .B1(n17330), .B2(n17340), .C1(
        n12132), .C2(n17337), .ZN(P2_U3215) );
  INV_X1 U19391 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n17331) );
  OAI222_X1 U19392 ( .A1(n17339), .A2(n12138), .B1(n17331), .B2(n17340), .C1(
        n12135), .C2(n17337), .ZN(P2_U3216) );
  INV_X1 U19393 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19806) );
  OAI222_X1 U19394 ( .A1(n17339), .A2(n12146), .B1(n19806), .B2(n17340), .C1(
        n12138), .C2(n17337), .ZN(P2_U3217) );
  INV_X1 U19395 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19808) );
  OAI222_X1 U19396 ( .A1(n17339), .A2(n12349), .B1(n19808), .B2(n17340), .C1(
        n12146), .C2(n17337), .ZN(P2_U3218) );
  INV_X1 U19397 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19810) );
  OAI222_X1 U19398 ( .A1(n17339), .A2(n12157), .B1(n19810), .B2(n17340), .C1(
        n12349), .C2(n17337), .ZN(P2_U3219) );
  INV_X1 U19399 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19812) );
  OAI222_X1 U19400 ( .A1(n17337), .A2(n12157), .B1(n19812), .B2(n17340), .C1(
        n12160), .C2(n17339), .ZN(P2_U3220) );
  INV_X1 U19401 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19814) );
  OAI222_X1 U19402 ( .A1(n17337), .A2(n12160), .B1(n19814), .B2(n17340), .C1(
        n12163), .C2(n17339), .ZN(P2_U3221) );
  INV_X1 U19403 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19816) );
  OAI222_X1 U19404 ( .A1(n17337), .A2(n12163), .B1(n19816), .B2(n17340), .C1(
        n12419), .C2(n17339), .ZN(P2_U3222) );
  INV_X1 U19405 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19818) );
  OAI222_X1 U19406 ( .A1(n17337), .A2(n12419), .B1(n19818), .B2(n17340), .C1(
        n12171), .C2(n17339), .ZN(P2_U3223) );
  INV_X1 U19407 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19820) );
  OAI222_X1 U19408 ( .A1(n17337), .A2(n12171), .B1(n19820), .B2(n17340), .C1(
        n12177), .C2(n17339), .ZN(P2_U3224) );
  INV_X1 U19409 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19822) );
  OAI222_X1 U19410 ( .A1(n17337), .A2(n12177), .B1(n19822), .B2(n17340), .C1(
        n16534), .C2(n17339), .ZN(P2_U3225) );
  INV_X1 U19411 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19824) );
  OAI222_X1 U19412 ( .A1(n17337), .A2(n16534), .B1(n19824), .B2(n17340), .C1(
        n16743), .C2(n17339), .ZN(P2_U3226) );
  INV_X1 U19413 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19826) );
  OAI222_X1 U19414 ( .A1(n17337), .A2(n16743), .B1(n19826), .B2(n17340), .C1(
        n18405), .C2(n17339), .ZN(P2_U3227) );
  INV_X1 U19415 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19828) );
  OAI222_X1 U19416 ( .A1(n17337), .A2(n18405), .B1(n19828), .B2(n17340), .C1(
        n18417), .C2(n17339), .ZN(P2_U3228) );
  INV_X1 U19417 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19830) );
  OAI222_X1 U19418 ( .A1(n17339), .A2(n16483), .B1(n19830), .B2(n17340), .C1(
        n18417), .C2(n17337), .ZN(P2_U3229) );
  INV_X1 U19419 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n17332) );
  OAI222_X1 U19420 ( .A1(n17337), .A2(n16483), .B1(n17332), .B2(n17340), .C1(
        n18437), .C2(n17339), .ZN(P2_U3230) );
  INV_X1 U19421 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n17333) );
  OAI222_X1 U19422 ( .A1(n17339), .A2(n12207), .B1(n17333), .B2(n17340), .C1(
        n18437), .C2(n17337), .ZN(P2_U3231) );
  INV_X1 U19423 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19834) );
  OAI222_X1 U19424 ( .A1(n17339), .A2(n16433), .B1(n19834), .B2(n17340), .C1(
        n12207), .C2(n17337), .ZN(P2_U3232) );
  INV_X1 U19425 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19836) );
  OAI222_X1 U19426 ( .A1(n17339), .A2(n16423), .B1(n19836), .B2(n17340), .C1(
        n16433), .C2(n17337), .ZN(P2_U3233) );
  INV_X1 U19427 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19838) );
  OAI222_X1 U19428 ( .A1(n17339), .A2(n16413), .B1(n19838), .B2(n17340), .C1(
        n16423), .C2(n17337), .ZN(P2_U3234) );
  INV_X1 U19429 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19840) );
  OAI222_X1 U19430 ( .A1(n17339), .A2(n17334), .B1(n19840), .B2(n17340), .C1(
        n16413), .C2(n17337), .ZN(P2_U3235) );
  INV_X1 U19431 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19842) );
  OAI222_X1 U19432 ( .A1(n17337), .A2(n17334), .B1(n19842), .B2(n17340), .C1(
        n17335), .C2(n17339), .ZN(P2_U3236) );
  INV_X1 U19433 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19844) );
  OAI222_X1 U19434 ( .A1(n17339), .A2(n18511), .B1(n19844), .B2(n17340), .C1(
        n17335), .C2(n17337), .ZN(P2_U3237) );
  INV_X1 U19435 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19846) );
  OAI222_X1 U19436 ( .A1(n17337), .A2(n18511), .B1(n19846), .B2(n17340), .C1(
        n16372), .C2(n17339), .ZN(P2_U3238) );
  INV_X1 U19437 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19848) );
  OAI222_X1 U19438 ( .A1(n17337), .A2(n16372), .B1(n19848), .B2(n17340), .C1(
        n17336), .C2(n17339), .ZN(P2_U3239) );
  INV_X1 U19439 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19850) );
  OAI222_X1 U19440 ( .A1(n17337), .A2(n17336), .B1(n19850), .B2(n17340), .C1(
        n17338), .C2(n17339), .ZN(P2_U3240) );
  INV_X1 U19441 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19854) );
  OAI222_X1 U19442 ( .A1(n17339), .A2(n18550), .B1(n19854), .B2(n17340), .C1(
        n17338), .C2(n17337), .ZN(P2_U3241) );
  OAI22_X1 U19443 ( .A1(n17343), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n17340), .ZN(n17341) );
  INV_X1 U19444 ( .A(n17341), .ZN(P2_U3588) );
  OAI22_X1 U19445 ( .A1(n17343), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n17340), .ZN(n17342) );
  INV_X1 U19446 ( .A(n17342), .ZN(P2_U3587) );
  MUX2_X1 U19447 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n17343), .Z(P2_U3586) );
  OAI22_X1 U19448 ( .A1(n17343), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n17340), .ZN(n17344) );
  INV_X1 U19449 ( .A(n17344), .ZN(P2_U3585) );
  NOR3_X1 U19450 ( .A1(n20661), .A2(n17346), .A3(n17345), .ZN(n17347) );
  OAI21_X1 U19451 ( .B1(n17348), .B2(n17347), .A(n21221), .ZN(n20558) );
  NOR3_X1 U19452 ( .A1(n19007), .A2(n19057), .A3(n20558), .ZN(n17740) );
  INV_X1 U19453 ( .A(n17740), .ZN(n17734) );
  INV_X1 U19454 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n20556) );
  INV_X1 U19455 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n20148) );
  NOR2_X1 U19456 ( .A1(n20556), .A2(n20148), .ZN(n17353) );
  NAND4_X1 U19457 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .A4(n17353), .ZN(n17379) );
  NOR2_X1 U19458 ( .A1(n17734), .A2(n17379), .ZN(n17375) );
  NAND2_X1 U19459 ( .A1(n20722), .A2(n17375), .ZN(n17428) );
  INV_X1 U19460 ( .A(n17428), .ZN(n17372) );
  AND2_X1 U19461 ( .A1(n20661), .A2(n17740), .ZN(n17738) );
  INV_X2 U19462 ( .A(n17738), .ZN(n17736) );
  NOR2_X1 U19463 ( .A1(n20661), .A2(n17734), .ZN(n17737) );
  NAND3_X1 U19464 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17353), .A3(n17737), .ZN(
        n17350) );
  NOR2_X1 U19465 ( .A1(n20175), .A2(n17350), .ZN(n17352) );
  AOI21_X1 U19466 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17736), .A(n17352), .ZN(
        n17349) );
  INV_X1 U19467 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18917) );
  OAI22_X1 U19468 ( .A1(n17372), .A2(n17349), .B1(n18917), .B2(n17736), .ZN(
        P3_U2699) );
  INV_X1 U19469 ( .A(n17350), .ZN(n17355) );
  AOI21_X1 U19470 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17736), .A(n17355), .ZN(
        n17351) );
  OAI22_X1 U19471 ( .A1(n17352), .A2(n17351), .B1(n18958), .B2(n17736), .ZN(
        P3_U2700) );
  AOI22_X1 U19472 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17736), .B1(n17353), .B2(
        n17737), .ZN(n17354) );
  INV_X1 U19473 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19002) );
  OAI22_X1 U19474 ( .A1(n17355), .A2(n17354), .B1(n19002), .B2(n17736), .ZN(
        P3_U2701) );
  AOI22_X1 U19475 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17585), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17360) );
  AOI22_X1 U19476 ( .A1(n17719), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17590), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17359) );
  AOI22_X1 U19477 ( .A1(n17683), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n13463), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17358) );
  AOI22_X1 U19478 ( .A1(n13934), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17357) );
  NAND4_X1 U19479 ( .A1(n17360), .A2(n17359), .A3(n17358), .A4(n17357), .ZN(
        n17367) );
  AOI22_X1 U19480 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17535), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17365) );
  AOI22_X1 U19481 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17364) );
  AOI22_X1 U19482 ( .A1(n17703), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17363) );
  AOI22_X1 U19483 ( .A1(n17689), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17362) );
  NAND4_X1 U19484 ( .A1(n17365), .A2(n17364), .A3(n17363), .A4(n17362), .ZN(
        n17366) );
  NOR2_X1 U19485 ( .A1(n17367), .A2(n17366), .ZN(n20733) );
  NAND2_X1 U19486 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .ZN(n17377) );
  NOR3_X1 U19487 ( .A1(n17734), .A2(n17377), .A3(n17379), .ZN(n17369) );
  NAND3_X1 U19488 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .A3(n17369), .ZN(n17485) );
  OAI221_X1 U19489 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(P3_EBX_REG_7__SCAN_IN), 
        .C1(P3_EBX_REG_8__SCAN_IN), .C2(n17369), .A(n17485), .ZN(n17368) );
  AOI22_X1 U19490 ( .A1(n17738), .A2(n20733), .B1(n17368), .B2(n17736), .ZN(
        P3_U2695) );
  OR2_X1 U19491 ( .A1(n20231), .A2(n17369), .ZN(n17371) );
  OR3_X1 U19492 ( .A1(n17377), .A2(n17428), .A3(P3_EBX_REG_7__SCAN_IN), .ZN(
        n17370) );
  OAI221_X1 U19493 ( .B1(n17738), .B2(n17371), .C1(n17736), .C2(n18793), .A(
        n17370), .ZN(P3_U2696) );
  NAND2_X1 U19494 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17372), .ZN(n17374) );
  INV_X1 U19495 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18835) );
  NAND3_X1 U19496 ( .A1(n17374), .A2(P3_EBX_REG_6__SCAN_IN), .A3(n17736), .ZN(
        n17373) );
  OAI221_X1 U19497 ( .B1(n17374), .B2(P3_EBX_REG_6__SCAN_IN), .C1(n17736), 
        .C2(n18835), .A(n17373), .ZN(P3_U2697) );
  OAI211_X1 U19498 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n17375), .A(n17374), .B(
        n17736), .ZN(n17376) );
  OAI21_X1 U19499 ( .B1(n17736), .B2(n18876), .A(n17376), .ZN(P3_U2698) );
  INV_X1 U19500 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n20243) );
  NOR4_X1 U19501 ( .A1(n20252), .A2(n20243), .A3(n20231), .A4(n17377), .ZN(
        n17378) );
  NAND3_X1 U19502 ( .A1(P3_EBX_REG_11__SCAN_IN), .A2(P3_EBX_REG_10__SCAN_IN), 
        .A3(n17378), .ZN(n17429) );
  NOR2_X1 U19503 ( .A1(n17429), .A2(n17379), .ZN(n17406) );
  NAND4_X1 U19504 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(P3_EBX_REG_12__SCAN_IN), .A4(n17406), .ZN(n17401) );
  NOR2_X1 U19505 ( .A1(n20336), .A2(n17401), .ZN(n17489) );
  NAND2_X1 U19506 ( .A1(n17489), .A2(n17737), .ZN(n17402) );
  AOI22_X1 U19507 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17383) );
  AOI22_X1 U19508 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17382) );
  AOI22_X1 U19509 ( .A1(n13934), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n20181), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17381) );
  AOI22_X1 U19510 ( .A1(n17356), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17380) );
  NAND4_X1 U19511 ( .A1(n17383), .A2(n17382), .A3(n17381), .A4(n17380), .ZN(
        n17389) );
  AOI22_X1 U19512 ( .A1(n17688), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17387) );
  AOI22_X1 U19513 ( .A1(n17689), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17502), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17386) );
  AOI22_X1 U19514 ( .A1(n17585), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17535), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17385) );
  AOI22_X1 U19515 ( .A1(n13897), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17384) );
  NAND4_X1 U19516 ( .A1(n17387), .A2(n17386), .A3(n17385), .A4(n17384), .ZN(
        n17388) );
  NOR2_X1 U19517 ( .A1(n17389), .A2(n17388), .ZN(n20714) );
  NAND3_X1 U19518 ( .A1(n17402), .A2(P3_EBX_REG_16__SCAN_IN), .A3(n17736), 
        .ZN(n17390) );
  OAI221_X1 U19519 ( .B1(n17402), .B2(P3_EBX_REG_16__SCAN_IN), .C1(n17736), 
        .C2(n20714), .A(n17390), .ZN(P3_U2687) );
  AOI22_X1 U19520 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17590), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17400) );
  AOI22_X1 U19521 ( .A1(n17688), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17399) );
  AOI22_X1 U19522 ( .A1(n17585), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17535), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17391) );
  OAI21_X1 U19523 ( .B1(n11009), .B2(n18793), .A(n17391), .ZN(n17397) );
  AOI22_X1 U19524 ( .A1(n13897), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17502), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17395) );
  AOI22_X1 U19525 ( .A1(n17689), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17394) );
  AOI22_X1 U19526 ( .A1(n13934), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n13463), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17393) );
  AOI22_X1 U19527 ( .A1(n17683), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17392) );
  NAND4_X1 U19528 ( .A1(n17395), .A2(n17394), .A3(n17393), .A4(n17392), .ZN(
        n17396) );
  AOI211_X1 U19529 ( .C1(n17465), .C2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n17397), .B(n17396), .ZN(n17398) );
  NAND3_X1 U19530 ( .A1(n17400), .A2(n17399), .A3(n17398), .ZN(n20723) );
  INV_X1 U19531 ( .A(n20723), .ZN(n17405) );
  OAI21_X1 U19532 ( .B1(n17734), .B2(n17401), .A(n20336), .ZN(n17403) );
  NAND3_X1 U19533 ( .A1(n17403), .A2(n17402), .A3(n17736), .ZN(n17404) );
  OAI21_X1 U19534 ( .B1(n17405), .B2(n17736), .A(n17404), .ZN(P3_U2688) );
  NAND2_X1 U19535 ( .A1(n17737), .A2(n20308), .ZN(n17433) );
  NAND2_X1 U19536 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17406), .ZN(n17417) );
  AOI22_X1 U19537 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17410) );
  AOI22_X1 U19538 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17409) );
  AOI22_X1 U19539 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n13463), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17408) );
  AOI22_X1 U19540 ( .A1(n17683), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17407) );
  NAND4_X1 U19541 ( .A1(n17410), .A2(n17409), .A3(n17408), .A4(n17407), .ZN(
        n17416) );
  AOI22_X1 U19542 ( .A1(n13897), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17502), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17414) );
  AOI22_X1 U19543 ( .A1(n17689), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17535), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17413) );
  AOI22_X1 U19544 ( .A1(n17590), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17585), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17412) );
  AOI22_X1 U19545 ( .A1(n17719), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17411) );
  NAND4_X1 U19546 ( .A1(n17414), .A2(n17413), .A3(n17412), .A4(n17411), .ZN(
        n17415) );
  NOR2_X1 U19547 ( .A1(n17416), .A2(n17415), .ZN(n20568) );
  AOI21_X1 U19548 ( .B1(n20722), .B2(n17417), .A(n17734), .ZN(n17434) );
  OAI222_X1 U19549 ( .A1(n17433), .A2(n17417), .B1(n17736), .B2(n20568), .C1(
        n20308), .C2(n17434), .ZN(P3_U2690) );
  INV_X1 U19550 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17435) );
  AOI22_X1 U19551 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17535), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17427) );
  AOI22_X1 U19552 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17585), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17426) );
  INV_X1 U19553 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17654) );
  AOI22_X1 U19554 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17418) );
  OAI21_X1 U19555 ( .B1(n10964), .B2(n17654), .A(n17418), .ZN(n17424) );
  AOI22_X1 U19556 ( .A1(n17689), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17502), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17422) );
  AOI22_X1 U19557 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17421) );
  AOI22_X1 U19558 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17420) );
  AOI22_X1 U19559 ( .A1(n17683), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n13463), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17419) );
  NAND4_X1 U19560 ( .A1(n17422), .A2(n17421), .A3(n17420), .A4(n17419), .ZN(
        n17423) );
  AOI211_X1 U19561 ( .C1(n17688), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n17424), .B(n17423), .ZN(n17425) );
  NAND3_X1 U19562 ( .A1(n17427), .A2(n17426), .A3(n17425), .ZN(n20717) );
  INV_X1 U19563 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17430) );
  OR2_X1 U19564 ( .A1(n17429), .A2(n17428), .ZN(n17457) );
  NOR4_X1 U19565 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n20308), .A3(n17430), .A4(
        n17457), .ZN(n17431) );
  AOI21_X1 U19566 ( .B1(n17738), .B2(n20717), .A(n17431), .ZN(n17432) );
  OAI221_X1 U19567 ( .B1(n17435), .B2(n17434), .C1(n17435), .C2(n17433), .A(
        n17432), .ZN(P3_U2689) );
  AOI22_X1 U19568 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17535), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17439) );
  AOI22_X1 U19569 ( .A1(n17719), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17689), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17438) );
  AOI22_X1 U19570 ( .A1(n17356), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17437) );
  AOI22_X1 U19571 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n20181), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17436) );
  NAND4_X1 U19572 ( .A1(n17439), .A2(n17438), .A3(n17437), .A4(n17436), .ZN(
        n17445) );
  AOI22_X1 U19573 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17443) );
  AOI22_X1 U19574 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17442) );
  AOI22_X1 U19575 ( .A1(n17703), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17441) );
  AOI22_X1 U19576 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17440) );
  NAND4_X1 U19577 ( .A1(n17443), .A2(n17442), .A3(n17441), .A4(n17440), .ZN(
        n17444) );
  NOR2_X1 U19578 ( .A1(n17445), .A2(n17444), .ZN(n20572) );
  NAND3_X1 U19579 ( .A1(n17457), .A2(P3_EBX_REG_12__SCAN_IN), .A3(n17736), 
        .ZN(n17446) );
  OAI221_X1 U19580 ( .B1(n17457), .B2(P3_EBX_REG_12__SCAN_IN), .C1(n17736), 
        .C2(n20572), .A(n17446), .ZN(P3_U2691) );
  AOI22_X1 U19581 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17456) );
  AOI22_X1 U19582 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17455) );
  AOI22_X1 U19583 ( .A1(n17689), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17502), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17447) );
  OAI21_X1 U19584 ( .B1(n11009), .B2(n18958), .A(n17447), .ZN(n17453) );
  AOI22_X1 U19585 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17535), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17451) );
  AOI22_X1 U19586 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17585), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17450) );
  AOI22_X1 U19587 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n13463), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17449) );
  AOI22_X1 U19588 ( .A1(n17683), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17448) );
  NAND4_X1 U19589 ( .A1(n17451), .A2(n17450), .A3(n17449), .A4(n17448), .ZN(
        n17452) );
  AOI211_X1 U19590 ( .C1(n10966), .C2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n17453), .B(n17452), .ZN(n17454) );
  NAND3_X1 U19591 ( .A1(n17456), .A2(n17455), .A3(n17454), .ZN(n20577) );
  INV_X1 U19592 ( .A(n20577), .ZN(n17460) );
  NOR2_X1 U19593 ( .A1(n20252), .A2(n17485), .ZN(n17473) );
  AOI21_X1 U19594 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17473), .A(
        P3_EBX_REG_11__SCAN_IN), .ZN(n17459) );
  NAND2_X1 U19595 ( .A1(n17736), .A2(n17457), .ZN(n17458) );
  OAI22_X1 U19596 ( .A1(n17460), .A2(n17736), .B1(n17459), .B2(n17458), .ZN(
        P3_U2692) );
  AOI22_X1 U19597 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17535), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17464) );
  AOI22_X1 U19598 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17689), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17463) );
  AOI22_X1 U19599 ( .A1(n17683), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17462) );
  AOI22_X1 U19600 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n13463), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17461) );
  NAND4_X1 U19601 ( .A1(n17464), .A2(n17463), .A3(n17462), .A4(n17461), .ZN(
        n17471) );
  AOI22_X1 U19602 ( .A1(n17719), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17502), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17469) );
  AOI22_X1 U19603 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17468) );
  AOI22_X1 U19604 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17585), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17467) );
  AOI22_X1 U19605 ( .A1(n17698), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17466) );
  NAND4_X1 U19606 ( .A1(n17469), .A2(n17468), .A3(n17467), .A4(n17466), .ZN(
        n17470) );
  NOR2_X1 U19607 ( .A1(n17471), .A2(n17470), .ZN(n20580) );
  NOR2_X1 U19608 ( .A1(n17738), .A2(n17473), .ZN(n17486) );
  NOR2_X1 U19609 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n20661), .ZN(n17472) );
  AOI22_X1 U19610 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17486), .B1(n17473), 
        .B2(n17472), .ZN(n17474) );
  OAI21_X1 U19611 ( .B1(n20580), .B2(n17736), .A(n17474), .ZN(P3_U2693) );
  AOI22_X1 U19612 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17478) );
  AOI22_X1 U19613 ( .A1(n17689), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n17722), .ZN(n17477) );
  AOI22_X1 U19614 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17714), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n20181), .ZN(n17476) );
  AOI22_X1 U19615 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n17713), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17554), .ZN(n17475) );
  NAND4_X1 U19616 ( .A1(n17478), .A2(n17477), .A3(n17476), .A4(n17475), .ZN(
        n17484) );
  AOI22_X1 U19617 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17719), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17482) );
  AOI22_X1 U19618 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17688), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17481) );
  AOI22_X1 U19619 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17503), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17703), .ZN(n17480) );
  AOI22_X1 U19620 ( .A1(n17585), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17479) );
  NAND4_X1 U19621 ( .A1(n17482), .A2(n17481), .A3(n17480), .A4(n17479), .ZN(
        n17483) );
  NOR2_X1 U19622 ( .A1(n17484), .A2(n17483), .ZN(n20586) );
  INV_X1 U19623 ( .A(n17485), .ZN(n17487) );
  OAI21_X1 U19624 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17487), .A(n17486), .ZN(
        n17488) );
  OAI21_X1 U19625 ( .B1(n20586), .B2(n17736), .A(n17488), .ZN(P3_U2694) );
  INV_X1 U19626 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n20455) );
  NAND2_X1 U19627 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n17619) );
  INV_X1 U19628 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17681) );
  NAND2_X1 U19629 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17489), .ZN(n17731) );
  NOR2_X1 U19630 ( .A1(n20378), .A2(n17731), .ZN(n17730) );
  AND2_X1 U19631 ( .A1(n17740), .A2(n17730), .ZN(n17696) );
  NAND2_X1 U19632 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17711), .ZN(n17680) );
  NOR2_X1 U19633 ( .A1(n17681), .A2(n17680), .ZN(n17600) );
  NAND4_X1 U19634 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(P3_EBX_REG_21__SCAN_IN), .A4(n17600), .ZN(n17490) );
  NOR4_X1 U19635 ( .A1(n20524), .A2(n20455), .A3(n17619), .A4(n17490), .ZN(
        n17491) );
  NAND3_X1 U19636 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(n17491), .ZN(n17494) );
  NOR2_X1 U19637 ( .A1(n17495), .A2(n17494), .ZN(n17599) );
  NAND2_X1 U19638 ( .A1(n17736), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n17493) );
  NAND2_X1 U19639 ( .A1(n17599), .A2(n20722), .ZN(n17492) );
  OAI22_X1 U19640 ( .A1(n17599), .A2(n17493), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n17492), .ZN(P3_U2672) );
  NAND2_X1 U19641 ( .A1(n17495), .A2(n17494), .ZN(n17496) );
  NAND2_X1 U19642 ( .A1(n17496), .A2(n17736), .ZN(n17598) );
  AOI22_X1 U19643 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n17501) );
  AOI22_X1 U19644 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17500) );
  AOI22_X1 U19645 ( .A1(n17683), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n13463), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17499) );
  AOI22_X1 U19646 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17498) );
  NAND4_X1 U19647 ( .A1(n17501), .A2(n17500), .A3(n17499), .A4(n17498), .ZN(
        n17509) );
  AOI22_X1 U19648 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17502), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17507) );
  AOI22_X1 U19649 ( .A1(n17719), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17506) );
  AOI22_X1 U19650 ( .A1(n17698), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17535), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17505) );
  AOI22_X1 U19651 ( .A1(n17689), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17585), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17504) );
  NAND4_X1 U19652 ( .A1(n17507), .A2(n17506), .A3(n17505), .A4(n17504), .ZN(
        n17508) );
  NOR2_X1 U19653 ( .A1(n17509), .A2(n17508), .ZN(n17618) );
  AOI22_X1 U19654 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17535), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17514) );
  AOI22_X1 U19655 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17703), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17513) );
  AOI22_X1 U19656 ( .A1(n17713), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17512) );
  AOI22_X1 U19657 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n20181), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17511) );
  NAND4_X1 U19658 ( .A1(n17514), .A2(n17513), .A3(n17512), .A4(n17511), .ZN(
        n17520) );
  AOI22_X1 U19659 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17518) );
  AOI22_X1 U19660 ( .A1(n17719), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17689), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17517) );
  AOI22_X1 U19661 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17516) );
  AOI22_X1 U19662 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17585), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17515) );
  NAND4_X1 U19663 ( .A1(n17518), .A2(n17517), .A3(n17516), .A4(n17515), .ZN(
        n17519) );
  NOR2_X1 U19664 ( .A1(n17520), .A2(n17519), .ZN(n17614) );
  AOI22_X1 U19665 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17585), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17524) );
  AOI22_X1 U19666 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17703), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17523) );
  AOI22_X1 U19667 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n13463), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17522) );
  AOI22_X1 U19668 ( .A1(n20181), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17521) );
  NAND4_X1 U19669 ( .A1(n17524), .A2(n17523), .A3(n17522), .A4(n17521), .ZN(
        n17530) );
  AOI22_X1 U19670 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17528) );
  AOI22_X1 U19671 ( .A1(n17561), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17527) );
  AOI22_X1 U19672 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17689), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17526) );
  AOI22_X1 U19673 ( .A1(n17698), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17535), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17525) );
  NAND4_X1 U19674 ( .A1(n17528), .A2(n17527), .A3(n17526), .A4(n17525), .ZN(
        n17529) );
  NOR2_X1 U19675 ( .A1(n17530), .A2(n17529), .ZN(n17637) );
  AOI22_X1 U19676 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17534) );
  AOI22_X1 U19677 ( .A1(n17703), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17533) );
  AOI22_X1 U19678 ( .A1(n20181), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13463), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17532) );
  AOI22_X1 U19679 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17531) );
  NAND4_X1 U19680 ( .A1(n17534), .A2(n17533), .A3(n17532), .A4(n17531), .ZN(
        n17541) );
  AOI22_X1 U19681 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17535), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17539) );
  AOI22_X1 U19682 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17689), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17538) );
  AOI22_X1 U19683 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17585), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17537) );
  AOI22_X1 U19684 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17536) );
  NAND4_X1 U19685 ( .A1(n17539), .A2(n17538), .A3(n17537), .A4(n17536), .ZN(
        n17540) );
  NOR2_X1 U19686 ( .A1(n17541), .A2(n17540), .ZN(n17647) );
  AOI22_X1 U19687 ( .A1(n17719), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17689), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17545) );
  AOI22_X1 U19688 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17703), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n17544) );
  AOI22_X1 U19689 ( .A1(n20181), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17543) );
  AOI22_X1 U19690 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13463), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n17542) );
  NAND4_X1 U19691 ( .A1(n17545), .A2(n17544), .A3(n17543), .A4(n17542), .ZN(
        n17552) );
  AOI22_X1 U19692 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17550) );
  AOI22_X1 U19693 ( .A1(n17546), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17549) );
  AOI22_X1 U19694 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17548) );
  AOI22_X1 U19695 ( .A1(n17720), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17722), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17547) );
  NAND4_X1 U19696 ( .A1(n17550), .A2(n17549), .A3(n17548), .A4(n17547), .ZN(
        n17551) );
  NOR2_X1 U19697 ( .A1(n17552), .A2(n17551), .ZN(n17648) );
  NOR2_X1 U19698 ( .A1(n17647), .A2(n17648), .ZN(n17646) );
  AOI22_X1 U19699 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n17722), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17698), .ZN(n17564) );
  AOI22_X1 U19700 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17719), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17563) );
  AOI22_X1 U19701 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17720), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17503), .ZN(n17553) );
  OAI21_X1 U19702 ( .B1(n19049), .B2(n17655), .A(n17553), .ZN(n17560) );
  AOI22_X1 U19703 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17688), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17558) );
  AOI22_X1 U19704 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17689), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17557) );
  AOI22_X1 U19705 ( .A1(n20181), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n13463), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17556) );
  AOI22_X1 U19706 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n17714), .ZN(n17555) );
  NAND4_X1 U19707 ( .A1(n17558), .A2(n17557), .A3(n17556), .A4(n17555), .ZN(
        n17559) );
  AOI211_X1 U19708 ( .C1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .C2(n17561), .A(
        n17560), .B(n17559), .ZN(n17562) );
  NAND3_X1 U19709 ( .A1(n17564), .A2(n17563), .A3(n17562), .ZN(n17642) );
  NAND2_X1 U19710 ( .A1(n17646), .A2(n17642), .ZN(n17641) );
  NOR2_X1 U19711 ( .A1(n17637), .A2(n17641), .ZN(n17636) );
  AOI22_X1 U19712 ( .A1(n17585), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17722), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17574) );
  AOI22_X1 U19713 ( .A1(n17719), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17573) );
  AOI22_X1 U19714 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17565) );
  OAI21_X1 U19715 ( .B1(n17655), .B2(n18958), .A(n17565), .ZN(n17571) );
  AOI22_X1 U19716 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n17569) );
  AOI22_X1 U19717 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17689), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17568) );
  AOI22_X1 U19718 ( .A1(n17713), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17567) );
  AOI22_X1 U19719 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n20181), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17566) );
  NAND4_X1 U19720 ( .A1(n17569), .A2(n17568), .A3(n17567), .A4(n17566), .ZN(
        n17570) );
  AOI211_X1 U19721 ( .C1(n17688), .C2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n17571), .B(n17570), .ZN(n17572) );
  NAND3_X1 U19722 ( .A1(n17574), .A2(n17573), .A3(n17572), .ZN(n17630) );
  NAND2_X1 U19723 ( .A1(n17636), .A2(n17630), .ZN(n17629) );
  NOR2_X1 U19724 ( .A1(n17614), .A2(n17629), .ZN(n17625) );
  AOI22_X1 U19725 ( .A1(n17688), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17584) );
  AOI22_X1 U19726 ( .A1(n17698), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17583) );
  AOI22_X1 U19727 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17722), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17575) );
  OAI21_X1 U19728 ( .B1(n17655), .B2(n18876), .A(n17575), .ZN(n17581) );
  AOI22_X1 U19729 ( .A1(n17689), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17585), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17579) );
  AOI22_X1 U19730 ( .A1(n17719), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17590), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17578) );
  AOI22_X1 U19731 ( .A1(n20181), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17577) );
  AOI22_X1 U19732 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17713), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17576) );
  NAND4_X1 U19733 ( .A1(n17579), .A2(n17578), .A3(n17577), .A4(n17576), .ZN(
        n17580) );
  AOI211_X1 U19734 ( .C1(n17465), .C2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n17581), .B(n17580), .ZN(n17582) );
  NAND3_X1 U19735 ( .A1(n17584), .A2(n17583), .A3(n17582), .ZN(n17624) );
  NAND2_X1 U19736 ( .A1(n17625), .A2(n17624), .ZN(n17623) );
  NOR2_X1 U19737 ( .A1(n17618), .A2(n17623), .ZN(n17617) );
  AOI22_X1 U19738 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17589) );
  AOI22_X1 U19739 ( .A1(n17585), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17588) );
  AOI22_X1 U19740 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n20181), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17587) );
  AOI22_X1 U19741 ( .A1(n17356), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17586) );
  NAND4_X1 U19742 ( .A1(n17589), .A2(n17588), .A3(n17587), .A4(n17586), .ZN(
        n17596) );
  AOI22_X1 U19743 ( .A1(n17703), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17722), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n17594) );
  AOI22_X1 U19744 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17689), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17593) );
  AOI22_X1 U19745 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17590), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n17592) );
  AOI22_X1 U19746 ( .A1(n17688), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17591) );
  NAND4_X1 U19747 ( .A1(n17594), .A2(n17593), .A3(n17592), .A4(n17591), .ZN(
        n17595) );
  NOR2_X1 U19748 ( .A1(n17596), .A2(n17595), .ZN(n17597) );
  XOR2_X1 U19749 ( .A(n17617), .B(n17597), .Z(n20675) );
  OAI22_X1 U19750 ( .A1(n17599), .A2(n17598), .B1(n20675), .B2(n17736), .ZN(
        P3_U2673) );
  NAND2_X1 U19751 ( .A1(n20722), .A2(n17600), .ZN(n17613) );
  OR2_X1 U19752 ( .A1(n17738), .A2(n17600), .ZN(n17682) );
  AOI22_X1 U19753 ( .A1(n17689), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n17604) );
  AOI22_X1 U19754 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17603) );
  AOI22_X1 U19755 ( .A1(n20181), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17713), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n17602) );
  AOI22_X1 U19756 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17601) );
  NAND4_X1 U19757 ( .A1(n17604), .A2(n17603), .A3(n17602), .A4(n17601), .ZN(
        n17610) );
  AOI22_X1 U19758 ( .A1(n17688), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17608) );
  AOI22_X1 U19759 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17607) );
  AOI22_X1 U19760 ( .A1(n17719), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17502), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17606) );
  AOI22_X1 U19761 ( .A1(n17698), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17722), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17605) );
  NAND4_X1 U19762 ( .A1(n17608), .A2(n17607), .A3(n17606), .A4(n17605), .ZN(
        n17609) );
  NOR2_X1 U19763 ( .A1(n17610), .A2(n17609), .ZN(n20627) );
  OAI22_X1 U19764 ( .A1(n20418), .A2(n17682), .B1(n17736), .B2(n20627), .ZN(
        n17611) );
  INV_X1 U19765 ( .A(n17611), .ZN(n17612) );
  OAI21_X1 U19766 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n17613), .A(n17612), .ZN(
        P3_U2682) );
  NOR2_X1 U19767 ( .A1(n20418), .A2(n17613), .ZN(n17652) );
  NAND2_X1 U19768 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n17652), .ZN(n17645) );
  NOR2_X1 U19769 ( .A1(n20448), .A2(n17645), .ZN(n17651) );
  NAND2_X1 U19770 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17651), .ZN(n17640) );
  NAND3_X1 U19771 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n17644), .ZN(n17631) );
  AOI21_X1 U19772 ( .B1(n17614), .B2(n17629), .A(n17625), .ZN(n20693) );
  INV_X1 U19773 ( .A(n20693), .ZN(n17616) );
  NAND3_X1 U19774 ( .A1(n17631), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17736), 
        .ZN(n17615) );
  OAI221_X1 U19775 ( .B1(n17631), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17736), 
        .C2(n17616), .A(n17615), .ZN(P3_U2676) );
  NAND2_X1 U19776 ( .A1(n17736), .A2(n17631), .ZN(n17632) );
  INV_X1 U19777 ( .A(n17632), .ZN(n17626) );
  AOI21_X1 U19778 ( .B1(n17737), .B2(n17619), .A(n17626), .ZN(n17622) );
  AOI21_X1 U19779 ( .B1(n17618), .B2(n17623), .A(n17617), .ZN(n20680) );
  NOR3_X1 U19780 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n17631), .A3(n17619), .ZN(
        n17620) );
  AOI21_X1 U19781 ( .B1(n17738), .B2(n20680), .A(n17620), .ZN(n17621) );
  OAI21_X1 U19782 ( .B1(n17622), .B2(n20524), .A(n17621), .ZN(P3_U2674) );
  OAI21_X1 U19783 ( .B1(n17625), .B2(n17624), .A(n17623), .ZN(n20686) );
  OAI221_X1 U19784 ( .B1(n17626), .B2(n17737), .C1(n17626), .C2(n20497), .A(
        P3_EBX_REG_28__SCAN_IN), .ZN(n17628) );
  OR3_X1 U19785 ( .A1(n20497), .A2(n17631), .A3(P3_EBX_REG_28__SCAN_IN), .ZN(
        n17627) );
  OAI211_X1 U19786 ( .C1(n17736), .C2(n20686), .A(n17628), .B(n17627), .ZN(
        P3_U2675) );
  OAI21_X1 U19787 ( .B1(n17636), .B2(n17630), .A(n17629), .ZN(n20668) );
  NAND2_X1 U19788 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n17644), .ZN(n17635) );
  INV_X1 U19789 ( .A(n17631), .ZN(n17634) );
  INV_X1 U19790 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n17633) );
  OAI222_X1 U19791 ( .A1(n17736), .A2(n20668), .B1(n17635), .B2(n17634), .C1(
        n17633), .C2(n17632), .ZN(P3_U2677) );
  AOI21_X1 U19792 ( .B1(n17637), .B2(n17641), .A(n17636), .ZN(n20657) );
  INV_X1 U19793 ( .A(n20657), .ZN(n17639) );
  NAND3_X1 U19794 ( .A1(n17640), .A2(P3_EBX_REG_25__SCAN_IN), .A3(n17736), 
        .ZN(n17638) );
  OAI221_X1 U19795 ( .B1(n17640), .B2(P3_EBX_REG_25__SCAN_IN), .C1(n17736), 
        .C2(n17639), .A(n17638), .ZN(P3_U2678) );
  AOI21_X1 U19796 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17736), .A(n17651), .ZN(
        n17643) );
  OAI21_X1 U19797 ( .B1(n17646), .B2(n17642), .A(n17641), .ZN(n20700) );
  OAI22_X1 U19798 ( .A1(n17644), .A2(n17643), .B1(n20700), .B2(n17736), .ZN(
        P3_U2679) );
  INV_X1 U19799 ( .A(n17645), .ZN(n17668) );
  AOI21_X1 U19800 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17736), .A(n17668), .ZN(
        n17650) );
  AOI21_X1 U19801 ( .B1(n17648), .B2(n17647), .A(n17646), .ZN(n20701) );
  INV_X1 U19802 ( .A(n20701), .ZN(n17649) );
  OAI22_X1 U19803 ( .A1(n17651), .A2(n17650), .B1(n17649), .B2(n17736), .ZN(
        P3_U2680) );
  AOI21_X1 U19804 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17736), .A(n17652), .ZN(
        n17667) );
  AOI22_X1 U19805 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17665) );
  AOI22_X1 U19806 ( .A1(n17719), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17664) );
  AOI22_X1 U19807 ( .A1(n17689), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17653) );
  OAI21_X1 U19808 ( .B1(n17655), .B2(n17654), .A(n17653), .ZN(n17662) );
  AOI22_X1 U19809 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17722), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17660) );
  AOI22_X1 U19810 ( .A1(n17656), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17723), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17659) );
  AOI22_X1 U19811 ( .A1(n20181), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17713), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n17658) );
  AOI22_X1 U19812 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17657) );
  NAND4_X1 U19813 ( .A1(n17660), .A2(n17659), .A3(n17658), .A4(n17657), .ZN(
        n17661) );
  AOI211_X1 U19814 ( .C1(n17688), .C2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n17662), .B(n17661), .ZN(n17663) );
  NAND3_X1 U19815 ( .A1(n17665), .A2(n17664), .A3(n17663), .ZN(n20634) );
  INV_X1 U19816 ( .A(n20634), .ZN(n17666) );
  OAI22_X1 U19817 ( .A1(n17668), .A2(n17667), .B1(n17666), .B2(n17736), .ZN(
        P3_U2681) );
  AOI22_X1 U19818 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17689), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17678) );
  AOI22_X1 U19819 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17561), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17677) );
  AOI22_X1 U19820 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17669) );
  OAI21_X1 U19821 ( .B1(n10964), .B2(n18917), .A(n17669), .ZN(n17675) );
  AOI22_X1 U19822 ( .A1(n17703), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17722), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17673) );
  AOI22_X1 U19823 ( .A1(n17719), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17672) );
  AOI22_X1 U19824 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17713), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17671) );
  AOI22_X1 U19825 ( .A1(n20181), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17670) );
  NAND4_X1 U19826 ( .A1(n17673), .A2(n17672), .A3(n17671), .A4(n17670), .ZN(
        n17674) );
  AOI211_X1 U19827 ( .C1(n17688), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n17675), .B(n17674), .ZN(n17676) );
  NAND3_X1 U19828 ( .A1(n17678), .A2(n17677), .A3(n17676), .ZN(n20630) );
  NAND2_X1 U19829 ( .A1(n17738), .A2(n20630), .ZN(n17679) );
  OAI221_X1 U19830 ( .B1(n17682), .B2(n17681), .C1(n17682), .C2(n17680), .A(
        n17679), .ZN(P3_U2683) );
  AOI22_X1 U19831 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17687) );
  AOI22_X1 U19832 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10966), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17686) );
  AOI22_X1 U19833 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n13463), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17685) );
  AOI22_X1 U19834 ( .A1(n17683), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17684) );
  NAND4_X1 U19835 ( .A1(n17687), .A2(n17686), .A3(n17685), .A4(n17684), .ZN(
        n17695) );
  AOI22_X1 U19836 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17688), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17693) );
  AOI22_X1 U19837 ( .A1(n17719), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17692) );
  AOI22_X1 U19838 ( .A1(n17689), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17502), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17691) );
  AOI22_X1 U19839 ( .A1(n17698), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17722), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17690) );
  NAND4_X1 U19840 ( .A1(n17693), .A2(n17692), .A3(n17691), .A4(n17690), .ZN(
        n17694) );
  NOR2_X1 U19841 ( .A1(n17695), .A2(n17694), .ZN(n20651) );
  NOR2_X1 U19842 ( .A1(n17738), .A2(n17711), .ZN(n17710) );
  OAI21_X1 U19843 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17696), .A(n17710), .ZN(
        n17697) );
  OAI21_X1 U19844 ( .B1(n20651), .B2(n17736), .A(n17697), .ZN(P3_U2685) );
  AOI22_X1 U19845 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17720), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17702) );
  AOI22_X1 U19846 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17698), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17701) );
  AOI22_X1 U19847 ( .A1(n20181), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17713), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17700) );
  AOI22_X1 U19848 ( .A1(n17554), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17497), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17699) );
  NAND4_X1 U19849 ( .A1(n17702), .A2(n17701), .A3(n17700), .A4(n17699), .ZN(
        n17709) );
  AOI22_X1 U19850 ( .A1(n17703), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17707) );
  AOI22_X1 U19851 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17689), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17706) );
  AOI22_X1 U19852 ( .A1(n17688), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17722), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17705) );
  AOI22_X1 U19853 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17704) );
  NAND4_X1 U19854 ( .A1(n17707), .A2(n17706), .A3(n17705), .A4(n17704), .ZN(
        n17708) );
  NOR2_X1 U19855 ( .A1(n17709), .A2(n17708), .ZN(n20645) );
  OAI222_X1 U19856 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n20722), .B1(
        P3_EBX_REG_19__SCAN_IN), .B2(n17711), .C1(n17710), .C2(n20390), .ZN(
        n17712) );
  OAI21_X1 U19857 ( .B1(n20645), .B2(n17736), .A(n17712), .ZN(P3_U2684) );
  AOI22_X1 U19858 ( .A1(n17465), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17503), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17718) );
  AOI22_X1 U19859 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17698), .B1(
        n17502), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17717) );
  AOI22_X1 U19860 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17713), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17554), .ZN(n17716) );
  AOI22_X1 U19861 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20181), .B1(
        P3_INSTQUEUE_REG_10__1__SCAN_IN), .B2(n17714), .ZN(n17715) );
  NAND4_X1 U19862 ( .A1(n17718), .A2(n17717), .A3(n17716), .A4(n17715), .ZN(
        n17729) );
  AOI22_X1 U19863 ( .A1(n17688), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n17719), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17727) );
  AOI22_X1 U19864 ( .A1(n10966), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17689), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17726) );
  AOI22_X1 U19865 ( .A1(n17721), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17720), .ZN(n17725) );
  AOI22_X1 U19866 ( .A1(n17723), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17722), .ZN(n17724) );
  NAND4_X1 U19867 ( .A1(n17727), .A2(n17726), .A3(n17725), .A4(n17724), .ZN(
        n17728) );
  NOR2_X1 U19868 ( .A1(n17729), .A2(n17728), .ZN(n20656) );
  AOI21_X1 U19869 ( .B1(n20378), .B2(n17731), .A(n17730), .ZN(n17732) );
  AOI22_X1 U19870 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17734), .B1(n17737), 
        .B2(n17732), .ZN(n17733) );
  OAI21_X1 U19871 ( .B1(n20656), .B2(n17736), .A(n17733), .ZN(P3_U2686) );
  NOR2_X1 U19872 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n20162) );
  AOI21_X1 U19873 ( .B1(P3_EBX_REG_1__SCAN_IN), .B2(P3_EBX_REG_0__SCAN_IN), 
        .A(n20162), .ZN(n20147) );
  AOI22_X1 U19874 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(n17734), .B1(n20147), .B2(
        n17737), .ZN(n17735) );
  OAI21_X1 U19875 ( .B1(n19049), .B2(n17736), .A(n17735), .ZN(P3_U2702) );
  AOI22_X1 U19876 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17738), .B1(
        n17737), .B2(n20556), .ZN(n17739) );
  OAI21_X1 U19877 ( .B1(n17740), .B2(n20556), .A(n17739), .ZN(P3_U2703) );
  NAND2_X1 U19878 ( .A1(n21098), .A2(n21232), .ZN(n17742) );
  OAI21_X1 U19879 ( .B1(n21193), .B2(n20104), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n17741) );
  OAI21_X1 U19880 ( .B1(n17742), .B2(n21225), .A(n17741), .ZN(P3_U2634) );
  NOR2_X1 U19881 ( .A1(n20097), .A2(n18145), .ZN(n17746) );
  AOI21_X1 U19882 ( .B1(n21248), .B2(n17744), .A(n17743), .ZN(n21238) );
  NOR2_X1 U19883 ( .A1(n21238), .A2(n18715), .ZN(n17745) );
  OAI22_X1 U19884 ( .A1(n21201), .A2(n17746), .B1(n18145), .B2(n17745), .ZN(
        P3_U2863) );
  INV_X1 U19885 ( .A(n17747), .ZN(n21185) );
  NOR2_X4 U19886 ( .A1(n20559), .A2(n21247), .ZN(n18128) );
  INV_X2 U19887 ( .A(n18128), .ZN(n18140) );
  OAI22_X1 U19888 ( .A1(n17865), .A2(n20906), .B1(n18140), .B2(n20907), .ZN(
        n18024) );
  NAND2_X1 U19889 ( .A1(n18024), .A2(n20950), .ZN(n17886) );
  INV_X2 U19890 ( .A(n17886), .ZN(n17976) );
  OAI22_X1 U19891 ( .A1(n17816), .A2(n17865), .B1(n21108), .B2(n18140), .ZN(
        n17793) );
  AOI21_X1 U19892 ( .B1(n17976), .B2(n17756), .A(n17793), .ZN(n17982) );
  INV_X1 U19893 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17762) );
  NOR2_X1 U19894 ( .A1(n17750), .A2(n20150), .ZN(n17979) );
  AOI21_X1 U19895 ( .B1(n18001), .B2(n17750), .A(n10977), .ZN(n17985) );
  OAI21_X1 U19896 ( .B1(n17979), .B2(n18135), .A(n17985), .ZN(n17768) );
  INV_X2 U19897 ( .A(n19005), .ZN(n19053) );
  AOI21_X2 U19898 ( .B1(n17925), .B2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n19053), .ZN(n17894) );
  NOR3_X1 U19899 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17894), .A3(
        n17750), .ZN(n17769) );
  INV_X1 U19900 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n21126) );
  NAND3_X2 U19901 ( .A1(n21612), .A2(n18136), .A3(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n17978) );
  INV_X1 U19902 ( .A(n17751), .ZN(n17752) );
  OAI21_X1 U19903 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17979), .A(
        n17752), .ZN(n20384) );
  OAI22_X1 U19904 ( .A1(n21176), .A2(n21126), .B1(n17978), .B2(n20384), .ZN(
        n17753) );
  AOI211_X1 U19905 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n17768), .A(
        n17769), .B(n17753), .ZN(n17758) );
  AOI21_X1 U19906 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n18010), .A(
        n17842), .ZN(n17755) );
  XNOR2_X1 U19907 ( .A(n17755), .B(n17759), .ZN(n21124) );
  NOR2_X1 U19908 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17756), .ZN(
        n21123) );
  AOI22_X1 U19909 ( .A1(n18038), .A2(n21124), .B1(n17976), .B2(n21123), .ZN(
        n17757) );
  OAI211_X1 U19910 ( .C1(n17982), .C2(n17762), .A(n17758), .B(n17757), .ZN(
        P3_U2812) );
  NOR2_X1 U19911 ( .A1(n17760), .A2(n17759), .ZN(n17833) );
  NOR3_X1 U19912 ( .A1(n17923), .A2(n17762), .A3(n17761), .ZN(n17841) );
  NOR2_X1 U19913 ( .A1(n17833), .A2(n17841), .ZN(n17763) );
  XOR2_X1 U19914 ( .A(n17763), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Z(
        n21096) );
  NOR2_X1 U19915 ( .A1(n17764), .A2(n17886), .ZN(n17850) );
  INV_X1 U19916 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17844) );
  NOR3_X1 U19917 ( .A1(n17764), .A2(n17844), .A3(n20964), .ZN(n21092) );
  NOR2_X1 U19918 ( .A1(n17764), .A2(n17844), .ZN(n17765) );
  NAND2_X1 U19919 ( .A1(n21108), .A2(n17765), .ZN(n21089) );
  INV_X1 U19920 ( .A(n21089), .ZN(n17766) );
  OAI22_X1 U19921 ( .A1(n21092), .A2(n17865), .B1(n17766), .B2(n18140), .ZN(
        n17851) );
  NOR3_X1 U19922 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17894), .A3(
        n11054), .ZN(n17767) );
  AOI221_X1 U19923 ( .B1(n17769), .B2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C1(
        n17768), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17767), .ZN(
        n17770) );
  NAND2_X1 U19924 ( .A1(n21137), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n21094) );
  OAI211_X1 U19925 ( .C1(n17978), .C2(n20399), .A(n17770), .B(n21094), .ZN(
        n17771) );
  AOI221_X1 U19926 ( .B1(n17850), .B2(n17844), .C1(n17851), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n17771), .ZN(n17772) );
  OAI21_X1 U19927 ( .B1(n21096), .B2(n18055), .A(n17772), .ZN(P3_U2811) );
  INV_X1 U19928 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17811) );
  NAND3_X1 U19929 ( .A1(n17773), .A2(n18010), .A3(n20912), .ZN(n18029) );
  INV_X1 U19930 ( .A(n18029), .ZN(n18014) );
  NAND2_X1 U19931 ( .A1(n20923), .A2(n18014), .ZN(n17810) );
  NOR2_X1 U19932 ( .A1(n17811), .A2(n17810), .ZN(n17774) );
  NAND2_X1 U19933 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17774), .ZN(
        n17995) );
  OAI22_X1 U19934 ( .A1(n20938), .A2(n17995), .B1(n17776), .B2(n18030), .ZN(
        n17777) );
  XOR2_X1 U19935 ( .A(n20958), .B(n17777), .Z(n20971) );
  NOR2_X1 U19936 ( .A1(n17894), .A2(n17778), .ZN(n17789) );
  NOR2_X1 U19937 ( .A1(n17778), .A2(n20150), .ZN(n17988) );
  AOI21_X1 U19938 ( .B1(n18001), .B2(n17778), .A(n10977), .ZN(n17991) );
  OAI21_X1 U19939 ( .B1(n17988), .B2(n18135), .A(n17991), .ZN(n17787) );
  NAND2_X1 U19940 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17988), .ZN(
        n20349) );
  OAI21_X1 U19941 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17988), .A(
        n20349), .ZN(n20335) );
  NAND2_X1 U19942 ( .A1(n21137), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n20969) );
  OAI21_X1 U19943 ( .B1(n17978), .B2(n20335), .A(n20969), .ZN(n17779) );
  AOI221_X1 U19944 ( .B1(n17789), .B2(n20339), .C1(n17787), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17779), .ZN(n17783) );
  NOR2_X1 U19945 ( .A1(n17816), .A2(n17865), .ZN(n17781) );
  OAI21_X1 U19946 ( .B1(n20962), .B2(n18140), .A(n20958), .ZN(n17780) );
  AOI22_X1 U19947 ( .A1(n20959), .A2(n17781), .B1(n17793), .B2(n17780), .ZN(
        n17782) );
  OAI211_X1 U19948 ( .C1(n20971), .C2(n18055), .A(n17783), .B(n17782), .ZN(
        P3_U2815) );
  AOI22_X1 U19949 ( .A1(n18010), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n21135), .B2(n17923), .ZN(n17784) );
  XNOR2_X1 U19950 ( .A(n17785), .B(n17784), .ZN(n21143) );
  INV_X1 U19951 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n20365) );
  INV_X1 U19952 ( .A(n17978), .ZN(n17961) );
  NAND2_X1 U19953 ( .A1(n17974), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17980) );
  INV_X1 U19954 ( .A(n17980), .ZN(n17786) );
  AOI21_X1 U19955 ( .B1(n20357), .B2(n20349), .A(n17786), .ZN(n20361) );
  AOI22_X1 U19956 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17787), .B1(
        n17961), .B2(n20361), .ZN(n17791) );
  OAI211_X1 U19957 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17789), .B(n17788), .ZN(n17790) );
  OAI211_X1 U19958 ( .C1(n20365), .C2(n21176), .A(n17791), .B(n17790), .ZN(
        n17792) );
  AOI221_X1 U19959 ( .B1(n17976), .B2(n21135), .C1(n17793), .C2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n17792), .ZN(n17794) );
  OAI21_X1 U19960 ( .B1(n18055), .B2(n21143), .A(n17794), .ZN(P3_U2814) );
  NOR2_X1 U19961 ( .A1(n20906), .A2(n20937), .ZN(n20924) );
  NOR2_X1 U19962 ( .A1(n20907), .A2(n20937), .ZN(n20928) );
  OAI22_X1 U19963 ( .A1(n17865), .A2(n20924), .B1(n18140), .B2(n20928), .ZN(
        n17813) );
  INV_X1 U19964 ( .A(n17813), .ZN(n17803) );
  NOR2_X1 U19965 ( .A1(n17894), .A2(n17795), .ZN(n17805) );
  INV_X1 U19966 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n20291) );
  NOR2_X1 U19967 ( .A1(n17795), .A2(n20150), .ZN(n18002) );
  INV_X1 U19968 ( .A(n18135), .ZN(n17898) );
  AOI21_X1 U19969 ( .B1(n18001), .B2(n17795), .A(n17898), .ZN(n17796) );
  OAI21_X1 U19970 ( .B1(n18002), .B2(n17796), .A(n18136), .ZN(n17808) );
  NAND2_X1 U19971 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n18002), .ZN(
        n17804) );
  OAI21_X1 U19972 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18002), .A(
        n17804), .ZN(n20296) );
  NAND2_X1 U19973 ( .A1(n21137), .A2(P3_REIP_REG_12__SCAN_IN), .ZN(n20932) );
  OAI21_X1 U19974 ( .B1(n17978), .B2(n20296), .A(n20932), .ZN(n17797) );
  AOI221_X1 U19975 ( .B1(n17805), .B2(n20291), .C1(n17808), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17797), .ZN(n17802) );
  INV_X1 U19976 ( .A(n18024), .ZN(n18042) );
  NOR2_X1 U19977 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18042), .ZN(
        n17800) );
  INV_X1 U19978 ( .A(n17810), .ZN(n17798) );
  NOR3_X1 U19979 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18025), .A3(
        n18030), .ZN(n17809) );
  NOR2_X1 U19980 ( .A1(n17798), .A2(n17809), .ZN(n17799) );
  XOR2_X1 U19981 ( .A(n17811), .B(n17799), .Z(n20931) );
  AOI22_X1 U19982 ( .A1(n20923), .A2(n17800), .B1(n18038), .B2(n20931), .ZN(
        n17801) );
  OAI211_X1 U19983 ( .C1(n17803), .C2(n17811), .A(n17802), .B(n17801), .ZN(
        P3_U2818) );
  INV_X1 U19984 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n21149) );
  NAND2_X1 U19985 ( .A1(n20929), .A2(n21149), .ZN(n21156) );
  NOR2_X1 U19986 ( .A1(n21176), .A2(n20344), .ZN(n21152) );
  INV_X1 U19987 ( .A(n17804), .ZN(n20302) );
  NAND2_X1 U19988 ( .A1(n17990), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17989) );
  OAI21_X1 U19989 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n20302), .A(
        n17989), .ZN(n20317) );
  OAI211_X1 U19990 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17805), .B(n20313), .ZN(n17806) );
  OAI21_X1 U19991 ( .B1(n17978), .B2(n20317), .A(n17806), .ZN(n17807) );
  AOI211_X1 U19992 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n17808), .A(
        n21152), .B(n17807), .ZN(n17815) );
  NAND2_X1 U19993 ( .A1(n17809), .A2(n17811), .ZN(n17996) );
  OAI21_X1 U19994 ( .B1(n17811), .B2(n17810), .A(n17996), .ZN(n17812) );
  XOR2_X1 U19995 ( .A(n17812), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n21154) );
  AOI22_X1 U19996 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17813), .B1(
        n18038), .B2(n21154), .ZN(n17814) );
  OAI211_X1 U19997 ( .C1(n18042), .C2(n21156), .A(n17815), .B(n17814), .ZN(
        P3_U2817) );
  NAND2_X1 U19998 ( .A1(n17817), .A2(n17976), .ZN(n17829) );
  NAND2_X1 U19999 ( .A1(n17817), .A2(n17816), .ZN(n20802) );
  NAND2_X1 U20000 ( .A1(n17817), .A2(n21108), .ZN(n20803) );
  AOI22_X1 U20001 ( .A1(n18052), .A2(n20802), .B1(n18128), .B2(n20803), .ZN(
        n17839) );
  INV_X1 U20002 ( .A(n17818), .ZN(n17819) );
  OAI21_X1 U20003 ( .B1(n17820), .B2(n17819), .A(n17840), .ZN(n17854) );
  XOR2_X1 U20004 ( .A(n20974), .B(n17854), .Z(n20978) );
  INV_X1 U20005 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17822) );
  INV_X1 U20006 ( .A(n17894), .ZN(n17936) );
  NAND2_X1 U20007 ( .A1(n13386), .A2(n17936), .ZN(n17830) );
  AOI221_X1 U20008 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C1(n17822), .C2(n17821), .A(
        n17830), .ZN(n17827) );
  OAI22_X1 U20009 ( .A1(n17823), .A2(n18135), .B1(n13386), .B2(n18096), .ZN(
        n17824) );
  NOR2_X1 U20010 ( .A1(n10977), .A2(n17824), .ZN(n17845) );
  OAI21_X1 U20011 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17977), .A(
        n17845), .ZN(n17832) );
  AOI22_X1 U20012 ( .A1(n21137), .A2(P3_REIP_REG_22__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n17832), .ZN(n17825) );
  OAI21_X1 U20013 ( .B1(n20435), .B2(n17978), .A(n17825), .ZN(n17826) );
  AOI211_X1 U20014 ( .C1(n20978), .C2(n18038), .A(n17827), .B(n17826), .ZN(
        n17828) );
  OAI221_X1 U20015 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17829), 
        .C1(n20974), .C2(n17839), .A(n17828), .ZN(P3_U2808) );
  INV_X1 U20016 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n20425) );
  NOR2_X1 U20017 ( .A1(n21176), .A2(n20425), .ZN(n20810) );
  OAI22_X1 U20018 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n17830), .B1(
        n17978), .B2(n20417), .ZN(n17831) );
  AOI211_X1 U20019 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(n17832), .A(
        n20810), .B(n17831), .ZN(n17838) );
  INV_X1 U20020 ( .A(n20806), .ZN(n17835) );
  NOR2_X1 U20021 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17834) );
  AOI22_X1 U20022 ( .A1(n17835), .A2(n17841), .B1(n17834), .B2(n17833), .ZN(
        n17836) );
  XOR2_X1 U20023 ( .A(n20807), .B(n17836), .Z(n20797) );
  NOR2_X1 U20024 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n20806), .ZN(
        n20811) );
  AOI22_X1 U20025 ( .A1(n18038), .A2(n20797), .B1(n20811), .B2(n17850), .ZN(
        n17837) );
  OAI211_X1 U20026 ( .C1(n17839), .C2(n20807), .A(n17838), .B(n17837), .ZN(
        P3_U2809) );
  OAI221_X1 U20027 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17842), 
        .C1(n17844), .C2(n17841), .A(n17840), .ZN(n17843) );
  XOR2_X1 U20028 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17843), .Z(
        n21107) );
  NOR2_X1 U20029 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17844), .ZN(
        n21103) );
  AOI221_X1 U20030 ( .B1(n17847), .B2(n17846), .C1(n19005), .C2(n17846), .A(
        n17845), .ZN(n17849) );
  NAND2_X1 U20031 ( .A1(n21137), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n21105) );
  OAI221_X1 U20032 ( .B1(n20410), .B2(n17978), .C1(n20410), .C2(n17977), .A(
        n21105), .ZN(n17848) );
  AOI211_X1 U20033 ( .C1(n21103), .C2(n17850), .A(n17849), .B(n17848), .ZN(
        n17853) );
  NAND2_X1 U20034 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17851), .ZN(
        n17852) );
  OAI211_X1 U20035 ( .C1(n21107), .C2(n18055), .A(n17853), .B(n17852), .ZN(
        P3_U2810) );
  AOI221_X1 U20036 ( .B1(n17923), .B2(n17855), .C1(n20974), .C2(n17855), .A(
        n17854), .ZN(n17856) );
  XOR2_X1 U20037 ( .A(n21071), .B(n17856), .Z(n21078) );
  NOR3_X1 U20038 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17894), .A3(
        n17857), .ZN(n17862) );
  OAI21_X1 U20039 ( .B1(n17872), .B2(n19005), .A(n18136), .ZN(n17858) );
  AOI21_X1 U20040 ( .B1(n17898), .B2(n17859), .A(n17858), .ZN(n17871) );
  OAI22_X1 U20041 ( .A1(n17871), .A2(n17860), .B1(n20444), .B2(n17978), .ZN(
        n17861) );
  AOI211_X1 U20042 ( .C1(P3_REIP_REG_23__SCAN_IN), .C2(n21137), .A(n17862), 
        .B(n17861), .ZN(n17869) );
  NAND2_X1 U20043 ( .A1(n18052), .A2(n21066), .ZN(n17863) );
  NAND2_X1 U20044 ( .A1(n18128), .A2(n21068), .ZN(n17864) );
  OAI22_X1 U20045 ( .A1(n17863), .A2(n20802), .B1(n17864), .B2(n20803), .ZN(
        n17867) );
  OAI21_X1 U20046 ( .B1(n17866), .B2(n17865), .A(n17864), .ZN(n17890) );
  AOI22_X1 U20047 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17867), .B1(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17890), .ZN(n17868) );
  OAI211_X1 U20048 ( .C1(n18055), .C2(n21078), .A(n17869), .B(n17868), .ZN(
        P3_U2807) );
  XOR2_X1 U20049 ( .A(n20986), .B(n17870), .Z(n20987) );
  OAI21_X1 U20050 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n18135), .A(
        n17871), .ZN(n17885) );
  INV_X1 U20051 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n20468) );
  NAND2_X1 U20052 ( .A1(n17872), .A2(n17936), .ZN(n17882) );
  AOI221_X1 U20053 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C1(n20468), .C2(n20454), .A(
        n17882), .ZN(n17874) );
  OAI22_X1 U20054 ( .A1(n21176), .A2(n20471), .B1(n20477), .B2(n17978), .ZN(
        n17873) );
  AOI211_X1 U20055 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17885), .A(
        n17874), .B(n17873), .ZN(n17879) );
  XOR2_X1 U20056 ( .A(n20986), .B(n17875), .Z(n20990) );
  INV_X1 U20057 ( .A(n17876), .ZN(n17921) );
  OAI21_X1 U20058 ( .B1(n17923), .B2(n17922), .A(n17921), .ZN(n17877) );
  XOR2_X1 U20059 ( .A(n17877), .B(n20986), .Z(n20991) );
  AOI22_X1 U20060 ( .A1(n18052), .A2(n20990), .B1(n18038), .B2(n20991), .ZN(
        n17878) );
  OAI211_X1 U20061 ( .C1(n18140), .C2(n20987), .A(n17879), .B(n17878), .ZN(
        P3_U2805) );
  AOI21_X1 U20062 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17881), .A(
        n17880), .ZN(n21087) );
  INV_X1 U20063 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n20465) );
  NOR2_X1 U20064 ( .A1(n21176), .A2(n20465), .ZN(n17884) );
  OAI22_X1 U20065 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n17882), .B1(
        n17978), .B2(n20462), .ZN(n17883) );
  AOI211_X1 U20066 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(n17885), .A(
        n17884), .B(n17883), .ZN(n17892) );
  NOR2_X1 U20067 ( .A1(n17887), .A2(n17886), .ZN(n17889) );
  AOI22_X1 U20068 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17890), .B1(
        n17889), .B2(n17888), .ZN(n17891) );
  OAI211_X1 U20069 ( .C1(n21087), .C2(n18055), .A(n17892), .B(n17891), .ZN(
        P3_U2806) );
  NOR3_X1 U20070 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17894), .A3(
        n17893), .ZN(n17916) );
  OAI21_X1 U20071 ( .B1(n17895), .B2(n18096), .A(n18136), .ZN(n17896) );
  AOI21_X1 U20072 ( .B1(n17898), .B2(n17897), .A(n17896), .ZN(n17926) );
  OAI21_X1 U20073 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17977), .A(
        n17926), .ZN(n17914) );
  NAND2_X1 U20074 ( .A1(n21137), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17901) );
  INV_X1 U20075 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n20510) );
  NAND3_X1 U20076 ( .A1(n17899), .A2(n20510), .A3(n17936), .ZN(n17900) );
  OAI211_X1 U20077 ( .C1(n20516), .C2(n17978), .A(n17901), .B(n17900), .ZN(
        n17902) );
  AOI221_X1 U20078 ( .B1(n17916), .B2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C1(
        n17914), .C2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17902), .ZN(
        n17912) );
  AOI22_X1 U20079 ( .A1(n18052), .A2(n21009), .B1(n18128), .B2(n21011), .ZN(
        n17928) );
  NAND2_X1 U20080 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17928), .ZN(
        n17917) );
  OAI211_X1 U20081 ( .C1(n18052), .C2(n18128), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n17917), .ZN(n17911) );
  NAND3_X1 U20082 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17903), .A3(
        n17976), .ZN(n17927) );
  NOR2_X1 U20083 ( .A1(n17904), .A2(n17927), .ZN(n17951) );
  NAND3_X1 U20084 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17951), .A3(
        n17905), .ZN(n17910) );
  OAI211_X1 U20085 ( .C1(n17908), .C2(n17907), .A(n18038), .B(n17906), .ZN(
        n17909) );
  NAND4_X1 U20086 ( .A1(n17912), .A2(n17911), .A3(n17910), .A4(n17909), .ZN(
        P3_U2802) );
  AOI22_X1 U20087 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17914), .B1(
        n17913), .B2(n17961), .ZN(n17920) );
  OAI21_X1 U20088 ( .B1(n18010), .B2(n11008), .A(n17915), .ZN(n21018) );
  AOI21_X1 U20089 ( .B1(n18038), .B2(n21018), .A(n17916), .ZN(n17919) );
  OAI21_X1 U20090 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17951), .A(
        n17917), .ZN(n17918) );
  NAND2_X1 U20091 ( .A1(n21137), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n21019) );
  NAND4_X1 U20092 ( .A1(n17920), .A2(n17919), .A3(n17918), .A4(n21019), .ZN(
        P3_U2803) );
  OAI221_X1 U20093 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17923), 
        .C1(n20986), .C2(n17922), .A(n17921), .ZN(n17924) );
  XOR2_X1 U20094 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n17924), .Z(
        n21007) );
  INV_X1 U20095 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n20493) );
  NOR2_X1 U20096 ( .A1(n21176), .A2(n20493), .ZN(n21005) );
  AOI21_X1 U20097 ( .B1(n17978), .B2(n17977), .A(n20490), .ZN(n17933) );
  AOI221_X1 U20098 ( .B1(n11061), .B2(n20485), .C1(n19005), .C2(n20485), .A(
        n17926), .ZN(n17932) );
  NOR2_X1 U20099 ( .A1(n20986), .A2(n17927), .ZN(n17930) );
  INV_X1 U20100 ( .A(n17928), .ZN(n17929) );
  MUX2_X1 U20101 ( .A(n17930), .B(n17929), .S(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .Z(n17931) );
  NOR4_X1 U20102 ( .A1(n21005), .A2(n17933), .A3(n17932), .A4(n17931), .ZN(
        n17934) );
  OAI21_X1 U20103 ( .B1(n18055), .B2(n21007), .A(n17934), .ZN(P3_U2804) );
  INV_X1 U20104 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n21052) );
  INV_X1 U20105 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n21033) );
  INV_X1 U20106 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21049) );
  NOR2_X1 U20107 ( .A1(n21033), .A2(n21049), .ZN(n21053) );
  NAND2_X1 U20108 ( .A1(n21053), .A2(n21030), .ZN(n17935) );
  XNOR2_X1 U20109 ( .A(n21052), .B(n17935), .ZN(n21057) );
  NAND2_X1 U20110 ( .A1(n21137), .A2(P3_REIP_REG_31__SCAN_IN), .ZN(n21063) );
  INV_X1 U20111 ( .A(n21063), .ZN(n17943) );
  NAND2_X1 U20112 ( .A1(n17937), .A2(n17936), .ZN(n17956) );
  XOR2_X1 U20113 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(n20538), .Z(
        n17941) );
  NOR2_X1 U20114 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17977), .ZN(
        n17960) );
  OAI22_X1 U20115 ( .A1(n18135), .A2(n17938), .B1(n19005), .B2(n17937), .ZN(
        n17939) );
  OR2_X1 U20116 ( .A1(n17939), .A2(n10977), .ZN(n17971) );
  NOR2_X1 U20117 ( .A1(n17960), .A2(n17971), .ZN(n17955) );
  OAI22_X1 U20118 ( .A1(n17956), .A2(n17941), .B1(n17940), .B2(n17955), .ZN(
        n17942) );
  AOI211_X1 U20119 ( .C1(n10967), .C2(n17961), .A(n17943), .B(n17942), .ZN(
        n17949) );
  NAND2_X1 U20120 ( .A1(n17945), .A2(n17944), .ZN(n17965) );
  OAI33_X1 U20121 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n17965), .B1(n21049), .B2(
        n17964), .B3(n21033), .ZN(n17946) );
  XNOR2_X1 U20122 ( .A(n21052), .B(n17946), .ZN(n21061) );
  AND2_X1 U20123 ( .A1(n17963), .A2(n21053), .ZN(n17947) );
  XNOR2_X1 U20124 ( .A(n21052), .B(n17947), .ZN(n21060) );
  AOI22_X1 U20125 ( .A1(n18038), .A2(n21061), .B1(n18052), .B2(n21060), .ZN(
        n17948) );
  OAI211_X1 U20126 ( .C1(n21057), .C2(n18140), .A(n17949), .B(n17948), .ZN(
        P3_U2799) );
  NOR2_X1 U20127 ( .A1(n17950), .A2(n21033), .ZN(n21039) );
  NAND2_X1 U20128 ( .A1(n21039), .A2(n17951), .ZN(n17959) );
  NAND2_X1 U20129 ( .A1(n17952), .A2(n21039), .ZN(n21022) );
  AOI22_X1 U20130 ( .A1(n18052), .A2(n21022), .B1(n18128), .B2(n21023), .ZN(
        n17968) );
  AOI22_X1 U20131 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n17964), .B1(
        n17965), .B2(n21033), .ZN(n17953) );
  XOR2_X1 U20132 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n17953), .Z(
        n21047) );
  INV_X1 U20133 ( .A(n21176), .ZN(n21167) );
  AOI22_X1 U20134 ( .A1(n21167), .A2(P3_REIP_REG_30__SCAN_IN), .B1(n20536), 
        .B2(n17961), .ZN(n17954) );
  OAI221_X1 U20135 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n17956), .C1(
        n20538), .C2(n17955), .A(n17954), .ZN(n17957) );
  AOI21_X1 U20136 ( .B1(n18038), .B2(n21047), .A(n17957), .ZN(n17958) );
  OAI221_X1 U20137 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n17959), 
        .C1(n21049), .C2(n17968), .A(n17958), .ZN(P3_U2800) );
  NOR2_X1 U20138 ( .A1(n17961), .A2(n17960), .ZN(n17973) );
  OAI21_X1 U20139 ( .B1(n17962), .B2(n19005), .A(n20523), .ZN(n17970) );
  INV_X1 U20140 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n20528) );
  NOR2_X1 U20141 ( .A1(n21176), .A2(n20528), .ZN(n21025) );
  AOI211_X1 U20142 ( .C1(n21030), .C2(n18128), .A(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B(n17963), .ZN(n17967) );
  NAND2_X1 U20143 ( .A1(n17965), .A2(n17964), .ZN(n17966) );
  XOR2_X1 U20144 ( .A(n17966), .B(n21033), .Z(n21036) );
  OAI22_X1 U20145 ( .A1(n17968), .A2(n17967), .B1(n21036), .B2(n18055), .ZN(
        n17969) );
  AOI211_X1 U20146 ( .C1(n17971), .C2(n17970), .A(n21025), .B(n17969), .ZN(
        n17972) );
  OAI21_X1 U20147 ( .B1(n20531), .B2(n17973), .A(n17972), .ZN(P3_U2801) );
  AOI21_X1 U20148 ( .B1(n17974), .B2(n19053), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17986) );
  OAI21_X1 U20149 ( .B1(n11053), .B2(n21121), .A(n17975), .ZN(n21130) );
  AOI21_X1 U20150 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17976), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17981) );
  AOI21_X1 U20151 ( .B1(n11133), .B2(n17980), .A(n17979), .ZN(n20371) );
  INV_X1 U20152 ( .A(n20371), .ZN(n20369) );
  OAI22_X1 U20153 ( .A1(n17982), .A2(n17981), .B1(n18122), .B2(n20369), .ZN(
        n17983) );
  AOI21_X1 U20154 ( .B1(n18038), .B2(n21130), .A(n17983), .ZN(n17984) );
  NAND2_X1 U20155 ( .A1(n21137), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n21133) );
  OAI211_X1 U20156 ( .C1(n17986), .C2(n17985), .A(n17984), .B(n21133), .ZN(
        P3_U2813) );
  OAI21_X1 U20157 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17987), .A(
        n20962), .ZN(n20941) );
  INV_X1 U20158 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n20331) );
  AOI21_X1 U20159 ( .B1(n20331), .B2(n17989), .A(n17988), .ZN(n20324) );
  AOI21_X1 U20160 ( .B1(n17990), .B2(n19053), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17992) );
  NAND2_X1 U20161 ( .A1(n21137), .A2(P3_REIP_REG_14__SCAN_IN), .ZN(n20947) );
  OAI21_X1 U20162 ( .B1(n17992), .B2(n17991), .A(n20947), .ZN(n17993) );
  AOI21_X1 U20163 ( .B1(n20324), .B2(n18129), .A(n17993), .ZN(n17999) );
  AOI21_X1 U20164 ( .B1(n20938), .B2(n17994), .A(n20959), .ZN(n20945) );
  OAI21_X1 U20165 ( .B1(n17996), .B2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n17995), .ZN(n17997) );
  XOR2_X1 U20166 ( .A(n17997), .B(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(
        n20946) );
  AOI22_X1 U20167 ( .A1(n18052), .A2(n20945), .B1(n18038), .B2(n20946), .ZN(
        n17998) );
  OAI211_X1 U20168 ( .C1(n18140), .C2(n20941), .A(n17999), .B(n17998), .ZN(
        P3_U2816) );
  AOI22_X1 U20169 ( .A1(n20907), .A2(n18128), .B1(n18052), .B2(n20906), .ZN(
        n18040) );
  OAI22_X1 U20170 ( .A1(n20916), .A2(n18029), .B1(n18025), .B2(n18030), .ZN(
        n18000) );
  XOR2_X1 U20171 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18000), .Z(
        n20918) );
  AOI211_X1 U20172 ( .C1(n20916), .C2(n18009), .A(n18042), .B(n20923), .ZN(
        n18007) );
  NAND2_X1 U20173 ( .A1(n20264), .A2(n19053), .ZN(n18017) );
  NOR2_X1 U20174 ( .A1(n10977), .A2(n18001), .ZN(n18069) );
  INV_X1 U20175 ( .A(n18069), .ZN(n18130) );
  NAND3_X1 U20176 ( .A1(n18130), .A2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A3(
        n18017), .ZN(n18005) );
  INV_X1 U20177 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n18003) );
  NAND2_X1 U20178 ( .A1(n20264), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18018) );
  AOI21_X1 U20179 ( .B1(n18003), .B2(n18018), .A(n18002), .ZN(n20278) );
  AOI22_X1 U20180 ( .A1(n21137), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n20278), 
        .B2(n18129), .ZN(n18004) );
  OAI211_X1 U20181 ( .C1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n18017), .A(
        n18005), .B(n18004), .ZN(n18006) );
  AOI211_X1 U20182 ( .C1(n18038), .C2(n20918), .A(n18007), .B(n18006), .ZN(
        n18008) );
  OAI21_X1 U20183 ( .B1(n18040), .B2(n18009), .A(n18008), .ZN(P3_U2819) );
  NAND2_X1 U20184 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18028), .ZN(
        n21164) );
  OAI21_X1 U20185 ( .B1(n18010), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n18029), .ZN(n18011) );
  OAI211_X1 U20186 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18012), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n18011), .ZN(n18013) );
  OAI21_X1 U20187 ( .B1(n18014), .B2(n21164), .A(n18013), .ZN(n18015) );
  AOI21_X1 U20188 ( .B1(n18016), .B2(n18030), .A(n18015), .ZN(n21157) );
  NOR2_X1 U20189 ( .A1(n21176), .A2(n20263), .ZN(n18023) );
  INV_X1 U20190 ( .A(n18017), .ZN(n18021) );
  INV_X1 U20191 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n18034) );
  NOR2_X1 U20192 ( .A1(n18046), .A2(n19005), .ZN(n18057) );
  NAND3_X1 U20193 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(n18057), .ZN(n18033) );
  NOR2_X1 U20194 ( .A1(n18034), .A2(n18033), .ZN(n18032) );
  AOI21_X1 U20195 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18130), .A(
        n18032), .ZN(n18020) );
  NAND3_X1 U20196 ( .A1(n18047), .A2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20250) );
  NOR2_X1 U20197 ( .A1(n18034), .A2(n20250), .ZN(n18019) );
  OAI21_X1 U20198 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18019), .A(
        n18018), .ZN(n20268) );
  OAI22_X1 U20199 ( .A1(n18021), .A2(n18020), .B1(n18122), .B2(n20268), .ZN(
        n18022) );
  AOI211_X1 U20200 ( .C1(n21157), .C2(n18038), .A(n18023), .B(n18022), .ZN(
        n18027) );
  NAND3_X1 U20201 ( .A1(n20916), .A2(n18025), .A3(n18024), .ZN(n18026) );
  OAI211_X1 U20202 ( .C1(n18040), .C2(n18028), .A(n18027), .B(n18026), .ZN(
        P3_U2820) );
  NAND2_X1 U20203 ( .A1(n18030), .A2(n18029), .ZN(n18031) );
  XNOR2_X1 U20204 ( .A(n18041), .B(n18031), .ZN(n21165) );
  AOI211_X1 U20205 ( .C1(n18033), .C2(n18034), .A(n18069), .B(n18032), .ZN(
        n18037) );
  INV_X1 U20206 ( .A(n20250), .ZN(n18035) );
  AOI22_X1 U20207 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n20250), .B1(
        n18035), .B2(n18034), .ZN(n20258) );
  INV_X1 U20208 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18221) );
  OAI22_X1 U20209 ( .A1(n18122), .A2(n20258), .B1(n21176), .B2(n18221), .ZN(
        n18036) );
  AOI211_X1 U20210 ( .C1(n18038), .C2(n21165), .A(n18037), .B(n18036), .ZN(
        n18039) );
  OAI221_X1 U20211 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18042), .C1(
        n18041), .C2(n18040), .A(n18039), .ZN(P3_U2821) );
  OAI21_X1 U20212 ( .B1(n18045), .B2(n18044), .A(n18043), .ZN(n20902) );
  OAI21_X1 U20213 ( .B1(n11136), .B2(n18096), .A(n18136), .ZN(n18064) );
  NOR2_X1 U20214 ( .A1(n21176), .A2(n20239), .ZN(n20896) );
  INV_X1 U20215 ( .A(n18047), .ZN(n20236) );
  NOR2_X1 U20216 ( .A1(n20236), .A2(n20150), .ZN(n18056) );
  OAI21_X1 U20217 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18056), .A(
        n20250), .ZN(n20238) );
  INV_X1 U20218 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n20242) );
  OAI221_X1 U20219 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18047), .C1(
        n20242), .C2(n20235), .A(n19053), .ZN(n18048) );
  OAI21_X1 U20220 ( .B1(n18122), .B2(n20238), .A(n18048), .ZN(n18049) );
  AOI211_X1 U20221 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n18064), .A(
        n20896), .B(n18049), .ZN(n18054) );
  AOI21_X1 U20222 ( .B1(n18051), .B2(n21172), .A(n18050), .ZN(n20897) );
  AOI22_X1 U20223 ( .A1(n18052), .A2(n20902), .B1(n18128), .B2(n20897), .ZN(
        n18053) );
  OAI211_X1 U20224 ( .C1(n18055), .C2(n20902), .A(n18054), .B(n18053), .ZN(
        P3_U2822) );
  INV_X1 U20225 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n20225) );
  NAND2_X1 U20226 ( .A1(n11136), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n20219) );
  AOI21_X1 U20227 ( .B1(n20235), .B2(n20219), .A(n18056), .ZN(n20221) );
  AOI22_X1 U20228 ( .A1(n20221), .A2(n18129), .B1(n18057), .B2(n20235), .ZN(
        n18066) );
  INV_X1 U20229 ( .A(n18081), .ZN(n18139) );
  OAI21_X1 U20230 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n18059), .A(
        n18058), .ZN(n20892) );
  NAND2_X1 U20231 ( .A1(n18061), .A2(n18060), .ZN(n18062) );
  XOR2_X1 U20232 ( .A(n18062), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n20887) );
  OAI22_X1 U20233 ( .A1(n18139), .A2(n20892), .B1(n18140), .B2(n20887), .ZN(
        n18063) );
  AOI21_X1 U20234 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18064), .A(
        n18063), .ZN(n18065) );
  OAI211_X1 U20235 ( .C1(n21176), .C2(n20225), .A(n18066), .B(n18065), .ZN(
        P3_U2823) );
  NAND2_X1 U20236 ( .A1(n18070), .A2(n19053), .ZN(n18078) );
  AOI21_X1 U20237 ( .B1(n20884), .B2(n18068), .A(n18067), .ZN(n20877) );
  AOI22_X1 U20238 ( .A1(n21137), .A2(P3_REIP_REG_6__SCAN_IN), .B1(n18128), 
        .B2(n20877), .ZN(n18077) );
  AOI21_X1 U20239 ( .B1(n19053), .B2(n18070), .A(n18069), .ZN(n18087) );
  NAND2_X1 U20240 ( .A1(n18070), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18079) );
  INV_X1 U20241 ( .A(n18079), .ZN(n18071) );
  OAI21_X1 U20242 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18071), .A(
        n20219), .ZN(n20208) );
  OAI21_X1 U20243 ( .B1(n18074), .B2(n18073), .A(n18072), .ZN(n20882) );
  OAI22_X1 U20244 ( .A1(n18122), .A2(n20208), .B1(n18139), .B2(n20882), .ZN(
        n18075) );
  AOI21_X1 U20245 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18087), .A(
        n18075), .ZN(n18076) );
  OAI211_X1 U20246 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n18078), .A(
        n18077), .B(n18076), .ZN(P3_U2824) );
  NOR2_X1 U20247 ( .A1(n18085), .A2(n20150), .ZN(n18090) );
  OAI21_X1 U20248 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n18090), .A(
        n18079), .ZN(n20198) );
  XOR2_X1 U20249 ( .A(n18080), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(
        n20869) );
  AOI22_X1 U20250 ( .A1(n21137), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18081), 
        .B2(n20869), .ZN(n18089) );
  AOI21_X1 U20251 ( .B1(n18084), .B2(n18083), .A(n18082), .ZN(n20868) );
  OAI21_X1 U20252 ( .B1(n10977), .B2(n18085), .A(n20206), .ZN(n18086) );
  AOI22_X1 U20253 ( .A1(n18128), .A2(n20868), .B1(n18087), .B2(n18086), .ZN(
        n18088) );
  OAI211_X1 U20254 ( .C1(n18122), .C2(n20198), .A(n18089), .B(n18088), .ZN(
        P3_U2825) );
  AND2_X1 U20255 ( .A1(n18097), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n18109) );
  INV_X1 U20256 ( .A(n18090), .ZN(n20188) );
  OAI21_X1 U20257 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18109), .A(
        n20188), .ZN(n20191) );
  NOR2_X1 U20258 ( .A1(n19005), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n18095) );
  OAI21_X1 U20259 ( .B1(n18093), .B2(n18092), .A(n18091), .ZN(n20856) );
  OAI22_X1 U20260 ( .A1(n21176), .A2(n20186), .B1(n18139), .B2(n20856), .ZN(
        n18094) );
  AOI21_X1 U20261 ( .B1(n18095), .B2(n18097), .A(n18094), .ZN(n18102) );
  OAI21_X1 U20262 ( .B1(n18097), .B2(n18096), .A(n18136), .ZN(n18113) );
  AOI21_X1 U20263 ( .B1(n18100), .B2(n18099), .A(n18098), .ZN(n20857) );
  AOI22_X1 U20264 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n18113), .B1(
        n18128), .B2(n20857), .ZN(n18101) );
  OAI211_X1 U20265 ( .C1(n18122), .C2(n20191), .A(n18102), .B(n18101), .ZN(
        P3_U2826) );
  OAI21_X1 U20266 ( .B1(n18105), .B2(n18104), .A(n18103), .ZN(n20851) );
  AOI21_X1 U20267 ( .B1(n18108), .B2(n18107), .A(n18106), .ZN(n20848) );
  AOI22_X1 U20268 ( .A1(n21167), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n18128), 
        .B2(n20848), .ZN(n18115) );
  NAND2_X1 U20269 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20160) );
  AOI21_X1 U20270 ( .B1(n18110), .B2(n20160), .A(n18109), .ZN(n20172) );
  OAI21_X1 U20271 ( .B1(n10977), .B2(n20157), .A(n18110), .ZN(n18112) );
  AOI22_X1 U20272 ( .A1(n20172), .A2(n18129), .B1(n18113), .B2(n18112), .ZN(
        n18114) );
  OAI211_X1 U20273 ( .C1(n18139), .C2(n20851), .A(n18115), .B(n18114), .ZN(
        P3_U2827) );
  AOI21_X1 U20274 ( .B1(n18118), .B2(n18117), .A(n18116), .ZN(n20838) );
  INV_X1 U20275 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n20156) );
  NOR2_X1 U20276 ( .A1(n21176), .A2(n20156), .ZN(n20839) );
  OAI21_X1 U20277 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n20160), .ZN(n20168) );
  OAI21_X1 U20278 ( .B1(n18121), .B2(n18120), .A(n18119), .ZN(n20835) );
  OAI22_X1 U20279 ( .A1(n18122), .A2(n20168), .B1(n18139), .B2(n20835), .ZN(
        n18123) );
  AOI211_X1 U20280 ( .C1(n18128), .C2(n20838), .A(n20839), .B(n18123), .ZN(
        n18124) );
  OAI221_X1 U20281 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n19005), .C1(
        n20157), .C2(n18136), .A(n18124), .ZN(P3_U2828) );
  OAI21_X1 U20282 ( .B1(n18126), .B2(n18133), .A(n18125), .ZN(n20823) );
  NAND2_X1 U20283 ( .A1(n20827), .A2(n18134), .ZN(n18127) );
  XNOR2_X1 U20284 ( .A(n18127), .B(n18126), .ZN(n20820) );
  AOI22_X1 U20285 ( .A1(n21167), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18128), 
        .B2(n20820), .ZN(n18132) );
  AOI22_X1 U20286 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n18130), .B1(
        n18129), .B2(n20150), .ZN(n18131) );
  OAI211_X1 U20287 ( .C1(n18139), .C2(n20823), .A(n18132), .B(n18131), .ZN(
        P3_U2829) );
  AOI21_X1 U20288 ( .B1(n18134), .B2(n20827), .A(n18133), .ZN(n20818) );
  INV_X1 U20289 ( .A(n20818), .ZN(n20817) );
  NAND3_X1 U20290 ( .A1(n20754), .A2(n18136), .A3(n18135), .ZN(n18137) );
  AOI22_X1 U20291 ( .A1(n21167), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18137), .ZN(n18138) );
  OAI221_X1 U20292 ( .B1(n20818), .B2(n18140), .C1(n20817), .C2(n18139), .A(
        n18138), .ZN(P3_U2830) );
  NOR2_X1 U20293 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18714), .ZN(
        n18742) );
  INV_X1 U20294 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n21213) );
  NOR2_X1 U20295 ( .A1(n21210), .A2(n21213), .ZN(n18725) );
  NAND2_X1 U20296 ( .A1(n21210), .A2(n21213), .ZN(n18776) );
  INV_X1 U20297 ( .A(n18776), .ZN(n18778) );
  NOR3_X1 U20298 ( .A1(n18725), .A2(n18778), .A3(n18771), .ZN(n18141) );
  AOI21_X1 U20299 ( .B1(n18742), .B2(n18142), .A(n18141), .ZN(n18144) );
  OAI22_X1 U20300 ( .A1(n18145), .A2(n18144), .B1(n18143), .B2(n21213), .ZN(
        P3_U2866) );
  NOR4_X1 U20301 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18149) );
  NOR4_X1 U20302 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n18148) );
  NOR4_X1 U20303 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18147) );
  NOR4_X1 U20304 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18146) );
  NAND4_X1 U20305 ( .A1(n18149), .A2(n18148), .A3(n18147), .A4(n18146), .ZN(
        n18155) );
  NOR4_X1 U20306 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_28__SCAN_IN), .A3(P3_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n18153) );
  AOI211_X1 U20307 ( .C1(P3_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A(P3_DATAWIDTH_REG_31__SCAN_IN), .B(
        P3_DATAWIDTH_REG_30__SCAN_IN), .ZN(n18152) );
  NOR4_X1 U20308 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18151) );
  NOR4_X1 U20309 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18150) );
  NAND4_X1 U20310 ( .A1(n18153), .A2(n18152), .A3(n18151), .A4(n18150), .ZN(
        n18154) );
  NOR2_X1 U20311 ( .A1(n18155), .A2(n18154), .ZN(n18166) );
  INV_X1 U20312 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18157) );
  OAI21_X1 U20313 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18166), .ZN(n18156) );
  OAI21_X1 U20314 ( .B1(n18166), .B2(n18157), .A(n18156), .ZN(P3_U3293) );
  INV_X1 U20315 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18160) );
  AOI21_X1 U20316 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18158) );
  INV_X1 U20317 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n20826) );
  OAI221_X1 U20318 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n18158), .C1(n20826), 
        .C2(P3_REIP_REG_0__SCAN_IN), .A(n18166), .ZN(n18159) );
  OAI21_X1 U20319 ( .B1(n18166), .B2(n18160), .A(n18159), .ZN(P3_U3292) );
  INV_X1 U20320 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18162) );
  NOR3_X1 U20321 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n18163) );
  OAI21_X1 U20322 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n18163), .A(n18166), .ZN(
        n18161) );
  OAI21_X1 U20323 ( .B1(n18166), .B2(n18162), .A(n18161), .ZN(P3_U2638) );
  INV_X1 U20324 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18165) );
  INV_X1 U20325 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21614) );
  OAI211_X1 U20326 ( .C1(n18163), .C2(n20826), .A(n21614), .B(n18166), .ZN(
        n18164) );
  OAI21_X1 U20327 ( .B1(n18166), .B2(n18165), .A(n18164), .ZN(P3_U2639) );
  INV_X1 U20328 ( .A(n18235), .ZN(n18228) );
  INV_X1 U20329 ( .A(P3_M_IO_N_REG_SCAN_IN), .ZN(n18237) );
  AOI22_X1 U20330 ( .A1(n18228), .A2(n18167), .B1(n18237), .B2(n18235), .ZN(
        P3_U3297) );
  OAI22_X1 U20331 ( .A1(n18235), .A2(n18168), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n21621), .ZN(n18169) );
  INV_X1 U20332 ( .A(n18169), .ZN(P3_U3294) );
  AOI21_X1 U20333 ( .B1(n21666), .B2(n21618), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n18170) );
  AOI22_X1 U20334 ( .A1(n18228), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n18170), 
        .B2(n18235), .ZN(P3_U2635) );
  INV_X1 U20335 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n20744) );
  AOI22_X1 U20336 ( .A1(n20098), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n18211), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n18171) );
  OAI21_X1 U20337 ( .B1(n20744), .B2(n18191), .A(n18171), .ZN(P3_U2767) );
  INV_X1 U20338 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n20591) );
  AOI22_X1 U20339 ( .A1(n20098), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n18211), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n18172) );
  OAI21_X1 U20340 ( .B1(n20591), .B2(n18191), .A(n18172), .ZN(P3_U2766) );
  INV_X1 U20341 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n20618) );
  AOI22_X1 U20342 ( .A1(n20098), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n18211), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n18173) );
  OAI21_X1 U20343 ( .B1(n20618), .B2(n18191), .A(n18173), .ZN(P3_U2765) );
  INV_X1 U20344 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n20614) );
  AOI22_X1 U20345 ( .A1(n20098), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n18203), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n18174) );
  OAI21_X1 U20346 ( .B1(n20614), .B2(n18191), .A(n18174), .ZN(P3_U2764) );
  INV_X1 U20347 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n18176) );
  AOI22_X1 U20348 ( .A1(n20098), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n18203), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n18175) );
  OAI21_X1 U20349 ( .B1(n18176), .B2(n18191), .A(n18175), .ZN(P3_U2763) );
  INV_X1 U20350 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n20564) );
  AOI22_X1 U20351 ( .A1(n20098), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n18203), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n18177) );
  OAI21_X1 U20352 ( .B1(n20564), .B2(n18191), .A(n18177), .ZN(P3_U2762) );
  INV_X1 U20353 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n20592) );
  AOI22_X1 U20354 ( .A1(n20098), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n18203), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n18178) );
  OAI21_X1 U20355 ( .B1(n20592), .B2(n18191), .A(n18178), .ZN(P3_U2761) );
  INV_X1 U20356 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n18180) );
  AOI22_X1 U20357 ( .A1(n20098), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n18211), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n18179) );
  OAI21_X1 U20358 ( .B1(n18180), .B2(n18191), .A(n18179), .ZN(P3_U2760) );
  INV_X1 U20359 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n20132) );
  AOI22_X1 U20360 ( .A1(n20098), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n18211), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n18181) );
  OAI21_X1 U20361 ( .B1(n20132), .B2(n18191), .A(n18181), .ZN(P3_U2759) );
  INV_X1 U20362 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n20584) );
  AOI22_X1 U20363 ( .A1(n20098), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n18211), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n18182) );
  OAI21_X1 U20364 ( .B1(n20584), .B2(n18191), .A(n18182), .ZN(P3_U2758) );
  INV_X1 U20365 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n18184) );
  AOI22_X1 U20366 ( .A1(n20098), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n18211), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n18183) );
  OAI21_X1 U20367 ( .B1(n18184), .B2(n18191), .A(n18183), .ZN(P3_U2757) );
  INV_X1 U20368 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n20620) );
  AOI22_X1 U20369 ( .A1(n20098), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n18211), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n18185) );
  OAI21_X1 U20370 ( .B1(n20620), .B2(n18191), .A(n18185), .ZN(P3_U2756) );
  INV_X1 U20371 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n20567) );
  AOI22_X1 U20372 ( .A1(n20098), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n18211), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n18186) );
  OAI21_X1 U20373 ( .B1(n20567), .B2(n18191), .A(n18186), .ZN(P3_U2755) );
  INV_X1 U20374 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n18188) );
  AOI22_X1 U20375 ( .A1(n20098), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n18211), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n18187) );
  OAI21_X1 U20376 ( .B1(n18188), .B2(n18191), .A(n18187), .ZN(P3_U2754) );
  INV_X1 U20377 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n20719) );
  AOI22_X1 U20378 ( .A1(n20098), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n18211), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n18189) );
  OAI21_X1 U20379 ( .B1(n20719), .B2(n18191), .A(n18189), .ZN(P3_U2753) );
  INV_X1 U20380 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n20726) );
  AOI22_X1 U20381 ( .A1(n20098), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n18211), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n18190) );
  OAI21_X1 U20382 ( .B1(n20726), .B2(n18191), .A(n18190), .ZN(P3_U2752) );
  INV_X1 U20383 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n18194) );
  NAND2_X1 U20384 ( .A1(n18192), .A2(n11096), .ZN(n18213) );
  AOI22_X1 U20385 ( .A1(n20098), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n18211), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n18193) );
  OAI21_X1 U20386 ( .B1(n18194), .B2(n18213), .A(n18193), .ZN(P3_U2751) );
  INV_X1 U20387 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n20623) );
  AOI22_X1 U20388 ( .A1(n20098), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n18211), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n18195) );
  OAI21_X1 U20389 ( .B1(n20623), .B2(n18213), .A(n18195), .ZN(P3_U2750) );
  INV_X1 U20390 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n20647) );
  AOI22_X1 U20391 ( .A1(n20098), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n18211), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n18196) );
  OAI21_X1 U20392 ( .B1(n20647), .B2(n18213), .A(n18196), .ZN(P3_U2749) );
  INV_X1 U20393 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n20109) );
  AOI22_X1 U20394 ( .A1(n20098), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n18203), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n18197) );
  OAI21_X1 U20395 ( .B1(n20109), .B2(n18213), .A(n18197), .ZN(P3_U2748) );
  INV_X1 U20396 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n20660) );
  AOI22_X1 U20397 ( .A1(n20098), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n18203), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n18198) );
  OAI21_X1 U20398 ( .B1(n20660), .B2(n18213), .A(n18198), .ZN(P3_U2747) );
  INV_X1 U20399 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n20638) );
  AOI22_X1 U20400 ( .A1(n20098), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n18203), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n18199) );
  OAI21_X1 U20401 ( .B1(n20638), .B2(n18213), .A(n18199), .ZN(P3_U2746) );
  INV_X1 U20402 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n20659) );
  AOI22_X1 U20403 ( .A1(n20098), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n18203), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n18200) );
  OAI21_X1 U20404 ( .B1(n20659), .B2(n18213), .A(n18200), .ZN(P3_U2745) );
  INV_X1 U20405 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n18202) );
  AOI22_X1 U20406 ( .A1(n20098), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n18203), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n18201) );
  OAI21_X1 U20407 ( .B1(n18202), .B2(n18213), .A(n18201), .ZN(P3_U2744) );
  AOI22_X1 U20408 ( .A1(n20098), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n18203), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n18204) );
  OAI21_X1 U20409 ( .B1(n11089), .B2(n18213), .A(n18204), .ZN(P3_U2743) );
  INV_X1 U20410 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n20662) );
  AOI22_X1 U20411 ( .A1(n20098), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n18211), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n18205) );
  OAI21_X1 U20412 ( .B1(n20662), .B2(n18213), .A(n18205), .ZN(P3_U2742) );
  AOI22_X1 U20413 ( .A1(n20098), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n18211), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n18206) );
  OAI21_X1 U20414 ( .B1(n11090), .B2(n18213), .A(n18206), .ZN(P3_U2741) );
  INV_X1 U20415 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n20689) );
  AOI22_X1 U20416 ( .A1(n20098), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n18211), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n18207) );
  OAI21_X1 U20417 ( .B1(n20689), .B2(n18213), .A(n18207), .ZN(P3_U2740) );
  INV_X1 U20418 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n18209) );
  AOI22_X1 U20419 ( .A1(n20098), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n18211), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n18208) );
  OAI21_X1 U20420 ( .B1(n18209), .B2(n18213), .A(n18208), .ZN(P3_U2739) );
  INV_X1 U20421 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n20677) );
  AOI22_X1 U20422 ( .A1(n20098), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n18211), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n18210) );
  OAI21_X1 U20423 ( .B1(n20677), .B2(n18213), .A(n18210), .ZN(P3_U2738) );
  INV_X1 U20424 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n20121) );
  AOI22_X1 U20425 ( .A1(n20098), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n18211), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n18212) );
  OAI21_X1 U20426 ( .B1(n20121), .B2(n18213), .A(n18212), .ZN(P3_U2737) );
  NOR2_X1 U20427 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(n18214), .ZN(n18215) );
  NOR2_X1 U20428 ( .A1(n21621), .A2(n18215), .ZN(P3_U2633) );
  NOR2_X1 U20429 ( .A1(n18235), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n21660) );
  INV_X1 U20430 ( .A(n21660), .ZN(n18229) );
  CLKBUF_X1 U20431 ( .A(n18229), .Z(n18226) );
  AOI22_X1 U20432 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n18230), .B1(
        P3_ADDRESS_REG_0__SCAN_IN), .B2(n18235), .ZN(n18216) );
  OAI21_X1 U20433 ( .B1(n20156), .B2(n18226), .A(n18216), .ZN(P3_U3032) );
  INV_X1 U20434 ( .A(n18230), .ZN(n18227) );
  AOI22_X1 U20435 ( .A1(n21660), .A2(P3_REIP_REG_3__SCAN_IN), .B1(
        P3_ADDRESS_REG_1__SCAN_IN), .B2(n18235), .ZN(n18217) );
  OAI21_X1 U20436 ( .B1(n18227), .B2(n20156), .A(n18217), .ZN(P3_U3033) );
  AOI22_X1 U20437 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n18230), .B1(
        P3_ADDRESS_REG_2__SCAN_IN), .B2(n18235), .ZN(n18218) );
  OAI21_X1 U20438 ( .B1(n20186), .B2(n18226), .A(n18218), .ZN(P3_U3034) );
  AOI22_X1 U20439 ( .A1(n21660), .A2(P3_REIP_REG_5__SCAN_IN), .B1(
        P3_ADDRESS_REG_3__SCAN_IN), .B2(n18235), .ZN(n18219) );
  OAI21_X1 U20440 ( .B1(n18227), .B2(n20186), .A(n18219), .ZN(P3_U3035) );
  AOI22_X1 U20441 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n18230), .B1(
        P3_ADDRESS_REG_4__SCAN_IN), .B2(n18235), .ZN(n18220) );
  OAI21_X1 U20442 ( .B1(n20875), .B2(n18226), .A(n18220), .ZN(P3_U3036) );
  INV_X1 U20443 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n19807) );
  OAI222_X1 U20444 ( .A1(n18226), .A2(n20225), .B1(n19807), .B2(n18228), .C1(
        n20875), .C2(n18227), .ZN(P3_U3037) );
  INV_X1 U20445 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n19809) );
  OAI222_X1 U20446 ( .A1(n18229), .A2(n20239), .B1(n19809), .B2(n18228), .C1(
        n20225), .C2(n18227), .ZN(P3_U3038) );
  INV_X1 U20447 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n19811) );
  OAI222_X1 U20448 ( .A1(n18229), .A2(n18221), .B1(n19811), .B2(n18228), .C1(
        n20239), .C2(n18227), .ZN(P3_U3039) );
  INV_X1 U20449 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n19813) );
  OAI222_X1 U20450 ( .A1(n18226), .A2(n20263), .B1(n19813), .B2(n18228), .C1(
        n18221), .C2(n18227), .ZN(P3_U3040) );
  INV_X1 U20451 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n19815) );
  OAI222_X1 U20452 ( .A1(n20263), .A2(n18227), .B1(n19815), .B2(n18228), .C1(
        n20920), .C2(n18226), .ZN(P3_U3041) );
  INV_X1 U20453 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n20299) );
  INV_X1 U20454 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n19817) );
  OAI222_X1 U20455 ( .A1(n18226), .A2(n20299), .B1(n19817), .B2(n18228), .C1(
        n20920), .C2(n18227), .ZN(P3_U3042) );
  INV_X1 U20456 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n19819) );
  OAI222_X1 U20457 ( .A1(n18226), .A2(n20344), .B1(n19819), .B2(n18228), .C1(
        n20299), .C2(n18227), .ZN(P3_U3043) );
  INV_X1 U20458 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n19821) );
  OAI222_X1 U20459 ( .A1(n20344), .A2(n18227), .B1(n19821), .B2(n18228), .C1(
        n20343), .C2(n18226), .ZN(P3_U3044) );
  INV_X1 U20460 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n20346) );
  INV_X1 U20461 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n19823) );
  OAI222_X1 U20462 ( .A1(n18226), .A2(n20346), .B1(n19823), .B2(n18228), .C1(
        n20343), .C2(n18227), .ZN(P3_U3045) );
  INV_X1 U20463 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n19825) );
  OAI222_X1 U20464 ( .A1(n18226), .A2(n20365), .B1(n19825), .B2(n18228), .C1(
        n20346), .C2(n18227), .ZN(P3_U3046) );
  INV_X1 U20465 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n19827) );
  OAI222_X1 U20466 ( .A1(n18226), .A2(n20366), .B1(n19827), .B2(n18228), .C1(
        n20365), .C2(n18227), .ZN(P3_U3047) );
  INV_X1 U20467 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n19829) );
  OAI222_X1 U20468 ( .A1(n18229), .A2(n21126), .B1(n19829), .B2(n18228), .C1(
        n20366), .C2(n18227), .ZN(P3_U3048) );
  INV_X1 U20469 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n19831) );
  OAI222_X1 U20470 ( .A1(n18229), .A2(n18223), .B1(n19831), .B2(n18228), .C1(
        n21126), .C2(n18227), .ZN(P3_U3049) );
  AOI22_X1 U20471 ( .A1(n21660), .A2(P3_REIP_REG_20__SCAN_IN), .B1(
        P3_ADDRESS_REG_18__SCAN_IN), .B2(n18235), .ZN(n18222) );
  OAI21_X1 U20472 ( .B1(n18227), .B2(n18223), .A(n18222), .ZN(P3_U3050) );
  AOI22_X1 U20473 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n18230), .B1(
        P3_ADDRESS_REG_19__SCAN_IN), .B2(n18235), .ZN(n18224) );
  OAI21_X1 U20474 ( .B1(n20425), .B2(n18226), .A(n18224), .ZN(P3_U3051) );
  INV_X1 U20475 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n20430) );
  INV_X1 U20476 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n19835) );
  OAI222_X1 U20477 ( .A1(n18229), .A2(n20430), .B1(n19835), .B2(n18228), .C1(
        n20425), .C2(n18227), .ZN(P3_U3052) );
  INV_X1 U20478 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18225) );
  INV_X1 U20479 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n19837) );
  OAI222_X1 U20480 ( .A1(n18229), .A2(n18225), .B1(n19837), .B2(n18228), .C1(
        n20430), .C2(n18227), .ZN(P3_U3053) );
  INV_X1 U20481 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n19839) );
  OAI222_X1 U20482 ( .A1(n18226), .A2(n20465), .B1(n19839), .B2(n18228), .C1(
        n18225), .C2(n18227), .ZN(P3_U3054) );
  INV_X1 U20483 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n19841) );
  OAI222_X1 U20484 ( .A1(n18226), .A2(n20471), .B1(n19841), .B2(n18228), .C1(
        n20465), .C2(n18227), .ZN(P3_U3055) );
  INV_X1 U20485 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n19843) );
  OAI222_X1 U20486 ( .A1(n18229), .A2(n20493), .B1(n19843), .B2(n18228), .C1(
        n20471), .C2(n18227), .ZN(P3_U3056) );
  INV_X1 U20487 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n20506) );
  INV_X1 U20488 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n19845) );
  OAI222_X1 U20489 ( .A1(n18226), .A2(n20506), .B1(n19845), .B2(n18228), .C1(
        n20493), .C2(n18227), .ZN(P3_U3057) );
  INV_X1 U20490 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n19847) );
  OAI222_X1 U20491 ( .A1(n18226), .A2(n20519), .B1(n19847), .B2(n18228), .C1(
        n20506), .C2(n18227), .ZN(P3_U3058) );
  INV_X1 U20492 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n19849) );
  OAI222_X1 U20493 ( .A1(n20519), .A2(n18227), .B1(n19849), .B2(n18228), .C1(
        n20528), .C2(n18226), .ZN(P3_U3059) );
  INV_X1 U20494 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n19851) );
  OAI222_X1 U20495 ( .A1(n18229), .A2(n21037), .B1(n19851), .B2(n18228), .C1(
        n20528), .C2(n18227), .ZN(P3_U3060) );
  AOI222_X1 U20496 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n18230), .B1(
        P3_ADDRESS_REG_29__SCAN_IN), .B2(n18235), .C1(P3_REIP_REG_31__SCAN_IN), 
        .C2(n21660), .ZN(n18231) );
  INV_X1 U20497 ( .A(n18231), .ZN(P3_U3061) );
  OAI22_X1 U20498 ( .A1(n18235), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n21621), .ZN(n18232) );
  INV_X1 U20499 ( .A(n18232), .ZN(P3_U3277) );
  OAI22_X1 U20500 ( .A1(n18235), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n21621), .ZN(n18233) );
  INV_X1 U20501 ( .A(n18233), .ZN(P3_U3276) );
  OAI22_X1 U20502 ( .A1(n18235), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n21621), .ZN(n18234) );
  INV_X1 U20503 ( .A(n18234), .ZN(P3_U3275) );
  OAI22_X1 U20504 ( .A1(n18235), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n21621), .ZN(n18236) );
  INV_X1 U20505 ( .A(n18236), .ZN(P3_U3274) );
  NOR4_X1 U20506 ( .A1(P3_BE_N_REG_1__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_BE_N_REG_2__SCAN_IN), .A4(P3_BE_N_REG_0__SCAN_IN), .ZN(n18239)
         );
  NOR4_X1 U20507 ( .A1(P3_ADS_N_REG_SCAN_IN), .A2(P3_D_C_N_REG_SCAN_IN), .A3(
        P3_W_R_N_REG_SCAN_IN), .A4(n18237), .ZN(n18238) );
  NAND3_X1 U20508 ( .A1(n18239), .A2(n18238), .A3(U215), .ZN(U213) );
  NOR2_X1 U20509 ( .A1(n21639), .A2(n18247), .ZN(n18245) );
  INV_X1 U20510 ( .A(n21645), .ZN(n18241) );
  OAI21_X1 U20511 ( .B1(n18241), .B2(n21607), .A(n18240), .ZN(n18243) );
  NAND3_X1 U20512 ( .A1(n18241), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n19686), 
        .ZN(n18242) );
  MUX2_X1 U20513 ( .A(n18243), .B(n18242), .S(n11774), .Z(n18244) );
  OAI21_X1 U20514 ( .B1(n18245), .B2(n18667), .A(n18244), .ZN(n18252) );
  NOR3_X1 U20515 ( .A1(n21639), .A2(n18247), .A3(n18246), .ZN(n18249) );
  AOI211_X1 U20516 ( .C1(n18250), .C2(n18657), .A(n18249), .B(n18248), .ZN(
        n18251) );
  MUX2_X1 U20517 ( .A(n18252), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n18251), 
        .Z(P2_U3610) );
  AOI22_X1 U20518 ( .A1(n18254), .A2(n18539), .B1(n18538), .B2(
        P2_EBX_REG_0__SCAN_IN), .ZN(n18257) );
  AOI22_X1 U20519 ( .A1(n18536), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n18534), 
        .B2(n18255), .ZN(n18256) );
  OAI211_X1 U20520 ( .C1(n18258), .C2(n18447), .A(n18257), .B(n18256), .ZN(
        n18259) );
  AOI21_X1 U20521 ( .B1(n18260), .B2(n18269), .A(n18259), .ZN(n18262) );
  NAND2_X1 U20522 ( .A1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18537), .ZN(
        n18261) );
  OAI211_X1 U20523 ( .C1(n13795), .C2(n18663), .A(n18262), .B(n18261), .ZN(
        P2_U2855) );
  INV_X1 U20524 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n18263) );
  OAI21_X1 U20525 ( .B1(n18263), .B2(n18554), .A(n18582), .ZN(n18265) );
  OAI22_X1 U20526 ( .A1(n18567), .A2(n19454), .B1(n12132), .B2(n18551), .ZN(
        n18264) );
  AOI211_X1 U20527 ( .C1(P2_EBX_REG_4__SCAN_IN), .C2(n18538), .A(n18265), .B(
        n18264), .ZN(n18266) );
  OAI21_X1 U20528 ( .B1(n18267), .B2(n18552), .A(n18266), .ZN(n18268) );
  AOI21_X1 U20529 ( .B1(n19393), .B2(n18269), .A(n18268), .ZN(n18276) );
  INV_X1 U20530 ( .A(n18270), .ZN(n18274) );
  NOR2_X1 U20531 ( .A1(n18361), .A2(n18271), .ZN(n18273) );
  AOI21_X1 U20532 ( .B1(n18274), .B2(n18273), .A(n18663), .ZN(n18272) );
  OAI21_X1 U20533 ( .B1(n18274), .B2(n18273), .A(n18272), .ZN(n18275) );
  OAI211_X1 U20534 ( .C1(n18277), .C2(n18447), .A(n18276), .B(n18275), .ZN(
        P2_U2851) );
  OAI21_X1 U20535 ( .B1(n12135), .B2(n18551), .A(n18583), .ZN(n18281) );
  OAI22_X1 U20536 ( .A1(n18279), .A2(n18552), .B1(n18278), .B2(n18557), .ZN(
        n18280) );
  AOI211_X1 U20537 ( .C1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n18537), .A(
        n18281), .B(n18280), .ZN(n18288) );
  NAND2_X1 U20538 ( .A1(n18562), .A2(n18282), .ZN(n18283) );
  XNOR2_X1 U20539 ( .A(n18284), .B(n18283), .ZN(n18285) );
  AOI22_X1 U20540 ( .A1(n18560), .A2(n18286), .B1(n18564), .B2(n18285), .ZN(
        n18287) );
  OAI211_X1 U20541 ( .C1(n18567), .C2(n19394), .A(n18288), .B(n18287), .ZN(
        P2_U2850) );
  OAI21_X1 U20542 ( .B1(n12138), .B2(n18551), .A(n18583), .ZN(n18292) );
  INV_X1 U20543 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n18289) );
  OAI22_X1 U20544 ( .A1(n18290), .A2(n18552), .B1(n18289), .B2(n18557), .ZN(
        n18291) );
  AOI211_X1 U20545 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n18524), .A(
        n18292), .B(n18291), .ZN(n18299) );
  NOR2_X1 U20546 ( .A1(n18361), .A2(n18293), .ZN(n18295) );
  XNOR2_X1 U20547 ( .A(n18295), .B(n18294), .ZN(n18296) );
  AOI22_X1 U20548 ( .A1(n18560), .A2(n18297), .B1(n18564), .B2(n18296), .ZN(
        n18298) );
  OAI211_X1 U20549 ( .C1(n18567), .C2(n19350), .A(n18299), .B(n18298), .ZN(
        P2_U2849) );
  NAND2_X1 U20550 ( .A1(n18562), .A2(n18300), .ZN(n18302) );
  XOR2_X1 U20551 ( .A(n18302), .B(n18301), .Z(n18311) );
  INV_X1 U20552 ( .A(n18303), .ZN(n18309) );
  AOI22_X1 U20553 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n18524), .B1(
        n18304), .B2(n18534), .ZN(n18305) );
  OAI211_X1 U20554 ( .C1(n18557), .C2(n14966), .A(n18305), .B(n18583), .ZN(
        n18306) );
  AOI21_X1 U20555 ( .B1(n18536), .B2(P2_REIP_REG_7__SCAN_IN), .A(n18306), .ZN(
        n18307) );
  OAI21_X1 U20556 ( .B1(n19185), .B2(n18567), .A(n18307), .ZN(n18308) );
  AOI21_X1 U20557 ( .B1(n18309), .B2(n18560), .A(n18308), .ZN(n18310) );
  OAI21_X1 U20558 ( .B1(n18311), .B2(n18663), .A(n18310), .ZN(P2_U2848) );
  AOI22_X1 U20559 ( .A1(n18538), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18537), .ZN(n18312) );
  OAI21_X1 U20560 ( .B1(n18313), .B2(n18552), .A(n18312), .ZN(n18314) );
  AOI211_X1 U20561 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n18536), .A(n18382), .B(
        n18314), .ZN(n18320) );
  NOR2_X1 U20562 ( .A1(n18361), .A2(n18315), .ZN(n18317) );
  XNOR2_X1 U20563 ( .A(n18317), .B(n18316), .ZN(n18318) );
  AOI22_X1 U20564 ( .A1(n18539), .A2(n19180), .B1(n18564), .B2(n18318), .ZN(
        n18319) );
  OAI211_X1 U20565 ( .C1(n18447), .C2(n18321), .A(n18320), .B(n18319), .ZN(
        P2_U2847) );
  AOI22_X1 U20566 ( .A1(n18322), .A2(n18534), .B1(P2_EBX_REG_9__SCAN_IN), .B2(
        n18538), .ZN(n18323) );
  OAI211_X1 U20567 ( .C1(n12157), .C2(n18551), .A(n18323), .B(n18582), .ZN(
        n18324) );
  AOI21_X1 U20568 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18524), .A(
        n18324), .ZN(n18330) );
  NAND2_X1 U20569 ( .A1(n18562), .A2(n18325), .ZN(n18326) );
  XNOR2_X1 U20570 ( .A(n18327), .B(n18326), .ZN(n18328) );
  AOI22_X1 U20571 ( .A1(n18539), .A2(n19177), .B1(n18564), .B2(n18328), .ZN(
        n18329) );
  OAI211_X1 U20572 ( .C1(n18447), .C2(n18331), .A(n18330), .B(n18329), .ZN(
        P2_U2846) );
  NOR2_X1 U20573 ( .A1(n18361), .A2(n18332), .ZN(n18333) );
  XOR2_X1 U20574 ( .A(n18334), .B(n18333), .Z(n18343) );
  INV_X1 U20575 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n18337) );
  AOI22_X1 U20576 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n18524), .B1(
        n18335), .B2(n18534), .ZN(n18336) );
  OAI211_X1 U20577 ( .C1(n18557), .C2(n18337), .A(n18336), .B(n18583), .ZN(
        n18338) );
  AOI21_X1 U20578 ( .B1(n18536), .B2(P2_REIP_REG_10__SCAN_IN), .A(n18338), 
        .ZN(n18339) );
  OAI21_X1 U20579 ( .B1(n19174), .B2(n18567), .A(n18339), .ZN(n18340) );
  AOI21_X1 U20580 ( .B1(n18341), .B2(n18560), .A(n18340), .ZN(n18342) );
  OAI21_X1 U20581 ( .B1(n18663), .B2(n18343), .A(n18342), .ZN(P2_U2845) );
  OAI21_X1 U20582 ( .B1(n12163), .B2(n18551), .A(n18583), .ZN(n18347) );
  INV_X1 U20583 ( .A(n18344), .ZN(n18345) );
  OAI22_X1 U20584 ( .A1(n18345), .A2(n18552), .B1(n11576), .B2(n18557), .ZN(
        n18346) );
  AOI211_X1 U20585 ( .C1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .C2(n18537), .A(
        n18347), .B(n18346), .ZN(n18354) );
  NAND2_X1 U20586 ( .A1(n18562), .A2(n18348), .ZN(n18349) );
  XNOR2_X1 U20587 ( .A(n18350), .B(n18349), .ZN(n18351) );
  AOI22_X1 U20588 ( .A1(n18560), .A2(n18352), .B1(n18564), .B2(n18351), .ZN(
        n18353) );
  OAI211_X1 U20589 ( .C1(n18567), .C2(n19171), .A(n18354), .B(n18353), .ZN(
        P2_U2844) );
  AOI22_X1 U20590 ( .A1(n18538), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18537), .ZN(n18355) );
  OAI21_X1 U20591 ( .B1(n18356), .B2(n18552), .A(n18355), .ZN(n18357) );
  AOI211_X1 U20592 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n18536), .A(n18382), 
        .B(n18357), .ZN(n18366) );
  AOI21_X1 U20593 ( .B1(n18359), .B2(n16777), .A(n18358), .ZN(n19166) );
  NOR2_X1 U20594 ( .A1(n18361), .A2(n18360), .ZN(n18363) );
  XNOR2_X1 U20595 ( .A(n18363), .B(n18362), .ZN(n18364) );
  AOI22_X1 U20596 ( .A1(n18539), .A2(n19166), .B1(n18564), .B2(n18364), .ZN(
        n18365) );
  OAI211_X1 U20597 ( .C1(n18447), .C2(n18367), .A(n18366), .B(n18365), .ZN(
        P2_U2843) );
  AOI22_X1 U20598 ( .A1(n18538), .A2(P2_EBX_REG_14__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n18537), .ZN(n18368) );
  OAI21_X1 U20599 ( .B1(n18369), .B2(n18552), .A(n18368), .ZN(n18370) );
  AOI211_X1 U20600 ( .C1(P2_REIP_REG_14__SCAN_IN), .C2(n18536), .A(n18382), 
        .B(n18370), .ZN(n18379) );
  NAND2_X1 U20601 ( .A1(n18372), .A2(n18371), .ZN(n18373) );
  AOI22_X1 U20602 ( .A1(n18539), .A2(n19159), .B1(n18560), .B2(n18577), .ZN(
        n18378) );
  OAI211_X1 U20603 ( .C1(n18376), .C2(n18375), .A(n18564), .B(n18374), .ZN(
        n18377) );
  NAND3_X1 U20604 ( .A1(n18379), .A2(n18378), .A3(n18377), .ZN(P2_U2841) );
  OAI22_X1 U20605 ( .A1(n18380), .A2(n18552), .B1(n11580), .B2(n18557), .ZN(
        n18381) );
  AOI211_X1 U20606 ( .C1(P2_REIP_REG_15__SCAN_IN), .C2(n18536), .A(n18382), 
        .B(n18381), .ZN(n18387) );
  OAI211_X1 U20607 ( .C1(n18385), .C2(n18384), .A(n18564), .B(n18383), .ZN(
        n18386) );
  OAI211_X1 U20608 ( .C1(n18554), .C2(n11151), .A(n18387), .B(n18386), .ZN(
        n18388) );
  AOI21_X1 U20609 ( .B1(n18560), .B2(n18389), .A(n18388), .ZN(n18390) );
  OAI21_X1 U20610 ( .B1(n18567), .B2(n19157), .A(n18390), .ZN(P2_U2840) );
  INV_X1 U20611 ( .A(n19675), .ZN(n18396) );
  AOI21_X1 U20612 ( .B1(P2_REIP_REG_16__SCAN_IN), .B2(n18536), .A(n18382), 
        .ZN(n18393) );
  AOI22_X1 U20613 ( .A1(n18391), .A2(n18534), .B1(P2_EBX_REG_16__SCAN_IN), 
        .B2(n18538), .ZN(n18392) );
  OAI211_X1 U20614 ( .C1(n18394), .C2(n18554), .A(n18393), .B(n18392), .ZN(
        n18395) );
  AOI21_X1 U20615 ( .B1(n18539), .B2(n18396), .A(n18395), .ZN(n18401) );
  OAI211_X1 U20616 ( .C1(n18399), .C2(n18398), .A(n18564), .B(n18397), .ZN(
        n18400) );
  OAI211_X1 U20617 ( .C1(n18402), .C2(n18447), .A(n18401), .B(n18400), .ZN(
        P2_U2839) );
  AOI22_X1 U20618 ( .A1(n18403), .A2(n18534), .B1(P2_EBX_REG_17__SCAN_IN), 
        .B2(n18538), .ZN(n18404) );
  OAI211_X1 U20619 ( .C1(n18405), .C2(n18551), .A(n18404), .B(n18582), .ZN(
        n18409) );
  OAI22_X1 U20620 ( .A1(n18567), .A2(n18407), .B1(n18447), .B2(n18406), .ZN(
        n18408) );
  AOI211_X1 U20621 ( .C1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(n18524), .A(
        n18409), .B(n18408), .ZN(n18414) );
  OAI211_X1 U20622 ( .C1(n18412), .C2(n18411), .A(n18564), .B(n18410), .ZN(
        n18413) );
  NAND2_X1 U20623 ( .A1(n18414), .A2(n18413), .ZN(P2_U2838) );
  AOI22_X1 U20624 ( .A1(n18415), .A2(n18534), .B1(P2_EBX_REG_18__SCAN_IN), 
        .B2(n18538), .ZN(n18416) );
  OAI211_X1 U20625 ( .C1(n18417), .C2(n18551), .A(n18416), .B(n18582), .ZN(
        n18421) );
  OAI22_X1 U20626 ( .A1(n18567), .A2(n18419), .B1(n18447), .B2(n18418), .ZN(
        n18420) );
  AOI211_X1 U20627 ( .C1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n18537), .A(
        n18421), .B(n18420), .ZN(n18426) );
  OAI211_X1 U20628 ( .C1(n18424), .C2(n18423), .A(n18564), .B(n18422), .ZN(
        n18425) );
  NAND2_X1 U20629 ( .A1(n18426), .A2(n18425), .ZN(P2_U2837) );
  AOI22_X1 U20630 ( .A1(n11964), .A2(n18534), .B1(P2_EBX_REG_19__SCAN_IN), 
        .B2(n18538), .ZN(n18427) );
  OAI211_X1 U20631 ( .C1(n16483), .C2(n18551), .A(n18427), .B(n18582), .ZN(
        n18428) );
  AOI21_X1 U20632 ( .B1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n18524), .A(
        n18428), .ZN(n18435) );
  INV_X1 U20633 ( .A(n18429), .ZN(n18602) );
  AOI22_X1 U20634 ( .A1(n18539), .A2(n18600), .B1(n18560), .B2(n18602), .ZN(
        n18434) );
  OAI211_X1 U20635 ( .C1(n18432), .C2(n18431), .A(n18564), .B(n18430), .ZN(
        n18433) );
  NAND3_X1 U20636 ( .A1(n18435), .A2(n18434), .A3(n18433), .ZN(P2_U2836) );
  INV_X1 U20637 ( .A(n19440), .ZN(n18441) );
  OAI22_X1 U20638 ( .A1(n11148), .A2(n18554), .B1(n18436), .B2(n18552), .ZN(
        n18440) );
  OAI22_X1 U20639 ( .A1(n18557), .A2(n18438), .B1(n18437), .B2(n18551), .ZN(
        n18439) );
  AOI211_X1 U20640 ( .C1(n18539), .C2(n18441), .A(n18440), .B(n18439), .ZN(
        n18446) );
  OAI211_X1 U20641 ( .C1(n18444), .C2(n18443), .A(n18564), .B(n18442), .ZN(
        n18445) );
  OAI211_X1 U20642 ( .C1(n18448), .C2(n18447), .A(n18446), .B(n18445), .ZN(
        P2_U2835) );
  AOI22_X1 U20643 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n18524), .B1(
        P2_REIP_REG_21__SCAN_IN), .B2(n18536), .ZN(n18457) );
  AOI22_X1 U20644 ( .A1(n11962), .A2(n18534), .B1(P2_EBX_REG_21__SCAN_IN), 
        .B2(n18538), .ZN(n18456) );
  AOI22_X1 U20645 ( .A1(n18450), .A2(n18560), .B1(n18449), .B2(n18539), .ZN(
        n18455) );
  OAI211_X1 U20646 ( .C1(n18453), .C2(n18452), .A(n18564), .B(n18451), .ZN(
        n18454) );
  NAND4_X1 U20647 ( .A1(n18457), .A2(n18456), .A3(n18455), .A4(n18454), .ZN(
        P2_U2834) );
  AOI22_X1 U20648 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18537), .B1(
        n18458), .B2(n18534), .ZN(n18466) );
  AOI22_X1 U20649 ( .A1(n18536), .A2(P2_REIP_REG_22__SCAN_IN), .B1(n18538), 
        .B2(P2_EBX_REG_22__SCAN_IN), .ZN(n18465) );
  AOI22_X1 U20650 ( .A1(n18539), .A2(n19343), .B1(n18560), .B2(n18459), .ZN(
        n18464) );
  OAI211_X1 U20651 ( .C1(n18462), .C2(n18461), .A(n18564), .B(n18460), .ZN(
        n18463) );
  NAND4_X1 U20652 ( .A1(n18466), .A2(n18465), .A3(n18464), .A4(n18463), .ZN(
        P2_U2833) );
  OAI22_X1 U20653 ( .A1(n16423), .A2(n18551), .B1(n18467), .B2(n18552), .ZN(
        n18471) );
  INV_X1 U20654 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n18468) );
  OAI22_X1 U20655 ( .A1(n18557), .A2(n18469), .B1(n18468), .B2(n18554), .ZN(
        n18470) );
  AOI211_X1 U20656 ( .C1(n18560), .C2(n18472), .A(n18471), .B(n18470), .ZN(
        n18477) );
  OAI211_X1 U20657 ( .C1(n18475), .C2(n18474), .A(n18564), .B(n18473), .ZN(
        n18476) );
  OAI211_X1 U20658 ( .C1(n18478), .C2(n18567), .A(n18477), .B(n18476), .ZN(
        P2_U2832) );
  AOI22_X1 U20659 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n18536), .B1(n18479), 
        .B2(n18534), .ZN(n18488) );
  AOI22_X1 U20660 ( .A1(n18538), .A2(P2_EBX_REG_24__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n18524), .ZN(n18487) );
  INV_X1 U20661 ( .A(n18480), .ZN(n18481) );
  AOI22_X1 U20662 ( .A1(n18539), .A2(n11367), .B1(n18560), .B2(n18481), .ZN(
        n18486) );
  OAI211_X1 U20663 ( .C1(n18484), .C2(n18483), .A(n18564), .B(n18482), .ZN(
        n18485) );
  NAND4_X1 U20664 ( .A1(n18488), .A2(n18487), .A3(n18486), .A4(n18485), .ZN(
        P2_U2831) );
  AOI22_X1 U20665 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n18536), .B1(n18489), 
        .B2(n18534), .ZN(n18498) );
  AOI22_X1 U20666 ( .A1(n18538), .A2(P2_EBX_REG_25__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18524), .ZN(n18497) );
  AOI22_X1 U20667 ( .A1(n18539), .A2(n18491), .B1(n18560), .B2(n18490), .ZN(
        n18496) );
  OAI211_X1 U20668 ( .C1(n18494), .C2(n18493), .A(n18564), .B(n18492), .ZN(
        n18495) );
  NAND4_X1 U20669 ( .A1(n18498), .A2(n18497), .A3(n18496), .A4(n18495), .ZN(
        P2_U2830) );
  AOI22_X1 U20670 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n18536), .B1(n18499), 
        .B2(n18534), .ZN(n18509) );
  AOI22_X1 U20671 ( .A1(n18538), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18537), .ZN(n18508) );
  INV_X1 U20672 ( .A(n18500), .ZN(n18502) );
  AOI22_X1 U20673 ( .A1(n18502), .A2(n18560), .B1(n18501), .B2(n18539), .ZN(
        n18507) );
  OAI211_X1 U20674 ( .C1(n18505), .C2(n18504), .A(n18564), .B(n18503), .ZN(
        n18506) );
  NAND4_X1 U20675 ( .A1(n18509), .A2(n18508), .A3(n18507), .A4(n18506), .ZN(
        P2_U2829) );
  OAI22_X1 U20676 ( .A1(n18511), .A2(n18551), .B1(n18510), .B2(n18552), .ZN(
        n18515) );
  OAI22_X1 U20677 ( .A1(n18557), .A2(n18513), .B1(n18512), .B2(n18554), .ZN(
        n18514) );
  AOI211_X1 U20678 ( .C1(n18516), .C2(n18560), .A(n18515), .B(n18514), .ZN(
        n18521) );
  OAI211_X1 U20679 ( .C1(n18519), .C2(n18518), .A(n18564), .B(n18517), .ZN(
        n18520) );
  OAI211_X1 U20680 ( .C1(n18567), .C2(n18522), .A(n18521), .B(n18520), .ZN(
        P2_U2828) );
  AOI22_X1 U20681 ( .A1(P2_REIP_REG_28__SCAN_IN), .A2(n18536), .B1(n18523), 
        .B2(n18534), .ZN(n18533) );
  AOI22_X1 U20682 ( .A1(n18538), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n18524), .ZN(n18532) );
  AOI22_X1 U20683 ( .A1(n18526), .A2(n18560), .B1(n18525), .B2(n18539), .ZN(
        n18531) );
  OAI211_X1 U20684 ( .C1(n18529), .C2(n18528), .A(n18564), .B(n18527), .ZN(
        n18530) );
  NAND4_X1 U20685 ( .A1(n18533), .A2(n18532), .A3(n18531), .A4(n18530), .ZN(
        P2_U2827) );
  AOI22_X1 U20686 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n18536), .B1(n18535), 
        .B2(n18534), .ZN(n18548) );
  AOI22_X1 U20687 ( .A1(n18538), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n18537), .ZN(n18547) );
  AOI22_X1 U20688 ( .A1(n18541), .A2(n18560), .B1(n18540), .B2(n18539), .ZN(
        n18546) );
  OAI211_X1 U20689 ( .C1(n18544), .C2(n18543), .A(n18564), .B(n18542), .ZN(
        n18545) );
  NAND4_X1 U20690 ( .A1(n18548), .A2(n18547), .A3(n18546), .A4(n18545), .ZN(
        P2_U2826) );
  INV_X1 U20691 ( .A(n18549), .ZN(n18553) );
  OAI22_X1 U20692 ( .A1(n18553), .A2(n18552), .B1(n18551), .B2(n18550), .ZN(
        n18559) );
  INV_X1 U20693 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n18555) );
  OAI22_X1 U20694 ( .A1(n18557), .A2(n18556), .B1(n18555), .B2(n18554), .ZN(
        n18558) );
  NAND4_X1 U20695 ( .A1(n18564), .A2(n18563), .A3(n18562), .A4(n18561), .ZN(
        n18565) );
  OAI211_X1 U20696 ( .C1(n16279), .C2(n18567), .A(n18566), .B(n18565), .ZN(
        P2_U2824) );
  INV_X1 U20697 ( .A(n18568), .ZN(n18569) );
  NOR3_X1 U20698 ( .A1(n18570), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n18569), .ZN(n18574) );
  AOI21_X1 U20699 ( .B1(n18585), .B2(n18572), .A(n18571), .ZN(n18573) );
  AOI211_X1 U20700 ( .C1(n18601), .C2(n19159), .A(n18574), .B(n18573), .ZN(
        n18581) );
  NAND2_X1 U20701 ( .A1(n18603), .A2(n18577), .ZN(n18578) );
  OAI211_X1 U20702 ( .C1(n12177), .C2(n18582), .A(n18581), .B(n18580), .ZN(
        P2_U3032) );
  NOR2_X1 U20703 ( .A1(n18583), .A2(n12419), .ZN(n18588) );
  INV_X1 U20704 ( .A(n18584), .ZN(n18586) );
  AOI21_X1 U20705 ( .B1(n17253), .B2(n18586), .A(n18585), .ZN(n18587) );
  AOI211_X1 U20706 ( .C1(n18601), .C2(n19166), .A(n18588), .B(n18587), .ZN(
        n18592) );
  AOI22_X1 U20707 ( .A1(n18590), .A2(n18604), .B1(n18603), .B2(n18589), .ZN(
        n18591) );
  OAI211_X1 U20708 ( .C1(n18609), .C2(n18593), .A(n18592), .B(n18591), .ZN(
        P2_U3034) );
  NAND2_X1 U20709 ( .A1(P2_REIP_REG_19__SCAN_IN), .A2(n18382), .ZN(n18594) );
  OAI21_X1 U20710 ( .B1(n18596), .B2(n18595), .A(n18594), .ZN(n18599) );
  NOR2_X1 U20711 ( .A1(n18597), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n18598) );
  AOI211_X1 U20712 ( .C1(n18601), .C2(n18600), .A(n18599), .B(n18598), .ZN(
        n18607) );
  AOI22_X1 U20713 ( .A1(n18605), .A2(n18604), .B1(n18603), .B2(n18602), .ZN(
        n18606) );
  OAI211_X1 U20714 ( .C1(n18609), .C2(n18608), .A(n18607), .B(n18606), .ZN(
        P2_U3027) );
  INV_X1 U20715 ( .A(n18611), .ZN(n18623) );
  AOI22_X1 U20716 ( .A1(n18611), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n18610), .B2(n18623), .ZN(n18651) );
  MUX2_X1 U20717 ( .A(n18612), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n18611), .Z(n18622) );
  INV_X1 U20718 ( .A(n18622), .ZN(n18650) );
  INV_X1 U20719 ( .A(n18617), .ZN(n18615) );
  INV_X1 U20720 ( .A(n18613), .ZN(n18614) );
  OAI211_X1 U20721 ( .C1(n18615), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n18614), .ZN(n18616) );
  OAI211_X1 U20722 ( .C1(n18617), .C2(n19294), .A(n18616), .B(n18623), .ZN(
        n18618) );
  AOI222_X1 U20723 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18651), 
        .B1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18618), .C1(n18651), 
        .C2(n18618), .ZN(n18621) );
  NOR2_X1 U20724 ( .A1(n18650), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18620) );
  OAI221_X1 U20725 ( .B1(n18622), .B2(n19213), .C1(n18621), .C2(n18620), .A(
        n18619), .ZN(n18649) );
  NOR2_X1 U20726 ( .A1(n18623), .A2(n14646), .ZN(n18647) );
  INV_X1 U20727 ( .A(n18624), .ZN(n18633) );
  NAND2_X1 U20728 ( .A1(n18626), .A2(n18625), .ZN(n18632) );
  INV_X1 U20729 ( .A(n18627), .ZN(n18629) );
  AOI22_X1 U20730 ( .A1(n18641), .A2(n18630), .B1(n18629), .B2(n18628), .ZN(
        n18631) );
  OAI211_X1 U20731 ( .C1(n18634), .C2(n18633), .A(n18632), .B(n18631), .ZN(
        n18635) );
  AOI21_X1 U20732 ( .B1(n18637), .B2(n18636), .A(n18635), .ZN(n18685) );
  INV_X1 U20733 ( .A(n18685), .ZN(n18646) );
  NAND4_X1 U20734 ( .A1(n18641), .A2(n18640), .A3(n18639), .A4(n18638), .ZN(
        n18682) );
  NOR2_X1 U20735 ( .A1(P2_FLUSH_REG_SCAN_IN), .A2(P2_MORE_REG_SCAN_IN), .ZN(
        n18643) );
  OAI22_X1 U20736 ( .A1(n18682), .A2(n18643), .B1(n11774), .B2(n18642), .ZN(
        n18644) );
  NOR4_X1 U20737 ( .A1(n18647), .A2(n18646), .A3(n18645), .A4(n18644), .ZN(
        n18648) );
  OAI211_X1 U20738 ( .C1(n18651), .C2(n18650), .A(n18649), .B(n18648), .ZN(
        n18678) );
  OAI21_X1 U20739 ( .B1(n18678), .B2(n18653), .A(n18652), .ZN(n18655) );
  NAND2_X1 U20740 ( .A1(n18672), .A2(n18656), .ZN(n18670) );
  NAND2_X1 U20741 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n18675), .ZN(n18659) );
  OAI21_X1 U20742 ( .B1(n18659), .B2(n18658), .A(n18657), .ZN(n18662) );
  NAND2_X1 U20743 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n21639), .ZN(n18660) );
  AOI21_X1 U20744 ( .B1(n18676), .B2(n18670), .A(n18660), .ZN(n18661) );
  AOI21_X1 U20745 ( .B1(n18670), .B2(n18662), .A(n18661), .ZN(n18664) );
  NAND2_X1 U20746 ( .A1(n18664), .A2(n18663), .ZN(P2_U3177) );
  AOI221_X1 U20747 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n18669), .C1(
        P2_STATE2_REG_3__SCAN_IN), .C2(n18672), .A(n18665), .ZN(n18666) );
  INV_X1 U20748 ( .A(n18666), .ZN(P2_U3593) );
  AOI21_X1 U20749 ( .B1(n18669), .B2(n18668), .A(n18667), .ZN(n18681) );
  INV_X1 U20750 ( .A(n18670), .ZN(n18680) );
  OAI21_X1 U20751 ( .B1(n18672), .B2(n18671), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n18673) );
  OAI211_X1 U20752 ( .C1(n18676), .C2(n18675), .A(n18674), .B(n18673), .ZN(
        n18677) );
  AOI21_X1 U20753 ( .B1(n18683), .B2(n18678), .A(n18677), .ZN(n18679) );
  OAI221_X1 U20754 ( .B1(n18681), .B2(n21639), .C1(n18681), .C2(n18680), .A(
        n18679), .ZN(P2_U3176) );
  NAND2_X1 U20755 ( .A1(n18683), .A2(n18682), .ZN(n18687) );
  NAND2_X1 U20756 ( .A1(n18687), .A2(P2_MORE_REG_SCAN_IN), .ZN(n18684) );
  OAI21_X1 U20757 ( .B1(n18687), .B2(n18685), .A(n18684), .ZN(P2_U3609) );
  AOI21_X1 U20758 ( .B1(n18687), .B2(P2_FLUSH_REG_SCAN_IN), .A(n18686), .ZN(
        n18688) );
  INV_X1 U20759 ( .A(n18688), .ZN(P2_U2819) );
  INV_X1 U20760 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n20089) );
  AOI22_X1 U20761 ( .A1(n19050), .A2(n20089), .B1(n16283), .B2(U215), .ZN(U282) );
  OAI22_X1 U20762 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19050), .ZN(n18689) );
  INV_X1 U20763 ( .A(n18689), .ZN(U281) );
  OAI22_X1 U20764 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19050), .ZN(n18690) );
  INV_X1 U20765 ( .A(n18690), .ZN(U280) );
  OAI22_X1 U20766 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n19050), .ZN(n18691) );
  INV_X1 U20767 ( .A(n18691), .ZN(U279) );
  OAI22_X1 U20768 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19050), .ZN(n18692) );
  INV_X1 U20769 ( .A(n18692), .ZN(U278) );
  OAI22_X1 U20770 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19050), .ZN(n18693) );
  INV_X1 U20771 ( .A(n18693), .ZN(U277) );
  OAI22_X1 U20772 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19050), .ZN(n18694) );
  INV_X1 U20773 ( .A(n18694), .ZN(U276) );
  OAI22_X1 U20774 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19050), .ZN(n18695) );
  INV_X1 U20775 ( .A(n18695), .ZN(U275) );
  OAI22_X1 U20776 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19050), .ZN(n18696) );
  INV_X1 U20777 ( .A(n18696), .ZN(U274) );
  OAI22_X1 U20778 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19050), .ZN(n18697) );
  INV_X1 U20779 ( .A(n18697), .ZN(U273) );
  OAI22_X1 U20780 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19050), .ZN(n18698) );
  INV_X1 U20781 ( .A(n18698), .ZN(U272) );
  OAI22_X1 U20782 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19050), .ZN(n18699) );
  INV_X1 U20783 ( .A(n18699), .ZN(U271) );
  OAI22_X1 U20784 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n18712), .ZN(n18700) );
  INV_X1 U20785 ( .A(n18700), .ZN(U270) );
  OAI22_X1 U20786 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19050), .ZN(n18701) );
  INV_X1 U20787 ( .A(n18701), .ZN(U269) );
  OAI22_X1 U20788 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n18712), .ZN(n18702) );
  INV_X1 U20789 ( .A(n18702), .ZN(U268) );
  OAI22_X1 U20790 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19050), .ZN(n18703) );
  INV_X1 U20791 ( .A(n18703), .ZN(U267) );
  OAI22_X1 U20792 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n18712), .ZN(n18704) );
  INV_X1 U20793 ( .A(n18704), .ZN(U266) );
  OAI22_X1 U20794 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n19050), .ZN(n18705) );
  INV_X1 U20795 ( .A(n18705), .ZN(U265) );
  OAI22_X1 U20796 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n18712), .ZN(n18706) );
  INV_X1 U20797 ( .A(n18706), .ZN(U264) );
  OAI22_X1 U20798 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n18712), .ZN(n18707) );
  INV_X1 U20799 ( .A(n18707), .ZN(U263) );
  OAI22_X1 U20800 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n18712), .ZN(n18708) );
  INV_X1 U20801 ( .A(n18708), .ZN(U262) );
  OAI22_X1 U20802 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n18712), .ZN(n18709) );
  INV_X1 U20803 ( .A(n18709), .ZN(U261) );
  OAI22_X1 U20804 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n18712), .ZN(n18710) );
  INV_X1 U20805 ( .A(n18710), .ZN(U260) );
  OAI22_X1 U20806 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n18712), .ZN(n18711) );
  INV_X1 U20807 ( .A(n18711), .ZN(U259) );
  OAI22_X1 U20808 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n18712), .ZN(n18713) );
  INV_X1 U20809 ( .A(n18713), .ZN(U258) );
  NAND2_X1 U20810 ( .A1(n21204), .A2(n18725), .ZN(n18724) );
  NOR2_X2 U20811 ( .A1(n18724), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19072) );
  INV_X1 U20812 ( .A(n19072), .ZN(n18966) );
  NAND2_X1 U20813 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n19053), .ZN(n18768) );
  INV_X1 U20814 ( .A(n18724), .ZN(n18716) );
  NAND2_X1 U20815 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18716), .ZN(
        n19154) );
  INV_X1 U20816 ( .A(n19154), .ZN(n19066) );
  NAND2_X1 U20817 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19053), .ZN(n18775) );
  INV_X1 U20818 ( .A(n18775), .ZN(n18789) );
  NOR2_X1 U20819 ( .A1(n21213), .A2(n18714), .ZN(n18780) );
  AND2_X1 U20820 ( .A1(n18770), .A2(n18780), .ZN(n19055) );
  INV_X1 U20821 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n20595) );
  NOR2_X2 U20822 ( .A1(n20595), .A2(n19054), .ZN(n18787) );
  AOI22_X1 U20823 ( .A1(n19066), .A2(n18789), .B1(n19055), .B2(n18787), .ZN(
        n18720) );
  NOR2_X1 U20824 ( .A1(n18715), .A2(n19054), .ZN(n18734) );
  AOI22_X1 U20825 ( .A1(n19053), .A2(n18716), .B1(n18780), .B2(n18734), .ZN(
        n19058) );
  NAND2_X1 U20826 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18780), .ZN(
        n19135) );
  INV_X1 U20827 ( .A(n19135), .ZN(n19137) );
  NAND2_X1 U20828 ( .A1(n18718), .A2(n18717), .ZN(n19056) );
  NOR2_X2 U20829 ( .A1(n20722), .A2(n19056), .ZN(n18790) );
  AOI22_X1 U20830 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19058), .B1(
        n19137), .B2(n18790), .ZN(n18719) );
  OAI211_X1 U20831 ( .C1(n18966), .C2(n18768), .A(n18720), .B(n18719), .ZN(
        P3_U2995) );
  NOR2_X1 U20832 ( .A1(n21213), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18741) );
  NAND2_X1 U20833 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18741), .ZN(
        n18732) );
  NOR2_X2 U20834 ( .A1(n21201), .A2(n18732), .ZN(n19077) );
  INV_X1 U20835 ( .A(n19077), .ZN(n19070) );
  INV_X1 U20836 ( .A(n18770), .ZN(n21224) );
  NAND2_X1 U20837 ( .A1(n21201), .A2(n18780), .ZN(n19142) );
  INV_X1 U20838 ( .A(n19142), .ZN(n19146) );
  NOR2_X1 U20839 ( .A1(n19066), .A2(n19146), .ZN(n18785) );
  NOR2_X1 U20840 ( .A1(n21224), .A2(n18785), .ZN(n19061) );
  AOI22_X1 U20841 ( .A1(n19072), .A2(n18789), .B1(n18787), .B2(n19061), .ZN(
        n18723) );
  NAND2_X1 U20842 ( .A1(n18966), .A2(n19070), .ZN(n18729) );
  INV_X1 U20843 ( .A(n18729), .ZN(n18728) );
  OAI21_X1 U20844 ( .B1(n18728), .B2(n18771), .A(n18785), .ZN(n18721) );
  OAI211_X1 U20845 ( .C1(n19146), .C2(n21232), .A(n19006), .B(n18721), .ZN(
        n19062) );
  AOI22_X1 U20846 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19062), .B1(
        n18790), .B2(n19146), .ZN(n18722) );
  OAI211_X1 U20847 ( .C1(n18768), .C2(n19070), .A(n18723), .B(n18722), .ZN(
        P3_U2987) );
  INV_X1 U20848 ( .A(n18768), .ZN(n18788) );
  INV_X1 U20849 ( .A(n18732), .ZN(n18733) );
  NAND2_X1 U20850 ( .A1(n21201), .A2(n18733), .ZN(n18971) );
  INV_X1 U20851 ( .A(n18971), .ZN(n19083) );
  NOR2_X1 U20852 ( .A1(n21224), .A2(n18724), .ZN(n19065) );
  AOI22_X1 U20853 ( .A1(n18788), .A2(n19083), .B1(n18787), .B2(n19065), .ZN(
        n18727) );
  AND2_X1 U20854 ( .A1(n21204), .A2(n18734), .ZN(n18779) );
  AOI22_X1 U20855 ( .A1(n19053), .A2(n18733), .B1(n18725), .B2(n18779), .ZN(
        n19067) );
  AOI22_X1 U20856 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19067), .B1(
        n18790), .B2(n19066), .ZN(n18726) );
  OAI211_X1 U20857 ( .C1(n18775), .C2(n19070), .A(n18727), .B(n18726), .ZN(
        P3_U2979) );
  NOR2_X1 U20858 ( .A1(n21201), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18759) );
  NAND2_X1 U20859 ( .A1(n18741), .A2(n18759), .ZN(n19081) );
  INV_X1 U20860 ( .A(n19081), .ZN(n19089) );
  NOR2_X1 U20861 ( .A1(n21224), .A2(n18728), .ZN(n19071) );
  AOI22_X1 U20862 ( .A1(n18788), .A2(n19089), .B1(n18787), .B2(n19071), .ZN(
        n18731) );
  NAND2_X1 U20863 ( .A1(n18971), .A2(n19081), .ZN(n18737) );
  OAI21_X1 U20864 ( .B1(n21232), .B2(n21201), .A(n19006), .ZN(n18784) );
  INV_X1 U20865 ( .A(n18784), .ZN(n18761) );
  AOI22_X1 U20866 ( .A1(n19053), .A2(n18737), .B1(n18761), .B2(n18729), .ZN(
        n19073) );
  AOI22_X1 U20867 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19073), .B1(
        n19072), .B2(n18790), .ZN(n18730) );
  OAI211_X1 U20868 ( .C1(n18775), .C2(n18971), .A(n18731), .B(n18730), .ZN(
        P3_U2971) );
  NAND2_X1 U20869 ( .A1(n21204), .A2(n21201), .ZN(n21206) );
  INV_X1 U20870 ( .A(n18741), .ZN(n18740) );
  NOR2_X2 U20871 ( .A1(n21206), .A2(n18740), .ZN(n19094) );
  INV_X1 U20872 ( .A(n19094), .ZN(n19087) );
  NOR2_X1 U20873 ( .A1(n21224), .A2(n18732), .ZN(n19076) );
  AOI22_X1 U20874 ( .A1(n18789), .A2(n19089), .B1(n18787), .B2(n19076), .ZN(
        n18736) );
  AOI22_X1 U20875 ( .A1(n19053), .A2(n18741), .B1(n18734), .B2(n18733), .ZN(
        n19078) );
  AOI22_X1 U20876 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19078), .B1(
        n18790), .B2(n19077), .ZN(n18735) );
  OAI211_X1 U20877 ( .C1(n18768), .C2(n19087), .A(n18736), .B(n18735), .ZN(
        P3_U2963) );
  INV_X1 U20878 ( .A(n18742), .ZN(n18749) );
  NOR2_X2 U20879 ( .A1(n21201), .A2(n18749), .ZN(n19100) );
  INV_X1 U20880 ( .A(n19100), .ZN(n19022) );
  AND2_X1 U20881 ( .A1(n18770), .A2(n18737), .ZN(n19082) );
  AOI22_X1 U20882 ( .A1(n18789), .A2(n19094), .B1(n18787), .B2(n19082), .ZN(
        n18739) );
  NAND2_X1 U20883 ( .A1(n19087), .A2(n19022), .ZN(n18746) );
  AOI22_X1 U20884 ( .A1(n19053), .A2(n18746), .B1(n18761), .B2(n18737), .ZN(
        n19084) );
  AOI22_X1 U20885 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19084), .B1(
        n18790), .B2(n19083), .ZN(n18738) );
  OAI211_X1 U20886 ( .C1(n18768), .C2(n19022), .A(n18739), .B(n18738), .ZN(
        P3_U2955) );
  NOR2_X2 U20887 ( .A1(n18749), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19106) );
  INV_X1 U20888 ( .A(n19106), .ZN(n19098) );
  NAND2_X1 U20889 ( .A1(n21204), .A2(n18770), .ZN(n18777) );
  NOR2_X1 U20890 ( .A1(n18740), .A2(n18777), .ZN(n19088) );
  AOI22_X1 U20891 ( .A1(n18789), .A2(n19100), .B1(n18787), .B2(n19088), .ZN(
        n18744) );
  AOI22_X1 U20892 ( .A1(n19053), .A2(n18742), .B1(n18741), .B2(n18779), .ZN(
        n19090) );
  AOI22_X1 U20893 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19090), .B1(
        n18790), .B2(n19089), .ZN(n18743) );
  OAI211_X1 U20894 ( .C1(n18768), .C2(n19098), .A(n18744), .B(n18743), .ZN(
        P3_U2947) );
  INV_X1 U20895 ( .A(n18759), .ZN(n18745) );
  NAND2_X1 U20896 ( .A1(n21213), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18755) );
  NOR2_X2 U20897 ( .A1(n18745), .A2(n18755), .ZN(n19112) );
  INV_X1 U20898 ( .A(n19112), .ZN(n19104) );
  AND2_X1 U20899 ( .A1(n18770), .A2(n18746), .ZN(n19093) );
  AOI22_X1 U20900 ( .A1(n18789), .A2(n19106), .B1(n18787), .B2(n19093), .ZN(
        n18748) );
  NAND2_X1 U20901 ( .A1(n19098), .A2(n19104), .ZN(n18752) );
  AOI22_X1 U20902 ( .A1(n19053), .A2(n18752), .B1(n18761), .B2(n18746), .ZN(
        n19095) );
  AOI22_X1 U20903 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19095), .B1(
        n18790), .B2(n19094), .ZN(n18747) );
  OAI211_X1 U20904 ( .C1(n18768), .C2(n19104), .A(n18748), .B(n18747), .ZN(
        P3_U2939) );
  INV_X1 U20905 ( .A(n19117), .ZN(n19110) );
  NOR2_X1 U20906 ( .A1(n21224), .A2(n18749), .ZN(n19099) );
  AOI22_X1 U20907 ( .A1(n18789), .A2(n19112), .B1(n18787), .B2(n19099), .ZN(
        n18751) );
  INV_X1 U20908 ( .A(n18755), .ZN(n18756) );
  AOI21_X1 U20909 ( .B1(n21204), .B2(n18771), .A(n19054), .ZN(n18764) );
  OAI211_X1 U20910 ( .C1(n19100), .C2(n21232), .A(n18756), .B(n18764), .ZN(
        n19101) );
  AOI22_X1 U20911 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19101), .B1(
        n18790), .B2(n19100), .ZN(n18750) );
  OAI211_X1 U20912 ( .C1(n18768), .C2(n19110), .A(n18751), .B(n18750), .ZN(
        P3_U2931) );
  NOR2_X1 U20913 ( .A1(n21204), .A2(n18776), .ZN(n18765) );
  NAND2_X1 U20914 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18765), .ZN(
        n19031) );
  INV_X1 U20915 ( .A(n19031), .ZN(n19125) );
  AND2_X1 U20916 ( .A1(n18770), .A2(n18752), .ZN(n19105) );
  AOI22_X1 U20917 ( .A1(n18788), .A2(n19125), .B1(n18787), .B2(n19105), .ZN(
        n18754) );
  NAND2_X1 U20918 ( .A1(n19110), .A2(n19031), .ZN(n18760) );
  AOI22_X1 U20919 ( .A1(n19053), .A2(n18760), .B1(n18761), .B2(n18752), .ZN(
        n19107) );
  AOI22_X1 U20920 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19107), .B1(
        n18790), .B2(n19106), .ZN(n18753) );
  OAI211_X1 U20921 ( .C1(n18775), .C2(n19110), .A(n18754), .B(n18753), .ZN(
        P3_U2923) );
  NAND2_X1 U20922 ( .A1(n21201), .A2(n18765), .ZN(n19121) );
  INV_X1 U20923 ( .A(n19121), .ZN(n19131) );
  NOR2_X1 U20924 ( .A1(n18777), .A2(n18755), .ZN(n19111) );
  AOI22_X1 U20925 ( .A1(n18788), .A2(n19131), .B1(n18787), .B2(n19111), .ZN(
        n18758) );
  AOI22_X1 U20926 ( .A1(n19053), .A2(n18765), .B1(n18779), .B2(n18756), .ZN(
        n19113) );
  AOI22_X1 U20927 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19113), .B1(
        n18790), .B2(n19112), .ZN(n18757) );
  OAI211_X1 U20928 ( .C1(n18775), .C2(n19031), .A(n18758), .B(n18757), .ZN(
        P3_U2915) );
  INV_X1 U20929 ( .A(n18790), .ZN(n18783) );
  NAND2_X1 U20930 ( .A1(n18759), .A2(n18778), .ZN(n19129) );
  INV_X1 U20931 ( .A(n19129), .ZN(n19138) );
  AND2_X1 U20932 ( .A1(n18770), .A2(n18760), .ZN(n19116) );
  AOI22_X1 U20933 ( .A1(n18788), .A2(n19138), .B1(n18787), .B2(n19116), .ZN(
        n18763) );
  NAND2_X1 U20934 ( .A1(n19121), .A2(n19129), .ZN(n18769) );
  AOI22_X1 U20935 ( .A1(n19053), .A2(n18769), .B1(n18761), .B2(n18760), .ZN(
        n19118) );
  AOI22_X1 U20936 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19118), .B1(
        n18789), .B2(n19131), .ZN(n18762) );
  OAI211_X1 U20937 ( .C1(n18783), .C2(n19110), .A(n18763), .B(n18762), .ZN(
        P3_U2907) );
  NOR2_X2 U20938 ( .A1(n21206), .A2(n18776), .ZN(n19149) );
  INV_X1 U20939 ( .A(n19149), .ZN(n19037) );
  OAI211_X1 U20940 ( .C1(n19125), .C2(n21232), .A(n18778), .B(n18764), .ZN(
        n19123) );
  AND2_X1 U20941 ( .A1(n18770), .A2(n18765), .ZN(n19122) );
  AOI22_X1 U20942 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19123), .B1(
        n18787), .B2(n19122), .ZN(n18767) );
  AOI22_X1 U20943 ( .A1(n18790), .A2(n19125), .B1(n18789), .B2(n19138), .ZN(
        n18766) );
  OAI211_X1 U20944 ( .C1(n18768), .C2(n19037), .A(n18767), .B(n18766), .ZN(
        P3_U2899) );
  AND2_X1 U20945 ( .A1(n18770), .A2(n18769), .ZN(n19130) );
  AOI22_X1 U20946 ( .A1(n18788), .A2(n19137), .B1(n18787), .B2(n19130), .ZN(
        n18774) );
  NOR2_X1 U20947 ( .A1(n19137), .A2(n19149), .ZN(n18786) );
  OAI22_X1 U20948 ( .A1(P3_STATE2_REG_3__SCAN_IN), .A2(n19129), .B1(n18786), 
        .B2(n18771), .ZN(n18772) );
  OAI21_X1 U20949 ( .B1(n19131), .B2(n18772), .A(n19006), .ZN(n19132) );
  AOI22_X1 U20950 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19132), .B1(
        n18790), .B2(n19131), .ZN(n18773) );
  OAI211_X1 U20951 ( .C1(n18775), .C2(n19037), .A(n18774), .B(n18773), .ZN(
        P3_U2891) );
  NOR2_X1 U20952 ( .A1(n18777), .A2(n18776), .ZN(n19136) );
  AOI22_X1 U20953 ( .A1(n19137), .A2(n18789), .B1(n18787), .B2(n19136), .ZN(
        n18782) );
  AOI22_X1 U20954 ( .A1(n19053), .A2(n18780), .B1(n18779), .B2(n18778), .ZN(
        n19139) );
  AOI22_X1 U20955 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19139), .B1(
        n18788), .B2(n19146), .ZN(n18781) );
  OAI211_X1 U20956 ( .C1(n18783), .C2(n19129), .A(n18782), .B(n18781), .ZN(
        P3_U2883) );
  OAI22_X1 U20957 ( .A1(n18785), .A2(n19005), .B1(n18786), .B2(n18784), .ZN(
        n19147) );
  NOR2_X1 U20958 ( .A1(n21224), .A2(n18786), .ZN(n19144) );
  AOI22_X1 U20959 ( .A1(n18788), .A2(n19066), .B1(n18787), .B2(n19144), .ZN(
        n18792) );
  AOI22_X1 U20960 ( .A1(n18790), .A2(n19149), .B1(n18789), .B2(n19146), .ZN(
        n18791) );
  OAI211_X1 U20961 ( .C1(n18793), .C2(n19147), .A(n18792), .B(n18791), .ZN(
        P3_U2875) );
  OAI22_X1 U20962 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n19050), .ZN(n18794) );
  INV_X1 U20963 ( .A(n18794), .ZN(U257) );
  INV_X1 U20964 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n18795) );
  NOR2_X1 U20965 ( .A1(n18795), .A2(n19005), .ZN(n18832) );
  INV_X1 U20966 ( .A(n18832), .ZN(n18823) );
  NAND2_X1 U20967 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19053), .ZN(n18828) );
  INV_X1 U20968 ( .A(n18828), .ZN(n18830) );
  NOR2_X2 U20969 ( .A1(n20600), .A2(n19054), .ZN(n18829) );
  AOI22_X1 U20970 ( .A1(n19072), .A2(n18830), .B1(n19055), .B2(n18829), .ZN(
        n18798) );
  NOR2_X2 U20971 ( .A1(n18796), .A2(n19056), .ZN(n18831) );
  AOI22_X1 U20972 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19058), .B1(
        n19137), .B2(n18831), .ZN(n18797) );
  OAI211_X1 U20973 ( .C1(n19154), .C2(n18823), .A(n18798), .B(n18797), .ZN(
        P3_U2994) );
  AOI22_X1 U20974 ( .A1(n19077), .A2(n18830), .B1(n19061), .B2(n18829), .ZN(
        n18800) );
  AOI22_X1 U20975 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19062), .B1(
        n19146), .B2(n18831), .ZN(n18799) );
  OAI211_X1 U20976 ( .C1(n18966), .C2(n18823), .A(n18800), .B(n18799), .ZN(
        P3_U2986) );
  AOI22_X1 U20977 ( .A1(n19077), .A2(n18832), .B1(n19065), .B2(n18829), .ZN(
        n18802) );
  AOI22_X1 U20978 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19067), .B1(
        n19066), .B2(n18831), .ZN(n18801) );
  OAI211_X1 U20979 ( .C1(n18971), .C2(n18828), .A(n18802), .B(n18801), .ZN(
        P3_U2978) );
  AOI22_X1 U20980 ( .A1(n19083), .A2(n18832), .B1(n19071), .B2(n18829), .ZN(
        n18804) );
  AOI22_X1 U20981 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19073), .B1(
        n19072), .B2(n18831), .ZN(n18803) );
  OAI211_X1 U20982 ( .C1(n19081), .C2(n18828), .A(n18804), .B(n18803), .ZN(
        P3_U2970) );
  AOI22_X1 U20983 ( .A1(n19089), .A2(n18832), .B1(n19076), .B2(n18829), .ZN(
        n18806) );
  AOI22_X1 U20984 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19078), .B1(
        n19077), .B2(n18831), .ZN(n18805) );
  OAI211_X1 U20985 ( .C1(n19087), .C2(n18828), .A(n18806), .B(n18805), .ZN(
        P3_U2962) );
  AOI22_X1 U20986 ( .A1(n19100), .A2(n18830), .B1(n19082), .B2(n18829), .ZN(
        n18808) );
  AOI22_X1 U20987 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19084), .B1(
        n19083), .B2(n18831), .ZN(n18807) );
  OAI211_X1 U20988 ( .C1(n19087), .C2(n18823), .A(n18808), .B(n18807), .ZN(
        P3_U2954) );
  AOI22_X1 U20989 ( .A1(n19100), .A2(n18832), .B1(n19088), .B2(n18829), .ZN(
        n18810) );
  AOI22_X1 U20990 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19090), .B1(
        n19089), .B2(n18831), .ZN(n18809) );
  OAI211_X1 U20991 ( .C1(n19098), .C2(n18828), .A(n18810), .B(n18809), .ZN(
        P3_U2946) );
  AOI22_X1 U20992 ( .A1(n19106), .A2(n18832), .B1(n19093), .B2(n18829), .ZN(
        n18812) );
  AOI22_X1 U20993 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19095), .B1(
        n19094), .B2(n18831), .ZN(n18811) );
  OAI211_X1 U20994 ( .C1(n19104), .C2(n18828), .A(n18812), .B(n18811), .ZN(
        P3_U2938) );
  AOI22_X1 U20995 ( .A1(n19117), .A2(n18830), .B1(n19099), .B2(n18829), .ZN(
        n18814) );
  AOI22_X1 U20996 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19101), .B1(
        n19100), .B2(n18831), .ZN(n18813) );
  OAI211_X1 U20997 ( .C1(n19104), .C2(n18823), .A(n18814), .B(n18813), .ZN(
        P3_U2930) );
  AOI22_X1 U20998 ( .A1(n19125), .A2(n18830), .B1(n19105), .B2(n18829), .ZN(
        n18816) );
  AOI22_X1 U20999 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19107), .B1(
        n19106), .B2(n18831), .ZN(n18815) );
  OAI211_X1 U21000 ( .C1(n19110), .C2(n18823), .A(n18816), .B(n18815), .ZN(
        P3_U2922) );
  AOI22_X1 U21001 ( .A1(n19111), .A2(n18829), .B1(n19131), .B2(n18830), .ZN(
        n18818) );
  AOI22_X1 U21002 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19113), .B1(
        n19112), .B2(n18831), .ZN(n18817) );
  OAI211_X1 U21003 ( .C1(n19031), .C2(n18823), .A(n18818), .B(n18817), .ZN(
        P3_U2914) );
  AOI22_X1 U21004 ( .A1(n19131), .A2(n18832), .B1(n19116), .B2(n18829), .ZN(
        n18820) );
  AOI22_X1 U21005 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19118), .B1(
        n19117), .B2(n18831), .ZN(n18819) );
  OAI211_X1 U21006 ( .C1(n19129), .C2(n18828), .A(n18820), .B(n18819), .ZN(
        P3_U2906) );
  AOI22_X1 U21007 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19123), .B1(
        n19122), .B2(n18829), .ZN(n18822) );
  AOI22_X1 U21008 ( .A1(n19125), .A2(n18831), .B1(n19149), .B2(n18830), .ZN(
        n18821) );
  OAI211_X1 U21009 ( .C1(n19129), .C2(n18823), .A(n18822), .B(n18821), .ZN(
        P3_U2898) );
  AOI22_X1 U21010 ( .A1(n19149), .A2(n18832), .B1(n19130), .B2(n18829), .ZN(
        n18825) );
  AOI22_X1 U21011 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19132), .B1(
        n19131), .B2(n18831), .ZN(n18824) );
  OAI211_X1 U21012 ( .C1(n19135), .C2(n18828), .A(n18825), .B(n18824), .ZN(
        P3_U2890) );
  AOI22_X1 U21013 ( .A1(n19137), .A2(n18832), .B1(n19136), .B2(n18829), .ZN(
        n18827) );
  AOI22_X1 U21014 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19139), .B1(
        n19138), .B2(n18831), .ZN(n18826) );
  OAI211_X1 U21015 ( .C1(n19142), .C2(n18828), .A(n18827), .B(n18826), .ZN(
        P3_U2882) );
  AOI22_X1 U21016 ( .A1(n19066), .A2(n18830), .B1(n19144), .B2(n18829), .ZN(
        n18834) );
  AOI22_X1 U21017 ( .A1(n19146), .A2(n18832), .B1(n19149), .B2(n18831), .ZN(
        n18833) );
  OAI211_X1 U21018 ( .C1(n18835), .C2(n19147), .A(n18834), .B(n18833), .ZN(
        P3_U2874) );
  OAI22_X1 U21019 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n19050), .ZN(n18836) );
  INV_X1 U21020 ( .A(n18836), .ZN(U256) );
  INV_X1 U21021 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n20626) );
  NOR2_X1 U21022 ( .A1(n20626), .A2(n19005), .ZN(n18873) );
  INV_X1 U21023 ( .A(n18873), .ZN(n18869) );
  NAND2_X1 U21024 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19053), .ZN(n18862) );
  INV_X1 U21025 ( .A(n18862), .ZN(n18871) );
  INV_X1 U21026 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n20605) );
  NOR2_X2 U21027 ( .A1(n20605), .A2(n19054), .ZN(n18870) );
  AOI22_X1 U21028 ( .A1(n19072), .A2(n18871), .B1(n19055), .B2(n18870), .ZN(
        n18839) );
  NOR2_X2 U21029 ( .A1(n18837), .A2(n19056), .ZN(n18872) );
  AOI22_X1 U21030 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19058), .B1(
        n19137), .B2(n18872), .ZN(n18838) );
  OAI211_X1 U21031 ( .C1(n19154), .C2(n18869), .A(n18839), .B(n18838), .ZN(
        P3_U2993) );
  AOI22_X1 U21032 ( .A1(n19072), .A2(n18873), .B1(n19061), .B2(n18870), .ZN(
        n18841) );
  AOI22_X1 U21033 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19062), .B1(
        n19146), .B2(n18872), .ZN(n18840) );
  OAI211_X1 U21034 ( .C1(n19070), .C2(n18862), .A(n18841), .B(n18840), .ZN(
        P3_U2985) );
  AOI22_X1 U21035 ( .A1(n19077), .A2(n18873), .B1(n19065), .B2(n18870), .ZN(
        n18843) );
  AOI22_X1 U21036 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19067), .B1(
        n19066), .B2(n18872), .ZN(n18842) );
  OAI211_X1 U21037 ( .C1(n18971), .C2(n18862), .A(n18843), .B(n18842), .ZN(
        P3_U2977) );
  AOI22_X1 U21038 ( .A1(n19089), .A2(n18871), .B1(n19071), .B2(n18870), .ZN(
        n18845) );
  AOI22_X1 U21039 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19073), .B1(
        n19072), .B2(n18872), .ZN(n18844) );
  OAI211_X1 U21040 ( .C1(n18971), .C2(n18869), .A(n18845), .B(n18844), .ZN(
        P3_U2969) );
  AOI22_X1 U21041 ( .A1(n19089), .A2(n18873), .B1(n19076), .B2(n18870), .ZN(
        n18847) );
  AOI22_X1 U21042 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19078), .B1(
        n19077), .B2(n18872), .ZN(n18846) );
  OAI211_X1 U21043 ( .C1(n19087), .C2(n18862), .A(n18847), .B(n18846), .ZN(
        P3_U2961) );
  AOI22_X1 U21044 ( .A1(n19100), .A2(n18871), .B1(n19082), .B2(n18870), .ZN(
        n18849) );
  AOI22_X1 U21045 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19084), .B1(
        n19083), .B2(n18872), .ZN(n18848) );
  OAI211_X1 U21046 ( .C1(n19087), .C2(n18869), .A(n18849), .B(n18848), .ZN(
        P3_U2953) );
  AOI22_X1 U21047 ( .A1(n19100), .A2(n18873), .B1(n19088), .B2(n18870), .ZN(
        n18851) );
  AOI22_X1 U21048 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19090), .B1(
        n19089), .B2(n18872), .ZN(n18850) );
  OAI211_X1 U21049 ( .C1(n19098), .C2(n18862), .A(n18851), .B(n18850), .ZN(
        P3_U2945) );
  AOI22_X1 U21050 ( .A1(n19112), .A2(n18871), .B1(n19093), .B2(n18870), .ZN(
        n18853) );
  AOI22_X1 U21051 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19095), .B1(
        n19094), .B2(n18872), .ZN(n18852) );
  OAI211_X1 U21052 ( .C1(n19098), .C2(n18869), .A(n18853), .B(n18852), .ZN(
        P3_U2937) );
  AOI22_X1 U21053 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19101), .B1(
        n19099), .B2(n18870), .ZN(n18855) );
  AOI22_X1 U21054 ( .A1(n19100), .A2(n18872), .B1(n19117), .B2(n18871), .ZN(
        n18854) );
  OAI211_X1 U21055 ( .C1(n19104), .C2(n18869), .A(n18855), .B(n18854), .ZN(
        P3_U2929) );
  AOI22_X1 U21056 ( .A1(n19117), .A2(n18873), .B1(n19105), .B2(n18870), .ZN(
        n18857) );
  AOI22_X1 U21057 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19107), .B1(
        n19106), .B2(n18872), .ZN(n18856) );
  OAI211_X1 U21058 ( .C1(n19031), .C2(n18862), .A(n18857), .B(n18856), .ZN(
        P3_U2921) );
  AOI22_X1 U21059 ( .A1(n19125), .A2(n18873), .B1(n19111), .B2(n18870), .ZN(
        n18859) );
  AOI22_X1 U21060 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19113), .B1(
        n19112), .B2(n18872), .ZN(n18858) );
  OAI211_X1 U21061 ( .C1(n19121), .C2(n18862), .A(n18859), .B(n18858), .ZN(
        P3_U2913) );
  AOI22_X1 U21062 ( .A1(n19131), .A2(n18873), .B1(n19116), .B2(n18870), .ZN(
        n18861) );
  AOI22_X1 U21063 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19118), .B1(
        n19117), .B2(n18872), .ZN(n18860) );
  OAI211_X1 U21064 ( .C1(n19129), .C2(n18862), .A(n18861), .B(n18860), .ZN(
        P3_U2905) );
  AOI22_X1 U21065 ( .A1(n19149), .A2(n18871), .B1(n19122), .B2(n18870), .ZN(
        n18864) );
  AOI22_X1 U21066 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19123), .B1(
        n19125), .B2(n18872), .ZN(n18863) );
  OAI211_X1 U21067 ( .C1(n19129), .C2(n18869), .A(n18864), .B(n18863), .ZN(
        P3_U2897) );
  AOI22_X1 U21068 ( .A1(n19137), .A2(n18871), .B1(n19130), .B2(n18870), .ZN(
        n18866) );
  AOI22_X1 U21069 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19132), .B1(
        n19131), .B2(n18872), .ZN(n18865) );
  OAI211_X1 U21070 ( .C1(n19037), .C2(n18869), .A(n18866), .B(n18865), .ZN(
        P3_U2889) );
  AOI22_X1 U21071 ( .A1(n19146), .A2(n18871), .B1(n19136), .B2(n18870), .ZN(
        n18868) );
  AOI22_X1 U21072 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19139), .B1(
        n19138), .B2(n18872), .ZN(n18867) );
  OAI211_X1 U21073 ( .C1(n19135), .C2(n18869), .A(n18868), .B(n18867), .ZN(
        P3_U2881) );
  AOI22_X1 U21074 ( .A1(n19066), .A2(n18871), .B1(n19144), .B2(n18870), .ZN(
        n18875) );
  AOI22_X1 U21075 ( .A1(n19146), .A2(n18873), .B1(n19149), .B2(n18872), .ZN(
        n18874) );
  OAI211_X1 U21076 ( .C1(n18876), .C2(n19147), .A(n18875), .B(n18874), .ZN(
        P3_U2873) );
  OAI22_X1 U21077 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n19050), .ZN(n18877) );
  INV_X1 U21078 ( .A(n18877), .ZN(U255) );
  INV_X1 U21079 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n19463) );
  NOR2_X1 U21080 ( .A1(n19463), .A2(n19005), .ZN(n18912) );
  INV_X1 U21081 ( .A(n18912), .ZN(n18910) );
  NAND2_X1 U21082 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19053), .ZN(n18907) );
  INV_X1 U21083 ( .A(n18907), .ZN(n18914) );
  NOR2_X2 U21084 ( .A1(n20611), .A2(n19054), .ZN(n18911) );
  AOI22_X1 U21085 ( .A1(n19072), .A2(n18914), .B1(n19055), .B2(n18911), .ZN(
        n18880) );
  NOR2_X2 U21086 ( .A1(n18878), .A2(n19056), .ZN(n18913) );
  AOI22_X1 U21087 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19058), .B1(
        n19137), .B2(n18913), .ZN(n18879) );
  OAI211_X1 U21088 ( .C1(n19154), .C2(n18910), .A(n18880), .B(n18879), .ZN(
        P3_U2992) );
  AOI22_X1 U21089 ( .A1(n19077), .A2(n18914), .B1(n19061), .B2(n18911), .ZN(
        n18882) );
  AOI22_X1 U21090 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19062), .B1(
        n19146), .B2(n18913), .ZN(n18881) );
  OAI211_X1 U21091 ( .C1(n18966), .C2(n18910), .A(n18882), .B(n18881), .ZN(
        P3_U2984) );
  AOI22_X1 U21092 ( .A1(n19065), .A2(n18911), .B1(n19083), .B2(n18914), .ZN(
        n18884) );
  AOI22_X1 U21093 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19067), .B1(
        n19066), .B2(n18913), .ZN(n18883) );
  OAI211_X1 U21094 ( .C1(n19070), .C2(n18910), .A(n18884), .B(n18883), .ZN(
        P3_U2976) );
  AOI22_X1 U21095 ( .A1(n19089), .A2(n18914), .B1(n19071), .B2(n18911), .ZN(
        n18886) );
  AOI22_X1 U21096 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19073), .B1(
        n19072), .B2(n18913), .ZN(n18885) );
  OAI211_X1 U21097 ( .C1(n18971), .C2(n18910), .A(n18886), .B(n18885), .ZN(
        P3_U2968) );
  AOI22_X1 U21098 ( .A1(n19089), .A2(n18912), .B1(n19076), .B2(n18911), .ZN(
        n18888) );
  AOI22_X1 U21099 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19078), .B1(
        n19077), .B2(n18913), .ZN(n18887) );
  OAI211_X1 U21100 ( .C1(n19087), .C2(n18907), .A(n18888), .B(n18887), .ZN(
        P3_U2960) );
  AOI22_X1 U21101 ( .A1(n19094), .A2(n18912), .B1(n19082), .B2(n18911), .ZN(
        n18890) );
  AOI22_X1 U21102 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19084), .B1(
        n19083), .B2(n18913), .ZN(n18889) );
  OAI211_X1 U21103 ( .C1(n19022), .C2(n18907), .A(n18890), .B(n18889), .ZN(
        P3_U2952) );
  AOI22_X1 U21104 ( .A1(n19100), .A2(n18912), .B1(n19088), .B2(n18911), .ZN(
        n18892) );
  AOI22_X1 U21105 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19090), .B1(
        n19089), .B2(n18913), .ZN(n18891) );
  OAI211_X1 U21106 ( .C1(n19098), .C2(n18907), .A(n18892), .B(n18891), .ZN(
        P3_U2944) );
  AOI22_X1 U21107 ( .A1(n19106), .A2(n18912), .B1(n19093), .B2(n18911), .ZN(
        n18894) );
  AOI22_X1 U21108 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19095), .B1(
        n19094), .B2(n18913), .ZN(n18893) );
  OAI211_X1 U21109 ( .C1(n19104), .C2(n18907), .A(n18894), .B(n18893), .ZN(
        P3_U2936) );
  AOI22_X1 U21110 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19101), .B1(
        n19099), .B2(n18911), .ZN(n18896) );
  AOI22_X1 U21111 ( .A1(n19100), .A2(n18913), .B1(n19112), .B2(n18912), .ZN(
        n18895) );
  OAI211_X1 U21112 ( .C1(n19110), .C2(n18907), .A(n18896), .B(n18895), .ZN(
        P3_U2928) );
  AOI22_X1 U21113 ( .A1(n19125), .A2(n18914), .B1(n19105), .B2(n18911), .ZN(
        n18898) );
  AOI22_X1 U21114 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19107), .B1(
        n19106), .B2(n18913), .ZN(n18897) );
  OAI211_X1 U21115 ( .C1(n19110), .C2(n18910), .A(n18898), .B(n18897), .ZN(
        P3_U2920) );
  AOI22_X1 U21116 ( .A1(n19111), .A2(n18911), .B1(n19131), .B2(n18914), .ZN(
        n18900) );
  AOI22_X1 U21117 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19113), .B1(
        n19112), .B2(n18913), .ZN(n18899) );
  OAI211_X1 U21118 ( .C1(n19031), .C2(n18910), .A(n18900), .B(n18899), .ZN(
        P3_U2912) );
  AOI22_X1 U21119 ( .A1(n19138), .A2(n18914), .B1(n19116), .B2(n18911), .ZN(
        n18902) );
  AOI22_X1 U21120 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19118), .B1(
        n19117), .B2(n18913), .ZN(n18901) );
  OAI211_X1 U21121 ( .C1(n19121), .C2(n18910), .A(n18902), .B(n18901), .ZN(
        P3_U2904) );
  AOI22_X1 U21122 ( .A1(n19149), .A2(n18914), .B1(n19122), .B2(n18911), .ZN(
        n18904) );
  AOI22_X1 U21123 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19123), .B1(
        n19125), .B2(n18913), .ZN(n18903) );
  OAI211_X1 U21124 ( .C1(n19129), .C2(n18910), .A(n18904), .B(n18903), .ZN(
        P3_U2896) );
  AOI22_X1 U21125 ( .A1(n19149), .A2(n18912), .B1(n19130), .B2(n18911), .ZN(
        n18906) );
  AOI22_X1 U21126 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19132), .B1(
        n19131), .B2(n18913), .ZN(n18905) );
  OAI211_X1 U21127 ( .C1(n19135), .C2(n18907), .A(n18906), .B(n18905), .ZN(
        P3_U2888) );
  AOI22_X1 U21128 ( .A1(n19146), .A2(n18914), .B1(n19136), .B2(n18911), .ZN(
        n18909) );
  AOI22_X1 U21129 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19139), .B1(
        n19138), .B2(n18913), .ZN(n18908) );
  OAI211_X1 U21130 ( .C1(n19135), .C2(n18910), .A(n18909), .B(n18908), .ZN(
        P3_U2880) );
  AOI22_X1 U21131 ( .A1(n19146), .A2(n18912), .B1(n19144), .B2(n18911), .ZN(
        n18916) );
  AOI22_X1 U21132 ( .A1(n19066), .A2(n18914), .B1(n19149), .B2(n18913), .ZN(
        n18915) );
  OAI211_X1 U21133 ( .C1(n18917), .C2(n19147), .A(n18916), .B(n18915), .ZN(
        P3_U2872) );
  OAI22_X1 U21134 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n19050), .ZN(n18918) );
  INV_X1 U21135 ( .A(n18918), .ZN(U254) );
  NAND2_X1 U21136 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19053), .ZN(n18951) );
  NAND2_X1 U21137 ( .A1(BUF2_REG_19__SCAN_IN), .A2(n19053), .ZN(n18946) );
  INV_X1 U21138 ( .A(n18946), .ZN(n18953) );
  AND2_X1 U21139 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n19006), .ZN(n18952) );
  AOI22_X1 U21140 ( .A1(n19066), .A2(n18953), .B1(n19055), .B2(n18952), .ZN(
        n18921) );
  NOR2_X2 U21141 ( .A1(n18919), .A2(n19056), .ZN(n18954) );
  AOI22_X1 U21142 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19058), .B1(
        n19137), .B2(n18954), .ZN(n18920) );
  OAI211_X1 U21143 ( .C1(n18966), .C2(n18951), .A(n18921), .B(n18920), .ZN(
        P3_U2991) );
  INV_X1 U21144 ( .A(n18951), .ZN(n18955) );
  AOI22_X1 U21145 ( .A1(n19077), .A2(n18955), .B1(n19061), .B2(n18952), .ZN(
        n18923) );
  AOI22_X1 U21146 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19062), .B1(
        n19146), .B2(n18954), .ZN(n18922) );
  OAI211_X1 U21147 ( .C1(n18966), .C2(n18946), .A(n18923), .B(n18922), .ZN(
        P3_U2983) );
  AOI22_X1 U21148 ( .A1(n19065), .A2(n18952), .B1(n19083), .B2(n18955), .ZN(
        n18925) );
  AOI22_X1 U21149 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19067), .B1(
        n19066), .B2(n18954), .ZN(n18924) );
  OAI211_X1 U21150 ( .C1(n19070), .C2(n18946), .A(n18925), .B(n18924), .ZN(
        P3_U2975) );
  AOI22_X1 U21151 ( .A1(n19083), .A2(n18953), .B1(n19071), .B2(n18952), .ZN(
        n18927) );
  AOI22_X1 U21152 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19073), .B1(
        n19072), .B2(n18954), .ZN(n18926) );
  OAI211_X1 U21153 ( .C1(n19081), .C2(n18951), .A(n18927), .B(n18926), .ZN(
        P3_U2967) );
  AOI22_X1 U21154 ( .A1(n19094), .A2(n18955), .B1(n19076), .B2(n18952), .ZN(
        n18929) );
  AOI22_X1 U21155 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19078), .B1(
        n19077), .B2(n18954), .ZN(n18928) );
  OAI211_X1 U21156 ( .C1(n19081), .C2(n18946), .A(n18929), .B(n18928), .ZN(
        P3_U2959) );
  AOI22_X1 U21157 ( .A1(n19094), .A2(n18953), .B1(n19082), .B2(n18952), .ZN(
        n18931) );
  AOI22_X1 U21158 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19084), .B1(
        n19083), .B2(n18954), .ZN(n18930) );
  OAI211_X1 U21159 ( .C1(n19022), .C2(n18951), .A(n18931), .B(n18930), .ZN(
        P3_U2951) );
  AOI22_X1 U21160 ( .A1(n19106), .A2(n18955), .B1(n19088), .B2(n18952), .ZN(
        n18933) );
  AOI22_X1 U21161 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19090), .B1(
        n19089), .B2(n18954), .ZN(n18932) );
  OAI211_X1 U21162 ( .C1(n19022), .C2(n18946), .A(n18933), .B(n18932), .ZN(
        P3_U2943) );
  AOI22_X1 U21163 ( .A1(n19106), .A2(n18953), .B1(n19093), .B2(n18952), .ZN(
        n18935) );
  AOI22_X1 U21164 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19095), .B1(
        n19094), .B2(n18954), .ZN(n18934) );
  OAI211_X1 U21165 ( .C1(n19104), .C2(n18951), .A(n18935), .B(n18934), .ZN(
        P3_U2935) );
  AOI22_X1 U21166 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19101), .B1(
        n19099), .B2(n18952), .ZN(n18937) );
  AOI22_X1 U21167 ( .A1(n19100), .A2(n18954), .B1(n19117), .B2(n18955), .ZN(
        n18936) );
  OAI211_X1 U21168 ( .C1(n19104), .C2(n18946), .A(n18937), .B(n18936), .ZN(
        P3_U2927) );
  AOI22_X1 U21169 ( .A1(n19125), .A2(n18955), .B1(n19105), .B2(n18952), .ZN(
        n18939) );
  AOI22_X1 U21170 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19107), .B1(
        n19106), .B2(n18954), .ZN(n18938) );
  OAI211_X1 U21171 ( .C1(n19110), .C2(n18946), .A(n18939), .B(n18938), .ZN(
        P3_U2919) );
  AOI22_X1 U21172 ( .A1(n19111), .A2(n18952), .B1(n19131), .B2(n18955), .ZN(
        n18941) );
  AOI22_X1 U21173 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19113), .B1(
        n19112), .B2(n18954), .ZN(n18940) );
  OAI211_X1 U21174 ( .C1(n19031), .C2(n18946), .A(n18941), .B(n18940), .ZN(
        P3_U2911) );
  AOI22_X1 U21175 ( .A1(n19131), .A2(n18953), .B1(n19116), .B2(n18952), .ZN(
        n18943) );
  AOI22_X1 U21176 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19118), .B1(
        n19117), .B2(n18954), .ZN(n18942) );
  OAI211_X1 U21177 ( .C1(n19129), .C2(n18951), .A(n18943), .B(n18942), .ZN(
        P3_U2903) );
  AOI22_X1 U21178 ( .A1(n19149), .A2(n18955), .B1(n19122), .B2(n18952), .ZN(
        n18945) );
  AOI22_X1 U21179 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19123), .B1(
        n19125), .B2(n18954), .ZN(n18944) );
  OAI211_X1 U21180 ( .C1(n19129), .C2(n18946), .A(n18945), .B(n18944), .ZN(
        P3_U2895) );
  AOI22_X1 U21181 ( .A1(n19149), .A2(n18953), .B1(n19130), .B2(n18952), .ZN(
        n18948) );
  AOI22_X1 U21182 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19132), .B1(
        n19131), .B2(n18954), .ZN(n18947) );
  OAI211_X1 U21183 ( .C1(n19135), .C2(n18951), .A(n18948), .B(n18947), .ZN(
        P3_U2887) );
  AOI22_X1 U21184 ( .A1(n19137), .A2(n18953), .B1(n19136), .B2(n18952), .ZN(
        n18950) );
  AOI22_X1 U21185 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19139), .B1(
        n19138), .B2(n18954), .ZN(n18949) );
  OAI211_X1 U21186 ( .C1(n19142), .C2(n18951), .A(n18950), .B(n18949), .ZN(
        P3_U2879) );
  AOI22_X1 U21187 ( .A1(n19146), .A2(n18953), .B1(n19144), .B2(n18952), .ZN(
        n18957) );
  AOI22_X1 U21188 ( .A1(n19066), .A2(n18955), .B1(n19149), .B2(n18954), .ZN(
        n18956) );
  OAI211_X1 U21189 ( .C1(n18958), .C2(n19147), .A(n18957), .B(n18956), .ZN(
        P3_U2871) );
  OAI22_X1 U21190 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n19050), .ZN(n18959) );
  INV_X1 U21191 ( .A(n18959), .ZN(U253) );
  INV_X1 U21192 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n18960) );
  NOR2_X1 U21193 ( .A1(n19005), .A2(n18960), .ZN(n18999) );
  INV_X1 U21194 ( .A(n18999), .ZN(n18992) );
  NAND2_X1 U21195 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19053), .ZN(n18995) );
  INV_X1 U21196 ( .A(n18995), .ZN(n18997) );
  AND2_X1 U21197 ( .A1(n19006), .A2(BUF2_REG_2__SCAN_IN), .ZN(n18996) );
  AOI22_X1 U21198 ( .A1(n19072), .A2(n18997), .B1(n19055), .B2(n18996), .ZN(
        n18963) );
  NOR2_X2 U21199 ( .A1(n18961), .A2(n19056), .ZN(n18998) );
  AOI22_X1 U21200 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19058), .B1(
        n19137), .B2(n18998), .ZN(n18962) );
  OAI211_X1 U21201 ( .C1(n19154), .C2(n18992), .A(n18963), .B(n18962), .ZN(
        P3_U2990) );
  AOI22_X1 U21202 ( .A1(n19077), .A2(n18997), .B1(n19061), .B2(n18996), .ZN(
        n18965) );
  AOI22_X1 U21203 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19062), .B1(
        n19146), .B2(n18998), .ZN(n18964) );
  OAI211_X1 U21204 ( .C1(n18966), .C2(n18992), .A(n18965), .B(n18964), .ZN(
        P3_U2982) );
  AOI22_X1 U21205 ( .A1(n19065), .A2(n18996), .B1(n19083), .B2(n18997), .ZN(
        n18968) );
  AOI22_X1 U21206 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19067), .B1(
        n19066), .B2(n18998), .ZN(n18967) );
  OAI211_X1 U21207 ( .C1(n19070), .C2(n18992), .A(n18968), .B(n18967), .ZN(
        P3_U2974) );
  AOI22_X1 U21208 ( .A1(n19089), .A2(n18997), .B1(n19071), .B2(n18996), .ZN(
        n18970) );
  AOI22_X1 U21209 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19073), .B1(
        n19072), .B2(n18998), .ZN(n18969) );
  OAI211_X1 U21210 ( .C1(n18971), .C2(n18992), .A(n18970), .B(n18969), .ZN(
        P3_U2966) );
  AOI22_X1 U21211 ( .A1(n19089), .A2(n18999), .B1(n19076), .B2(n18996), .ZN(
        n18973) );
  AOI22_X1 U21212 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19078), .B1(
        n19077), .B2(n18998), .ZN(n18972) );
  OAI211_X1 U21213 ( .C1(n19087), .C2(n18995), .A(n18973), .B(n18972), .ZN(
        P3_U2958) );
  AOI22_X1 U21214 ( .A1(n19094), .A2(n18999), .B1(n19082), .B2(n18996), .ZN(
        n18975) );
  AOI22_X1 U21215 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19084), .B1(
        n19083), .B2(n18998), .ZN(n18974) );
  OAI211_X1 U21216 ( .C1(n19022), .C2(n18995), .A(n18975), .B(n18974), .ZN(
        P3_U2950) );
  AOI22_X1 U21217 ( .A1(n19100), .A2(n18999), .B1(n19088), .B2(n18996), .ZN(
        n18977) );
  AOI22_X1 U21218 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19090), .B1(
        n19089), .B2(n18998), .ZN(n18976) );
  OAI211_X1 U21219 ( .C1(n19098), .C2(n18995), .A(n18977), .B(n18976), .ZN(
        P3_U2942) );
  AOI22_X1 U21220 ( .A1(n19112), .A2(n18997), .B1(n19093), .B2(n18996), .ZN(
        n18979) );
  AOI22_X1 U21221 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19095), .B1(
        n19094), .B2(n18998), .ZN(n18978) );
  OAI211_X1 U21222 ( .C1(n19098), .C2(n18992), .A(n18979), .B(n18978), .ZN(
        P3_U2934) );
  AOI22_X1 U21223 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19101), .B1(
        n19099), .B2(n18996), .ZN(n18981) );
  AOI22_X1 U21224 ( .A1(n19100), .A2(n18998), .B1(n19112), .B2(n18999), .ZN(
        n18980) );
  OAI211_X1 U21225 ( .C1(n19110), .C2(n18995), .A(n18981), .B(n18980), .ZN(
        P3_U2926) );
  AOI22_X1 U21226 ( .A1(n19125), .A2(n18997), .B1(n19105), .B2(n18996), .ZN(
        n18983) );
  AOI22_X1 U21227 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19107), .B1(
        n19106), .B2(n18998), .ZN(n18982) );
  OAI211_X1 U21228 ( .C1(n19110), .C2(n18992), .A(n18983), .B(n18982), .ZN(
        P3_U2918) );
  AOI22_X1 U21229 ( .A1(n19111), .A2(n18996), .B1(n19131), .B2(n18997), .ZN(
        n18985) );
  AOI22_X1 U21230 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19113), .B1(
        n19112), .B2(n18998), .ZN(n18984) );
  OAI211_X1 U21231 ( .C1(n19031), .C2(n18992), .A(n18985), .B(n18984), .ZN(
        P3_U2910) );
  AOI22_X1 U21232 ( .A1(n19131), .A2(n18999), .B1(n19116), .B2(n18996), .ZN(
        n18987) );
  AOI22_X1 U21233 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19118), .B1(
        n19117), .B2(n18998), .ZN(n18986) );
  OAI211_X1 U21234 ( .C1(n19129), .C2(n18995), .A(n18987), .B(n18986), .ZN(
        P3_U2902) );
  AOI22_X1 U21235 ( .A1(n19138), .A2(n18999), .B1(n19122), .B2(n18996), .ZN(
        n18989) );
  AOI22_X1 U21236 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19123), .B1(
        n19125), .B2(n18998), .ZN(n18988) );
  OAI211_X1 U21237 ( .C1(n19037), .C2(n18995), .A(n18989), .B(n18988), .ZN(
        P3_U2894) );
  AOI22_X1 U21238 ( .A1(n19137), .A2(n18997), .B1(n19130), .B2(n18996), .ZN(
        n18991) );
  AOI22_X1 U21239 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19132), .B1(
        n19131), .B2(n18998), .ZN(n18990) );
  OAI211_X1 U21240 ( .C1(n19037), .C2(n18992), .A(n18991), .B(n18990), .ZN(
        P3_U2886) );
  AOI22_X1 U21241 ( .A1(n19137), .A2(n18999), .B1(n19136), .B2(n18996), .ZN(
        n18994) );
  AOI22_X1 U21242 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19139), .B1(
        n19138), .B2(n18998), .ZN(n18993) );
  OAI211_X1 U21243 ( .C1(n19142), .C2(n18995), .A(n18994), .B(n18993), .ZN(
        P3_U2878) );
  AOI22_X1 U21244 ( .A1(n19066), .A2(n18997), .B1(n19144), .B2(n18996), .ZN(
        n19001) );
  AOI22_X1 U21245 ( .A1(n19146), .A2(n18999), .B1(n19149), .B2(n18998), .ZN(
        n19000) );
  OAI211_X1 U21246 ( .C1(n19002), .C2(n19147), .A(n19001), .B(n19000), .ZN(
        P3_U2870) );
  OAI22_X1 U21247 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n19050), .ZN(n19003) );
  INV_X1 U21248 ( .A(n19003), .ZN(U252) );
  INV_X1 U21249 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n19004) );
  NOR2_X1 U21250 ( .A1(n19005), .A2(n19004), .ZN(n19046) );
  INV_X1 U21251 ( .A(n19046), .ZN(n19034) );
  NAND2_X1 U21252 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19053), .ZN(n19042) );
  INV_X1 U21253 ( .A(n19042), .ZN(n19044) );
  AND2_X1 U21254 ( .A1(n19006), .A2(BUF2_REG_1__SCAN_IN), .ZN(n19043) );
  AOI22_X1 U21255 ( .A1(n19072), .A2(n19044), .B1(n19055), .B2(n19043), .ZN(
        n19009) );
  NOR2_X2 U21256 ( .A1(n19007), .A2(n19056), .ZN(n19045) );
  AOI22_X1 U21257 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19058), .B1(
        n19137), .B2(n19045), .ZN(n19008) );
  OAI211_X1 U21258 ( .C1(n19154), .C2(n19034), .A(n19009), .B(n19008), .ZN(
        P3_U2989) );
  AOI22_X1 U21259 ( .A1(n19072), .A2(n19046), .B1(n19061), .B2(n19043), .ZN(
        n19011) );
  AOI22_X1 U21260 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19062), .B1(
        n19146), .B2(n19045), .ZN(n19010) );
  OAI211_X1 U21261 ( .C1(n19070), .C2(n19042), .A(n19011), .B(n19010), .ZN(
        P3_U2981) );
  AOI22_X1 U21262 ( .A1(n19065), .A2(n19043), .B1(n19083), .B2(n19044), .ZN(
        n19013) );
  AOI22_X1 U21263 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19067), .B1(
        n19066), .B2(n19045), .ZN(n19012) );
  OAI211_X1 U21264 ( .C1(n19070), .C2(n19034), .A(n19013), .B(n19012), .ZN(
        P3_U2973) );
  AOI22_X1 U21265 ( .A1(n19083), .A2(n19046), .B1(n19071), .B2(n19043), .ZN(
        n19015) );
  AOI22_X1 U21266 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19073), .B1(
        n19072), .B2(n19045), .ZN(n19014) );
  OAI211_X1 U21267 ( .C1(n19081), .C2(n19042), .A(n19015), .B(n19014), .ZN(
        P3_U2965) );
  AOI22_X1 U21268 ( .A1(n19094), .A2(n19044), .B1(n19076), .B2(n19043), .ZN(
        n19017) );
  AOI22_X1 U21269 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19078), .B1(
        n19077), .B2(n19045), .ZN(n19016) );
  OAI211_X1 U21270 ( .C1(n19081), .C2(n19034), .A(n19017), .B(n19016), .ZN(
        P3_U2957) );
  AOI22_X1 U21271 ( .A1(n19094), .A2(n19046), .B1(n19082), .B2(n19043), .ZN(
        n19019) );
  AOI22_X1 U21272 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19084), .B1(
        n19083), .B2(n19045), .ZN(n19018) );
  OAI211_X1 U21273 ( .C1(n19022), .C2(n19042), .A(n19019), .B(n19018), .ZN(
        P3_U2949) );
  AOI22_X1 U21274 ( .A1(n19106), .A2(n19044), .B1(n19088), .B2(n19043), .ZN(
        n19021) );
  AOI22_X1 U21275 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19090), .B1(
        n19089), .B2(n19045), .ZN(n19020) );
  OAI211_X1 U21276 ( .C1(n19022), .C2(n19034), .A(n19021), .B(n19020), .ZN(
        P3_U2941) );
  AOI22_X1 U21277 ( .A1(n19112), .A2(n19044), .B1(n19093), .B2(n19043), .ZN(
        n19024) );
  AOI22_X1 U21278 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19095), .B1(
        n19094), .B2(n19045), .ZN(n19023) );
  OAI211_X1 U21279 ( .C1(n19098), .C2(n19034), .A(n19024), .B(n19023), .ZN(
        P3_U2933) );
  AOI22_X1 U21280 ( .A1(n19112), .A2(n19046), .B1(n19099), .B2(n19043), .ZN(
        n19026) );
  AOI22_X1 U21281 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19101), .B1(
        n19100), .B2(n19045), .ZN(n19025) );
  OAI211_X1 U21282 ( .C1(n19110), .C2(n19042), .A(n19026), .B(n19025), .ZN(
        P3_U2925) );
  AOI22_X1 U21283 ( .A1(n19125), .A2(n19044), .B1(n19105), .B2(n19043), .ZN(
        n19028) );
  AOI22_X1 U21284 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19107), .B1(
        n19106), .B2(n19045), .ZN(n19027) );
  OAI211_X1 U21285 ( .C1(n19110), .C2(n19034), .A(n19028), .B(n19027), .ZN(
        P3_U2917) );
  AOI22_X1 U21286 ( .A1(n19111), .A2(n19043), .B1(n19131), .B2(n19044), .ZN(
        n19030) );
  AOI22_X1 U21287 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19113), .B1(
        n19112), .B2(n19045), .ZN(n19029) );
  OAI211_X1 U21288 ( .C1(n19031), .C2(n19034), .A(n19030), .B(n19029), .ZN(
        P3_U2909) );
  AOI22_X1 U21289 ( .A1(n19138), .A2(n19044), .B1(n19116), .B2(n19043), .ZN(
        n19033) );
  AOI22_X1 U21290 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19118), .B1(
        n19117), .B2(n19045), .ZN(n19032) );
  OAI211_X1 U21291 ( .C1(n19121), .C2(n19034), .A(n19033), .B(n19032), .ZN(
        P3_U2901) );
  AOI22_X1 U21292 ( .A1(n19138), .A2(n19046), .B1(n19122), .B2(n19043), .ZN(
        n19036) );
  AOI22_X1 U21293 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19123), .B1(
        n19125), .B2(n19045), .ZN(n19035) );
  OAI211_X1 U21294 ( .C1(n19037), .C2(n19042), .A(n19036), .B(n19035), .ZN(
        P3_U2893) );
  AOI22_X1 U21295 ( .A1(n19149), .A2(n19046), .B1(n19130), .B2(n19043), .ZN(
        n19039) );
  AOI22_X1 U21296 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19132), .B1(
        n19131), .B2(n19045), .ZN(n19038) );
  OAI211_X1 U21297 ( .C1(n19135), .C2(n19042), .A(n19039), .B(n19038), .ZN(
        P3_U2885) );
  AOI22_X1 U21298 ( .A1(n19137), .A2(n19046), .B1(n19136), .B2(n19043), .ZN(
        n19041) );
  AOI22_X1 U21299 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19139), .B1(
        n19138), .B2(n19045), .ZN(n19040) );
  OAI211_X1 U21300 ( .C1(n19142), .C2(n19042), .A(n19041), .B(n19040), .ZN(
        P3_U2877) );
  AOI22_X1 U21301 ( .A1(n19066), .A2(n19044), .B1(n19144), .B2(n19043), .ZN(
        n19048) );
  AOI22_X1 U21302 ( .A1(n19146), .A2(n19046), .B1(n19149), .B2(n19045), .ZN(
        n19047) );
  OAI211_X1 U21303 ( .C1(n19049), .C2(n19147), .A(n19048), .B(n19047), .ZN(
        P3_U2869) );
  OAI22_X1 U21304 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n19050), .ZN(n19051) );
  INV_X1 U21305 ( .A(n19051), .ZN(U251) );
  INV_X1 U21306 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n19052) );
  NOR2_X1 U21307 ( .A1(n19005), .A2(n19052), .ZN(n19145) );
  INV_X1 U21308 ( .A(n19145), .ZN(n19128) );
  NAND2_X1 U21309 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19053), .ZN(n19153) );
  INV_X1 U21310 ( .A(n19153), .ZN(n19124) );
  INV_X1 U21311 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n20123) );
  NOR2_X2 U21312 ( .A1(n19054), .A2(n20123), .ZN(n19143) );
  AOI22_X1 U21313 ( .A1(n19072), .A2(n19124), .B1(n19055), .B2(n19143), .ZN(
        n19060) );
  NOR2_X2 U21314 ( .A1(n19057), .A2(n19056), .ZN(n19148) );
  AOI22_X1 U21315 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19058), .B1(
        n19137), .B2(n19148), .ZN(n19059) );
  OAI211_X1 U21316 ( .C1(n19154), .C2(n19128), .A(n19060), .B(n19059), .ZN(
        P3_U2988) );
  AOI22_X1 U21317 ( .A1(n19072), .A2(n19145), .B1(n19061), .B2(n19143), .ZN(
        n19064) );
  AOI22_X1 U21318 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19062), .B1(
        n19146), .B2(n19148), .ZN(n19063) );
  OAI211_X1 U21319 ( .C1(n19070), .C2(n19153), .A(n19064), .B(n19063), .ZN(
        P3_U2980) );
  AOI22_X1 U21320 ( .A1(n19065), .A2(n19143), .B1(n19083), .B2(n19124), .ZN(
        n19069) );
  AOI22_X1 U21321 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19067), .B1(
        n19066), .B2(n19148), .ZN(n19068) );
  OAI211_X1 U21322 ( .C1(n19070), .C2(n19128), .A(n19069), .B(n19068), .ZN(
        P3_U2972) );
  AOI22_X1 U21323 ( .A1(n19083), .A2(n19145), .B1(n19071), .B2(n19143), .ZN(
        n19075) );
  AOI22_X1 U21324 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19073), .B1(
        n19072), .B2(n19148), .ZN(n19074) );
  OAI211_X1 U21325 ( .C1(n19081), .C2(n19153), .A(n19075), .B(n19074), .ZN(
        P3_U2964) );
  AOI22_X1 U21326 ( .A1(n19094), .A2(n19124), .B1(n19076), .B2(n19143), .ZN(
        n19080) );
  AOI22_X1 U21327 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19078), .B1(
        n19077), .B2(n19148), .ZN(n19079) );
  OAI211_X1 U21328 ( .C1(n19081), .C2(n19128), .A(n19080), .B(n19079), .ZN(
        P3_U2956) );
  AOI22_X1 U21329 ( .A1(n19100), .A2(n19124), .B1(n19082), .B2(n19143), .ZN(
        n19086) );
  AOI22_X1 U21330 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19084), .B1(
        n19083), .B2(n19148), .ZN(n19085) );
  OAI211_X1 U21331 ( .C1(n19087), .C2(n19128), .A(n19086), .B(n19085), .ZN(
        P3_U2948) );
  AOI22_X1 U21332 ( .A1(n19100), .A2(n19145), .B1(n19088), .B2(n19143), .ZN(
        n19092) );
  AOI22_X1 U21333 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19090), .B1(
        n19089), .B2(n19148), .ZN(n19091) );
  OAI211_X1 U21334 ( .C1(n19098), .C2(n19153), .A(n19092), .B(n19091), .ZN(
        P3_U2940) );
  AOI22_X1 U21335 ( .A1(n19112), .A2(n19124), .B1(n19093), .B2(n19143), .ZN(
        n19097) );
  AOI22_X1 U21336 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19095), .B1(
        n19094), .B2(n19148), .ZN(n19096) );
  OAI211_X1 U21337 ( .C1(n19098), .C2(n19128), .A(n19097), .B(n19096), .ZN(
        P3_U2932) );
  AOI22_X1 U21338 ( .A1(n19117), .A2(n19124), .B1(n19099), .B2(n19143), .ZN(
        n19103) );
  AOI22_X1 U21339 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19101), .B1(
        n19100), .B2(n19148), .ZN(n19102) );
  OAI211_X1 U21340 ( .C1(n19104), .C2(n19128), .A(n19103), .B(n19102), .ZN(
        P3_U2924) );
  AOI22_X1 U21341 ( .A1(n19125), .A2(n19124), .B1(n19105), .B2(n19143), .ZN(
        n19109) );
  AOI22_X1 U21342 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19107), .B1(
        n19106), .B2(n19148), .ZN(n19108) );
  OAI211_X1 U21343 ( .C1(n19110), .C2(n19128), .A(n19109), .B(n19108), .ZN(
        P3_U2916) );
  AOI22_X1 U21344 ( .A1(n19125), .A2(n19145), .B1(n19111), .B2(n19143), .ZN(
        n19115) );
  AOI22_X1 U21345 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19113), .B1(
        n19112), .B2(n19148), .ZN(n19114) );
  OAI211_X1 U21346 ( .C1(n19121), .C2(n19153), .A(n19115), .B(n19114), .ZN(
        P3_U2908) );
  AOI22_X1 U21347 ( .A1(n19138), .A2(n19124), .B1(n19116), .B2(n19143), .ZN(
        n19120) );
  AOI22_X1 U21348 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19118), .B1(
        n19117), .B2(n19148), .ZN(n19119) );
  OAI211_X1 U21349 ( .C1(n19121), .C2(n19128), .A(n19120), .B(n19119), .ZN(
        P3_U2900) );
  AOI22_X1 U21350 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19123), .B1(
        n19122), .B2(n19143), .ZN(n19127) );
  AOI22_X1 U21351 ( .A1(n19125), .A2(n19148), .B1(n19149), .B2(n19124), .ZN(
        n19126) );
  OAI211_X1 U21352 ( .C1(n19129), .C2(n19128), .A(n19127), .B(n19126), .ZN(
        P3_U2892) );
  AOI22_X1 U21353 ( .A1(n19149), .A2(n19145), .B1(n19130), .B2(n19143), .ZN(
        n19134) );
  AOI22_X1 U21354 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19132), .B1(
        n19131), .B2(n19148), .ZN(n19133) );
  OAI211_X1 U21355 ( .C1(n19135), .C2(n19153), .A(n19134), .B(n19133), .ZN(
        P3_U2884) );
  AOI22_X1 U21356 ( .A1(n19137), .A2(n19145), .B1(n19136), .B2(n19143), .ZN(
        n19141) );
  AOI22_X1 U21357 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19139), .B1(
        n19138), .B2(n19148), .ZN(n19140) );
  OAI211_X1 U21358 ( .C1(n19142), .C2(n19153), .A(n19141), .B(n19140), .ZN(
        P3_U2876) );
  AOI22_X1 U21359 ( .A1(n19146), .A2(n19145), .B1(n19144), .B2(n19143), .ZN(
        n19152) );
  INV_X1 U21360 ( .A(n19147), .ZN(n19150) );
  AOI22_X1 U21361 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19150), .B1(
        n19149), .B2(n19148), .ZN(n19151) );
  OAI211_X1 U21362 ( .C1(n19154), .C2(n19153), .A(n19152), .B(n19151), .ZN(
        P3_U2868) );
  OAI222_X1 U21363 ( .A1(n19157), .A2(n19349), .B1(n19156), .B2(n19508), .C1(
        n19155), .C2(n19619), .ZN(P2_U2904) );
  AOI22_X1 U21364 ( .A1(n19159), .A2(n19396), .B1(n19158), .B2(n19175), .ZN(
        n19160) );
  OAI21_X1 U21365 ( .B1(n19508), .B2(n19161), .A(n19160), .ZN(P2_U2905) );
  OAI222_X1 U21366 ( .A1(n19164), .A2(n19349), .B1(n19163), .B2(n19508), .C1(
        n19619), .C2(n19162), .ZN(P2_U2906) );
  AOI22_X1 U21367 ( .A1(n19166), .A2(n19396), .B1(n19165), .B2(n19175), .ZN(
        n19167) );
  OAI21_X1 U21368 ( .B1(n19508), .B2(n19168), .A(n19167), .ZN(P2_U2907) );
  OAI222_X1 U21369 ( .A1(n19171), .A2(n19349), .B1(n19170), .B2(n19508), .C1(
        n19619), .C2(n19169), .ZN(P2_U2908) );
  AOI22_X1 U21370 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19670), .B1(n19172), 
        .B2(n19175), .ZN(n19173) );
  OAI21_X1 U21371 ( .B1(n19349), .B2(n19174), .A(n19173), .ZN(P2_U2909) );
  AOI22_X1 U21372 ( .A1(n19177), .A2(n19396), .B1(n19176), .B2(n19175), .ZN(
        n19178) );
  OAI21_X1 U21373 ( .B1(n19508), .B2(n19179), .A(n19178), .ZN(P2_U2910) );
  AOI22_X1 U21374 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19670), .B1(n19180), .B2(
        n19396), .ZN(n19181) );
  OAI21_X1 U21375 ( .B1(n19182), .B2(n19619), .A(n19181), .ZN(P2_U2911) );
  OAI222_X1 U21376 ( .A1(n19185), .A2(n19349), .B1(n19184), .B2(n19508), .C1(
        n19619), .C2(n19183), .ZN(P2_U2912) );
  OAI21_X1 U21377 ( .B1(n11835), .B2(n19687), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19186) );
  OAI21_X1 U21378 ( .B1(n19187), .B2(n19326), .A(n19186), .ZN(n19688) );
  AOI22_X1 U21379 ( .A1(n19688), .A2(n15206), .B1(n19687), .B2(n19328), .ZN(
        n19194) );
  NOR2_X1 U21380 ( .A1(n19198), .A2(n19255), .ZN(n19192) );
  INV_X1 U21381 ( .A(n11835), .ZN(n19189) );
  OAI21_X1 U21382 ( .B1(n19292), .B2(n19687), .A(n19312), .ZN(n19188) );
  OAI21_X1 U21383 ( .B1(n19189), .B2(n19297), .A(n19188), .ZN(n19190) );
  OAI21_X1 U21384 ( .B1(n19192), .B2(n19191), .A(n19190), .ZN(n19691) );
  AOI22_X1 U21385 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19691), .B1(
        n19789), .B2(n19338), .ZN(n19193) );
  OAI211_X1 U21386 ( .C1(n19341), .C2(n19699), .A(n19194), .B(n19193), .ZN(
        P2_U3175) );
  NOR2_X2 U21387 ( .A1(n19198), .A2(n19195), .ZN(n19709) );
  INV_X1 U21388 ( .A(n19709), .ZN(n19706) );
  OAI21_X1 U21389 ( .B1(n11831), .B2(n19700), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19196) );
  OAI21_X1 U21390 ( .B1(n19209), .B2(n19326), .A(n19196), .ZN(n19701) );
  AOI22_X1 U21391 ( .A1(n19701), .A2(n15206), .B1(n19328), .B2(n19700), .ZN(
        n19204) );
  OAI21_X1 U21392 ( .B1(n19198), .B2(n19197), .A(n19209), .ZN(n19202) );
  INV_X1 U21393 ( .A(n11831), .ZN(n19200) );
  OAI211_X1 U21394 ( .C1(n19200), .C2(n19297), .A(n19326), .B(n19199), .ZN(
        n19201) );
  NAND3_X1 U21395 ( .A1(n19202), .A2(n19312), .A3(n19201), .ZN(n19703) );
  AOI22_X1 U21396 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19703), .B1(
        n19702), .B2(n19338), .ZN(n19203) );
  OAI211_X1 U21397 ( .C1(n19341), .C2(n19706), .A(n19204), .B(n19203), .ZN(
        P2_U3159) );
  INV_X1 U21398 ( .A(n19205), .ZN(n19211) );
  INV_X1 U21399 ( .A(n19206), .ZN(n19208) );
  INV_X1 U21400 ( .A(n19270), .ZN(n19207) );
  NAND2_X1 U21401 ( .A1(n19208), .A2(n19207), .ZN(n19281) );
  NOR2_X1 U21402 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19209), .ZN(
        n19707) );
  OAI21_X1 U21403 ( .B1(n11812), .B2(n19707), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19210) );
  OAI21_X1 U21404 ( .B1(n19211), .B2(n19281), .A(n19210), .ZN(n19708) );
  AOI22_X1 U21405 ( .A1(n19708), .A2(n15206), .B1(n19328), .B2(n19707), .ZN(
        n19219) );
  OAI21_X1 U21406 ( .B1(n19630), .B2(n19709), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19212) );
  OAI21_X1 U21407 ( .B1(n19281), .B2(n19213), .A(n19212), .ZN(n19217) );
  OAI21_X1 U21408 ( .B1(n19295), .B2(n19707), .A(n19312), .ZN(n19214) );
  OAI21_X1 U21409 ( .B1(n19215), .B2(n19297), .A(n19214), .ZN(n19216) );
  NAND2_X1 U21410 ( .A1(n19217), .A2(n19216), .ZN(n19710) );
  AOI22_X1 U21411 ( .A1(n19710), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n19338), .B2(n19709), .ZN(n19218) );
  OAI211_X1 U21412 ( .C1(n19341), .C2(n19718), .A(n19219), .B(n19218), .ZN(
        P2_U3151) );
  NAND3_X1 U21413 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19221), .ZN(n19231) );
  NOR2_X1 U21414 ( .A1(n19263), .A2(n19231), .ZN(n19713) );
  OAI21_X1 U21415 ( .B1(n11832), .B2(n19713), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19222) );
  OAI21_X1 U21416 ( .B1(n19231), .B2(n19326), .A(n19222), .ZN(n19714) );
  AOI22_X1 U21417 ( .A1(n19714), .A2(n15206), .B1(n19328), .B2(n19713), .ZN(
        n19228) );
  OAI21_X1 U21418 ( .B1(n19453), .B2(n19293), .A(n19231), .ZN(n19226) );
  INV_X1 U21419 ( .A(n11832), .ZN(n19224) );
  OAI21_X1 U21420 ( .B1(n19292), .B2(n19713), .A(n19312), .ZN(n19223) );
  OAI21_X1 U21421 ( .B1(n19224), .B2(n19297), .A(n19223), .ZN(n19225) );
  NAND2_X1 U21422 ( .A1(n19226), .A2(n19225), .ZN(n19715) );
  AOI22_X1 U21423 ( .A1(n19338), .A2(n19630), .B1(
        P2_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n19715), .ZN(n19227) );
  OAI211_X1 U21424 ( .C1(n19341), .C2(n19633), .A(n19228), .B(n19227), .ZN(
        P2_U3143) );
  AOI21_X1 U21425 ( .B1(n19229), .B2(n19633), .A(n21607), .ZN(n19230) );
  NOR2_X1 U21426 ( .A1(n19230), .A2(n19326), .ZN(n19235) );
  NOR2_X1 U21427 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19231), .ZN(
        n19719) );
  NOR2_X1 U21428 ( .A1(n19719), .A2(n19726), .ZN(n19237) );
  AOI211_X1 U21429 ( .C1(n19232), .C2(n19233), .A(n19295), .B(n19719), .ZN(
        n19234) );
  AOI22_X1 U21430 ( .A1(n19319), .A2(n19727), .B1(n19328), .B2(n19719), .ZN(
        n19240) );
  INV_X1 U21431 ( .A(n19235), .ZN(n19238) );
  OAI21_X1 U21432 ( .B1(n19232), .B2(n19719), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19236) );
  AOI22_X1 U21433 ( .A1(n15206), .A2(n19721), .B1(n19720), .B2(n19338), .ZN(
        n19239) );
  OAI211_X1 U21434 ( .C1(n19725), .C2(n19241), .A(n19240), .B(n19239), .ZN(
        P2_U3135) );
  NOR2_X1 U21435 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19242), .ZN(
        n19733) );
  AOI22_X1 U21436 ( .A1(n19338), .A2(n19734), .B1(n19328), .B2(n19733), .ZN(
        n19252) );
  OAI21_X1 U21437 ( .B1(n19734), .B2(n19742), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19243) );
  NAND2_X1 U21438 ( .A1(n19243), .A2(n19295), .ZN(n19250) );
  NOR2_X1 U21439 ( .A1(n19291), .A2(n19266), .ZN(n19740) );
  NOR2_X1 U21440 ( .A1(n19250), .A2(n19740), .ZN(n19244) );
  AOI211_X1 U21441 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19245), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19244), .ZN(n19246) );
  OAI21_X1 U21442 ( .B1(n19733), .B2(n19246), .A(n19312), .ZN(n19736) );
  NOR2_X1 U21443 ( .A1(n19740), .A2(n19733), .ZN(n19249) );
  OAI21_X1 U21444 ( .B1(n19247), .B2(n19733), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19248) );
  AOI22_X1 U21445 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19736), .B1(
        n19735), .B2(n15206), .ZN(n19251) );
  OAI211_X1 U21446 ( .C1(n19341), .C2(n19739), .A(n19252), .B(n19251), .ZN(
        P2_U3119) );
  NAND2_X1 U21447 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19269), .ZN(
        n19254) );
  OAI21_X1 U21448 ( .B1(n11834), .B2(n19740), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19253) );
  OAI21_X1 U21449 ( .B1(n19254), .B2(n19326), .A(n19253), .ZN(n19741) );
  AOI22_X1 U21450 ( .A1(n19741), .A2(n15206), .B1(n19328), .B2(n19740), .ZN(
        n19262) );
  OAI22_X1 U21451 ( .A1(n19256), .A2(n19255), .B1(n19266), .B2(n19294), .ZN(
        n19260) );
  INV_X1 U21452 ( .A(n11834), .ZN(n19258) );
  INV_X1 U21453 ( .A(n19740), .ZN(n19257) );
  OAI211_X1 U21454 ( .C1(n19258), .C2(n19297), .A(n19326), .B(n19257), .ZN(
        n19259) );
  NAND3_X1 U21455 ( .A1(n19260), .A2(n19312), .A3(n19259), .ZN(n19743) );
  AOI22_X1 U21456 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19743), .B1(
        n19742), .B2(n19338), .ZN(n19261) );
  OAI211_X1 U21457 ( .C1(n19341), .C2(n19752), .A(n19262), .B(n19261), .ZN(
        P2_U3111) );
  NAND2_X1 U21458 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19263), .ZN(
        n19311) );
  NOR2_X1 U21459 ( .A1(n19311), .A2(n19266), .ZN(n19746) );
  OAI21_X1 U21460 ( .B1(n19264), .B2(n19746), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19265) );
  OAI21_X1 U21461 ( .B1(n19318), .B2(n19266), .A(n19265), .ZN(n19747) );
  AOI22_X1 U21462 ( .A1(n19747), .A2(n15206), .B1(n19328), .B2(n19746), .ZN(
        n19275) );
  OAI21_X1 U21463 ( .B1(n19295), .B2(n19746), .A(n19312), .ZN(n19267) );
  OAI21_X1 U21464 ( .B1(n19268), .B2(n19297), .A(n19267), .ZN(n19273) );
  NAND2_X1 U21465 ( .A1(n19270), .A2(n19269), .ZN(n19271) );
  OAI221_X1 U21466 ( .B1(n21607), .B2(n19758), .C1(n21607), .C2(n19752), .A(
        n19271), .ZN(n19272) );
  AOI22_X1 U21467 ( .A1(n19338), .A2(n19645), .B1(
        P2_INSTQUEUE_REG_6__7__SCAN_IN), .B2(n19748), .ZN(n19274) );
  OAI211_X1 U21468 ( .C1(n19341), .C2(n19758), .A(n19275), .B(n19274), .ZN(
        P2_U3103) );
  INV_X1 U21469 ( .A(n19308), .ZN(n19278) );
  INV_X1 U21470 ( .A(n19276), .ZN(n19277) );
  NOR2_X1 U21471 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19279), .ZN(
        n19759) );
  AOI22_X1 U21472 ( .A1(n19338), .A2(n19760), .B1(n19328), .B2(n19759), .ZN(
        n19289) );
  OAI21_X1 U21473 ( .B1(n19760), .B2(n19653), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19280) );
  NAND2_X1 U21474 ( .A1(n19280), .A2(n19295), .ZN(n19287) );
  NOR2_X1 U21475 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19281), .ZN(
        n19284) );
  OAI21_X1 U21476 ( .B1(n19295), .B2(n19759), .A(n19312), .ZN(n19282) );
  OAI21_X1 U21477 ( .B1(n11825), .B2(n19297), .A(n19282), .ZN(n19283) );
  INV_X1 U21478 ( .A(n19284), .ZN(n19286) );
  OAI21_X1 U21479 ( .B1(n11813), .B2(n19759), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19285) );
  AOI22_X1 U21480 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19762), .B1(
        n15206), .B2(n19761), .ZN(n19288) );
  OAI211_X1 U21481 ( .C1(n19341), .C2(n19770), .A(n19289), .B(n19288), .ZN(
        P2_U3087) );
  NOR2_X2 U21482 ( .A1(n19308), .A2(n19290), .ZN(n19774) );
  INV_X1 U21483 ( .A(n19774), .ZN(n19656) );
  NOR2_X1 U21484 ( .A1(n19291), .A2(n19323), .ZN(n19765) );
  AOI22_X1 U21485 ( .A1(n19338), .A2(n19653), .B1(n19328), .B2(n19765), .ZN(
        n19306) );
  OAI21_X1 U21486 ( .B1(n19330), .B2(n19293), .A(n19292), .ZN(n19304) );
  NOR2_X1 U21487 ( .A1(n19294), .A2(n19323), .ZN(n19300) );
  INV_X1 U21488 ( .A(n19301), .ZN(n19298) );
  OAI21_X1 U21489 ( .B1(n19295), .B2(n19765), .A(n19312), .ZN(n19296) );
  OAI21_X1 U21490 ( .B1(n19298), .B2(n19297), .A(n19296), .ZN(n19299) );
  OAI21_X1 U21491 ( .B1(n19304), .B2(n19300), .A(n19299), .ZN(n19767) );
  INV_X1 U21492 ( .A(n19300), .ZN(n19303) );
  OAI21_X1 U21493 ( .B1(n19301), .B2(n19765), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19302) );
  OAI21_X1 U21494 ( .B1(n19304), .B2(n19303), .A(n19302), .ZN(n19766) );
  AOI22_X1 U21495 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19767), .B1(
        n15206), .B2(n19766), .ZN(n19305) );
  OAI211_X1 U21496 ( .C1(n19341), .C2(n19656), .A(n19306), .B(n19305), .ZN(
        P2_U3079) );
  NOR2_X2 U21497 ( .A1(n19308), .A2(n19307), .ZN(n19781) );
  NOR2_X1 U21498 ( .A1(n19318), .A2(n19323), .ZN(n19309) );
  AOI221_X1 U21499 ( .B1(n19781), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19774), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19309), .ZN(n19315) );
  NOR2_X1 U21500 ( .A1(n19310), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19313) );
  NOR2_X1 U21501 ( .A1(n19311), .A2(n19323), .ZN(n19772) );
  OAI211_X1 U21502 ( .C1(n19313), .C2(n19772), .A(n19326), .B(n19312), .ZN(
        n19314) );
  OAI21_X1 U21503 ( .B1(n19316), .B2(n19772), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19317) );
  OAI21_X1 U21504 ( .B1(n19323), .B2(n19318), .A(n19317), .ZN(n19773) );
  AOI22_X1 U21505 ( .A1(n19773), .A2(n15206), .B1(n19328), .B2(n19772), .ZN(
        n19321) );
  AOI22_X1 U21506 ( .A1(n19774), .A2(n19338), .B1(n19781), .B2(n19319), .ZN(
        n19320) );
  OAI211_X1 U21507 ( .C1(n19778), .C2(n19322), .A(n19321), .B(n19320), .ZN(
        P2_U3071) );
  NOR2_X1 U21508 ( .A1(n19324), .A2(n19323), .ZN(n19779) );
  OAI21_X1 U21509 ( .B1(n11830), .B2(n19779), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19325) );
  OAI21_X1 U21510 ( .B1(n19327), .B2(n19326), .A(n19325), .ZN(n19780) );
  AOI22_X1 U21511 ( .A1(n19780), .A2(n15206), .B1(n19328), .B2(n19779), .ZN(
        n19340) );
  NOR2_X1 U21512 ( .A1(n19330), .A2(n19329), .ZN(n19337) );
  INV_X1 U21513 ( .A(n19779), .ZN(n19334) );
  NAND2_X1 U21514 ( .A1(n11830), .A2(n19331), .ZN(n19333) );
  OAI211_X1 U21515 ( .C1(n19683), .C2(n19334), .A(n19333), .B(n19332), .ZN(
        n19335) );
  OAI21_X1 U21516 ( .B1(n19337), .B2(n19336), .A(n19335), .ZN(n19782) );
  AOI22_X1 U21517 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19782), .B1(
        n19781), .B2(n19338), .ZN(n19339) );
  OAI211_X1 U21518 ( .C1(n19341), .C2(n19785), .A(n19340), .B(n19339), .ZN(
        P2_U3063) );
  AOI22_X1 U21519 ( .A1(n19672), .A2(n19342), .B1(P2_EAX_REG_22__SCAN_IN), 
        .B2(n19670), .ZN(n19347) );
  AOI22_X1 U21520 ( .A1(n19674), .A2(BUF2_REG_22__SCAN_IN), .B1(n19673), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n19346) );
  AOI22_X1 U21521 ( .A1(n19344), .A2(n19561), .B1(n19612), .B2(n19343), .ZN(
        n19345) );
  NAND3_X1 U21522 ( .A1(n19347), .A2(n19346), .A3(n19345), .ZN(P2_U2897) );
  OAI222_X1 U21523 ( .A1(n19350), .A2(n19349), .B1(n19348), .B2(n19508), .C1(
        n19619), .C2(n19351), .ZN(P2_U2913) );
  AOI22_X1 U21524 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n19689), .B1(
        BUF1_REG_30__SCAN_IN), .B2(n19690), .ZN(n19386) );
  NOR2_X2 U21525 ( .A1(n11684), .A2(n19685), .ZN(n19387) );
  AOI22_X1 U21526 ( .A1(n19688), .A2(n19352), .B1(n19687), .B2(n19387), .ZN(
        n19354) );
  AOI22_X1 U21527 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19690), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19689), .ZN(n19381) );
  AOI22_X1 U21528 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19691), .B1(
        n19789), .B2(n19389), .ZN(n19353) );
  OAI211_X1 U21529 ( .C1(n19386), .C2(n19699), .A(n19354), .B(n19353), .ZN(
        P2_U3174) );
  AOI22_X1 U21530 ( .A1(n19566), .A2(n19389), .B1(n19694), .B2(n19387), .ZN(
        n19356) );
  AOI22_X1 U21531 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19696), .B1(
        n19352), .B2(n19695), .ZN(n19355) );
  OAI211_X1 U21532 ( .C1(n19386), .C2(n19574), .A(n19356), .B(n19355), .ZN(
        P2_U3166) );
  AOI22_X1 U21533 ( .A1(n19701), .A2(n19352), .B1(n19387), .B2(n19700), .ZN(
        n19358) );
  INV_X1 U21534 ( .A(n19386), .ZN(n19388) );
  AOI22_X1 U21535 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19703), .B1(
        n19709), .B2(n19388), .ZN(n19357) );
  OAI211_X1 U21536 ( .C1(n19381), .C2(n19574), .A(n19358), .B(n19357), .ZN(
        P2_U3158) );
  AOI22_X1 U21537 ( .A1(n19708), .A2(n19352), .B1(n19387), .B2(n19707), .ZN(
        n19360) );
  AOI22_X1 U21538 ( .A1(n19710), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n19709), .B2(n19389), .ZN(n19359) );
  OAI211_X1 U21539 ( .C1(n19386), .C2(n19718), .A(n19360), .B(n19359), .ZN(
        P2_U3150) );
  AOI22_X1 U21540 ( .A1(n19714), .A2(n19352), .B1(n19387), .B2(n19713), .ZN(
        n19362) );
  AOI22_X1 U21541 ( .A1(n19630), .A2(n19389), .B1(
        P2_INSTQUEUE_REG_11__6__SCAN_IN), .B2(n19715), .ZN(n19361) );
  OAI211_X1 U21542 ( .C1(n19386), .C2(n19633), .A(n19362), .B(n19361), .ZN(
        P2_U3142) );
  AOI22_X1 U21543 ( .A1(n19388), .A2(n19727), .B1(n19387), .B2(n19719), .ZN(
        n19364) );
  AOI22_X1 U21544 ( .A1(n19352), .A2(n19721), .B1(n19720), .B2(n19389), .ZN(
        n19363) );
  OAI211_X1 U21545 ( .C1(n19725), .C2(n11893), .A(n19364), .B(n19363), .ZN(
        P2_U3134) );
  INV_X1 U21546 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n19367) );
  AOI22_X1 U21547 ( .A1(n19388), .A2(n19734), .B1(n19726), .B2(n19387), .ZN(
        n19366) );
  AOI22_X1 U21548 ( .A1(n19352), .A2(n19728), .B1(n19727), .B2(n19389), .ZN(
        n19365) );
  OAI211_X1 U21549 ( .C1(n19732), .C2(n19367), .A(n19366), .B(n19365), .ZN(
        P2_U3126) );
  AOI22_X1 U21550 ( .A1(n19734), .A2(n19389), .B1(n19387), .B2(n19733), .ZN(
        n19369) );
  AOI22_X1 U21551 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19736), .B1(
        n19735), .B2(n19352), .ZN(n19368) );
  OAI211_X1 U21552 ( .C1(n19386), .C2(n19739), .A(n19369), .B(n19368), .ZN(
        P2_U3118) );
  AOI22_X1 U21553 ( .A1(n19741), .A2(n19352), .B1(n19740), .B2(n19387), .ZN(
        n19371) );
  AOI22_X1 U21554 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19743), .B1(
        n19742), .B2(n19389), .ZN(n19370) );
  OAI211_X1 U21555 ( .C1(n19386), .C2(n19752), .A(n19371), .B(n19370), .ZN(
        P2_U3110) );
  AOI22_X1 U21556 ( .A1(n19747), .A2(n19352), .B1(n19387), .B2(n19746), .ZN(
        n19373) );
  AOI22_X1 U21557 ( .A1(n19645), .A2(n19389), .B1(
        P2_INSTQUEUE_REG_6__6__SCAN_IN), .B2(n19748), .ZN(n19372) );
  OAI211_X1 U21558 ( .C1(n19386), .C2(n19758), .A(n19373), .B(n19372), .ZN(
        P2_U3102) );
  AOI22_X1 U21559 ( .A1(n19388), .A2(n19760), .B1(n19753), .B2(n19387), .ZN(
        n19375) );
  AOI22_X1 U21560 ( .A1(n19352), .A2(n19754), .B1(n19749), .B2(n19389), .ZN(
        n19374) );
  OAI211_X1 U21561 ( .C1(n19376), .C2(n11541), .A(n19375), .B(n19374), .ZN(
        P2_U3094) );
  AOI22_X1 U21562 ( .A1(n19760), .A2(n19389), .B1(n19759), .B2(n19387), .ZN(
        n19378) );
  AOI22_X1 U21563 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19762), .B1(
        n19352), .B2(n19761), .ZN(n19377) );
  OAI211_X1 U21564 ( .C1(n19386), .C2(n19770), .A(n19378), .B(n19377), .ZN(
        P2_U3086) );
  AOI22_X1 U21565 ( .A1(n19388), .A2(n19774), .B1(n19765), .B2(n19387), .ZN(
        n19380) );
  AOI22_X1 U21566 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19767), .B1(
        n19352), .B2(n19766), .ZN(n19379) );
  OAI211_X1 U21567 ( .C1(n19381), .C2(n19770), .A(n19380), .B(n19379), .ZN(
        P2_U3078) );
  AOI22_X1 U21568 ( .A1(n19773), .A2(n19352), .B1(n19387), .B2(n19772), .ZN(
        n19383) );
  AOI22_X1 U21569 ( .A1(n19774), .A2(n19389), .B1(n19781), .B2(n19388), .ZN(
        n19382) );
  OAI211_X1 U21570 ( .C1(n19778), .C2(n14186), .A(n19383), .B(n19382), .ZN(
        P2_U3070) );
  AOI22_X1 U21571 ( .A1(n19780), .A2(n19352), .B1(n19387), .B2(n19779), .ZN(
        n19385) );
  AOI22_X1 U21572 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19782), .B1(
        n19781), .B2(n19389), .ZN(n19384) );
  OAI211_X1 U21573 ( .C1(n19386), .C2(n19785), .A(n19385), .B(n19384), .ZN(
        P2_U3062) );
  AOI22_X1 U21574 ( .A1(n19388), .A2(n19789), .B1(n19788), .B2(n19387), .ZN(
        n19391) );
  AOI22_X1 U21575 ( .A1(n19794), .A2(n19389), .B1(n19792), .B2(n19352), .ZN(
        n19390) );
  OAI211_X1 U21576 ( .C1(n19798), .C2(n19392), .A(n19391), .B(n19390), .ZN(
        P2_U3054) );
  INV_X1 U21577 ( .A(n19454), .ZN(n19446) );
  NAND2_X1 U21578 ( .A1(n19393), .A2(n19446), .ZN(n19456) );
  OAI21_X1 U21579 ( .B1(n19456), .B2(n19677), .A(n19394), .ZN(n19395) );
  AOI22_X1 U21580 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19670), .B1(n19396), .B2(
        n19395), .ZN(n19397) );
  OAI21_X1 U21581 ( .B1(n19398), .B2(n19619), .A(n19397), .ZN(P2_U2914) );
  AOI22_X1 U21582 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19690), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19689), .ZN(n19428) );
  NOR2_X2 U21583 ( .A1(n19400), .A2(n19685), .ZN(n19434) );
  AOI22_X1 U21584 ( .A1(n19688), .A2(n19399), .B1(n19687), .B2(n19434), .ZN(
        n19402) );
  AOI22_X1 U21585 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19690), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19689), .ZN(n19433) );
  AOI22_X1 U21586 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19691), .B1(
        n19566), .B2(n19435), .ZN(n19401) );
  OAI211_X1 U21587 ( .C1(n19428), .C2(n19569), .A(n19402), .B(n19401), .ZN(
        P2_U3173) );
  AOI22_X1 U21588 ( .A1(n19435), .A2(n19702), .B1(n19694), .B2(n19434), .ZN(
        n19404) );
  AOI22_X1 U21589 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19696), .B1(
        n19399), .B2(n19695), .ZN(n19403) );
  OAI211_X1 U21590 ( .C1(n19428), .C2(n19699), .A(n19404), .B(n19403), .ZN(
        P2_U3165) );
  AOI22_X1 U21591 ( .A1(n19701), .A2(n19399), .B1(n19434), .B2(n19700), .ZN(
        n19406) );
  AOI22_X1 U21592 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19703), .B1(
        n19709), .B2(n19435), .ZN(n19405) );
  OAI211_X1 U21593 ( .C1(n19428), .C2(n19574), .A(n19406), .B(n19405), .ZN(
        P2_U3157) );
  AOI22_X1 U21594 ( .A1(n19708), .A2(n19399), .B1(n19434), .B2(n19707), .ZN(
        n19408) );
  AOI22_X1 U21595 ( .A1(n19710), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n19709), .B2(n19436), .ZN(n19407) );
  OAI211_X1 U21596 ( .C1(n19433), .C2(n19718), .A(n19408), .B(n19407), .ZN(
        P2_U3149) );
  AOI22_X1 U21597 ( .A1(n19714), .A2(n19399), .B1(n19434), .B2(n19713), .ZN(
        n19410) );
  AOI22_X1 U21598 ( .A1(n19630), .A2(n19436), .B1(
        P2_INSTQUEUE_REG_11__5__SCAN_IN), .B2(n19715), .ZN(n19409) );
  OAI211_X1 U21599 ( .C1(n19433), .C2(n19633), .A(n19410), .B(n19409), .ZN(
        P2_U3141) );
  AOI22_X1 U21600 ( .A1(n19720), .A2(n19436), .B1(n19434), .B2(n19719), .ZN(
        n19412) );
  AOI22_X1 U21601 ( .A1(n19399), .A2(n19721), .B1(n19727), .B2(n19435), .ZN(
        n19411) );
  OAI211_X1 U21602 ( .C1(n19725), .C2(n11843), .A(n19412), .B(n19411), .ZN(
        P2_U3133) );
  INV_X1 U21603 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n19415) );
  AOI22_X1 U21604 ( .A1(n19435), .A2(n19734), .B1(n19726), .B2(n19434), .ZN(
        n19414) );
  AOI22_X1 U21605 ( .A1(n19399), .A2(n19728), .B1(n19727), .B2(n19436), .ZN(
        n19413) );
  OAI211_X1 U21606 ( .C1(n19732), .C2(n19415), .A(n19414), .B(n19413), .ZN(
        P2_U3125) );
  AOI22_X1 U21607 ( .A1(n19734), .A2(n19436), .B1(n19434), .B2(n19733), .ZN(
        n19417) );
  AOI22_X1 U21608 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19736), .B1(
        n19735), .B2(n19399), .ZN(n19416) );
  OAI211_X1 U21609 ( .C1(n19433), .C2(n19739), .A(n19417), .B(n19416), .ZN(
        P2_U3117) );
  AOI22_X1 U21610 ( .A1(n19741), .A2(n19399), .B1(n19740), .B2(n19434), .ZN(
        n19419) );
  AOI22_X1 U21611 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19743), .B1(
        n19742), .B2(n19436), .ZN(n19418) );
  OAI211_X1 U21612 ( .C1(n19433), .C2(n19752), .A(n19419), .B(n19418), .ZN(
        P2_U3109) );
  AOI22_X1 U21613 ( .A1(n19747), .A2(n19399), .B1(n19434), .B2(n19746), .ZN(
        n19421) );
  AOI22_X1 U21614 ( .A1(n19435), .A2(n19749), .B1(
        P2_INSTQUEUE_REG_6__5__SCAN_IN), .B2(n19748), .ZN(n19420) );
  OAI211_X1 U21615 ( .C1(n19428), .C2(n19752), .A(n19421), .B(n19420), .ZN(
        P2_U3101) );
  AOI22_X1 U21616 ( .A1(n19436), .A2(n19749), .B1(n19753), .B2(n19434), .ZN(
        n19423) );
  AOI22_X1 U21617 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19755), .B1(
        n19399), .B2(n19754), .ZN(n19422) );
  OAI211_X1 U21618 ( .C1(n19433), .C2(n19650), .A(n19423), .B(n19422), .ZN(
        P2_U3093) );
  AOI22_X1 U21619 ( .A1(n19760), .A2(n19436), .B1(n19759), .B2(n19434), .ZN(
        n19425) );
  AOI22_X1 U21620 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19762), .B1(
        n19399), .B2(n19761), .ZN(n19424) );
  OAI211_X1 U21621 ( .C1(n19433), .C2(n19770), .A(n19425), .B(n19424), .ZN(
        P2_U3085) );
  AOI22_X1 U21622 ( .A1(n19435), .A2(n19774), .B1(n19765), .B2(n19434), .ZN(
        n19427) );
  AOI22_X1 U21623 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19767), .B1(
        n19399), .B2(n19766), .ZN(n19426) );
  OAI211_X1 U21624 ( .C1(n19428), .C2(n19770), .A(n19427), .B(n19426), .ZN(
        P2_U3077) );
  AOI22_X1 U21625 ( .A1(n19773), .A2(n19399), .B1(n19434), .B2(n19772), .ZN(
        n19430) );
  AOI22_X1 U21626 ( .A1(n19774), .A2(n19436), .B1(n19781), .B2(n19435), .ZN(
        n19429) );
  OAI211_X1 U21627 ( .C1(n19778), .C2(n14177), .A(n19430), .B(n19429), .ZN(
        P2_U3069) );
  AOI22_X1 U21628 ( .A1(n19780), .A2(n19399), .B1(n19434), .B2(n19779), .ZN(
        n19432) );
  AOI22_X1 U21629 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19782), .B1(
        n19781), .B2(n19436), .ZN(n19431) );
  OAI211_X1 U21630 ( .C1(n19433), .C2(n19785), .A(n19432), .B(n19431), .ZN(
        P2_U3061) );
  AOI22_X1 U21631 ( .A1(n19435), .A2(n19789), .B1(n19788), .B2(n19434), .ZN(
        n19438) );
  AOI22_X1 U21632 ( .A1(n19794), .A2(n19436), .B1(n19792), .B2(n19399), .ZN(
        n19437) );
  OAI211_X1 U21633 ( .C1(n19798), .C2(n14932), .A(n19438), .B(n19437), .ZN(
        P2_U3053) );
  AOI22_X1 U21634 ( .A1(n19672), .A2(n19439), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n19670), .ZN(n19445) );
  AOI22_X1 U21635 ( .A1(n19674), .A2(BUF2_REG_20__SCAN_IN), .B1(n19673), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n19444) );
  OAI22_X1 U21636 ( .A1(n19441), .A2(n19677), .B1(n19676), .B2(n19440), .ZN(
        n19442) );
  INV_X1 U21637 ( .A(n19442), .ZN(n19443) );
  NAND3_X1 U21638 ( .A1(n19445), .A2(n19444), .A3(n19443), .ZN(P2_U2899) );
  AOI22_X1 U21639 ( .A1(n19612), .A2(n19446), .B1(n19670), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n19460) );
  XNOR2_X1 U21640 ( .A(n19447), .B(n19611), .ZN(n19615) );
  NOR2_X1 U21641 ( .A1(n19615), .A2(n19614), .ZN(n19613) );
  AOI21_X1 U21642 ( .B1(n19449), .B2(n19448), .A(n19613), .ZN(n19450) );
  XNOR2_X1 U21643 ( .A(n19450), .B(n19558), .ZN(n19560) );
  NAND2_X1 U21644 ( .A1(n19450), .A2(n19558), .ZN(n19451) );
  OAI21_X1 U21645 ( .B1(n19560), .B2(n19452), .A(n19451), .ZN(n19512) );
  XNOR2_X1 U21646 ( .A(n19453), .B(n19509), .ZN(n19513) );
  NOR2_X1 U21647 ( .A1(n19512), .A2(n19513), .ZN(n19511) );
  AOI21_X1 U21648 ( .B1(n19509), .B2(n19453), .A(n19511), .ZN(n19458) );
  NAND2_X1 U21649 ( .A1(n19455), .A2(n19454), .ZN(n19457) );
  OAI211_X1 U21650 ( .C1(n19458), .C2(n19457), .A(n19456), .B(n19561), .ZN(
        n19459) );
  OAI211_X1 U21651 ( .C1(n19461), .C2(n19619), .A(n19460), .B(n19459), .ZN(
        P2_U2915) );
  NOR2_X2 U21652 ( .A1(n19461), .A2(n19683), .ZN(n19503) );
  NOR2_X2 U21653 ( .A1(n11331), .A2(n19685), .ZN(n19501) );
  AOI22_X1 U21654 ( .A1(n19688), .A2(n19503), .B1(n19687), .B2(n19501), .ZN(
        n19466) );
  OAI22_X2 U21655 ( .A1(n20066), .A2(n19464), .B1(n19463), .B2(n19462), .ZN(
        n19504) );
  AOI22_X1 U21656 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19691), .B1(
        n19789), .B2(n19504), .ZN(n19465) );
  OAI211_X1 U21657 ( .C1(n19500), .C2(n19699), .A(n19466), .B(n19465), .ZN(
        P2_U3172) );
  INV_X1 U21658 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n19470) );
  AOI22_X1 U21659 ( .A1(n19504), .A2(n19566), .B1(n19694), .B2(n19501), .ZN(
        n19468) );
  INV_X1 U21660 ( .A(n19500), .ZN(n19502) );
  AOI22_X1 U21661 ( .A1(n19503), .A2(n19695), .B1(n19702), .B2(n19502), .ZN(
        n19467) );
  OAI211_X1 U21662 ( .C1(n19470), .C2(n19469), .A(n19468), .B(n19467), .ZN(
        P2_U3164) );
  AOI22_X1 U21663 ( .A1(n19701), .A2(n19503), .B1(n19501), .B2(n19700), .ZN(
        n19472) );
  AOI22_X1 U21664 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19703), .B1(
        n19702), .B2(n19504), .ZN(n19471) );
  OAI211_X1 U21665 ( .C1(n19500), .C2(n19706), .A(n19472), .B(n19471), .ZN(
        P2_U3156) );
  AOI22_X1 U21666 ( .A1(n19708), .A2(n19503), .B1(n19501), .B2(n19707), .ZN(
        n19474) );
  AOI22_X1 U21667 ( .A1(n19710), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n19709), .B2(n19504), .ZN(n19473) );
  OAI211_X1 U21668 ( .C1(n19500), .C2(n19718), .A(n19474), .B(n19473), .ZN(
        P2_U3148) );
  AOI22_X1 U21669 ( .A1(n19714), .A2(n19503), .B1(n19501), .B2(n19713), .ZN(
        n19476) );
  AOI22_X1 U21670 ( .A1(n19504), .A2(n19630), .B1(
        P2_INSTQUEUE_REG_11__4__SCAN_IN), .B2(n19715), .ZN(n19475) );
  OAI211_X1 U21671 ( .C1(n19500), .C2(n19633), .A(n19476), .B(n19475), .ZN(
        P2_U3140) );
  INV_X1 U21672 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n19479) );
  AOI22_X1 U21673 ( .A1(n19502), .A2(n19727), .B1(n19501), .B2(n19719), .ZN(
        n19478) );
  AOI22_X1 U21674 ( .A1(n19503), .A2(n19721), .B1(n19720), .B2(n19504), .ZN(
        n19477) );
  OAI211_X1 U21675 ( .C1(n19725), .C2(n19479), .A(n19478), .B(n19477), .ZN(
        P2_U3132) );
  INV_X1 U21676 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n19482) );
  AOI22_X1 U21677 ( .A1(n19504), .A2(n19727), .B1(n19726), .B2(n19501), .ZN(
        n19481) );
  AOI22_X1 U21678 ( .A1(n19734), .A2(n19502), .B1(n19503), .B2(n19728), .ZN(
        n19480) );
  OAI211_X1 U21679 ( .C1(n19732), .C2(n19482), .A(n19481), .B(n19480), .ZN(
        P2_U3124) );
  AOI22_X1 U21680 ( .A1(n19504), .A2(n19734), .B1(n19501), .B2(n19733), .ZN(
        n19484) );
  AOI22_X1 U21681 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19736), .B1(
        n19735), .B2(n19503), .ZN(n19483) );
  OAI211_X1 U21682 ( .C1(n19500), .C2(n19739), .A(n19484), .B(n19483), .ZN(
        P2_U3116) );
  AOI22_X1 U21683 ( .A1(n19741), .A2(n19503), .B1(n19740), .B2(n19501), .ZN(
        n19486) );
  AOI22_X1 U21684 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19743), .B1(
        n19742), .B2(n19504), .ZN(n19485) );
  OAI211_X1 U21685 ( .C1(n19500), .C2(n19752), .A(n19486), .B(n19485), .ZN(
        P2_U3108) );
  AOI22_X1 U21686 ( .A1(n19747), .A2(n19503), .B1(n19501), .B2(n19746), .ZN(
        n19488) );
  AOI22_X1 U21687 ( .A1(n19504), .A2(n19645), .B1(
        P2_INSTQUEUE_REG_6__4__SCAN_IN), .B2(n19748), .ZN(n19487) );
  OAI211_X1 U21688 ( .C1(n19500), .C2(n19758), .A(n19488), .B(n19487), .ZN(
        P2_U3100) );
  AOI22_X1 U21689 ( .A1(n19504), .A2(n19749), .B1(n19753), .B2(n19501), .ZN(
        n19490) );
  AOI22_X1 U21690 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19755), .B1(
        n19503), .B2(n19754), .ZN(n19489) );
  OAI211_X1 U21691 ( .C1(n19500), .C2(n19650), .A(n19490), .B(n19489), .ZN(
        P2_U3092) );
  AOI22_X1 U21692 ( .A1(n19504), .A2(n19760), .B1(n19501), .B2(n19759), .ZN(
        n19492) );
  AOI22_X1 U21693 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19762), .B1(
        n19503), .B2(n19761), .ZN(n19491) );
  OAI211_X1 U21694 ( .C1(n19500), .C2(n19770), .A(n19492), .B(n19491), .ZN(
        P2_U3084) );
  AOI22_X1 U21695 ( .A1(n19504), .A2(n19653), .B1(n19765), .B2(n19501), .ZN(
        n19494) );
  AOI22_X1 U21696 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19767), .B1(
        n19503), .B2(n19766), .ZN(n19493) );
  OAI211_X1 U21697 ( .C1(n19500), .C2(n19656), .A(n19494), .B(n19493), .ZN(
        P2_U3076) );
  INV_X1 U21698 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n19497) );
  AOI22_X1 U21699 ( .A1(n19773), .A2(n19503), .B1(n19501), .B2(n19772), .ZN(
        n19496) );
  AOI22_X1 U21700 ( .A1(n19774), .A2(n19504), .B1(n19781), .B2(n19502), .ZN(
        n19495) );
  OAI211_X1 U21701 ( .C1(n19778), .C2(n19497), .A(n19496), .B(n19495), .ZN(
        P2_U3068) );
  AOI22_X1 U21702 ( .A1(n19780), .A2(n19503), .B1(n19501), .B2(n19779), .ZN(
        n19499) );
  AOI22_X1 U21703 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19782), .B1(
        n19781), .B2(n19504), .ZN(n19498) );
  OAI211_X1 U21704 ( .C1(n19500), .C2(n19785), .A(n19499), .B(n19498), .ZN(
        P2_U3060) );
  INV_X1 U21705 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n19507) );
  AOI22_X1 U21706 ( .A1(n19502), .A2(n19789), .B1(n19788), .B2(n19501), .ZN(
        n19506) );
  AOI22_X1 U21707 ( .A1(n19794), .A2(n19504), .B1(n19792), .B2(n19503), .ZN(
        n19505) );
  OAI211_X1 U21708 ( .C1(n19798), .C2(n19507), .A(n19506), .B(n19505), .ZN(
        P2_U3052) );
  OAI22_X1 U21709 ( .A1(n19509), .A2(n19676), .B1(n19508), .B2(n17302), .ZN(
        n19510) );
  INV_X1 U21710 ( .A(n19510), .ZN(n19516) );
  AOI21_X1 U21711 ( .B1(n19513), .B2(n19512), .A(n19511), .ZN(n19514) );
  OR2_X1 U21712 ( .A1(n19514), .A2(n19677), .ZN(n19515) );
  OAI211_X1 U21713 ( .C1(n19517), .C2(n19619), .A(n19516), .B(n19515), .ZN(
        P2_U2916) );
  AOI22_X1 U21714 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19690), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19689), .ZN(n19545) );
  NOR2_X2 U21715 ( .A1(n19517), .A2(n19683), .ZN(n19553) );
  NOR2_X2 U21716 ( .A1(n11245), .A2(n19685), .ZN(n19551) );
  AOI22_X1 U21717 ( .A1(n19688), .A2(n19553), .B1(n19687), .B2(n19551), .ZN(
        n19519) );
  AOI22_X1 U21718 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19689), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19690), .ZN(n19550) );
  INV_X1 U21719 ( .A(n19550), .ZN(n19552) );
  AOI22_X1 U21720 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19691), .B1(
        n19566), .B2(n19552), .ZN(n19518) );
  OAI211_X1 U21721 ( .C1(n19545), .C2(n19569), .A(n19519), .B(n19518), .ZN(
        P2_U3171) );
  AOI22_X1 U21722 ( .A1(n19566), .A2(n19554), .B1(n19694), .B2(n19551), .ZN(
        n19521) );
  AOI22_X1 U21723 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19696), .B1(
        n19553), .B2(n19695), .ZN(n19520) );
  OAI211_X1 U21724 ( .C1(n19550), .C2(n19574), .A(n19521), .B(n19520), .ZN(
        P2_U3163) );
  AOI22_X1 U21725 ( .A1(n19701), .A2(n19553), .B1(n19551), .B2(n19700), .ZN(
        n19523) );
  AOI22_X1 U21726 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19703), .B1(
        n19709), .B2(n19552), .ZN(n19522) );
  OAI211_X1 U21727 ( .C1(n19545), .C2(n19574), .A(n19523), .B(n19522), .ZN(
        P2_U3155) );
  AOI22_X1 U21728 ( .A1(n19708), .A2(n19553), .B1(n19551), .B2(n19707), .ZN(
        n19525) );
  AOI22_X1 U21729 ( .A1(n19710), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n19709), .B2(n19554), .ZN(n19524) );
  OAI211_X1 U21730 ( .C1(n19550), .C2(n19718), .A(n19525), .B(n19524), .ZN(
        P2_U3147) );
  AOI22_X1 U21731 ( .A1(n19714), .A2(n19553), .B1(n19551), .B2(n19713), .ZN(
        n19527) );
  AOI22_X1 U21732 ( .A1(n19630), .A2(n19554), .B1(
        P2_INSTQUEUE_REG_11__3__SCAN_IN), .B2(n19715), .ZN(n19526) );
  OAI211_X1 U21733 ( .C1(n19550), .C2(n19633), .A(n19527), .B(n19526), .ZN(
        P2_U3139) );
  AOI22_X1 U21734 ( .A1(n19720), .A2(n19554), .B1(n19551), .B2(n19719), .ZN(
        n19529) );
  AOI22_X1 U21735 ( .A1(n19553), .A2(n19721), .B1(n19727), .B2(n19552), .ZN(
        n19528) );
  OAI211_X1 U21736 ( .C1(n19725), .C2(n19530), .A(n19529), .B(n19528), .ZN(
        P2_U3131) );
  AOI22_X1 U21737 ( .A1(n19727), .A2(n19554), .B1(n19726), .B2(n19551), .ZN(
        n19532) );
  AOI22_X1 U21738 ( .A1(n19734), .A2(n19552), .B1(n19553), .B2(n19728), .ZN(
        n19531) );
  OAI211_X1 U21739 ( .C1(n19732), .C2(n11483), .A(n19532), .B(n19531), .ZN(
        P2_U3123) );
  AOI22_X1 U21740 ( .A1(n19734), .A2(n19554), .B1(n19551), .B2(n19733), .ZN(
        n19534) );
  AOI22_X1 U21741 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19736), .B1(
        n19735), .B2(n19553), .ZN(n19533) );
  OAI211_X1 U21742 ( .C1(n19550), .C2(n19739), .A(n19534), .B(n19533), .ZN(
        P2_U3115) );
  AOI22_X1 U21743 ( .A1(n19741), .A2(n19553), .B1(n19740), .B2(n19551), .ZN(
        n19536) );
  AOI22_X1 U21744 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19743), .B1(
        n19742), .B2(n19554), .ZN(n19535) );
  OAI211_X1 U21745 ( .C1(n19550), .C2(n19752), .A(n19536), .B(n19535), .ZN(
        P2_U3107) );
  AOI22_X1 U21746 ( .A1(n19747), .A2(n19553), .B1(n19551), .B2(n19746), .ZN(
        n19538) );
  AOI22_X1 U21747 ( .A1(n19554), .A2(n19645), .B1(
        P2_INSTQUEUE_REG_6__3__SCAN_IN), .B2(n19748), .ZN(n19537) );
  OAI211_X1 U21748 ( .C1(n19550), .C2(n19758), .A(n19538), .B(n19537), .ZN(
        P2_U3099) );
  AOI22_X1 U21749 ( .A1(n19554), .A2(n19749), .B1(n19753), .B2(n19551), .ZN(
        n19540) );
  AOI22_X1 U21750 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19755), .B1(
        n19553), .B2(n19754), .ZN(n19539) );
  OAI211_X1 U21751 ( .C1(n19550), .C2(n19650), .A(n19540), .B(n19539), .ZN(
        P2_U3091) );
  AOI22_X1 U21752 ( .A1(n19760), .A2(n19554), .B1(n19759), .B2(n19551), .ZN(
        n19542) );
  AOI22_X1 U21753 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19762), .B1(
        n19553), .B2(n19761), .ZN(n19541) );
  OAI211_X1 U21754 ( .C1(n19550), .C2(n19770), .A(n19542), .B(n19541), .ZN(
        P2_U3083) );
  AOI22_X1 U21755 ( .A1(n19552), .A2(n19774), .B1(n19765), .B2(n19551), .ZN(
        n19544) );
  AOI22_X1 U21756 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19767), .B1(
        n19553), .B2(n19766), .ZN(n19543) );
  OAI211_X1 U21757 ( .C1(n19545), .C2(n19770), .A(n19544), .B(n19543), .ZN(
        P2_U3075) );
  AOI22_X1 U21758 ( .A1(n19773), .A2(n19553), .B1(n19551), .B2(n19772), .ZN(
        n19547) );
  AOI22_X1 U21759 ( .A1(n19774), .A2(n19554), .B1(n19781), .B2(n19552), .ZN(
        n19546) );
  OAI211_X1 U21760 ( .C1(n19778), .C2(n11814), .A(n19547), .B(n19546), .ZN(
        P2_U3067) );
  AOI22_X1 U21761 ( .A1(n19780), .A2(n19553), .B1(n19551), .B2(n19779), .ZN(
        n19549) );
  AOI22_X1 U21762 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19782), .B1(
        n19781), .B2(n19554), .ZN(n19548) );
  OAI211_X1 U21763 ( .C1(n19550), .C2(n19785), .A(n19549), .B(n19548), .ZN(
        P2_U3059) );
  AOI22_X1 U21764 ( .A1(n19552), .A2(n19789), .B1(n19788), .B2(n19551), .ZN(
        n19556) );
  AOI22_X1 U21765 ( .A1(n19794), .A2(n19554), .B1(n19792), .B2(n19553), .ZN(
        n19555) );
  OAI211_X1 U21766 ( .C1(n19798), .C2(n19557), .A(n19556), .B(n19555), .ZN(
        P2_U3051) );
  AOI22_X1 U21767 ( .A1(n19558), .A2(n19612), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19670), .ZN(n19564) );
  XNOR2_X1 U21768 ( .A(n19560), .B(n19559), .ZN(n19562) );
  NAND2_X1 U21769 ( .A1(n19562), .A2(n19561), .ZN(n19563) );
  OAI211_X1 U21770 ( .C1(n19565), .C2(n19619), .A(n19564), .B(n19563), .ZN(
        P2_U2917) );
  AOI22_X1 U21771 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19690), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19689), .ZN(n19597) );
  NOR2_X2 U21772 ( .A1(n19565), .A2(n19683), .ZN(n19606) );
  AOI22_X1 U21773 ( .A1(n19688), .A2(n19606), .B1(n19687), .B2(n19604), .ZN(
        n19568) );
  AOI22_X1 U21774 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19690), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19689), .ZN(n19603) );
  AOI22_X1 U21775 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19691), .B1(
        n19566), .B2(n19605), .ZN(n19567) );
  OAI211_X1 U21776 ( .C1(n19597), .C2(n19569), .A(n19568), .B(n19567), .ZN(
        P2_U3170) );
  AOI22_X1 U21777 ( .A1(n19702), .A2(n19605), .B1(n19694), .B2(n19604), .ZN(
        n19571) );
  AOI22_X1 U21778 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19696), .B1(
        n19606), .B2(n19695), .ZN(n19570) );
  OAI211_X1 U21779 ( .C1(n19597), .C2(n19699), .A(n19571), .B(n19570), .ZN(
        P2_U3162) );
  AOI22_X1 U21780 ( .A1(n19701), .A2(n19606), .B1(n19604), .B2(n19700), .ZN(
        n19573) );
  AOI22_X1 U21781 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19703), .B1(
        n19709), .B2(n19605), .ZN(n19572) );
  OAI211_X1 U21782 ( .C1(n19597), .C2(n19574), .A(n19573), .B(n19572), .ZN(
        P2_U3154) );
  AOI22_X1 U21783 ( .A1(n19708), .A2(n19606), .B1(n19604), .B2(n19707), .ZN(
        n19576) );
  AOI22_X1 U21784 ( .A1(n19710), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n19709), .B2(n19607), .ZN(n19575) );
  OAI211_X1 U21785 ( .C1(n19603), .C2(n19718), .A(n19576), .B(n19575), .ZN(
        P2_U3146) );
  AOI22_X1 U21786 ( .A1(n19714), .A2(n19606), .B1(n19604), .B2(n19713), .ZN(
        n19578) );
  AOI22_X1 U21787 ( .A1(n19720), .A2(n19605), .B1(
        P2_INSTQUEUE_REG_11__2__SCAN_IN), .B2(n19715), .ZN(n19577) );
  OAI211_X1 U21788 ( .C1(n19597), .C2(n19718), .A(n19578), .B(n19577), .ZN(
        P2_U3138) );
  INV_X1 U21789 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n19581) );
  AOI22_X1 U21790 ( .A1(n19607), .A2(n19720), .B1(n19604), .B2(n19719), .ZN(
        n19580) );
  AOI22_X1 U21791 ( .A1(n19606), .A2(n19721), .B1(n19727), .B2(n19605), .ZN(
        n19579) );
  OAI211_X1 U21792 ( .C1(n19725), .C2(n19581), .A(n19580), .B(n19579), .ZN(
        P2_U3130) );
  INV_X1 U21793 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n19584) );
  AOI22_X1 U21794 ( .A1(n19734), .A2(n19605), .B1(n19726), .B2(n19604), .ZN(
        n19583) );
  AOI22_X1 U21795 ( .A1(n19606), .A2(n19728), .B1(n19727), .B2(n19607), .ZN(
        n19582) );
  OAI211_X1 U21796 ( .C1(n19732), .C2(n19584), .A(n19583), .B(n19582), .ZN(
        P2_U3122) );
  AOI22_X1 U21797 ( .A1(n19607), .A2(n19734), .B1(n19604), .B2(n19733), .ZN(
        n19586) );
  AOI22_X1 U21798 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19736), .B1(
        n19735), .B2(n19606), .ZN(n19585) );
  OAI211_X1 U21799 ( .C1(n19603), .C2(n19739), .A(n19586), .B(n19585), .ZN(
        P2_U3114) );
  AOI22_X1 U21800 ( .A1(n19741), .A2(n19606), .B1(n19740), .B2(n19604), .ZN(
        n19588) );
  AOI22_X1 U21801 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19743), .B1(
        n19645), .B2(n19605), .ZN(n19587) );
  OAI211_X1 U21802 ( .C1(n19597), .C2(n19739), .A(n19588), .B(n19587), .ZN(
        P2_U3106) );
  AOI22_X1 U21803 ( .A1(n19747), .A2(n19606), .B1(n19604), .B2(n19746), .ZN(
        n19590) );
  AOI22_X1 U21804 ( .A1(n19605), .A2(n19749), .B1(
        P2_INSTQUEUE_REG_6__2__SCAN_IN), .B2(n19748), .ZN(n19589) );
  OAI211_X1 U21805 ( .C1(n19597), .C2(n19752), .A(n19590), .B(n19589), .ZN(
        P2_U3098) );
  AOI22_X1 U21806 ( .A1(n19607), .A2(n19749), .B1(n19753), .B2(n19604), .ZN(
        n19592) );
  AOI22_X1 U21807 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19755), .B1(
        n19606), .B2(n19754), .ZN(n19591) );
  OAI211_X1 U21808 ( .C1(n19603), .C2(n19650), .A(n19592), .B(n19591), .ZN(
        P2_U3090) );
  AOI22_X1 U21809 ( .A1(n19607), .A2(n19760), .B1(n19759), .B2(n19604), .ZN(
        n19594) );
  AOI22_X1 U21810 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19762), .B1(
        n19606), .B2(n19761), .ZN(n19593) );
  OAI211_X1 U21811 ( .C1(n19603), .C2(n19770), .A(n19594), .B(n19593), .ZN(
        P2_U3082) );
  AOI22_X1 U21812 ( .A1(n19605), .A2(n19774), .B1(n19765), .B2(n19604), .ZN(
        n19596) );
  AOI22_X1 U21813 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19767), .B1(
        n19606), .B2(n19766), .ZN(n19595) );
  OAI211_X1 U21814 ( .C1(n19597), .C2(n19770), .A(n19596), .B(n19595), .ZN(
        P2_U3074) );
  INV_X1 U21815 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n19600) );
  AOI22_X1 U21816 ( .A1(n19773), .A2(n19606), .B1(n19604), .B2(n19772), .ZN(
        n19599) );
  AOI22_X1 U21817 ( .A1(n19774), .A2(n19607), .B1(n19781), .B2(n19605), .ZN(
        n19598) );
  OAI211_X1 U21818 ( .C1(n19778), .C2(n19600), .A(n19599), .B(n19598), .ZN(
        P2_U3066) );
  AOI22_X1 U21819 ( .A1(n19780), .A2(n19606), .B1(n19604), .B2(n19779), .ZN(
        n19602) );
  AOI22_X1 U21820 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19782), .B1(
        n19781), .B2(n19607), .ZN(n19601) );
  OAI211_X1 U21821 ( .C1(n19603), .C2(n19785), .A(n19602), .B(n19601), .ZN(
        P2_U3058) );
  INV_X1 U21822 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n19610) );
  AOI22_X1 U21823 ( .A1(n19789), .A2(n19605), .B1(n19788), .B2(n19604), .ZN(
        n19609) );
  AOI22_X1 U21824 ( .A1(n19794), .A2(n19607), .B1(n19792), .B2(n19606), .ZN(
        n19608) );
  OAI211_X1 U21825 ( .C1(n19798), .C2(n19610), .A(n19609), .B(n19608), .ZN(
        P2_U3050) );
  AOI22_X1 U21826 ( .A1(n19612), .A2(n19611), .B1(n19670), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19618) );
  AOI21_X1 U21827 ( .B1(n19615), .B2(n19614), .A(n19613), .ZN(n19616) );
  OR2_X1 U21828 ( .A1(n19616), .A2(n19677), .ZN(n19617) );
  OAI211_X1 U21829 ( .C1(n19620), .C2(n19619), .A(n19618), .B(n19617), .ZN(
        P2_U2918) );
  AOI22_X1 U21830 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19690), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19689), .ZN(n19662) );
  NOR2_X2 U21831 ( .A1(n19620), .A2(n19683), .ZN(n19665) );
  NOR2_X2 U21832 ( .A1(n19621), .A2(n19685), .ZN(n19663) );
  AOI22_X1 U21833 ( .A1(n19688), .A2(n19665), .B1(n19687), .B2(n19663), .ZN(
        n19623) );
  AOI22_X1 U21834 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19690), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19689), .ZN(n19644) );
  AOI22_X1 U21835 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19691), .B1(
        n19789), .B2(n19666), .ZN(n19622) );
  OAI211_X1 U21836 ( .C1(n19662), .C2(n19699), .A(n19623), .B(n19622), .ZN(
        P2_U3169) );
  INV_X1 U21837 ( .A(n19662), .ZN(n19664) );
  AOI22_X1 U21838 ( .A1(n19664), .A2(n19702), .B1(n19694), .B2(n19663), .ZN(
        n19625) );
  AOI22_X1 U21839 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19696), .B1(
        n19665), .B2(n19695), .ZN(n19624) );
  OAI211_X1 U21840 ( .C1(n19644), .C2(n19699), .A(n19625), .B(n19624), .ZN(
        P2_U3161) );
  AOI22_X1 U21841 ( .A1(n19701), .A2(n19665), .B1(n19663), .B2(n19700), .ZN(
        n19627) );
  AOI22_X1 U21842 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19703), .B1(
        n19702), .B2(n19666), .ZN(n19626) );
  OAI211_X1 U21843 ( .C1(n19662), .C2(n19706), .A(n19627), .B(n19626), .ZN(
        P2_U3153) );
  AOI22_X1 U21844 ( .A1(n19708), .A2(n19665), .B1(n19663), .B2(n19707), .ZN(
        n19629) );
  AOI22_X1 U21845 ( .A1(n19710), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n19709), .B2(n19666), .ZN(n19628) );
  OAI211_X1 U21846 ( .C1(n19662), .C2(n19718), .A(n19629), .B(n19628), .ZN(
        P2_U3145) );
  AOI22_X1 U21847 ( .A1(n19714), .A2(n19665), .B1(n19663), .B2(n19713), .ZN(
        n19632) );
  AOI22_X1 U21848 ( .A1(n19630), .A2(n19666), .B1(
        P2_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n19715), .ZN(n19631) );
  OAI211_X1 U21849 ( .C1(n19662), .C2(n19633), .A(n19632), .B(n19631), .ZN(
        P2_U3137) );
  INV_X1 U21850 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n19636) );
  AOI22_X1 U21851 ( .A1(n19664), .A2(n19727), .B1(n19663), .B2(n19719), .ZN(
        n19635) );
  AOI22_X1 U21852 ( .A1(n19665), .A2(n19721), .B1(n19720), .B2(n19666), .ZN(
        n19634) );
  OAI211_X1 U21853 ( .C1(n19725), .C2(n19636), .A(n19635), .B(n19634), .ZN(
        P2_U3129) );
  INV_X1 U21854 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n19639) );
  AOI22_X1 U21855 ( .A1(n19727), .A2(n19666), .B1(n19726), .B2(n19663), .ZN(
        n19638) );
  AOI22_X1 U21856 ( .A1(n19734), .A2(n19664), .B1(n19665), .B2(n19728), .ZN(
        n19637) );
  OAI211_X1 U21857 ( .C1(n19732), .C2(n19639), .A(n19638), .B(n19637), .ZN(
        P2_U3121) );
  AOI22_X1 U21858 ( .A1(n19734), .A2(n19666), .B1(n19663), .B2(n19733), .ZN(
        n19641) );
  AOI22_X1 U21859 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19736), .B1(
        n19735), .B2(n19665), .ZN(n19640) );
  OAI211_X1 U21860 ( .C1(n19662), .C2(n19739), .A(n19641), .B(n19640), .ZN(
        P2_U3113) );
  AOI22_X1 U21861 ( .A1(n19741), .A2(n19665), .B1(n19740), .B2(n19663), .ZN(
        n19643) );
  AOI22_X1 U21862 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19743), .B1(
        n19645), .B2(n19664), .ZN(n19642) );
  OAI211_X1 U21863 ( .C1(n19644), .C2(n19739), .A(n19643), .B(n19642), .ZN(
        P2_U3105) );
  AOI22_X1 U21864 ( .A1(n19747), .A2(n19665), .B1(n19663), .B2(n19746), .ZN(
        n19647) );
  AOI22_X1 U21865 ( .A1(n19645), .A2(n19666), .B1(
        P2_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n19748), .ZN(n19646) );
  OAI211_X1 U21866 ( .C1(n19662), .C2(n19758), .A(n19647), .B(n19646), .ZN(
        P2_U3097) );
  AOI22_X1 U21867 ( .A1(n19749), .A2(n19666), .B1(n19753), .B2(n19663), .ZN(
        n19649) );
  AOI22_X1 U21868 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19755), .B1(
        n19665), .B2(n19754), .ZN(n19648) );
  OAI211_X1 U21869 ( .C1(n19662), .C2(n19650), .A(n19649), .B(n19648), .ZN(
        P2_U3089) );
  AOI22_X1 U21870 ( .A1(n19760), .A2(n19666), .B1(n19663), .B2(n19759), .ZN(
        n19652) );
  AOI22_X1 U21871 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19762), .B1(
        n19665), .B2(n19761), .ZN(n19651) );
  OAI211_X1 U21872 ( .C1(n19662), .C2(n19770), .A(n19652), .B(n19651), .ZN(
        P2_U3081) );
  AOI22_X1 U21873 ( .A1(n19653), .A2(n19666), .B1(n19765), .B2(n19663), .ZN(
        n19655) );
  AOI22_X1 U21874 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19767), .B1(
        n19665), .B2(n19766), .ZN(n19654) );
  OAI211_X1 U21875 ( .C1(n19662), .C2(n19656), .A(n19655), .B(n19654), .ZN(
        P2_U3073) );
  INV_X1 U21876 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n19659) );
  AOI22_X1 U21877 ( .A1(n19773), .A2(n19665), .B1(n19663), .B2(n19772), .ZN(
        n19658) );
  AOI22_X1 U21878 ( .A1(n19774), .A2(n19666), .B1(n19781), .B2(n19664), .ZN(
        n19657) );
  OAI211_X1 U21879 ( .C1(n19778), .C2(n19659), .A(n19658), .B(n19657), .ZN(
        P2_U3065) );
  AOI22_X1 U21880 ( .A1(n19780), .A2(n19665), .B1(n19663), .B2(n19779), .ZN(
        n19661) );
  AOI22_X1 U21881 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19782), .B1(
        n19781), .B2(n19666), .ZN(n19660) );
  OAI211_X1 U21882 ( .C1(n19662), .C2(n19785), .A(n19661), .B(n19660), .ZN(
        P2_U3057) );
  AOI22_X1 U21883 ( .A1(n19664), .A2(n19789), .B1(n19788), .B2(n19663), .ZN(
        n19668) );
  AOI22_X1 U21884 ( .A1(n19794), .A2(n19666), .B1(n19792), .B2(n19665), .ZN(
        n19667) );
  OAI211_X1 U21885 ( .C1(n19798), .C2(n19669), .A(n19668), .B(n19667), .ZN(
        P2_U3049) );
  INV_X1 U21886 ( .A(n19684), .ZN(n19671) );
  AOI22_X1 U21887 ( .A1(n19672), .A2(n19671), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n19670), .ZN(n19682) );
  AOI22_X1 U21888 ( .A1(n19674), .A2(BUF2_REG_16__SCAN_IN), .B1(n19673), .B2(
        BUF1_REG_16__SCAN_IN), .ZN(n19681) );
  OAI22_X1 U21889 ( .A1(n19678), .A2(n19677), .B1(n19676), .B2(n19675), .ZN(
        n19679) );
  INV_X1 U21890 ( .A(n19679), .ZN(n19680) );
  NAND3_X1 U21891 ( .A1(n19682), .A2(n19681), .A3(n19680), .ZN(P2_U2903) );
  AOI22_X1 U21892 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19690), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19689), .ZN(n19786) );
  NOR2_X2 U21893 ( .A1(n19684), .A2(n19683), .ZN(n19791) );
  NOR2_X2 U21894 ( .A1(n19686), .A2(n19685), .ZN(n19787) );
  AOI22_X1 U21895 ( .A1(n19688), .A2(n19791), .B1(n19687), .B2(n19787), .ZN(
        n19693) );
  AOI22_X1 U21896 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19690), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19689), .ZN(n19771) );
  AOI22_X1 U21897 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19691), .B1(
        n19789), .B2(n19793), .ZN(n19692) );
  OAI211_X1 U21898 ( .C1(n19786), .C2(n19699), .A(n19693), .B(n19692), .ZN(
        P2_U3168) );
  AOI22_X1 U21899 ( .A1(n19790), .A2(n19702), .B1(n19694), .B2(n19787), .ZN(
        n19698) );
  AOI22_X1 U21900 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19696), .B1(
        n19791), .B2(n19695), .ZN(n19697) );
  OAI211_X1 U21901 ( .C1(n19771), .C2(n19699), .A(n19698), .B(n19697), .ZN(
        P2_U3160) );
  AOI22_X1 U21902 ( .A1(n19701), .A2(n19791), .B1(n19787), .B2(n19700), .ZN(
        n19705) );
  AOI22_X1 U21903 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19703), .B1(
        n19702), .B2(n19793), .ZN(n19704) );
  OAI211_X1 U21904 ( .C1(n19786), .C2(n19706), .A(n19705), .B(n19704), .ZN(
        P2_U3152) );
  AOI22_X1 U21905 ( .A1(n19708), .A2(n19791), .B1(n19787), .B2(n19707), .ZN(
        n19712) );
  AOI22_X1 U21906 ( .A1(n19710), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n19709), .B2(n19793), .ZN(n19711) );
  OAI211_X1 U21907 ( .C1(n19786), .C2(n19718), .A(n19712), .B(n19711), .ZN(
        P2_U3144) );
  AOI22_X1 U21908 ( .A1(n19714), .A2(n19791), .B1(n19787), .B2(n19713), .ZN(
        n19717) );
  AOI22_X1 U21909 ( .A1(n19790), .A2(n19720), .B1(
        P2_INSTQUEUE_REG_11__0__SCAN_IN), .B2(n19715), .ZN(n19716) );
  OAI211_X1 U21910 ( .C1(n19771), .C2(n19718), .A(n19717), .B(n19716), .ZN(
        P2_U3136) );
  INV_X1 U21911 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n19724) );
  AOI22_X1 U21912 ( .A1(n19720), .A2(n19793), .B1(n19787), .B2(n19719), .ZN(
        n19723) );
  AOI22_X1 U21913 ( .A1(n19791), .A2(n19721), .B1(n19727), .B2(n19790), .ZN(
        n19722) );
  OAI211_X1 U21914 ( .C1(n19725), .C2(n19724), .A(n19723), .B(n19722), .ZN(
        P2_U3128) );
  INV_X1 U21915 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n19731) );
  AOI22_X1 U21916 ( .A1(n19790), .A2(n19734), .B1(n19726), .B2(n19787), .ZN(
        n19730) );
  AOI22_X1 U21917 ( .A1(n19791), .A2(n19728), .B1(n19727), .B2(n19793), .ZN(
        n19729) );
  OAI211_X1 U21918 ( .C1(n19732), .C2(n19731), .A(n19730), .B(n19729), .ZN(
        P2_U3120) );
  AOI22_X1 U21919 ( .A1(n19734), .A2(n19793), .B1(n19787), .B2(n19733), .ZN(
        n19738) );
  AOI22_X1 U21920 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19736), .B1(
        n19735), .B2(n19791), .ZN(n19737) );
  OAI211_X1 U21921 ( .C1(n19786), .C2(n19739), .A(n19738), .B(n19737), .ZN(
        P2_U3112) );
  AOI22_X1 U21922 ( .A1(n19741), .A2(n19791), .B1(n19740), .B2(n19787), .ZN(
        n19745) );
  AOI22_X1 U21923 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19743), .B1(
        n19742), .B2(n19793), .ZN(n19744) );
  OAI211_X1 U21924 ( .C1(n19786), .C2(n19752), .A(n19745), .B(n19744), .ZN(
        P2_U3104) );
  AOI22_X1 U21925 ( .A1(n19747), .A2(n19791), .B1(n19787), .B2(n19746), .ZN(
        n19751) );
  AOI22_X1 U21926 ( .A1(n19790), .A2(n19749), .B1(
        P2_INSTQUEUE_REG_6__0__SCAN_IN), .B2(n19748), .ZN(n19750) );
  OAI211_X1 U21927 ( .C1(n19771), .C2(n19752), .A(n19751), .B(n19750), .ZN(
        P2_U3096) );
  AOI22_X1 U21928 ( .A1(n19790), .A2(n19760), .B1(n19753), .B2(n19787), .ZN(
        n19757) );
  AOI22_X1 U21929 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19755), .B1(
        n19791), .B2(n19754), .ZN(n19756) );
  OAI211_X1 U21930 ( .C1(n19771), .C2(n19758), .A(n19757), .B(n19756), .ZN(
        P2_U3088) );
  AOI22_X1 U21931 ( .A1(n19760), .A2(n19793), .B1(n19759), .B2(n19787), .ZN(
        n19764) );
  AOI22_X1 U21932 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19762), .B1(
        n19791), .B2(n19761), .ZN(n19763) );
  OAI211_X1 U21933 ( .C1(n19786), .C2(n19770), .A(n19764), .B(n19763), .ZN(
        P2_U3080) );
  AOI22_X1 U21934 ( .A1(n19790), .A2(n19774), .B1(n19765), .B2(n19787), .ZN(
        n19769) );
  AOI22_X1 U21935 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19767), .B1(
        n19791), .B2(n19766), .ZN(n19768) );
  OAI211_X1 U21936 ( .C1(n19771), .C2(n19770), .A(n19769), .B(n19768), .ZN(
        P2_U3072) );
  INV_X1 U21937 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n19777) );
  AOI22_X1 U21938 ( .A1(n19773), .A2(n19791), .B1(n19787), .B2(n19772), .ZN(
        n19776) );
  AOI22_X1 U21939 ( .A1(n19774), .A2(n19793), .B1(n19781), .B2(n19790), .ZN(
        n19775) );
  OAI211_X1 U21940 ( .C1(n19778), .C2(n19777), .A(n19776), .B(n19775), .ZN(
        P2_U3064) );
  AOI22_X1 U21941 ( .A1(n19780), .A2(n19791), .B1(n19787), .B2(n19779), .ZN(
        n19784) );
  AOI22_X1 U21942 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19782), .B1(
        n19781), .B2(n19793), .ZN(n19783) );
  OAI211_X1 U21943 ( .C1(n19786), .C2(n19785), .A(n19784), .B(n19783), .ZN(
        P2_U3056) );
  AOI22_X1 U21944 ( .A1(n19790), .A2(n19789), .B1(n19788), .B2(n19787), .ZN(
        n19796) );
  AOI22_X1 U21945 ( .A1(n19794), .A2(n19793), .B1(n19792), .B2(n19791), .ZN(
        n19795) );
  OAI211_X1 U21946 ( .C1(n19798), .C2(n19797), .A(n19796), .B(n19795), .ZN(
        P2_U3048) );
  INV_X1 U21947 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n20086) );
  INV_X1 U21948 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n19799) );
  AOI222_X1 U21949 ( .A1(n20086), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n20089), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n19799), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n19800) );
  INV_X1 U21950 ( .A(n19853), .ZN(n19852) );
  OAI22_X1 U21951 ( .A1(n19853), .A2(P3_ADDRESS_REG_0__SCAN_IN), .B1(
        P2_ADDRESS_REG_0__SCAN_IN), .B2(n19852), .ZN(n19801) );
  INV_X1 U21952 ( .A(n19801), .ZN(U376) );
  OAI22_X1 U21953 ( .A1(n19853), .A2(P3_ADDRESS_REG_1__SCAN_IN), .B1(
        P2_ADDRESS_REG_1__SCAN_IN), .B2(n19852), .ZN(n19802) );
  INV_X1 U21954 ( .A(n19802), .ZN(U365) );
  OAI22_X1 U21955 ( .A1(n19853), .A2(P3_ADDRESS_REG_2__SCAN_IN), .B1(
        P2_ADDRESS_REG_2__SCAN_IN), .B2(n19852), .ZN(n19803) );
  INV_X1 U21956 ( .A(n19803), .ZN(U354) );
  OAI22_X1 U21957 ( .A1(n19853), .A2(P3_ADDRESS_REG_3__SCAN_IN), .B1(
        P2_ADDRESS_REG_3__SCAN_IN), .B2(n19852), .ZN(n19804) );
  INV_X1 U21958 ( .A(n19804), .ZN(U353) );
  OAI22_X1 U21959 ( .A1(n19853), .A2(P3_ADDRESS_REG_4__SCAN_IN), .B1(
        P2_ADDRESS_REG_4__SCAN_IN), .B2(n19852), .ZN(n19805) );
  INV_X1 U21960 ( .A(n19805), .ZN(U352) );
  INV_X1 U21961 ( .A(n19853), .ZN(n19856) );
  AOI22_X1 U21962 ( .A1(n19856), .A2(n19807), .B1(n19806), .B2(n19853), .ZN(
        U351) );
  AOI22_X1 U21963 ( .A1(n19856), .A2(n19809), .B1(n19808), .B2(n19853), .ZN(
        U350) );
  AOI22_X1 U21964 ( .A1(n19856), .A2(n19811), .B1(n19810), .B2(n19853), .ZN(
        U349) );
  AOI22_X1 U21965 ( .A1(n19856), .A2(n19813), .B1(n19812), .B2(n19853), .ZN(
        U348) );
  AOI22_X1 U21966 ( .A1(n19856), .A2(n19815), .B1(n19814), .B2(n19853), .ZN(
        U347) );
  AOI22_X1 U21967 ( .A1(n19856), .A2(n19817), .B1(n19816), .B2(n19853), .ZN(
        U375) );
  AOI22_X1 U21968 ( .A1(n19856), .A2(n19819), .B1(n19818), .B2(n19853), .ZN(
        U374) );
  AOI22_X1 U21969 ( .A1(n19856), .A2(n19821), .B1(n19820), .B2(n19853), .ZN(
        U373) );
  AOI22_X1 U21970 ( .A1(n19856), .A2(n19823), .B1(n19822), .B2(n19853), .ZN(
        U372) );
  AOI22_X1 U21971 ( .A1(n19856), .A2(n19825), .B1(n19824), .B2(n19853), .ZN(
        U371) );
  AOI22_X1 U21972 ( .A1(n19856), .A2(n19827), .B1(n19826), .B2(n19853), .ZN(
        U370) );
  AOI22_X1 U21973 ( .A1(n19856), .A2(n19829), .B1(n19828), .B2(n19853), .ZN(
        U369) );
  AOI22_X1 U21974 ( .A1(n19856), .A2(n19831), .B1(n19830), .B2(n19853), .ZN(
        U368) );
  OAI22_X1 U21975 ( .A1(n19853), .A2(P3_ADDRESS_REG_18__SCAN_IN), .B1(
        P2_ADDRESS_REG_18__SCAN_IN), .B2(n19856), .ZN(n19832) );
  INV_X1 U21976 ( .A(n19832), .ZN(U367) );
  OAI22_X1 U21977 ( .A1(n19853), .A2(P3_ADDRESS_REG_19__SCAN_IN), .B1(
        P2_ADDRESS_REG_19__SCAN_IN), .B2(n19852), .ZN(n19833) );
  INV_X1 U21978 ( .A(n19833), .ZN(U366) );
  AOI22_X1 U21979 ( .A1(n19856), .A2(n19835), .B1(n19834), .B2(n19853), .ZN(
        U364) );
  AOI22_X1 U21980 ( .A1(n19856), .A2(n19837), .B1(n19836), .B2(n19853), .ZN(
        U363) );
  AOI22_X1 U21981 ( .A1(n19856), .A2(n19839), .B1(n19838), .B2(n19853), .ZN(
        U362) );
  AOI22_X1 U21982 ( .A1(n19856), .A2(n19841), .B1(n19840), .B2(n19853), .ZN(
        U361) );
  AOI22_X1 U21983 ( .A1(n19852), .A2(n19843), .B1(n19842), .B2(n19853), .ZN(
        U360) );
  AOI22_X1 U21984 ( .A1(n19856), .A2(n19845), .B1(n19844), .B2(n19853), .ZN(
        U359) );
  AOI22_X1 U21985 ( .A1(n19856), .A2(n19847), .B1(n19846), .B2(n19853), .ZN(
        U358) );
  AOI22_X1 U21986 ( .A1(n19856), .A2(n19849), .B1(n19848), .B2(n19853), .ZN(
        U357) );
  AOI22_X1 U21987 ( .A1(n19852), .A2(n19851), .B1(n19850), .B2(n19853), .ZN(
        U356) );
  INV_X1 U21988 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n19855) );
  AOI22_X1 U21989 ( .A1(n19856), .A2(n19855), .B1(n19854), .B2(n19853), .ZN(
        U355) );
  AOI22_X1 U21990 ( .A1(n21257), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19858) );
  OAI21_X1 U21991 ( .B1(n21680), .B2(n19877), .A(n19858), .ZN(P1_U2936) );
  AOI22_X1 U21992 ( .A1(n19868), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19859) );
  OAI21_X1 U21993 ( .B1(n21685), .B2(n19877), .A(n19859), .ZN(P1_U2935) );
  AOI22_X1 U21994 ( .A1(n19868), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19860) );
  OAI21_X1 U21995 ( .B1(n21691), .B2(n19877), .A(n19860), .ZN(P1_U2934) );
  AOI22_X1 U21996 ( .A1(n19868), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19861) );
  OAI21_X1 U21997 ( .B1(n19862), .B2(n19877), .A(n19861), .ZN(P1_U2933) );
  AOI22_X1 U21998 ( .A1(n21257), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19863) );
  OAI21_X1 U21999 ( .B1(n21700), .B2(n19877), .A(n19863), .ZN(P1_U2932) );
  AOI22_X1 U22000 ( .A1(n19868), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19864) );
  OAI21_X1 U22001 ( .B1(n12875), .B2(n19877), .A(n19864), .ZN(P1_U2931) );
  AOI22_X1 U22002 ( .A1(n19868), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19866) );
  OAI21_X1 U22003 ( .B1(n21711), .B2(n19877), .A(n19866), .ZN(P1_U2930) );
  AOI22_X1 U22004 ( .A1(n21257), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19867) );
  OAI21_X1 U22005 ( .B1(n15264), .B2(n19877), .A(n19867), .ZN(P1_U2929) );
  INV_X1 U22006 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n21723) );
  AOI22_X1 U22007 ( .A1(n19868), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19869) );
  OAI21_X1 U22008 ( .B1(n21723), .B2(n19877), .A(n19869), .ZN(P1_U2928) );
  INV_X1 U22009 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n21731) );
  AOI22_X1 U22010 ( .A1(n21257), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19870) );
  OAI21_X1 U22011 ( .B1(n21731), .B2(n19877), .A(n19870), .ZN(P1_U2927) );
  INV_X1 U22012 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n21738) );
  AOI22_X1 U22013 ( .A1(n21257), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19871) );
  OAI21_X1 U22014 ( .B1(n21738), .B2(n19877), .A(n19871), .ZN(P1_U2926) );
  INV_X1 U22015 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n21744) );
  AOI22_X1 U22016 ( .A1(n21257), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19872) );
  OAI21_X1 U22017 ( .B1(n21744), .B2(n19877), .A(n19872), .ZN(P1_U2925) );
  INV_X1 U22018 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n21751) );
  AOI22_X1 U22019 ( .A1(n21257), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19873) );
  OAI21_X1 U22020 ( .B1(n21751), .B2(n19877), .A(n19873), .ZN(P1_U2924) );
  INV_X1 U22021 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n21758) );
  AOI22_X1 U22022 ( .A1(n21257), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19874) );
  OAI21_X1 U22023 ( .B1(n21758), .B2(n19877), .A(n19874), .ZN(P1_U2923) );
  INV_X1 U22024 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n21767) );
  AOI22_X1 U22025 ( .A1(n21257), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19875) );
  OAI21_X1 U22026 ( .B1(n21767), .B2(n19877), .A(n19875), .ZN(P1_U2922) );
  AOI22_X1 U22027 ( .A1(n21257), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n19865), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19876) );
  OAI21_X1 U22028 ( .B1(n19878), .B2(n19877), .A(n19876), .ZN(P1_U2921) );
  OR2_X1 U22029 ( .A1(n12613), .A2(n22308), .ZN(n21627) );
  INV_X1 U22030 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n19880) );
  OR2_X1 U22031 ( .A1(n22308), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n19899) );
  OAI222_X1 U22032 ( .A1(n21627), .A2(n21418), .B1(n19879), .B2(n22307), .C1(
        n19880), .C2(n19899), .ZN(P1_U3197) );
  INV_X1 U22033 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n19881) );
  OAI222_X1 U22034 ( .A1(n19899), .A2(n14961), .B1(n19881), .B2(n22307), .C1(
        n19880), .C2(n21627), .ZN(P1_U3198) );
  INV_X1 U22035 ( .A(n19899), .ZN(n19912) );
  INV_X1 U22036 ( .A(n22307), .ZN(n19913) );
  INV_X1 U22037 ( .A(n21627), .ZN(n19914) );
  AOI222_X1 U22038 ( .A1(n19912), .A2(P1_REIP_REG_4__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n19913), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n19914), .ZN(n19882) );
  INV_X1 U22039 ( .A(n19882), .ZN(P1_U3199) );
  AOI222_X1 U22040 ( .A1(n19912), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n19913), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n19914), .ZN(n19883) );
  INV_X1 U22041 ( .A(n19883), .ZN(P1_U3200) );
  AOI222_X1 U22042 ( .A1(n19914), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n19913), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n19912), .ZN(n19884) );
  INV_X1 U22043 ( .A(n19884), .ZN(P1_U3201) );
  AOI22_X1 U22044 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19912), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n22308), .ZN(n19885) );
  OAI21_X1 U22045 ( .B1(n19886), .B2(n21627), .A(n19885), .ZN(P1_U3202) );
  AOI22_X1 U22046 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19914), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n22308), .ZN(n19887) );
  OAI21_X1 U22047 ( .B1(n21487), .B2(n19899), .A(n19887), .ZN(P1_U3203) );
  AOI222_X1 U22048 ( .A1(n19912), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n19913), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n19914), .ZN(n19888) );
  INV_X1 U22049 ( .A(n19888), .ZN(P1_U3204) );
  AOI222_X1 U22050 ( .A1(n19912), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n19913), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n19914), .ZN(n19889) );
  INV_X1 U22051 ( .A(n19889), .ZN(P1_U3205) );
  AOI22_X1 U22052 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n19912), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n22308), .ZN(n19890) );
  OAI21_X1 U22053 ( .B1(n21496), .B2(n21627), .A(n19890), .ZN(P1_U3206) );
  AOI22_X1 U22054 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n19914), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n19913), .ZN(n19891) );
  OAI21_X1 U22055 ( .B1(n21313), .B2(n19899), .A(n19891), .ZN(P1_U3207) );
  AOI22_X1 U22056 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n19912), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n19913), .ZN(n19892) );
  OAI21_X1 U22057 ( .B1(n21313), .B2(n21627), .A(n19892), .ZN(P1_U3208) );
  AOI22_X1 U22058 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n19914), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n19913), .ZN(n19893) );
  OAI21_X1 U22059 ( .B1(n19894), .B2(n19899), .A(n19893), .ZN(P1_U3209) );
  AOI222_X1 U22060 ( .A1(n19912), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n19913), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n19914), .ZN(n19895) );
  INV_X1 U22061 ( .A(n19895), .ZN(P1_U3210) );
  AOI222_X1 U22062 ( .A1(n19914), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n19913), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n19912), .ZN(n19896) );
  INV_X1 U22063 ( .A(n19896), .ZN(P1_U3211) );
  AOI22_X1 U22064 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n19912), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n19913), .ZN(n19897) );
  OAI21_X1 U22065 ( .B1(n21359), .B2(n21627), .A(n19897), .ZN(P1_U3212) );
  AOI22_X1 U22066 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(n19914), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n19913), .ZN(n19898) );
  OAI21_X1 U22067 ( .B1(n21576), .B2(n19899), .A(n19898), .ZN(P1_U3213) );
  AOI222_X1 U22068 ( .A1(n19912), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n19913), .C1(P1_REIP_REG_18__SCAN_IN), 
        .C2(n19914), .ZN(n19900) );
  INV_X1 U22069 ( .A(n19900), .ZN(P1_U3214) );
  AOI222_X1 U22070 ( .A1(n19912), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n19913), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n19914), .ZN(n19901) );
  INV_X1 U22071 ( .A(n19901), .ZN(P1_U3215) );
  AOI222_X1 U22072 ( .A1(n19912), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n19913), .C1(P1_REIP_REG_20__SCAN_IN), 
        .C2(n19914), .ZN(n19902) );
  INV_X1 U22073 ( .A(n19902), .ZN(P1_U3216) );
  AOI222_X1 U22074 ( .A1(n19912), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n19913), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n19914), .ZN(n19903) );
  INV_X1 U22075 ( .A(n19903), .ZN(P1_U3217) );
  AOI222_X1 U22076 ( .A1(n19914), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n19913), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n19912), .ZN(n19904) );
  INV_X1 U22077 ( .A(n19904), .ZN(P1_U3218) );
  AOI222_X1 U22078 ( .A1(n19914), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n19913), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n19912), .ZN(n19905) );
  INV_X1 U22079 ( .A(n19905), .ZN(P1_U3219) );
  AOI222_X1 U22080 ( .A1(n19912), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n19913), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n19914), .ZN(n19906) );
  INV_X1 U22081 ( .A(n19906), .ZN(P1_U3220) );
  AOI222_X1 U22082 ( .A1(n19912), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n19913), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n19914), .ZN(n19907) );
  INV_X1 U22083 ( .A(n19907), .ZN(P1_U3221) );
  AOI222_X1 U22084 ( .A1(n19914), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n19913), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n19912), .ZN(n19908) );
  INV_X1 U22085 ( .A(n19908), .ZN(P1_U3222) );
  AOI222_X1 U22086 ( .A1(n19912), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n19913), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n19914), .ZN(n19909) );
  INV_X1 U22087 ( .A(n19909), .ZN(P1_U3223) );
  AOI222_X1 U22088 ( .A1(n19914), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n19913), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n19912), .ZN(n19910) );
  INV_X1 U22089 ( .A(n19910), .ZN(P1_U3224) );
  AOI222_X1 U22090 ( .A1(n19914), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n19913), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n19912), .ZN(n19911) );
  INV_X1 U22091 ( .A(n19911), .ZN(P1_U3225) );
  AOI222_X1 U22092 ( .A1(n19914), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n19913), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n19912), .ZN(n19915) );
  INV_X1 U22093 ( .A(n19915), .ZN(P1_U3226) );
  OAI22_X1 U22094 ( .A1(n22308), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n22307), .ZN(n19916) );
  INV_X1 U22095 ( .A(n19916), .ZN(P1_U3458) );
  AOI221_X1 U22096 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(P1_REIP_REG_1__SCAN_IN), 
        .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(P1_REIP_REG_1__SCAN_IN), .A(
        P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19927) );
  NOR4_X1 U22097 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19920) );
  NOR4_X1 U22098 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19919) );
  NOR4_X1 U22099 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A3(P1_DATAWIDTH_REG_3__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_2__SCAN_IN), .ZN(n19918) );
  NOR4_X1 U22100 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_7__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19917) );
  NAND4_X1 U22101 ( .A1(n19920), .A2(n19919), .A3(n19918), .A4(n19917), .ZN(
        n19926) );
  NOR4_X1 U22102 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_27__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n19924) );
  AOI211_X1 U22103 ( .C1(P1_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A(P1_DATAWIDTH_REG_31__SCAN_IN), .B(
        P1_DATAWIDTH_REG_30__SCAN_IN), .ZN(n19923) );
  NOR4_X1 U22104 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_19__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19922) );
  NOR4_X1 U22105 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_24__SCAN_IN), .A3(P1_DATAWIDTH_REG_23__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_22__SCAN_IN), .ZN(n19921) );
  NAND4_X1 U22106 ( .A1(n19924), .A2(n19923), .A3(n19922), .A4(n19921), .ZN(
        n19925) );
  NOR2_X1 U22107 ( .A1(n19926), .A2(n19925), .ZN(n19939) );
  MUX2_X1 U22108 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .B(n19927), .S(n19939), 
        .Z(P1_U2808) );
  OAI22_X1 U22109 ( .A1(n22308), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n22307), .ZN(n19928) );
  INV_X1 U22110 ( .A(n19928), .ZN(P1_U3459) );
  AOI21_X1 U22111 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n19929) );
  OAI221_X1 U22112 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19929), .C1(n21418), 
        .C2(P1_REIP_REG_0__SCAN_IN), .A(n19939), .ZN(n19930) );
  OAI21_X1 U22113 ( .B1(n19939), .B2(n19931), .A(n19930), .ZN(P1_U3481) );
  OAI22_X1 U22114 ( .A1(n22308), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n22307), .ZN(n19932) );
  INV_X1 U22115 ( .A(n19932), .ZN(P1_U3460) );
  NOR3_X1 U22116 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19933) );
  OAI21_X1 U22117 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19933), .A(n19939), .ZN(
        n19934) );
  OAI21_X1 U22118 ( .B1(n19939), .B2(n19935), .A(n19934), .ZN(P1_U2807) );
  OAI22_X1 U22119 ( .A1(n22308), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n22307), .ZN(n19936) );
  INV_X1 U22120 ( .A(n19936), .ZN(P1_U3461) );
  OAI21_X1 U22121 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n19939), .ZN(n19937) );
  OAI21_X1 U22122 ( .B1(n19939), .B2(n19938), .A(n19937), .ZN(P1_U3482) );
  AOI22_X1 U22123 ( .A1(n19943), .A2(n19942), .B1(n19941), .B2(n19940), .ZN(
        n19944) );
  OAI21_X1 U22124 ( .B1(n19946), .B2(n19945), .A(n19944), .ZN(P1_U2863) );
  INV_X1 U22125 ( .A(n19947), .ZN(n19949) );
  AOI21_X1 U22126 ( .B1(n19949), .B2(n21400), .A(n19948), .ZN(n21405) );
  NOR2_X1 U22127 ( .A1(n21378), .A2(n19950), .ZN(n21403) );
  INV_X1 U22128 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19951) );
  AOI21_X1 U22129 ( .B1(n19952), .B2(n19983), .A(n19951), .ZN(n19953) );
  AOI211_X1 U22130 ( .C1(n21405), .C2(n20020), .A(n21403), .B(n19953), .ZN(
        n19954) );
  OAI21_X1 U22131 ( .B1(n19957), .B2(n19955), .A(n19954), .ZN(P1_U2999) );
  INV_X1 U22132 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n21440) );
  OAI22_X1 U22133 ( .A1(n21449), .A2(n19957), .B1(n21452), .B2(n20025), .ZN(
        n19958) );
  AOI21_X1 U22134 ( .B1(n20020), .B2(n21293), .A(n19958), .ZN(n19960) );
  INV_X1 U22135 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n21443) );
  NOR2_X1 U22136 ( .A1(n21378), .A2(n21443), .ZN(n21299) );
  INV_X1 U22137 ( .A(n21299), .ZN(n19959) );
  OAI211_X1 U22138 ( .C1(n19983), .C2(n21440), .A(n19960), .B(n19959), .ZN(
        P1_U2994) );
  INV_X1 U22139 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n21472) );
  INV_X1 U22140 ( .A(n21478), .ZN(n19961) );
  AOI222_X1 U22141 ( .A1(n19962), .A2(n20020), .B1(n20021), .B2(n21475), .C1(
        n19961), .C2(n20000), .ZN(n19964) );
  OAI211_X1 U22142 ( .C1(n19983), .C2(n21472), .A(n19964), .B(n19963), .ZN(
        P1_U2992) );
  MUX2_X1 U22143 ( .A(n19965), .B(n19974), .S(n19975), .Z(n19967) );
  INV_X1 U22144 ( .A(n19967), .ZN(n19969) );
  INV_X1 U22145 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n19966) );
  NOR2_X1 U22146 ( .A1(n19967), .A2(n19966), .ZN(n19977) );
  INV_X1 U22147 ( .A(n19977), .ZN(n19968) );
  OAI21_X1 U22148 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n19969), .A(
        n19968), .ZN(n21306) );
  AOI22_X1 U22149 ( .A1(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n20015), .B1(
        n21390), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n19973) );
  INV_X1 U22150 ( .A(n19970), .ZN(n21505) );
  INV_X1 U22151 ( .A(n19971), .ZN(n21504) );
  AOI22_X1 U22152 ( .A1(n21505), .A2(n20021), .B1(n20000), .B2(n21504), .ZN(
        n19972) );
  OAI211_X1 U22153 ( .C1(n21578), .C2(n21306), .A(n19973), .B(n19972), .ZN(
        P1_U2989) );
  INV_X1 U22154 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n19982) );
  NOR2_X1 U22155 ( .A1(n19977), .A2(n19974), .ZN(n19976) );
  MUX2_X1 U22156 ( .A(n19977), .B(n19976), .S(n19975), .Z(n19978) );
  XNOR2_X1 U22157 ( .A(n19978), .B(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n21328) );
  OAI22_X1 U22158 ( .A1(n21328), .A2(n21578), .B1(n20025), .B2(n21515), .ZN(
        n19979) );
  AOI21_X1 U22159 ( .B1(n20021), .B2(n19980), .A(n19979), .ZN(n19981) );
  NAND2_X1 U22160 ( .A1(n21390), .A2(P1_REIP_REG_11__SCAN_IN), .ZN(n21321) );
  OAI211_X1 U22161 ( .C1(n19983), .C2(n19982), .A(n19981), .B(n21321), .ZN(
        P1_U2988) );
  AOI21_X1 U22162 ( .B1(n19986), .B2(n19985), .A(n19984), .ZN(n21320) );
  AOI22_X1 U22163 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n20015), .B1(
        n21390), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n19989) );
  INV_X1 U22164 ( .A(n19987), .ZN(n21524) );
  AOI22_X1 U22165 ( .A1(n20000), .A2(n21525), .B1(n20021), .B2(n21524), .ZN(
        n19988) );
  OAI211_X1 U22166 ( .C1(n21320), .C2(n21578), .A(n19989), .B(n19988), .ZN(
        P1_U2987) );
  NOR2_X1 U22167 ( .A1(n19991), .A2(n19990), .ZN(n19994) );
  INV_X1 U22168 ( .A(n19992), .ZN(n19993) );
  AOI21_X1 U22169 ( .B1(n19995), .B2(n19994), .A(n19993), .ZN(n19997) );
  XNOR2_X1 U22170 ( .A(n20009), .B(n21272), .ZN(n19996) );
  XNOR2_X1 U22171 ( .A(n19997), .B(n19996), .ZN(n21275) );
  AOI22_X1 U22172 ( .A1(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n20015), .B1(
        n21390), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n20003) );
  INV_X1 U22173 ( .A(n19998), .ZN(n20001) );
  AOI22_X1 U22174 ( .A1(n20001), .A2(n20021), .B1(n20000), .B2(n19999), .ZN(
        n20002) );
  OAI211_X1 U22175 ( .C1(n21275), .C2(n21578), .A(n20003), .B(n20002), .ZN(
        P1_U2985) );
  AOI22_X1 U22176 ( .A1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n20015), .B1(
        n21390), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n20013) );
  AOI21_X1 U22177 ( .B1(n20006), .B2(n20005), .A(n20004), .ZN(n20011) );
  INV_X1 U22178 ( .A(n20007), .ZN(n20008) );
  AOI21_X1 U22179 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n20009), .A(
        n20008), .ZN(n20010) );
  XNOR2_X1 U22180 ( .A(n20011), .B(n20010), .ZN(n21364) );
  AOI22_X1 U22181 ( .A1(n21542), .A2(n20021), .B1(n21364), .B2(n20020), .ZN(
        n20012) );
  OAI211_X1 U22182 ( .C1(n20025), .C2(n20014), .A(n20013), .B(n20012), .ZN(
        P1_U2983) );
  AOI22_X1 U22183 ( .A1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n20015), .B1(
        n21390), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n20024) );
  INV_X1 U22184 ( .A(n21572), .ZN(n20022) );
  OAI21_X1 U22185 ( .B1(n20018), .B2(n20017), .A(n20016), .ZN(n20019) );
  INV_X1 U22186 ( .A(n20019), .ZN(n21349) );
  AOI22_X1 U22187 ( .A1(n20022), .A2(n20021), .B1(n20020), .B2(n21349), .ZN(
        n20023) );
  OAI211_X1 U22188 ( .C1(n20025), .C2(n21564), .A(n20024), .B(n20023), .ZN(
        P1_U2981) );
  OAI21_X1 U22189 ( .B1(n21625), .B2(P1_D_C_N_REG_SCAN_IN), .A(n22308), .ZN(
        n20026) );
  OAI21_X1 U22190 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n22308), .A(n20026), 
        .ZN(P1_U2804) );
  AOI22_X1 U22191 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n10968), .ZN(n20028) );
  OAI21_X1 U22192 ( .B1(n14950), .B2(n20088), .A(n20028), .ZN(U247) );
  AOI22_X1 U22193 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n10968), .ZN(n20029) );
  OAI21_X1 U22194 ( .B1(n20030), .B2(n20088), .A(n20029), .ZN(U246) );
  AOI22_X1 U22195 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n10968), .ZN(n20031) );
  OAI21_X1 U22196 ( .B1(n20032), .B2(n20088), .A(n20031), .ZN(U245) );
  AOI22_X1 U22197 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n10968), .ZN(n20033) );
  OAI21_X1 U22198 ( .B1(n20034), .B2(n20088), .A(n20033), .ZN(U244) );
  AOI22_X1 U22199 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n10968), .ZN(n20035) );
  OAI21_X1 U22200 ( .B1(n20036), .B2(n20088), .A(n20035), .ZN(U243) );
  AOI22_X1 U22201 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n10968), .ZN(n20037) );
  OAI21_X1 U22202 ( .B1(n20038), .B2(n20088), .A(n20037), .ZN(U242) );
  AOI22_X1 U22203 ( .A1(P1_DATAO_REG_6__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_6__SCAN_IN), .B2(n10968), .ZN(n20039) );
  OAI21_X1 U22204 ( .B1(n20040), .B2(n20088), .A(n20039), .ZN(U241) );
  AOI22_X1 U22205 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n10968), .ZN(n20041) );
  OAI21_X1 U22206 ( .B1(n20042), .B2(n20088), .A(n20041), .ZN(U240) );
  INV_X1 U22207 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n20044) );
  AOI22_X1 U22208 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n10968), .ZN(n20043) );
  OAI21_X1 U22209 ( .B1(n20044), .B2(n20088), .A(n20043), .ZN(U239) );
  AOI22_X1 U22210 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n10968), .ZN(n20045) );
  OAI21_X1 U22211 ( .B1(n20046), .B2(n20088), .A(n20045), .ZN(U238) );
  AOI22_X1 U22212 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n10968), .ZN(n20047) );
  OAI21_X1 U22213 ( .B1(n20048), .B2(n20088), .A(n20047), .ZN(U237) );
  INV_X1 U22214 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n20050) );
  AOI22_X1 U22215 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n10968), .ZN(n20049) );
  OAI21_X1 U22216 ( .B1(n20050), .B2(n20088), .A(n20049), .ZN(U236) );
  AOI22_X1 U22217 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n10968), .ZN(n20051) );
  OAI21_X1 U22218 ( .B1(n20052), .B2(n20088), .A(n20051), .ZN(U235) );
  INV_X1 U22219 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n20054) );
  AOI22_X1 U22220 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n10968), .ZN(n20053) );
  OAI21_X1 U22221 ( .B1(n20054), .B2(n20088), .A(n20053), .ZN(U234) );
  AOI22_X1 U22222 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n10968), .ZN(n20055) );
  OAI21_X1 U22223 ( .B1(n14399), .B2(n20088), .A(n20055), .ZN(U233) );
  AOI22_X1 U22224 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n10968), .ZN(n20056) );
  OAI21_X1 U22225 ( .B1(n14797), .B2(n20088), .A(n20056), .ZN(U232) );
  AOI22_X1 U22226 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n10968), .ZN(n20057) );
  OAI21_X1 U22227 ( .B1(n20058), .B2(n20088), .A(n20057), .ZN(U231) );
  AOI22_X1 U22228 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n10968), .ZN(n20059) );
  OAI21_X1 U22229 ( .B1(n20060), .B2(n20088), .A(n20059), .ZN(U230) );
  AOI22_X1 U22230 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n10968), .ZN(n20061) );
  OAI21_X1 U22231 ( .B1(n20062), .B2(n20088), .A(n20061), .ZN(U229) );
  AOI22_X1 U22232 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n10968), .ZN(n20063) );
  OAI21_X1 U22233 ( .B1(n20064), .B2(n20088), .A(n20063), .ZN(U228) );
  AOI22_X1 U22234 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n10968), .ZN(n20065) );
  OAI21_X1 U22235 ( .B1(n20066), .B2(n20088), .A(n20065), .ZN(U227) );
  AOI22_X1 U22236 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n10968), .ZN(n20067) );
  OAI21_X1 U22237 ( .B1(n20068), .B2(n20088), .A(n20067), .ZN(U226) );
  INV_X1 U22238 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n22153) );
  AOI22_X1 U22239 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n10968), .ZN(n20069) );
  OAI21_X1 U22240 ( .B1(n22153), .B2(n20088), .A(n20069), .ZN(U225) );
  AOI22_X1 U22241 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n10968), .ZN(n20070) );
  OAI21_X1 U22242 ( .B1(n20071), .B2(n20088), .A(n20070), .ZN(U224) );
  AOI22_X1 U22243 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n10968), .ZN(n20072) );
  OAI21_X1 U22244 ( .B1(n20073), .B2(n20088), .A(n20072), .ZN(U223) );
  AOI22_X1 U22245 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n10968), .ZN(n20074) );
  OAI21_X1 U22246 ( .B1(n20075), .B2(n20088), .A(n20074), .ZN(U222) );
  AOI22_X1 U22247 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n10968), .ZN(n20076) );
  OAI21_X1 U22248 ( .B1(n20077), .B2(n20088), .A(n20076), .ZN(U221) );
  AOI22_X1 U22249 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n10968), .ZN(n20079) );
  OAI21_X1 U22250 ( .B1(n20080), .B2(n20088), .A(n20079), .ZN(U220) );
  AOI22_X1 U22251 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n10968), .ZN(n20081) );
  OAI21_X1 U22252 ( .B1(n20082), .B2(n20088), .A(n20081), .ZN(U219) );
  AOI22_X1 U22253 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n10968), .ZN(n20083) );
  OAI21_X1 U22254 ( .B1(n20084), .B2(n20088), .A(n20083), .ZN(U218) );
  INV_X1 U22255 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n22147) );
  AOI22_X1 U22256 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n20078), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n10968), .ZN(n20085) );
  OAI21_X1 U22257 ( .B1(n22147), .B2(n20088), .A(n20085), .ZN(U217) );
  OAI222_X1 U22258 ( .A1(U212), .A2(n20089), .B1(n20088), .B2(n20087), .C1(
        U214), .C2(n20086), .ZN(U216) );
  AOI22_X1 U22259 ( .A1(n22307), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20090), 
        .B2(n22308), .ZN(P1_U3483) );
  OAI21_X1 U22260 ( .B1(P3_STATEBS16_REG_SCAN_IN), .B2(n20559), .A(n20091), 
        .ZN(n20092) );
  AOI211_X1 U22261 ( .C1(n20093), .C2(n20092), .A(n21619), .B(n21098), .ZN(
        n20096) );
  OAI21_X1 U22262 ( .B1(n20096), .B2(n20095), .A(n20094), .ZN(n20102) );
  AOI22_X1 U22263 ( .A1(n20098), .A2(n21659), .B1(n20097), .B2(n21244), .ZN(
        n20100) );
  NAND2_X1 U22264 ( .A1(n20100), .A2(n20099), .ZN(n20101) );
  MUX2_X1 U22265 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .B(n20102), .S(n20101), 
        .Z(P3_U3296) );
  NOR2_X2 U22266 ( .A1(n21222), .A2(n20104), .ZN(n20137) );
  AOI22_X1 U22267 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n20137), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n20140), .ZN(n20105) );
  OAI21_X1 U22268 ( .B1(n20123), .B2(n20139), .A(n20105), .ZN(P3_U2768) );
  INV_X1 U22269 ( .A(n20137), .ZN(n20145) );
  AOI22_X1 U22270 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20143), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n20142), .ZN(n20106) );
  OAI21_X1 U22271 ( .B1(n20623), .B2(n20145), .A(n20106), .ZN(P3_U2769) );
  AOI22_X1 U22272 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20143), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n20142), .ZN(n20107) );
  OAI21_X1 U22273 ( .B1(n20647), .B2(n20145), .A(n20107), .ZN(P3_U2770) );
  AOI22_X1 U22274 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20143), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n20142), .ZN(n20108) );
  OAI21_X1 U22275 ( .B1(n20109), .B2(n20145), .A(n20108), .ZN(P3_U2771) );
  AOI22_X1 U22276 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n20137), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n20140), .ZN(n20110) );
  OAI21_X1 U22277 ( .B1(n20611), .B2(n20139), .A(n20110), .ZN(P3_U2772) );
  AOI22_X1 U22278 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n20137), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n20140), .ZN(n20111) );
  OAI21_X1 U22279 ( .B1(n20605), .B2(n20139), .A(n20111), .ZN(P3_U2773) );
  AOI22_X1 U22280 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n20137), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n20140), .ZN(n20112) );
  OAI21_X1 U22281 ( .B1(n20600), .B2(n20139), .A(n20112), .ZN(P3_U2774) );
  AOI22_X1 U22282 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n20137), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n20140), .ZN(n20113) );
  OAI21_X1 U22283 ( .B1(n20595), .B2(n20139), .A(n20113), .ZN(P3_U2775) );
  AOI22_X1 U22284 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20143), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n20140), .ZN(n20114) );
  OAI21_X1 U22285 ( .B1(n11089), .B2(n20145), .A(n20114), .ZN(P3_U2776) );
  INV_X1 U22286 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n20589) );
  AOI22_X1 U22287 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n20137), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n20140), .ZN(n20115) );
  OAI21_X1 U22288 ( .B1(n20589), .B2(n20139), .A(n20115), .ZN(P3_U2777) );
  INV_X1 U22289 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n20583) );
  AOI22_X1 U22290 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n20137), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n20140), .ZN(n20116) );
  OAI21_X1 U22291 ( .B1(n20583), .B2(n20139), .A(n20116), .ZN(P3_U2778) );
  AOI22_X1 U22292 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20143), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n20140), .ZN(n20117) );
  OAI21_X1 U22293 ( .B1(n20689), .B2(n20145), .A(n20117), .ZN(P3_U2779) );
  INV_X1 U22294 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n20575) );
  AOI22_X1 U22295 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n20137), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n20142), .ZN(n20118) );
  OAI21_X1 U22296 ( .B1(n20575), .B2(n20139), .A(n20118), .ZN(P3_U2780) );
  INV_X1 U22297 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n20570) );
  AOI22_X1 U22298 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n20137), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n20142), .ZN(n20119) );
  OAI21_X1 U22299 ( .B1(n20570), .B2(n20139), .A(n20119), .ZN(P3_U2781) );
  AOI22_X1 U22300 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20143), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n20142), .ZN(n20120) );
  OAI21_X1 U22301 ( .B1(n20121), .B2(n20145), .A(n20120), .ZN(P3_U2782) );
  AOI22_X1 U22302 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n20137), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n20142), .ZN(n20122) );
  OAI21_X1 U22303 ( .B1(n20123), .B2(n20139), .A(n20122), .ZN(P3_U2783) );
  AOI22_X1 U22304 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20143), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n20142), .ZN(n20124) );
  OAI21_X1 U22305 ( .B1(n20591), .B2(n20145), .A(n20124), .ZN(P3_U2784) );
  AOI22_X1 U22306 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20143), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n20142), .ZN(n20125) );
  OAI21_X1 U22307 ( .B1(n20618), .B2(n20145), .A(n20125), .ZN(P3_U2785) );
  AOI22_X1 U22308 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20143), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n20142), .ZN(n20126) );
  OAI21_X1 U22309 ( .B1(n20614), .B2(n20145), .A(n20126), .ZN(P3_U2786) );
  AOI22_X1 U22310 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n20137), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n20142), .ZN(n20127) );
  OAI21_X1 U22311 ( .B1(n20611), .B2(n20139), .A(n20127), .ZN(P3_U2787) );
  AOI22_X1 U22312 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n20137), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n20142), .ZN(n20128) );
  OAI21_X1 U22313 ( .B1(n20605), .B2(n20139), .A(n20128), .ZN(P3_U2788) );
  AOI22_X1 U22314 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n20137), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n20142), .ZN(n20129) );
  OAI21_X1 U22315 ( .B1(n20600), .B2(n20139), .A(n20129), .ZN(P3_U2789) );
  AOI22_X1 U22316 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n20137), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n20142), .ZN(n20130) );
  OAI21_X1 U22317 ( .B1(n20595), .B2(n20139), .A(n20130), .ZN(P3_U2790) );
  AOI22_X1 U22318 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20143), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n20142), .ZN(n20131) );
  OAI21_X1 U22319 ( .B1(n20132), .B2(n20145), .A(n20131), .ZN(P3_U2791) );
  AOI22_X1 U22320 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n20137), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n20142), .ZN(n20133) );
  OAI21_X1 U22321 ( .B1(n20589), .B2(n20139), .A(n20133), .ZN(P3_U2792) );
  AOI22_X1 U22322 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n20137), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n20142), .ZN(n20134) );
  OAI21_X1 U22323 ( .B1(n20583), .B2(n20139), .A(n20134), .ZN(P3_U2793) );
  AOI22_X1 U22324 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20143), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n20140), .ZN(n20135) );
  OAI21_X1 U22325 ( .B1(n20620), .B2(n20145), .A(n20135), .ZN(P3_U2794) );
  AOI22_X1 U22326 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n20137), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n20142), .ZN(n20136) );
  OAI21_X1 U22327 ( .B1(n20575), .B2(n20139), .A(n20136), .ZN(P3_U2795) );
  AOI22_X1 U22328 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n20137), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n20142), .ZN(n20138) );
  OAI21_X1 U22329 ( .B1(n20570), .B2(n20139), .A(n20138), .ZN(P3_U2796) );
  AOI22_X1 U22330 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20143), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n20140), .ZN(n20141) );
  OAI21_X1 U22331 ( .B1(n20719), .B2(n20145), .A(n20141), .ZN(P3_U2797) );
  AOI22_X1 U22332 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n20143), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n20142), .ZN(n20144) );
  OAI21_X1 U22333 ( .B1(n20726), .B2(n20145), .A(n20144), .ZN(P3_U2798) );
  NAND2_X1 U22334 ( .A1(n20146), .A2(n20775), .ZN(n20753) );
  INV_X1 U22335 ( .A(n20550), .ZN(n20154) );
  AOI22_X1 U22336 ( .A1(n20546), .A2(n20147), .B1(P3_REIP_REG_1__SCAN_IN), 
        .B2(n20552), .ZN(n20153) );
  NOR2_X1 U22337 ( .A1(n21229), .A2(n20332), .ZN(n20314) );
  INV_X1 U22338 ( .A(n20314), .ZN(n20218) );
  OAI21_X1 U22339 ( .B1(n20553), .B2(n20218), .A(n20537), .ZN(n20151) );
  NOR2_X1 U22340 ( .A1(n21229), .A2(n10967), .ZN(n20300) );
  NOR2_X1 U22341 ( .A1(n21229), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n20301) );
  NOR2_X1 U22342 ( .A1(n20300), .A2(n20301), .ZN(n20249) );
  INV_X1 U22343 ( .A(n20249), .ZN(n20213) );
  OAI22_X1 U22344 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n20549), .B1(n20525), 
        .B2(n20148), .ZN(n20149) );
  AOI221_X1 U22345 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20151), .C1(
        n20150), .C2(n20213), .A(n20149), .ZN(n20152) );
  OAI211_X1 U22346 ( .C1(n20753), .C2(n20154), .A(n20153), .B(n20152), .ZN(
        P3_U2670) );
  INV_X1 U22347 ( .A(n20300), .ZN(n20347) );
  INV_X1 U22348 ( .A(n20775), .ZN(n20765) );
  OAI21_X1 U22349 ( .B1(n20765), .B2(n20764), .A(n20155), .ZN(n20768) );
  NOR2_X1 U22350 ( .A1(n20156), .A2(n20826), .ZN(n20170) );
  AOI211_X1 U22351 ( .C1(n20156), .C2(n20826), .A(n20170), .B(n20549), .ZN(
        n20159) );
  OAI22_X1 U22352 ( .A1(n20157), .A2(n20537), .B1(n20156), .B2(n20548), .ZN(
        n20158) );
  AOI211_X1 U22353 ( .C1(n20550), .C2(n20768), .A(n20159), .B(n20158), .ZN(
        n20167) );
  INV_X1 U22354 ( .A(n20168), .ZN(n20161) );
  OAI21_X1 U22355 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20160), .A(
        n10967), .ZN(n20171) );
  AOI211_X1 U22356 ( .C1(n20161), .C2(n20312), .A(n21229), .B(n20171), .ZN(
        n20165) );
  INV_X1 U22357 ( .A(n20162), .ZN(n20163) );
  AOI211_X1 U22358 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n20163), .A(n20176), .B(
        n20508), .ZN(n20164) );
  AOI211_X1 U22359 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n20547), .A(n20165), .B(
        n20164), .ZN(n20166) );
  OAI211_X1 U22360 ( .C1(n20168), .C2(n20347), .A(n20167), .B(n20166), .ZN(
        P3_U2669) );
  AOI22_X1 U22361 ( .A1(n20547), .A2(P3_EBX_REG_3__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n20450), .ZN(n20180) );
  NAND2_X1 U22362 ( .A1(n20182), .A2(n20440), .ZN(n20173) );
  INV_X1 U22363 ( .A(n20173), .ZN(n20169) );
  NOR2_X1 U22364 ( .A1(n20759), .A2(n20764), .ZN(n20781) );
  AOI21_X1 U22365 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20781), .A(
        n20795), .ZN(n20783) );
  OR2_X1 U22366 ( .A1(n17497), .A2(n20783), .ZN(n20792) );
  AOI22_X1 U22367 ( .A1(n20170), .A2(n20169), .B1(n20550), .B2(n20792), .ZN(
        n20179) );
  INV_X1 U22368 ( .A(n21229), .ZN(n20542) );
  XNOR2_X1 U22369 ( .A(n20172), .B(n20171), .ZN(n20174) );
  NAND2_X1 U22370 ( .A1(n20548), .A2(n20173), .ZN(n20185) );
  AOI22_X1 U22371 ( .A1(n20542), .A2(n20174), .B1(P3_REIP_REG_3__SCAN_IN), 
        .B2(n20185), .ZN(n20178) );
  OAI211_X1 U22372 ( .C1(n20176), .C2(n20175), .A(n20546), .B(n20183), .ZN(
        n20177) );
  NAND4_X1 U22373 ( .A1(n20180), .A2(n20179), .A3(n20178), .A4(n20177), .ZN(
        P3_U2668) );
  AOI22_X1 U22374 ( .A1(n20547), .A2(P3_EBX_REG_4__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n20450), .ZN(n20195) );
  AOI221_X1 U22375 ( .B1(n20181), .B2(n20550), .C1(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n20550), .A(n21167), .ZN(
        n20194) );
  NOR2_X1 U22376 ( .A1(n20549), .A2(n20182), .ZN(n20187) );
  AOI211_X1 U22377 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n20183), .A(n20203), .B(
        n20508), .ZN(n20184) );
  AOI221_X1 U22378 ( .B1(n20187), .B2(n20186), .C1(n20185), .C2(
        P3_REIP_REG_4__SCAN_IN), .A(n20184), .ZN(n20193) );
  INV_X1 U22379 ( .A(n20301), .ZN(n20348) );
  OAI21_X1 U22380 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n20348), .A(
        n20347), .ZN(n20190) );
  OAI21_X1 U22381 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20188), .A(
        n10967), .ZN(n20197) );
  OAI21_X1 U22382 ( .B1(n21229), .B2(n20197), .A(n20191), .ZN(n20189) );
  OAI21_X1 U22383 ( .B1(n20191), .B2(n20190), .A(n20189), .ZN(n20192) );
  NAND4_X1 U22384 ( .A1(n20195), .A2(n20194), .A3(n20193), .A4(n20192), .ZN(
        P3_U2667) );
  AOI21_X1 U22385 ( .B1(n20440), .B2(n20196), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n20200) );
  AOI21_X1 U22386 ( .B1(n20440), .B2(n20207), .A(n20552), .ZN(n20224) );
  XNOR2_X1 U22387 ( .A(n20198), .B(n20197), .ZN(n20199) );
  OAI22_X1 U22388 ( .A1(n20200), .A2(n20224), .B1(n21229), .B2(n20199), .ZN(
        n20201) );
  AOI211_X1 U22389 ( .C1(n20547), .C2(P3_EBX_REG_5__SCAN_IN), .A(n21167), .B(
        n20201), .ZN(n20205) );
  OAI211_X1 U22390 ( .C1(n20203), .C2(n20202), .A(n20546), .B(n20209), .ZN(
        n20204) );
  OAI211_X1 U22391 ( .C1(n20537), .C2(n20206), .A(n20205), .B(n20204), .ZN(
        P3_U2666) );
  OAI21_X1 U22392 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20219), .A(
        n20208), .ZN(n20217) );
  NOR3_X1 U22393 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n20549), .A3(n20207), .ZN(
        n20222) );
  AOI211_X1 U22394 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n20450), .A(
        n21167), .B(n20222), .ZN(n20216) );
  AOI21_X1 U22395 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n20347), .A(
        n20208), .ZN(n20214) );
  AOI211_X1 U22396 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n20209), .A(n20232), .B(
        n20508), .ZN(n20212) );
  INV_X1 U22397 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n20210) );
  OAI22_X1 U22398 ( .A1(n20525), .A2(n20210), .B1(n20875), .B2(n20224), .ZN(
        n20211) );
  AOI211_X1 U22399 ( .C1(n20214), .C2(n20213), .A(n20212), .B(n20211), .ZN(
        n20215) );
  OAI211_X1 U22400 ( .C1(n20218), .C2(n20217), .A(n20216), .B(n20215), .ZN(
        P3_U2665) );
  OAI21_X1 U22401 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20219), .A(
        n10967), .ZN(n20220) );
  XNOR2_X1 U22402 ( .A(n20221), .B(n20220), .ZN(n20230) );
  INV_X1 U22403 ( .A(n20222), .ZN(n20223) );
  AOI21_X1 U22404 ( .B1(n20224), .B2(n20223), .A(n20225), .ZN(n20229) );
  NAND3_X1 U22405 ( .A1(n20440), .A2(n20226), .A3(n20225), .ZN(n20227) );
  OAI211_X1 U22406 ( .C1(n20525), .C2(n20231), .A(n21176), .B(n20227), .ZN(
        n20228) );
  AOI211_X1 U22407 ( .C1(n20542), .C2(n20230), .A(n20229), .B(n20228), .ZN(
        n20234) );
  OAI211_X1 U22408 ( .C1(n20232), .C2(n20231), .A(n20546), .B(n20241), .ZN(
        n20233) );
  OAI211_X1 U22409 ( .C1(n20537), .C2(n20235), .A(n20234), .B(n20233), .ZN(
        P3_U2664) );
  OAI21_X1 U22410 ( .B1(n20236), .B2(n20312), .A(n10967), .ZN(n20237) );
  XNOR2_X1 U22411 ( .A(n20238), .B(n20237), .ZN(n20248) );
  OAI21_X1 U22412 ( .B1(n20257), .B2(n20549), .A(n20548), .ZN(n20272) );
  OAI21_X1 U22413 ( .B1(n20549), .B2(n20240), .A(n20239), .ZN(n20246) );
  AOI211_X1 U22414 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n20241), .A(n20251), .B(
        n20508), .ZN(n20245) );
  OAI22_X1 U22415 ( .A1(n20525), .A2(n20243), .B1(n20242), .B2(n20537), .ZN(
        n20244) );
  AOI211_X1 U22416 ( .C1(n20272), .C2(n20246), .A(n20245), .B(n20244), .ZN(
        n20247) );
  OAI211_X1 U22417 ( .C1(n20248), .C2(n21229), .A(n20247), .B(n21176), .ZN(
        P3_U2663) );
  AOI22_X1 U22418 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n20450), .B1(
        P3_REIP_REG_9__SCAN_IN), .B2(n20272), .ZN(n20261) );
  NOR2_X1 U22419 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n20549), .ZN(n20273) );
  AOI211_X1 U22420 ( .C1(n20250), .C2(n20347), .A(n20249), .B(n20258), .ZN(
        n20256) );
  AOI21_X1 U22421 ( .B1(n20546), .B2(n20251), .A(n20547), .ZN(n20254) );
  OR2_X1 U22422 ( .A1(n20508), .A2(n20251), .ZN(n20253) );
  AOI22_X1 U22423 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(n20254), .B1(n20253), .B2(
        n20252), .ZN(n20255) );
  AOI211_X1 U22424 ( .C1(n20257), .C2(n20273), .A(n20256), .B(n20255), .ZN(
        n20260) );
  OAI211_X1 U22425 ( .C1(n20312), .C2(n20265), .A(n20314), .B(n20258), .ZN(
        n20259) );
  NAND4_X1 U22426 ( .A1(n20261), .A2(n20260), .A3(n21176), .A4(n20259), .ZN(
        P3_U2662) );
  NOR2_X1 U22427 ( .A1(n20549), .A2(n20262), .ZN(n20279) );
  AOI22_X1 U22428 ( .A1(n20547), .A2(P3_EBX_REG_10__SCAN_IN), .B1(n20279), 
        .B2(n20263), .ZN(n20276) );
  OAI21_X1 U22429 ( .B1(n11138), .B2(n20312), .A(n10967), .ZN(n20277) );
  NOR2_X1 U22430 ( .A1(n20265), .A2(n20312), .ZN(n20266) );
  OAI21_X1 U22431 ( .B1(n20266), .B2(n20268), .A(n20542), .ZN(n20267) );
  AOI22_X1 U22432 ( .A1(n20268), .A2(n20277), .B1(n20347), .B2(n20267), .ZN(
        n20271) );
  AOI211_X1 U22433 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n20269), .A(n20284), .B(
        n20508), .ZN(n20270) );
  AOI211_X1 U22434 ( .C1(n20450), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n20271), .B(n20270), .ZN(n20275) );
  OAI21_X1 U22435 ( .B1(n20273), .B2(n20272), .A(P3_REIP_REG_10__SCAN_IN), 
        .ZN(n20274) );
  NAND4_X1 U22436 ( .A1(n20276), .A2(n20275), .A3(n21176), .A4(n20274), .ZN(
        P3_U2661) );
  AOI22_X1 U22437 ( .A1(n20547), .A2(P3_EBX_REG_11__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n20450), .ZN(n20287) );
  XNOR2_X1 U22438 ( .A(n20278), .B(n20277), .ZN(n20282) );
  OAI21_X1 U22439 ( .B1(n20290), .B2(n20549), .A(n20548), .ZN(n20288) );
  AOI21_X1 U22440 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n20279), .A(
        P3_REIP_REG_11__SCAN_IN), .ZN(n20280) );
  INV_X1 U22441 ( .A(n20280), .ZN(n20281) );
  AOI22_X1 U22442 ( .A1(n20542), .A2(n20282), .B1(n20288), .B2(n20281), .ZN(
        n20286) );
  OAI211_X1 U22443 ( .C1(n20284), .C2(n20283), .A(n20546), .B(n20289), .ZN(
        n20285) );
  NAND4_X1 U22444 ( .A1(n20287), .A2(n20286), .A3(n21176), .A4(n20285), .ZN(
        P3_U2660) );
  INV_X1 U22445 ( .A(n20288), .ZN(n20304) );
  AOI211_X1 U22446 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n20289), .A(n20305), .B(
        n20508), .ZN(n20293) );
  NAND3_X1 U22447 ( .A1(n20440), .A2(n20290), .A3(n20299), .ZN(n20303) );
  OAI211_X1 U22448 ( .C1(n20291), .C2(n20537), .A(n21176), .B(n20303), .ZN(
        n20292) );
  AOI211_X1 U22449 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n20547), .A(n20293), .B(
        n20292), .ZN(n20298) );
  OAI21_X1 U22450 ( .B1(n17795), .B2(n20312), .A(n10967), .ZN(n20295) );
  AOI21_X1 U22451 ( .B1(n20296), .B2(n20295), .A(n21229), .ZN(n20294) );
  OAI21_X1 U22452 ( .B1(n20296), .B2(n20295), .A(n20294), .ZN(n20297) );
  OAI211_X1 U22453 ( .C1(n20304), .C2(n20299), .A(n20298), .B(n20297), .ZN(
        P3_U2659) );
  AOI21_X1 U22454 ( .B1(n20302), .B2(n20301), .A(n20300), .ZN(n20318) );
  NOR2_X1 U22455 ( .A1(n20549), .A2(n20342), .ZN(n20311) );
  NAND2_X1 U22456 ( .A1(n20304), .A2(n20303), .ZN(n20310) );
  AOI21_X1 U22457 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n20450), .A(
        n21167), .ZN(n20307) );
  OAI211_X1 U22458 ( .C1(n20305), .C2(n20308), .A(n20546), .B(n20319), .ZN(
        n20306) );
  OAI211_X1 U22459 ( .C1(n20308), .C2(n20525), .A(n20307), .B(n20306), .ZN(
        n20309) );
  AOI221_X1 U22460 ( .B1(n20311), .B2(n20344), .C1(n20310), .C2(
        P3_REIP_REG_13__SCAN_IN), .A(n20309), .ZN(n20316) );
  OR3_X1 U22461 ( .A1(n17795), .A2(n20313), .A3(n20312), .ZN(n20330) );
  NAND3_X1 U22462 ( .A1(n20314), .A2(n20317), .A3(n20330), .ZN(n20315) );
  OAI211_X1 U22463 ( .C1(n20318), .C2(n20317), .A(n20316), .B(n20315), .ZN(
        P3_U2658) );
  AOI211_X1 U22464 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n20319), .A(n20337), .B(
        n20508), .ZN(n20328) );
  OAI21_X1 U22465 ( .B1(n20549), .B2(n20320), .A(n20548), .ZN(n20321) );
  INV_X1 U22466 ( .A(n20321), .ZN(n20364) );
  NOR3_X1 U22467 ( .A1(n20549), .A2(n20344), .A3(n20342), .ZN(n20322) );
  NOR2_X1 U22468 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n20322), .ZN(n20326) );
  NAND2_X1 U22469 ( .A1(n10967), .A2(n20330), .ZN(n20323) );
  XOR2_X1 U22470 ( .A(n20324), .B(n20323), .Z(n20325) );
  OAI22_X1 U22471 ( .A1(n20364), .A2(n20326), .B1(n21229), .B2(n20325), .ZN(
        n20327) );
  AOI211_X1 U22472 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n20547), .A(n20328), .B(
        n20327), .ZN(n20329) );
  OAI211_X1 U22473 ( .C1(n20331), .C2(n20537), .A(n20329), .B(n21176), .ZN(
        P3_U2657) );
  NOR2_X1 U22474 ( .A1(n20331), .A2(n20330), .ZN(n20350) );
  OR2_X1 U22475 ( .A1(n20350), .A2(n20332), .ZN(n20334) );
  OAI21_X1 U22476 ( .B1(n20335), .B2(n20334), .A(n20542), .ZN(n20333) );
  AOI21_X1 U22477 ( .B1(n20335), .B2(n20334), .A(n20333), .ZN(n20341) );
  OAI211_X1 U22478 ( .C1(n20337), .C2(n20336), .A(n20546), .B(n20353), .ZN(
        n20338) );
  OAI211_X1 U22479 ( .C1(n20339), .C2(n20537), .A(n21176), .B(n20338), .ZN(
        n20340) );
  AOI211_X1 U22480 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n20547), .A(n20341), .B(
        n20340), .ZN(n20345) );
  NOR4_X1 U22481 ( .A1(n20549), .A2(n20344), .A3(n20343), .A4(n20342), .ZN(
        n20352) );
  NAND2_X1 U22482 ( .A1(n20352), .A2(n20346), .ZN(n20363) );
  OAI211_X1 U22483 ( .C1(n20364), .C2(n20346), .A(n20345), .B(n20363), .ZN(
        P3_U2656) );
  OAI21_X1 U22484 ( .B1(n20349), .B2(n20348), .A(n20347), .ZN(n20360) );
  NAND2_X1 U22485 ( .A1(n20351), .A2(n20350), .ZN(n20382) );
  NAND2_X1 U22486 ( .A1(n10967), .A2(n20382), .ZN(n20368) );
  NOR3_X1 U22487 ( .A1(n20361), .A2(n21229), .A3(n20368), .ZN(n20359) );
  AND3_X1 U22488 ( .A1(n20365), .A2(P3_REIP_REG_15__SCAN_IN), .A3(n20352), 
        .ZN(n20355) );
  AOI211_X1 U22489 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n20353), .A(n20372), .B(
        n20508), .ZN(n20354) );
  AOI211_X1 U22490 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n20547), .A(n20355), .B(
        n20354), .ZN(n20356) );
  OAI211_X1 U22491 ( .C1(n20357), .C2(n20537), .A(n20356), .B(n21176), .ZN(
        n20358) );
  AOI211_X1 U22492 ( .C1(n20361), .C2(n20360), .A(n20359), .B(n20358), .ZN(
        n20362) );
  OAI221_X1 U22493 ( .B1(n20365), .B2(n20364), .C1(n20365), .C2(n20363), .A(
        n20362), .ZN(P3_U2655) );
  OAI21_X1 U22494 ( .B1(n20381), .B2(n20549), .A(n20548), .ZN(n20396) );
  OAI21_X1 U22495 ( .B1(n20549), .B2(n20367), .A(n20366), .ZN(n20376) );
  INV_X1 U22496 ( .A(n20368), .ZN(n20370) );
  OAI221_X1 U22497 ( .B1(n20371), .B2(n20370), .C1(n20369), .C2(n20368), .A(
        n20542), .ZN(n20374) );
  OAI211_X1 U22498 ( .C1(n20372), .C2(n20378), .A(n20546), .B(n20379), .ZN(
        n20373) );
  OAI211_X1 U22499 ( .C1(n20537), .C2(n11133), .A(n20374), .B(n20373), .ZN(
        n20375) );
  AOI21_X1 U22500 ( .B1(n20396), .B2(n20376), .A(n20375), .ZN(n20377) );
  OAI211_X1 U22501 ( .C1(n20525), .C2(n20378), .A(n20377), .B(n21176), .ZN(
        P3_U2654) );
  AOI211_X1 U22502 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n20379), .A(n20389), .B(
        n20508), .ZN(n20380) );
  AOI21_X1 U22503 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n20547), .A(n20380), .ZN(
        n20388) );
  NOR2_X1 U22504 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n20549), .ZN(n20395) );
  AOI22_X1 U22505 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n20450), .B1(
        n20381), .B2(n20395), .ZN(n20387) );
  OAI21_X1 U22506 ( .B1(n11133), .B2(n20382), .A(n10967), .ZN(n20383) );
  XOR2_X1 U22507 ( .A(n20384), .B(n20383), .Z(n20385) );
  AOI22_X1 U22508 ( .A1(n20542), .A2(n20385), .B1(P3_REIP_REG_18__SCAN_IN), 
        .B2(n20396), .ZN(n20386) );
  NAND4_X1 U22509 ( .A1(n20388), .A2(n20387), .A3(n20386), .A4(n21176), .ZN(
        P3_U2653) );
  AOI22_X1 U22510 ( .A1(n20547), .A2(P3_EBX_REG_19__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n20450), .ZN(n20403) );
  OAI21_X1 U22511 ( .B1(n20390), .B2(n20389), .A(n20546), .ZN(n20391) );
  INV_X1 U22512 ( .A(n20391), .ZN(n20394) );
  NOR3_X1 U22513 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n20549), .A3(n20392), 
        .ZN(n20393) );
  AOI211_X1 U22514 ( .C1(n20394), .C2(n20405), .A(n21167), .B(n20393), .ZN(
        n20402) );
  OAI21_X1 U22515 ( .B1(n20396), .B2(n20395), .A(P3_REIP_REG_19__SCAN_IN), 
        .ZN(n20401) );
  OAI211_X1 U22516 ( .C1(n20399), .C2(n20398), .A(n20542), .B(n20397), .ZN(
        n20400) );
  NAND4_X1 U22517 ( .A1(n20403), .A2(n20402), .A3(n20401), .A4(n20400), .ZN(
        P3_U2652) );
  AOI22_X1 U22518 ( .A1(n20547), .A2(P3_EBX_REG_20__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20450), .ZN(n20413) );
  OAI21_X1 U22519 ( .B1(n20404), .B2(n20549), .A(n20548), .ZN(n20431) );
  AND2_X1 U22520 ( .A1(n20440), .A2(n20414), .ZN(n20407) );
  AOI211_X1 U22521 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n20405), .A(n20419), .B(
        n20508), .ZN(n20406) );
  AOI221_X1 U22522 ( .B1(P3_REIP_REG_20__SCAN_IN), .B2(n20431), .C1(n20407), 
        .C2(n20431), .A(n20406), .ZN(n20412) );
  OAI211_X1 U22523 ( .C1(n20410), .C2(n20409), .A(n20542), .B(n20408), .ZN(
        n20411) );
  NAND3_X1 U22524 ( .A1(n20413), .A2(n20412), .A3(n20411), .ZN(P3_U2651) );
  AOI22_X1 U22525 ( .A1(n20547), .A2(P3_EBX_REG_21__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n20450), .ZN(n20423) );
  NAND3_X1 U22526 ( .A1(n20440), .A2(P3_REIP_REG_20__SCAN_IN), .A3(n20414), 
        .ZN(n20424) );
  NOR2_X1 U22527 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n20424), .ZN(n20432) );
  AOI21_X1 U22528 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n20431), .A(n20432), 
        .ZN(n20422) );
  OAI211_X1 U22529 ( .C1(n20417), .C2(n20416), .A(n20542), .B(n20415), .ZN(
        n20421) );
  OAI211_X1 U22530 ( .C1(n20419), .C2(n20418), .A(n20546), .B(n20426), .ZN(
        n20420) );
  NAND4_X1 U22531 ( .A1(n20423), .A2(n20422), .A3(n20421), .A4(n20420), .ZN(
        P3_U2650) );
  NOR2_X1 U22532 ( .A1(n20425), .A2(n20424), .ZN(n20441) );
  AOI211_X1 U22533 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n20426), .A(n20445), .B(
        n20508), .ZN(n20429) );
  AOI22_X1 U22534 ( .A1(n20547), .A2(P3_EBX_REG_22__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20450), .ZN(n20427) );
  INV_X1 U22535 ( .A(n20427), .ZN(n20428) );
  AOI211_X1 U22536 ( .C1(n20441), .C2(n20430), .A(n20429), .B(n20428), .ZN(
        n20438) );
  OAI21_X1 U22537 ( .B1(n20432), .B2(n20431), .A(P3_REIP_REG_22__SCAN_IN), 
        .ZN(n20437) );
  OAI211_X1 U22538 ( .C1(n20435), .C2(n20434), .A(n20542), .B(n20433), .ZN(
        n20436) );
  NAND3_X1 U22539 ( .A1(n20438), .A2(n20437), .A3(n20436), .ZN(P3_U2649) );
  AOI21_X1 U22540 ( .B1(n20440), .B2(n20439), .A(n20552), .ZN(n20467) );
  AOI21_X1 U22541 ( .B1(P3_REIP_REG_22__SCAN_IN), .B2(n20441), .A(
        P3_REIP_REG_23__SCAN_IN), .ZN(n20452) );
  OAI211_X1 U22542 ( .C1(n20444), .C2(n20443), .A(n20542), .B(n20442), .ZN(
        n20447) );
  OAI211_X1 U22543 ( .C1(n20445), .C2(n20448), .A(n20546), .B(n20453), .ZN(
        n20446) );
  OAI211_X1 U22544 ( .C1(n20448), .C2(n20525), .A(n20447), .B(n20446), .ZN(
        n20449) );
  AOI21_X1 U22545 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n20450), .A(
        n20449), .ZN(n20451) );
  OAI21_X1 U22546 ( .B1(n20467), .B2(n20452), .A(n20451), .ZN(P3_U2648) );
  NOR2_X1 U22547 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n20549), .ZN(n20459) );
  AOI211_X1 U22548 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n20453), .A(n20474), .B(
        n20508), .ZN(n20457) );
  OAI22_X1 U22549 ( .A1(n20525), .A2(n20455), .B1(n20454), .B2(n20537), .ZN(
        n20456) );
  AOI211_X1 U22550 ( .C1(n20459), .C2(n20458), .A(n20457), .B(n20456), .ZN(
        n20464) );
  OAI211_X1 U22551 ( .C1(n20462), .C2(n20461), .A(n20542), .B(n20460), .ZN(
        n20463) );
  OAI211_X1 U22552 ( .C1(n20467), .C2(n20465), .A(n20464), .B(n20463), .ZN(
        P3_U2647) );
  NOR2_X1 U22553 ( .A1(n20549), .A2(n20466), .ZN(n20472) );
  OAI21_X1 U22554 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n20549), .A(n20467), 
        .ZN(n20470) );
  OAI22_X1 U22555 ( .A1(n20525), .A2(n20473), .B1(n20468), .B2(n20537), .ZN(
        n20469) );
  AOI221_X1 U22556 ( .B1(n20472), .B2(n20471), .C1(n20470), .C2(
        P3_REIP_REG_25__SCAN_IN), .A(n20469), .ZN(n20480) );
  OAI211_X1 U22557 ( .C1(n20474), .C2(n20473), .A(n20546), .B(n20481), .ZN(
        n20479) );
  OAI211_X1 U22558 ( .C1(n20477), .C2(n20476), .A(n20542), .B(n20475), .ZN(
        n20478) );
  NAND3_X1 U22559 ( .A1(n20480), .A2(n20479), .A3(n20478), .ZN(P3_U2646) );
  INV_X1 U22560 ( .A(n20505), .ZN(n20494) );
  AOI211_X1 U22561 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n20481), .A(n20498), .B(
        n20508), .ZN(n20487) );
  INV_X1 U22562 ( .A(n20482), .ZN(n20484) );
  OAI22_X1 U22563 ( .A1(n20485), .A2(n20537), .B1(n20484), .B2(n20483), .ZN(
        n20486) );
  AOI211_X1 U22564 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n20547), .A(n20487), .B(
        n20486), .ZN(n20492) );
  OAI211_X1 U22565 ( .C1(n20490), .C2(n20489), .A(n20542), .B(n20488), .ZN(
        n20491) );
  OAI211_X1 U22566 ( .C1(n20494), .C2(n20493), .A(n20492), .B(n20491), .ZN(
        P3_U2645) );
  OAI22_X1 U22567 ( .A1(n20525), .A2(n20497), .B1(n20495), .B2(n20537), .ZN(
        n20496) );
  AOI221_X1 U22568 ( .B1(n20507), .B2(n20506), .C1(n20505), .C2(
        P3_REIP_REG_27__SCAN_IN), .A(n20496), .ZN(n20504) );
  OAI211_X1 U22569 ( .C1(n20498), .C2(n20497), .A(n20546), .B(n20509), .ZN(
        n20503) );
  OAI211_X1 U22570 ( .C1(n20501), .C2(n20500), .A(n20542), .B(n20499), .ZN(
        n20502) );
  NAND3_X1 U22571 ( .A1(n20504), .A2(n20503), .A3(n20502), .ZN(P3_U2644) );
  AOI21_X1 U22572 ( .B1(n20507), .B2(n20506), .A(n20505), .ZN(n20520) );
  AOI211_X1 U22573 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n20509), .A(n20521), .B(
        n20508), .ZN(n20513) );
  OAI22_X1 U22574 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n20511), .B1(n20537), 
        .B2(n20510), .ZN(n20512) );
  AOI211_X1 U22575 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n20547), .A(n20513), .B(
        n20512), .ZN(n20518) );
  OAI211_X1 U22576 ( .C1(n20516), .C2(n20515), .A(n20542), .B(n20514), .ZN(
        n20517) );
  OAI211_X1 U22577 ( .C1(n20520), .C2(n20519), .A(n20518), .B(n20517), .ZN(
        P3_U2643) );
  NOR2_X1 U22578 ( .A1(n20521), .A2(n20524), .ZN(n20534) );
  NAND2_X1 U22579 ( .A1(n20546), .A2(n20522), .ZN(n20545) );
  OAI22_X1 U22580 ( .A1(n20525), .A2(n20524), .B1(n20523), .B2(n20537), .ZN(
        n20526) );
  AOI221_X1 U22581 ( .B1(n20529), .B2(n20528), .C1(n20527), .C2(
        P3_REIP_REG_29__SCAN_IN), .A(n20526), .ZN(n20533) );
  OAI211_X1 U22582 ( .C1(n20531), .C2(n20530), .A(n20542), .B(n20535), .ZN(
        n20532) );
  OAI211_X1 U22583 ( .C1(n20534), .C2(n20545), .A(n20533), .B(n20532), .ZN(
        P3_U2642) );
  OAI22_X1 U22584 ( .A1(n20539), .A2(n21037), .B1(n20538), .B2(n20537), .ZN(
        n20540) );
  OAI21_X1 U22585 ( .B1(n20547), .B2(n20543), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n20544) );
  NOR2_X1 U22586 ( .A1(n20547), .A2(n20546), .ZN(n20557) );
  NAND2_X1 U22587 ( .A1(n20549), .A2(n20548), .ZN(n20551) );
  AOI22_X1 U22588 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n20551), .B1(n20550), 
        .B2(n20748), .ZN(n20555) );
  OR3_X1 U22589 ( .A1(n20553), .A2(n20552), .A3(n20791), .ZN(n20554) );
  OAI211_X1 U22590 ( .C1(n20557), .C2(n20556), .A(n20555), .B(n20554), .ZN(
        P3_U2671) );
  NOR3_X1 U22591 ( .A1(n20559), .A2(n11096), .A3(n20558), .ZN(n20560) );
  INV_X1 U22592 ( .A(n20565), .ZN(n20590) );
  NAND2_X1 U22593 ( .A1(n20590), .A2(n20563), .ZN(n20610) );
  NAND2_X1 U22594 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .ZN(n20621) );
  NAND2_X1 U22595 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_10__SCAN_IN), 
        .ZN(n20576) );
  OR3_X1 U22596 ( .A1(n20661), .A2(n20728), .A3(n20576), .ZN(n20579) );
  NOR2_X1 U22597 ( .A1(n20620), .A2(n20579), .ZN(n20571) );
  INV_X1 U22598 ( .A(n20571), .ZN(n20566) );
  NOR2_X1 U22599 ( .A1(n20621), .A2(n20566), .ZN(n20715) );
  NOR2_X1 U22600 ( .A1(n20567), .A2(n20566), .ZN(n20574) );
  AOI21_X1 U22601 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n20736), .A(n20574), .ZN(
        n20569) );
  OAI222_X1 U22602 ( .A1(n20610), .A2(n20570), .B1(n20715), .B2(n20569), .C1(
        n20732), .C2(n20568), .ZN(P3_U2722) );
  AOI21_X1 U22603 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n20736), .A(n20571), .ZN(
        n20573) );
  OAI222_X1 U22604 ( .A1(n20610), .A2(n20575), .B1(n20574), .B2(n20573), .C1(
        n20732), .C2(n20572), .ZN(P3_U2723) );
  NAND2_X1 U22605 ( .A1(n20736), .A2(n20622), .ZN(n20582) );
  AOI22_X1 U22606 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20741), .B1(n20740), .B2(
        n20577), .ZN(n20578) );
  OAI221_X1 U22607 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n20579), .C1(n20620), 
        .C2(n20582), .A(n20578), .ZN(P3_U2724) );
  NOR2_X1 U22608 ( .A1(n20661), .A2(n20728), .ZN(n20585) );
  AOI21_X1 U22609 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n20585), .A(
        P3_EAX_REG_10__SCAN_IN), .ZN(n20581) );
  OAI222_X1 U22610 ( .A1(n20610), .A2(n20583), .B1(n20582), .B2(n20581), .C1(
        n20732), .C2(n20580), .ZN(P3_U2725) );
  NOR2_X1 U22611 ( .A1(n20728), .A2(n20584), .ZN(n20588) );
  AOI21_X1 U22612 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n20736), .A(n20585), .ZN(
        n20587) );
  OAI222_X1 U22613 ( .A1(n20610), .A2(n20589), .B1(n20588), .B2(n20587), .C1(
        n20732), .C2(n20586), .ZN(P3_U2726) );
  NAND2_X1 U22614 ( .A1(n20722), .A2(n20590), .ZN(n20743) );
  NOR2_X1 U22615 ( .A1(n20614), .A2(n20615), .ZN(n20606) );
  NAND2_X1 U22616 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n20609), .ZN(n20596) );
  NOR2_X1 U22617 ( .A1(n20592), .A2(n20596), .ZN(n20599) );
  AOI21_X1 U22618 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n20736), .A(n20599), .ZN(
        n20594) );
  OAI222_X1 U22619 ( .A1(n20610), .A2(n20595), .B1(n20729), .B2(n20594), .C1(
        n20732), .C2(n20593), .ZN(P3_U2728) );
  INV_X1 U22620 ( .A(n20596), .ZN(n20604) );
  AOI21_X1 U22621 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n20736), .A(n20604), .ZN(
        n20598) );
  OAI222_X1 U22622 ( .A1(n20600), .A2(n20610), .B1(n20599), .B2(n20598), .C1(
        n20732), .C2(n20597), .ZN(P3_U2729) );
  AOI21_X1 U22623 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n20736), .A(n20609), .ZN(
        n20603) );
  INV_X1 U22624 ( .A(n20601), .ZN(n20602) );
  OAI222_X1 U22625 ( .A1(n20605), .A2(n20610), .B1(n20604), .B2(n20603), .C1(
        n20732), .C2(n20602), .ZN(P3_U2730) );
  AOI21_X1 U22626 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n20736), .A(n20606), .ZN(
        n20608) );
  OAI222_X1 U22627 ( .A1(n20611), .A2(n20610), .B1(n20609), .B2(n20608), .C1(
        n20732), .C2(n20607), .ZN(P3_U2731) );
  NAND2_X1 U22628 ( .A1(n20736), .A2(n20615), .ZN(n20619) );
  AOI22_X1 U22629 ( .A1(n20741), .A2(BUF2_REG_3__SCAN_IN), .B1(n20740), .B2(
        n20612), .ZN(n20613) );
  OAI221_X1 U22630 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n20615), .C1(n20614), 
        .C2(n20619), .A(n20613), .ZN(P3_U2732) );
  AOI22_X1 U22631 ( .A1(n20741), .A2(BUF2_REG_2__SCAN_IN), .B1(n20740), .B2(
        n20616), .ZN(n20617) );
  OAI221_X1 U22632 ( .B1(n20619), .B2(n20735), .C1(n20619), .C2(n20618), .A(
        n20617), .ZN(P3_U2733) );
  INV_X1 U22633 ( .A(n20721), .ZN(n20716) );
  NAND2_X1 U22634 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n20646), .ZN(n20642) );
  NAND2_X1 U22635 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n20631), .ZN(n20637) );
  NAND2_X1 U22636 ( .A1(n20736), .A2(n20637), .ZN(n20635) );
  NOR2_X2 U22637 ( .A1(n20624), .A2(n20736), .ZN(n20709) );
  NAND2_X1 U22638 ( .A1(n20625), .A2(n20690), .ZN(n20707) );
  OAI22_X1 U22639 ( .A1(n20627), .A2(n20732), .B1(n20626), .B2(n20707), .ZN(
        n20628) );
  AOI21_X1 U22640 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n20709), .A(n20628), .ZN(
        n20629) );
  OAI221_X1 U22641 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n20637), .C1(n20638), 
        .C2(n20635), .A(n20629), .ZN(P3_U2714) );
  AOI22_X1 U22642 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n20708), .B1(n20740), .B2(
        n20630), .ZN(n20633) );
  AOI22_X1 U22643 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n20709), .B1(n20631), .B2(
        n20660), .ZN(n20632) );
  OAI211_X1 U22644 ( .C1(n20660), .C2(n20635), .A(n20633), .B(n20632), .ZN(
        P3_U2715) );
  AOI22_X1 U22645 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n20708), .B1(n20740), .B2(
        n20634), .ZN(n20641) );
  OAI21_X1 U22646 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n20743), .A(n20635), .ZN(
        n20636) );
  AOI22_X1 U22647 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n20709), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n20636), .ZN(n20640) );
  OR3_X1 U22648 ( .A1(n20638), .A2(n20637), .A3(P3_EAX_REG_22__SCAN_IN), .ZN(
        n20639) );
  NAND3_X1 U22649 ( .A1(n20641), .A2(n20640), .A3(n20639), .ZN(P3_U2713) );
  AOI22_X1 U22650 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n20709), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n20708), .ZN(n20644) );
  OAI211_X1 U22651 ( .C1(n20646), .C2(P3_EAX_REG_19__SCAN_IN), .A(n20736), .B(
        n20642), .ZN(n20643) );
  OAI211_X1 U22652 ( .C1(n20645), .C2(n20732), .A(n20644), .B(n20643), .ZN(
        P3_U2716) );
  AOI22_X1 U22653 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n20709), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n20708), .ZN(n20650) );
  AOI211_X1 U22654 ( .C1(n20647), .C2(n20652), .A(n20646), .B(n20690), .ZN(
        n20648) );
  INV_X1 U22655 ( .A(n20648), .ZN(n20649) );
  OAI211_X1 U22656 ( .C1(n20651), .C2(n20732), .A(n20650), .B(n20649), .ZN(
        P3_U2717) );
  AOI22_X1 U22657 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n20709), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n20708), .ZN(n20655) );
  INV_X1 U22658 ( .A(n20710), .ZN(n20653) );
  OAI211_X1 U22659 ( .C1(n20653), .C2(P3_EAX_REG_17__SCAN_IN), .A(n20736), .B(
        n20652), .ZN(n20654) );
  OAI211_X1 U22660 ( .C1(n20656), .C2(n20732), .A(n20655), .B(n20654), .ZN(
        P3_U2718) );
  AOI22_X1 U22661 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n20708), .B1(n20740), .B2(
        n20657), .ZN(n20658) );
  INV_X1 U22662 ( .A(n20658), .ZN(n20664) );
  AOI211_X1 U22663 ( .C1(n20662), .C2(n20696), .A(n11013), .B(n20690), .ZN(
        n20663) );
  AOI211_X1 U22664 ( .C1(n20709), .C2(BUF2_REG_9__SCAN_IN), .A(n20664), .B(
        n20663), .ZN(n20665) );
  INV_X1 U22665 ( .A(n20665), .ZN(P3_U2710) );
  AOI22_X1 U22666 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n20709), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n20708), .ZN(n20667) );
  OAI211_X1 U22667 ( .C1(n11013), .C2(P3_EAX_REG_26__SCAN_IN), .A(n20736), .B(
        n20688), .ZN(n20666) );
  OAI211_X1 U22668 ( .C1(n20668), .C2(n20732), .A(n20667), .B(n20666), .ZN(
        P3_U2709) );
  NAND2_X1 U22669 ( .A1(n20687), .A2(P3_EAX_REG_28__SCAN_IN), .ZN(n20683) );
  NOR2_X2 U22670 ( .A1(n20683), .A2(n20677), .ZN(n20676) );
  NAND2_X1 U22671 ( .A1(n20676), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n20672) );
  AND2_X1 U22672 ( .A1(n20708), .A2(BUF2_REG_31__SCAN_IN), .ZN(n20669) );
  OAI21_X1 U22673 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n20672), .A(n20671), .ZN(
        P3_U2704) );
  AOI22_X1 U22674 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20709), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n20708), .ZN(n20674) );
  OAI211_X1 U22675 ( .C1(n20676), .C2(P3_EAX_REG_30__SCAN_IN), .A(n20736), .B(
        n20672), .ZN(n20673) );
  OAI211_X1 U22676 ( .C1(n20675), .C2(n20732), .A(n20674), .B(n20673), .ZN(
        P3_U2705) );
  INV_X1 U22677 ( .A(n20676), .ZN(n20679) );
  OAI21_X1 U22678 ( .B1(n20690), .B2(n20677), .A(n20683), .ZN(n20678) );
  AOI22_X1 U22679 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n20708), .B1(n20679), .B2(
        n20678), .ZN(n20682) );
  AOI22_X1 U22680 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n20709), .B1(n20740), .B2(
        n20680), .ZN(n20681) );
  NAND2_X1 U22681 ( .A1(n20682), .A2(n20681), .ZN(P3_U2706) );
  AOI22_X1 U22682 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n20709), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n20708), .ZN(n20685) );
  OAI211_X1 U22683 ( .C1(n20687), .C2(P3_EAX_REG_28__SCAN_IN), .A(n20736), .B(
        n20683), .ZN(n20684) );
  OAI211_X1 U22684 ( .C1(n20686), .C2(n20732), .A(n20685), .B(n20684), .ZN(
        P3_U2707) );
  INV_X1 U22685 ( .A(n20687), .ZN(n20692) );
  OAI21_X1 U22686 ( .B1(n20690), .B2(n20689), .A(n20688), .ZN(n20691) );
  AOI22_X1 U22687 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n20708), .B1(n20692), .B2(
        n20691), .ZN(n20695) );
  AOI22_X1 U22688 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n20709), .B1(n20740), .B2(
        n20693), .ZN(n20694) );
  NAND2_X1 U22689 ( .A1(n20695), .A2(n20694), .ZN(P3_U2708) );
  AOI22_X1 U22690 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20709), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n20708), .ZN(n20699) );
  OAI211_X1 U22691 ( .C1(n20697), .C2(P3_EAX_REG_24__SCAN_IN), .A(n20736), .B(
        n20696), .ZN(n20698) );
  OAI211_X1 U22692 ( .C1(n20700), .C2(n20732), .A(n20699), .B(n20698), .ZN(
        P3_U2711) );
  AOI22_X1 U22693 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n20709), .B1(n20740), .B2(
        n20701), .ZN(n20705) );
  OAI211_X1 U22694 ( .C1(n20703), .C2(P3_EAX_REG_23__SCAN_IN), .A(n20736), .B(
        n20702), .ZN(n20704) );
  OAI211_X1 U22695 ( .C1(n20707), .C2(n20706), .A(n20705), .B(n20704), .ZN(
        P3_U2712) );
  AOI22_X1 U22696 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n20709), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n20708), .ZN(n20713) );
  OAI211_X1 U22697 ( .C1(n20711), .C2(P3_EAX_REG_16__SCAN_IN), .A(n20736), .B(
        n20710), .ZN(n20712) );
  OAI211_X1 U22698 ( .C1(n20714), .C2(n20732), .A(n20713), .B(n20712), .ZN(
        P3_U2719) );
  INV_X1 U22699 ( .A(n20715), .ZN(n20720) );
  NAND2_X1 U22700 ( .A1(n20736), .A2(n20716), .ZN(n20725) );
  AOI22_X1 U22701 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n20741), .B1(n20740), .B2(
        n20717), .ZN(n20718) );
  OAI221_X1 U22702 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n20720), .C1(n20719), 
        .C2(n20725), .A(n20718), .ZN(P3_U2721) );
  NAND2_X1 U22703 ( .A1(n20722), .A2(n20721), .ZN(n20727) );
  AOI22_X1 U22704 ( .A1(n20740), .A2(n20723), .B1(BUF2_REG_15__SCAN_IN), .B2(
        n20741), .ZN(n20724) );
  OAI221_X1 U22705 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(n20727), .C1(n20726), 
        .C2(n20725), .A(n20724), .ZN(P3_U2720) );
  OAI211_X1 U22706 ( .C1(n20729), .C2(P3_EAX_REG_8__SCAN_IN), .A(n20736), .B(
        n20728), .ZN(n20731) );
  NAND2_X1 U22707 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n20741), .ZN(n20730) );
  OAI211_X1 U22708 ( .C1(n20733), .C2(n20732), .A(n20731), .B(n20730), .ZN(
        P3_U2727) );
  AOI22_X1 U22709 ( .A1(n20741), .A2(BUF2_REG_1__SCAN_IN), .B1(n20740), .B2(
        n20734), .ZN(n20738) );
  OAI211_X1 U22710 ( .C1(n20745), .C2(P3_EAX_REG_1__SCAN_IN), .A(n20736), .B(
        n20735), .ZN(n20737) );
  NAND2_X1 U22711 ( .A1(n20738), .A2(n20737), .ZN(P3_U2734) );
  AOI22_X1 U22712 ( .A1(n20741), .A2(BUF2_REG_0__SCAN_IN), .B1(n20740), .B2(
        n20739), .ZN(n20742) );
  OAI221_X1 U22713 ( .B1(n20745), .B2(n20744), .C1(n20745), .C2(n20743), .A(
        n20742), .ZN(P3_U2735) );
  NOR2_X1 U22714 ( .A1(n20746), .A2(n21171), .ZN(n20752) );
  AOI22_X1 U22715 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n21175), .B1(
        n20752), .B2(n20748), .ZN(n21205) );
  AOI222_X1 U22716 ( .A1(n20827), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n21205), 
        .B2(n20791), .C1(n20748), .C2(n21234), .ZN(n20747) );
  AOI22_X1 U22717 ( .A1(n20796), .A2(n20748), .B1(n20747), .B2(n20793), .ZN(
        P3_U3290) );
  AOI21_X1 U22718 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n21171), .A(
        n20749), .ZN(n20790) );
  NAND2_X1 U22719 ( .A1(n20790), .A2(n20750), .ZN(n20758) );
  INV_X1 U22720 ( .A(n20758), .ZN(n20751) );
  OAI22_X1 U22721 ( .A1(n20752), .A2(n20753), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n20751), .ZN(n21203) );
  INV_X1 U22722 ( .A(n20753), .ZN(n20756) );
  OAI22_X1 U22723 ( .A1(n20832), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n21052), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20771) );
  INV_X1 U22724 ( .A(n20771), .ZN(n20755) );
  NOR2_X1 U22725 ( .A1(n20754), .A2(n20827), .ZN(n20770) );
  AOI222_X1 U22726 ( .A1(n21203), .A2(n20791), .B1(n20756), .B2(n21234), .C1(
        n20755), .C2(n20770), .ZN(n20757) );
  AOI22_X1 U22727 ( .A1(n20796), .A2(n20759), .B1(n20757), .B2(n20793), .ZN(
        P3_U3289) );
  OAI221_X1 U22728 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C1(n20764), .C2(n20759), .A(
        n20758), .ZN(n20767) );
  INV_X1 U22729 ( .A(n20760), .ZN(n20830) );
  OAI22_X1 U22730 ( .A1(n20763), .A2(n20762), .B1(n20830), .B2(n20761), .ZN(
        n20784) );
  NOR2_X1 U22731 ( .A1(n20765), .A2(n20764), .ZN(n20772) );
  OAI21_X1 U22732 ( .B1(n20779), .B2(n20784), .A(n20772), .ZN(n20766) );
  OAI211_X1 U22733 ( .C1(n21119), .C2(n20768), .A(n20767), .B(n20766), .ZN(
        n21200) );
  AOI222_X1 U22734 ( .A1(n21200), .A2(n20791), .B1(n20771), .B2(n20770), .C1(
        n20769), .C2(n21234), .ZN(n20774) );
  AOI22_X1 U22735 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n20796), .B1(
        n21234), .B2(n20772), .ZN(n20773) );
  OAI21_X1 U22736 ( .B1(n20796), .B2(n20774), .A(n20773), .ZN(P3_U3288) );
  NOR2_X1 U22737 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20795), .ZN(
        n20780) );
  AOI211_X1 U22738 ( .C1(n20776), .C2(n20775), .A(n13934), .B(n21119), .ZN(
        n20778) );
  AOI22_X1 U22739 ( .A1(n20780), .A2(n20779), .B1(n20778), .B2(n20777), .ZN(
        n20788) );
  OR2_X1 U22740 ( .A1(n20830), .A2(n20831), .ZN(n20786) );
  OR2_X1 U22741 ( .A1(n20795), .A2(n20781), .ZN(n20782) );
  OAI21_X1 U22742 ( .B1(n20830), .B2(n20789), .A(n20782), .ZN(n20785) );
  AOI22_X1 U22743 ( .A1(n20786), .A2(n20785), .B1(n20784), .B2(n20783), .ZN(
        n20787) );
  OAI211_X1 U22744 ( .C1(n20790), .C2(n20789), .A(n20788), .B(n20787), .ZN(
        n21198) );
  AOI22_X1 U22745 ( .A1(n21234), .A2(n20792), .B1(n20791), .B2(n21198), .ZN(
        n20794) );
  AOI22_X1 U22746 ( .A1(n20796), .A2(n20795), .B1(n20794), .B2(n20793), .ZN(
        P3_U3285) );
  INV_X1 U22747 ( .A(n20797), .ZN(n20813) );
  NOR2_X1 U22748 ( .A1(n20973), .A2(n21080), .ZN(n21104) );
  NOR2_X1 U22749 ( .A1(n20827), .A2(n20904), .ZN(n21168) );
  OAI221_X1 U22750 ( .B1(n20951), .B2(n20798), .C1(n20951), .C2(n21168), .A(
        n21151), .ZN(n21088) );
  AOI21_X1 U22751 ( .B1(n20799), .B2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n21175), .ZN(n20800) );
  AOI21_X1 U22752 ( .B1(n21184), .B2(n20801), .A(n20800), .ZN(n21091) );
  INV_X1 U22753 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n21097) );
  AOI22_X1 U22754 ( .A1(n21184), .A2(n20806), .B1(n20903), .B2(n21097), .ZN(
        n20805) );
  AOI22_X1 U22755 ( .A1(n21183), .A2(n20803), .B1(n21067), .B2(n20802), .ZN(
        n20804) );
  NAND3_X1 U22756 ( .A1(n21091), .A2(n20805), .A3(n20804), .ZN(n20976) );
  AOI211_X1 U22757 ( .C1(n21171), .C2(n20806), .A(n21088), .B(n20976), .ZN(
        n20808) );
  NOR3_X1 U22758 ( .A1(n21167), .A2(n20808), .A3(n20807), .ZN(n20809) );
  AOI211_X1 U22759 ( .C1(n20811), .C2(n21104), .A(n20810), .B(n20809), .ZN(
        n20812) );
  OAI21_X1 U22760 ( .B1(n20813), .B2(n21144), .A(n20812), .ZN(P3_U2841) );
  NAND2_X1 U22761 ( .A1(n21151), .A2(n21183), .ZN(n20888) );
  INV_X1 U22762 ( .A(n20870), .ZN(n20893) );
  AND2_X1 U22763 ( .A1(n21137), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n20815) );
  NOR2_X1 U22764 ( .A1(n21184), .A2(n21171), .ZN(n21100) );
  AOI221_X1 U22765 ( .B1(n21100), .B2(n20827), .C1(n21175), .C2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n21080), .ZN(n20814) );
  AOI211_X1 U22766 ( .C1(n21062), .C2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n20815), .B(n20814), .ZN(n20816) );
  OAI221_X1 U22767 ( .B1(n20818), .B2(n20888), .C1(n20817), .C2(n20893), .A(
        n20816), .ZN(P3_U2862) );
  NOR2_X1 U22768 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n21100), .ZN(
        n20819) );
  AOI22_X1 U22769 ( .A1(n21183), .A2(n20820), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20819), .ZN(n20822) );
  OAI211_X1 U22770 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n20903), .A(
        n20832), .B(n21140), .ZN(n20821) );
  OAI211_X1 U22771 ( .C1(n20823), .C2(n21190), .A(n20822), .B(n20821), .ZN(
        n20824) );
  AOI22_X1 U22772 ( .A1(n21151), .A2(n20824), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n21062), .ZN(n20825) );
  OAI21_X1 U22773 ( .B1(n21176), .B2(n20826), .A(n20825), .ZN(P3_U2861) );
  NOR3_X1 U22774 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n20842), .A3(
        n20832), .ZN(n20837) );
  NOR2_X1 U22775 ( .A1(n20832), .A2(n20827), .ZN(n20828) );
  OAI221_X1 U22776 ( .B1(n20843), .B2(n20828), .C1(n20843), .C2(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(n21184), .ZN(n20834) );
  NOR2_X1 U22777 ( .A1(n20951), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n21115) );
  NOR3_X1 U22778 ( .A1(n20831), .A2(n20830), .A3(n20829), .ZN(n21112) );
  INV_X1 U22779 ( .A(n21112), .ZN(n21170) );
  OAI211_X1 U22780 ( .C1(n21115), .C2(n20832), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n21170), .ZN(n20833) );
  OAI211_X1 U22781 ( .C1(n20835), .C2(n21190), .A(n20834), .B(n20833), .ZN(
        n20836) );
  AOI211_X1 U22782 ( .C1(n20838), .C2(n21183), .A(n20837), .B(n20836), .ZN(
        n20841) );
  AOI21_X1 U22783 ( .B1(n21062), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n20839), .ZN(n20840) );
  OAI21_X1 U22784 ( .B1(n20841), .B2(n21080), .A(n20840), .ZN(P3_U2860) );
  AOI22_X1 U22785 ( .A1(n21137), .A2(P3_REIP_REG_3__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n21062), .ZN(n20850) );
  OAI22_X1 U22786 ( .A1(n21119), .A2(n20843), .B1(n20844), .B2(n20842), .ZN(
        n20853) );
  INV_X1 U22787 ( .A(n20853), .ZN(n20879) );
  AOI21_X1 U22788 ( .B1(n20879), .B2(n20865), .A(n21080), .ZN(n20847) );
  OAI21_X1 U22789 ( .B1(n21115), .B2(n20844), .A(n21170), .ZN(n20845) );
  OAI211_X1 U22790 ( .C1(n21119), .C2(n20846), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n20845), .ZN(n20852) );
  AOI22_X1 U22791 ( .A1(n21012), .A2(n20848), .B1(n20847), .B2(n20852), .ZN(
        n20849) );
  OAI211_X1 U22792 ( .C1(n20893), .C2(n20851), .A(n20850), .B(n20849), .ZN(
        P3_U2859) );
  NAND3_X1 U22793 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n21140), .A3(
        n20852), .ZN(n20855) );
  NAND3_X1 U22794 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n20866), .A3(
        n20853), .ZN(n20854) );
  OAI211_X1 U22795 ( .C1(n20856), .C2(n21190), .A(n20855), .B(n20854), .ZN(
        n20858) );
  AOI22_X1 U22796 ( .A1(n21151), .A2(n20858), .B1(n21012), .B2(n20857), .ZN(
        n20860) );
  NAND2_X1 U22797 ( .A1(n21137), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n20859) );
  OAI211_X1 U22798 ( .C1(n21074), .C2(n20866), .A(n20860), .B(n20859), .ZN(
        P3_U2858) );
  INV_X1 U22799 ( .A(n20861), .ZN(n20862) );
  AOI21_X1 U22800 ( .B1(n21184), .B2(n20862), .A(n21115), .ZN(n20883) );
  OAI211_X1 U22801 ( .C1(n20863), .C2(n21112), .A(n21151), .B(n20883), .ZN(
        n20864) );
  NAND2_X1 U22802 ( .A1(n21176), .A2(n20864), .ZN(n20874) );
  NOR4_X1 U22803 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20879), .A3(
        n20866), .A4(n20865), .ZN(n20867) );
  AOI22_X1 U22804 ( .A1(n21167), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n21151), 
        .B2(n20867), .ZN(n20872) );
  AOI22_X1 U22805 ( .A1(n20870), .A2(n20869), .B1(n21012), .B2(n20868), .ZN(
        n20871) );
  OAI211_X1 U22806 ( .C1(n20873), .C2(n20874), .A(n20872), .B(n20871), .ZN(
        P3_U2857) );
  OAI22_X1 U22807 ( .A1(n21176), .A2(n20875), .B1(n20884), .B2(n20874), .ZN(
        n20876) );
  AOI21_X1 U22808 ( .B1(n21012), .B2(n20877), .A(n20876), .ZN(n20881) );
  NOR2_X1 U22809 ( .A1(n20879), .A2(n20878), .ZN(n20886) );
  NAND3_X1 U22810 ( .A1(n21151), .A2(n20886), .A3(n20884), .ZN(n20880) );
  OAI211_X1 U22811 ( .C1(n20882), .C2(n20893), .A(n20881), .B(n20880), .ZN(
        P3_U2856) );
  OAI211_X1 U22812 ( .C1(n21174), .C2(n21112), .A(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B(n20883), .ZN(n20885) );
  OAI221_X1 U22813 ( .B1(n20885), .B2(n21184), .C1(n20885), .C2(n20884), .A(
        n21151), .ZN(n20894) );
  AOI21_X1 U22814 ( .B1(n21074), .B2(n20894), .A(n20898), .ZN(n20890) );
  NAND2_X1 U22815 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n20886), .ZN(
        n20913) );
  OAI22_X1 U22816 ( .A1(n20888), .A2(n20887), .B1(n20913), .B2(n20894), .ZN(
        n20889) );
  AOI211_X1 U22817 ( .C1(P3_REIP_REG_7__SCAN_IN), .C2(n21137), .A(n20890), .B(
        n20889), .ZN(n20891) );
  OAI21_X1 U22818 ( .B1(n20893), .B2(n20892), .A(n20891), .ZN(P3_U2855) );
  AOI221_X1 U22819 ( .B1(n21051), .B2(n21074), .C1(n20894), .C2(n21074), .A(
        n21172), .ZN(n20895) );
  AOI211_X1 U22820 ( .C1(n20897), .C2(n21012), .A(n20896), .B(n20895), .ZN(
        n20901) );
  NOR3_X1 U22821 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n20898), .A3(
        n20913), .ZN(n20899) );
  OAI221_X1 U22822 ( .B1(n20899), .B2(n21067), .C1(n20899), .C2(n20902), .A(
        n21151), .ZN(n20900) );
  OAI211_X1 U22823 ( .C1(n20902), .C2(n21144), .A(n20901), .B(n20900), .ZN(
        P3_U2854) );
  OAI21_X1 U22824 ( .B1(n20916), .B2(n20904), .A(n20903), .ZN(n20905) );
  OAI21_X1 U22825 ( .B1(n20923), .B2(n21119), .A(n20905), .ZN(n20925) );
  NAND2_X1 U22826 ( .A1(n21056), .A2(n21110), .ZN(n21117) );
  AOI21_X1 U22827 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n21168), .A(
        n20951), .ZN(n20910) );
  AOI22_X1 U22828 ( .A1(n21183), .A2(n20907), .B1(n21067), .B2(n20906), .ZN(
        n20909) );
  NAND2_X1 U22829 ( .A1(n21184), .A2(n20908), .ZN(n20954) );
  NAND3_X1 U22830 ( .A1(n20909), .A2(n21074), .A3(n20954), .ZN(n21178) );
  AOI211_X1 U22831 ( .C1(n20916), .C2(n21117), .A(n20910), .B(n21178), .ZN(
        n21158) );
  OAI21_X1 U22832 ( .B1(n20951), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n21158), .ZN(n20911) );
  OAI21_X1 U22833 ( .B1(n20925), .B2(n20911), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n20921) );
  INV_X1 U22834 ( .A(n20912), .ZN(n20914) );
  NOR2_X1 U22835 ( .A1(n20914), .A2(n20913), .ZN(n20956) );
  OR2_X1 U22836 ( .A1(n20956), .A2(n20915), .ZN(n20922) );
  NOR3_X1 U22837 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n20916), .A3(
        n21181), .ZN(n20917) );
  AOI21_X1 U22838 ( .B1(n21166), .B2(n20918), .A(n20917), .ZN(n20919) );
  OAI221_X1 U22839 ( .B1(n21167), .B2(n20921), .C1(n21176), .C2(n20920), .A(
        n20919), .ZN(P3_U2851) );
  AOI21_X1 U22840 ( .B1(n20923), .B2(n20922), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n20935) );
  INV_X1 U22841 ( .A(n20924), .ZN(n20926) );
  AOI21_X1 U22842 ( .B1(n21067), .B2(n20926), .A(n20925), .ZN(n20927) );
  OAI21_X1 U22843 ( .B1(n20928), .B2(n21056), .A(n20927), .ZN(n21145) );
  INV_X1 U22844 ( .A(n20954), .ZN(n20930) );
  AOI21_X1 U22845 ( .B1(n20929), .B2(n21168), .A(n20951), .ZN(n21146) );
  NOR2_X1 U22846 ( .A1(n20930), .A2(n21146), .ZN(n20940) );
  OAI211_X1 U22847 ( .C1(n21175), .C2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B(n20940), .ZN(n21148) );
  OAI21_X1 U22848 ( .B1(n21145), .B2(n21148), .A(n21151), .ZN(n20934) );
  AOI22_X1 U22849 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n21062), .B1(
        n21166), .B2(n20931), .ZN(n20933) );
  OAI211_X1 U22850 ( .C1(n20935), .C2(n20934), .A(n20933), .B(n20932), .ZN(
        P3_U2850) );
  NOR2_X1 U22851 ( .A1(n21175), .A2(n21113), .ZN(n21161) );
  OAI22_X1 U22852 ( .A1(n21175), .A2(n20957), .B1(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n21100), .ZN(n20936) );
  AOI211_X1 U22853 ( .C1(n21184), .C2(n20937), .A(n21161), .B(n20936), .ZN(
        n20939) );
  AOI21_X1 U22854 ( .B1(n20940), .B2(n20939), .A(n20938), .ZN(n20944) );
  NAND2_X1 U22855 ( .A1(n20957), .A2(n20956), .ZN(n20942) );
  OAI22_X1 U22856 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n20942), .B1(
        n21056), .B2(n20941), .ZN(n20943) );
  AOI211_X1 U22857 ( .C1(n21067), .C2(n20945), .A(n20944), .B(n20943), .ZN(
        n20949) );
  AOI22_X1 U22858 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n21062), .B1(
        n21166), .B2(n20946), .ZN(n20948) );
  OAI211_X1 U22859 ( .C1(n20949), .C2(n21080), .A(n20948), .B(n20947), .ZN(
        P3_U2848) );
  OR2_X1 U22860 ( .A1(n21056), .A2(n21108), .ZN(n20963) );
  AOI22_X1 U22861 ( .A1(n20951), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20950), .B2(n21168), .ZN(n20952) );
  AOI211_X1 U22862 ( .C1(n21147), .C2(n20953), .A(n20952), .B(n21161), .ZN(
        n20955) );
  NAND2_X1 U22863 ( .A1(n20955), .A2(n20954), .ZN(n20966) );
  NAND4_X1 U22864 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n20957), .A3(
        n20956), .A4(n20966), .ZN(n20961) );
  NAND3_X1 U22865 ( .A1(n21067), .A2(n20959), .A3(n20958), .ZN(n20960) );
  OAI211_X1 U22866 ( .C1(n20963), .C2(n20962), .A(n20961), .B(n20960), .ZN(
        n20968) );
  NAND2_X1 U22867 ( .A1(n21067), .A2(n20964), .ZN(n20965) );
  OAI211_X1 U22868 ( .C1(n21108), .C2(n21056), .A(n21151), .B(n20965), .ZN(
        n21139) );
  NOR2_X1 U22869 ( .A1(n20966), .A2(n21139), .ZN(n20967) );
  NOR2_X1 U22870 ( .A1(n21167), .A2(n20967), .ZN(n21138) );
  AOI22_X1 U22871 ( .A1(n21151), .A2(n20968), .B1(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n21138), .ZN(n20970) );
  OAI211_X1 U22872 ( .C1(n20971), .C2(n21144), .A(n20970), .B(n20969), .ZN(
        P3_U2847) );
  NOR2_X1 U22873 ( .A1(n20973), .A2(n20972), .ZN(n21082) );
  INV_X1 U22874 ( .A(n21147), .ZN(n21159) );
  OAI22_X1 U22875 ( .A1(n21115), .A2(n20983), .B1(n21171), .B2(n20974), .ZN(
        n20975) );
  OAI21_X1 U22876 ( .B1(n21159), .B2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n20975), .ZN(n20977) );
  OAI22_X1 U22877 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n21082), .B1(
        n20977), .B2(n20976), .ZN(n20981) );
  AOI22_X1 U22878 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n21062), .B1(
        n21166), .B2(n20978), .ZN(n20980) );
  NAND2_X1 U22879 ( .A1(n21137), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n20979) );
  OAI211_X1 U22880 ( .C1(n21080), .C2(n20981), .A(n20980), .B(n20979), .ZN(
        P3_U2840) );
  INV_X1 U22881 ( .A(n20999), .ZN(n20985) );
  NAND2_X1 U22882 ( .A1(n21029), .A2(n21026), .ZN(n20982) );
  NOR3_X1 U22883 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n20985), .A3(
        n20982), .ZN(n20989) );
  OAI21_X1 U22884 ( .B1(n21115), .B2(n20983), .A(n21170), .ZN(n21069) );
  NAND2_X1 U22885 ( .A1(n21073), .A2(n21069), .ZN(n20984) );
  OAI21_X1 U22886 ( .B1(n20985), .B2(n20984), .A(n21140), .ZN(n20996) );
  OAI22_X1 U22887 ( .A1(n21056), .A2(n20987), .B1(n20986), .B2(n20996), .ZN(
        n20988) );
  AOI211_X1 U22888 ( .C1(n20990), .C2(n21067), .A(n20989), .B(n20988), .ZN(
        n20994) );
  AOI22_X1 U22889 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n21062), .B1(
        n21166), .B2(n20991), .ZN(n20993) );
  NAND2_X1 U22890 ( .A1(n21137), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n20992) );
  OAI211_X1 U22891 ( .C1(n20994), .C2(n21080), .A(n20993), .B(n20992), .ZN(
        P3_U2837) );
  NAND2_X1 U22892 ( .A1(n21012), .A2(n21011), .ZN(n21003) );
  NAND2_X1 U22893 ( .A1(n21067), .A2(n21009), .ZN(n20995) );
  OAI211_X1 U22894 ( .C1(n21051), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n20996), .B(n20995), .ZN(n20997) );
  OAI21_X1 U22895 ( .B1(n20998), .B2(n20997), .A(n21151), .ZN(n21002) );
  NOR2_X1 U22896 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n21001) );
  AOI21_X1 U22897 ( .B1(n21075), .B2(n20999), .A(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n21000) );
  AOI211_X1 U22898 ( .C1(n21003), .C2(n21002), .A(n21001), .B(n21000), .ZN(
        n21004) );
  AOI211_X1 U22899 ( .C1(n21062), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n21005), .B(n21004), .ZN(n21006) );
  OAI21_X1 U22900 ( .B1(n21144), .B2(n21007), .A(n21006), .ZN(P3_U2836) );
  AOI211_X1 U22901 ( .C1(n21067), .C2(n21009), .A(n21015), .B(n21008), .ZN(
        n21010) );
  OAI211_X1 U22902 ( .C1(n21028), .C2(n21112), .A(n21010), .B(n21069), .ZN(
        n21013) );
  AOI22_X1 U22903 ( .A1(n21151), .A2(n21013), .B1(n21012), .B2(n21011), .ZN(
        n21016) );
  AOI222_X1 U22904 ( .A1(n21016), .A2(n21015), .B1(n21016), .B2(n21074), .C1(
        n21015), .C2(n21014), .ZN(n21017) );
  AOI21_X1 U22905 ( .B1(n21166), .B2(n21018), .A(n21017), .ZN(n21020) );
  NAND2_X1 U22906 ( .A1(n21020), .A2(n21019), .ZN(P3_U2835) );
  AOI21_X1 U22907 ( .B1(n21027), .B2(n21021), .A(n21175), .ZN(n21041) );
  AOI22_X1 U22908 ( .A1(n21183), .A2(n21023), .B1(n21067), .B2(n21022), .ZN(
        n21044) );
  NAND4_X1 U22909 ( .A1(n21029), .A2(n21028), .A3(n21027), .A4(n21026), .ZN(
        n21054) );
  NAND2_X1 U22910 ( .A1(n21183), .A2(n21030), .ZN(n21031) );
  OAI211_X1 U22911 ( .C1(n21032), .C2(n21110), .A(n21054), .B(n21031), .ZN(
        n21042) );
  NAND3_X1 U22912 ( .A1(n21151), .A2(n21033), .A3(n21042), .ZN(n21034) );
  OAI211_X1 U22913 ( .C1(n21036), .C2(n21144), .A(n21035), .B(n21034), .ZN(
        P3_U2833) );
  NOR2_X1 U22914 ( .A1(n21176), .A2(n21037), .ZN(n21046) );
  OAI211_X1 U22915 ( .C1(n21051), .C2(n21039), .A(n21038), .B(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21040) );
  NOR2_X1 U22916 ( .A1(n21041), .A2(n21040), .ZN(n21050) );
  AOI21_X1 U22917 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n21042), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21043) );
  AOI211_X1 U22918 ( .C1(n21044), .C2(n21050), .A(n21080), .B(n21043), .ZN(
        n21045) );
  AOI211_X1 U22919 ( .C1(n21166), .C2(n21047), .A(n21046), .B(n21045), .ZN(
        n21048) );
  OAI21_X1 U22920 ( .B1(n21074), .B2(n21049), .A(n21048), .ZN(P3_U2832) );
  NOR3_X1 U22921 ( .A1(n21051), .A2(n21050), .A3(n21052), .ZN(n21059) );
  NAND2_X1 U22922 ( .A1(n21053), .A2(n21052), .ZN(n21055) );
  OAI22_X1 U22923 ( .A1(n21057), .A2(n21056), .B1(n21055), .B2(n21054), .ZN(
        n21058) );
  AOI211_X1 U22924 ( .C1(n21067), .C2(n21060), .A(n21059), .B(n21058), .ZN(
        n21065) );
  AOI22_X1 U22925 ( .A1(n21062), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n21166), .B2(n21061), .ZN(n21064) );
  OAI211_X1 U22926 ( .C1(n21065), .C2(n21080), .A(n21064), .B(n21063), .ZN(
        P3_U2831) );
  NAND2_X1 U22927 ( .A1(n21137), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n21077) );
  AOI22_X1 U22928 ( .A1(n21183), .A2(n21068), .B1(n21067), .B2(n21066), .ZN(
        n21070) );
  NAND3_X1 U22929 ( .A1(n21070), .A2(n21074), .A3(n21069), .ZN(n21084) );
  NOR2_X1 U22930 ( .A1(n21071), .A2(n21084), .ZN(n21072) );
  AOI21_X1 U22931 ( .B1(n21073), .B2(n21072), .A(n21167), .ZN(n21083) );
  OAI221_X1 U22932 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n21075), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n21074), .A(n21083), .ZN(
        n21076) );
  OAI211_X1 U22933 ( .C1(n21078), .C2(n21144), .A(n21077), .B(n21076), .ZN(
        P3_U2839) );
  NOR3_X1 U22934 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n21080), .A3(
        n21079), .ZN(n21081) );
  AOI22_X1 U22935 ( .A1(n21167), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n21082), 
        .B2(n21081), .ZN(n21086) );
  OAI211_X1 U22936 ( .C1(n21140), .C2(n21084), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n21083), .ZN(n21085) );
  OAI211_X1 U22937 ( .C1(n21087), .C2(n21144), .A(n21086), .B(n21085), .ZN(
        P3_U2838) );
  AOI21_X1 U22938 ( .B1(n21183), .B2(n21089), .A(n21088), .ZN(n21090) );
  OAI211_X1 U22939 ( .C1(n21092), .C2(n21110), .A(n21091), .B(n21090), .ZN(
        n21093) );
  NAND2_X1 U22940 ( .A1(n21176), .A2(n21093), .ZN(n21099) );
  NAND2_X1 U22941 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21099), .ZN(
        n21101) );
  OAI21_X1 U22942 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n21104), .A(
        n21101), .ZN(n21095) );
  OAI211_X1 U22943 ( .C1(n21096), .C2(n21144), .A(n21095), .B(n21094), .ZN(
        P3_U2843) );
  AOI221_X1 U22944 ( .B1(n21100), .B2(n21099), .C1(n21098), .C2(n21099), .A(
        n21097), .ZN(n21102) );
  AOI22_X1 U22945 ( .A1(n21104), .A2(n21103), .B1(n21102), .B2(n21101), .ZN(
        n21106) );
  OAI211_X1 U22946 ( .C1(n21144), .C2(n21107), .A(n21106), .B(n21105), .ZN(
        P3_U2842) );
  OAI211_X1 U22947 ( .C1(n21111), .C2(n21110), .A(n21109), .B(n21108), .ZN(
        n21116) );
  NOR2_X1 U22948 ( .A1(n21122), .A2(n21135), .ZN(n21129) );
  AOI21_X1 U22949 ( .B1(n21113), .B2(n21129), .A(n21112), .ZN(n21114) );
  AOI211_X1 U22950 ( .C1(n21117), .C2(n21116), .A(n21115), .B(n21114), .ZN(
        n21118) );
  OAI211_X1 U22951 ( .C1(n21120), .C2(n21119), .A(n21151), .B(n21118), .ZN(
        n21131) );
  OAI221_X1 U22952 ( .B1(n21131), .B2(n21121), .C1(n21131), .C2(n21170), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n21127) );
  NOR2_X1 U22953 ( .A1(n21122), .A2(n21181), .ZN(n21136) );
  AOI22_X1 U22954 ( .A1(n21166), .A2(n21124), .B1(n21136), .B2(n21123), .ZN(
        n21125) );
  OAI221_X1 U22955 ( .B1(n21137), .B2(n21127), .C1(n21176), .C2(n21126), .A(
        n21125), .ZN(P3_U2844) );
  NOR2_X1 U22956 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n21181), .ZN(
        n21128) );
  AOI22_X1 U22957 ( .A1(n21166), .A2(n21130), .B1(n21129), .B2(n21128), .ZN(
        n21134) );
  NAND3_X1 U22958 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n21176), .A3(
        n21131), .ZN(n21132) );
  NAND3_X1 U22959 ( .A1(n21134), .A2(n21133), .A3(n21132), .ZN(P3_U2845) );
  AOI22_X1 U22960 ( .A1(n21137), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n21136), 
        .B2(n21135), .ZN(n21142) );
  OAI211_X1 U22961 ( .C1(n21140), .C2(n21139), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n21138), .ZN(n21141) );
  OAI211_X1 U22962 ( .C1(n21144), .C2(n21143), .A(n21142), .B(n21141), .ZN(
        P3_U2846) );
  AOI211_X1 U22963 ( .C1(n21148), .C2(n21147), .A(n21146), .B(n21145), .ZN(
        n21150) );
  AOI211_X1 U22964 ( .C1(n21151), .C2(n21150), .A(n21167), .B(n21149), .ZN(
        n21153) );
  AOI211_X1 U22965 ( .C1(n21166), .C2(n21154), .A(n21153), .B(n21152), .ZN(
        n21155) );
  OAI21_X1 U22966 ( .B1(n21181), .B2(n21156), .A(n21155), .ZN(P3_U2849) );
  AOI22_X1 U22967 ( .A1(n21167), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n21166), 
        .B2(n21157), .ZN(n21163) );
  OAI21_X1 U22968 ( .B1(n21159), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n21158), .ZN(n21160) );
  OAI211_X1 U22969 ( .C1(n21161), .C2(n21160), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n21176), .ZN(n21162) );
  OAI211_X1 U22970 ( .C1(n21164), .C2(n21181), .A(n21163), .B(n21162), .ZN(
        P3_U2852) );
  AOI22_X1 U22971 ( .A1(n21167), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n21166), 
        .B2(n21165), .ZN(n21180) );
  INV_X1 U22972 ( .A(n21168), .ZN(n21169) );
  OAI211_X1 U22973 ( .C1(n21172), .C2(n21171), .A(n21170), .B(n21169), .ZN(
        n21173) );
  OAI221_X1 U22974 ( .B1(n21175), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(
        n21175), .C2(n21174), .A(n21173), .ZN(n21177) );
  OAI211_X1 U22975 ( .C1(n21178), .C2(n21177), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n21176), .ZN(n21179) );
  OAI211_X1 U22976 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n21181), .A(
        n21180), .B(n21179), .ZN(P3_U2853) );
  NAND2_X1 U22977 ( .A1(n21619), .A2(n20098), .ZN(n21228) );
  INV_X1 U22978 ( .A(n21182), .ZN(n21227) );
  NOR2_X1 U22979 ( .A1(n21184), .A2(n21183), .ZN(n21186) );
  OAI222_X1 U22980 ( .A1(n21190), .A2(n21189), .B1(n21188), .B2(n21187), .C1(
        n21186), .C2(n21185), .ZN(n21246) );
  INV_X1 U22981 ( .A(n21191), .ZN(n21194) );
  NOR3_X1 U22982 ( .A1(n21194), .A2(n21193), .A3(n21192), .ZN(n21245) );
  OAI21_X1 U22983 ( .B1(P3_FLUSH_REG_SCAN_IN), .B2(P3_MORE_REG_SCAN_IN), .A(
        n21245), .ZN(n21195) );
  OAI211_X1 U22984 ( .C1(n21197), .C2(n21199), .A(n21196), .B(n21195), .ZN(
        n21219) );
  AOI22_X1 U22985 ( .A1(n21208), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n21198), .B2(n21199), .ZN(n21217) );
  MUX2_X1 U22986 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n21200), .S(
        n21199), .Z(n21212) );
  OR3_X1 U22987 ( .A1(n21205), .A2(n21204), .A3(n21201), .ZN(n21202) );
  AOI22_X1 U22988 ( .A1(n21205), .A2(n21204), .B1(n21203), .B2(n21202), .ZN(
        n21207) );
  OAI21_X1 U22989 ( .B1(n21208), .B2(n21207), .A(n21206), .ZN(n21211) );
  AND2_X1 U22990 ( .A1(n21212), .A2(n21211), .ZN(n21209) );
  OAI221_X1 U22991 ( .B1(n21212), .B2(n21211), .C1(n21210), .C2(n21209), .A(
        n21214), .ZN(n21216) );
  AOI21_X1 U22992 ( .B1(n21214), .B2(n21213), .A(n21212), .ZN(n21215) );
  AOI222_X1 U22993 ( .A1(n21217), .A2(n21216), .B1(n21217), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n21216), .C2(n21215), .ZN(
        n21218) );
  NOR4_X1 U22994 ( .A1(n21220), .A2(n21246), .A3(n21219), .A4(n21218), .ZN(
        n21243) );
  OAI211_X1 U22995 ( .C1(n21223), .C2(n21222), .A(n21221), .B(n21243), .ZN(
        n21231) );
  OAI21_X1 U22996 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n21659), .A(n21231), 
        .ZN(n21237) );
  OR3_X1 U22997 ( .A1(n21225), .A2(n21237), .A3(n21224), .ZN(n21226) );
  NAND4_X1 U22998 ( .A1(n21229), .A2(n21228), .A3(n21227), .A4(n21226), .ZN(
        P3_U2997) );
  OAI221_X1 U22999 ( .B1(n21232), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n21232), 
        .C2(n21231), .A(n21230), .ZN(P3_U3282) );
  AOI22_X1 U23000 ( .A1(n21235), .A2(n21234), .B1(n21619), .B2(n20098), .ZN(
        n21236) );
  INV_X1 U23001 ( .A(n21236), .ZN(n21240) );
  NOR2_X1 U23002 ( .A1(n21238), .A2(n21237), .ZN(n21239) );
  MUX2_X1 U23003 ( .A(n21240), .B(n21239), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n21242) );
  OAI211_X1 U23004 ( .C1(n21243), .C2(n21244), .A(n21242), .B(n21241), .ZN(
        P3_U2996) );
  NOR2_X1 U23005 ( .A1(n21245), .A2(n21244), .ZN(n21249) );
  MUX2_X1 U23006 ( .A(P3_MORE_REG_SCAN_IN), .B(n21246), .S(n21249), .Z(
        P3_U3295) );
  OAI21_X1 U23007 ( .B1(n21249), .B2(n21248), .A(n21247), .ZN(P3_U2637) );
  OAI211_X1 U23008 ( .C1(n21250), .C2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .B(n21622), .ZN(n21251) );
  OAI21_X1 U23009 ( .B1(n21252), .B2(n21251), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n21254) );
  NAND2_X1 U23010 ( .A1(n21254), .A2(n21253), .ZN(n21259) );
  AOI211_X1 U23011 ( .C1(n21257), .C2(n21622), .A(n21256), .B(n21255), .ZN(
        n21258) );
  MUX2_X1 U23012 ( .A(n21259), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n21258), 
        .Z(P1_U3485) );
  INV_X1 U23013 ( .A(n21402), .ZN(n21260) );
  OAI221_X1 U23014 ( .B1(n21271), .B2(n21260), .C1(n21271), .C2(n21331), .A(
        n21274), .ZN(n21270) );
  AOI22_X1 U23015 ( .A1(n21262), .A2(n21406), .B1(n21394), .B2(n21261), .ZN(
        n21269) );
  NAND2_X1 U23016 ( .A1(n21390), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n21268) );
  AOI21_X1 U23017 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n21331), .A(
        n21402), .ZN(n21263) );
  AOI211_X1 U23018 ( .C1(n21265), .C2(n21264), .A(n21263), .B(n21334), .ZN(
        n21266) );
  OAI21_X1 U23019 ( .B1(n21333), .B2(n21332), .A(n21266), .ZN(n21277) );
  NAND2_X1 U23020 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n21277), .ZN(
        n21267) );
  NAND4_X1 U23021 ( .A1(n21270), .A2(n21269), .A3(n21268), .A4(n21267), .ZN(
        P1_U3018) );
  AND2_X1 U23022 ( .A1(n21274), .A2(n21271), .ZN(n21278) );
  NAND2_X1 U23023 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n21303) );
  NOR2_X1 U23024 ( .A1(n21303), .A2(n21305), .ZN(n21325) );
  NAND4_X1 U23025 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(n21325), .A4(n21272), .ZN(
        n21273) );
  OAI22_X1 U23026 ( .A1(n21275), .A2(n21327), .B1(n21274), .B2(n21273), .ZN(
        n21276) );
  AOI221_X1 U23027 ( .B1(n21278), .B2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), 
        .C1(n21277), .C2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A(n21276), .ZN(
        n21280) );
  NAND2_X1 U23028 ( .A1(n21390), .A2(P1_REIP_REG_14__SCAN_IN), .ZN(n21279) );
  OAI211_X1 U23029 ( .C1(n21409), .C2(n21281), .A(n21280), .B(n21279), .ZN(
        P1_U3017) );
  AOI221_X1 U23030 ( .B1(n21284), .B2(n21337), .C1(n21283), .C2(n21337), .A(
        n21282), .ZN(n21302) );
  INV_X1 U23031 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21301) );
  NAND2_X1 U23032 ( .A1(n21301), .A2(n21285), .ZN(n21291) );
  OAI22_X1 U23033 ( .A1(n21287), .A2(n21327), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n21286), .ZN(n21288) );
  AOI211_X1 U23034 ( .C1(n21394), .C2(n21453), .A(n21289), .B(n21288), .ZN(
        n21290) );
  OAI221_X1 U23035 ( .B1(n21292), .B2(n21302), .C1(n21292), .C2(n21291), .A(
        n21290), .ZN(P1_U3025) );
  INV_X1 U23036 ( .A(n21293), .ZN(n21297) );
  NAND2_X1 U23037 ( .A1(n21294), .A2(n21301), .ZN(n21296) );
  OAI22_X1 U23038 ( .A1(n21297), .A2(n21327), .B1(n21296), .B2(n21295), .ZN(
        n21298) );
  AOI211_X1 U23039 ( .C1(n21394), .C2(n21438), .A(n21299), .B(n21298), .ZN(
        n21300) );
  OAI21_X1 U23040 ( .B1(n21302), .B2(n21301), .A(n21300), .ZN(P1_U3026) );
  OAI21_X1 U23041 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n21303), .ZN(n21304) );
  OAI22_X1 U23042 ( .A1(n21327), .A2(n21306), .B1(n21305), .B2(n21304), .ZN(
        n21307) );
  AOI21_X1 U23043 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n21308), .A(
        n21307), .ZN(n21310) );
  NAND2_X1 U23044 ( .A1(n21390), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n21309) );
  OAI211_X1 U23045 ( .C1(n21409), .C2(n21499), .A(n21310), .B(n21309), .ZN(
        P1_U3021) );
  NOR2_X1 U23046 ( .A1(n21324), .A2(n21311), .ZN(n21317) );
  OAI21_X1 U23047 ( .B1(n21347), .B2(n21317), .A(n21312), .ZN(n21323) );
  OAI22_X1 U23048 ( .A1(n21378), .A2(n21313), .B1(n21409), .B2(n21522), .ZN(
        n21314) );
  AOI21_X1 U23049 ( .B1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n21323), .A(
        n21314), .ZN(n21319) );
  NAND3_X1 U23050 ( .A1(n21317), .A2(n21316), .A3(n21315), .ZN(n21318) );
  OAI211_X1 U23051 ( .C1(n21320), .C2(n21327), .A(n21319), .B(n21318), .ZN(
        P1_U3019) );
  OAI21_X1 U23052 ( .B1(n21409), .B2(n21512), .A(n21321), .ZN(n21322) );
  AOI221_X1 U23053 ( .B1(n21325), .B2(n21324), .C1(n21323), .C2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n21322), .ZN(n21326) );
  OAI21_X1 U23054 ( .B1(n21328), .B2(n21327), .A(n21326), .ZN(P1_U3020) );
  AOI22_X1 U23055 ( .A1(n21394), .A2(n21330), .B1(n21406), .B2(n21329), .ZN(
        n21341) );
  NAND3_X1 U23056 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(n21331), .ZN(n21336) );
  AOI21_X1 U23057 ( .B1(n21344), .B2(n21333), .A(n21332), .ZN(n21335) );
  AOI211_X1 U23058 ( .C1(n21337), .C2(n21336), .A(n21335), .B(n21334), .ZN(
        n21346) );
  INV_X1 U23059 ( .A(n21346), .ZN(n21365) );
  NAND2_X1 U23060 ( .A1(n21344), .A2(n21342), .ZN(n21360) );
  NOR2_X1 U23061 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n21360), .ZN(
        n21366) );
  NOR2_X1 U23062 ( .A1(n21378), .A2(n21338), .ZN(n21339) );
  AOI211_X1 U23063 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n21365), .A(
        n21366), .B(n21339), .ZN(n21340) );
  NAND2_X1 U23064 ( .A1(n21341), .A2(n21340), .ZN(P1_U3016) );
  AND4_X1 U23065 ( .A1(n21348), .A2(n21344), .A3(n21343), .A4(n21342), .ZN(
        n21345) );
  AOI21_X1 U23066 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n21390), .A(n21345), 
        .ZN(n21351) );
  OAI21_X1 U23067 ( .B1(n21348), .B2(n21347), .A(n21346), .ZN(n21355) );
  AOI22_X1 U23068 ( .A1(n21349), .A2(n21406), .B1(
        P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n21355), .ZN(n21350) );
  OAI211_X1 U23069 ( .C1(n21409), .C2(n21563), .A(n21351), .B(n21350), .ZN(
        P1_U3013) );
  OAI21_X1 U23070 ( .B1(n21353), .B2(n21360), .A(n21352), .ZN(n21354) );
  AOI22_X1 U23071 ( .A1(n21406), .A2(n21356), .B1(n21355), .B2(n21354), .ZN(
        n21358) );
  NAND2_X1 U23072 ( .A1(n21390), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n21357) );
  OAI211_X1 U23073 ( .C1(n21409), .C2(n21557), .A(n21358), .B(n21357), .ZN(
        P1_U3014) );
  NOR2_X1 U23074 ( .A1(n21378), .A2(n21359), .ZN(n21363) );
  NOR3_X1 U23075 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n21361), .A3(
        n21360), .ZN(n21362) );
  AOI211_X1 U23076 ( .C1(n21406), .C2(n21364), .A(n21363), .B(n21362), .ZN(
        n21368) );
  OAI21_X1 U23077 ( .B1(n21366), .B2(n21365), .A(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n21367) );
  OAI211_X1 U23078 ( .C1(n21409), .C2(n21544), .A(n21368), .B(n21367), .ZN(
        P1_U3015) );
  INV_X1 U23079 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n21379) );
  INV_X1 U23080 ( .A(n21369), .ZN(n21372) );
  INV_X1 U23081 ( .A(n21370), .ZN(n21371) );
  AOI22_X1 U23082 ( .A1(n21372), .A2(n21406), .B1(n21394), .B2(n21371), .ZN(
        n21377) );
  INV_X1 U23083 ( .A(n21399), .ZN(n21374) );
  AOI22_X1 U23084 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n21375), .B1(
        n21374), .B2(n21373), .ZN(n21376) );
  OAI211_X1 U23085 ( .C1(n21379), .C2(n21378), .A(n21377), .B(n21376), .ZN(
        P1_U3012) );
  INV_X1 U23086 ( .A(n21380), .ZN(n21384) );
  NOR3_X1 U23087 ( .A1(n21399), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n21381), .ZN(n21382) );
  AOI211_X1 U23088 ( .C1(n21384), .C2(n21406), .A(n21383), .B(n21382), .ZN(
        n21388) );
  OAI21_X1 U23089 ( .B1(n21386), .B2(n21385), .A(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n21387) );
  OAI211_X1 U23090 ( .C1(n21409), .C2(n21389), .A(n21388), .B(n21387), .ZN(
        P1_U3009) );
  AOI22_X1 U23091 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n21391), .B1(
        n21390), .B2(P1_REIP_REG_23__SCAN_IN), .ZN(n21397) );
  INV_X1 U23092 ( .A(n21392), .ZN(n21395) );
  AOI22_X1 U23093 ( .A1(n21395), .A2(n21406), .B1(n21394), .B2(n21393), .ZN(
        n21396) );
  OAI211_X1 U23094 ( .C1(n21399), .C2(n21398), .A(n21397), .B(n21396), .ZN(
        P1_U3008) );
  AOI21_X1 U23095 ( .B1(n21402), .B2(n21401), .A(n21400), .ZN(n21404) );
  AOI211_X1 U23096 ( .C1(n21406), .C2(n21405), .A(n21404), .B(n21403), .ZN(
        n21408) );
  OAI211_X1 U23097 ( .C1(n21410), .C2(n21409), .A(n21408), .B(n21407), .ZN(
        P1_U3031) );
  INV_X1 U23098 ( .A(n21411), .ZN(n21458) );
  NOR2_X1 U23099 ( .A1(n21559), .A2(n21412), .ZN(n21414) );
  AOI211_X1 U23100 ( .C1(n21415), .C2(n21469), .A(n21414), .B(n21413), .ZN(
        n21417) );
  NAND2_X1 U23101 ( .A1(n21938), .A2(n21423), .ZN(n21416) );
  OAI211_X1 U23102 ( .C1(n21458), .C2(n21418), .A(n21417), .B(n21416), .ZN(
        n21421) );
  NOR2_X1 U23103 ( .A1(n21448), .A2(n21419), .ZN(n21420) );
  AOI211_X1 U23104 ( .C1(n21536), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n21421), .B(n21420), .ZN(n21422) );
  OAI21_X1 U23105 ( .B1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n21565), .A(
        n21422), .ZN(P1_U2839) );
  INV_X1 U23106 ( .A(n21448), .ZN(n21431) );
  AOI21_X1 U23107 ( .B1(n21424), .B2(n21423), .A(n21532), .ZN(n21426) );
  NAND2_X1 U23108 ( .A1(n21533), .A2(P1_EBX_REG_4__SCAN_IN), .ZN(n21425) );
  OAI211_X1 U23109 ( .C1(n21427), .C2(n21562), .A(n21426), .B(n21425), .ZN(
        n21430) );
  NOR2_X1 U23110 ( .A1(n21566), .A2(n21428), .ZN(n21429) );
  AOI211_X1 U23111 ( .C1(n21432), .C2(n21431), .A(n21430), .B(n21429), .ZN(
        n21436) );
  NOR3_X1 U23112 ( .A1(n21433), .A2(n14961), .A3(n21459), .ZN(n21434) );
  NAND2_X1 U23113 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n21434), .ZN(n21442) );
  OAI211_X1 U23114 ( .C1(P1_REIP_REG_4__SCAN_IN), .C2(n21434), .A(n21442), .B(
        n21552), .ZN(n21435) );
  OAI211_X1 U23115 ( .C1(n21565), .C2(n21437), .A(n21436), .B(n21435), .ZN(
        P1_U2836) );
  AOI22_X1 U23116 ( .A1(n21438), .A2(n21469), .B1(n21533), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n21439) );
  OAI211_X1 U23117 ( .C1(n21566), .C2(n21440), .A(n21439), .B(n21560), .ZN(
        n21441) );
  INV_X1 U23118 ( .A(n21441), .ZN(n21447) );
  OAI21_X1 U23119 ( .B1(n21495), .B2(n21443), .A(n21442), .ZN(n21445) );
  NOR2_X1 U23120 ( .A1(n21443), .A2(n21442), .ZN(n21460) );
  INV_X1 U23121 ( .A(n21460), .ZN(n21444) );
  NAND2_X1 U23122 ( .A1(n21445), .A2(n21444), .ZN(n21446) );
  OAI211_X1 U23123 ( .C1(n21449), .C2(n21448), .A(n21447), .B(n21446), .ZN(
        n21450) );
  INV_X1 U23124 ( .A(n21450), .ZN(n21451) );
  OAI21_X1 U23125 ( .B1(n21452), .B2(n21565), .A(n21451), .ZN(P1_U2835) );
  AOI22_X1 U23126 ( .A1(n21453), .A2(n21469), .B1(n21533), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n21454) );
  OAI211_X1 U23127 ( .C1(n21566), .C2(n21455), .A(n21454), .B(n21560), .ZN(
        n21456) );
  AOI21_X1 U23128 ( .B1(n21457), .B2(n21541), .A(n21456), .ZN(n21462) );
  OAI21_X1 U23129 ( .B1(n21465), .B2(n21459), .A(n21458), .ZN(n21474) );
  OAI21_X1 U23130 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(n21460), .A(n21474), .ZN(
        n21461) );
  OAI211_X1 U23131 ( .C1(n21565), .C2(n21463), .A(n21462), .B(n21461), .ZN(
        P1_U2834) );
  INV_X1 U23132 ( .A(n21464), .ZN(n21470) );
  NAND2_X1 U23133 ( .A1(n21465), .A2(n21483), .ZN(n21466) );
  OAI22_X1 U23134 ( .A1(n21559), .A2(n21467), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n21466), .ZN(n21468) );
  AOI21_X1 U23135 ( .B1(n21470), .B2(n21469), .A(n21468), .ZN(n21471) );
  OAI211_X1 U23136 ( .C1(n21566), .C2(n21472), .A(n21471), .B(n21560), .ZN(
        n21473) );
  INV_X1 U23137 ( .A(n21473), .ZN(n21477) );
  AOI22_X1 U23138 ( .A1(n21475), .A2(n21541), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n21474), .ZN(n21476) );
  OAI211_X1 U23139 ( .C1(n21478), .C2(n21565), .A(n21477), .B(n21476), .ZN(
        P1_U2833) );
  OAI22_X1 U23140 ( .A1(n21565), .A2(n21480), .B1(n21479), .B2(n21559), .ZN(
        n21481) );
  INV_X1 U23141 ( .A(n21481), .ZN(n21492) );
  NAND2_X1 U23142 ( .A1(n21483), .A2(n21482), .ZN(n21484) );
  OAI21_X1 U23143 ( .B1(n21485), .B2(n21484), .A(n21560), .ZN(n21490) );
  OAI22_X1 U23144 ( .A1(n21488), .A2(n21571), .B1(n21487), .B2(n21486), .ZN(
        n21489) );
  AOI211_X1 U23145 ( .C1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n21536), .A(
        n21490), .B(n21489), .ZN(n21491) );
  OAI211_X1 U23146 ( .C1(n21562), .C2(n21493), .A(n21492), .B(n21491), .ZN(
        P1_U2832) );
  OAI21_X1 U23147 ( .B1(n21496), .B2(n21495), .A(n21494), .ZN(n21497) );
  INV_X1 U23148 ( .A(n21497), .ZN(n21508) );
  OAI22_X1 U23149 ( .A1(n21499), .A2(n21562), .B1(n21559), .B2(n21498), .ZN(
        n21500) );
  INV_X1 U23150 ( .A(n21500), .ZN(n21501) );
  OAI211_X1 U23151 ( .C1(n21566), .C2(n21502), .A(n21501), .B(n21560), .ZN(
        n21503) );
  INV_X1 U23152 ( .A(n21503), .ZN(n21507) );
  AOI22_X1 U23153 ( .A1(n21505), .A2(n21541), .B1(n21535), .B2(n21504), .ZN(
        n21506) );
  OAI211_X1 U23154 ( .C1(n21510), .C2(n21508), .A(n21507), .B(n21506), .ZN(
        P1_U2830) );
  INV_X1 U23155 ( .A(n21509), .ZN(n21520) );
  AOI21_X1 U23156 ( .B1(P1_REIP_REG_11__SCAN_IN), .B2(n21552), .A(n21510), 
        .ZN(n21519) );
  INV_X1 U23157 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n21511) );
  OAI22_X1 U23158 ( .A1(n21512), .A2(n21562), .B1(n21511), .B2(n21559), .ZN(
        n21513) );
  AOI211_X1 U23159 ( .C1(n21536), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n21532), .B(n21513), .ZN(n21518) );
  OAI22_X1 U23160 ( .A1(n21515), .A2(n21565), .B1(n21571), .B2(n21514), .ZN(
        n21516) );
  INV_X1 U23161 ( .A(n21516), .ZN(n21517) );
  OAI211_X1 U23162 ( .C1(n21520), .C2(n21519), .A(n21518), .B(n21517), .ZN(
        P1_U2829) );
  AOI21_X1 U23163 ( .B1(P1_REIP_REG_12__SCAN_IN), .B2(n21552), .A(n21520), 
        .ZN(n21528) );
  OAI22_X1 U23164 ( .A1(n21522), .A2(n21562), .B1(n21521), .B2(n21559), .ZN(
        n21523) );
  AOI211_X1 U23165 ( .C1(n21536), .C2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n21532), .B(n21523), .ZN(n21527) );
  AOI22_X1 U23166 ( .A1(n21525), .A2(n21535), .B1(n21541), .B2(n21524), .ZN(
        n21526) );
  OAI211_X1 U23167 ( .C1(n21529), .C2(n21528), .A(n21527), .B(n21526), .ZN(
        P1_U2828) );
  INV_X1 U23168 ( .A(n21530), .ZN(n21531) );
  AOI21_X1 U23169 ( .B1(n21552), .B2(P1_REIP_REG_16__SCAN_IN), .A(n21531), 
        .ZN(n21539) );
  AOI21_X1 U23170 ( .B1(n21533), .B2(P1_EBX_REG_16__SCAN_IN), .A(n21532), .ZN(
        n21538) );
  AOI22_X1 U23171 ( .A1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n21536), .B1(
        n21535), .B2(n21534), .ZN(n21537) );
  OAI211_X1 U23172 ( .C1(n21539), .C2(n21554), .A(n21538), .B(n21537), .ZN(
        n21540) );
  AOI21_X1 U23173 ( .B1(n21542), .B2(n21541), .A(n21540), .ZN(n21543) );
  OAI21_X1 U23174 ( .B1(n21562), .B2(n21544), .A(n21543), .ZN(P1_U2824) );
  OAI22_X1 U23175 ( .A1(n21546), .A2(n21565), .B1(n21566), .B2(n21545), .ZN(
        n21548) );
  OAI21_X1 U23176 ( .B1(n21559), .B2(n15825), .A(n21560), .ZN(n21547) );
  NOR2_X1 U23177 ( .A1(n21548), .A2(n21547), .ZN(n21549) );
  OAI21_X1 U23178 ( .B1(n21550), .B2(n21571), .A(n21549), .ZN(n21551) );
  INV_X1 U23179 ( .A(n21551), .ZN(n21556) );
  NAND2_X1 U23180 ( .A1(n21552), .A2(n21577), .ZN(n21575) );
  INV_X1 U23181 ( .A(n21575), .ZN(n21553) );
  OAI21_X1 U23182 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(n21554), .A(n21553), 
        .ZN(n21555) );
  OAI211_X1 U23183 ( .C1(n21557), .C2(n21562), .A(n21556), .B(n21555), .ZN(
        P1_U2823) );
  OR2_X1 U23184 ( .A1(n21559), .A2(n21558), .ZN(n21561) );
  OAI211_X1 U23185 ( .C1(n21563), .C2(n21562), .A(n21561), .B(n21560), .ZN(
        n21569) );
  INV_X1 U23186 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n21567) );
  OAI22_X1 U23187 ( .A1(n21567), .A2(n21566), .B1(n21565), .B2(n21564), .ZN(
        n21568) );
  NOR2_X1 U23188 ( .A1(n21569), .A2(n21568), .ZN(n21570) );
  OAI21_X1 U23189 ( .B1(n21572), .B2(n21571), .A(n21570), .ZN(n21573) );
  INV_X1 U23190 ( .A(n21573), .ZN(n21574) );
  OAI221_X1 U23191 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n21577), .C1(n21576), 
        .C2(n21575), .A(n21574), .ZN(P1_U2822) );
  OAI21_X1 U23192 ( .B1(n21579), .B2(n14903), .A(n21578), .ZN(P1_U2806) );
  AOI22_X1 U23193 ( .A1(n21581), .A2(n21580), .B1(n21850), .B2(n21925), .ZN(
        n21586) );
  INV_X1 U23194 ( .A(n21582), .ZN(n21584) );
  NOR2_X1 U23195 ( .A1(n21584), .A2(n21583), .ZN(n21600) );
  NOR2_X1 U23196 ( .A1(n21587), .A2(n21600), .ZN(n21585) );
  AOI22_X1 U23197 ( .A1(n21915), .A2(n21587), .B1(n21586), .B2(n21585), .ZN(
        P1_U3478) );
  AOI21_X1 U23198 ( .B1(n21588), .B2(n21622), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n21590) );
  OAI21_X1 U23199 ( .B1(n21592), .B2(n21590), .A(n21589), .ZN(P1_U3163) );
  INV_X1 U23200 ( .A(n21591), .ZN(n21595) );
  AOI211_X1 U23201 ( .C1(P1_STATE2_REG_3__SCAN_IN), .C2(n21595), .A(n21593), 
        .B(n21592), .ZN(n21594) );
  INV_X1 U23202 ( .A(n21594), .ZN(P1_U3466) );
  AOI21_X1 U23203 ( .B1(n21597), .B2(n21596), .A(n21595), .ZN(n21598) );
  OAI22_X1 U23204 ( .A1(n21600), .A2(n21599), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n21598), .ZN(n21601) );
  OAI21_X1 U23205 ( .B1(n21602), .B2(n22310), .A(n21601), .ZN(P1_U3161) );
  OAI21_X1 U23206 ( .B1(n21605), .B2(n21936), .A(n21603), .ZN(P1_U2805) );
  INV_X1 U23207 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n21604) );
  OAI21_X1 U23208 ( .B1(n21605), .B2(n21604), .A(n21603), .ZN(P1_U3465) );
  INV_X1 U23209 ( .A(n21606), .ZN(n21608) );
  OAI21_X1 U23210 ( .B1(n21610), .B2(n21607), .A(n21608), .ZN(P2_U2818) );
  OAI21_X1 U23211 ( .B1(n21610), .B2(n21609), .A(n21608), .ZN(P2_U3592) );
  INV_X1 U23212 ( .A(n21611), .ZN(n21613) );
  OAI21_X1 U23213 ( .B1(n21615), .B2(n21612), .A(n21613), .ZN(P3_U2636) );
  OAI21_X1 U23214 ( .B1(n21615), .B2(n21614), .A(n21613), .ZN(P3_U3281) );
  INV_X1 U23215 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21616) );
  AOI21_X1 U23216 ( .B1(HOLD), .B2(n21617), .A(n21616), .ZN(n21620) );
  AOI21_X1 U23217 ( .B1(n21619), .B2(P3_STATE_REG_1__SCAN_IN), .A(n21618), 
        .ZN(n21672) );
  AOI21_X1 U23218 ( .B1(n21658), .B2(NA), .A(n21666), .ZN(n21670) );
  OAI22_X1 U23219 ( .A1(n21621), .A2(n21620), .B1(n21672), .B2(n21670), .ZN(
        P3_U3029) );
  INV_X1 U23220 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21630) );
  OAI21_X1 U23221 ( .B1(NA), .B2(n21622), .A(n21631), .ZN(n21623) );
  OAI211_X1 U23222 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n21630), .A(
        P1_STATE_REG_0__SCAN_IN), .B(n21623), .ZN(n21629) );
  NAND2_X1 U23223 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n21624), .ZN(n21632) );
  INV_X1 U23224 ( .A(n21632), .ZN(n21635) );
  AOI221_X1 U23225 ( .B1(n21630), .B2(P1_STATE_REG_0__SCAN_IN), .C1(n21632), 
        .C2(P1_STATE_REG_0__SCAN_IN), .A(n21625), .ZN(n21626) );
  AOI22_X1 U23226 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n21635), .B1(n21626), 
        .B2(n21667), .ZN(n21628) );
  OAI211_X1 U23227 ( .C1(n21629), .C2(n21665), .A(n21628), .B(n21627), .ZN(
        P1_U3196) );
  AOI21_X1 U23228 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(HOLD), .A(n21630), .ZN(
        n21638) );
  AOI22_X1 U23229 ( .A1(n21631), .A2(HOLD), .B1(P1_STATE_REG_0__SCAN_IN), .B2(
        n21638), .ZN(n21634) );
  NAND3_X1 U23230 ( .A1(n21634), .A2(n21633), .A3(n21632), .ZN(P1_U3195) );
  AOI22_X1 U23231 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(NA), .B2(
        n13632), .ZN(n21637) );
  OAI21_X1 U23232 ( .B1(n21635), .B2(n13632), .A(n12613), .ZN(n21636) );
  OAI221_X1 U23233 ( .B1(n22307), .B2(n21638), .C1(n22307), .C2(n21637), .A(
        n21636), .ZN(P1_U3194) );
  OAI21_X1 U23234 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(P2_STATE_REG_1__SCAN_IN), 
        .A(HOLD), .ZN(n21643) );
  NAND2_X1 U23235 ( .A1(n21639), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n21649) );
  NAND2_X1 U23236 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n21649), .ZN(n21653) );
  INV_X1 U23237 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21644) );
  AOI22_X1 U23238 ( .A1(n21640), .A2(n21653), .B1(n21644), .B2(n17337), .ZN(
        n21642) );
  NAND2_X1 U23239 ( .A1(n21641), .A2(NA), .ZN(n21652) );
  OAI211_X1 U23240 ( .C1(n17340), .C2(n21643), .A(n21642), .B(n21652), .ZN(
        P2_U3209) );
  NAND2_X1 U23241 ( .A1(n21665), .A2(n21644), .ZN(n21651) );
  AOI211_X1 U23242 ( .C1(P2_STATE_REG_2__SCAN_IN), .C2(HOLD), .A(n21655), .B(
        n21644), .ZN(n21646) );
  AOI211_X1 U23243 ( .C1(n21647), .C2(n21651), .A(n21646), .B(n21645), .ZN(
        n21648) );
  NAND2_X1 U23244 ( .A1(n21648), .A2(n21649), .ZN(P2_U3210) );
  OAI22_X1 U23245 ( .A1(NA), .A2(n21649), .B1(P2_STATE_REG_1__SCAN_IN), .B2(
        P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n21650) );
  AOI22_X1 U23246 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(HOLD), .B1(n21651), .B2(
        n21650), .ZN(n21656) );
  NAND3_X1 U23247 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n21653), .A3(n21652), 
        .ZN(n21654) );
  OAI21_X1 U23248 ( .B1(n21656), .B2(n21655), .A(n21654), .ZN(P2_U3211) );
  OAI211_X1 U23249 ( .C1(n21666), .C2(n21665), .A(P3_STATE_REG_0__SCAN_IN), 
        .B(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21663) );
  NOR2_X1 U23250 ( .A1(HOLD), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n21674)
         );
  NAND2_X1 U23251 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n21666), .ZN(n21657) );
  NOR2_X1 U23252 ( .A1(n21674), .A2(n21657), .ZN(n21661) );
  NOR2_X1 U23253 ( .A1(n21659), .A2(n21658), .ZN(n21668) );
  AOI211_X1 U23254 ( .C1(n21661), .C2(n21664), .A(n21660), .B(n21668), .ZN(
        n21662) );
  OAI211_X1 U23255 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(n21664), .A(n21663), 
        .B(n21662), .ZN(P3_U3030) );
  OAI22_X1 U23256 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(n21666), .B2(n21665), .ZN(n21669)
         );
  OAI221_X1 U23257 ( .B1(n21669), .B2(n21668), .C1(n21669), .C2(n21667), .A(
        P3_STATE_REG_0__SCAN_IN), .ZN(n21673) );
  INV_X1 U23258 ( .A(n21670), .ZN(n21671) );
  OAI22_X1 U23259 ( .A1(n21674), .A2(n21673), .B1(n21672), .B2(n21671), .ZN(
        P3_U3031) );
  NOR2_X1 U23260 ( .A1(n21761), .A2(n21675), .ZN(n21678) );
  AOI21_X1 U23261 ( .B1(P1_UWORD_REG_0__SCAN_IN), .B2(n21729), .A(n21678), 
        .ZN(n21676) );
  OAI21_X1 U23262 ( .B1(n21677), .B2(n21766), .A(n21676), .ZN(P1_U2937) );
  AOI21_X1 U23263 ( .B1(P1_LWORD_REG_0__SCAN_IN), .B2(n21729), .A(n21678), 
        .ZN(n21679) );
  OAI21_X1 U23264 ( .B1(n21680), .B2(n21766), .A(n21679), .ZN(P1_U2952) );
  NOR2_X1 U23265 ( .A1(n21761), .A2(n21681), .ZN(n21683) );
  AOI21_X1 U23266 ( .B1(P1_UWORD_REG_1__SCAN_IN), .B2(n21729), .A(n21683), 
        .ZN(n21682) );
  OAI21_X1 U23267 ( .B1(n13042), .B2(n21766), .A(n21682), .ZN(P1_U2938) );
  AOI21_X1 U23268 ( .B1(P1_LWORD_REG_1__SCAN_IN), .B2(n21729), .A(n21683), 
        .ZN(n21684) );
  OAI21_X1 U23269 ( .B1(n21685), .B2(n21766), .A(n21684), .ZN(P1_U2953) );
  NOR2_X1 U23270 ( .A1(n21761), .A2(n21686), .ZN(n21689) );
  AOI21_X1 U23271 ( .B1(P1_UWORD_REG_2__SCAN_IN), .B2(n21729), .A(n21689), 
        .ZN(n21687) );
  OAI21_X1 U23272 ( .B1(n21688), .B2(n21766), .A(n21687), .ZN(P1_U2939) );
  AOI21_X1 U23273 ( .B1(P1_LWORD_REG_2__SCAN_IN), .B2(n21729), .A(n21689), 
        .ZN(n21690) );
  OAI21_X1 U23274 ( .B1(n21691), .B2(n21766), .A(n21690), .ZN(P1_U2954) );
  AOI22_X1 U23275 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n21729), .B1(n21692), 
        .B2(P1_EAX_REG_3__SCAN_IN), .ZN(n21694) );
  NAND2_X1 U23276 ( .A1(n21694), .A2(n21693), .ZN(P1_U2955) );
  NOR2_X1 U23277 ( .A1(n21761), .A2(n21695), .ZN(n21698) );
  AOI21_X1 U23278 ( .B1(P1_UWORD_REG_4__SCAN_IN), .B2(n21729), .A(n21698), 
        .ZN(n21696) );
  OAI21_X1 U23279 ( .B1(n21697), .B2(n21766), .A(n21696), .ZN(P1_U2941) );
  AOI21_X1 U23280 ( .B1(P1_LWORD_REG_4__SCAN_IN), .B2(n21729), .A(n21698), 
        .ZN(n21699) );
  OAI21_X1 U23281 ( .B1(n21700), .B2(n21766), .A(n21699), .ZN(P1_U2956) );
  NOR2_X1 U23282 ( .A1(n21761), .A2(n21701), .ZN(n21704) );
  AOI21_X1 U23283 ( .B1(P1_UWORD_REG_5__SCAN_IN), .B2(n21729), .A(n21704), 
        .ZN(n21702) );
  OAI21_X1 U23284 ( .B1(n21703), .B2(n21766), .A(n21702), .ZN(P1_U2942) );
  AOI21_X1 U23285 ( .B1(P1_LWORD_REG_5__SCAN_IN), .B2(n21729), .A(n21704), 
        .ZN(n21705) );
  OAI21_X1 U23286 ( .B1(n12875), .B2(n21766), .A(n21705), .ZN(P1_U2957) );
  NOR2_X1 U23287 ( .A1(n21761), .A2(n21706), .ZN(n21709) );
  AOI21_X1 U23288 ( .B1(P1_UWORD_REG_6__SCAN_IN), .B2(n21729), .A(n21709), 
        .ZN(n21707) );
  OAI21_X1 U23289 ( .B1(n21708), .B2(n21766), .A(n21707), .ZN(P1_U2943) );
  AOI21_X1 U23290 ( .B1(P1_LWORD_REG_6__SCAN_IN), .B2(n21729), .A(n21709), 
        .ZN(n21710) );
  OAI21_X1 U23291 ( .B1(n21711), .B2(n21766), .A(n21710), .ZN(P1_U2958) );
  NOR2_X1 U23292 ( .A1(n21761), .A2(n21712), .ZN(n21715) );
  AOI21_X1 U23293 ( .B1(P1_UWORD_REG_7__SCAN_IN), .B2(n21729), .A(n21715), 
        .ZN(n21713) );
  OAI21_X1 U23294 ( .B1(n21714), .B2(n21766), .A(n21713), .ZN(P1_U2944) );
  AOI21_X1 U23295 ( .B1(P1_LWORD_REG_7__SCAN_IN), .B2(n21729), .A(n21715), 
        .ZN(n21716) );
  OAI21_X1 U23296 ( .B1(n15264), .B2(n21766), .A(n21716), .ZN(P1_U2959) );
  INV_X1 U23297 ( .A(n21717), .ZN(n21718) );
  NOR2_X1 U23298 ( .A1(n21761), .A2(n21718), .ZN(n21721) );
  AOI21_X1 U23299 ( .B1(P1_UWORD_REG_8__SCAN_IN), .B2(n21729), .A(n21721), 
        .ZN(n21719) );
  OAI21_X1 U23300 ( .B1(n21720), .B2(n21766), .A(n21719), .ZN(P1_U2945) );
  AOI21_X1 U23301 ( .B1(P1_LWORD_REG_8__SCAN_IN), .B2(n21729), .A(n21721), 
        .ZN(n21722) );
  OAI21_X1 U23302 ( .B1(n21723), .B2(n21766), .A(n21722), .ZN(P1_U2960) );
  INV_X1 U23303 ( .A(n21724), .ZN(n21725) );
  NOR2_X1 U23304 ( .A1(n21761), .A2(n21725), .ZN(n21728) );
  AOI21_X1 U23305 ( .B1(P1_UWORD_REG_9__SCAN_IN), .B2(n21729), .A(n21728), 
        .ZN(n21726) );
  OAI21_X1 U23306 ( .B1(n21727), .B2(n21766), .A(n21726), .ZN(P1_U2946) );
  AOI21_X1 U23307 ( .B1(P1_LWORD_REG_9__SCAN_IN), .B2(n21729), .A(n21728), 
        .ZN(n21730) );
  OAI21_X1 U23308 ( .B1(n21731), .B2(n21766), .A(n21730), .ZN(P1_U2961) );
  INV_X1 U23309 ( .A(n21732), .ZN(n21733) );
  NOR2_X1 U23310 ( .A1(n21761), .A2(n21733), .ZN(n21736) );
  AOI21_X1 U23311 ( .B1(P1_UWORD_REG_10__SCAN_IN), .B2(n21729), .A(n21736), 
        .ZN(n21734) );
  OAI21_X1 U23312 ( .B1(n21735), .B2(n21766), .A(n21734), .ZN(P1_U2947) );
  AOI21_X1 U23313 ( .B1(P1_LWORD_REG_10__SCAN_IN), .B2(n21729), .A(n21736), 
        .ZN(n21737) );
  OAI21_X1 U23314 ( .B1(n21738), .B2(n21766), .A(n21737), .ZN(P1_U2962) );
  INV_X1 U23315 ( .A(n21739), .ZN(n21740) );
  NOR2_X1 U23316 ( .A1(n21761), .A2(n21740), .ZN(n21742) );
  AOI21_X1 U23317 ( .B1(P1_UWORD_REG_11__SCAN_IN), .B2(n21729), .A(n21742), 
        .ZN(n21741) );
  OAI21_X1 U23318 ( .B1(n13231), .B2(n21766), .A(n21741), .ZN(P1_U2948) );
  AOI21_X1 U23319 ( .B1(P1_LWORD_REG_11__SCAN_IN), .B2(n21729), .A(n21742), 
        .ZN(n21743) );
  OAI21_X1 U23320 ( .B1(n21744), .B2(n21766), .A(n21743), .ZN(P1_U2963) );
  INV_X1 U23321 ( .A(n21745), .ZN(n21746) );
  NOR2_X1 U23322 ( .A1(n21761), .A2(n21746), .ZN(n21749) );
  AOI21_X1 U23323 ( .B1(P1_UWORD_REG_12__SCAN_IN), .B2(n21729), .A(n21749), 
        .ZN(n21747) );
  OAI21_X1 U23324 ( .B1(n21748), .B2(n21766), .A(n21747), .ZN(P1_U2949) );
  AOI21_X1 U23325 ( .B1(P1_LWORD_REG_12__SCAN_IN), .B2(n21729), .A(n21749), 
        .ZN(n21750) );
  OAI21_X1 U23326 ( .B1(n21751), .B2(n21766), .A(n21750), .ZN(P1_U2964) );
  INV_X1 U23327 ( .A(n21752), .ZN(n21753) );
  NOR2_X1 U23328 ( .A1(n21761), .A2(n21753), .ZN(n21756) );
  AOI21_X1 U23329 ( .B1(P1_UWORD_REG_13__SCAN_IN), .B2(n21729), .A(n21756), 
        .ZN(n21754) );
  OAI21_X1 U23330 ( .B1(n21755), .B2(n21766), .A(n21754), .ZN(P1_U2950) );
  AOI21_X1 U23331 ( .B1(P1_LWORD_REG_13__SCAN_IN), .B2(n21729), .A(n21756), 
        .ZN(n21757) );
  OAI21_X1 U23332 ( .B1(n21758), .B2(n21766), .A(n21757), .ZN(P1_U2965) );
  INV_X1 U23333 ( .A(n21759), .ZN(n21760) );
  NOR2_X1 U23334 ( .A1(n21761), .A2(n21760), .ZN(n21764) );
  AOI21_X1 U23335 ( .B1(P1_UWORD_REG_14__SCAN_IN), .B2(n21729), .A(n21764), 
        .ZN(n21762) );
  OAI21_X1 U23336 ( .B1(n21763), .B2(n21766), .A(n21762), .ZN(P1_U2951) );
  AOI21_X1 U23337 ( .B1(P1_LWORD_REG_14__SCAN_IN), .B2(n21729), .A(n21764), 
        .ZN(n21765) );
  OAI21_X1 U23338 ( .B1(n21767), .B2(n21766), .A(n21765), .ZN(P1_U2966) );
  INV_X1 U23339 ( .A(n22207), .ZN(n21768) );
  NAND2_X1 U23340 ( .A1(n21768), .A2(n21925), .ZN(n21770) );
  NOR2_X1 U23341 ( .A1(n21919), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n21894) );
  INV_X1 U23342 ( .A(n21894), .ZN(n21837) );
  OAI21_X1 U23343 ( .B1(n21770), .B2(n22214), .A(n21837), .ZN(n21777) );
  OR2_X1 U23344 ( .A1(n21821), .A2(n21771), .ZN(n21793) );
  NOR2_X1 U23345 ( .A1(n21793), .A2(n21938), .ZN(n21774) );
  NOR2_X1 U23346 ( .A1(n21772), .A2(n21917), .ZN(n21863) );
  INV_X1 U23347 ( .A(n21903), .ZN(n21896) );
  OR2_X1 U23348 ( .A1(n21904), .A2(n21896), .ZN(n21822) );
  INV_X1 U23349 ( .A(n21822), .ZN(n21779) );
  AOI22_X1 U23350 ( .A1(n21777), .A2(n21774), .B1(n21863), .B2(n21779), .ZN(
        n22211) );
  INV_X1 U23351 ( .A(n21935), .ZN(n21913) );
  NOR3_X1 U23352 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21788) );
  NAND2_X1 U23353 ( .A1(n21915), .A2(n21788), .ZN(n21775) );
  INV_X1 U23354 ( .A(n21775), .ZN(n22206) );
  AOI22_X1 U23355 ( .A1(n22207), .A2(n21944), .B1(n21934), .B2(n22206), .ZN(
        n21781) );
  INV_X1 U23356 ( .A(n21772), .ZN(n21773) );
  NOR2_X1 U23357 ( .A1(n21773), .A2(n21917), .ZN(n21839) );
  INV_X1 U23358 ( .A(n21774), .ZN(n21776) );
  AOI22_X1 U23359 ( .A1(n21777), .A2(n21776), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n21775), .ZN(n21778) );
  OAI211_X1 U23360 ( .C1(n21779), .C2(n21917), .A(n21886), .B(n21778), .ZN(
        n22208) );
  AOI22_X1 U23361 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n22208), .B1(
        n22214), .B2(n21901), .ZN(n21780) );
  OAI211_X1 U23362 ( .C1(n22211), .C2(n21913), .A(n21781), .B(n21780), .ZN(
        P1_U3033) );
  INV_X1 U23363 ( .A(n21793), .ZN(n21805) );
  INV_X1 U23364 ( .A(n21783), .ZN(n21916) );
  INV_X1 U23365 ( .A(n21788), .ZN(n21784) );
  NOR2_X1 U23366 ( .A1(n21915), .A2(n21784), .ZN(n22212) );
  AOI21_X1 U23367 ( .B1(n21805), .B2(n21916), .A(n22212), .ZN(n21785) );
  OAI22_X1 U23368 ( .A1(n21785), .A2(n21919), .B1(n21784), .B2(n21917), .ZN(
        n22213) );
  AOI22_X1 U23369 ( .A1(n21935), .A2(n22213), .B1(n21934), .B2(n22212), .ZN(
        n21790) );
  INV_X1 U23370 ( .A(n21809), .ZN(n21786) );
  OAI211_X1 U23371 ( .C1(n21786), .C2(n21936), .A(n21925), .B(n21785), .ZN(
        n21787) );
  OAI211_X1 U23372 ( .C1(n21925), .C2(n21788), .A(n21923), .B(n21787), .ZN(
        n22215) );
  AOI22_X1 U23373 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n22215), .B1(
        n22214), .B2(n21944), .ZN(n21789) );
  OAI211_X1 U23374 ( .C1(n21947), .C2(n22219), .A(n21790), .B(n21789), .ZN(
        P1_U3041) );
  NAND2_X1 U23375 ( .A1(n22219), .A2(n21925), .ZN(n21792) );
  OAI21_X1 U23376 ( .B1(n21792), .B2(n22226), .A(n21837), .ZN(n21796) );
  NOR2_X1 U23377 ( .A1(n21793), .A2(n14906), .ZN(n21798) );
  NOR2_X1 U23378 ( .A1(n21903), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21840) );
  AOI22_X1 U23379 ( .A1(n21796), .A2(n21798), .B1(n21840), .B2(n21863), .ZN(
        n22224) );
  INV_X1 U23380 ( .A(n21944), .ZN(n21881) );
  NOR3_X1 U23381 ( .A1(n21794), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n21811) );
  NAND2_X1 U23382 ( .A1(n21915), .A2(n21811), .ZN(n22218) );
  OAI22_X1 U23383 ( .A1(n22219), .A2(n21881), .B1(n21880), .B2(n22218), .ZN(
        n21795) );
  INV_X1 U23384 ( .A(n21795), .ZN(n21801) );
  INV_X1 U23385 ( .A(n21796), .ZN(n21799) );
  NOR2_X1 U23386 ( .A1(n21840), .A2(n21917), .ZN(n21843) );
  AOI21_X1 U23387 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n22218), .A(n21843), 
        .ZN(n21797) );
  OAI211_X1 U23388 ( .C1(n21799), .C2(n21798), .A(n21797), .B(n21886), .ZN(
        n22221) );
  AOI22_X1 U23389 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n22221), .B1(
        n22226), .B2(n21901), .ZN(n21800) );
  OAI211_X1 U23390 ( .C1(n22224), .C2(n21913), .A(n21801), .B(n21800), .ZN(
        P1_U3049) );
  INV_X1 U23391 ( .A(n21811), .ZN(n21806) );
  INV_X1 U23392 ( .A(n21802), .ZN(n21803) );
  NAND2_X1 U23393 ( .A1(n21809), .A2(n21803), .ZN(n21804) );
  NAND2_X1 U23394 ( .A1(n21804), .A2(n21925), .ZN(n21810) );
  NOR2_X1 U23395 ( .A1(n21915), .A2(n21806), .ZN(n22225) );
  AOI21_X1 U23396 ( .B1(n21805), .B2(n21853), .A(n22225), .ZN(n21813) );
  OAI22_X1 U23397 ( .A1(n21917), .A2(n21806), .B1(n21810), .B2(n21813), .ZN(
        n21807) );
  AOI22_X1 U23398 ( .A1(n22233), .A2(n21901), .B1(n21934), .B2(n22225), .ZN(
        n21817) );
  INV_X1 U23399 ( .A(n21810), .ZN(n21814) );
  OAI21_X1 U23400 ( .B1(n21876), .B2(n21811), .A(n21923), .ZN(n21812) );
  AOI21_X1 U23401 ( .B1(n21814), .B2(n21813), .A(n21812), .ZN(n21815) );
  AOI22_X1 U23402 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n22227), .B1(
        n22226), .B2(n21944), .ZN(n21816) );
  OAI211_X1 U23403 ( .C1(n22230), .C2(n21913), .A(n21817), .B(n21816), .ZN(
        P1_U3057) );
  NAND2_X1 U23404 ( .A1(n21819), .A2(n21818), .ZN(n21831) );
  OR2_X1 U23405 ( .A1(n21831), .A2(n21850), .ZN(n22243) );
  NAND2_X1 U23406 ( .A1(n21854), .A2(n14906), .ZN(n21823) );
  INV_X1 U23407 ( .A(n21839), .ZN(n21928) );
  OAI22_X1 U23408 ( .A1(n21823), .A2(n21919), .B1(n21928), .B2(n21822), .ZN(
        n22232) );
  NOR3_X1 U23409 ( .A1(n21900), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21833) );
  INV_X1 U23410 ( .A(n21833), .ZN(n21829) );
  NOR2_X1 U23411 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21829), .ZN(
        n22231) );
  AOI22_X1 U23412 ( .A1(n21935), .A2(n22232), .B1(n21934), .B2(n22231), .ZN(
        n21828) );
  OAI21_X1 U23413 ( .B1(n22166), .B2(n22233), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n21824) );
  AOI21_X1 U23414 ( .B1(n21824), .B2(n21823), .A(P1_STATE2_REG_3__SCAN_IN), 
        .ZN(n21826) );
  AOI22_X1 U23415 ( .A1(n22234), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n21944), .B2(n22233), .ZN(n21827) );
  OAI211_X1 U23416 ( .C1(n21947), .C2(n22243), .A(n21828), .B(n21827), .ZN(
        P1_U3065) );
  NOR2_X1 U23417 ( .A1(n21915), .A2(n21829), .ZN(n22237) );
  AOI21_X1 U23418 ( .B1(n21854), .B2(n21916), .A(n22237), .ZN(n21830) );
  OAI22_X1 U23419 ( .A1(n21830), .A2(n21919), .B1(n21829), .B2(n21917), .ZN(
        n22238) );
  AOI22_X1 U23420 ( .A1(n21935), .A2(n22238), .B1(n21934), .B2(n22237), .ZN(
        n21835) );
  OAI21_X1 U23421 ( .B1(n21831), .B2(n21936), .A(n21830), .ZN(n21832) );
  OAI221_X1 U23422 ( .B1(n21925), .B2(n21833), .C1(n21919), .C2(n21832), .A(
        n21923), .ZN(n22240) );
  AOI22_X1 U23423 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n22240), .B1(
        n22166), .B2(n21944), .ZN(n21834) );
  OAI211_X1 U23424 ( .C1(n21947), .C2(n22245), .A(n21835), .B(n21834), .ZN(
        P1_U3073) );
  NAND2_X1 U23425 ( .A1(n22245), .A2(n21925), .ZN(n21838) );
  OAI21_X1 U23426 ( .B1(n22253), .B2(n21838), .A(n21837), .ZN(n21845) );
  AND2_X1 U23427 ( .A1(n21854), .A2(n21938), .ZN(n21842) );
  AOI22_X1 U23428 ( .A1(n21845), .A2(n21842), .B1(n21840), .B2(n21839), .ZN(
        n22250) );
  NOR3_X1 U23429 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n21932), .ZN(n21847) );
  INV_X1 U23430 ( .A(n21847), .ZN(n22244) );
  OAI22_X1 U23431 ( .A1(n22245), .A2(n21881), .B1(n21880), .B2(n22244), .ZN(
        n21841) );
  INV_X1 U23432 ( .A(n21841), .ZN(n21849) );
  INV_X1 U23433 ( .A(n21842), .ZN(n21844) );
  AOI21_X1 U23434 ( .B1(n21845), .B2(n21844), .A(n21843), .ZN(n21846) );
  OAI211_X1 U23435 ( .C1(n21847), .C2(n21902), .A(n21942), .B(n21846), .ZN(
        n22247) );
  AOI22_X1 U23436 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n22247), .B1(
        n22253), .B2(n21901), .ZN(n21848) );
  OAI211_X1 U23437 ( .C1(n22250), .C2(n21913), .A(n21849), .B(n21848), .ZN(
        P1_U3081) );
  INV_X1 U23438 ( .A(n21852), .ZN(n22251) );
  AOI21_X1 U23439 ( .B1(n21854), .B2(n21853), .A(n22251), .ZN(n21856) );
  NOR2_X1 U23440 ( .A1(n21932), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21859) );
  INV_X1 U23441 ( .A(n21859), .ZN(n21855) );
  OAI22_X1 U23442 ( .A1(n21856), .A2(n21919), .B1(n21855), .B2(n21917), .ZN(
        n22252) );
  AOI22_X1 U23443 ( .A1(n21935), .A2(n22252), .B1(n22251), .B2(n21934), .ZN(
        n21861) );
  NAND2_X1 U23444 ( .A1(n21857), .A2(n21856), .ZN(n21858) );
  OAI221_X1 U23445 ( .B1(n21925), .B2(n21859), .C1(n21919), .C2(n21858), .A(
        n21923), .ZN(n22254) );
  AOI22_X1 U23446 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n22254), .B1(
        n22253), .B2(n21944), .ZN(n21860) );
  OAI211_X1 U23447 ( .C1(n21947), .C2(n22257), .A(n21861), .B(n21860), .ZN(
        P1_U3089) );
  INV_X1 U23448 ( .A(n21884), .ZN(n21864) );
  INV_X1 U23449 ( .A(n21863), .ZN(n21888) );
  INV_X1 U23450 ( .A(n21904), .ZN(n21897) );
  OAI33_X1 U23451 ( .A1(n21919), .A2(n21938), .A3(n21864), .B1(n21888), .B2(
        n21896), .B3(n21897), .ZN(n22259) );
  NOR3_X1 U23452 ( .A1(n21933), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21875) );
  INV_X1 U23453 ( .A(n21875), .ZN(n21871) );
  NOR2_X1 U23454 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21871), .ZN(
        n22258) );
  AOI22_X1 U23455 ( .A1(n21935), .A2(n11071), .B1(n21934), .B2(n22258), .ZN(
        n21869) );
  AOI21_X1 U23456 ( .B1(n22270), .B2(n22257), .A(n21936), .ZN(n21865) );
  AOI21_X1 U23457 ( .B1(n21884), .B2(n14906), .A(n21865), .ZN(n21866) );
  NOR2_X1 U23458 ( .A1(n21866), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21867) );
  AOI22_X1 U23459 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n22261), .B1(
        n22260), .B2(n21944), .ZN(n21868) );
  OAI211_X1 U23460 ( .C1(n21947), .C2(n22270), .A(n21869), .B(n21868), .ZN(
        P1_U3097) );
  NOR2_X1 U23461 ( .A1(n21915), .A2(n21871), .ZN(n22264) );
  AOI21_X1 U23462 ( .B1(n21884), .B2(n21916), .A(n22264), .ZN(n21872) );
  OAI22_X1 U23463 ( .A1(n21872), .A2(n21919), .B1(n21871), .B2(n21917), .ZN(
        n22265) );
  AOI22_X1 U23464 ( .A1(n21935), .A2(n22265), .B1(n21934), .B2(n22264), .ZN(
        n21878) );
  OAI21_X1 U23465 ( .B1(n21873), .B2(n21936), .A(n21872), .ZN(n21874) );
  OAI221_X1 U23466 ( .B1(n21876), .B2(n21875), .C1(n21919), .C2(n21874), .A(
        n21923), .ZN(n22267) );
  INV_X1 U23467 ( .A(n22270), .ZN(n22176) );
  AOI22_X1 U23468 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n22267), .B1(
        n22176), .B2(n21944), .ZN(n21877) );
  OAI211_X1 U23469 ( .C1(n21947), .C2(n22279), .A(n21878), .B(n21877), .ZN(
        P1_U3105) );
  NAND2_X1 U23470 ( .A1(n21915), .A2(n21879), .ZN(n22271) );
  OAI22_X1 U23471 ( .A1(n22279), .A2(n21881), .B1(n21880), .B2(n22271), .ZN(
        n21882) );
  INV_X1 U23472 ( .A(n21882), .ZN(n21892) );
  NAND2_X1 U23473 ( .A1(n22273), .A2(n22279), .ZN(n21883) );
  AOI21_X1 U23474 ( .B1(n21883), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n21919), 
        .ZN(n21887) );
  NAND2_X1 U23475 ( .A1(n21884), .A2(n21938), .ZN(n21889) );
  AOI22_X1 U23476 ( .A1(n21887), .A2(n21889), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n22271), .ZN(n21885) );
  NAND2_X1 U23477 ( .A1(n21896), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n21929) );
  NAND2_X1 U23478 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n21929), .ZN(n21941) );
  NAND3_X1 U23479 ( .A1(n21886), .A2(n21885), .A3(n21941), .ZN(n22276) );
  INV_X1 U23480 ( .A(n21887), .ZN(n21890) );
  OAI22_X1 U23481 ( .A1(n21890), .A2(n21889), .B1(n21888), .B2(n21929), .ZN(
        n22275) );
  AOI22_X1 U23482 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n22276), .B1(
        n21935), .B2(n22275), .ZN(n21891) );
  OAI211_X1 U23483 ( .C1(n21947), .C2(n22273), .A(n21892), .B(n21891), .ZN(
        P1_U3113) );
  NOR2_X2 U23484 ( .A1(n21921), .A2(n21893), .ZN(n22291) );
  NOR2_X1 U23485 ( .A1(n22291), .A2(n21919), .ZN(n21895) );
  AOI21_X1 U23486 ( .B1(n21895), .B2(n21910), .A(n21894), .ZN(n21909) );
  INV_X1 U23487 ( .A(n21909), .ZN(n21899) );
  NOR2_X1 U23488 ( .A1(n21931), .A2(n21938), .ZN(n21908) );
  NOR3_X1 U23489 ( .A1(n21928), .A2(n21897), .A3(n21896), .ZN(n21898) );
  NOR3_X1 U23490 ( .A1(n21900), .A2(n21933), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n21924) );
  INV_X1 U23491 ( .A(n21924), .ZN(n21918) );
  NOR2_X1 U23492 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21918), .ZN(
        n22281) );
  AOI22_X1 U23493 ( .A1(n22291), .A2(n21901), .B1(n21934), .B2(n22281), .ZN(
        n21912) );
  INV_X1 U23494 ( .A(n22281), .ZN(n21906) );
  AOI21_X1 U23495 ( .B1(n21904), .B2(n21903), .A(n21917), .ZN(n21905) );
  AOI21_X1 U23496 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n21906), .A(n21905), 
        .ZN(n21907) );
  OAI211_X1 U23497 ( .C1(n21909), .C2(n21908), .A(n21942), .B(n21907), .ZN(
        n22284) );
  AOI22_X1 U23498 ( .A1(n22284), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n21944), .B2(n22283), .ZN(n21911) );
  OAI211_X1 U23499 ( .C1(n22288), .C2(n21913), .A(n21912), .B(n21911), .ZN(
        P1_U3129) );
  INV_X1 U23500 ( .A(n21931), .ZN(n21939) );
  NOR2_X1 U23501 ( .A1(n21915), .A2(n21918), .ZN(n22289) );
  AOI21_X1 U23502 ( .B1(n21939), .B2(n21916), .A(n22289), .ZN(n21920) );
  OAI22_X1 U23503 ( .A1(n21920), .A2(n21919), .B1(n21918), .B2(n21917), .ZN(
        n22290) );
  AOI22_X1 U23504 ( .A1(n21935), .A2(n22290), .B1(n21934), .B2(n22289), .ZN(
        n21927) );
  OAI211_X1 U23505 ( .C1(n21921), .C2(n21936), .A(n21925), .B(n21920), .ZN(
        n21922) );
  OAI211_X1 U23506 ( .C1(n21925), .C2(n21924), .A(n21923), .B(n21922), .ZN(
        n22292) );
  AOI22_X1 U23507 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n22292), .B1(
        n22291), .B2(n21944), .ZN(n21926) );
  OAI211_X1 U23508 ( .C1(n21947), .C2(n22295), .A(n21927), .B(n21926), .ZN(
        P1_U3137) );
  NAND2_X1 U23509 ( .A1(n21938), .A2(n21925), .ZN(n21930) );
  OAI22_X1 U23510 ( .A1(n21931), .A2(n21930), .B1(n21929), .B2(n21928), .ZN(
        n22298) );
  NOR3_X2 U23511 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n21933), .A3(
        n21932), .ZN(n22296) );
  AOI22_X1 U23512 ( .A1(n21935), .A2(n22298), .B1(n21934), .B2(n22296), .ZN(
        n21946) );
  AOI21_X1 U23513 ( .B1(n22305), .B2(n22295), .A(n21936), .ZN(n21937) );
  AOI21_X1 U23514 ( .B1(n21939), .B2(n21938), .A(n21937), .ZN(n21940) );
  NOR2_X1 U23515 ( .A1(n21940), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n21943) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n22302), .B1(
        n22301), .B2(n21944), .ZN(n21945) );
  OAI211_X1 U23517 ( .C1(n21947), .C2(n22305), .A(n21946), .B(n21945), .ZN(
        P1_U3145) );
  AOI22_X1 U23518 ( .A1(n22207), .A2(n21985), .B1(n21984), .B2(n22206), .ZN(
        n21949) );
  AOI22_X1 U23519 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n22208), .B1(
        n22214), .B2(n21977), .ZN(n21948) );
  OAI211_X1 U23520 ( .C1(n22211), .C2(n21980), .A(n21949), .B(n21948), .ZN(
        P1_U3034) );
  INV_X1 U23521 ( .A(n21977), .ZN(n21988) );
  AOI22_X1 U23522 ( .A1(n21984), .A2(n22212), .B1(n22213), .B2(n21983), .ZN(
        n21951) );
  AOI22_X1 U23523 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n22215), .B1(
        n22214), .B2(n21985), .ZN(n21950) );
  OAI211_X1 U23524 ( .C1(n21988), .C2(n22219), .A(n21951), .B(n21950), .ZN(
        P1_U3042) );
  INV_X1 U23525 ( .A(n21985), .ZN(n21976) );
  INV_X1 U23526 ( .A(n21984), .ZN(n21970) );
  OAI22_X1 U23527 ( .A1(n22219), .A2(n21976), .B1(n21970), .B2(n22218), .ZN(
        n21952) );
  INV_X1 U23528 ( .A(n21952), .ZN(n21954) );
  AOI22_X1 U23529 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n22221), .B1(
        n22226), .B2(n21977), .ZN(n21953) );
  OAI211_X1 U23530 ( .C1(n22224), .C2(n21980), .A(n21954), .B(n21953), .ZN(
        P1_U3050) );
  AOI22_X1 U23531 ( .A1(n22226), .A2(n21985), .B1(n21984), .B2(n22225), .ZN(
        n21956) );
  AOI22_X1 U23532 ( .A1(n22227), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n22233), .B2(n21977), .ZN(n21955) );
  OAI211_X1 U23533 ( .C1(n22230), .C2(n21980), .A(n21956), .B(n21955), .ZN(
        P1_U3058) );
  AOI22_X1 U23534 ( .A1(n21984), .A2(n22231), .B1(n21983), .B2(n22232), .ZN(
        n21958) );
  AOI22_X1 U23535 ( .A1(n22234), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n22233), .B2(n21985), .ZN(n21957) );
  OAI211_X1 U23536 ( .C1(n21988), .C2(n22243), .A(n21958), .B(n21957), .ZN(
        P1_U3066) );
  AOI22_X1 U23537 ( .A1(n21984), .A2(n22237), .B1(n21983), .B2(n22238), .ZN(
        n21960) );
  AOI22_X1 U23538 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n22240), .B1(
        n22166), .B2(n21985), .ZN(n21959) );
  OAI211_X1 U23539 ( .C1(n21988), .C2(n22245), .A(n21960), .B(n21959), .ZN(
        P1_U3074) );
  OAI22_X1 U23540 ( .A1(n22245), .A2(n21976), .B1(n21970), .B2(n22244), .ZN(
        n21961) );
  INV_X1 U23541 ( .A(n21961), .ZN(n21963) );
  AOI22_X1 U23542 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n22247), .B1(
        n22253), .B2(n21977), .ZN(n21962) );
  OAI211_X1 U23543 ( .C1(n22250), .C2(n21980), .A(n21963), .B(n21962), .ZN(
        P1_U3082) );
  AOI22_X1 U23544 ( .A1(n21984), .A2(n22251), .B1(n21983), .B2(n22252), .ZN(
        n21965) );
  AOI22_X1 U23545 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n22254), .B1(
        n22253), .B2(n21985), .ZN(n21964) );
  OAI211_X1 U23546 ( .C1(n21988), .C2(n22257), .A(n21965), .B(n21964), .ZN(
        P1_U3090) );
  AOI22_X1 U23547 ( .A1(n11071), .A2(n21983), .B1(n21984), .B2(n22258), .ZN(
        n21967) );
  AOI22_X1 U23548 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n22261), .B1(
        n22260), .B2(n21985), .ZN(n21966) );
  OAI211_X1 U23549 ( .C1(n21988), .C2(n22270), .A(n21967), .B(n21966), .ZN(
        P1_U3098) );
  AOI22_X1 U23550 ( .A1(n21984), .A2(n22264), .B1(n21983), .B2(n22265), .ZN(
        n21969) );
  INV_X1 U23551 ( .A(n22279), .ZN(n22266) );
  AOI22_X1 U23552 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n22267), .B1(
        n22266), .B2(n21977), .ZN(n21968) );
  OAI211_X1 U23553 ( .C1(n21976), .C2(n22270), .A(n21969), .B(n21968), .ZN(
        P1_U3106) );
  OAI22_X1 U23554 ( .A1(n22273), .A2(n21988), .B1(n21970), .B2(n22271), .ZN(
        n21971) );
  INV_X1 U23555 ( .A(n21971), .ZN(n21973) );
  AOI22_X1 U23556 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n22276), .B1(
        n21983), .B2(n22275), .ZN(n21972) );
  OAI211_X1 U23557 ( .C1(n21976), .C2(n22279), .A(n21973), .B(n21972), .ZN(
        P1_U3114) );
  AOI22_X1 U23558 ( .A1(n21984), .A2(n22183), .B1(n21983), .B2(n22184), .ZN(
        n21975) );
  AOI22_X1 U23559 ( .A1(n22185), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n22283), .B2(n21977), .ZN(n21974) );
  OAI211_X1 U23560 ( .C1(n21976), .C2(n22273), .A(n21975), .B(n21974), .ZN(
        P1_U3122) );
  AOI22_X1 U23561 ( .A1(n22291), .A2(n21977), .B1(n21984), .B2(n22281), .ZN(
        n21979) );
  AOI22_X1 U23562 ( .A1(n22284), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n21985), .B2(n22283), .ZN(n21978) );
  OAI211_X1 U23563 ( .C1(n22288), .C2(n21980), .A(n21979), .B(n21978), .ZN(
        P1_U3130) );
  AOI22_X1 U23564 ( .A1(n21984), .A2(n22289), .B1(n21983), .B2(n22290), .ZN(
        n21982) );
  AOI22_X1 U23565 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n22292), .B1(
        n22291), .B2(n21985), .ZN(n21981) );
  OAI211_X1 U23566 ( .C1(n21988), .C2(n22295), .A(n21982), .B(n21981), .ZN(
        P1_U3138) );
  AOI22_X1 U23567 ( .A1(n21984), .A2(n22296), .B1(n21983), .B2(n22298), .ZN(
        n21987) );
  AOI22_X1 U23568 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n22302), .B1(
        n22301), .B2(n21985), .ZN(n21986) );
  OAI211_X1 U23569 ( .C1(n21988), .C2(n22305), .A(n21987), .B(n21986), .ZN(
        P1_U3146) );
  AOI22_X1 U23570 ( .A1(n22207), .A2(n22024), .B1(n22023), .B2(n22206), .ZN(
        n21990) );
  AOI22_X1 U23571 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n22208), .B1(
        n22214), .B2(n22016), .ZN(n21989) );
  OAI211_X1 U23572 ( .C1(n22211), .C2(n22019), .A(n21990), .B(n21989), .ZN(
        P1_U3035) );
  AOI22_X1 U23573 ( .A1(n22023), .A2(n22212), .B1(n22213), .B2(n22022), .ZN(
        n21992) );
  AOI22_X1 U23574 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n22215), .B1(
        n22214), .B2(n22024), .ZN(n21991) );
  OAI211_X1 U23575 ( .C1(n22027), .C2(n22219), .A(n21992), .B(n21991), .ZN(
        P1_U3043) );
  INV_X1 U23576 ( .A(n22024), .ZN(n22015) );
  INV_X1 U23577 ( .A(n22023), .ZN(n22011) );
  OAI22_X1 U23578 ( .A1(n22219), .A2(n22015), .B1(n22011), .B2(n22218), .ZN(
        n21993) );
  INV_X1 U23579 ( .A(n21993), .ZN(n21995) );
  AOI22_X1 U23580 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n22221), .B1(
        n22226), .B2(n22016), .ZN(n21994) );
  OAI211_X1 U23581 ( .C1(n22224), .C2(n22019), .A(n21995), .B(n21994), .ZN(
        P1_U3051) );
  AOI22_X1 U23582 ( .A1(n22226), .A2(n22024), .B1(n22023), .B2(n22225), .ZN(
        n21997) );
  AOI22_X1 U23583 ( .A1(n22227), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n22233), .B2(n22016), .ZN(n21996) );
  OAI211_X1 U23584 ( .C1(n22230), .C2(n22019), .A(n21997), .B(n21996), .ZN(
        P1_U3059) );
  AOI22_X1 U23585 ( .A1(n22023), .A2(n22231), .B1(n22022), .B2(n22232), .ZN(
        n21999) );
  AOI22_X1 U23586 ( .A1(n22234), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n22233), .B2(n22024), .ZN(n21998) );
  OAI211_X1 U23587 ( .C1(n22027), .C2(n22243), .A(n21999), .B(n21998), .ZN(
        P1_U3067) );
  AOI22_X1 U23588 ( .A1(n22023), .A2(n22237), .B1(n22022), .B2(n22238), .ZN(
        n22001) );
  AOI22_X1 U23589 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n22240), .B1(
        n22166), .B2(n22024), .ZN(n22000) );
  OAI211_X1 U23590 ( .C1(n22027), .C2(n22245), .A(n22001), .B(n22000), .ZN(
        P1_U3075) );
  OAI22_X1 U23591 ( .A1(n22245), .A2(n22015), .B1(n22011), .B2(n22244), .ZN(
        n22002) );
  INV_X1 U23592 ( .A(n22002), .ZN(n22004) );
  AOI22_X1 U23593 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n22247), .B1(
        n22253), .B2(n22016), .ZN(n22003) );
  OAI211_X1 U23594 ( .C1(n22250), .C2(n22019), .A(n22004), .B(n22003), .ZN(
        P1_U3083) );
  AOI22_X1 U23595 ( .A1(n22023), .A2(n22251), .B1(n22022), .B2(n22252), .ZN(
        n22006) );
  AOI22_X1 U23596 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n22254), .B1(
        n22253), .B2(n22024), .ZN(n22005) );
  OAI211_X1 U23597 ( .C1(n22027), .C2(n22257), .A(n22006), .B(n22005), .ZN(
        P1_U3091) );
  AOI22_X1 U23598 ( .A1(n11071), .A2(n22022), .B1(n22023), .B2(n22258), .ZN(
        n22008) );
  AOI22_X1 U23599 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n22261), .B1(
        n22260), .B2(n22024), .ZN(n22007) );
  OAI211_X1 U23600 ( .C1(n22027), .C2(n22270), .A(n22008), .B(n22007), .ZN(
        P1_U3099) );
  AOI22_X1 U23601 ( .A1(n22023), .A2(n22264), .B1(n22022), .B2(n22265), .ZN(
        n22010) );
  AOI22_X1 U23602 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n22267), .B1(
        n22176), .B2(n22024), .ZN(n22009) );
  OAI211_X1 U23603 ( .C1(n22027), .C2(n22279), .A(n22010), .B(n22009), .ZN(
        P1_U3107) );
  OAI22_X1 U23604 ( .A1(n22273), .A2(n22027), .B1(n22011), .B2(n22271), .ZN(
        n22012) );
  INV_X1 U23605 ( .A(n22012), .ZN(n22014) );
  AOI22_X1 U23606 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n22276), .B1(
        n22022), .B2(n22275), .ZN(n22013) );
  OAI211_X1 U23607 ( .C1(n22015), .C2(n22279), .A(n22014), .B(n22013), .ZN(
        P1_U3115) );
  AOI22_X1 U23608 ( .A1(n22291), .A2(n22016), .B1(n22023), .B2(n22281), .ZN(
        n22018) );
  AOI22_X1 U23609 ( .A1(n22284), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n22024), .B2(n22283), .ZN(n22017) );
  OAI211_X1 U23610 ( .C1(n22288), .C2(n22019), .A(n22018), .B(n22017), .ZN(
        P1_U3131) );
  AOI22_X1 U23611 ( .A1(n22023), .A2(n22289), .B1(n22022), .B2(n22290), .ZN(
        n22021) );
  AOI22_X1 U23612 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n22292), .B1(
        n22291), .B2(n22024), .ZN(n22020) );
  OAI211_X1 U23613 ( .C1(n22027), .C2(n22295), .A(n22021), .B(n22020), .ZN(
        P1_U3139) );
  AOI22_X1 U23614 ( .A1(n22023), .A2(n22296), .B1(n22022), .B2(n22298), .ZN(
        n22026) );
  AOI22_X1 U23615 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n22302), .B1(
        n22301), .B2(n22024), .ZN(n22025) );
  OAI211_X1 U23616 ( .C1(n22027), .C2(n22305), .A(n22026), .B(n22025), .ZN(
        P1_U3147) );
  AOI22_X1 U23617 ( .A1(n22207), .A2(n22062), .B1(n22061), .B2(n22206), .ZN(
        n22029) );
  AOI22_X1 U23618 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n22208), .B1(
        n22214), .B2(n22054), .ZN(n22028) );
  OAI211_X1 U23619 ( .C1(n22211), .C2(n22057), .A(n22029), .B(n22028), .ZN(
        P1_U3036) );
  AOI22_X1 U23620 ( .A1(n22061), .A2(n22212), .B1(n22213), .B2(n22060), .ZN(
        n22031) );
  AOI22_X1 U23621 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n22215), .B1(
        n22214), .B2(n22062), .ZN(n22030) );
  OAI211_X1 U23622 ( .C1(n22065), .C2(n22219), .A(n22031), .B(n22030), .ZN(
        P1_U3044) );
  INV_X1 U23623 ( .A(n22218), .ZN(n22158) );
  AOI22_X1 U23624 ( .A1(n22226), .A2(n22054), .B1(n22061), .B2(n22158), .ZN(
        n22033) );
  INV_X1 U23625 ( .A(n22219), .ZN(n22159) );
  AOI22_X1 U23626 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n22221), .B1(
        n22159), .B2(n22062), .ZN(n22032) );
  OAI211_X1 U23627 ( .C1(n22224), .C2(n22057), .A(n22033), .B(n22032), .ZN(
        P1_U3052) );
  AOI22_X1 U23628 ( .A1(n22233), .A2(n22054), .B1(n22061), .B2(n22225), .ZN(
        n22035) );
  AOI22_X1 U23629 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n22227), .B1(
        n22226), .B2(n22062), .ZN(n22034) );
  OAI211_X1 U23630 ( .C1(n22230), .C2(n22057), .A(n22035), .B(n22034), .ZN(
        P1_U3060) );
  AOI22_X1 U23631 ( .A1(n22061), .A2(n22231), .B1(n22060), .B2(n22232), .ZN(
        n22037) );
  AOI22_X1 U23632 ( .A1(n22234), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n22233), .B2(n22062), .ZN(n22036) );
  OAI211_X1 U23633 ( .C1(n22065), .C2(n22243), .A(n22037), .B(n22036), .ZN(
        P1_U3068) );
  AOI22_X1 U23634 ( .A1(n22061), .A2(n22237), .B1(n22060), .B2(n22238), .ZN(
        n22039) );
  AOI22_X1 U23635 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n22240), .B1(
        n22166), .B2(n22062), .ZN(n22038) );
  OAI211_X1 U23636 ( .C1(n22065), .C2(n22245), .A(n22039), .B(n22038), .ZN(
        P1_U3076) );
  INV_X1 U23637 ( .A(n22062), .ZN(n22053) );
  INV_X1 U23638 ( .A(n22061), .ZN(n22049) );
  OAI22_X1 U23639 ( .A1(n22245), .A2(n22053), .B1(n22049), .B2(n22244), .ZN(
        n22040) );
  INV_X1 U23640 ( .A(n22040), .ZN(n22042) );
  AOI22_X1 U23641 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n22247), .B1(
        n22253), .B2(n22054), .ZN(n22041) );
  OAI211_X1 U23642 ( .C1(n22250), .C2(n22057), .A(n22042), .B(n22041), .ZN(
        P1_U3084) );
  AOI22_X1 U23643 ( .A1(n22061), .A2(n22251), .B1(n22060), .B2(n22252), .ZN(
        n22044) );
  AOI22_X1 U23644 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n22254), .B1(
        n22253), .B2(n22062), .ZN(n22043) );
  OAI211_X1 U23645 ( .C1(n22065), .C2(n22257), .A(n22044), .B(n22043), .ZN(
        P1_U3092) );
  AOI22_X1 U23646 ( .A1(n11071), .A2(n22060), .B1(n22061), .B2(n22258), .ZN(
        n22046) );
  AOI22_X1 U23647 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n22261), .B1(
        n22260), .B2(n22062), .ZN(n22045) );
  OAI211_X1 U23648 ( .C1(n22065), .C2(n22270), .A(n22046), .B(n22045), .ZN(
        P1_U3100) );
  AOI22_X1 U23649 ( .A1(n22061), .A2(n22264), .B1(n22060), .B2(n22265), .ZN(
        n22048) );
  AOI22_X1 U23650 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n22267), .B1(
        n22176), .B2(n22062), .ZN(n22047) );
  OAI211_X1 U23651 ( .C1(n22065), .C2(n22279), .A(n22048), .B(n22047), .ZN(
        P1_U3108) );
  OAI22_X1 U23652 ( .A1(n22273), .A2(n22065), .B1(n22049), .B2(n22271), .ZN(
        n22050) );
  INV_X1 U23653 ( .A(n22050), .ZN(n22052) );
  AOI22_X1 U23654 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n22276), .B1(
        n22060), .B2(n22275), .ZN(n22051) );
  OAI211_X1 U23655 ( .C1(n22053), .C2(n22279), .A(n22052), .B(n22051), .ZN(
        P1_U3116) );
  AOI22_X1 U23656 ( .A1(n22291), .A2(n22054), .B1(n22061), .B2(n22281), .ZN(
        n22056) );
  AOI22_X1 U23657 ( .A1(n22284), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n22062), .B2(n22283), .ZN(n22055) );
  OAI211_X1 U23658 ( .C1(n22288), .C2(n22057), .A(n22056), .B(n22055), .ZN(
        P1_U3132) );
  AOI22_X1 U23659 ( .A1(n22061), .A2(n22289), .B1(n22060), .B2(n22290), .ZN(
        n22059) );
  AOI22_X1 U23660 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n22292), .B1(
        n22291), .B2(n22062), .ZN(n22058) );
  OAI211_X1 U23661 ( .C1(n22065), .C2(n22295), .A(n22059), .B(n22058), .ZN(
        P1_U3140) );
  AOI22_X1 U23662 ( .A1(n22061), .A2(n22296), .B1(n22060), .B2(n22298), .ZN(
        n22064) );
  AOI22_X1 U23663 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n22302), .B1(
        n22301), .B2(n22062), .ZN(n22063) );
  OAI211_X1 U23664 ( .C1(n22065), .C2(n22305), .A(n22064), .B(n22063), .ZN(
        P1_U3148) );
  AOI22_X1 U23665 ( .A1(n22207), .A2(n22096), .B1(n22100), .B2(n22206), .ZN(
        n22067) );
  AOI22_X1 U23666 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n22208), .B1(
        n22214), .B2(n22102), .ZN(n22066) );
  OAI211_X1 U23667 ( .C1(n22211), .C2(n22093), .A(n22067), .B(n22066), .ZN(
        P1_U3037) );
  AOI22_X1 U23668 ( .A1(n22101), .A2(n22213), .B1(n22100), .B2(n22212), .ZN(
        n22069) );
  AOI22_X1 U23669 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n22215), .B1(
        n22214), .B2(n22096), .ZN(n22068) );
  OAI211_X1 U23670 ( .C1(n22099), .C2(n22219), .A(n22069), .B(n22068), .ZN(
        P1_U3045) );
  AOI22_X1 U23671 ( .A1(n22226), .A2(n22102), .B1(n22100), .B2(n22158), .ZN(
        n22071) );
  AOI22_X1 U23672 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n22221), .B1(
        n22159), .B2(n22096), .ZN(n22070) );
  OAI211_X1 U23673 ( .C1(n22224), .C2(n22093), .A(n22071), .B(n22070), .ZN(
        P1_U3053) );
  AOI22_X1 U23674 ( .A1(n22233), .A2(n22102), .B1(n22100), .B2(n22225), .ZN(
        n22073) );
  AOI22_X1 U23675 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n22227), .B1(
        n22226), .B2(n22096), .ZN(n22072) );
  OAI211_X1 U23676 ( .C1(n22230), .C2(n22093), .A(n22073), .B(n22072), .ZN(
        P1_U3061) );
  AOI22_X1 U23677 ( .A1(n22101), .A2(n22232), .B1(n22100), .B2(n22231), .ZN(
        n22075) );
  AOI22_X1 U23678 ( .A1(n22234), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n22233), .B2(n22096), .ZN(n22074) );
  OAI211_X1 U23679 ( .C1(n22099), .C2(n22243), .A(n22075), .B(n22074), .ZN(
        P1_U3069) );
  AOI22_X1 U23680 ( .A1(n22101), .A2(n22238), .B1(n22100), .B2(n22237), .ZN(
        n22077) );
  AOI22_X1 U23681 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n22240), .B1(
        n22166), .B2(n22096), .ZN(n22076) );
  OAI211_X1 U23682 ( .C1(n22099), .C2(n22245), .A(n22077), .B(n22076), .ZN(
        P1_U3077) );
  INV_X1 U23683 ( .A(n22096), .ZN(n22105) );
  INV_X1 U23684 ( .A(n22100), .ZN(n22087) );
  OAI22_X1 U23685 ( .A1(n22245), .A2(n22105), .B1(n22087), .B2(n22244), .ZN(
        n22078) );
  INV_X1 U23686 ( .A(n22078), .ZN(n22080) );
  AOI22_X1 U23687 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n22247), .B1(
        n22253), .B2(n22102), .ZN(n22079) );
  OAI211_X1 U23688 ( .C1(n22250), .C2(n22093), .A(n22080), .B(n22079), .ZN(
        P1_U3085) );
  AOI22_X1 U23689 ( .A1(n22101), .A2(n22252), .B1(n22251), .B2(n22100), .ZN(
        n22082) );
  AOI22_X1 U23690 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n22254), .B1(
        n22253), .B2(n22096), .ZN(n22081) );
  OAI211_X1 U23691 ( .C1(n22099), .C2(n22257), .A(n22082), .B(n22081), .ZN(
        P1_U3093) );
  AOI22_X1 U23692 ( .A1(n11071), .A2(n22101), .B1(n22100), .B2(n22258), .ZN(
        n22084) );
  AOI22_X1 U23693 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n22261), .B1(
        n22260), .B2(n22096), .ZN(n22083) );
  OAI211_X1 U23694 ( .C1(n22099), .C2(n22270), .A(n22084), .B(n22083), .ZN(
        P1_U3101) );
  AOI22_X1 U23695 ( .A1(n22101), .A2(n22265), .B1(n22100), .B2(n22264), .ZN(
        n22086) );
  AOI22_X1 U23696 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n22267), .B1(
        n22266), .B2(n22102), .ZN(n22085) );
  OAI211_X1 U23697 ( .C1(n22105), .C2(n22270), .A(n22086), .B(n22085), .ZN(
        P1_U3109) );
  OAI22_X1 U23698 ( .A1(n22273), .A2(n22099), .B1(n22087), .B2(n22271), .ZN(
        n22088) );
  INV_X1 U23699 ( .A(n22088), .ZN(n22090) );
  AOI22_X1 U23700 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n22276), .B1(
        n22101), .B2(n22275), .ZN(n22089) );
  OAI211_X1 U23701 ( .C1(n22105), .C2(n22279), .A(n22090), .B(n22089), .ZN(
        P1_U3117) );
  AOI22_X1 U23702 ( .A1(n22291), .A2(n22102), .B1(n22100), .B2(n22281), .ZN(
        n22092) );
  AOI22_X1 U23703 ( .A1(n22284), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n22096), .B2(n22283), .ZN(n22091) );
  OAI211_X1 U23704 ( .C1(n22288), .C2(n22093), .A(n22092), .B(n22091), .ZN(
        P1_U3133) );
  AOI22_X1 U23705 ( .A1(n22101), .A2(n22290), .B1(n22100), .B2(n22289), .ZN(
        n22095) );
  AOI22_X1 U23706 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n22292), .B1(
        n22291), .B2(n22096), .ZN(n22094) );
  OAI211_X1 U23707 ( .C1(n22099), .C2(n22295), .A(n22095), .B(n22094), .ZN(
        P1_U3141) );
  AOI22_X1 U23708 ( .A1(n22101), .A2(n22298), .B1(n22100), .B2(n22296), .ZN(
        n22098) );
  AOI22_X1 U23709 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n22302), .B1(
        n22301), .B2(n22096), .ZN(n22097) );
  OAI211_X1 U23710 ( .C1(n22099), .C2(n22305), .A(n22098), .B(n22097), .ZN(
        P1_U3149) );
  AOI22_X1 U23711 ( .A1(n22101), .A2(n22199), .B1(n22197), .B2(n22100), .ZN(
        n22104) );
  AOI22_X1 U23712 ( .A1(n22202), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n22207), .B2(n22102), .ZN(n22103) );
  OAI211_X1 U23713 ( .C1(n22105), .C2(n22305), .A(n22104), .B(n22103), .ZN(
        P1_U3157) );
  AOI22_X1 U23714 ( .A1(n22207), .A2(n22140), .B1(n22139), .B2(n22206), .ZN(
        n22107) );
  AOI22_X1 U23715 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n22208), .B1(
        n22214), .B2(n22132), .ZN(n22106) );
  OAI211_X1 U23716 ( .C1(n22211), .C2(n22135), .A(n22107), .B(n22106), .ZN(
        P1_U3038) );
  AOI22_X1 U23717 ( .A1(n22139), .A2(n22212), .B1(n22213), .B2(n22138), .ZN(
        n22109) );
  AOI22_X1 U23718 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n22215), .B1(
        n22214), .B2(n22140), .ZN(n22108) );
  OAI211_X1 U23719 ( .C1(n22143), .C2(n22219), .A(n22109), .B(n22108), .ZN(
        P1_U3046) );
  AOI22_X1 U23720 ( .A1(n22226), .A2(n22132), .B1(n22139), .B2(n22158), .ZN(
        n22111) );
  AOI22_X1 U23721 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n22221), .B1(
        n22159), .B2(n22140), .ZN(n22110) );
  OAI211_X1 U23722 ( .C1(n22224), .C2(n22135), .A(n22111), .B(n22110), .ZN(
        P1_U3054) );
  AOI22_X1 U23723 ( .A1(n22226), .A2(n22140), .B1(n22139), .B2(n22225), .ZN(
        n22113) );
  AOI22_X1 U23724 ( .A1(n22227), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n22233), .B2(n22132), .ZN(n22112) );
  OAI211_X1 U23725 ( .C1(n22230), .C2(n22135), .A(n22113), .B(n22112), .ZN(
        P1_U3062) );
  AOI22_X1 U23726 ( .A1(n22139), .A2(n22231), .B1(n22138), .B2(n22232), .ZN(
        n22115) );
  AOI22_X1 U23727 ( .A1(n22234), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n22233), .B2(n22140), .ZN(n22114) );
  OAI211_X1 U23728 ( .C1(n22143), .C2(n22243), .A(n22115), .B(n22114), .ZN(
        P1_U3070) );
  INV_X1 U23729 ( .A(n22140), .ZN(n22131) );
  AOI22_X1 U23730 ( .A1(n22139), .A2(n22237), .B1(n22138), .B2(n22238), .ZN(
        n22117) );
  INV_X1 U23731 ( .A(n22245), .ZN(n22239) );
  AOI22_X1 U23732 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n22240), .B1(
        n22239), .B2(n22132), .ZN(n22116) );
  OAI211_X1 U23733 ( .C1(n22131), .C2(n22243), .A(n22117), .B(n22116), .ZN(
        P1_U3078) );
  INV_X1 U23734 ( .A(n22139), .ZN(n22127) );
  OAI22_X1 U23735 ( .A1(n22245), .A2(n22131), .B1(n22127), .B2(n22244), .ZN(
        n22118) );
  INV_X1 U23736 ( .A(n22118), .ZN(n22120) );
  AOI22_X1 U23737 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n22247), .B1(
        n22253), .B2(n22132), .ZN(n22119) );
  OAI211_X1 U23738 ( .C1(n22250), .C2(n22135), .A(n22120), .B(n22119), .ZN(
        P1_U3086) );
  AOI22_X1 U23739 ( .A1(n22139), .A2(n22251), .B1(n22138), .B2(n22252), .ZN(
        n22122) );
  AOI22_X1 U23740 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n22254), .B1(
        n22253), .B2(n22140), .ZN(n22121) );
  OAI211_X1 U23741 ( .C1(n22143), .C2(n22257), .A(n22122), .B(n22121), .ZN(
        P1_U3094) );
  AOI22_X1 U23742 ( .A1(n11071), .A2(n22138), .B1(n22258), .B2(n22139), .ZN(
        n22124) );
  AOI22_X1 U23743 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n22261), .B1(
        n22260), .B2(n22140), .ZN(n22123) );
  OAI211_X1 U23744 ( .C1(n22143), .C2(n22270), .A(n22124), .B(n22123), .ZN(
        P1_U3102) );
  AOI22_X1 U23745 ( .A1(n22139), .A2(n22264), .B1(n22138), .B2(n22265), .ZN(
        n22126) );
  AOI22_X1 U23746 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n22267), .B1(
        n22266), .B2(n22132), .ZN(n22125) );
  OAI211_X1 U23747 ( .C1(n22131), .C2(n22270), .A(n22126), .B(n22125), .ZN(
        P1_U3110) );
  OAI22_X1 U23748 ( .A1(n22273), .A2(n22143), .B1(n22127), .B2(n22271), .ZN(
        n22128) );
  INV_X1 U23749 ( .A(n22128), .ZN(n22130) );
  AOI22_X1 U23750 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n22276), .B1(
        n22138), .B2(n22275), .ZN(n22129) );
  OAI211_X1 U23751 ( .C1(n22131), .C2(n22279), .A(n22130), .B(n22129), .ZN(
        P1_U3118) );
  AOI22_X1 U23752 ( .A1(n22291), .A2(n22132), .B1(n22139), .B2(n22281), .ZN(
        n22134) );
  AOI22_X1 U23753 ( .A1(n22284), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n22140), .B2(n22283), .ZN(n22133) );
  OAI211_X1 U23754 ( .C1(n22288), .C2(n22135), .A(n22134), .B(n22133), .ZN(
        P1_U3134) );
  AOI22_X1 U23755 ( .A1(n22139), .A2(n22289), .B1(n22138), .B2(n22290), .ZN(
        n22137) );
  AOI22_X1 U23756 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n22292), .B1(
        n22291), .B2(n22140), .ZN(n22136) );
  OAI211_X1 U23757 ( .C1(n22143), .C2(n22295), .A(n22137), .B(n22136), .ZN(
        P1_U3142) );
  AOI22_X1 U23758 ( .A1(n22139), .A2(n22296), .B1(n22138), .B2(n22298), .ZN(
        n22142) );
  AOI22_X1 U23759 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n22302), .B1(
        n22301), .B2(n22140), .ZN(n22141) );
  OAI211_X1 U23760 ( .C1(n22143), .C2(n22305), .A(n22142), .B(n22141), .ZN(
        P1_U3150) );
  NAND2_X1 U23761 ( .A1(n22149), .A2(n22148), .ZN(n22179) );
  AOI22_X1 U23762 ( .A1(n22207), .A2(n22193), .B1(n22198), .B2(n22206), .ZN(
        n22155) );
  INV_X1 U23763 ( .A(DATAI_22_), .ZN(n22151) );
  OAI22_X1 U23764 ( .A1(n22153), .A2(n22152), .B1(n22151), .B2(n22150), .ZN(
        n22201) );
  AOI22_X1 U23765 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n22208), .B1(
        n22214), .B2(n22201), .ZN(n22154) );
  OAI211_X1 U23766 ( .C1(n22211), .C2(n22190), .A(n22155), .B(n22154), .ZN(
        P1_U3039) );
  INV_X1 U23767 ( .A(n22201), .ZN(n22196) );
  AOI22_X1 U23768 ( .A1(n22200), .A2(n22213), .B1(n22198), .B2(n22212), .ZN(
        n22157) );
  AOI22_X1 U23769 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n22215), .B1(
        n22214), .B2(n22193), .ZN(n22156) );
  OAI211_X1 U23770 ( .C1(n22196), .C2(n22219), .A(n22157), .B(n22156), .ZN(
        P1_U3047) );
  AOI22_X1 U23771 ( .A1(n22226), .A2(n22201), .B1(n22158), .B2(n22198), .ZN(
        n22161) );
  AOI22_X1 U23772 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n22221), .B1(
        n22159), .B2(n22193), .ZN(n22160) );
  OAI211_X1 U23773 ( .C1(n22224), .C2(n22190), .A(n22161), .B(n22160), .ZN(
        P1_U3055) );
  AOI22_X1 U23774 ( .A1(n22226), .A2(n22193), .B1(n22225), .B2(n22198), .ZN(
        n22163) );
  AOI22_X1 U23775 ( .A1(n22227), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n22233), .B2(n22201), .ZN(n22162) );
  OAI211_X1 U23776 ( .C1(n22230), .C2(n22190), .A(n22163), .B(n22162), .ZN(
        P1_U3063) );
  AOI22_X1 U23777 ( .A1(n22200), .A2(n22232), .B1(n22198), .B2(n22231), .ZN(
        n22165) );
  AOI22_X1 U23778 ( .A1(n22234), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n22233), .B2(n22193), .ZN(n22164) );
  OAI211_X1 U23779 ( .C1(n22196), .C2(n22243), .A(n22165), .B(n22164), .ZN(
        P1_U3071) );
  AOI22_X1 U23780 ( .A1(n22200), .A2(n22238), .B1(n22198), .B2(n22237), .ZN(
        n22168) );
  AOI22_X1 U23781 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n22240), .B1(
        n22166), .B2(n22193), .ZN(n22167) );
  OAI211_X1 U23782 ( .C1(n22196), .C2(n22245), .A(n22168), .B(n22167), .ZN(
        P1_U3079) );
  INV_X1 U23783 ( .A(n22193), .ZN(n22205) );
  OAI22_X1 U23784 ( .A1(n22245), .A2(n22205), .B1(n22179), .B2(n22244), .ZN(
        n22169) );
  INV_X1 U23785 ( .A(n22169), .ZN(n22171) );
  AOI22_X1 U23786 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n22247), .B1(
        n22253), .B2(n22201), .ZN(n22170) );
  OAI211_X1 U23787 ( .C1(n22250), .C2(n22190), .A(n22171), .B(n22170), .ZN(
        P1_U3087) );
  AOI22_X1 U23788 ( .A1(n22200), .A2(n22252), .B1(n22198), .B2(n22251), .ZN(
        n22173) );
  AOI22_X1 U23789 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n22254), .B1(
        n22253), .B2(n22193), .ZN(n22172) );
  OAI211_X1 U23790 ( .C1(n22196), .C2(n22257), .A(n22173), .B(n22172), .ZN(
        P1_U3095) );
  AOI22_X1 U23791 ( .A1(n11071), .A2(n22200), .B1(n22198), .B2(n22258), .ZN(
        n22175) );
  AOI22_X1 U23792 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n22261), .B1(
        n22260), .B2(n22193), .ZN(n22174) );
  OAI211_X1 U23793 ( .C1(n22196), .C2(n22270), .A(n22175), .B(n22174), .ZN(
        P1_U3103) );
  AOI22_X1 U23794 ( .A1(n22200), .A2(n22265), .B1(n22198), .B2(n22264), .ZN(
        n22178) );
  AOI22_X1 U23795 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n22267), .B1(
        n22176), .B2(n22193), .ZN(n22177) );
  OAI211_X1 U23796 ( .C1(n22196), .C2(n22279), .A(n22178), .B(n22177), .ZN(
        P1_U3111) );
  OAI22_X1 U23797 ( .A1(n22273), .A2(n22196), .B1(n22179), .B2(n22271), .ZN(
        n22180) );
  INV_X1 U23798 ( .A(n22180), .ZN(n22182) );
  AOI22_X1 U23799 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n22276), .B1(
        n22200), .B2(n22275), .ZN(n22181) );
  OAI211_X1 U23800 ( .C1(n22205), .C2(n22279), .A(n22182), .B(n22181), .ZN(
        P1_U3119) );
  AOI22_X1 U23801 ( .A1(n22200), .A2(n22184), .B1(n22198), .B2(n22183), .ZN(
        n22187) );
  AOI22_X1 U23802 ( .A1(n22185), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n22283), .B2(n22201), .ZN(n22186) );
  OAI211_X1 U23803 ( .C1(n22205), .C2(n22273), .A(n22187), .B(n22186), .ZN(
        P1_U3127) );
  AOI22_X1 U23804 ( .A1(n22291), .A2(n22201), .B1(n22198), .B2(n22281), .ZN(
        n22189) );
  AOI22_X1 U23805 ( .A1(n22284), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n22193), .B2(n22283), .ZN(n22188) );
  OAI211_X1 U23806 ( .C1(n22288), .C2(n22190), .A(n22189), .B(n22188), .ZN(
        P1_U3135) );
  AOI22_X1 U23807 ( .A1(n22200), .A2(n22290), .B1(n22198), .B2(n22289), .ZN(
        n22192) );
  AOI22_X1 U23808 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n22292), .B1(
        n22291), .B2(n22193), .ZN(n22191) );
  OAI211_X1 U23809 ( .C1(n22196), .C2(n22295), .A(n22192), .B(n22191), .ZN(
        P1_U3143) );
  AOI22_X1 U23810 ( .A1(n22200), .A2(n22298), .B1(n22198), .B2(n22296), .ZN(
        n22195) );
  AOI22_X1 U23811 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n22302), .B1(
        n22301), .B2(n22193), .ZN(n22194) );
  OAI211_X1 U23812 ( .C1(n22196), .C2(n22305), .A(n22195), .B(n22194), .ZN(
        P1_U3151) );
  AOI22_X1 U23813 ( .A1(n22200), .A2(n22199), .B1(n22198), .B2(n22197), .ZN(
        n22204) );
  AOI22_X1 U23814 ( .A1(n22202), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n22201), .B2(n22207), .ZN(n22203) );
  OAI211_X1 U23815 ( .C1(n22205), .C2(n22305), .A(n22204), .B(n22203), .ZN(
        P1_U3159) );
  AOI22_X1 U23816 ( .A1(n22207), .A2(n22300), .B1(n22297), .B2(n22206), .ZN(
        n22210) );
  AOI22_X1 U23817 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n22208), .B1(
        n22214), .B2(n22282), .ZN(n22209) );
  OAI211_X1 U23818 ( .C1(n22211), .C2(n22287), .A(n22210), .B(n22209), .ZN(
        P1_U3040) );
  AOI22_X1 U23819 ( .A1(n22299), .A2(n22213), .B1(n22297), .B2(n22212), .ZN(
        n22217) );
  AOI22_X1 U23820 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n22215), .B1(
        n22214), .B2(n22300), .ZN(n22216) );
  OAI211_X1 U23821 ( .C1(n22306), .C2(n22219), .A(n22217), .B(n22216), .ZN(
        P1_U3048) );
  OAI22_X1 U23822 ( .A1(n22219), .A2(n22280), .B1(n22272), .B2(n22218), .ZN(
        n22220) );
  INV_X1 U23823 ( .A(n22220), .ZN(n22223) );
  AOI22_X1 U23824 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n22221), .B1(
        n22226), .B2(n22282), .ZN(n22222) );
  OAI211_X1 U23825 ( .C1(n22224), .C2(n22287), .A(n22223), .B(n22222), .ZN(
        P1_U3056) );
  AOI22_X1 U23826 ( .A1(n22233), .A2(n22282), .B1(n22297), .B2(n22225), .ZN(
        n22229) );
  AOI22_X1 U23827 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n22227), .B1(
        n22226), .B2(n22300), .ZN(n22228) );
  OAI211_X1 U23828 ( .C1(n22230), .C2(n22287), .A(n22229), .B(n22228), .ZN(
        P1_U3064) );
  AOI22_X1 U23829 ( .A1(n22299), .A2(n22232), .B1(n22297), .B2(n22231), .ZN(
        n22236) );
  AOI22_X1 U23830 ( .A1(n22234), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n22233), .B2(n22300), .ZN(n22235) );
  OAI211_X1 U23831 ( .C1(n22306), .C2(n22243), .A(n22236), .B(n22235), .ZN(
        P1_U3072) );
  AOI22_X1 U23832 ( .A1(n22299), .A2(n22238), .B1(n22297), .B2(n22237), .ZN(
        n22242) );
  AOI22_X1 U23833 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n22240), .B1(
        n22239), .B2(n22282), .ZN(n22241) );
  OAI211_X1 U23834 ( .C1(n22280), .C2(n22243), .A(n22242), .B(n22241), .ZN(
        P1_U3080) );
  OAI22_X1 U23835 ( .A1(n22245), .A2(n22280), .B1(n22272), .B2(n22244), .ZN(
        n22246) );
  INV_X1 U23836 ( .A(n22246), .ZN(n22249) );
  AOI22_X1 U23837 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n22247), .B1(
        n22253), .B2(n22282), .ZN(n22248) );
  OAI211_X1 U23838 ( .C1(n22250), .C2(n22287), .A(n22249), .B(n22248), .ZN(
        P1_U3088) );
  AOI22_X1 U23839 ( .A1(n22299), .A2(n22252), .B1(n22251), .B2(n22297), .ZN(
        n22256) );
  AOI22_X1 U23840 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n22254), .B1(
        n22253), .B2(n22300), .ZN(n22255) );
  OAI211_X1 U23841 ( .C1(n22306), .C2(n22257), .A(n22256), .B(n22255), .ZN(
        P1_U3096) );
  AOI22_X1 U23842 ( .A1(n11071), .A2(n22299), .B1(n22297), .B2(n22258), .ZN(
        n22263) );
  AOI22_X1 U23843 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n22261), .B1(
        n22260), .B2(n22300), .ZN(n22262) );
  OAI211_X1 U23844 ( .C1(n22306), .C2(n22270), .A(n22263), .B(n22262), .ZN(
        P1_U3104) );
  AOI22_X1 U23845 ( .A1(n22299), .A2(n22265), .B1(n22297), .B2(n22264), .ZN(
        n22269) );
  AOI22_X1 U23846 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n22267), .B1(
        n22266), .B2(n22282), .ZN(n22268) );
  OAI211_X1 U23847 ( .C1(n22280), .C2(n22270), .A(n22269), .B(n22268), .ZN(
        P1_U3112) );
  OAI22_X1 U23848 ( .A1(n22273), .A2(n22306), .B1(n22272), .B2(n22271), .ZN(
        n22274) );
  INV_X1 U23849 ( .A(n22274), .ZN(n22278) );
  AOI22_X1 U23850 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n22276), .B1(
        n22299), .B2(n22275), .ZN(n22277) );
  OAI211_X1 U23851 ( .C1(n22280), .C2(n22279), .A(n22278), .B(n22277), .ZN(
        P1_U3120) );
  AOI22_X1 U23852 ( .A1(n22291), .A2(n22282), .B1(n22297), .B2(n22281), .ZN(
        n22286) );
  AOI22_X1 U23853 ( .A1(n22284), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n22300), .B2(n22283), .ZN(n22285) );
  OAI211_X1 U23854 ( .C1(n22288), .C2(n22287), .A(n22286), .B(n22285), .ZN(
        P1_U3136) );
  AOI22_X1 U23855 ( .A1(n22299), .A2(n22290), .B1(n22297), .B2(n22289), .ZN(
        n22294) );
  AOI22_X1 U23856 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n22292), .B1(
        n22291), .B2(n22300), .ZN(n22293) );
  OAI211_X1 U23857 ( .C1(n22306), .C2(n22295), .A(n22294), .B(n22293), .ZN(
        P1_U3144) );
  AOI22_X1 U23858 ( .A1(n22299), .A2(n22298), .B1(n22297), .B2(n22296), .ZN(
        n22304) );
  AOI22_X1 U23859 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n22302), .B1(
        n22301), .B2(n22300), .ZN(n22303) );
  OAI211_X1 U23860 ( .C1(n22306), .C2(n22305), .A(n22304), .B(n22303), .ZN(
        P1_U3152) );
  OAI22_X1 U23861 ( .A1(n22308), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n22307), .ZN(n22309) );
  INV_X1 U23862 ( .A(n22309), .ZN(P1_U3486) );
  OAI21_X1 U23863 ( .B1(n22311), .B2(n22310), .A(P1_MEMORYFETCH_REG_SCAN_IN), 
        .ZN(n22313) );
  NAND2_X1 U23864 ( .A1(n22313), .A2(n22312), .ZN(P1_U2801) );
  INV_X1 U12886 ( .A(n14367), .ZN(n14360) );
  INV_X2 U11099 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11613) );
  AND2_X2 U14056 ( .A1(n12518), .A2(n14900), .ZN(n12735) );
  AND2_X2 U11390 ( .A1(n14749), .A2(n11215), .ZN(n12736) );
  NAND2_X1 U12544 ( .A1(n12639), .A2(n15596), .ZN(n12618) );
  CLKBUF_X1 U11084 ( .A(n12696), .Z(n12728) );
  INV_X2 U11197 ( .A(n17655), .ZN(n17703) );
  XNOR2_X1 U15424 ( .A(n13680), .B(n13679), .ZN(n14842) );
  AND2_X1 U12480 ( .A1(n15787), .A2(n11049), .ZN(n15740) );
  CLKBUF_X1 U11112 ( .A(n12761), .Z(n12672) );
  AND2_X2 U11131 ( .A1(n11215), .A2(n14895), .ZN(n12696) );
  CLKBUF_X1 U11138 ( .A(n12385), .Z(n14233) );
  CLKBUF_X1 U11139 ( .A(n11643), .Z(n10971) );
  NOR2_X2 U11170 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15321) );
  INV_X2 U11179 ( .A(n14446), .ZN(n14411) );
  CLKBUF_X1 U11184 ( .A(n11721), .Z(n11722) );
  CLKBUF_X1 U11185 ( .A(n13534), .Z(n10976) );
  CLKBUF_X1 U11186 ( .A(n12513), .Z(n14731) );
  CLKBUF_X1 U11360 ( .A(n12621), .Z(n15245) );
  CLKBUF_X1 U11845 ( .A(n14819), .Z(n10980) );
  CLKBUF_X1 U11869 ( .A(n11681), .Z(n12246) );
  CLKBUF_X1 U12076 ( .A(n15740), .Z(n15741) );
  CLKBUF_X1 U12167 ( .A(n17307), .Z(n17320) );
  CLKBUF_X1 U13178 ( .A(n20140), .Z(n20142) );
  CLKBUF_X1 U14052 ( .A(n18111), .Z(n10977) );
  INV_X2 U14202 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15576) );
  CLKBUF_X1 U14205 ( .A(n11749), .Z(n18258) );
  CLKBUF_X1 U17863 ( .A(n12736), .Z(n12671) );
endmodule

