

module b17_C_2inp_gates_syn ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, 
        DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, 
        DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, 
        DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, 
        DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, 
        DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, 
        READY1, READY2, P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN, 
        P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN, 
        P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN, 
        P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN, 
        P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN, 
        P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN, 
        P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN, 
        P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN, 
        P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN, 
        P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN, 
        P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN, 
        P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN, 
        P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN, 
        P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN, 
        P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN, 
        P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN, 
        P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN, 
        P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, 
        P1_REIP_REG_6__SCAN_IN, P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, 
        P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, 
        P1_REIP_REG_0__SCAN_IN, P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, 
        P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, 
        P1_EBX_REG_26__SCAN_IN, P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, 
        P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, 
        P1_EBX_REG_20__SCAN_IN, P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, 
        P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, 
        P1_EBX_REG_14__SCAN_IN, P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, 
        P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, 
        P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, 
        P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, 
        P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, 
        P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, 
        P1_EAX_REG_28__SCAN_IN, P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, 
        P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, 
        P1_EAX_REG_22__SCAN_IN, P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, 
        P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, 
        P1_EAX_REG_16__SCAN_IN, P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, 
        P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, 
        P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, 
        P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, 
        P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, 
        P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput127, keyinput126, keyinput125,
         keyinput124, keyinput123, keyinput122, keyinput121, keyinput120,
         keyinput119, keyinput118, keyinput117, keyinput116, keyinput115,
         keyinput114, keyinput113, keyinput112, keyinput111, keyinput110,
         keyinput109, keyinput108, keyinput107, keyinput106, keyinput105,
         keyinput104, keyinput103, keyinput102, keyinput101, keyinput100,
         keyinput99, keyinput98, keyinput97, keyinput96, keyinput95,
         keyinput94, keyinput93, keyinput92, keyinput91, keyinput90,
         keyinput89, keyinput88, keyinput87, keyinput86, keyinput85,
         keyinput84, keyinput83, keyinput82, keyinput81, keyinput80,
         keyinput79, keyinput78, keyinput77, keyinput76, keyinput75,
         keyinput74, keyinput73, keyinput72, keyinput71, keyinput70,
         keyinput69, keyinput68, keyinput67, keyinput66, keyinput65,
         keyinput64, keyinput63, keyinput62, keyinput61, keyinput60,
         keyinput59, keyinput58, keyinput57, keyinput56, keyinput55,
         keyinput54, keyinput53, keyinput52, keyinput51, keyinput50,
         keyinput49, keyinput48, keyinput47, keyinput46, keyinput45,
         keyinput44, keyinput43, keyinput42, keyinput41, keyinput40,
         keyinput39, keyinput38, keyinput37, keyinput36, keyinput35,
         keyinput34, keyinput33, keyinput32, keyinput31, keyinput30,
         keyinput29, keyinput28, keyinput27, keyinput26, keyinput25,
         keyinput24, keyinput23, keyinput22, keyinput21, keyinput20,
         keyinput19, keyinput18, keyinput17, keyinput16, keyinput15,
         keyinput14, keyinput13, keyinput12, keyinput11, keyinput10, keyinput9,
         keyinput8, keyinput7, keyinput6, keyinput5, keyinput4, keyinput3,
         keyinput2, keyinput1, keyinput0;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9725, n9726, n9727,
         n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737,
         n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747,
         n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757,
         n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767,
         n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777,
         n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787,
         n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797,
         n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807,
         n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817,
         n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857,
         n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867,
         n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877,
         n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887,
         n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897,
         n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907,
         n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
         n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
         n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
         n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
         n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
         n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
         n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
         n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
         n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
         n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
         n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014,
         n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022,
         n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
         n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038,
         n10039, n10040, n10041, n10042, n10043, n10044, n10045, n10046,
         n10047, n10048, n10049, n10050, n10051, n10052, n10053, n10054,
         n10055, n10056, n10057, n10058, n10059, n10060, n10061, n10062,
         n10063, n10064, n10065, n10066, n10067, n10068, n10069, n10070,
         n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
         n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086,
         n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
         n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102,
         n10103, n10104, n10105, n10106, n10107, n10108, n10109, n10110,
         n10111, n10112, n10113, n10114, n10115, n10116, n10117, n10118,
         n10119, n10120, n10121, n10122, n10123, n10124, n10125, n10126,
         n10127, n10128, n10129, n10130, n10131, n10132, n10133, n10134,
         n10135, n10136, n10137, n10138, n10139, n10140, n10141, n10142,
         n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
         n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
         n10167, n10168, n10169, n10170, n10171, n10172, n10173, n10174,
         n10175, n10176, n10177, n10178, n10179, n10180, n10181, n10182,
         n10183, n10184, n10185, n10186, n10187, n10188, n10189, n10190,
         n10191, n10192, n10193, n10194, n10195, n10196, n10197, n10198,
         n10199, n10200, n10201, n10202, n10203, n10204, n10205, n10206,
         n10207, n10208, n10209, n10210, n10211, n10212, n10213, n10214,
         n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
         n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238,
         n10239, n10240, n10241, n10242, n10243, n10244, n10245, n10246,
         n10247, n10248, n10249, n10250, n10251, n10252, n10253, n10254,
         n10255, n10256, n10257, n10258, n10259, n10260, n10261, n10262,
         n10263, n10264, n10265, n10266, n10267, n10268, n10269, n10270,
         n10271, n10272, n10273, n10274, n10275, n10276, n10277, n10278,
         n10279, n10280, n10281, n10282, n10283, n10284, n10285, n10286,
         n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
         n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302,
         n10303, n10304, n10305, n10306, n10307, n10308, n10309, n10310,
         n10311, n10312, n10313, n10314, n10315, n10316, n10317, n10318,
         n10319, n10320, n10321, n10322, n10323, n10324, n10325, n10326,
         n10327, n10328, n10329, n10330, n10331, n10332, n10333, n10334,
         n10335, n10336, n10337, n10338, n10339, n10340, n10341, n10342,
         n10343, n10344, n10345, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10355, n10356, n10357, n10358,
         n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
         n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374,
         n10375, n10376, n10377, n10378, n10379, n10380, n10381, n10382,
         n10383, n10384, n10385, n10386, n10387, n10388, n10389, n10390,
         n10391, n10392, n10393, n10394, n10395, n10396, n10397, n10398,
         n10399, n10400, n10401, n10402, n10403, n10404, n10405, n10406,
         n10407, n10408, n10409, n10410, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
         n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438,
         n10439, n10440, n10441, n10442, n10443, n10444, n10445, n10446,
         n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710,
         n10711, n10712, n10713, n10714, n10715, n10716, n10717, n10718,
         n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726,
         n10727, n10728, n10729, n10730, n10731, n10732, n10733, n10734,
         n10735, n10736, n10737, n10738, n10739, n10740, n10741, n10742,
         n10743, n10744, n10745, n10746, n10747, n10748, n10749, n10750,
         n10751, n10752, n10753, n10754, n10755, n10756, n10757, n10758,
         n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
         n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774,
         n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
         n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790,
         n10791, n10792, n10793, n10794, n10795, n10796, n10797, n10798,
         n10799, n10800, n10801, n10802, n10803, n10804, n10805, n10806,
         n10807, n10808, n10809, n10810, n10811, n10812, n10813, n10814,
         n10815, n10816, n10817, n10818, n10819, n10820, n10821, n10822,
         n10823, n10824, n10825, n10826, n10827, n10828, n10829, n10830,
         n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
         n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
         n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862,
         n10863, n10864, n10865, n10866, n10867, n10868, n10869, n10870,
         n10871, n10872, n10873, n10874, n10875, n10876, n10877, n10878,
         n10879, n10880, n10881, n10882, n10883, n10884, n10885, n10886,
         n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
         n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902,
         n10903, n10904, n10905, n10906, n10907, n10908, n10909, n10910,
         n10911, n10912, n10913, n10914, n10915, n10916, n10917, n10918,
         n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
         n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934,
         n10935, n10936, n10937, n10938, n10939, n10940, n10941, n10942,
         n10943, n10944, n10945, n10946, n10947, n10948, n10949, n10950,
         n10951, n10952, n10953, n10954, n10955, n10956, n10957, n10958,
         n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
         n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974,
         n10975, n10976, n10977, n10978, n10979, n10980, n10981, n10982,
         n10983, n10984, n10985, n10986, n10987, n10988, n10989, n10990,
         n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
         n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
         n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030,
         n11031, n11032, n11033, n11034, n11035, n11036, n11037, n11038,
         n11039, n11040, n11041, n11042, n11043, n11044, n11045, n11046,
         n11047, n11048, n11049, n11050, n11051, n11052, n11053, n11054,
         n11055, n11056, n11057, n11058, n11059, n11060, n11061, n11062,
         n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078,
         n11079, n11080, n11081, n11082, n11083, n11084, n11085, n11086,
         n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
         n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102,
         n11103, n11104, n11105, n11106, n11107, n11108, n11109, n11110,
         n11111, n11112, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11121, n11122, n11123, n11124, n11125, n11126,
         n11127, n11128, n11129, n11130, n11131, n11132, n11133, n11134,
         n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
         n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150,
         n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
         n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166,
         n11167, n11168, n11169, n11170, n11171, n11172, n11173, n11174,
         n11175, n11176, n11177, n11178, n11179, n11180, n11181, n11182,
         n11183, n11184, n11185, n11186, n11187, n11188, n11189, n11190,
         n11191, n11192, n11193, n11194, n11195, n11196, n11197, n11198,
         n11199, n11200, n11201, n11202, n11203, n11204, n11205, n11206,
         n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
         n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222,
         n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11230,
         n11231, n11232, n11233, n11234, n11235, n11236, n11237, n11238,
         n11239, n11240, n11241, n11242, n11243, n11244, n11245, n11246,
         n11247, n11248, n11249, n11250, n11251, n11252, n11253, n11254,
         n11255, n11256, n11257, n11258, n11259, n11260, n11261, n11262,
         n11263, n11264, n11265, n11266, n11267, n11268, n11269, n11270,
         n11271, n11272, n11273, n11274, n11275, n11276, n11277, n11278,
         n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
         n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
         n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302,
         n11303, n11304, n11305, n11306, n11307, n11308, n11309, n11310,
         n11311, n11312, n11313, n11314, n11315, n11316, n11317, n11318,
         n11319, n11320, n11321, n11322, n11323, n11324, n11325, n11326,
         n11327, n11328, n11329, n11330, n11331, n11332, n11333, n11334,
         n11335, n11336, n11337, n11338, n11339, n11340, n11341, n11342,
         n11343, n11344, n11345, n11346, n11347, n11348, n11349, n11350,
         n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
         n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366,
         n11367, n11368, n11369, n11370, n11371, n11372, n11373, n11374,
         n11375, n11376, n11377, n11378, n11379, n11380, n11381, n11382,
         n11383, n11384, n11385, n11386, n11387, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11397, n11398,
         n11399, n11400, n11401, n11402, n11403, n11404, n11405, n11406,
         n11407, n11408, n11409, n11410, n11411, n11412, n11413, n11414,
         n11415, n11416, n11417, n11418, n11419, n11420, n11421, n11422,
         n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
         n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438,
         n11439, n11440, n11441, n11442, n11443, n11444, n11445, n11446,
         n11447, n11448, n11449, n11450, n11451, n11452, n11453, n11454,
         n11455, n11456, n11457, n11458, n11459, n11460, n11461, n11462,
         n11463, n11464, n11465, n11466, n11467, n11468, n11469, n11470,
         n11471, n11472, n11473, n11474, n11475, n11476, n11477, n11478,
         n11479, n11480, n11481, n11482, n11483, n11484, n11485, n11486,
         n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
         n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
         n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510,
         n11511, n11512, n11513, n11514, n11515, n11516, n11517, n11518,
         n11519, n11520, n11521, n11522, n11523, n11524, n11525, n11526,
         n11527, n11528, n11529, n11530, n11531, n11532, n11533, n11534,
         n11535, n11536, n11537, n11538, n11539, n11540, n11541, n11542,
         n11543, n11544, n11545, n11546, n11547, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11555, n11556, n11557, n11558,
         n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
         n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
         n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582,
         n11583, n11584, n11585, n11586, n11587, n11588, n11589, n11590,
         n11591, n11592, n11593, n11594, n11595, n11596, n11597, n11598,
         n11599, n11600, n11601, n11602, n11603, n11604, n11605, n11606,
         n11607, n11608, n11609, n11610, n11611, n11612, n11613, n11614,
         n11615, n11616, n11617, n11618, n11619, n11620, n11621, n11622,
         n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
         n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638,
         n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
         n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654,
         n11655, n11656, n11657, n11658, n11659, n11660, n11661, n11662,
         n11663, n11664, n11665, n11666, n11667, n11668, n11669, n11670,
         n11671, n11672, n11673, n11674, n11675, n11676, n11677, n11678,
         n11679, n11680, n11681, n11682, n11683, n11684, n11685, n11686,
         n11687, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
         n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702,
         n11703, n11704, n11705, n11706, n11707, n11708, n11709, n11710,
         n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
         n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726,
         n11727, n11728, n11729, n11730, n11731, n11732, n11733, n11734,
         n11735, n11736, n11737, n11738, n11739, n11740, n11741, n11742,
         n11743, n11744, n11745, n11746, n11747, n11748, n11749, n11750,
         n11751, n11752, n11753, n11754, n11755, n11756, n11757, n11758,
         n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
         n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774,
         n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
         n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790,
         n11791, n11792, n11793, n11794, n11795, n11796, n11797, n11798,
         n11799, n11800, n11801, n11802, n11803, n11804, n11805, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11813, n11814,
         n11815, n11816, n11817, n11818, n11819, n11820, n11821, n11822,
         n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
         n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838,
         n11839, n11840, n11841, n11842, n11843, n11844, n11845, n11846,
         n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
         n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862,
         n11863, n11864, n11865, n11866, n11867, n11868, n11869, n11870,
         n11871, n11872, n11873, n11874, n11875, n11876, n11877, n11878,
         n11879, n11880, n11881, n11882, n11883, n11884, n11885, n11886,
         n11887, n11888, n11889, n11890, n11891, n11892, n11893, n11894,
         n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
         n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
         n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,
         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
         n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650,
         n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,
         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
         n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
         n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
         n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
         n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
         n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722,
         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
         n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,
         n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
         n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
         n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
         n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834,
         n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
         n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
         n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
         n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866,
         n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
         n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882,
         n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890,
         n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
         n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906,
         n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914,
         n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922,
         n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
         n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938,
         n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946,
         n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954,
         n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962,
         n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970,
         n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978,
         n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986,
         n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994,
         n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002,
         n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010,
         n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018,
         n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026,
         n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034,
         n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042,
         n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050,
         n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058,
         n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066,
         n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074,
         n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082,
         n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
         n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098,
         n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
         n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114,
         n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122,
         n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130,
         n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
         n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146,
         n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154,
         n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
         n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
         n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178,
         n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186,
         n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194,
         n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202,
         n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
         n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218,
         n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226,
         n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
         n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
         n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250,
         n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258,
         n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266,
         n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274,
         n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282,
         n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290,
         n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298,
         n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
         n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314,
         n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322,
         n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330,
         n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338,
         n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346,
         n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354,
         n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362,
         n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370,
         n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
         n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386,
         n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394,
         n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402,
         n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410,
         n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418,
         n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
         n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434,
         n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442,
         n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
         n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458,
         n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466,
         n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474,
         n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
         n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490,
         n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
         n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506,
         n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
         n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522,
         n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530,
         n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538,
         n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546,
         n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554,
         n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562,
         n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570,
         n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578,
         n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586,
         n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
         n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602,
         n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610,
         n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618,
         n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
         n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
         n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642,
         n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650,
         n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658,
         n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666,
         n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674,
         n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682,
         n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690,
         n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698,
         n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
         n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
         n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722,
         n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730,
         n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
         n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746,
         n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754,
         n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762,
         n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770,
         n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
         n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
         n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794,
         n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802,
         n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
         n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818,
         n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
         n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834,
         n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
         n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
         n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
         n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906,
         n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914,
         n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
         n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
         n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938,
         n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
         n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954,
         n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962,
         n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970,
         n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978,
         n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986,
         n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
         n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
         n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
         n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018,
         n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
         n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034,
         n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
         n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
         n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
         n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
         n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
         n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
         n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
         n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
         n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
         n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
         n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
         n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162,
         n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
         n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178,
         n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
         n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
         n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202,
         n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
         n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
         n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226,
         n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250,
         n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
         n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
         n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274,
         n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282,
         n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
         n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298,
         n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306,
         n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314,
         n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322,
         n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
         n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338,
         n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
         n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
         n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
         n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370,
         n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378,
         n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
         n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
         n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
         n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
         n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
         n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
         n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
         n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442,
         n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450,
         n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
         n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
         n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
         n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482,
         n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490,
         n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
         n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
         n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514,
         n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
         n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
         n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
         n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
         n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554,
         n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562,
         n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
         n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
         n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
         n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610,
         n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
         n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626,
         n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634,
         n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
         n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
         n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
         n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
         n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
         n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
         n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
         n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
         n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
         n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754,
         n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
         n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770,
         n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778,
         n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
         n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
         n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
         n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
         n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
         n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
         n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842,
         n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
         n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
         n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
         n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874,
         n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
         n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
         n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
         n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
         n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946,
         n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
         n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
         n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970,
         n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
         n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986,
         n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994,
         n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
         n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
         n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018,
         n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026,
         n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034,
         n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
         n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050,
         n21051;

  INV_X1 U11161 ( .A(n19993), .ZN(n19965) );
  NOR2_X1 U11163 ( .A1(n12728), .A2(n15277), .ZN(n15032) );
  NOR2_X1 U11164 ( .A1(n19815), .A2(n19357), .ZN(n19448) );
  AND2_X1 U11165 ( .A1(n13969), .A2(n13968), .ZN(n15233) );
  OR2_X1 U11166 ( .A1(n16052), .A2(n13845), .ZN(n13866) );
  INV_X2 U11167 ( .A(n16758), .ZN(n16820) );
  CLKBUF_X1 U11168 ( .A(n9763), .Z(n9719) );
  AND2_X2 U11169 ( .A1(n11932), .A2(n19385), .ZN(n10267) );
  OR2_X1 U11170 ( .A1(n11929), .A2(n11928), .ZN(n19601) );
  NAND2_X1 U11171 ( .A1(n11296), .A2(n11295), .ZN(n20097) );
  AND2_X1 U11172 ( .A1(n11922), .A2(n11921), .ZN(n12007) );
  AND2_X1 U11173 ( .A1(n11920), .A2(n11926), .ZN(n12030) );
  AND2_X1 U11174 ( .A1(n11920), .A2(n11921), .ZN(n19433) );
  AND2_X1 U11175 ( .A1(n11922), .A2(n11926), .ZN(n19262) );
  AND2_X1 U11176 ( .A1(n11911), .A2(n11917), .ZN(n12009) );
  CLKBUF_X2 U11177 ( .A(n11916), .Z(n15591) );
  CLKBUF_X2 U11178 ( .A(n16992), .Z(n17118) );
  BUF_X2 U11179 ( .A(n12836), .Z(n17192) );
  CLKBUF_X2 U11180 ( .A(n12994), .Z(n17097) );
  CLKBUF_X1 U11181 ( .A(n12994), .Z(n17191) );
  CLKBUF_X1 U11182 ( .A(n16992), .Z(n17057) );
  AND3_X1 U11183 ( .A1(n13394), .A2(n11173), .A3(n11172), .ZN(n10055) );
  AND2_X1 U11184 ( .A1(n10662), .A2(n10809), .ZN(n12518) );
  AND2_X1 U11185 ( .A1(n12542), .A2(n10239), .ZN(n12524) );
  CLKBUF_X2 U11186 ( .A(n11136), .Z(n11636) );
  AND2_X1 U11187 ( .A1(n10661), .A2(n10809), .ZN(n12517) );
  CLKBUF_X2 U11188 ( .A(n11090), .Z(n9721) );
  INV_X1 U11189 ( .A(n10368), .ZN(n12528) );
  NAND2_X2 U11190 ( .A1(n18827), .A2(n21023), .ZN(n16826) );
  BUF_X1 U11191 ( .A(n11114), .Z(n13196) );
  CLKBUF_X2 U11192 ( .A(n11156), .Z(n13568) );
  NAND2_X1 U11193 ( .A1(n10752), .A2(n10690), .ZN(n12221) );
  CLKBUF_X1 U11194 ( .A(n11165), .Z(n11782) );
  INV_X1 U11195 ( .A(n11730), .ZN(n20139) );
  CLKBUF_X3 U11196 ( .A(n10741), .Z(n19237) );
  NAND2_X1 U11197 ( .A1(n19228), .A2(n10735), .ZN(n10758) );
  INV_X1 U11199 ( .A(n10725), .ZN(n10742) );
  AND2_X1 U11200 ( .A1(n10926), .A2(n10929), .ZN(n9752) );
  AND2_X2 U11201 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10929) );
  NOR2_X2 U11202 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13468) );
  AND2_X2 U11203 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10930) );
  AND2_X2 U11204 ( .A1(n10238), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9744) );
  AND3_X1 U11205 ( .A1(n10198), .A2(n9737), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9746) );
  AND2_X2 U11206 ( .A1(n15580), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10662) );
  INV_X1 U11207 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10198) );
  AND2_X2 U11208 ( .A1(n9906), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15579) );
  CLKBUF_X1 U11209 ( .A(n18112), .Z(n9717) );
  NOR3_X1 U11210 ( .A1(n16337), .A2(n18679), .A3(n18185), .ZN(n18112) );
  AND2_X2 U11211 ( .A1(n9728), .A2(n9729), .ZN(n14156) );
  NOR2_X2 U11212 ( .A1(n10759), .A2(n10758), .ZN(n12703) );
  AND2_X1 U11213 ( .A1(n13468), .A2(n10928), .ZN(n11107) );
  CLKBUF_X2 U11214 ( .A(n11107), .Z(n11616) );
  AND3_X1 U11215 ( .A1(n10198), .A2(n10197), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9761) );
  AND4_X1 U11216 ( .A1(n11144), .A2(n11143), .A3(n11142), .A4(n11141), .ZN(
        n11155) );
  NAND2_X1 U11217 ( .A1(n11222), .A2(n11730), .ZN(n11733) );
  BUF_X1 U11218 ( .A(n12540), .Z(n12686) );
  OAI21_X1 U11219 ( .B1(n9763), .B2(n15558), .A(n10781), .ZN(n10783) );
  OR2_X1 U11220 ( .A1(n11929), .A2(n11906), .ZN(n11960) );
  NAND2_X1 U11221 ( .A1(n18827), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12789) );
  NAND2_X1 U11222 ( .A1(n18812), .A2(n18820), .ZN(n12783) );
  OR2_X1 U11223 ( .A1(n11101), .A2(n11100), .ZN(n13445) );
  OR2_X1 U11224 ( .A1(n12138), .A2(n12137), .ZN(n12152) );
  AND2_X1 U11225 ( .A1(n10660), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10366) );
  AND2_X1 U11226 ( .A1(n9745), .A2(n10809), .ZN(n12523) );
  INV_X1 U11227 ( .A(n12481), .ZN(n12534) );
  BUF_X1 U11228 ( .A(n10314), .Z(n9757) );
  AND2_X1 U11230 ( .A1(n12753), .A2(n10120), .ZN(n10119) );
  AND2_X1 U11231 ( .A1(n11922), .A2(n11918), .ZN(n12002) );
  AND2_X1 U11232 ( .A1(n11919), .A2(n11921), .ZN(n12000) );
  NAND2_X1 U11233 ( .A1(n9722), .A2(n13748), .ZN(n20721) );
  INV_X1 U11234 ( .A(n13445), .ZN(n20125) );
  NOR2_X2 U11235 ( .A1(n12152), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n12157) );
  OAI21_X1 U11236 ( .B1(n15033), .B2(n15034), .A(n12765), .ZN(n12770) );
  OR2_X1 U11237 ( .A1(n12147), .A2(n12146), .ZN(n12148) );
  XNOR2_X1 U11238 ( .A(n13277), .B(n10284), .ZN(n13341) );
  NOR2_X1 U11240 ( .A1(n17800), .A2(n17811), .ZN(n17777) );
  INV_X1 U11241 ( .A(n11879), .ZN(n14191) );
  INV_X1 U11242 ( .A(n19969), .ZN(n19982) );
  NAND2_X1 U11243 ( .A1(n10724), .A2(n12247), .ZN(n12180) );
  INV_X1 U11244 ( .A(n19173), .ZN(n19180) );
  INV_X1 U11246 ( .A(n17877), .ZN(n17864) );
  INV_X1 U11247 ( .A(n19932), .ZN(n15894) );
  XOR2_X1 U11248 ( .A(n15133), .B(n15132), .Z(n15372) );
  INV_X1 U11249 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14108) );
  AND2_X1 U11250 ( .A1(n10927), .A2(n13460), .ZN(n11136) );
  OR2_X1 U11251 ( .A1(n18813), .A2(n17872), .ZN(n9718) );
  AND2_X2 U11252 ( .A1(n10238), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9745) );
  AND3_X2 U11253 ( .A1(n10689), .A2(n10758), .A3(n10737), .ZN(n10752) );
  NAND2_X2 U11254 ( .A1(n12302), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9763) );
  NAND2_X2 U11255 ( .A1(n15057), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15058) );
  NAND2_X2 U11256 ( .A1(n13250), .A2(n13249), .ZN(n13257) );
  NAND2_X2 U11257 ( .A1(n10031), .A2(n11175), .ZN(n11177) );
  NAND2_X2 U11259 ( .A1(n12401), .A2(n12400), .ZN(n13417) );
  OR2_X2 U11260 ( .A1(n14589), .A2(n16025), .ZN(n9942) );
  INV_X2 U11261 ( .A(n14952), .ZN(n12464) );
  NOR2_X4 U11262 ( .A1(n12792), .A2(n12783), .ZN(n12834) );
  OAI21_X2 U11263 ( .B1(n12327), .B2(n12762), .A(n19000), .ZN(n12054) );
  NOR2_X2 U11264 ( .A1(n12085), .A2(n12083), .ZN(n12102) );
  NAND2_X1 U11265 ( .A1(n20212), .A2(n11275), .ZN(n20377) );
  INV_X1 U11266 ( .A(n20212), .ZN(n11193) );
  NAND2_X2 U11267 ( .A1(n15251), .A2(n12335), .ZN(n12343) );
  NAND3_X2 U11268 ( .A1(n10093), .A2(n10092), .A3(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15251) );
  XNOR2_X2 U11269 ( .A(n13640), .B(n13549), .ZN(n13639) );
  NAND2_X2 U11270 ( .A1(n9876), .A2(n9874), .ZN(n13640) );
  NAND2_X2 U11271 ( .A1(n19193), .A2(n19209), .ZN(n19194) );
  XNOR2_X2 U11272 ( .A(n12322), .B(n12321), .ZN(n19193) );
  XNOR2_X2 U11273 ( .A(n12387), .B(n12385), .ZN(n13301) );
  NAND2_X2 U11274 ( .A1(n12375), .A2(n12374), .ZN(n12387) );
  NAND2_X2 U11275 ( .A1(n12320), .A2(n12319), .ZN(n12321) );
  NAND2_X2 U11276 ( .A1(n14929), .A2(n10132), .ZN(n14917) );
  XNOR2_X2 U11277 ( .A(n12024), .B(n12022), .ZN(n12325) );
  XNOR2_X2 U11278 ( .A(n13712), .B(n13660), .ZN(n13711) );
  NAND2_X2 U11279 ( .A1(n13642), .A2(n13641), .ZN(n13712) );
  NOR2_X4 U11280 ( .A1(n15068), .A2(n15056), .ZN(n15301) );
  NOR2_X2 U11281 ( .A1(n12991), .A2(n12990), .ZN(n18234) );
  OAI21_X2 U11282 ( .B1(n13478), .B2(n12396), .A(n12395), .ZN(n12397) );
  NOR3_X2 U11283 ( .A1(n17651), .A2(n17566), .A3(n17921), .ZN(n17558) );
  NOR2_X2 U11284 ( .A1(n17567), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17566) );
  NAND2_X1 U11285 ( .A1(n15159), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16175) );
  NOR2_X1 U11286 ( .A1(n14778), .A2(n14759), .ZN(n14760) );
  NOR2_X1 U11287 ( .A1(n12175), .A2(n10715), .ZN(n12758) );
  XNOR2_X1 U11288 ( .A(n12307), .B(n12306), .ZN(n12322) );
  NAND2_X1 U11289 ( .A1(n9856), .A2(n11934), .ZN(n11997) );
  AND2_X1 U11291 ( .A1(n11920), .A2(n11918), .ZN(n12008) );
  AND2_X1 U11292 ( .A1(n11920), .A2(n11917), .ZN(n19353) );
  AND2_X1 U11293 ( .A1(n11342), .A2(n11279), .ZN(n9804) );
  NAND2_X1 U11294 ( .A1(n11361), .A2(n11360), .ZN(n20182) );
  INV_X4 U11295 ( .A(n18654), .ZN(n18094) );
  NOR2_X1 U11296 ( .A1(n9891), .A2(n9890), .ZN(n15659) );
  CLKBUF_X2 U11297 ( .A(n10800), .Z(n10913) );
  AND2_X2 U11298 ( .A1(n12263), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10787) );
  CLKBUF_X1 U11299 ( .A(n11183), .Z(n11184) );
  AOI22_X1 U11300 ( .A1(n10030), .A2(n10029), .B1(n13445), .B2(n11733), .ZN(
        n10028) );
  INV_X1 U11301 ( .A(n13751), .ZN(n9722) );
  INV_X2 U11302 ( .A(n17330), .ZN(n18245) );
  NAND2_X2 U11303 ( .A1(n9945), .A2(n9793), .ZN(n13751) );
  NAND2_X2 U11304 ( .A1(n20125), .A2(n13360), .ZN(n11780) );
  INV_X2 U11305 ( .A(n10741), .ZN(n12150) );
  BUF_X2 U11306 ( .A(n11932), .Z(n9743) );
  AND2_X1 U11307 ( .A1(n11167), .A2(n11156), .ZN(n11102) );
  NOR2_X1 U11308 ( .A1(n12800), .A2(n12799), .ZN(n16337) );
  NAND2_X2 U11309 ( .A1(n16269), .A2(n11932), .ZN(n12247) );
  AND4_X1 U11310 ( .A1(n11036), .A2(n11035), .A3(n11034), .A4(n11033), .ZN(
        n11048) );
  AND4_X1 U11311 ( .A1(n11053), .A2(n11052), .A3(n11051), .A4(n11050), .ZN(
        n11069) );
  AND4_X1 U11312 ( .A1(n11057), .A2(n11056), .A3(n11055), .A4(n11054), .ZN(
        n11068) );
  INV_X1 U11313 ( .A(n17117), .ZN(n16869) );
  BUF_X2 U11314 ( .A(n11643), .Z(n9741) );
  CLKBUF_X2 U11315 ( .A(n12867), .Z(n17189) );
  CLKBUF_X2 U11316 ( .A(n11237), .Z(n11637) );
  CLKBUF_X2 U11317 ( .A(n11597), .Z(n14111) );
  INV_X4 U11318 ( .A(n16909), .ZN(n9720) );
  CLKBUF_X2 U11319 ( .A(n11260), .Z(n14112) );
  CLKBUF_X2 U11320 ( .A(n11253), .Z(n11635) );
  CLKBUF_X2 U11321 ( .A(n11095), .Z(n14117) );
  CLKBUF_X2 U11322 ( .A(n11252), .Z(n14119) );
  INV_X1 U11323 ( .A(n10128), .ZN(n17173) );
  NOR2_X2 U11324 ( .A1(n12783), .A2(n12789), .ZN(n12867) );
  AND2_X2 U11325 ( .A1(n14149), .A2(n14718), .ZN(n10928) );
  NOR2_X4 U11326 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15569) );
  INV_X4 U11327 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18812) );
  AOI21_X1 U11328 ( .B1(n15277), .B2(n12728), .A(n15053), .ZN(n15285) );
  AND2_X1 U11329 ( .A1(n15159), .A2(n15420), .ZN(n15172) );
  NOR2_X1 U11330 ( .A1(n15165), .A2(n15127), .ZN(n9873) );
  NAND2_X2 U11331 ( .A1(n14501), .A2(n14177), .ZN(n14443) );
  OAI21_X1 U11332 ( .B1(n14155), .B2(n14154), .A(n14153), .ZN(n14220) );
  AOI21_X1 U11333 ( .B1(n11723), .B2(n14241), .A(n14155), .ZN(n14441) );
  OAI21_X2 U11334 ( .B1(n15174), .B2(n12131), .A(n12130), .ZN(n15098) );
  OAI21_X1 U11335 ( .B1(n14256), .B2(n14258), .A(n14257), .ZN(n14465) );
  CLKBUF_X1 U11336 ( .A(n14240), .Z(n14257) );
  OAI21_X1 U11337 ( .B1(n15120), .B2(n12082), .A(n15122), .ZN(n15123) );
  OAI21_X1 U11338 ( .B1(n14507), .B2(n9851), .A(n14545), .ZN(n14501) );
  CLKBUF_X1 U11339 ( .A(n14255), .Z(n14256) );
  OR2_X1 U11340 ( .A1(n15748), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14507) );
  XNOR2_X1 U11341 ( .A(n12747), .B(n12746), .ZN(n12774) );
  AND2_X1 U11342 ( .A1(n12627), .A2(n12625), .ZN(n10144) );
  XNOR2_X1 U11343 ( .A(n14880), .B(n12740), .ZN(n15270) );
  OAI21_X1 U11344 ( .B1(n14168), .B2(n14160), .A(n9879), .ZN(n9880) );
  INV_X1 U11345 ( .A(n14881), .ZN(n14880) );
  AND3_X1 U11346 ( .A1(n15238), .A2(n15528), .A3(n15241), .ZN(n12058) );
  NAND3_X1 U11347 ( .A1(n14558), .A2(n14159), .A3(n14167), .ZN(n14168) );
  AND3_X1 U11348 ( .A1(n12333), .A2(n10095), .A3(n12330), .ZN(n10091) );
  NOR2_X1 U11349 ( .A1(n12764), .A2(n12763), .ZN(n12765) );
  AND2_X1 U11350 ( .A1(n10904), .A2(n10019), .ZN(n12300) );
  AND2_X1 U11351 ( .A1(n14587), .A2(n9940), .ZN(n9939) );
  NOR2_X1 U11352 ( .A1(n14897), .A2(n14898), .ZN(n10904) );
  AOI21_X1 U11353 ( .B1(n10119), .B2(n12754), .A(n12755), .ZN(n10117) );
  NOR2_X1 U11354 ( .A1(n10614), .A2(n10615), .ZN(n12736) );
  XNOR2_X1 U11355 ( .A(n12345), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n15231) );
  NAND2_X1 U11356 ( .A1(n12759), .A2(n9918), .ZN(n15035) );
  OR2_X1 U11357 ( .A1(n12566), .A2(n12586), .ZN(n10132) );
  OR2_X1 U11358 ( .A1(n17540), .A2(n12904), .ZN(n10103) );
  XNOR2_X1 U11359 ( .A(n12766), .B(n10716), .ZN(n12759) );
  OR2_X1 U11360 ( .A1(n12336), .A2(n12158), .ZN(n12345) );
  AND2_X1 U11361 ( .A1(n12326), .A2(n13970), .ZN(n13964) );
  OR2_X1 U11362 ( .A1(n16094), .A2(n12158), .ZN(n12172) );
  AND2_X1 U11363 ( .A1(n9966), .A2(n9965), .ZN(n9964) );
  NOR2_X1 U11364 ( .A1(n12024), .A2(n12023), .ZN(n12047) );
  NAND2_X1 U11365 ( .A1(n13894), .A2(n13893), .ZN(n15971) );
  NAND2_X1 U11366 ( .A1(n14795), .A2(n9781), .ZN(n14778) );
  XNOR2_X1 U11367 ( .A(n14209), .B(n14208), .ZN(n14588) );
  NAND2_X1 U11368 ( .A1(n10714), .A2(n12166), .ZN(n12175) );
  NAND2_X1 U11369 ( .A1(n13803), .A2(n13802), .ZN(n13891) );
  INV_X1 U11370 ( .A(n12329), .ZN(n12045) );
  INV_X1 U11371 ( .A(n13854), .ZN(n10020) );
  NAND2_X1 U11372 ( .A1(n17599), .A2(n12902), .ZN(n17567) );
  OR2_X1 U11373 ( .A1(n12140), .A2(n12158), .ZN(n12141) );
  AND2_X1 U11374 ( .A1(n12018), .A2(n12017), .ZN(n12022) );
  AND2_X1 U11375 ( .A1(n12044), .A2(n12043), .ZN(n12329) );
  NOR2_X1 U11376 ( .A1(n13573), .A2(n13674), .ZN(n13672) );
  NOR2_X1 U11377 ( .A1(n19439), .A2(n19609), .ZN(n19424) );
  OR2_X1 U11378 ( .A1(n12040), .A2(n12039), .ZN(n12044) );
  NOR2_X1 U11379 ( .A1(n19610), .A2(n19609), .ZN(n19664) );
  AND2_X1 U11380 ( .A1(n9732), .A2(n9785), .ZN(n13728) );
  OAI21_X1 U11381 ( .B1(n16508), .B2(n16498), .A(n9982), .ZN(n9985) );
  AND2_X2 U11382 ( .A1(n13417), .A2(n10024), .ZN(n9732) );
  AND2_X1 U11383 ( .A1(n13900), .A2(n13899), .ZN(n13901) );
  NAND2_X1 U11384 ( .A1(n9896), .A2(n9895), .ZN(n17664) );
  AND4_X1 U11385 ( .A1(n11914), .A2(n11925), .A3(n11924), .A4(n11912), .ZN(
        n9859) );
  OR2_X1 U11386 ( .A1(n17675), .A2(n18011), .ZN(n9896) );
  INV_X1 U11387 ( .A(n9718), .ZN(n9758) );
  OR2_X1 U11388 ( .A1(n16510), .A2(n17514), .ZN(n16508) );
  XNOR2_X1 U11389 ( .A(n13476), .B(n13477), .ZN(n19818) );
  OR2_X1 U11390 ( .A1(n14344), .A2(n14336), .ZN(n14334) );
  AOI211_X2 U11391 ( .C1(n19434), .C2(n10692), .A(n19734), .B(n9838), .ZN(
        n19455) );
  OR2_X1 U11392 ( .A1(n15843), .A2(n14342), .ZN(n14344) );
  NOR2_X1 U11393 ( .A1(n13629), .A2(n13630), .ZN(n13628) );
  NAND2_X1 U11394 ( .A1(n12134), .A2(n12155), .ZN(n12090) );
  NOR2_X1 U11395 ( .A1(n16519), .A2(n16518), .ZN(n16517) );
  NAND2_X1 U11396 ( .A1(n9798), .A2(n11375), .ZN(n13574) );
  NAND2_X1 U11397 ( .A1(n10833), .A2(n10832), .ZN(n13629) );
  XNOR2_X1 U11398 ( .A(n13895), .B(n11337), .ZN(n13905) );
  NAND2_X1 U11399 ( .A1(n11322), .A2(n9937), .ZN(n13895) );
  NAND2_X1 U11400 ( .A1(n10085), .A2(n10084), .ZN(n16195) );
  AND2_X1 U11401 ( .A1(n13256), .A2(n12384), .ZN(n13302) );
  NOR2_X2 U11402 ( .A1(n17448), .A2(n16439), .ZN(n17869) );
  NOR2_X2 U11403 ( .A1(n14071), .A2(n14072), .ZN(n14080) );
  NOR2_X1 U11404 ( .A1(n20249), .A2(n20147), .ZN(n20632) );
  NOR2_X1 U11405 ( .A1(n20249), .A2(n20143), .ZN(n20625) );
  NOR2_X1 U11406 ( .A1(n20249), .A2(n20138), .ZN(n20619) );
  NAND2_X2 U11407 ( .A1(n14409), .A2(n13569), .ZN(n14431) );
  NOR2_X1 U11408 ( .A1(n20249), .A2(n20134), .ZN(n20613) );
  NOR2_X1 U11409 ( .A1(n20249), .A2(n20129), .ZN(n20607) );
  OR2_X1 U11410 ( .A1(n14032), .A2(n14031), .ZN(n14071) );
  NOR2_X1 U11411 ( .A1(n20249), .A2(n20119), .ZN(n20595) );
  NOR2_X1 U11412 ( .A1(n20249), .A2(n20103), .ZN(n20584) );
  NOR2_X1 U11413 ( .A1(n20249), .A2(n20124), .ZN(n20601) );
  NAND2_X1 U11414 ( .A1(n9804), .A2(n20097), .ZN(n11377) );
  AOI21_X1 U11415 ( .B1(n11896), .B2(n9867), .A(n9797), .ZN(n13421) );
  OAI21_X1 U11416 ( .B1(n20182), .B2(n11525), .A(n11364), .ZN(n13498) );
  NAND2_X1 U11417 ( .A1(n15591), .A2(n12379), .ZN(n12375) );
  AND2_X1 U11418 ( .A1(n13258), .A2(n19038), .ZN(n11917) );
  AND2_X1 U11419 ( .A1(n15568), .A2(n19038), .ZN(n11918) );
  AND2_X1 U11420 ( .A1(n11909), .A2(n14102), .ZN(n11921) );
  NOR2_X1 U11421 ( .A1(n17568), .A2(n16555), .ZN(n16554) );
  NAND2_X1 U11422 ( .A1(n12378), .A2(n12377), .ZN(n14104) );
  AND2_X1 U11423 ( .A1(n14102), .A2(n11908), .ZN(n11926) );
  NAND2_X1 U11424 ( .A1(n16050), .A2(n16049), .ZN(n16052) );
  NAND2_X1 U11425 ( .A1(n12078), .A2(n12155), .ZN(n12073) );
  NOR2_X2 U11426 ( .A1(n19237), .A2(n19253), .ZN(n19238) );
  AND2_X1 U11427 ( .A1(n16561), .A2(n16469), .ZN(n16555) );
  AND2_X1 U11428 ( .A1(n13813), .A2(n13814), .ZN(n16050) );
  AOI21_X2 U11429 ( .B1(n12777), .B2(n18874), .A(n9993), .ZN(n19019) );
  NAND2_X1 U11430 ( .A1(n18651), .A2(n9889), .ZN(n18654) );
  INV_X2 U11431 ( .A(n17438), .ZN(n17439) );
  AOI21_X1 U11432 ( .B1(n18680), .B2(n10145), .A(n15672), .ZN(n15768) );
  NAND2_X1 U11433 ( .A1(n10777), .A2(n10776), .ZN(n10782) );
  AND2_X1 U11434 ( .A1(n16585), .A2(n16469), .ZN(n16576) );
  NAND2_X1 U11435 ( .A1(n11284), .A2(n11283), .ZN(n20244) );
  OR2_X1 U11436 ( .A1(n9802), .A2(n19237), .ZN(n12155) );
  NAND2_X1 U11437 ( .A1(n11205), .A2(n11204), .ZN(n11206) );
  NAND2_X1 U11438 ( .A1(n10806), .A2(n10805), .ZN(n10811) );
  NAND2_X1 U11439 ( .A1(n10757), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10807) );
  INV_X1 U11440 ( .A(n12020), .ZN(n9914) );
  NOR2_X1 U11441 ( .A1(n15661), .A2(n15664), .ZN(n18681) );
  OAI21_X1 U11442 ( .B1(n13024), .B2(n15669), .A(n13023), .ZN(n13032) );
  NAND2_X1 U11443 ( .A1(n10261), .A2(n10075), .ZN(n13275) );
  NOR2_X2 U11444 ( .A1(n16337), .A2(n12892), .ZN(n17782) );
  AOI21_X1 U11445 ( .B1(n12742), .B2(P2_REIP_REG_1__SCAN_IN), .A(n10780), .ZN(
        n10781) );
  AND4_X1 U11446 ( .A1(n10765), .A2(n10764), .A3(n10808), .A4(n10763), .ZN(
        n10766) );
  AND3_X1 U11447 ( .A1(n13022), .A2(n13021), .A3(n13020), .ZN(n13023) );
  AND2_X1 U11448 ( .A1(n11982), .A2(n11971), .ZN(n11993) );
  OR2_X1 U11449 ( .A1(n12308), .A2(n10528), .ZN(n10075) );
  INV_X2 U11450 ( .A(n10856), .ZN(n12741) );
  INV_X1 U11451 ( .A(n10787), .ZN(n10856) );
  AND2_X1 U11452 ( .A1(n13019), .A2(n13018), .ZN(n13020) );
  NOR2_X1 U11453 ( .A1(n11164), .A2(n13398), .ZN(n11173) );
  AND2_X1 U11454 ( .A1(n12211), .A2(n10736), .ZN(n12290) );
  AND2_X1 U11455 ( .A1(n17542), .A2(n9835), .ZN(n16321) );
  NAND2_X1 U11456 ( .A1(n12220), .A2(n10740), .ZN(n12251) );
  NOR2_X1 U11457 ( .A1(n12019), .A2(n9916), .ZN(n9915) );
  NAND2_X1 U11458 ( .A1(n12221), .A2(n10760), .ZN(n9863) );
  NOR2_X1 U11459 ( .A1(n13426), .A2(n14140), .ZN(n13405) );
  AND2_X1 U11460 ( .A1(n11879), .A2(n11803), .ZN(n13702) );
  INV_X1 U11461 ( .A(n20721), .ZN(n13955) );
  NAND2_X1 U11462 ( .A1(n11080), .A2(n11102), .ZN(n11114) );
  NAND2_X1 U11463 ( .A1(n11249), .A2(n13751), .ZN(n13746) );
  AND2_X1 U11464 ( .A1(n12222), .A2(n12707), .ZN(n10740) );
  AND3_X1 U11465 ( .A1(n12180), .A2(n12258), .A3(n10726), .ZN(n9799) );
  NOR2_X1 U11466 ( .A1(n17561), .A2(n17562), .ZN(n17542) );
  INV_X1 U11467 ( .A(n13751), .ZN(n20120) );
  NOR2_X1 U11468 ( .A1(n11780), .A2(n20148), .ZN(n11158) );
  AND2_X1 U11469 ( .A1(n15641), .A2(n18238), .ZN(n18648) );
  AND2_X1 U11470 ( .A1(n17330), .A2(n9888), .ZN(n13031) );
  AND2_X1 U11471 ( .A1(n12707), .A2(n19385), .ZN(n10281) );
  NAND3_X1 U11472 ( .A1(n13003), .A2(n13002), .A3(n13001), .ZN(n17330) );
  INV_X1 U11473 ( .A(n18217), .ZN(n17448) );
  AND2_X1 U11474 ( .A1(n12216), .A2(n9855), .ZN(n10734) );
  CLKBUF_X1 U11475 ( .A(n10761), .Z(n19245) );
  AND2_X1 U11476 ( .A1(n10721), .A2(n12707), .ZN(n12724) );
  NAND4_X1 U11477 ( .A1(n9811), .A2(n9764), .A3(n9765), .A4(n12843), .ZN(
        n13046) );
  INV_X1 U11478 ( .A(n10723), .ZN(n10724) );
  CLKBUF_X1 U11479 ( .A(n10725), .Z(n12215) );
  OR2_X1 U11480 ( .A1(n11232), .A2(n11231), .ZN(n13954) );
  AND2_X1 U11481 ( .A1(n10630), .A2(n10728), .ZN(n12216) );
  INV_X1 U11482 ( .A(n16269), .ZN(n10690) );
  NOR2_X2 U11483 ( .A1(n12923), .A2(n12922), .ZN(n18217) );
  NOR2_X1 U11484 ( .A1(n12878), .A2(n12877), .ZN(n17876) );
  CLKBUF_X1 U11485 ( .A(n11730), .Z(n14185) );
  CLKBUF_X1 U11486 ( .A(n10728), .Z(n10729) );
  NAND4_X2 U11487 ( .A1(n11049), .A2(n11048), .A3(n11047), .A4(n11046), .ZN(
        n11156) );
  NAND2_X1 U11488 ( .A1(n10642), .A2(n10641), .ZN(n10725) );
  OR2_X2 U11489 ( .A1(n11113), .A2(n11112), .ZN(n13360) );
  NAND2_X1 U11490 ( .A1(n10629), .A2(n10628), .ZN(n10728) );
  NAND2_X1 U11491 ( .A1(n10653), .A2(n10654), .ZN(n12201) );
  NAND4_X2 U11492 ( .A1(n11069), .A2(n11068), .A3(n11067), .A4(n11066), .ZN(
        n11165) );
  NAND2_X2 U11493 ( .A1(n11079), .A2(n9882), .ZN(n11730) );
  NAND2_X2 U11494 ( .A1(n10669), .A2(n10668), .ZN(n16269) );
  AND4_X1 U11495 ( .A1(n10429), .A2(n10428), .A3(n10427), .A4(n10426), .ZN(
        n10430) );
  AND4_X1 U11496 ( .A1(n11020), .A2(n11019), .A3(n11018), .A4(n11017), .ZN(
        n11026) );
  AND4_X1 U11497 ( .A1(n11045), .A2(n11044), .A3(n11043), .A4(n11042), .ZN(
        n11046) );
  AND4_X1 U11498 ( .A1(n11071), .A2(n11074), .A3(n11072), .A4(n11073), .ZN(
        n9882) );
  AND4_X1 U11499 ( .A1(n11118), .A2(n11117), .A3(n11116), .A4(n11115), .ZN(
        n11134) );
  AND4_X1 U11500 ( .A1(n11122), .A2(n11121), .A3(n11120), .A4(n11119), .ZN(
        n11133) );
  AND4_X1 U11501 ( .A1(n11040), .A2(n11039), .A3(n11038), .A4(n11037), .ZN(
        n11047) );
  AND4_X1 U11502 ( .A1(n11024), .A2(n11023), .A3(n11022), .A4(n11021), .ZN(
        n11025) );
  AND4_X1 U11503 ( .A1(n11061), .A2(n11060), .A3(n11059), .A4(n11058), .ZN(
        n11067) );
  AND4_X1 U11504 ( .A1(n11016), .A2(n11015), .A3(n11014), .A4(n11013), .ZN(
        n11027) );
  AND4_X1 U11505 ( .A1(n11130), .A2(n11129), .A3(n11128), .A4(n11127), .ZN(
        n11131) );
  NAND2_X2 U11506 ( .A1(n19879), .A2(n19760), .ZN(n19801) );
  INV_X2 U11507 ( .A(n20685), .ZN(n9723) );
  AND4_X1 U11508 ( .A1(n11078), .A2(n11077), .A3(n11076), .A4(n11075), .ZN(
        n11079) );
  AND4_X1 U11509 ( .A1(n11148), .A2(n11147), .A3(n11146), .A4(n11145), .ZN(
        n11154) );
  INV_X2 U11510 ( .A(n17187), .ZN(n17165) );
  NAND2_X2 U11511 ( .A1(n18842), .A2(n18737), .ZN(n18781) );
  NOR2_X2 U11512 ( .A1(n20107), .A2(n20106), .ZN(n20108) );
  AND4_X1 U11513 ( .A1(n11032), .A2(n11031), .A3(n11030), .A4(n11029), .ZN(
        n11049) );
  INV_X2 U11514 ( .A(n16424), .ZN(U215) );
  INV_X1 U11515 ( .A(n10957), .ZN(n9725) );
  BUF_X2 U11516 ( .A(n12539), .Z(n10380) );
  BUF_X2 U11517 ( .A(n12833), .Z(n17183) );
  BUF_X2 U11518 ( .A(n12836), .Z(n17167) );
  CLKBUF_X3 U11519 ( .A(n16864), .Z(n12992) );
  CLKBUF_X2 U11520 ( .A(n12833), .Z(n16891) );
  BUF_X2 U11521 ( .A(n12867), .Z(n17163) );
  INV_X1 U11522 ( .A(n12790), .ZN(n12868) );
  NOR2_X2 U11523 ( .A1(n18451), .A2(n18385), .ZN(n18437) );
  CLKBUF_X1 U11524 ( .A(n13225), .Z(n13830) );
  INV_X2 U11525 ( .A(n16426), .ZN(n16428) );
  NAND2_X2 U11526 ( .A1(n18877), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n19797) );
  AND2_X2 U11527 ( .A1(n12690), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10367) );
  OR2_X1 U11528 ( .A1(n12793), .A2(n18665), .ZN(n16791) );
  NAND2_X1 U11529 ( .A1(n13459), .A2(n10928), .ZN(n11041) );
  OAI21_X1 U11530 ( .B1(n12717), .B2(n12716), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13225) );
  AND2_X2 U11531 ( .A1(n13460), .A2(n10930), .ZN(n11643) );
  INV_X2 U11532 ( .A(n18193), .ZN(n9726) );
  OR2_X1 U11533 ( .A1(n18665), .A2(n12791), .ZN(n10128) );
  INV_X2 U11534 ( .A(n19864), .ZN(n9727) );
  AND2_X2 U11535 ( .A1(n14718), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10926) );
  AND2_X2 U11536 ( .A1(n10921), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13460) );
  NAND2_X1 U11537 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n21023), .ZN(
        n12792) );
  AND3_X2 U11538 ( .A1(n10198), .A2(n10197), .A3(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n12690) );
  AND2_X2 U11539 ( .A1(n15580), .A2(n10197), .ZN(n12550) );
  NAND2_X1 U11540 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18665) );
  INV_X2 U11541 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10197) );
  INV_X2 U11542 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n10692) );
  BUF_X4 U11543 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n16229) );
  NAND2_X2 U11544 ( .A1(n15526), .A2(n12344), .ZN(n15229) );
  NAND2_X1 U11545 ( .A1(n13903), .A2(n9731), .ZN(n9728) );
  OR2_X1 U11546 ( .A1(n9730), .A2(n10067), .ZN(n9729) );
  INV_X1 U11547 ( .A(n14017), .ZN(n9730) );
  AND2_X1 U11548 ( .A1(n9806), .A2(n14017), .ZN(n9731) );
  NAND2_X1 U11549 ( .A1(n12021), .A2(n19015), .ZN(n12052) );
  AOI21_X2 U11550 ( .B1(n15387), .B2(n15388), .A(n15129), .ZN(n15143) );
  AND2_X1 U11551 ( .A1(n15406), .A2(n15403), .ZN(n15387) );
  INV_X1 U11552 ( .A(n9732), .ZN(n13538) );
  INV_X1 U11553 ( .A(n11156), .ZN(n20148) );
  NAND2_X1 U11554 ( .A1(n9877), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14459) );
  NOR2_X2 U11555 ( .A1(n17468), .A2(n17277), .ZN(n17272) );
  NOR2_X2 U11556 ( .A1(n17427), .A2(n17355), .ZN(n17353) );
  NAND2_X1 U11557 ( .A1(n15229), .A2(n9736), .ZN(n9733) );
  AND2_X2 U11558 ( .A1(n9733), .A2(n9734), .ZN(n15137) );
  OR2_X1 U11559 ( .A1(n9735), .A2(n12347), .ZN(n9734) );
  INV_X1 U11560 ( .A(n9790), .ZN(n9735) );
  AND2_X1 U11561 ( .A1(n15231), .A2(n9790), .ZN(n9736) );
  NAND2_X4 U11562 ( .A1(n11276), .A2(n20377), .ZN(n13669) );
  INV_X1 U11563 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9737) );
  AND2_X2 U11564 ( .A1(n10238), .A2(n9737), .ZN(n12539) );
  AND2_X1 U11565 ( .A1(n15569), .A2(n10197), .ZN(n9756) );
  INV_X2 U11566 ( .A(n20095), .ZN(n13664) );
  NAND2_X2 U11567 ( .A1(n13162), .A2(n20120), .ZN(n13447) );
  AND2_X2 U11568 ( .A1(n11182), .A2(n11135), .ZN(n13162) );
  CLKBUF_X1 U11569 ( .A(n13800), .Z(n9738) );
  NAND2_X1 U11570 ( .A1(n13714), .A2(n13713), .ZN(n13800) );
  INV_X1 U11571 ( .A(n9739), .ZN(n15097) );
  AND2_X2 U11572 ( .A1(n13860), .A2(n13924), .ZN(n13923) );
  AND2_X2 U11573 ( .A1(n14322), .A2(n11659), .ZN(n14317) );
  NOR2_X2 U11574 ( .A1(n13819), .A2(n11421), .ZN(n13860) );
  NAND2_X1 U11575 ( .A1(n15971), .A2(n15973), .ZN(n13903) );
  OR2_X1 U11576 ( .A1(n14160), .A2(n14563), .ZN(n15946) );
  NAND2_X1 U11577 ( .A1(n11901), .A2(n11900), .ZN(n11899) );
  NAND2_X1 U11579 ( .A1(n9868), .A2(n9867), .ZN(n9866) );
  NAND2_X1 U11581 ( .A1(n9854), .A2(n9853), .ZN(n10700) );
  NAND2_X1 U11582 ( .A1(n9854), .A2(n9853), .ZN(n9740) );
  BUF_X8 U11583 ( .A(n11643), .Z(n9742) );
  NOR2_X2 U11584 ( .A1(n16269), .A2(n11932), .ZN(n10723) );
  XNOR2_X1 U11585 ( .A(n13480), .B(n20244), .ZN(n20349) );
  OR2_X1 U11586 ( .A1(n11192), .A2(n9932), .ZN(n9931) );
  INV_X2 U11587 ( .A(n10807), .ZN(n10795) );
  NAND2_X1 U11588 ( .A1(n11903), .A2(n11904), .ZN(n11908) );
  AND2_X2 U11589 ( .A1(n11165), .A2(n11156), .ZN(n11159) );
  INV_X2 U11590 ( .A(n10700), .ZN(n10741) );
  OAI21_X2 U11591 ( .B1(n10793), .B2(n9763), .A(n10792), .ZN(n10796) );
  NAND2_X1 U11592 ( .A1(n12302), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9762) );
  AND3_X1 U11593 ( .A1(n10630), .A2(n10742), .A3(n19228), .ZN(n10689) );
  INV_X2 U11594 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14718) );
  NOR2_X2 U11595 ( .A1(n10721), .A2(n9740), .ZN(n10727) );
  NAND2_X4 U11596 ( .A1(n10258), .A2(n10257), .ZN(n10721) );
  INV_X2 U11597 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10921) );
  OR2_X1 U11598 ( .A1(n11927), .A2(n11928), .ZN(n19494) );
  NAND2_X2 U11599 ( .A1(n15230), .A2(n12347), .ZN(n15159) );
  AND2_X1 U11600 ( .A1(n13468), .A2(n10928), .ZN(n9747) );
  AND2_X1 U11601 ( .A1(n13468), .A2(n10928), .ZN(n9748) );
  NAND2_X2 U11602 ( .A1(n9944), .A2(n14524), .ZN(n15928) );
  AND2_X1 U11603 ( .A1(n11157), .A2(n11180), .ZN(n13201) );
  AND2_X1 U11604 ( .A1(n11899), .A2(n11902), .ZN(n14102) );
  NOR2_X4 U11605 ( .A1(n18647), .A2(n18145), .ZN(n18052) );
  INV_X2 U11606 ( .A(n18656), .ZN(n18647) );
  AND2_X1 U11607 ( .A1(n10928), .A2(n10929), .ZN(n9749) );
  AND2_X1 U11608 ( .A1(n10928), .A2(n10929), .ZN(n9750) );
  NAND2_X2 U11609 ( .A1(n11180), .A2(n11730), .ZN(n11168) );
  INV_X4 U11610 ( .A(n11041), .ZN(n10968) );
  INV_X1 U11611 ( .A(n9762), .ZN(n10908) );
  AND2_X1 U11612 ( .A1(n10926), .A2(n10929), .ZN(n9759) );
  NOR2_X1 U11613 ( .A1(n12793), .A2(n16826), .ZN(n9753) );
  AND2_X1 U11614 ( .A1(n10927), .A2(n10929), .ZN(n9754) );
  AND2_X1 U11615 ( .A1(n10927), .A2(n10929), .ZN(n9755) );
  AND2_X1 U11616 ( .A1(n10927), .A2(n10929), .ZN(n11095) );
  NAND2_X2 U11617 ( .A1(n19194), .A2(n12324), .ZN(n13967) );
  INV_X2 U11618 ( .A(n11167), .ZN(n11222) );
  NAND2_X2 U11619 ( .A1(n15066), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15068) );
  OAI21_X2 U11620 ( .B1(n14894), .B2(n14887), .A(n12677), .ZN(n14878) );
  NOR2_X2 U11621 ( .A1(n14893), .A2(n14895), .ZN(n14894) );
  NOR2_X2 U11622 ( .A1(n13360), .A2(n13445), .ZN(n13470) );
  AND2_X2 U11623 ( .A1(n9739), .A2(n9850), .ZN(n15066) );
  AND2_X2 U11624 ( .A1(n15569), .A2(n9737), .ZN(n12540) );
  XNOR2_X1 U11625 ( .A(n13301), .B(n13302), .ZN(n19825) );
  INV_X1 U11628 ( .A(n14478), .ZN(n9877) );
  NAND3_X2 U11629 ( .A1(n9862), .A2(n15585), .A3(n9860), .ZN(n12302) );
  NAND2_X1 U11630 ( .A1(n10733), .A2(n16269), .ZN(n10760) );
  OAI21_X2 U11631 ( .B1(n13425), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11219), 
        .ZN(n11342) );
  NAND2_X2 U11632 ( .A1(n13480), .A2(n11208), .ZN(n13425) );
  AND2_X2 U11633 ( .A1(n10926), .A2(n10929), .ZN(n11149) );
  AND2_X1 U11634 ( .A1(n10927), .A2(n13460), .ZN(n9760) );
  OR2_X1 U11635 ( .A1(n11167), .A2(n20639), .ZN(n11270) );
  NAND2_X1 U11636 ( .A1(n10759), .A2(n19228), .ZN(n10743) );
  INV_X1 U11637 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10196) );
  NAND2_X1 U11638 ( .A1(n12046), .A2(n12045), .ZN(n12048) );
  NAND2_X1 U11639 ( .A1(n9796), .A2(n9768), .ZN(n12018) );
  NAND2_X1 U11640 ( .A1(n10732), .A2(n10731), .ZN(n9864) );
  NAND2_X1 U11641 ( .A1(n10727), .A2(n10730), .ZN(n10732) );
  NOR2_X1 U11642 ( .A1(n10729), .A2(n16269), .ZN(n10730) );
  NAND2_X1 U11643 ( .A1(n11322), .A2(n11385), .ZN(n11394) );
  OR2_X1 U11644 ( .A1(n13568), .A2(n20640), .ZN(n11354) );
  NOR2_X1 U11645 ( .A1(n11782), .A2(n20640), .ZN(n11413) );
  INV_X1 U11646 ( .A(n12049), .ZN(n9916) );
  NAND2_X1 U11647 ( .A1(n12464), .A2(n14953), .ZN(n14945) );
  NAND2_X1 U11648 ( .A1(n10023), .A2(n13856), .ZN(n10022) );
  INV_X1 U11649 ( .A(n13944), .ZN(n10023) );
  NAND2_X1 U11650 ( .A1(n12758), .A2(n12757), .ZN(n12766) );
  NOR2_X1 U11651 ( .A1(n9975), .A2(n9974), .ZN(n9973) );
  INV_X1 U11652 ( .A(n9976), .ZN(n9974) );
  NAND2_X1 U11653 ( .A1(n10087), .A2(n15513), .ZN(n10086) );
  INV_X1 U11654 ( .A(n14826), .ZN(n10087) );
  AND2_X1 U11655 ( .A1(n10011), .A2(n13485), .ZN(n10010) );
  INV_X1 U11656 ( .A(n13514), .ZN(n10011) );
  NAND2_X1 U11657 ( .A1(n9921), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13062) );
  NAND2_X1 U11658 ( .A1(n13738), .A2(n13737), .ZN(n19927) );
  INV_X1 U11659 ( .A(n11354), .ZN(n14137) );
  NAND2_X1 U11660 ( .A1(n11378), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11387) );
  AND3_X1 U11661 ( .A1(n14501), .A2(n14177), .A3(n9934), .ZN(n9933) );
  AND2_X1 U11662 ( .A1(n14178), .A2(n9935), .ZN(n9934) );
  NAND2_X1 U11663 ( .A1(n9877), .A2(n9791), .ZN(n14461) );
  NAND4_X1 U11664 ( .A1(n11191), .A2(n11190), .A3(n11189), .A4(n11188), .ZN(
        n11220) );
  NOR2_X1 U11665 ( .A1(n10193), .A2(n15049), .ZN(n10194) );
  AND2_X1 U11666 ( .A1(n15425), .A2(n12274), .ZN(n15556) );
  OR2_X1 U11667 ( .A1(n13254), .A2(n13253), .ZN(n13256) );
  NAND2_X1 U11668 ( .A1(n13059), .A2(n17804), .ZN(n17794) );
  AND2_X1 U11669 ( .A1(n10099), .A2(n17813), .ZN(n17803) );
  INV_X1 U11670 ( .A(n18684), .ZN(n18069) );
  NAND2_X1 U11671 ( .A1(n21051), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11937) );
  OR2_X1 U11672 ( .A1(n12930), .A2(n12931), .ZN(n12926) );
  INV_X1 U11673 ( .A(n11386), .ZN(n11322) );
  AND2_X1 U11674 ( .A1(n10090), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10368) );
  INV_X1 U11675 ( .A(n12233), .ZN(n10090) );
  NOR2_X1 U11676 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12542) );
  AOI21_X1 U11677 ( .B1(n10367), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n10089), .ZN(n10240) );
  AND2_X1 U11678 ( .A1(n10368), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n10089) );
  AOI22_X1 U11679 ( .A1(n12550), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10216) );
  AND2_X1 U11680 ( .A1(n12225), .A2(n12224), .ZN(n12267) );
  INV_X1 U11681 ( .A(n11927), .ZN(n11919) );
  NAND2_X1 U11682 ( .A1(n15591), .A2(n13777), .ZN(n11929) );
  AOI22_X1 U11683 ( .A1(n10660), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9745), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10621) );
  NAND2_X1 U11684 ( .A1(n12550), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(
        n10617) );
  NOR2_X1 U11686 ( .A1(n12201), .A2(n10725), .ZN(n9855) );
  INV_X1 U11687 ( .A(n18225), .ZN(n9888) );
  INV_X1 U11688 ( .A(n14270), .ZN(n10033) );
  OR2_X1 U11689 ( .A1(n10040), .A2(n10038), .ZN(n10037) );
  INV_X1 U11690 ( .A(n14341), .ZN(n10038) );
  OR2_X1 U11691 ( .A1(n10041), .A2(n14408), .ZN(n10040) );
  INV_X1 U11692 ( .A(n14130), .ZN(n11714) );
  NAND2_X1 U11693 ( .A1(n14716), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n14130) );
  AND2_X1 U11694 ( .A1(n10045), .A2(n9846), .ZN(n10044) );
  OR2_X1 U11695 ( .A1(n10047), .A2(n10046), .ZN(n10045) );
  AND2_X1 U11696 ( .A1(n13995), .A2(n14063), .ZN(n10046) );
  NAND2_X1 U11697 ( .A1(n13923), .A2(n10047), .ZN(n14064) );
  NAND2_X1 U11698 ( .A1(n14314), .A2(n14291), .ZN(n14271) );
  OR2_X1 U11699 ( .A1(n14326), .A2(n14320), .ZN(n9961) );
  NOR2_X1 U11700 ( .A1(n14534), .A2(n14536), .ZN(n14170) );
  NOR2_X1 U11701 ( .A1(n9958), .A2(n13865), .ZN(n9957) );
  INV_X1 U11702 ( .A(n13926), .ZN(n9958) );
  INV_X1 U11703 ( .A(n13866), .ZN(n9956) );
  INV_X1 U11704 ( .A(n13948), .ZN(n10068) );
  INV_X1 U11705 ( .A(n11823), .ZN(n11883) );
  INV_X1 U11706 ( .A(n11878), .ZN(n11888) );
  OR2_X1 U11707 ( .A1(n13950), .A2(n13520), .ZN(n11246) );
  AOI21_X1 U11708 ( .B1(n13596), .B2(n16064), .A(n15731), .ZN(n20104) );
  NOR2_X1 U11709 ( .A1(n11167), .A2(n11730), .ZN(n11157) );
  NAND2_X1 U11710 ( .A1(n9917), .A2(n9843), .ZN(n12111) );
  NAND2_X1 U11711 ( .A1(n12073), .A2(n10708), .ZN(n12085) );
  AND2_X1 U11712 ( .A1(n10386), .A2(n10385), .ZN(n12016) );
  OAI22_X1 U11713 ( .A1(n10807), .A2(n10809), .B1(n10808), .B2(n19824), .ZN(
        n10810) );
  INV_X1 U11714 ( .A(n15543), .ZN(n10072) );
  AND4_X1 U11715 ( .A1(n10404), .A2(n10403), .A3(n10402), .A4(n10401), .ZN(
        n10410) );
  NOR2_X1 U11716 ( .A1(n15059), .A2(n10005), .ZN(n10004) );
  INV_X1 U11717 ( .A(n14922), .ZN(n10016) );
  NOR2_X1 U11718 ( .A1(n14729), .A2(n10018), .ZN(n10017) );
  INV_X1 U11719 ( .A(n14744), .ZN(n10018) );
  INV_X1 U11720 ( .A(n15207), .ZN(n10113) );
  NAND2_X1 U11721 ( .A1(n10845), .A2(n10009), .ZN(n10008) );
  INV_X1 U11722 ( .A(n13697), .ZN(n10009) );
  NOR2_X1 U11723 ( .A1(n15220), .A2(n9977), .ZN(n9976) );
  INV_X1 U11724 ( .A(n10124), .ZN(n9977) );
  AND4_X1 U11725 ( .A1(n10425), .A2(n10424), .A3(n10423), .A4(n10422), .ZN(
        n10431) );
  AND4_X1 U11726 ( .A1(n10418), .A2(n10417), .A3(n10416), .A4(n10415), .ZN(
        n10432) );
  AND4_X1 U11727 ( .A1(n10351), .A2(n10350), .A3(n10349), .A4(n10348), .ZN(
        n10357) );
  NAND2_X1 U11728 ( .A1(n11970), .A2(n11969), .ZN(n11996) );
  CLKBUF_X2 U11729 ( .A(n10266), .Z(n12733) );
  NAND2_X1 U11730 ( .A1(n9799), .A2(n9864), .ZN(n15585) );
  INV_X1 U11731 ( .A(n10758), .ZN(n12258) );
  INV_X1 U11732 ( .A(n11926), .ZN(n11928) );
  INV_X1 U11733 ( .A(n19838), .ZN(n15608) );
  NOR2_X1 U11734 ( .A1(n18213), .A2(n15662), .ZN(n15661) );
  NAND2_X1 U11735 ( .A1(n9980), .A2(n9979), .ZN(n16531) );
  INV_X1 U11736 ( .A(n17543), .ZN(n9979) );
  OR2_X2 U11737 ( .A1(n12783), .A2(n16826), .ZN(n17083) );
  INV_X1 U11738 ( .A(n16910), .ZN(n17187) );
  NOR2_X1 U11739 ( .A1(n12783), .A2(n18665), .ZN(n12833) );
  NOR2_X1 U11740 ( .A1(n13029), .A2(n16430), .ZN(n15664) );
  NAND2_X1 U11741 ( .A1(n17801), .A2(n12891), .ZN(n12894) );
  NAND2_X1 U11742 ( .A1(n17781), .A2(n10104), .ZN(n17692) );
  NOR2_X1 U11743 ( .A1(n17819), .A2(n9920), .ZN(n13057) );
  AOI21_X1 U11744 ( .B1(n17820), .B2(n17821), .A(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n9920) );
  NOR2_X1 U11745 ( .A1(n15765), .A2(n18245), .ZN(n13025) );
  INV_X2 U11746 ( .A(n14086), .ZN(n17162) );
  INV_X1 U11747 ( .A(n13702), .ZN(n14207) );
  OR2_X1 U11748 ( .A1(n13376), .A2(n11781), .ZN(n13453) );
  INV_X1 U11749 ( .A(n11159), .ZN(n14140) );
  NAND2_X1 U11750 ( .A1(n13534), .A2(n11367), .ZN(n13575) );
  OR2_X1 U11751 ( .A1(n11695), .A2(n14275), .ZN(n11705) );
  NAND2_X1 U11752 ( .A1(n14173), .A2(n14160), .ZN(n14500) );
  AND2_X1 U11753 ( .A1(n15927), .A2(n10146), .ZN(n10069) );
  NOR2_X1 U11754 ( .A1(n11594), .A2(n15831), .ZN(n11613) );
  NAND2_X1 U11755 ( .A1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n11613), .ZN(
        n11630) );
  AOI21_X1 U11756 ( .B1(n13896), .B2(n11413), .A(n11400), .ZN(n13707) );
  AOI21_X1 U11757 ( .B1(n13715), .B2(n11413), .A(n11384), .ZN(n13674) );
  OR2_X1 U11758 ( .A1(n11778), .A2(n11777), .ZN(n13496) );
  AND2_X1 U11759 ( .A1(n14160), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14174) );
  AND2_X1 U11760 ( .A1(n14524), .A2(n14175), .ZN(n9943) );
  INV_X1 U11761 ( .A(n13912), .ZN(n9878) );
  INV_X1 U11762 ( .A(n14580), .ZN(n15995) );
  INV_X1 U11763 ( .A(n13408), .ZN(n13403) );
  NAND2_X1 U11764 ( .A1(n11349), .A2(n13904), .ZN(n10050) );
  NAND2_X1 U11765 ( .A1(n11176), .A2(n10056), .ZN(n10053) );
  NOR2_X1 U11766 ( .A1(n9949), .A2(n9946), .ZN(n9945) );
  INV_X1 U11767 ( .A(n20097), .ZN(n13665) );
  NOR2_X1 U11768 ( .A1(n20413), .A2(n20249), .ZN(n20556) );
  AOI21_X1 U11769 ( .B1(n20517), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20249), 
        .ZN(n20587) );
  OR2_X1 U11770 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20104), .ZN(n20249) );
  INV_X1 U11771 ( .A(n9917), .ZN(n12113) );
  NAND2_X1 U11772 ( .A1(n9914), .A2(n9915), .ZN(n12056) );
  NAND2_X1 U11773 ( .A1(n9871), .A2(n10799), .ZN(n9868) );
  INV_X1 U11774 ( .A(n12232), .ZN(n16273) );
  NAND2_X1 U11775 ( .A1(n12300), .A2(n14882), .ZN(n14881) );
  AND2_X1 U11776 ( .A1(n13416), .A2(n9847), .ZN(n10025) );
  NAND2_X1 U11777 ( .A1(n14985), .A2(n10081), .ZN(n10614) );
  NOR3_X1 U11778 ( .A1(n9840), .A2(n10082), .A3(n10083), .ZN(n10081) );
  INV_X1 U11779 ( .A(n14968), .ZN(n10083) );
  INV_X1 U11780 ( .A(n14986), .ZN(n10082) );
  NAND2_X1 U11781 ( .A1(n14928), .A2(n14930), .ZN(n14929) );
  NOR2_X1 U11782 ( .A1(n10022), .A2(n9845), .ZN(n10021) );
  NAND2_X1 U11783 ( .A1(n13973), .A2(n10074), .ZN(n10073) );
  INV_X1 U11784 ( .A(n14832), .ZN(n10074) );
  INV_X1 U11785 ( .A(n15035), .ZN(n12764) );
  INV_X1 U11786 ( .A(n15082), .ZN(n9966) );
  OR2_X1 U11787 ( .A1(n15363), .A2(n15367), .ZN(n15349) );
  NAND2_X1 U11788 ( .A1(n10866), .A2(n10865), .ZN(n13940) );
  INV_X1 U11789 ( .A(n13105), .ZN(n10865) );
  INV_X1 U11790 ( .A(n13104), .ZN(n10866) );
  NOR2_X1 U11791 ( .A1(n9822), .A2(n10088), .ZN(n10084) );
  INV_X1 U11792 ( .A(n14824), .ZN(n10085) );
  INV_X1 U11793 ( .A(n13117), .ZN(n10088) );
  NAND2_X1 U11794 ( .A1(n13419), .A2(n9809), .ZN(n13540) );
  INV_X1 U11795 ( .A(n13964), .ZN(n10095) );
  NAND2_X1 U11796 ( .A1(n10203), .A2(n10809), .ZN(n10210) );
  NAND2_X1 U11797 ( .A1(n10208), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10209) );
  AND2_X1 U11798 ( .A1(n19818), .A2(n19846), .ZN(n19296) );
  NAND2_X1 U11799 ( .A1(n19818), .A2(n19110), .ZN(n19439) );
  INV_X1 U11800 ( .A(n19547), .ZN(n19323) );
  OR2_X1 U11801 ( .A1(n19818), .A2(n19110), .ZN(n19631) );
  OR2_X1 U11802 ( .A1(n19818), .A2(n19846), .ZN(n19610) );
  INV_X1 U11803 ( .A(n19436), .ZN(n19680) );
  OR2_X1 U11804 ( .A1(n19825), .A2(n19838), .ZN(n19815) );
  NAND2_X1 U11805 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19680), .ZN(n19253) );
  NAND2_X1 U11806 ( .A1(n10659), .A2(n10809), .ZN(n10669) );
  NOR2_X1 U11807 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n19861) );
  AOI21_X1 U11808 ( .B1(n16820), .B2(n9983), .A(n16820), .ZN(n9982) );
  OR2_X1 U11809 ( .A1(n16541), .A2(n16820), .ZN(n9980) );
  AOI21_X1 U11810 ( .B1(n16469), .B2(n17605), .A(n17588), .ZN(n9991) );
  OR2_X1 U11811 ( .A1(n16576), .A2(n17605), .ZN(n9992) );
  NOR2_X2 U11812 ( .A1(n12793), .A2(n16826), .ZN(n16910) );
  NAND2_X1 U11813 ( .A1(n18213), .A2(n18217), .ZN(n15765) );
  AND2_X1 U11814 ( .A1(n16672), .A2(n9989), .ZN(n9988) );
  INV_X1 U11815 ( .A(n17715), .ZN(n9989) );
  AND2_X1 U11816 ( .A1(n16302), .A2(n9930), .ZN(n17721) );
  XNOR2_X1 U11817 ( .A(n12894), .B(n12893), .ZN(n17788) );
  INV_X1 U11818 ( .A(n12895), .ZN(n12893) );
  NAND2_X1 U11819 ( .A1(n17788), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17787) );
  OAI21_X1 U11820 ( .B1(n17782), .B2(n12911), .A(n12910), .ZN(n15740) );
  NOR2_X1 U11821 ( .A1(n17527), .A2(n12900), .ZN(n16338) );
  AOI21_X1 U11822 ( .B1(n16340), .B2(n18069), .A(n16339), .ZN(n16343) );
  NAND2_X1 U11823 ( .A1(n12906), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17527) );
  INV_X1 U11824 ( .A(n10103), .ZN(n12906) );
  OAI211_X1 U11825 ( .C1(n17558), .C2(n17886), .A(n9823), .B(n17557), .ZN(
        n17541) );
  NOR2_X1 U11826 ( .A1(n17541), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17540) );
  NAND2_X1 U11827 ( .A1(n17662), .A2(n12900), .ZN(n17599) );
  NOR2_X1 U11828 ( .A1(n17692), .A2(n17994), .ZN(n17675) );
  INV_X1 U11829 ( .A(n13073), .ZN(n18073) );
  INV_X1 U11830 ( .A(n17943), .ZN(n18072) );
  INV_X1 U11831 ( .A(n17795), .ZN(n9922) );
  NAND2_X1 U11832 ( .A1(n17833), .A2(n12888), .ZN(n17815) );
  NAND2_X1 U11833 ( .A1(n9893), .A2(n9892), .ZN(n17813) );
  INV_X1 U11834 ( .A(n17816), .ZN(n9892) );
  INV_X1 U11835 ( .A(n17815), .ZN(n9893) );
  INV_X1 U11836 ( .A(n15639), .ZN(n18683) );
  INV_X1 U11837 ( .A(n18853), .ZN(n18213) );
  AND2_X1 U11838 ( .A1(n14198), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13758) );
  NAND2_X1 U11839 ( .A1(n9941), .A2(n20070), .ZN(n9940) );
  INV_X1 U11840 ( .A(n14588), .ZN(n9941) );
  XNOR2_X1 U11841 ( .A(n14196), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14589) );
  NAND2_X1 U11842 ( .A1(n10060), .A2(n10057), .ZN(n14196) );
  INV_X1 U11843 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20517) );
  OR2_X1 U11844 ( .A1(n11359), .A2(n13367), .ZN(n11361) );
  NAND2_X1 U11845 ( .A1(n9800), .A2(n11207), .ZN(n11208) );
  INV_X1 U11846 ( .A(n20094), .ZN(n13689) );
  INV_X1 U11847 ( .A(n12759), .ZN(n12760) );
  NAND2_X1 U11848 ( .A1(n10195), .A2(n15039), .ZN(n16072) );
  NAND2_X1 U11849 ( .A1(n16078), .A2(n16079), .ZN(n16077) );
  INV_X1 U11850 ( .A(n19846), .ZN(n19110) );
  XNOR2_X1 U11851 ( .A(n10155), .B(n10154), .ZN(n12777) );
  NAND2_X1 U11852 ( .A1(n10194), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10155) );
  XNOR2_X1 U11853 ( .A(n12729), .B(n12745), .ZN(n12782) );
  INV_X1 U11854 ( .A(n16187), .ZN(n19205) );
  AND2_X1 U11855 ( .A1(n16194), .A2(n19831), .ZN(n19201) );
  NAND2_X1 U11856 ( .A1(n12774), .A2(n19212), .ZN(n12748) );
  NAND2_X1 U11857 ( .A1(n15260), .A2(n19208), .ZN(n15269) );
  INV_X1 U11858 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19824) );
  NAND2_X1 U11859 ( .A1(n14102), .A2(n12379), .ZN(n12378) );
  OR2_X1 U11860 ( .A1(n19439), .A2(n19323), .ZN(n19366) );
  INV_X1 U11861 ( .A(n16824), .ZN(n16838) );
  NAND2_X1 U11862 ( .A1(n17595), .A2(n16303), .ZN(n17534) );
  AOI21_X1 U11863 ( .B1(n16314), .B2(n16316), .A(n21009), .ZN(n9884) );
  NAND2_X1 U11864 ( .A1(n10110), .A2(n10108), .ZN(n16334) );
  NAND2_X1 U11865 ( .A1(n15739), .A2(n10111), .ZN(n10110) );
  OAI21_X1 U11866 ( .B1(n12908), .B2(n12909), .A(n9844), .ZN(n10108) );
  AND2_X1 U11867 ( .A1(n12912), .A2(n12913), .ZN(n10111) );
  AND2_X1 U11868 ( .A1(n17890), .A2(n9927), .ZN(n9926) );
  AND2_X1 U11869 ( .A1(n17907), .A2(n9928), .ZN(n9927) );
  AND2_X1 U11870 ( .A1(n17891), .A2(n17889), .ZN(n9928) );
  INV_X1 U11871 ( .A(n18191), .ZN(n18185) );
  INV_X1 U11872 ( .A(n18198), .ZN(n18184) );
  INV_X1 U11873 ( .A(n12022), .ZN(n12023) );
  INV_X1 U11874 ( .A(n12517), .ZN(n10393) );
  NAND2_X1 U11875 ( .A1(n10759), .A2(n10745), .ZN(n10746) );
  NAND2_X1 U11876 ( .A1(n11728), .A2(n11727), .ZN(n11750) );
  INV_X1 U11877 ( .A(n11749), .ZN(n11728) );
  AND2_X1 U11878 ( .A1(n11750), .A2(n11729), .ZN(n11758) );
  OR2_X1 U11879 ( .A1(n11672), .A2(n11671), .ZN(n11678) );
  AND2_X1 U11880 ( .A1(n13995), .A2(n14029), .ZN(n10047) );
  AOI21_X1 U11881 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20486), .A(
        n11757), .ZN(n11767) );
  AOI21_X1 U11882 ( .B1(n14545), .B2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9879) );
  NOR2_X1 U11883 ( .A1(n11393), .A2(n9938), .ZN(n9937) );
  INV_X1 U11884 ( .A(n11385), .ZN(n9938) );
  OR2_X1 U11885 ( .A1(n11307), .A2(n11306), .ZN(n13805) );
  OR2_X1 U11886 ( .A1(n13748), .A2(n20639), .ZN(n11251) );
  NAND2_X1 U11887 ( .A1(n11163), .A2(n11162), .ZN(n13398) );
  AOI22_X1 U11888 ( .A1(n11252), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11070), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11109) );
  NOR2_X1 U11889 ( .A1(n14718), .A2(n20639), .ZN(n10032) );
  NAND2_X1 U11890 ( .A1(n11937), .A2(n11936), .ZN(n11940) );
  AOI22_X1 U11891 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n12008), .B1(
        n12009), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11912) );
  AOI22_X1 U11892 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12030), .B1(
        n21051), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11913) );
  AOI22_X1 U11893 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19433), .B1(
        n12007), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11923) );
  AOI22_X1 U11894 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19262), .B1(
        n12010), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11915) );
  AND4_X1 U11895 ( .A1(n10328), .A2(n10327), .A3(n10326), .A4(n10325), .ZN(
        n10331) );
  AOI22_X1 U11896 ( .A1(n10660), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9745), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10646) );
  AOI22_X1 U11897 ( .A1(n10660), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9745), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10651) );
  AND2_X1 U11898 ( .A1(n12215), .A2(n12707), .ZN(n10726) );
  AOI22_X1 U11899 ( .A1(n12550), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10252) );
  AOI22_X1 U11900 ( .A1(n10660), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n9745), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10634) );
  AOI22_X1 U11901 ( .A1(n12550), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10636) );
  AOI22_X1 U11902 ( .A1(n10660), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9744), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10639) );
  XNOR2_X1 U11903 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10677) );
  AOI21_X1 U11904 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18659), .A(
        n12925), .ZN(n12931) );
  NAND2_X1 U11905 ( .A1(n18820), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12794) );
  NOR2_X1 U11906 ( .A1(n13041), .A2(n17876), .ZN(n13047) );
  NOR2_X1 U11907 ( .A1(n13026), .A2(n15665), .ZN(n13030) );
  AND2_X1 U11908 ( .A1(n10035), .A2(n11688), .ZN(n10034) );
  NOR2_X1 U11909 ( .A1(n14313), .A2(n10036), .ZN(n10035) );
  INV_X1 U11910 ( .A(n14318), .ZN(n10036) );
  NOR2_X1 U11911 ( .A1(n20853), .A2(n11630), .ZN(n11631) );
  NAND2_X1 U11912 ( .A1(n11563), .A2(n10042), .ZN(n10041) );
  INV_X1 U11913 ( .A(n14357), .ZN(n10042) );
  INV_X1 U11914 ( .A(n14136), .ZN(n11559) );
  NOR2_X1 U11915 ( .A1(n14160), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10064) );
  INV_X1 U11916 ( .A(n14054), .ZN(n9950) );
  NAND2_X1 U11917 ( .A1(n13895), .A2(n13904), .ZN(n13952) );
  AND2_X1 U11918 ( .A1(n14191), .A2(n11786), .ZN(n11878) );
  AND2_X1 U11919 ( .A1(n13200), .A2(n13389), .ZN(n13373) );
  NAND2_X1 U11920 ( .A1(n11161), .A2(n13447), .ZN(n11176) );
  NOR2_X1 U11921 ( .A1(n14149), .A2(n20639), .ZN(n10056) );
  OR2_X1 U11922 ( .A1(n11268), .A2(n11267), .ZN(n13521) );
  INV_X1 U11923 ( .A(n11764), .ZN(n11770) );
  AND2_X1 U11924 ( .A1(n11158), .A2(n13201), .ZN(n13439) );
  NAND2_X1 U11925 ( .A1(n11114), .A2(n13360), .ZN(n10027) );
  OAI21_X1 U11926 ( .B1(n12209), .B2(n12194), .A(n12193), .ZN(n12195) );
  NAND2_X1 U11927 ( .A1(n10151), .A2(n12155), .ZN(n10714) );
  OR2_X1 U11928 ( .A1(n12160), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10151) );
  NAND2_X1 U11929 ( .A1(n12157), .A2(n14915), .ZN(n12160) );
  NAND2_X1 U11930 ( .A1(n9908), .A2(n9907), .ZN(n12078) );
  INV_X1 U11931 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n9907) );
  INV_X1 U11932 ( .A(n12070), .ZN(n9908) );
  NOR2_X1 U11933 ( .A1(n12065), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12067) );
  NAND2_X1 U11934 ( .A1(n9914), .A2(n9912), .ZN(n12065) );
  AND2_X1 U11935 ( .A1(n9771), .A2(n10148), .ZN(n9912) );
  NAND2_X1 U11936 ( .A1(n9909), .A2(n10701), .ZN(n11984) );
  NAND2_X1 U11937 ( .A1(n19237), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10701) );
  NAND2_X1 U11938 ( .A1(n12205), .A2(n12150), .ZN(n9909) );
  CLKBUF_X1 U11939 ( .A(n12550), .Z(n12689) );
  AOI21_X1 U11940 ( .B1(n14917), .B2(n14920), .A(n12587), .ZN(n12608) );
  INV_X1 U11941 ( .A(n14797), .ZN(n10078) );
  NOR2_X1 U11942 ( .A1(n14768), .A2(n9999), .ZN(n9998) );
  NOR2_X1 U11943 ( .A1(n15188), .A2(n9996), .ZN(n9995) );
  INV_X1 U11944 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n9996) );
  NOR2_X1 U11945 ( .A1(n20749), .A2(n10003), .ZN(n10002) );
  INV_X1 U11946 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10003) );
  INV_X1 U11947 ( .A(n10714), .ZN(n12768) );
  NAND2_X1 U11948 ( .A1(n12172), .A2(n10121), .ZN(n10120) );
  OR2_X1 U11949 ( .A1(n16106), .A2(n12158), .ZN(n12164) );
  NOR2_X1 U11950 ( .A1(n15092), .A2(n10098), .ZN(n10097) );
  AND2_X1 U11951 ( .A1(n14784), .A2(n12762), .ZN(n12127) );
  NOR2_X1 U11952 ( .A1(n14954), .A2(n10014), .ZN(n10013) );
  INV_X1 U11953 ( .A(n14002), .ZN(n10080) );
  AND2_X1 U11954 ( .A1(n12063), .A2(n12066), .ZN(n10124) );
  NAND2_X1 U11955 ( .A1(n12346), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12347) );
  NAND2_X1 U11956 ( .A1(n12325), .A2(n12158), .ZN(n12021) );
  AND3_X1 U11957 ( .A1(n10306), .A2(n10305), .A3(n10304), .ZN(n12313) );
  AND4_X1 U11958 ( .A1(n10299), .A2(n10298), .A3(n10297), .A4(n10296), .ZN(
        n10305) );
  AND4_X1 U11959 ( .A1(n10303), .A2(n10302), .A3(n10301), .A4(n10300), .ZN(
        n10304) );
  NAND2_X1 U11960 ( .A1(n10785), .A2(n10784), .ZN(n11904) );
  INV_X1 U11961 ( .A(n10783), .ZN(n10784) );
  NOR2_X1 U11962 ( .A1(n10280), .A2(n10279), .ZN(n12310) );
  NOR2_X1 U11963 ( .A1(n10244), .A2(n10245), .ZN(n12308) );
  NAND2_X1 U11964 ( .A1(n10215), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9853) );
  NAND2_X1 U11965 ( .A1(n10220), .A2(n10809), .ZN(n9854) );
  INV_X1 U11966 ( .A(n12201), .ZN(n10735) );
  NAND2_X1 U11967 ( .A1(n19834), .A2(n19680), .ZN(n13829) );
  AND2_X1 U11968 ( .A1(n12376), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11976) );
  NOR2_X1 U11969 ( .A1(n21023), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n12935) );
  NAND2_X1 U11970 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12956) );
  INV_X1 U11971 ( .A(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n20743) );
  INV_X1 U11972 ( .A(n12788), .ZN(n16909) );
  NOR2_X1 U11973 ( .A1(n12794), .A2(n18665), .ZN(n12994) );
  INV_X1 U11974 ( .A(n12841), .ZN(n10101) );
  NOR2_X1 U11975 ( .A1(n12793), .A2(n12789), .ZN(n16864) );
  NOR2_X1 U11976 ( .A1(n12794), .A2(n12789), .ZN(n12790) );
  NOR2_X1 U11977 ( .A1(n12792), .A2(n12794), .ZN(n12788) );
  NAND2_X1 U11978 ( .A1(n17542), .A2(n9779), .ZN(n13069) );
  NAND2_X1 U11979 ( .A1(n10139), .A2(n12903), .ZN(n12904) );
  NOR2_X1 U11980 ( .A1(n17555), .A2(n17885), .ZN(n17521) );
  INV_X1 U11981 ( .A(n17391), .ZN(n13041) );
  XNOR2_X1 U11982 ( .A(n17391), .B(n17383), .ZN(n12880) );
  XNOR2_X1 U11983 ( .A(n13047), .B(n13046), .ZN(n13048) );
  INV_X1 U11984 ( .A(n13031), .ZN(n15665) );
  NAND2_X1 U11985 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18812), .ZN(
        n12793) );
  NAND2_X1 U11986 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12791) );
  INV_X1 U11987 ( .A(n17185), .ZN(n14086) );
  NAND2_X1 U11988 ( .A1(n9953), .A2(n9842), .ZN(n14204) );
  NAND2_X1 U11989 ( .A1(n11889), .A2(n14250), .ZN(n9952) );
  AND2_X1 U11990 ( .A1(n11795), .A2(n11794), .ZN(n13551) );
  NAND2_X1 U11991 ( .A1(n11722), .A2(n9826), .ZN(n14153) );
  AND2_X1 U11992 ( .A1(n11722), .A2(n11721), .ZN(n14155) );
  AND2_X1 U11993 ( .A1(n14468), .A2(n14135), .ZN(n11706) );
  OR2_X1 U11994 ( .A1(n11698), .A2(n11697), .ZN(n14270) );
  OR2_X1 U11995 ( .A1(n15807), .A2(n11423), .ZN(n11657) );
  AND2_X1 U11996 ( .A1(n11615), .A2(n11614), .ZN(n14333) );
  AND2_X1 U11997 ( .A1(n11596), .A2(n11595), .ZN(n14341) );
  CLKBUF_X1 U11998 ( .A(n14331), .Z(n14332) );
  NOR2_X1 U11999 ( .A1(n11558), .A2(n15849), .ZN(n11578) );
  NAND2_X1 U12000 ( .A1(n11578), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11594) );
  NOR2_X1 U12001 ( .A1(n11513), .A2(n15870), .ZN(n11545) );
  NAND2_X1 U12002 ( .A1(n11497), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11513) );
  AND2_X1 U12003 ( .A1(n10044), .A2(n14052), .ZN(n10043) );
  AND2_X1 U12004 ( .A1(n11493), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n11497) );
  AND2_X1 U12005 ( .A1(n11438), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11455) );
  NOR2_X1 U12006 ( .A1(n11422), .A2(n13931), .ZN(n11438) );
  NAND2_X1 U12007 ( .A1(n11416), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11422) );
  AND2_X1 U12008 ( .A1(n11395), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11397) );
  INV_X1 U12009 ( .A(n13707), .ZN(n11401) );
  INV_X1 U12010 ( .A(n13693), .ZN(n11402) );
  NOR2_X1 U12011 ( .A1(n11387), .A2(n20884), .ZN(n11395) );
  CLKBUF_X1 U12012 ( .A(n13672), .Z(n13673) );
  AND2_X1 U12013 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n11085), .ZN(
        n11378) );
  INV_X1 U12014 ( .A(n13532), .ZN(n11366) );
  NOR2_X1 U12015 ( .A1(n10063), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10061) );
  INV_X1 U12016 ( .A(n10064), .ZN(n10063) );
  NOR2_X1 U12017 ( .A1(n10062), .A2(n10059), .ZN(n10058) );
  INV_X1 U12018 ( .A(n14174), .ZN(n10059) );
  NOR2_X1 U12019 ( .A1(n10064), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10062) );
  AND2_X1 U12020 ( .A1(n9953), .A2(n9951), .ZN(n14248) );
  NOR2_X1 U12021 ( .A1(n14266), .A2(n9954), .ZN(n9951) );
  NOR2_X1 U12022 ( .A1(n14272), .A2(n14266), .ZN(n14265) );
  OR2_X1 U12023 ( .A1(n9962), .A2(n14315), .ZN(n9960) );
  AND2_X1 U12024 ( .A1(n11850), .A2(n11849), .ZN(n15844) );
  NAND2_X1 U12025 ( .A1(n14347), .A2(n15844), .ZN(n15843) );
  NAND2_X1 U12026 ( .A1(n9936), .A2(n14166), .ZN(n14523) );
  NOR2_X1 U12027 ( .A1(n15935), .A2(n14171), .ZN(n14524) );
  NAND2_X1 U12028 ( .A1(n14080), .A2(n9776), .ZN(n14061) );
  NAND2_X1 U12029 ( .A1(n14080), .A2(n14079), .ZN(n14082) );
  AND2_X1 U12030 ( .A1(n14160), .A2(n16022), .ZN(n14550) );
  INV_X1 U12031 ( .A(n14012), .ZN(n9955) );
  NAND2_X1 U12032 ( .A1(n9956), .A2(n9957), .ZN(n14013) );
  NOR2_X1 U12033 ( .A1(n13866), .A2(n13865), .ZN(n13927) );
  NAND2_X1 U12034 ( .A1(n13551), .A2(n13550), .ZN(n13653) );
  NAND2_X1 U12035 ( .A1(n9948), .A2(n9947), .ZN(n13850) );
  INV_X1 U12036 ( .A(n13652), .ZN(n9947) );
  INV_X1 U12037 ( .A(n13653), .ZN(n9948) );
  OAI21_X1 U12038 ( .B1(n11351), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11248), 
        .ZN(n11348) );
  OAI21_X1 U12039 ( .B1(n11246), .B2(n20639), .A(n11245), .ZN(n11247) );
  INV_X1 U12040 ( .A(n11360), .ZN(n11279) );
  INV_X1 U12041 ( .A(n11197), .ZN(n9932) );
  AND2_X1 U12042 ( .A1(n13453), .A2(n13452), .ZN(n15699) );
  NOR2_X1 U12043 ( .A1(n20182), .A2(n20181), .ZN(n20406) );
  INV_X1 U12044 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20486) );
  INV_X1 U12045 ( .A(n20460), .ZN(n20464) );
  OR3_X1 U12046 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20104), .A3(n20492), 
        .ZN(n20149) );
  AND2_X1 U12047 ( .A1(n14146), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15727) );
  NAND2_X1 U12048 ( .A1(n9911), .A2(n9910), .ZN(n12205) );
  NAND2_X1 U12049 ( .A1(n12247), .A2(n12187), .ZN(n9910) );
  NAND2_X1 U12050 ( .A1(n12313), .A2(n12194), .ZN(n9911) );
  NAND2_X1 U12051 ( .A1(n12088), .A2(n14944), .ZN(n12134) );
  NAND2_X1 U12052 ( .A1(n19019), .A2(n10134), .ZN(n14752) );
  NAND2_X1 U12053 ( .A1(n14752), .A2(n15113), .ZN(n14751) );
  NOR2_X1 U12054 ( .A1(n13109), .A2(n13984), .ZN(n14003) );
  NAND2_X1 U12055 ( .A1(n10170), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10171) );
  NAND2_X1 U12056 ( .A1(n12102), .A2(n10709), .ZN(n12104) );
  INV_X1 U12057 ( .A(n12299), .ZN(n10019) );
  INV_X1 U12058 ( .A(n10904), .ZN(n14900) );
  NOR2_X1 U12059 ( .A1(n13633), .A2(n13632), .ZN(n12403) );
  AND2_X1 U12060 ( .A1(n10821), .A2(n10820), .ZN(n13514) );
  XNOR2_X1 U12061 ( .A(n12736), .B(n12735), .ZN(n16069) );
  NAND2_X1 U12062 ( .A1(n14985), .A2(n14986), .ZN(n14978) );
  NOR2_X1 U12063 ( .A1(n14905), .A2(n14904), .ZN(n14903) );
  NAND2_X1 U12064 ( .A1(n12516), .A2(n14948), .ZN(n10026) );
  NAND2_X1 U12065 ( .A1(n10079), .A2(n10076), .ZN(n15016) );
  NOR2_X1 U12066 ( .A1(n9817), .A2(n10077), .ZN(n10076) );
  INV_X1 U12067 ( .A(n13109), .ZN(n10079) );
  NAND2_X1 U12068 ( .A1(n10078), .A2(n15015), .ZN(n10077) );
  CLKBUF_X1 U12069 ( .A(n14945), .Z(n14946) );
  AND4_X1 U12070 ( .A1(n12418), .A2(n12417), .A3(n12416), .A4(n12415), .ZN(
        n13944) );
  AND3_X1 U12071 ( .A1(n10584), .A2(n10583), .A3(n10582), .ZN(n13108) );
  AND3_X1 U12072 ( .A1(n10565), .A2(n10564), .A3(n10563), .ZN(n15465) );
  NAND2_X1 U12073 ( .A1(n10434), .A2(n10433), .ZN(n15532) );
  AOI21_X1 U12074 ( .B1(n10073), .B2(n10412), .A(n10072), .ZN(n10071) );
  INV_X1 U12075 ( .A(n18880), .ZN(n13249) );
  INV_X1 U12076 ( .A(n10739), .ZN(n12706) );
  NAND2_X1 U12077 ( .A1(n10337), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10265) );
  OAI21_X1 U12078 ( .B1(n19869), .B2(n15557), .A(n10262), .ZN(n10263) );
  INV_X1 U12079 ( .A(n13225), .ZN(n13828) );
  NAND2_X1 U12080 ( .A1(n10187), .A2(n9787), .ZN(n10193) );
  NAND2_X1 U12081 ( .A1(n10187), .A2(n10004), .ZN(n10191) );
  NAND2_X1 U12082 ( .A1(n10187), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10189) );
  AND2_X1 U12083 ( .A1(n10185), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10187) );
  NAND2_X1 U12084 ( .A1(n10175), .A2(n9788), .ZN(n10183) );
  NOR2_X1 U12085 ( .A1(n10183), .A2(n10182), .ZN(n10185) );
  NAND2_X1 U12086 ( .A1(n10175), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10176) );
  NOR2_X1 U12087 ( .A1(n10173), .A2(n18918), .ZN(n10175) );
  NOR2_X1 U12088 ( .A1(n10171), .A2(n15156), .ZN(n10174) );
  NAND2_X1 U12089 ( .A1(n10174), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10173) );
  OAI21_X1 U12090 ( .B1(n9873), .B2(n9872), .A(n15152), .ZN(n15406) );
  INV_X1 U12091 ( .A(n15128), .ZN(n9872) );
  AND2_X1 U12092 ( .A1(n10168), .A2(n9994), .ZN(n10170) );
  AND2_X1 U12093 ( .A1(n9778), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9994) );
  NAND2_X1 U12094 ( .A1(n10168), .A2(n9778), .ZN(n10169) );
  NAND2_X1 U12095 ( .A1(n10168), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10167) );
  INV_X1 U12096 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n15188) );
  NAND2_X1 U12097 ( .A1(n10166), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10165) );
  NOR2_X1 U12098 ( .A1(n15211), .A2(n10165), .ZN(n10168) );
  NAND2_X1 U12099 ( .A1(n10000), .A2(n10001), .ZN(n10163) );
  AND2_X1 U12100 ( .A1(n9780), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10000) );
  NOR2_X1 U12101 ( .A1(n10163), .A2(n16179), .ZN(n10166) );
  AND2_X1 U12102 ( .A1(n13419), .A2(n10010), .ZN(n13512) );
  AND2_X1 U12103 ( .A1(n10001), .A2(n9780), .ZN(n10164) );
  NAND2_X1 U12104 ( .A1(n10001), .A2(n10002), .ZN(n10161) );
  NOR2_X1 U12105 ( .A1(n10159), .A2(n20749), .ZN(n10162) );
  NAND2_X1 U12106 ( .A1(n13419), .A2(n13485), .ZN(n13513) );
  INV_X1 U12107 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13767) );
  NOR2_X1 U12108 ( .A1(n10158), .A2(n13767), .ZN(n10160) );
  NAND2_X1 U12109 ( .A1(n10115), .A2(n10114), .ZN(n15033) );
  AOI21_X1 U12110 ( .B1(n10118), .B2(n10117), .A(n10116), .ZN(n10115) );
  NAND2_X1 U12111 ( .A1(n12169), .A2(n10117), .ZN(n10114) );
  INV_X1 U12112 ( .A(n15045), .ZN(n10116) );
  NOR2_X1 U12113 ( .A1(n12158), .A2(n15261), .ZN(n9918) );
  AND2_X1 U12114 ( .A1(n12350), .A2(n9850), .ZN(n10096) );
  OAI21_X1 U12115 ( .B1(n12761), .B2(n12158), .A(n15277), .ZN(n15045) );
  NOR2_X1 U12116 ( .A1(n10119), .A2(n15278), .ZN(n10118) );
  AND2_X1 U12117 ( .A1(n9783), .A2(n14913), .ZN(n10015) );
  NAND2_X1 U12118 ( .A1(n12149), .A2(n9968), .ZN(n9967) );
  NOR2_X1 U12119 ( .A1(n15089), .A2(n15092), .ZN(n10127) );
  OR2_X1 U12120 ( .A1(n10126), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9965) );
  INV_X1 U12121 ( .A(n15089), .ZN(n10126) );
  NAND2_X1 U12122 ( .A1(n9794), .A2(n12762), .ZN(n15089) );
  NAND2_X1 U12123 ( .A1(n14760), .A2(n10017), .ZN(n14923) );
  OR2_X1 U12124 ( .A1(n15394), .A2(n12268), .ZN(n15363) );
  INV_X1 U12125 ( .A(n14764), .ZN(n14782) );
  NAND2_X1 U12126 ( .A1(n14795), .A2(n10013), .ZN(n14955) );
  NOR3_X1 U12127 ( .A1(n13109), .A2(n9817), .A3(n14797), .ZN(n15014) );
  NAND2_X1 U12128 ( .A1(n10007), .A2(n13724), .ZN(n10006) );
  INV_X1 U12129 ( .A(n10008), .ZN(n10007) );
  NAND2_X1 U12130 ( .A1(n10112), .A2(n9972), .ZN(n9971) );
  INV_X1 U12131 ( .A(n9795), .ZN(n9972) );
  NAND2_X1 U12132 ( .A1(n15204), .A2(n15207), .ZN(n15120) );
  NOR2_X1 U12133 ( .A1(n13676), .A2(n10008), .ZN(n13725) );
  INV_X1 U12134 ( .A(n15469), .ZN(n15498) );
  AND3_X1 U12135 ( .A1(n10493), .A2(n10492), .A3(n10491), .ZN(n14814) );
  OR2_X1 U12136 ( .A1(n14824), .A2(n10086), .ZN(n15514) );
  AND2_X1 U12137 ( .A1(n12077), .A2(n16207), .ZN(n15220) );
  INV_X1 U12138 ( .A(n13539), .ZN(n10832) );
  INV_X1 U12139 ( .A(n13540), .ZN(n10833) );
  AND3_X1 U12140 ( .A1(n10458), .A2(n10457), .A3(n10456), .ZN(n14826) );
  NAND2_X1 U12141 ( .A1(n9852), .A2(n11995), .ZN(n13969) );
  AND3_X1 U12142 ( .A1(n10361), .A2(n10360), .A3(n10359), .ZN(n14832) );
  NAND2_X1 U12143 ( .A1(n13761), .A2(n13763), .ZN(n9969) );
  OR2_X1 U12144 ( .A1(n12352), .A2(n15582), .ZN(n12274) );
  NAND2_X1 U12145 ( .A1(n9863), .A2(n19869), .ZN(n9862) );
  NAND2_X1 U12146 ( .A1(n12370), .A2(n19385), .ZN(n12394) );
  AND2_X2 U12147 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n15580) );
  OR2_X1 U12148 ( .A1(n14104), .A2(n12383), .ZN(n12384) );
  AND2_X1 U12149 ( .A1(n14097), .A2(n14096), .ZN(n16242) );
  INV_X1 U12150 ( .A(n19296), .ZN(n19357) );
  INV_X1 U12151 ( .A(n19494), .ZN(n19497) );
  AND2_X1 U12152 ( .A1(n19825), .A2(n15608), .ZN(n19547) );
  INV_X1 U12153 ( .A(n19252), .ZN(n19242) );
  NOR2_X2 U12154 ( .A1(n13828), .A2(n13829), .ZN(n19251) );
  NOR2_X2 U12155 ( .A1(n13830), .A2(n13829), .ZN(n19252) );
  INV_X1 U12156 ( .A(n10630), .ZN(n19254) );
  INV_X1 U12157 ( .A(n16242), .ZN(n16281) );
  INV_X1 U12158 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16280) );
  NAND2_X1 U12159 ( .A1(n17448), .A2(n18213), .ZN(n13029) );
  OR2_X1 U12160 ( .A1(n13027), .A2(n18221), .ZN(n16430) );
  INV_X1 U12161 ( .A(n18867), .ZN(n18856) );
  OAI22_X1 U12162 ( .A1(n18679), .A2(n18688), .B1(n15639), .B2(n18684), .ZN(
        n18689) );
  AND2_X1 U12163 ( .A1(n16531), .A2(n16469), .ZN(n16518) );
  OR2_X1 U12164 ( .A1(n16587), .A2(n17613), .ZN(n16585) );
  NOR2_X1 U12165 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16720), .ZN(n16708) );
  NOR2_X1 U12166 ( .A1(n17446), .A2(n17445), .ZN(n17447) );
  NAND2_X1 U12167 ( .A1(n17542), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17511) );
  NAND2_X1 U12168 ( .A1(n17585), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17561) );
  NOR2_X1 U12169 ( .A1(n17640), .A2(n17641), .ZN(n17629) );
  NAND2_X1 U12170 ( .A1(n17661), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17640) );
  AND2_X1 U12171 ( .A1(n9988), .A2(n17777), .ZN(n16467) );
  AOI21_X1 U12172 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n13068), .A(
        n18593), .ZN(n17714) );
  NAND2_X1 U12173 ( .A1(n17777), .A2(n16672), .ZN(n17713) );
  NAND2_X1 U12174 ( .A1(n13064), .A2(n17774), .ZN(n16302) );
  INV_X1 U12175 ( .A(n13062), .ZN(n13060) );
  NAND2_X1 U12176 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17828) );
  NOR2_X1 U12177 ( .A1(n21009), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n10109) );
  NOR2_X1 U12178 ( .A1(n10102), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10129) );
  OR2_X1 U12179 ( .A1(n17566), .A2(n17782), .ZN(n17557) );
  NOR2_X1 U12180 ( .A1(n18023), .A2(n17575), .ZN(n17926) );
  OR2_X1 U12181 ( .A1(n18107), .A2(n17448), .ZN(n18684) );
  NAND2_X1 U12182 ( .A1(n12901), .A2(n10130), .ZN(n12902) );
  AND2_X1 U12183 ( .A1(n17674), .A2(n9803), .ZN(n9895) );
  AND2_X1 U12184 ( .A1(n17721), .A2(n9929), .ZN(n17705) );
  NOR2_X1 U12185 ( .A1(n20828), .A2(n18034), .ZN(n9929) );
  INV_X1 U12186 ( .A(n17721), .ZN(n18047) );
  INV_X1 U12187 ( .A(n16302), .ZN(n18070) );
  AND2_X1 U12188 ( .A1(n12896), .A2(n9900), .ZN(n9899) );
  AOI21_X1 U12189 ( .B1(n12896), .B2(n18106), .A(n9900), .ZN(n9897) );
  NAND2_X1 U12190 ( .A1(n18114), .A2(n17782), .ZN(n17781) );
  NAND2_X1 U12191 ( .A1(n13061), .A2(n9924), .ZN(n17775) );
  AOI21_X1 U12192 ( .B1(n9921), .B2(n9828), .A(n9770), .ZN(n9924) );
  XNOR2_X1 U12193 ( .A(n13057), .B(n9919), .ZN(n17805) );
  INV_X1 U12194 ( .A(n13058), .ZN(n9919) );
  NAND2_X1 U12195 ( .A1(n17830), .A2(n13055), .ZN(n17820) );
  NOR2_X1 U12196 ( .A1(n17820), .A2(n17821), .ZN(n17819) );
  NAND2_X1 U12197 ( .A1(n17846), .A2(n12885), .ZN(n17834) );
  XNOR2_X1 U12198 ( .A(n9894), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17835) );
  INV_X1 U12199 ( .A(n12887), .ZN(n9894) );
  NAND2_X1 U12200 ( .A1(n17834), .A2(n17835), .ZN(n17833) );
  INV_X1 U12201 ( .A(n18685), .ZN(n18145) );
  XNOR2_X1 U12202 ( .A(n12880), .B(n12866), .ZN(n17859) );
  XNOR2_X1 U12203 ( .A(n13048), .B(n12866), .ZN(n17856) );
  NAND2_X1 U12204 ( .A1(n17855), .A2(n17856), .ZN(n17854) );
  NOR2_X1 U12205 ( .A1(n13027), .A2(n13032), .ZN(n15660) );
  NOR2_X1 U12206 ( .A1(n13028), .A2(n15640), .ZN(n9890) );
  INV_X1 U12207 ( .A(n13025), .ZN(n13028) );
  NAND2_X1 U12208 ( .A1(n18856), .A2(n15674), .ZN(n18685) );
  OR2_X1 U12209 ( .A1(n18827), .A2(n12791), .ZN(n15676) );
  NOR2_X1 U12210 ( .A1(n12950), .A2(n12949), .ZN(n18225) );
  NOR2_X1 U12211 ( .A1(n12981), .A2(n12980), .ZN(n18238) );
  INV_X1 U12212 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n20757) );
  INV_X1 U12213 ( .A(n20716), .ZN(n13734) );
  NAND2_X1 U12214 ( .A1(n13567), .A2(n13181), .ZN(n20716) );
  OR2_X1 U12215 ( .A1(n13755), .A2(n13754), .ZN(n19969) );
  INV_X1 U12216 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15849) );
  INV_X1 U12217 ( .A(n19986), .ZN(n19971) );
  INV_X1 U12218 ( .A(n19959), .ZN(n19987) );
  INV_X1 U12219 ( .A(n19953), .ZN(n19925) );
  OR2_X1 U12220 ( .A1(n19932), .A2(n13744), .ZN(n19996) );
  INV_X1 U12221 ( .A(n19927), .ZN(n19967) );
  AND2_X1 U12222 ( .A1(n19927), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19991) );
  CLKBUF_X1 U12223 ( .A(n14141), .Z(n14422) );
  INV_X1 U12224 ( .A(n14411), .ZN(n14421) );
  INV_X1 U12225 ( .A(n14429), .ZN(n14075) );
  AND2_X1 U12226 ( .A1(n13305), .A2(n15723), .ZN(n20023) );
  INV_X2 U12227 ( .A(n20017), .ZN(n20033) );
  XNOR2_X1 U12228 ( .A(n13742), .B(n13741), .ZN(n14198) );
  OR2_X1 U12229 ( .A1(n14110), .A2(n14181), .ZN(n13742) );
  INV_X1 U12230 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15831) );
  INV_X1 U12231 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15870) );
  AND2_X1 U12232 ( .A1(n14078), .A2(n14069), .ZN(n15958) );
  INV_X1 U12233 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20884) );
  NAND2_X1 U12234 ( .A1(n15962), .A2(n13501), .ZN(n15984) );
  AND2_X1 U12235 ( .A1(n15984), .A2(n20059), .ZN(n15979) );
  INV_X1 U12236 ( .A(n15984), .ZN(n20060) );
  XNOR2_X1 U12237 ( .A(n9881), .B(n14591), .ZN(n14590) );
  NAND2_X1 U12238 ( .A1(n10065), .A2(n10066), .ZN(n9881) );
  NAND2_X1 U12239 ( .A1(n14180), .A2(n14179), .ZN(n10066) );
  OR2_X1 U12240 ( .A1(n15985), .A2(n14570), .ZN(n14653) );
  NAND2_X1 U12241 ( .A1(n13949), .A2(n13948), .ZN(n14015) );
  NAND2_X1 U12242 ( .A1(n13903), .A2(n15972), .ZN(n13913) );
  INV_X1 U12243 ( .A(n13656), .ZN(n14577) );
  OR2_X1 U12244 ( .A1(n13409), .A2(n13404), .ZN(n14580) );
  OR2_X1 U12245 ( .A1(n13500), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20066) );
  NOR2_X1 U12246 ( .A1(n13408), .A2(n13406), .ZN(n20085) );
  INV_X1 U12247 ( .A(n20547), .ZN(n20581) );
  INV_X1 U12248 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20487) );
  OAI21_X1 U12249 ( .B1(n20097), .B2(n9804), .A(n11377), .ZN(n20096) );
  AND2_X1 U12250 ( .A1(n13597), .A2(n20249), .ZN(n20094) );
  NOR2_X1 U12251 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19883) );
  INV_X1 U12252 ( .A(n20222), .ZN(n20239) );
  INV_X1 U12253 ( .A(n20271), .ZN(n20238) );
  OAI21_X1 U12254 ( .B1(n20265), .B2(n20250), .A(n20556), .ZN(n20268) );
  INV_X1 U12255 ( .A(n20297), .ZN(n20267) );
  AND2_X1 U12256 ( .A1(n20328), .A2(n20406), .ZN(n20345) );
  OAI211_X1 U12257 ( .C1(n20371), .C2(n20492), .A(n20421), .B(n20356), .ZN(
        n20373) );
  INV_X1 U12258 ( .A(n20405), .ZN(n20384) );
  INV_X1 U12259 ( .A(n20516), .ZN(n20477) );
  INV_X1 U12260 ( .A(n20578), .ZN(n20536) );
  INV_X1 U12261 ( .A(n20539), .ZN(n20543) );
  NOR2_X1 U12262 ( .A1(n20517), .A2(n20580), .ZN(n20630) );
  AND2_X1 U12263 ( .A1(n20098), .A2(n20463), .ZN(n20634) );
  NOR2_X1 U12264 ( .A1(n13436), .A2(n20492), .ZN(n15731) );
  INV_X1 U12265 ( .A(n20715), .ZN(n20727) );
  AND2_X1 U12266 ( .A1(n10688), .A2(n16273), .ZN(n13134) );
  NAND2_X1 U12267 ( .A1(n16088), .A2(n16089), .ZN(n16087) );
  NAND2_X1 U12268 ( .A1(n16100), .A2(n16101), .ZN(n16099) );
  NAND2_X1 U12269 ( .A1(n16112), .A2(n16113), .ZN(n16111) );
  NAND2_X1 U12270 ( .A1(n16126), .A2(n16127), .ZN(n16125) );
  NAND2_X1 U12271 ( .A1(n16135), .A2(n16136), .ZN(n16134) );
  NAND2_X1 U12272 ( .A1(n14751), .A2(n19019), .ZN(n14732) );
  NAND2_X1 U12273 ( .A1(n14732), .A2(n15103), .ZN(n14731) );
  INV_X1 U12274 ( .A(n19014), .ZN(n19035) );
  AND2_X1 U12275 ( .A1(n12116), .A2(n12115), .ZN(n14790) );
  INV_X1 U12276 ( .A(n19019), .ZN(n19005) );
  INV_X1 U12277 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n15211) );
  NOR2_X1 U12278 ( .A1(n12020), .A2(n12019), .ZN(n12050) );
  INV_X1 U12279 ( .A(n19028), .ZN(n18999) );
  NAND2_X1 U12280 ( .A1(n9870), .A2(n9871), .ZN(n9869) );
  AND2_X1 U12281 ( .A1(n11895), .A2(n10799), .ZN(n9870) );
  OAI21_X1 U12282 ( .B1(n12300), .B2(n14882), .A(n14881), .ZN(n15275) );
  AND2_X1 U12283 ( .A1(n10025), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10024) );
  INV_X1 U12284 ( .A(n14966), .ZN(n14941) );
  OR2_X1 U12285 ( .A1(n13257), .A2(n19254), .ZN(n14966) );
  OAI21_X1 U12286 ( .B1(n14878), .B2(n14879), .A(n10133), .ZN(n12701) );
  XNOR2_X1 U12287 ( .A(n14878), .B(n14879), .ZN(n14973) );
  AND2_X1 U12288 ( .A1(n14940), .A2(n14939), .ZN(n16150) );
  NOR2_X1 U12289 ( .A1(n13339), .A2(n13830), .ZN(n19049) );
  NOR2_X1 U12290 ( .A1(n13339), .A2(n13828), .ZN(n19047) );
  NAND2_X1 U12291 ( .A1(n19072), .A2(n12708), .ZN(n16141) );
  OAI21_X1 U12292 ( .B1(n13775), .B2(n10073), .A(n10412), .ZN(n15544) );
  NOR2_X1 U12293 ( .A1(n19107), .A2(n19106), .ZN(n19086) );
  AND2_X1 U12294 ( .A1(n19072), .A2(n19254), .ZN(n19106) );
  INV_X1 U12295 ( .A(n13146), .ZN(n19187) );
  INV_X1 U12296 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16179) );
  INV_X1 U12297 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n20749) );
  INV_X1 U12298 ( .A(n13777), .ZN(n13478) );
  INV_X1 U12299 ( .A(n19197), .ZN(n16188) );
  INV_X1 U12300 ( .A(n16194), .ZN(n19190) );
  INV_X1 U12301 ( .A(n19201), .ZN(n16186) );
  INV_X1 U12302 ( .A(n9873), .ZN(n15150) );
  AND2_X1 U12303 ( .A1(n12278), .A2(n12277), .ZN(n16217) );
  AND2_X1 U12304 ( .A1(n10093), .A2(n10092), .ZN(n15252) );
  OR2_X1 U12305 ( .A1(n12352), .A2(n12293), .ZN(n16197) );
  OR2_X1 U12306 ( .A1(n12352), .A2(n12264), .ZN(n15425) );
  INV_X1 U12307 ( .A(n16197), .ZN(n19208) );
  INV_X1 U12308 ( .A(n15556), .ZN(n15426) );
  OR2_X1 U12309 ( .A1(n14104), .A2(n13248), .ZN(n19846) );
  INV_X1 U12310 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15764) );
  AND2_X1 U12311 ( .A1(n13256), .A2(n13255), .ZN(n19838) );
  NAND2_X1 U12312 ( .A1(n13827), .A2(n13826), .ZN(n19258) );
  OR2_X1 U12313 ( .A1(n13836), .A2(n13833), .ZN(n13827) );
  OAI21_X1 U12314 ( .B1(n13836), .B2(n13835), .A(n13834), .ZN(n19257) );
  OAI21_X1 U12315 ( .B1(n19363), .B2(n19362), .A(n19361), .ZN(n19382) );
  INV_X1 U12316 ( .A(n19560), .ZN(n19577) );
  INV_X1 U12317 ( .A(n19697), .ZN(n19581) );
  INV_X1 U12318 ( .A(n19630), .ZN(n19623) );
  INV_X1 U12319 ( .A(n19691), .ZN(n19646) );
  OAI22_X1 U12320 ( .A1(n20810), .A2(n19243), .B1(n19227), .B2(n19242), .ZN(
        n19653) );
  OAI21_X1 U12321 ( .B1(n19642), .B2(n19641), .A(n19640), .ZN(n19666) );
  INV_X1 U12322 ( .A(n19645), .ZN(n19682) );
  INV_X1 U12323 ( .A(n19270), .ZN(n19686) );
  INV_X1 U12324 ( .A(n19567), .ZN(n19711) );
  NOR2_X1 U12325 ( .A1(n19631), .A2(n19815), .ZN(n19718) );
  OAI22_X1 U12326 ( .A1(n19244), .A2(n19243), .B1(n20790), .B2(n19242), .ZN(
        n19717) );
  AND2_X1 U12327 ( .A1(n12391), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19724) );
  OR2_X1 U12328 ( .A1(n19741), .A2(n10692), .ZN(n18880) );
  OR2_X1 U12329 ( .A1(n16290), .A2(n16289), .ZN(n16291) );
  INV_X1 U12330 ( .A(n9985), .ZN(n16487) );
  INV_X1 U12331 ( .A(n9984), .ZN(n16497) );
  AND2_X1 U12332 ( .A1(n9984), .A2(n9983), .ZN(n16496) );
  INV_X1 U12333 ( .A(n9980), .ZN(n16533) );
  NOR2_X1 U12334 ( .A1(n16542), .A2(n17554), .ZN(n16541) );
  INV_X1 U12335 ( .A(n16807), .ZN(n16825) );
  AND2_X1 U12336 ( .A1(n9992), .A2(n16469), .ZN(n16563) );
  NOR2_X1 U12337 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16588), .ZN(n16574) );
  OAI21_X1 U12338 ( .B1(n17603), .B2(n16820), .A(n16645), .ZN(n16597) );
  NOR2_X1 U12339 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16772), .ZN(n16756) );
  NOR2_X2 U12340 ( .A1(n18808), .A2(n16834), .ZN(n16821) );
  AND2_X1 U12341 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n17026), .ZN(n17013) );
  NOR4_X2 U12342 ( .A1(n18217), .A2(n18213), .A3(n15766), .A4(n18708), .ZN(
        n17235) );
  INV_X1 U12343 ( .A(n17235), .ZN(n17237) );
  INV_X1 U12344 ( .A(n17258), .ZN(n17255) );
  NAND2_X1 U12345 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17272), .ZN(n17267) );
  NAND2_X1 U12346 ( .A1(n17318), .A2(n17244), .ZN(n17283) );
  NOR2_X1 U12347 ( .A1(n17389), .A2(n18238), .ZN(n17316) );
  NOR2_X1 U12348 ( .A1(n17329), .A2(n17504), .ZN(n17325) );
  AOI211_X1 U12349 ( .C1(n17184), .C2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n13000), .B(n12999), .ZN(n13001) );
  NAND2_X1 U12350 ( .A1(n17242), .A2(n17365), .ZN(n17355) );
  INV_X1 U12351 ( .A(n17389), .ZN(n17354) );
  NOR2_X1 U12352 ( .A1(n12810), .A2(n12809), .ZN(n17372) );
  INV_X1 U12353 ( .A(n17392), .ZN(n17384) );
  NAND2_X1 U12354 ( .A1(n15769), .A2(n17354), .ZN(n17387) );
  OAI21_X1 U12355 ( .B1(n15768), .B2(n15767), .A(n18849), .ZN(n17388) );
  INV_X1 U12356 ( .A(n17387), .ZN(n17393) );
  NOR2_X1 U12357 ( .A1(n17445), .A2(n17397), .ZN(n17443) );
  OAI21_X1 U12358 ( .B1(n18217), .B2(n18854), .A(n17447), .ZN(n17505) );
  NAND2_X1 U12359 ( .A1(n18217), .A2(n17447), .ZN(n17508) );
  NOR2_X1 U12360 ( .A1(n17606), .A2(n17607), .ZN(n17585) );
  NOR2_X1 U12361 ( .A1(n17773), .A2(n17994), .ZN(n17658) );
  AND3_X1 U12362 ( .A1(n9988), .A2(n9986), .A3(n17777), .ZN(n17661) );
  NOR2_X1 U12363 ( .A1(n17680), .A2(n9987), .ZN(n9986) );
  NOR2_X1 U12364 ( .A1(n13073), .A2(n17994), .ZN(n17940) );
  AND2_X1 U12365 ( .A1(n9887), .A2(n9886), .ZN(n17773) );
  NAND2_X1 U12366 ( .A1(n17869), .A2(n16302), .ZN(n9886) );
  NAND2_X1 U12367 ( .A1(n17784), .A2(n18073), .ZN(n9887) );
  INV_X1 U12368 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17811) );
  NOR2_X1 U12369 ( .A1(n18217), .A2(n16439), .ZN(n17818) );
  NOR2_X1 U12370 ( .A1(n17828), .A2(n17841), .ZN(n17812) );
  INV_X1 U12371 ( .A(n18454), .ZN(n18593) );
  NAND2_X1 U12372 ( .A1(n17877), .A2(n17845), .ZN(n17872) );
  NAND2_X1 U12373 ( .A1(n17665), .A2(n9718), .ZN(n17871) );
  INV_X1 U12374 ( .A(n17869), .ZN(n17881) );
  OAI21_X1 U12375 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18848), .A(n16439), 
        .ZN(n17877) );
  INV_X1 U12376 ( .A(n17818), .ZN(n17880) );
  OAI21_X1 U12377 ( .B1(n17515), .B2(n16345), .A(n16344), .ZN(n9904) );
  AND2_X1 U12378 ( .A1(n16343), .A2(n16342), .ZN(n16344) );
  OR2_X1 U12379 ( .A1(n16338), .A2(n10131), .ZN(n16345) );
  NAND2_X1 U12380 ( .A1(n9774), .A2(n9848), .ZN(n9902) );
  AND2_X1 U12381 ( .A1(n9926), .A2(n9925), .ZN(n17893) );
  AOI21_X1 U12382 ( .B1(n18647), .B2(n17899), .A(n17892), .ZN(n9925) );
  NAND2_X1 U12383 ( .A1(n18094), .A2(n18052), .ZN(n18107) );
  NAND2_X1 U12384 ( .A1(n17705), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18023) );
  INV_X1 U12385 ( .A(n9921), .ZN(n17793) );
  NOR2_X2 U12386 ( .A1(n15660), .A2(n13034), .ZN(n18656) );
  INV_X1 U12387 ( .A(n15659), .ZN(n13034) );
  INV_X1 U12388 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18207) );
  AOI211_X1 U12389 ( .C1(n18849), .C2(n18677), .A(n18212), .B(n15675), .ZN(
        n18832) );
  INV_X1 U12390 ( .A(n18832), .ZN(n18830) );
  INV_X1 U12391 ( .A(n16823), .ZN(n18717) );
  INV_X1 U12392 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18808) );
  INV_X1 U12393 ( .A(n18793), .ZN(n18863) );
  NAND2_X1 U12395 ( .A1(n9942), .A2(n9939), .ZN(P1_U3000) );
  NAND2_X1 U12396 ( .A1(n10917), .A2(n10916), .ZN(n10918) );
  AOI21_X1 U12397 ( .B1(n12774), .B2(n19201), .A(n12778), .ZN(n12781) );
  NOR2_X1 U12398 ( .A1(n12305), .A2(n12304), .ZN(n12355) );
  AND2_X1 U12399 ( .A1(n16086), .A2(n19212), .ZN(n12304) );
  OR2_X1 U12400 ( .A1(n16502), .A2(P3_EBX_REG_30__SCAN_IN), .ZN(n9978) );
  INV_X1 U12401 ( .A(n13081), .ZN(n13082) );
  AOI21_X1 U12402 ( .B1(n16333), .B2(n17869), .A(n13080), .ZN(n13081) );
  OR3_X1 U12403 ( .A1(n17534), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n16304), .ZN(n9883) );
  NAND2_X1 U12404 ( .A1(n16310), .A2(n17783), .ZN(n9885) );
  NAND2_X1 U12405 ( .A1(n10107), .A2(n10105), .ZN(P3_U2831) );
  AOI21_X1 U12406 ( .B1(n16333), .B2(n18184), .A(n10106), .ZN(n10105) );
  OAI21_X1 U12407 ( .B1(n16336), .B2(n18044), .A(n16335), .ZN(n10106) );
  NAND2_X1 U12408 ( .A1(n9905), .A2(n9901), .ZN(P3_U2834) );
  AOI21_X1 U12409 ( .B1(n9904), .B2(n9903), .A(n9902), .ZN(n9901) );
  NAND2_X1 U12410 ( .A1(n16350), .A2(n12905), .ZN(n9905) );
  NOR2_X1 U12411 ( .A1(n9726), .A2(n12905), .ZN(n9903) );
  AND2_X1 U12412 ( .A1(n9926), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17900) );
  AND2_X1 U12413 ( .A1(n12842), .A2(n10101), .ZN(n9764) );
  NAND4_X1 U12414 ( .A1(n10742), .A2(n19254), .A3(n10741), .A4(n10721), .ZN(
        n10759) );
  AND4_X1 U12415 ( .A1(n12840), .A2(n12839), .A3(n12838), .A4(n12837), .ZN(
        n9765) );
  INV_X1 U12416 ( .A(n10039), .ZN(n14345) );
  NAND2_X2 U12417 ( .A1(n10210), .A2(n10209), .ZN(n11932) );
  INV_X2 U12418 ( .A(n11932), .ZN(n19869) );
  NAND2_X1 U12419 ( .A1(n9732), .A2(n9777), .ZN(n13683) );
  AND3_X1 U12420 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9766) );
  OR2_X1 U12421 ( .A1(n12792), .A2(n12793), .ZN(n9767) );
  NOR2_X1 U12422 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n15676), .ZN(
        n12836) );
  NAND2_X1 U12423 ( .A1(n15928), .A2(n15927), .ZN(n14508) );
  NAND2_X1 U12424 ( .A1(n14317), .A2(n14318), .ZN(n14311) );
  INV_X1 U12425 ( .A(n13748), .ZN(n11249) );
  NAND2_X1 U12426 ( .A1(n15159), .A2(n12348), .ZN(n15392) );
  NAND2_X1 U12427 ( .A1(n9739), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15091) );
  NAND2_X1 U12428 ( .A1(n10020), .A2(n13856), .ZN(n13855) );
  AND4_X1 U12429 ( .A1(n12015), .A2(n12014), .A3(n12013), .A4(n12012), .ZN(
        n9768) );
  INV_X1 U12430 ( .A(n11957), .ZN(n11999) );
  NOR2_X1 U12431 ( .A1(n14978), .A2(n9840), .ZN(n9769) );
  AND2_X1 U12432 ( .A1(n17795), .A2(n17794), .ZN(n9770) );
  AND2_X1 U12433 ( .A1(n9915), .A2(n9913), .ZN(n9771) );
  OR3_X1 U12434 ( .A1(n14334), .A2(n9962), .A3(n14326), .ZN(n9772) );
  NOR2_X1 U12435 ( .A1(n14058), .A2(n10041), .ZN(n10039) );
  AND2_X1 U12436 ( .A1(n9816), .A2(n14501), .ZN(n9773) );
  AND2_X1 U12437 ( .A1(n9864), .A2(n9814), .ZN(n10769) );
  NAND3_X1 U12438 ( .A1(n17526), .A2(n9717), .A3(n17516), .ZN(n9774) );
  NAND2_X1 U12439 ( .A1(n9732), .A2(n12403), .ZN(n13634) );
  NAND2_X1 U12440 ( .A1(n13417), .A2(n13416), .ZN(n13415) );
  NOR2_X1 U12441 ( .A1(n13775), .A2(n14832), .ZN(n9775) );
  AND2_X1 U12442 ( .A1(n14079), .A2(n9950), .ZN(n9776) );
  AND2_X1 U12443 ( .A1(n12403), .A2(n9831), .ZN(n9777) );
  AND2_X1 U12444 ( .A1(n9995), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9778) );
  AND2_X1 U12445 ( .A1(n9766), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9779) );
  AND2_X1 U12446 ( .A1(n10002), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9780) );
  AND2_X1 U12447 ( .A1(n10013), .A2(n10012), .ZN(n9781) );
  OR2_X1 U12448 ( .A1(n13676), .A2(n13122), .ZN(n9782) );
  AND2_X1 U12449 ( .A1(n10017), .A2(n10016), .ZN(n9783) );
  AND2_X1 U12450 ( .A1(n9776), .A2(n9830), .ZN(n9784) );
  AND2_X1 U12451 ( .A1(n9777), .A2(n9829), .ZN(n9785) );
  INV_X1 U12452 ( .A(n15520), .ZN(n19212) );
  INV_X1 U12453 ( .A(n9863), .ZN(n10722) );
  AND2_X1 U12454 ( .A1(n9998), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9786) );
  AND2_X1 U12455 ( .A1(n10004), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9787) );
  AND2_X1 U12456 ( .A1(n9786), .A2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9788) );
  AND2_X1 U12457 ( .A1(n12348), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n9789) );
  AND2_X1 U12458 ( .A1(n9789), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9790) );
  AND2_X1 U12459 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n14444), .ZN(
        n9791) );
  OR2_X1 U12460 ( .A1(n14735), .A2(n15326), .ZN(n9792) );
  NAND2_X1 U12461 ( .A1(n14558), .A2(n14159), .ZN(n14522) );
  AND2_X1 U12462 ( .A1(n12550), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12465) );
  AND4_X1 U12463 ( .A1(n11140), .A2(n11139), .A3(n11138), .A4(n11137), .ZN(
        n9793) );
  OR2_X1 U12464 ( .A1(n12233), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10570) );
  INV_X1 U12465 ( .A(n10104), .ZN(n12898) );
  NAND2_X1 U12466 ( .A1(n17787), .A2(n9899), .ZN(n10104) );
  INV_X1 U12467 ( .A(n10159), .ZN(n10001) );
  NOR2_X1 U12468 ( .A1(n12157), .A2(n12154), .ZN(n9794) );
  AND2_X1 U12469 ( .A1(n13751), .A2(n13360), .ZN(n11787) );
  INV_X1 U12470 ( .A(n11787), .ZN(n11879) );
  INV_X2 U12471 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10809) );
  AND2_X1 U12472 ( .A1(n14317), .A2(n10035), .ZN(n14283) );
  AND2_X1 U12473 ( .A1(n15159), .A2(n9789), .ZN(n15141) );
  NAND2_X1 U12474 ( .A1(n14317), .A2(n10034), .ZN(n14269) );
  NOR2_X1 U12475 ( .A1(n14058), .A2(n10040), .ZN(n14339) );
  AND2_X1 U12476 ( .A1(n9739), .A2(n10097), .ZN(n15077) );
  AND2_X1 U12477 ( .A1(n15121), .A2(n9825), .ZN(n9795) );
  AND2_X1 U12478 ( .A1(n13923), .A2(n13995), .ZN(n13993) );
  AND4_X1 U12479 ( .A1(n12006), .A2(n12005), .A3(n12004), .A4(n12003), .ZN(
        n9796) );
  NOR2_X1 U12480 ( .A1(n10811), .A2(n10810), .ZN(n9797) );
  OR2_X1 U12481 ( .A1(n20096), .A2(n11525), .ZN(n9798) );
  AND2_X1 U12482 ( .A1(n11276), .A2(n11197), .ZN(n9800) );
  AND2_X1 U12483 ( .A1(n10928), .A2(n10929), .ZN(n11070) );
  OAI21_X1 U12484 ( .B1(n12169), .B2(n10118), .A(n10117), .ZN(n15047) );
  NAND2_X1 U12485 ( .A1(n10125), .A2(n12063), .ZN(n15510) );
  NAND2_X1 U12486 ( .A1(n12149), .A2(n12148), .ZN(n15088) );
  NAND2_X1 U12487 ( .A1(n15120), .A2(n15121), .ZN(n15195) );
  NAND2_X1 U12488 ( .A1(n9967), .A2(n9965), .ZN(n15079) );
  XOR2_X1 U12489 ( .A(n12769), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .Z(
        n9801) );
  AND2_X1 U12490 ( .A1(n11922), .A2(n11917), .ZN(n12010) );
  NAND2_X1 U12491 ( .A1(n9914), .A2(n9771), .ZN(n9802) );
  XNOR2_X1 U12492 ( .A(n10811), .B(n10810), .ZN(n11895) );
  INV_X1 U12493 ( .A(n11895), .ZN(n9867) );
  NAND2_X1 U12494 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10158) );
  NOR2_X1 U12495 ( .A1(n14903), .A2(n10144), .ZN(n12647) );
  NAND2_X1 U12496 ( .A1(n12341), .A2(n12340), .ZN(n15525) );
  OR2_X1 U12497 ( .A1(n12900), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9803) );
  NAND2_X1 U12498 ( .A1(n12389), .A2(n12388), .ZN(n13477) );
  NOR2_X1 U12499 ( .A1(n14016), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9805) );
  AND2_X1 U12500 ( .A1(n15972), .A2(n9878), .ZN(n9806) );
  OR2_X1 U12501 ( .A1(n12169), .A2(n12172), .ZN(n9807) );
  NOR2_X1 U12502 ( .A1(n14240), .A2(n14242), .ZN(n11722) );
  AND2_X1 U12503 ( .A1(n12330), .A2(n12328), .ZN(n9808) );
  AND2_X1 U12504 ( .A1(n10010), .A2(n13491), .ZN(n9809) );
  INV_X1 U12505 ( .A(n12001), .ZN(n15614) );
  OR2_X1 U12506 ( .A1(n12608), .A2(n12607), .ZN(n9810) );
  NOR2_X1 U12507 ( .A1(n9792), .A2(n14991), .ZN(n14985) );
  NAND2_X1 U12508 ( .A1(n9967), .A2(n9964), .ZN(n15069) );
  INV_X1 U12509 ( .A(n10102), .ZN(n17526) );
  NAND2_X1 U12510 ( .A1(n10103), .A2(n17892), .ZN(n10102) );
  AND2_X1 U12511 ( .A1(n10125), .A2(n9976), .ZN(n15204) );
  INV_X1 U12512 ( .A(n10112), .ZN(n9975) );
  AOI21_X1 U12513 ( .B1(n9795), .B2(n10113), .A(n12082), .ZN(n10112) );
  NAND2_X1 U12514 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n9811) );
  AND3_X1 U12515 ( .A1(n11913), .A2(n11915), .A3(n11923), .ZN(n9812) );
  OR2_X1 U12516 ( .A1(n14978), .A2(n14979), .ZN(n9813) );
  AND2_X1 U12517 ( .A1(n12180), .A2(n10726), .ZN(n9814) );
  NOR2_X1 U12518 ( .A1(n16309), .A2(n9884), .ZN(n9815) );
  AND2_X1 U12519 ( .A1(n14177), .A2(n9935), .ZN(n9816) );
  NAND2_X1 U12520 ( .A1(n12048), .A2(n12336), .ZN(n12327) );
  OR2_X1 U12521 ( .A1(n12150), .A2(n10707), .ZN(n10148) );
  AND2_X1 U12522 ( .A1(n12159), .A2(n15316), .ZN(n15082) );
  NAND2_X1 U12523 ( .A1(n10233), .A2(n10281), .ZN(n10547) );
  INV_X1 U12524 ( .A(n14350), .ZN(n14337) );
  INV_X1 U12525 ( .A(n12158), .ZN(n12762) );
  OR2_X1 U12526 ( .A1(n10080), .A2(n13984), .ZN(n9817) );
  NOR2_X1 U12527 ( .A1(n13854), .A2(n10022), .ZN(n13943) );
  AND2_X1 U12528 ( .A1(n13923), .A2(n10044), .ZN(n14051) );
  AND2_X1 U12529 ( .A1(n14760), .A2(n9783), .ZN(n9818) );
  NAND2_X1 U12530 ( .A1(n13723), .A2(n13793), .ZN(n13104) );
  NAND2_X1 U12531 ( .A1(n14760), .A2(n14744), .ZN(n14728) );
  AND2_X1 U12532 ( .A1(n14795), .A2(n14794), .ZN(n9819) );
  AND2_X1 U12533 ( .A1(n10168), .A2(n9995), .ZN(n9820) );
  OR2_X1 U12534 ( .A1(n14058), .A2(n14357), .ZN(n9821) );
  INV_X1 U12535 ( .A(n11786), .ZN(n14206) );
  AND2_X1 U12536 ( .A1(n13751), .A2(n13748), .ZN(n11786) );
  INV_X1 U12537 ( .A(n14206), .ZN(n13381) );
  INV_X1 U12538 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20639) );
  AND2_X1 U12539 ( .A1(n13941), .A2(n14962), .ZN(n14795) );
  AND2_X1 U12540 ( .A1(n14760), .A2(n10015), .ZN(n14907) );
  NOR2_X1 U12541 ( .A1(n14824), .A2(n14826), .ZN(n14825) );
  NAND2_X1 U12542 ( .A1(n11402), .A2(n11401), .ZN(n13706) );
  AND3_X1 U12543 ( .A1(n11158), .A2(n13201), .A3(n13748), .ZN(n13153) );
  OR2_X1 U12544 ( .A1(n10086), .A2(n14814), .ZN(n9822) );
  XNOR2_X1 U12545 ( .A(n12052), .B(n13970), .ZN(n13968) );
  INV_X1 U12546 ( .A(n12055), .ZN(n9913) );
  NOR2_X1 U12547 ( .A1(n13676), .A2(n10006), .ZN(n13723) );
  NAND2_X1 U12548 ( .A1(n9969), .A2(n13762), .ZN(n19191) );
  OR2_X1 U12549 ( .A1(n12900), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9823) );
  AND2_X1 U12550 ( .A1(n13923), .A2(n10043), .ZN(n14050) );
  INV_X1 U12551 ( .A(n13643), .ZN(n13904) );
  NAND4_X1 U12552 ( .A1(n10358), .A2(n10357), .A3(n10356), .A4(n10355), .ZN(
        n12306) );
  NAND2_X1 U12553 ( .A1(n11879), .A2(n11786), .ZN(n11823) );
  AND2_X1 U12554 ( .A1(n10175), .A2(n9998), .ZN(n9824) );
  NAND2_X1 U12555 ( .A1(n18968), .A2(n12080), .ZN(n9825) );
  INV_X1 U12556 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11280) );
  AND2_X1 U12557 ( .A1(n14154), .A2(n11721), .ZN(n9826) );
  XNOR2_X1 U12558 ( .A(n14934), .B(n12586), .ZN(n14928) );
  AND2_X2 U12559 ( .A1(n10927), .A2(n13459), .ZN(n11260) );
  NOR2_X1 U12560 ( .A1(n14945), .A2(n12480), .ZN(n14933) );
  OR2_X1 U12561 ( .A1(n13109), .A2(n9817), .ZN(n9827) );
  INV_X1 U12562 ( .A(n13068), .ZN(n17665) );
  NOR2_X1 U12563 ( .A1(n18721), .A2(n17864), .ZN(n13068) );
  INV_X1 U12564 ( .A(n17784), .ZN(n17720) );
  AND2_X1 U12565 ( .A1(n17818), .A2(n16337), .ZN(n17784) );
  NOR2_X1 U12566 ( .A1(n13063), .A2(n18106), .ZN(n9828) );
  NOR2_X1 U12567 ( .A1(n15016), .A2(n14780), .ZN(n14764) );
  AND2_X1 U12568 ( .A1(n13730), .A2(n12404), .ZN(n9829) );
  NAND2_X1 U12569 ( .A1(n13107), .A2(n10585), .ZN(n13109) );
  NAND2_X1 U12570 ( .A1(n10125), .A2(n10124), .ZN(n15217) );
  AND2_X2 U12571 ( .A1(n13459), .A2(n10930), .ZN(n11253) );
  NOR2_X1 U12572 ( .A1(n13940), .A2(n13939), .ZN(n13941) );
  INV_X1 U12573 ( .A(n9953), .ZN(n14272) );
  NOR2_X1 U12574 ( .A1(n14271), .A2(n14273), .ZN(n9953) );
  AND2_X1 U12575 ( .A1(n14353), .A2(n14354), .ZN(n9830) );
  INV_X1 U12576 ( .A(n9959), .ZN(n14319) );
  NOR3_X1 U12577 ( .A1(n14334), .A2(n9961), .A3(n9962), .ZN(n9959) );
  INV_X1 U12578 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n20789) );
  AND2_X1 U12579 ( .A1(n13681), .A2(n13684), .ZN(n9831) );
  AND2_X1 U12580 ( .A1(n11334), .A2(n11333), .ZN(n11393) );
  AND2_X1 U12581 ( .A1(n18221), .A2(n18225), .ZN(n9832) );
  XNOR2_X1 U12582 ( .A(n12608), .B(n12607), .ZN(n14911) );
  AND2_X1 U12583 ( .A1(n9957), .A2(n9955), .ZN(n9833) );
  NAND2_X1 U12584 ( .A1(n9923), .A2(n9922), .ZN(n9921) );
  AND2_X1 U12585 ( .A1(n9784), .A2(n14348), .ZN(n9834) );
  AND2_X1 U12586 ( .A1(n9779), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9835) );
  AND2_X1 U12587 ( .A1(n10033), .A2(n10034), .ZN(n9836) );
  INV_X1 U12588 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n9987) );
  NOR2_X1 U12589 ( .A1(n11351), .A2(n20212), .ZN(n9837) );
  INV_X1 U12590 ( .A(n19215), .ZN(n16223) );
  NOR3_X1 U12591 ( .A1(n19433), .A2(n19467), .A3(n10692), .ZN(n9838) );
  AND2_X1 U12592 ( .A1(n13417), .A2(n10025), .ZN(n13490) );
  NAND2_X1 U12593 ( .A1(n15532), .A2(n15531), .ZN(n14824) );
  AND2_X1 U12594 ( .A1(n14080), .A2(n9784), .ZN(n9839) );
  NAND2_X1 U12595 ( .A1(n10175), .A2(n9786), .ZN(n10179) );
  OR2_X1 U12596 ( .A1(n14979), .A2(n12294), .ZN(n9840) );
  AND2_X1 U12597 ( .A1(n14080), .A2(n9834), .ZN(n14347) );
  NOR2_X1 U12598 ( .A1(n14824), .A2(n9822), .ZN(n9841) );
  INV_X1 U12599 ( .A(n20085), .ZN(n14712) );
  INV_X1 U12600 ( .A(n14712), .ZN(n20070) );
  OR2_X1 U12601 ( .A1(n12352), .A2(n19852), .ZN(n16227) );
  INV_X1 U12602 ( .A(n16227), .ZN(n19219) );
  AND2_X1 U12603 ( .A1(n13421), .A2(n13420), .ZN(n13419) );
  NOR2_X1 U12604 ( .A1(n13850), .A2(n13849), .ZN(n13813) );
  INV_X1 U12605 ( .A(n16498), .ZN(n9983) );
  NOR2_X1 U12606 ( .A1(n9952), .A2(n14266), .ZN(n9842) );
  OR2_X1 U12607 ( .A1(n12150), .A2(n10712), .ZN(n9843) );
  NOR2_X1 U12608 ( .A1(n12913), .A2(n10109), .ZN(n9844) );
  NAND2_X1 U12609 ( .A1(n14958), .A2(n14001), .ZN(n9845) );
  AND2_X1 U12610 ( .A1(n14067), .A2(n14076), .ZN(n9846) );
  AND2_X1 U12611 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n9847) );
  INV_X1 U12612 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n18874) );
  INV_X1 U12613 ( .A(n14794), .ZN(n10014) );
  INV_X1 U12614 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n9997) );
  OR2_X1 U12615 ( .A1(n18882), .A2(n19869), .ZN(n19198) );
  INV_X1 U12616 ( .A(n19198), .ZN(n16190) );
  INV_X1 U12617 ( .A(n14777), .ZN(n10012) );
  INV_X1 U12618 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9906) );
  INV_X1 U12619 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n9999) );
  INV_X1 U12620 ( .A(n17710), .ZN(n9930) );
  OR2_X1 U12621 ( .A1(n18193), .A2(n18789), .ZN(n9848) );
  INV_X1 U12622 ( .A(n12754), .ZN(n10121) );
  AND2_X1 U12623 ( .A1(n17542), .A2(n9766), .ZN(n9849) );
  AND2_X1 U12624 ( .A1(n10097), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9850) );
  NAND2_X1 U12625 ( .A1(n15749), .A2(n14675), .ZN(n9851) );
  INV_X1 U12626 ( .A(n15278), .ZN(n10123) );
  INV_X1 U12627 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10098) );
  INV_X1 U12628 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10005) );
  NAND3_X2 U12629 ( .A1(n18866), .A2(n20757), .A3(n18865), .ZN(n18193) );
  NAND2_X1 U12630 ( .A1(n13035), .A2(n15679), .ZN(n18679) );
  NAND4_X1 U12631 ( .A1(n18193), .A2(n18847), .A3(n18717), .A4(n18706), .ZN(
        n16783) );
  AOI22_X2 U12632 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20151), .B1(DATAI_26_), 
        .B2(n20108), .ZN(n20605) );
  AOI22_X2 U12633 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20151), .B1(DATAI_27_), 
        .B2(n20108), .ZN(n20611) );
  AOI22_X2 U12634 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20151), .B1(DATAI_28_), 
        .B2(n20108), .ZN(n20617) );
  AOI22_X2 U12635 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20151), .B1(DATAI_29_), 
        .B2(n20108), .ZN(n20623) );
  AOI22_X2 U12636 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20151), .B1(DATAI_30_), 
        .B2(n20108), .ZN(n20629) );
  NOR3_X2 U12637 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18713), .A3(
        n18293), .ZN(n18266) );
  NOR3_X2 U12638 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18713), .A3(
        n18427), .ZN(n18400) );
  NOR3_X2 U12639 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18713), .A3(
        n18479), .ZN(n18447) );
  NAND2_X1 U12640 ( .A1(n16334), .A2(n9717), .ZN(n10107) );
  NOR3_X4 U12641 ( .A1(n14428), .A2(n20148), .A3(n14185), .ZN(n14424) );
  INV_X1 U12642 ( .A(n14409), .ZN(n14428) );
  AOI22_X2 U12643 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20151), .B1(DATAI_25_), 
        .B2(n20108), .ZN(n20599) );
  NOR3_X2 U12644 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18713), .A3(
        n18385), .ZN(n18354) );
  NAND3_X1 U12645 ( .A1(n9969), .A2(n11994), .A3(n13762), .ZN(n9852) );
  OR2_X1 U12646 ( .A1(n11990), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13762) );
  NAND2_X1 U12647 ( .A1(n11990), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13761) );
  AND2_X2 U12648 ( .A1(n10734), .A2(n10727), .ZN(n10733) );
  NAND2_X2 U12649 ( .A1(n10231), .A2(n10232), .ZN(n10630) );
  INV_X1 U12650 ( .A(n11931), .ZN(n9858) );
  NAND2_X1 U12651 ( .A1(n9857), .A2(n9743), .ZN(n9856) );
  NAND3_X1 U12652 ( .A1(n9859), .A2(n9858), .A3(n9812), .ZN(n9857) );
  NAND2_X1 U12653 ( .A1(n9861), .A2(n19869), .ZN(n9860) );
  INV_X1 U12654 ( .A(n9865), .ZN(n9861) );
  NAND4_X1 U12655 ( .A1(n12724), .A2(n12258), .A3(n10723), .A4(n19237), .ZN(
        n9865) );
  NAND2_X1 U12656 ( .A1(n10722), .A2(n9865), .ZN(n10775) );
  NAND2_X2 U12657 ( .A1(n9869), .A2(n9866), .ZN(n13777) );
  NAND2_X2 U12658 ( .A1(n11898), .A2(n11897), .ZN(n9871) );
  NAND2_X1 U12659 ( .A1(n9871), .A2(n10799), .ZN(n11896) );
  NAND2_X1 U12660 ( .A1(n13530), .A2(n9875), .ZN(n9874) );
  INV_X1 U12661 ( .A(n20063), .ZN(n9875) );
  NAND2_X1 U12662 ( .A1(n13529), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n9876) );
  XNOR2_X1 U12663 ( .A(n13530), .B(n20063), .ZN(n13529) );
  OAI21_X2 U12664 ( .B1(n13669), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11278), 
        .ZN(n13367) );
  NAND2_X2 U12665 ( .A1(n11193), .A2(n11192), .ZN(n11276) );
  NAND2_X1 U12666 ( .A1(n13903), .A2(n9806), .ZN(n13949) );
  NAND2_X1 U12667 ( .A1(n14169), .A2(n9880), .ZN(n9944) );
  NAND3_X1 U12668 ( .A1(n9885), .A2(n9815), .A3(n9883), .ZN(P3_U2800) );
  INV_X4 U12669 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n21023) );
  NAND2_X1 U12670 ( .A1(n15659), .A2(n9832), .ZN(n9889) );
  AOI21_X1 U12671 ( .B1(n15659), .B2(n13033), .A(n13032), .ZN(n18651) );
  INV_X1 U12672 ( .A(n18681), .ZN(n9891) );
  OR2_X2 U12673 ( .A1(n17664), .A2(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17662) );
  OAI21_X2 U12674 ( .B1(n9898), .B2(n17788), .A(n9897), .ZN(n13073) );
  INV_X1 U12675 ( .A(n12896), .ZN(n9898) );
  AND2_X2 U12676 ( .A1(n13073), .A2(n10104), .ZN(n18114) );
  INV_X1 U12677 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n9900) );
  INV_X2 U12678 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18820) );
  AND2_X4 U12679 ( .A1(n15579), .A2(n14108), .ZN(n10660) );
  NOR2_X2 U12680 ( .A1(n11984), .A2(n11983), .ZN(n11982) );
  NOR2_X2 U12681 ( .A1(n12111), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12088) );
  NOR2_X2 U12682 ( .A1(n12104), .A2(n10711), .ZN(n9917) );
  INV_X1 U12683 ( .A(n17794), .ZN(n9923) );
  OAI211_X2 U12684 ( .C1(n11193), .C2(n9932), .A(n11206), .B(n9931), .ZN(
        n13480) );
  NAND2_X1 U12685 ( .A1(n14459), .A2(n9933), .ZN(n14434) );
  INV_X1 U12686 ( .A(n14448), .ZN(n9935) );
  NAND2_X1 U12687 ( .A1(n14533), .A2(n14170), .ZN(n9936) );
  NAND2_X1 U12688 ( .A1(n14164), .A2(n15946), .ZN(n14534) );
  NAND2_X1 U12689 ( .A1(n9944), .A2(n9943), .ZN(n15748) );
  NAND4_X1 U12690 ( .A1(n11153), .A2(n11151), .A3(n11150), .A4(n11152), .ZN(
        n9946) );
  NAND3_X1 U12691 ( .A1(n9804), .A2(n20097), .A3(n11376), .ZN(n11386) );
  NAND2_X1 U12692 ( .A1(n11155), .A2(n11154), .ZN(n9949) );
  NOR2_X1 U12693 ( .A1(n13748), .A2(n13751), .ZN(n11183) );
  INV_X1 U12694 ( .A(n14250), .ZN(n9954) );
  NAND2_X1 U12695 ( .A1(n9956), .A2(n9833), .ZN(n14032) );
  AND2_X2 U12696 ( .A1(n11280), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13459) );
  NOR3_X2 U12697 ( .A1(n14334), .A2(n9961), .A3(n9960), .ZN(n14314) );
  NOR2_X1 U12698 ( .A1(n14334), .A2(n14326), .ZN(n14660) );
  INV_X1 U12699 ( .A(n14659), .ZN(n9962) );
  XNOR2_X2 U12700 ( .A(n11997), .B(n11996), .ZN(n13765) );
  NAND2_X1 U12701 ( .A1(n13765), .A2(n12158), .ZN(n11974) );
  INV_X1 U12702 ( .A(n12148), .ZN(n9963) );
  NOR2_X1 U12703 ( .A1(n9963), .A2(n10127), .ZN(n9968) );
  NAND2_X1 U12704 ( .A1(n10125), .A2(n9973), .ZN(n9970) );
  NAND2_X1 U12705 ( .A1(n9970), .A2(n9971), .ZN(n15183) );
  NAND3_X1 U12706 ( .A1(n16495), .A2(n16494), .A3(n9978), .ZN(P3_U2641) );
  INV_X1 U12707 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n9981) );
  NAND2_X1 U12708 ( .A1(n16508), .A2(n16469), .ZN(n9984) );
  XNOR2_X1 U12709 ( .A(n9985), .B(n16488), .ZN(n16492) );
  NAND3_X1 U12710 ( .A1(n9988), .A2(n17777), .A3(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17679) );
  NAND2_X1 U12711 ( .A1(n16576), .A2(n16469), .ZN(n9990) );
  NAND2_X1 U12712 ( .A1(n9990), .A2(n9991), .ZN(n16561) );
  INV_X1 U12713 ( .A(n9992), .ZN(n16575) );
  AND2_X1 U12714 ( .A1(n12745), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9993) );
  NAND2_X1 U12715 ( .A1(n10020), .A2(n10021), .ZN(n14952) );
  NOR2_X2 U12716 ( .A1(n14945), .A2(n10026), .ZN(n14934) );
  NAND2_X1 U12717 ( .A1(n11102), .A2(n11180), .ZN(n10029) );
  OAI21_X1 U12718 ( .B1(n20139), .B2(n13445), .A(n11159), .ZN(n10030) );
  AND2_X2 U12719 ( .A1(n13468), .A2(n10926), .ZN(n11252) );
  NAND2_X1 U12720 ( .A1(n10054), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11198) );
  NAND2_X1 U12721 ( .A1(n10054), .A2(n10032), .ZN(n10031) );
  AND2_X2 U12722 ( .A1(n14317), .A2(n9836), .ZN(n14255) );
  NOR2_X2 U12723 ( .A1(n14058), .A2(n10037), .ZN(n14331) );
  OAI21_X1 U12724 ( .B1(n11348), .B2(n11349), .A(n11350), .ZN(n13363) );
  NAND2_X1 U12725 ( .A1(n11348), .A2(n11349), .ZN(n11350) );
  OAI211_X1 U12726 ( .C1(n11348), .C2(n10050), .A(n13362), .B(n10048), .ZN(
        n20061) );
  NAND2_X1 U12727 ( .A1(n11348), .A2(n10049), .ZN(n10048) );
  NOR2_X1 U12728 ( .A1(n11349), .A2(n13643), .ZN(n10049) );
  NAND2_X1 U12729 ( .A1(n10055), .A2(n11171), .ZN(n10051) );
  NAND2_X1 U12730 ( .A1(n10051), .A2(n10056), .ZN(n10052) );
  XNOR2_X1 U12731 ( .A(n11221), .B(n11220), .ZN(n11351) );
  NAND3_X1 U12732 ( .A1(n10053), .A2(n11178), .A3(n10052), .ZN(n11221) );
  NAND4_X1 U12733 ( .A1(n10055), .A2(n13447), .A3(n11171), .A4(n11161), .ZN(
        n10054) );
  NAND2_X1 U12734 ( .A1(n14433), .A2(n14174), .ZN(n10065) );
  NAND2_X1 U12735 ( .A1(n14433), .A2(n10058), .ZN(n10057) );
  NAND2_X1 U12736 ( .A1(n14180), .A2(n10061), .ZN(n10060) );
  NOR2_X1 U12737 ( .A1(n9805), .A2(n10068), .ZN(n10067) );
  NAND2_X2 U12738 ( .A1(n14157), .A2(n10141), .ZN(n14558) );
  NAND2_X1 U12739 ( .A1(n15928), .A2(n10069), .ZN(n14173) );
  NAND2_X1 U12740 ( .A1(n13775), .A2(n10412), .ZN(n10070) );
  NAND2_X1 U12741 ( .A1(n10070), .A2(n10071), .ZN(n10434) );
  AND2_X2 U12742 ( .A1(n13274), .A2(n13275), .ZN(n13277) );
  NAND2_X1 U12743 ( .A1(n10091), .A2(n10094), .ZN(n10092) );
  INV_X1 U12744 ( .A(n13967), .ZN(n10094) );
  NAND2_X2 U12745 ( .A1(n12332), .A2(n9808), .ZN(n10093) );
  OR2_X2 U12746 ( .A1(n13967), .A2(n13964), .ZN(n12332) );
  NAND2_X1 U12747 ( .A1(n9739), .A2(n10096), .ZN(n12728) );
  NAND2_X1 U12748 ( .A1(n10100), .A2(n20760), .ZN(n10099) );
  NAND2_X1 U12749 ( .A1(n17815), .A2(n17816), .ZN(n10100) );
  NAND3_X2 U12750 ( .A1(n10152), .A2(n12830), .A3(n10136), .ZN(n17391) );
  INV_X1 U12751 ( .A(n12169), .ZN(n12756) );
  INV_X1 U12752 ( .A(n12755), .ZN(n10122) );
  NAND3_X2 U12753 ( .A1(n12060), .A2(n12059), .A3(n12058), .ZN(n10125) );
  AND2_X1 U12754 ( .A1(n11998), .A2(n11997), .ZN(n12307) );
  NAND3_X1 U12755 ( .A1(n11998), .A2(n11997), .A3(n12306), .ZN(n12024) );
  NAND2_X1 U12756 ( .A1(n11919), .A2(n11918), .ZN(n12001) );
  INV_X1 U12757 ( .A(n11929), .ZN(n11911) );
  NAND2_X1 U12758 ( .A1(n11350), .A2(n11274), .ZN(n11359) );
  NAND2_X1 U12759 ( .A1(n14050), .A2(n14059), .ZN(n14058) );
  XNOR2_X1 U12760 ( .A(n11342), .B(n11360), .ZN(n13517) );
  NAND2_X1 U12761 ( .A1(n11221), .A2(n11220), .ZN(n11275) );
  NAND2_X1 U12762 ( .A1(n11974), .A2(n14849), .ZN(n11990) );
  INV_X1 U12763 ( .A(n13706), .ZN(n11403) );
  XNOR2_X1 U12764 ( .A(n12701), .B(n12700), .ZN(n14203) );
  NAND2_X1 U12765 ( .A1(n14331), .A2(n14333), .ZN(n14323) );
  AOI21_X2 U12766 ( .B1(n9760), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n11126), .ZN(n11132) );
  OR2_X1 U12767 ( .A1(n11901), .A2(n11900), .ZN(n11902) );
  AND2_X1 U12768 ( .A1(n10807), .A2(n10766), .ZN(n10767) );
  OR2_X1 U12769 ( .A1(n9762), .A2(n13972), .ZN(n10806) );
  XNOR2_X1 U12770 ( .A(n12627), .B(n12625), .ZN(n14905) );
  NOR2_X1 U12771 ( .A1(n12794), .A2(n16826), .ZN(n12835) );
  NOR2_X1 U12772 ( .A1(n16826), .A2(n12791), .ZN(n16992) );
  OR3_X1 U12773 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17600), .ZN(n10130) );
  OR2_X1 U12774 ( .A1(n18679), .A2(n16337), .ZN(n10131) );
  INV_X1 U12775 ( .A(n10352), .ZN(n12484) );
  OR2_X1 U12776 ( .A1(n12680), .A2(n12679), .ZN(n10133) );
  OR2_X1 U12777 ( .A1(n10178), .A2(n14762), .ZN(n10134) );
  AND4_X1 U12778 ( .A1(n10452), .A2(n10451), .A3(n10450), .A4(n10449), .ZN(
        n10135) );
  AND3_X1 U12779 ( .A1(n12827), .A2(n12826), .A3(n12825), .ZN(n10136) );
  INV_X1 U12780 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13931) );
  NOR2_X1 U12781 ( .A1(n13425), .A2(n20490), .ZN(n10137) );
  AND2_X1 U12782 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_22__SCAN_IN), 
        .ZN(n10138) );
  OR2_X1 U12783 ( .A1(n17558), .A2(n12900), .ZN(n10139) );
  AND2_X1 U12784 ( .A1(n11932), .A2(n19223), .ZN(n10140) );
  OR2_X1 U12785 ( .A1(n14160), .A2(n14158), .ZN(n10141) );
  INV_X1 U12786 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n12376) );
  AND2_X1 U12787 ( .A1(n12523), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n10142) );
  NOR2_X1 U12788 ( .A1(n20455), .A2(n20486), .ZN(n10143) );
  OR2_X1 U12789 ( .A1(n17446), .A2(n18217), .ZN(n10145) );
  NAND2_X1 U12790 ( .A1(n14350), .A2(n20148), .ZN(n20002) );
  INV_X1 U12791 ( .A(n20002), .ZN(n11892) );
  AND2_X2 U12792 ( .A1(n12686), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10287) );
  INV_X1 U12793 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14175) );
  INV_X1 U12794 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12371) );
  INV_X2 U12795 ( .A(n17238), .ZN(n17233) );
  AND2_X1 U12796 ( .A1(n14172), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10146) );
  INV_X1 U12797 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n14146) );
  AND2_X1 U12798 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(P3_EAX_REG_13__SCAN_IN), 
        .ZN(n10147) );
  INV_X1 U12799 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12905) );
  INV_X1 U12800 ( .A(n14954), .ZN(n10879) );
  NOR2_X1 U12801 ( .A1(n20455), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10149) );
  AND2_X1 U12802 ( .A1(n14778), .A2(n14759), .ZN(n10150) );
  INV_X1 U12803 ( .A(n13257), .ZN(n13251) );
  AND4_X1 U12804 ( .A1(n12824), .A2(n12823), .A3(n12822), .A4(n12821), .ZN(
        n10152) );
  INV_X1 U12805 ( .A(n12834), .ZN(n17132) );
  OR2_X1 U12806 ( .A1(n18452), .A2(n18359), .ZN(n18454) );
  INV_X1 U12807 ( .A(n12742), .ZN(n10800) );
  INV_X1 U12808 ( .A(n15975), .ZN(n20106) );
  INV_X1 U12809 ( .A(n14283), .ZN(n14312) );
  NOR2_X2 U12810 ( .A1(n14323), .A2(n14324), .ZN(n14322) );
  INV_X1 U12811 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n16287) );
  AND2_X1 U12812 ( .A1(n11124), .A2(n11123), .ZN(n10153) );
  INV_X1 U12813 ( .A(n11041), .ZN(n14118) );
  INV_X1 U12814 ( .A(n12257), .ZN(n10745) );
  NAND2_X1 U12815 ( .A1(n12009), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11936) );
  NAND2_X1 U12816 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20517), .ZN(
        n11739) );
  AND2_X1 U12817 ( .A1(n11742), .A2(n11725), .ZN(n11749) );
  INV_X1 U12818 ( .A(n14523), .ZN(n14167) );
  OR2_X1 U12819 ( .A1(n11332), .A2(n11331), .ZN(n13907) );
  OR2_X1 U12820 ( .A1(n11182), .A2(n13748), .ZN(n11171) );
  INV_X1 U12821 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10670) );
  NAND2_X1 U12822 ( .A1(n10739), .A2(n12215), .ZN(n12222) );
  NAND2_X1 U12823 ( .A1(n12706), .A2(n10729), .ZN(n10731) );
  INV_X1 U12824 ( .A(n12247), .ZN(n12194) );
  AND2_X1 U12825 ( .A1(n10617), .A2(n10616), .ZN(n10619) );
  XNOR2_X1 U12826 ( .A(n11280), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11759) );
  OR2_X1 U12827 ( .A1(n11740), .A2(n11739), .ZN(n11742) );
  INV_X1 U12828 ( .A(n11247), .ZN(n11248) );
  INV_X1 U12829 ( .A(n12518), .ZN(n10392) );
  NOR2_X1 U12830 ( .A1(n11758), .A2(n11759), .ZN(n11757) );
  INV_X1 U12831 ( .A(n11070), .ZN(n10957) );
  INV_X1 U12832 ( .A(n14346), .ZN(n11563) );
  INV_X1 U12833 ( .A(n13862), .ZN(n11421) );
  INV_X1 U12834 ( .A(n13820), .ZN(n11404) );
  OR2_X1 U12835 ( .A1(n11319), .A2(n11318), .ZN(n13808) );
  OR2_X1 U12836 ( .A1(n11243), .A2(n11242), .ZN(n13520) );
  OR2_X1 U12837 ( .A1(n11218), .A2(n11217), .ZN(n13522) );
  AOI22_X1 U12838 ( .A1(n10968), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9752), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11099) );
  AND4_X1 U12839 ( .A1(n11065), .A2(n11064), .A3(n11063), .A4(n11062), .ZN(
        n11066) );
  AOI21_X1 U12840 ( .B1(n10679), .B2(n10677), .A(n10675), .ZN(n10684) );
  OR2_X1 U12841 ( .A1(n12603), .A2(n12605), .ZN(n12609) );
  AND2_X1 U12842 ( .A1(n12559), .A2(n12564), .ZN(n12582) );
  AND4_X1 U12843 ( .A1(n10384), .A2(n10383), .A3(n10382), .A4(n10381), .ZN(
        n10385) );
  NAND3_X1 U12844 ( .A1(n11167), .A2(n13748), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11764) );
  INV_X1 U12845 ( .A(n14284), .ZN(n11688) );
  INV_X1 U12846 ( .A(n14391), .ZN(n11659) );
  INV_X1 U12847 ( .A(n11733), .ZN(n13386) );
  OAI21_X1 U12848 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n11196), .A(
        n11195), .ZN(n11197) );
  AND2_X1 U12849 ( .A1(n12179), .A2(n12178), .ZN(n12209) );
  INV_X1 U12850 ( .A(n12465), .ZN(n12497) );
  INV_X1 U12851 ( .A(n10263), .ZN(n10264) );
  INV_X1 U12852 ( .A(n15046), .ZN(n12763) );
  INV_X1 U12853 ( .A(n12752), .ZN(n12753) );
  OR2_X1 U12854 ( .A1(n13103), .A2(n12158), .ZN(n12122) );
  NAND2_X1 U12855 ( .A1(n10661), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12481) );
  NOR2_X1 U12856 ( .A1(n18238), .A2(n17248), .ZN(n15667) );
  INV_X1 U12857 ( .A(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n21022) );
  NOR2_X1 U12858 ( .A1(n17372), .A2(n12864), .ZN(n12889) );
  INV_X1 U12859 ( .A(n12882), .ZN(n12883) );
  INV_X1 U12860 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12866) );
  NAND2_X1 U12861 ( .A1(n11270), .A2(n11251), .ZN(n11775) );
  NAND2_X1 U12862 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11368) );
  NOR2_X1 U12863 ( .A1(n19967), .A2(n20640), .ZN(n13747) );
  AND2_X1 U12864 ( .A1(n11812), .A2(n11811), .ZN(n16049) );
  NOR2_X1 U12865 ( .A1(n11478), .A2(n15885), .ZN(n11493) );
  AND2_X1 U12866 ( .A1(n20640), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14136) );
  INV_X1 U12867 ( .A(n13531), .ZN(n11365) );
  AND2_X1 U12868 ( .A1(n14545), .A2(n14609), .ZN(n14178) );
  AND2_X1 U12869 ( .A1(n11829), .A2(n11828), .ZN(n14031) );
  OR2_X1 U12870 ( .A1(n11294), .A2(n11293), .ZN(n13645) );
  NAND2_X1 U12871 ( .A1(n11359), .A2(n13367), .ZN(n11360) );
  NAND2_X1 U12872 ( .A1(n10686), .A2(n10685), .ZN(n12197) );
  INV_X1 U12873 ( .A(n13122), .ZN(n10845) );
  NAND2_X1 U12874 ( .A1(n10265), .A2(n10264), .ZN(n13274) );
  OR3_X1 U12875 ( .A1(n14750), .A2(n12158), .A3(n15338), .ZN(n15110) );
  INV_X1 U12876 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19385) );
  NAND2_X1 U12877 ( .A1(n12202), .A2(n12199), .ZN(n16276) );
  NAND2_X1 U12878 ( .A1(n15667), .A2(n9832), .ZN(n15640) );
  AND2_X1 U12879 ( .A1(n17334), .A2(n10147), .ZN(n17243) );
  NAND2_X1 U12880 ( .A1(n13079), .A2(n13078), .ZN(n13080) );
  NOR2_X1 U12881 ( .A1(n13047), .A2(n13046), .ZN(n13044) );
  INV_X1 U12882 ( .A(n17782), .ZN(n12900) );
  NOR2_X1 U12883 ( .A1(n18679), .A2(n17362), .ZN(n17943) );
  NOR2_X1 U12884 ( .A1(n17380), .A2(n12865), .ZN(n12886) );
  INV_X1 U12885 ( .A(n18107), .ZN(n13035) );
  INV_X1 U12886 ( .A(n13153), .ZN(n13154) );
  OR2_X1 U12887 ( .A1(n11717), .A2(n11716), .ZN(n13739) );
  AND2_X1 U12888 ( .A1(n11664), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n11668) );
  INV_X1 U12889 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15885) );
  AND2_X1 U12890 ( .A1(n13748), .A2(n13747), .ZN(n13753) );
  AND2_X1 U12891 ( .A1(n11815), .A2(n11814), .ZN(n13845) );
  INV_X1 U12892 ( .A(n11413), .ZN(n11525) );
  OR2_X1 U12893 ( .A1(n11720), .A2(n11719), .ZN(n14242) );
  AND2_X1 U12894 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n11631), .ZN(
        n11664) );
  AND2_X1 U12895 ( .A1(n11562), .A2(n11561), .ZN(n14346) );
  NAND2_X1 U12896 ( .A1(n13403), .A2(n13384), .ZN(n15755) );
  INV_X1 U12897 ( .A(n13496), .ZN(n13436) );
  INV_X1 U12898 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20414) );
  INV_X1 U12899 ( .A(n13517), .ZN(n20095) );
  NOR2_X1 U12900 ( .A1(n20299), .A2(n20249), .ZN(n20421) );
  OR2_X1 U12901 ( .A1(n20096), .A2(n13664), .ZN(n20460) );
  INV_X1 U12902 ( .A(n13363), .ZN(n20181) );
  INV_X1 U12903 ( .A(n18957), .ZN(n19031) );
  OR2_X1 U12904 ( .A1(n15177), .A2(n15176), .ZN(n15448) );
  OR2_X1 U12905 ( .A1(n12352), .A2(n12303), .ZN(n15520) );
  AND2_X1 U12906 ( .A1(n16276), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n14103) );
  OR3_X1 U12907 ( .A1(n19353), .A2(n19379), .A3(n10692), .ZN(n19358) );
  INV_X1 U12908 ( .A(n19460), .ZN(n19491) );
  OR3_X1 U12909 ( .A1(n12009), .A2(n19594), .A3(n10692), .ZN(n15631) );
  OR2_X1 U12910 ( .A1(n19825), .A2(n15608), .ZN(n19609) );
  AOI21_X1 U12911 ( .B1(n12939), .B2(n12938), .A(n12937), .ZN(n18682) );
  NOR2_X1 U12912 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16612), .ZN(n16598) );
  NOR2_X1 U12913 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16679), .ZN(n16663) );
  INV_X1 U12914 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16702) );
  NOR2_X1 U12915 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16746), .ZN(n16732) );
  NOR2_X1 U12916 ( .A1(n20783), .A2(n17095), .ZN(n17077) );
  AND2_X1 U12917 ( .A1(n18648), .A2(n13030), .ZN(n15674) );
  NOR2_X1 U12918 ( .A1(n17283), .A2(n17464), .ZN(n17282) );
  NAND2_X1 U12919 ( .A1(n17353), .A2(n17243), .ZN(n17329) );
  INV_X1 U12920 ( .A(n18234), .ZN(n17248) );
  INV_X1 U12921 ( .A(n17871), .ZN(n17861) );
  INV_X1 U12922 ( .A(n17599), .ZN(n17625) );
  INV_X1 U12923 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18659) );
  INV_X1 U12924 ( .A(n15678), .ZN(n18221) );
  NOR2_X1 U12925 ( .A1(n13154), .A2(n19884), .ZN(n13155) );
  NAND2_X1 U12926 ( .A1(n11668), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11685) );
  AND2_X1 U12927 ( .A1(n19927), .A2(n13743), .ZN(n19932) );
  AND3_X1 U12928 ( .A1(n13753), .A2(n13749), .A3(n15724), .ZN(n19959) );
  AND2_X1 U12929 ( .A1(n19927), .A2(n13758), .ZN(n19993) );
  INV_X1 U12930 ( .A(n14599), .ZN(n11893) );
  NOR2_X1 U12931 ( .A1(n14428), .A2(n13569), .ZN(n14429) );
  INV_X1 U12932 ( .A(n13358), .ZN(n20043) );
  NAND2_X1 U12933 ( .A1(n11545), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11558) );
  NAND2_X1 U12934 ( .A1(n11455), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11478) );
  AND2_X1 U12935 ( .A1(n11397), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11416) );
  AND2_X1 U12936 ( .A1(n13496), .A2(n13495), .ZN(n20064) );
  AND2_X1 U12937 ( .A1(n13497), .A2(n20547), .ZN(n15975) );
  AND2_X1 U12938 ( .A1(n14641), .A2(n14567), .ZN(n15985) );
  AND2_X1 U12939 ( .A1(n13797), .A2(n14663), .ZN(n20078) );
  NAND2_X1 U12940 ( .A1(n13379), .A2(n13560), .ZN(n13408) );
  INV_X1 U12941 ( .A(n20180), .ZN(n20152) );
  INV_X1 U12942 ( .A(n20183), .ZN(n20207) );
  INV_X1 U12943 ( .A(n20191), .ZN(n20237) );
  AND2_X1 U12944 ( .A1(n20328), .A2(n20277), .ZN(n20319) );
  INV_X1 U12945 ( .A(n20376), .ZN(n20353) );
  NOR2_X1 U12946 ( .A1(n20517), .A2(n20323), .ZN(n20343) );
  AND2_X1 U12947 ( .A1(n13664), .A2(n13665), .ZN(n20328) );
  NOR2_X2 U12948 ( .A1(n20460), .A2(n20523), .ZN(n20450) );
  INV_X1 U12949 ( .A(n20480), .ZN(n20482) );
  NOR2_X1 U12950 ( .A1(n20182), .A2(n13363), .ZN(n20463) );
  INV_X1 U12951 ( .A(n20638), .ZN(n20574) );
  NAND2_X1 U12952 ( .A1(n20182), .A2(n20181), .ZN(n20523) );
  INV_X1 U12953 ( .A(n20682), .ZN(n20695) );
  INV_X1 U12954 ( .A(n19037), .ZN(n10916) );
  AND2_X1 U12955 ( .A1(n10697), .A2(n16288), .ZN(n18957) );
  INV_X1 U12956 ( .A(n19041), .ZN(n19003) );
  INV_X1 U12957 ( .A(n19026), .ZN(n19029) );
  AND3_X1 U12958 ( .A1(n10454), .A2(n10453), .A3(n10135), .ZN(n13633) );
  INV_X1 U12959 ( .A(n12699), .ZN(n12700) );
  AND2_X1 U12960 ( .A1(n9813), .A2(n14980), .ZN(n16097) );
  INV_X1 U12961 ( .A(n19082), .ZN(n19107) );
  INV_X1 U12962 ( .A(n13145), .ZN(n19185) );
  INV_X1 U12963 ( .A(n14890), .ZN(n16086) );
  AND2_X1 U12964 ( .A1(n16194), .A2(n13191), .ZN(n16187) );
  NAND2_X1 U12965 ( .A1(n12246), .A2(n13249), .ZN(n12352) );
  INV_X1 U12966 ( .A(n19636), .ZN(n19820) );
  INV_X1 U12967 ( .A(n19289), .ZN(n19281) );
  NOR2_X1 U12968 ( .A1(n19491), .A2(n19439), .ZN(n19319) );
  AND2_X1 U12969 ( .A1(n19296), .A2(n19547), .ZN(n19348) );
  INV_X1 U12970 ( .A(n19366), .ZN(n19381) );
  NOR2_X1 U12971 ( .A1(n19357), .A2(n19609), .ZN(n19401) );
  NOR2_X1 U12972 ( .A1(n19439), .A2(n19815), .ZN(n19486) );
  AND2_X1 U12973 ( .A1(n19825), .A2(n19838), .ZN(n19460) );
  NOR2_X2 U12974 ( .A1(n19610), .A2(n19491), .ZN(n19540) );
  NOR2_X1 U12975 ( .A1(n19631), .A2(n19323), .ZN(n19560) );
  INV_X1 U12976 ( .A(n19563), .ZN(n19596) );
  INV_X1 U12977 ( .A(n19631), .ZN(n19461) );
  AND2_X1 U12978 ( .A1(n12237), .A2(n19842), .ZN(n19853) );
  NOR3_X1 U12979 ( .A1(n19861), .A2(n10692), .A3(n16291), .ZN(n19737) );
  OR3_X1 U12980 ( .A1(n12961), .A2(n12960), .A3(n12959), .ZN(n18853) );
  INV_X1 U12981 ( .A(n16837), .ZN(n16827) );
  NOR2_X1 U12982 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16635), .ZN(n16617) );
  NOR2_X1 U12983 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16655), .ZN(n16639) );
  NOR2_X1 U12984 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16699), .ZN(n16684) );
  NOR2_X2 U12985 ( .A1(n18701), .A2(n16461), .ZN(n16807) );
  INV_X1 U12986 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n16801) );
  INV_X1 U12987 ( .A(n16783), .ZN(n16834) );
  AND2_X1 U12988 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17013), .ZN(n16987) );
  NOR2_X1 U12989 ( .A1(n17237), .A2(n16842), .ZN(n17115) );
  AOI21_X1 U12990 ( .B1(n18683), .B2(n15674), .A(n15642), .ZN(n15766) );
  NOR2_X1 U12991 ( .A1(n17472), .A2(n17267), .ZN(n17263) );
  OR2_X1 U12992 ( .A1(n17466), .A2(n17276), .ZN(n17277) );
  NOR2_X1 U12993 ( .A1(n17450), .A2(n17324), .ZN(n17318) );
  NAND2_X1 U12994 ( .A1(P3_EAX_REG_15__SCAN_IN), .A2(n17325), .ZN(n17324) );
  INV_X1 U12995 ( .A(n17460), .ZN(n17490) );
  INV_X1 U12996 ( .A(n17495), .ZN(n17506) );
  INV_X1 U12997 ( .A(n17761), .ZN(n17783) );
  AND2_X1 U12998 ( .A1(n17599), .A2(n17619), .ZN(n17651) );
  NOR2_X1 U12999 ( .A1(n9726), .A2(n18191), .ZN(n18187) );
  NAND2_X1 U13000 ( .A1(n20757), .A2(n18211), .ZN(n18452) );
  NOR2_X1 U13001 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18808), .ZN(
        n18828) );
  INV_X1 U13002 ( .A(n18708), .ZN(n18849) );
  INV_X1 U13003 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18728) );
  NAND2_X1 U13004 ( .A1(n13496), .A2(n13155), .ZN(n13567) );
  INV_X1 U13005 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20906) );
  INV_X1 U13006 ( .A(n19991), .ZN(n19956) );
  INV_X1 U13007 ( .A(n15958), .ZN(n15893) );
  OR2_X1 U13008 ( .A1(n20023), .A2(n20719), .ZN(n20017) );
  INV_X1 U13009 ( .A(n20023), .ZN(n20035) );
  NOR2_X1 U13010 ( .A1(n13567), .A2(n13323), .ZN(n13357) );
  INV_X1 U13011 ( .A(n15979), .ZN(n15978) );
  INV_X1 U13012 ( .A(n20064), .ZN(n15962) );
  OR2_X1 U13013 ( .A1(n16009), .A2(n15985), .ZN(n16006) );
  INV_X1 U13014 ( .A(n20082), .ZN(n16025) );
  INV_X1 U13015 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13484) );
  OR2_X1 U13016 ( .A1(n20217), .A2(n20488), .ZN(n20180) );
  OR2_X1 U13017 ( .A1(n20217), .A2(n20216), .ZN(n20271) );
  NAND2_X1 U13018 ( .A1(n20328), .A2(n20352), .ZN(n20297) );
  AOI22_X1 U13019 ( .A1(n20303), .A2(n20301), .B1(n20300), .B2(n20299), .ZN(
        n20736) );
  INV_X1 U13020 ( .A(n20345), .ZN(n20729) );
  NAND2_X1 U13021 ( .A1(n20328), .A2(n20463), .ZN(n20376) );
  NAND2_X1 U13022 ( .A1(n20464), .A2(n20352), .ZN(n20405) );
  AOI22_X1 U13023 ( .A1(n20419), .A2(n20416), .B1(n20413), .B2(n20412), .ZN(
        n20454) );
  NAND2_X1 U13024 ( .A1(n20464), .A2(n20406), .ZN(n20480) );
  NAND2_X1 U13025 ( .A1(n20464), .A2(n20463), .ZN(n20516) );
  OR2_X1 U13026 ( .A1(n20585), .A2(n20488), .ZN(n20539) );
  OR2_X1 U13027 ( .A1(n20585), .A2(n20523), .ZN(n20578) );
  OR2_X1 U13028 ( .A1(n20551), .A2(n20585), .ZN(n20638) );
  INV_X1 U13029 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20640) );
  INV_X1 U13030 ( .A(n20704), .ZN(n20643) );
  INV_X1 U13031 ( .A(n20713), .ZN(n20715) );
  OR2_X1 U13032 ( .A1(n16265), .A2(n18880), .ZN(n19863) );
  NAND2_X1 U13033 ( .A1(n18999), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19041) );
  NAND2_X1 U13034 ( .A1(n19072), .A2(n12706), .ZN(n19082) );
  AND2_X2 U13035 ( .A1(n12705), .A2(n13249), .ZN(n19072) );
  INV_X1 U13036 ( .A(n19074), .ZN(n19113) );
  OR2_X1 U13037 ( .A1(n19182), .A2(n19121), .ZN(n19149) );
  NAND2_X1 U13038 ( .A1(n19182), .A2(n19864), .ZN(n19173) );
  NAND2_X1 U13039 ( .A1(n19119), .A2(n19871), .ZN(n19182) );
  INV_X1 U13040 ( .A(n13178), .ZN(n19116) );
  AOI21_X1 U13041 ( .B1(n16086), .B2(n19201), .A(n12364), .ZN(n12368) );
  INV_X1 U13042 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n20775) );
  OR2_X1 U13043 ( .A1(n18882), .A2(n9743), .ZN(n19197) );
  NAND2_X1 U13044 ( .A1(n18882), .A2(n12360), .ZN(n16194) );
  INV_X1 U13045 ( .A(n14102), .ZN(n19038) );
  OR2_X1 U13046 ( .A1(n12352), .A2(n19854), .ZN(n19215) );
  INV_X1 U13047 ( .A(n19258), .ZN(n19250) );
  NAND2_X1 U13048 ( .A1(n19460), .A2(n19296), .ZN(n19289) );
  INV_X1 U13049 ( .A(n19319), .ZN(n19316) );
  INV_X1 U13050 ( .A(n19348), .ZN(n19346) );
  INV_X1 U13051 ( .A(n19401), .ZN(n19413) );
  INV_X1 U13052 ( .A(n19424), .ZN(n19432) );
  INV_X1 U13053 ( .A(n19448), .ZN(n19459) );
  INV_X1 U13054 ( .A(n19486), .ZN(n19484) );
  NAND2_X1 U13055 ( .A1(n19461), .A2(n19460), .ZN(n19521) );
  INV_X1 U13056 ( .A(n19540), .ZN(n19537) );
  INV_X1 U13057 ( .A(n19717), .ZN(n19571) );
  INV_X1 U13058 ( .A(n19597), .ZN(n19587) );
  NAND2_X1 U13059 ( .A1(n19461), .A2(n19604), .ZN(n19630) );
  INV_X1 U13060 ( .A(n19653), .ZN(n19703) );
  INV_X1 U13061 ( .A(n19718), .ZN(n19732) );
  INV_X1 U13062 ( .A(n19808), .ZN(n19742) );
  AND3_X1 U13063 ( .A1(n19747), .A2(n19797), .A3(n19754), .ZN(n19871) );
  AOI21_X1 U13064 ( .B1(n18681), .B2(n18680), .A(n17445), .ZN(n18868) );
  NAND2_X1 U13065 ( .A1(n18849), .A2(n18689), .ZN(n16439) );
  AOI211_X1 U13066 ( .C1(n16493), .C2(n16852), .A(n16482), .B(n16481), .ZN(
        n16483) );
  INV_X1 U13067 ( .A(n16457), .ZN(n16824) );
  INV_X1 U13068 ( .A(n16821), .ZN(n16804) );
  AND3_X1 U13069 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), 
        .A3(n16986), .ZN(n16976) );
  INV_X1 U13070 ( .A(n16980), .ZN(n16986) );
  INV_X1 U13071 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17232) );
  INV_X1 U13072 ( .A(n17316), .ZN(n17289) );
  NOR2_X1 U13073 ( .A1(n17425), .A2(n17348), .ZN(n17352) );
  NOR2_X1 U13074 ( .A1(n12820), .A2(n12819), .ZN(n17380) );
  INV_X1 U13075 ( .A(n17388), .ZN(n17242) );
  INV_X1 U13076 ( .A(n17408), .ZN(n17416) );
  NAND2_X1 U13077 ( .A1(n17410), .A2(n17442), .ZN(n17438) );
  INV_X1 U13078 ( .A(n17443), .ZN(n17442) );
  INV_X1 U13079 ( .A(n17505), .ZN(n17460) );
  NAND2_X1 U13080 ( .A1(n17448), .A2(n17460), .ZN(n17495) );
  AOI21_X1 U13081 ( .B1(n16334), .B2(n17783), .A(n13082), .ZN(n13083) );
  INV_X1 U13082 ( .A(n17658), .ZN(n17686) );
  NAND2_X1 U13083 ( .A1(n17362), .A2(n17818), .ZN(n17761) );
  INV_X1 U13084 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17841) );
  INV_X1 U13085 ( .A(n9717), .ZN(n18090) );
  INV_X1 U13086 ( .A(n18187), .ZN(n18165) );
  INV_X1 U13087 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n21027) );
  INV_X1 U13088 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18663) );
  INV_X1 U13089 ( .A(n18530), .ZN(n18603) );
  INV_X1 U13090 ( .A(n18805), .ZN(n18802) );
  INV_X1 U13091 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18744) );
  INV_X1 U13092 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18747) );
  INV_X1 U13093 ( .A(n18863), .ZN(n18842) );
  NOR2_X1 U13094 ( .A1(n18728), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18793) );
  INV_X1 U13095 ( .A(n16392), .ZN(n16397) );
  OAI21_X1 U13096 ( .B1(n14365), .B2(n14359), .A(n11894), .ZN(P1_U2843) );
  OR4_X1 U13097 ( .A1(n13115), .A2(n13114), .A3(n13113), .A4(n13112), .ZN(
        P2_U2840) );
  INV_X1 U13098 ( .A(n13083), .ZN(P3_U2799) );
  INV_X1 U13099 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12745) );
  NAND2_X1 U13100 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n10160), .ZN(
        n10159) );
  INV_X1 U13101 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15156) );
  INV_X1 U13102 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18918) );
  INV_X1 U13103 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14768) );
  INV_X1 U13104 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14737) );
  INV_X1 U13105 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10182) );
  INV_X1 U13106 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15059) );
  INV_X1 U13107 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10190) );
  INV_X1 U13108 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n15049) );
  INV_X1 U13109 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10154) );
  AOI21_X1 U13110 ( .B1(n18918), .B2(n10173), .A(n10175), .ZN(n18909) );
  AOI21_X1 U13111 ( .B1(n15156), .B2(n10171), .A(n10174), .ZN(n15155) );
  AOI21_X1 U13112 ( .B1(n20775), .B2(n10169), .A(n10170), .ZN(n16166) );
  AOI21_X1 U13113 ( .B1(n15188), .B2(n10167), .A(n9820), .ZN(n18959) );
  NAND2_X1 U13114 ( .A1(n10165), .A2(n15211), .ZN(n10157) );
  INV_X1 U13115 ( .A(n10168), .ZN(n10156) );
  AND2_X1 U13116 ( .A1(n10157), .A2(n10156), .ZN(n15213) );
  AOI21_X1 U13117 ( .B1(n16179), .B2(n10163), .A(n10166), .ZN(n18977) );
  AOI21_X1 U13118 ( .B1(n20789), .B2(n10161), .A(n10164), .ZN(n18988) );
  AOI21_X1 U13119 ( .B1(n20749), .B2(n10159), .A(n10162), .ZN(n19021) );
  AOI21_X1 U13120 ( .B1(n13767), .B2(n10158), .A(n10160), .ZN(n14845) );
  INV_X1 U13121 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15557) );
  INV_X1 U13122 ( .A(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n19039) );
  AOI22_X1 U13123 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15557), .B1(n19039), 
        .B2(n18874), .ZN(n14867) );
  INV_X1 U13124 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15558) );
  AOI22_X1 U13125 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15558), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18874), .ZN(n14866) );
  NOR2_X1 U13126 ( .A1(n14867), .A2(n14866), .ZN(n14865) );
  OAI21_X1 U13127 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n10158), .ZN(n14854) );
  NAND2_X1 U13128 ( .A1(n14865), .A2(n14854), .ZN(n14843) );
  NOR2_X1 U13129 ( .A1(n14845), .A2(n14843), .ZN(n14830) );
  OAI21_X1 U13130 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n10160), .A(
        n10159), .ZN(n19204) );
  NAND2_X1 U13131 ( .A1(n14830), .A2(n19204), .ZN(n19018) );
  NOR2_X1 U13132 ( .A1(n19021), .A2(n19018), .ZN(n19004) );
  OAI21_X1 U13133 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n10162), .A(
        n10161), .ZN(n19006) );
  NAND2_X1 U13134 ( .A1(n19004), .A2(n19006), .ZN(n18987) );
  NOR2_X1 U13135 ( .A1(n18988), .A2(n18987), .ZN(n14818) );
  OAI21_X1 U13136 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n10164), .A(
        n10163), .ZN(n15245) );
  NAND2_X1 U13137 ( .A1(n14818), .A2(n15245), .ZN(n18976) );
  NOR2_X1 U13138 ( .A1(n18977), .A2(n18976), .ZN(n14807) );
  OAI21_X1 U13139 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n10166), .A(
        n10165), .ZN(n15224) );
  NAND2_X1 U13140 ( .A1(n14807), .A2(n15224), .ZN(n13116) );
  NOR2_X1 U13141 ( .A1(n15213), .A2(n13116), .ZN(n18965) );
  OAI21_X1 U13142 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n10168), .A(
        n10167), .ZN(n18967) );
  NAND2_X1 U13143 ( .A1(n18965), .A2(n18967), .ZN(n18958) );
  NOR2_X1 U13144 ( .A1(n18959), .A2(n18958), .ZN(n18943) );
  OAI21_X1 U13145 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n9820), .A(
        n10169), .ZN(n18944) );
  NAND2_X1 U13146 ( .A1(n18943), .A2(n18944), .ZN(n13100) );
  NOR2_X1 U13147 ( .A1(n16166), .A2(n13100), .ZN(n18931) );
  OR2_X1 U13148 ( .A1(n10170), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10172) );
  NAND2_X1 U13149 ( .A1(n10172), .A2(n10171), .ZN(n18932) );
  NAND2_X1 U13150 ( .A1(n18931), .A2(n18932), .ZN(n18922) );
  NOR2_X1 U13151 ( .A1(n15155), .A2(n18922), .ZN(n14791) );
  OAI21_X1 U13152 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n10174), .A(
        n10173), .ZN(n16165) );
  NAND2_X1 U13153 ( .A1(n14791), .A2(n16165), .ZN(n18907) );
  OR2_X1 U13154 ( .A1(n18909), .A2(n18907), .ZN(n14775) );
  OAI21_X1 U13155 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n10175), .A(
        n10176), .ZN(n14776) );
  INV_X1 U13156 ( .A(n14776), .ZN(n15144) );
  NOR2_X1 U13157 ( .A1(n14775), .A2(n15144), .ZN(n14774) );
  INV_X1 U13158 ( .A(n14774), .ZN(n10178) );
  AND2_X1 U13159 ( .A1(n10176), .A2(n14768), .ZN(n10177) );
  OR2_X1 U13160 ( .A1(n10177), .A2(n9824), .ZN(n15135) );
  INV_X1 U13161 ( .A(n15135), .ZN(n14762) );
  OR2_X1 U13162 ( .A1(n9824), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10180) );
  NAND2_X1 U13163 ( .A1(n10179), .A2(n10180), .ZN(n15113) );
  NAND2_X1 U13164 ( .A1(n10179), .A2(n14737), .ZN(n10181) );
  NAND2_X1 U13165 ( .A1(n10183), .A2(n10181), .ZN(n15103) );
  NAND2_X1 U13166 ( .A1(n19019), .A2(n14731), .ZN(n16135) );
  AND2_X1 U13167 ( .A1(n10183), .A2(n10182), .ZN(n10184) );
  OR2_X1 U13168 ( .A1(n10184), .A2(n10185), .ZN(n16136) );
  NAND2_X1 U13169 ( .A1(n19019), .A2(n16134), .ZN(n16126) );
  NOR2_X1 U13170 ( .A1(n10185), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10186) );
  OR2_X1 U13171 ( .A1(n10187), .A2(n10186), .ZN(n16127) );
  NAND2_X1 U13172 ( .A1(n19019), .A2(n16125), .ZN(n16112) );
  OAI21_X1 U13173 ( .B1(n10187), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n10189), .ZN(n16113) );
  NAND2_X1 U13174 ( .A1(n19019), .A2(n16111), .ZN(n16100) );
  INV_X1 U13175 ( .A(n10191), .ZN(n10188) );
  AOI21_X1 U13176 ( .B1(n15059), .B2(n10189), .A(n10188), .ZN(n15062) );
  INV_X1 U13177 ( .A(n15062), .ZN(n16101) );
  NAND2_X1 U13178 ( .A1(n19019), .A2(n16099), .ZN(n16088) );
  NAND2_X1 U13179 ( .A1(n10191), .A2(n10190), .ZN(n10192) );
  NAND2_X1 U13180 ( .A1(n10193), .A2(n10192), .ZN(n16089) );
  NAND2_X1 U13181 ( .A1(n19019), .A2(n16087), .ZN(n16078) );
  AOI21_X1 U13182 ( .B1(n15049), .B2(n10193), .A(n10194), .ZN(n15052) );
  INV_X1 U13183 ( .A(n15052), .ZN(n16079) );
  NAND2_X1 U13184 ( .A1(n19019), .A2(n16077), .ZN(n10195) );
  XNOR2_X1 U13185 ( .A(n10194), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15039) );
  NOR3_X1 U13186 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15762) );
  NAND2_X1 U13187 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15762), .ZN(n19738) );
  INV_X2 U13188 ( .A(n19738), .ZN(n18915) );
  OAI211_X1 U13189 ( .C1(n10195), .C2(n15039), .A(n18915), .B(n16072), .ZN(
        n10920) );
  AND2_X2 U13190 ( .A1(n10196), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10238) );
  AOI22_X1 U13191 ( .A1(n10660), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9744), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10202) );
  AOI22_X1 U13192 ( .A1(n12539), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12690), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10201) );
  AND2_X4 U13193 ( .A1(n15579), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10661) );
  AOI22_X1 U13194 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12540), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10200) );
  AOI22_X1 U13195 ( .A1(n12550), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10199) );
  NAND4_X1 U13196 ( .A1(n10202), .A2(n10201), .A3(n10200), .A4(n10199), .ZN(
        n10203) );
  AOI22_X1 U13197 ( .A1(n10660), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10661), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10207) );
  AOI22_X1 U13198 ( .A1(n12539), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9761), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10206) );
  AOI22_X1 U13199 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9756), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10205) );
  AOI22_X1 U13200 ( .A1(n12550), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10204) );
  NAND4_X1 U13201 ( .A1(n10207), .A2(n10206), .A3(n10205), .A4(n10204), .ZN(
        n10208) );
  AOI22_X1 U13202 ( .A1(n10660), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12690), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10214) );
  AOI22_X1 U13203 ( .A1(n9745), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n10661), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10213) );
  AOI22_X1 U13204 ( .A1(n12539), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12540), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10212) );
  AOI22_X1 U13205 ( .A1(n12550), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10211) );
  NAND4_X1 U13206 ( .A1(n10214), .A2(n10213), .A3(n10212), .A4(n10211), .ZN(
        n10215) );
  AOI22_X1 U13207 ( .A1(n10660), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9744), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10219) );
  AOI22_X1 U13208 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12690), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10218) );
  AOI22_X1 U13209 ( .A1(n12539), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9756), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10217) );
  NAND4_X1 U13210 ( .A1(n10219), .A2(n10218), .A3(n10217), .A4(n10216), .ZN(
        n10220) );
  NOR2_X1 U13211 ( .A1(n11932), .A2(n12150), .ZN(n10233) );
  AOI22_X1 U13212 ( .A1(n10660), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9744), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10224) );
  AOI22_X1 U13213 ( .A1(n12539), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12690), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10223) );
  AOI22_X1 U13214 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12540), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10222) );
  AOI22_X1 U13215 ( .A1(n12550), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10221) );
  NAND4_X1 U13216 ( .A1(n10224), .A2(n10223), .A3(n10222), .A4(n10221), .ZN(
        n10225) );
  NAND2_X1 U13217 ( .A1(n10225), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10232) );
  AOI22_X1 U13218 ( .A1(n10660), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9744), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10229) );
  AOI22_X1 U13219 ( .A1(n12539), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12690), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10228) );
  AOI22_X1 U13220 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12540), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10227) );
  AOI22_X1 U13221 ( .A1(n12550), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10226) );
  NAND4_X1 U13222 ( .A1(n10229), .A2(n10228), .A3(n10227), .A4(n10226), .ZN(
        n10230) );
  NAND2_X1 U13223 ( .A1(n10230), .A2(n10809), .ZN(n10231) );
  NOR2_X1 U13224 ( .A1(n12707), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10266) );
  AOI222_X1 U13225 ( .A1(P2_REIP_REG_30__SCAN_IN), .A2(n10337), .B1(n12733), 
        .B2(P2_EAX_REG_30__SCAN_IN), .C1(n10267), .C2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10615) );
  AND2_X2 U13226 ( .A1(n10380), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10352) );
  AOI22_X1 U13227 ( .A1(n10352), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12465), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10237) );
  INV_X1 U13228 ( .A(n10287), .ZN(n12482) );
  NAND3_X1 U13229 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n16229), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12233) );
  AOI22_X1 U13230 ( .A1(n10287), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12525), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10236) );
  AOI22_X1 U13231 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12523), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10235) );
  INV_X1 U13232 ( .A(n10662), .ZN(n12541) );
  AOI22_X1 U13233 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12518), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10234) );
  NAND4_X1 U13234 ( .A1(n10237), .A2(n10236), .A3(n10235), .A4(n10234), .ZN(
        n10245) );
  AND2_X1 U13235 ( .A1(n10238), .A2(n12542), .ZN(n10292) );
  NOR2_X1 U13236 ( .A1(n14108), .A2(n16229), .ZN(n10239) );
  AOI22_X1 U13237 ( .A1(n10292), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10243) );
  AND2_X1 U13238 ( .A1(n12542), .A2(n15580), .ZN(n10442) );
  AND2_X1 U13239 ( .A1(n12542), .A2(n15569), .ZN(n10322) );
  AOI22_X1 U13240 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10322), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10242) );
  AND2_X2 U13241 ( .A1(n10660), .A2(n10809), .ZN(n10274) );
  AOI22_X1 U13242 ( .A1(n10366), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10274), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10241) );
  NAND4_X1 U13243 ( .A1(n10243), .A2(n10242), .A3(n10241), .A4(n10240), .ZN(
        n10244) );
  AND2_X1 U13244 ( .A1(n12150), .A2(n19385), .ZN(n10246) );
  AND2_X1 U13245 ( .A1(n10246), .A2(n19869), .ZN(n10314) );
  INV_X1 U13246 ( .A(n10314), .ZN(n10528) );
  AOI22_X1 U13247 ( .A1(n10660), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9745), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10250) );
  AOI22_X1 U13248 ( .A1(n12539), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12690), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10249) );
  AOI22_X1 U13249 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12540), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10248) );
  AOI22_X1 U13250 ( .A1(n12550), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10247) );
  NAND4_X1 U13251 ( .A1(n10250), .A2(n10249), .A3(n10248), .A4(n10247), .ZN(
        n10251) );
  NAND2_X1 U13252 ( .A1(n10251), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10258) );
  AOI22_X1 U13253 ( .A1(n10660), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9745), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10255) );
  AOI22_X1 U13254 ( .A1(n12539), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9746), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10254) );
  AOI22_X1 U13255 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12540), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n10253) );
  NAND4_X1 U13256 ( .A1(n10255), .A2(n10254), .A3(n10253), .A4(n10252), .ZN(
        n10256) );
  NAND2_X1 U13257 ( .A1(n10256), .A2(n10809), .ZN(n10257) );
  INV_X1 U13258 ( .A(n10721), .ZN(n10761) );
  NAND2_X2 U13259 ( .A1(n10761), .A2(n9740), .ZN(n10739) );
  NAND2_X1 U13260 ( .A1(n12706), .A2(n10267), .ZN(n10307) );
  INV_X1 U13261 ( .A(n10281), .ZN(n10259) );
  OAI21_X1 U13262 ( .B1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19385), .A(
        n10259), .ZN(n10260) );
  AND2_X1 U13263 ( .A1(n10307), .A2(n10260), .ZN(n10261) );
  INV_X2 U13264 ( .A(n10547), .ZN(n10337) );
  INV_X1 U13265 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18897) );
  AOI21_X1 U13266 ( .B1(n19254), .B2(P2_EAX_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10262) );
  AOI22_X1 U13267 ( .A1(n10266), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n10267), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10269) );
  NAND2_X1 U13268 ( .A1(n10337), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10268) );
  NAND2_X1 U13269 ( .A1(n10269), .A2(n10268), .ZN(n10284) );
  AOI22_X1 U13270 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n12517), .B1(
        n10366), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10273) );
  AOI22_X1 U13271 ( .A1(n12523), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n10368), .ZN(n10272) );
  AOI22_X1 U13272 ( .A1(n10287), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10367), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10271) );
  AOI22_X1 U13273 ( .A1(n10352), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n12525), .ZN(n10270) );
  NAND4_X1 U13274 ( .A1(n10273), .A2(n10272), .A3(n10271), .A4(n10270), .ZN(
        n10280) );
  AOI22_X1 U13275 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n10442), .B1(
        n10322), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10278) );
  AOI22_X1 U13276 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10292), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10277) );
  AOI22_X1 U13277 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n12518), .ZN(n10276) );
  AOI22_X1 U13278 ( .A1(n10274), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12465), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10275) );
  NAND4_X1 U13279 ( .A1(n10278), .A2(n10277), .A3(n10276), .A4(n10275), .ZN(
        n10279) );
  OR2_X1 U13280 ( .A1(n12310), .A2(n10528), .ZN(n10283) );
  AOI22_X1 U13281 ( .A1(n10739), .A2(n10281), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10282) );
  NAND2_X1 U13282 ( .A1(n10283), .A2(n10282), .ZN(n13340) );
  NOR2_X1 U13283 ( .A1(n13341), .A2(n13340), .ZN(n10286) );
  NOR2_X1 U13284 ( .A1(n13277), .A2(n10284), .ZN(n10285) );
  NOR2_X2 U13285 ( .A1(n10286), .A2(n10285), .ZN(n10312) );
  NAND2_X1 U13286 ( .A1(n10274), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n10290) );
  NAND2_X1 U13287 ( .A1(n10287), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10289) );
  NAND2_X1 U13288 ( .A1(n10352), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10288) );
  NAND3_X1 U13289 ( .A1(n10290), .A2(n10289), .A3(n10288), .ZN(n10291) );
  NOR2_X1 U13290 ( .A1(n10142), .A2(n10291), .ZN(n10306) );
  NAND2_X1 U13291 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10299) );
  NAND2_X1 U13292 ( .A1(n10366), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10298) );
  AOI22_X1 U13293 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10442), .B1(
        n10322), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10297) );
  INV_X1 U13294 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10294) );
  NAND2_X1 U13295 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n12525), .ZN(
        n10293) );
  OAI21_X1 U13296 ( .B1(n12528), .B2(n10294), .A(n10293), .ZN(n10295) );
  AOI21_X1 U13297 ( .B1(n10292), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n10295), .ZN(n10296) );
  NAND2_X1 U13298 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10303) );
  AOI22_X1 U13299 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10302) );
  NAND2_X1 U13300 ( .A1(n12518), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10301) );
  NAND2_X1 U13301 ( .A1(n12465), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10300) );
  NAND2_X1 U13302 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10308) );
  OAI211_X1 U13303 ( .C1(n10528), .C2(n12313), .A(n10308), .B(n10307), .ZN(
        n10311) );
  XNOR2_X1 U13304 ( .A(n10312), .B(n10311), .ZN(n13284) );
  AOI22_X1 U13305 ( .A1(n12733), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n10267), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10310) );
  NAND2_X1 U13306 ( .A1(n10337), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10309) );
  NAND2_X1 U13307 ( .A1(n10310), .A2(n10309), .ZN(n13283) );
  NOR2_X1 U13308 ( .A1(n13284), .A2(n13283), .ZN(n13285) );
  NOR2_X1 U13309 ( .A1(n10312), .A2(n10311), .ZN(n10313) );
  NOR2_X2 U13310 ( .A1(n13285), .A2(n10313), .ZN(n13774) );
  NAND2_X1 U13311 ( .A1(n10337), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U13312 ( .A1(n10267), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n10335) );
  INV_X1 U13313 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10316) );
  INV_X1 U13314 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10315) );
  OAI22_X1 U13315 ( .A1(n10393), .A2(n10316), .B1(n10392), .B2(n10315), .ZN(
        n10321) );
  INV_X1 U13316 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10319) );
  NAND2_X1 U13317 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n10318) );
  NAND2_X1 U13318 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10317) );
  OAI211_X1 U13319 ( .C1(n12497), .C2(n10319), .A(n10318), .B(n10317), .ZN(
        n10320) );
  NOR2_X1 U13320 ( .A1(n10321), .A2(n10320), .ZN(n10332) );
  NAND2_X1 U13321 ( .A1(n10366), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10328) );
  NAND2_X1 U13322 ( .A1(n12523), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n10327) );
  AOI22_X1 U13323 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10292), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10326) );
  INV_X1 U13324 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10323) );
  INV_X1 U13325 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n20820) );
  OAI22_X1 U13326 ( .A1(n12528), .A2(n10323), .B1(n10570), .B2(n20820), .ZN(
        n10324) );
  AOI21_X1 U13327 ( .B1(n10322), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A(
        n10324), .ZN(n10325) );
  AOI22_X1 U13328 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10274), .B1(
        n12534), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10330) );
  AOI22_X1 U13329 ( .A1(n10352), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n10287), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10329) );
  NAND4_X1 U13330 ( .A1(n10332), .A2(n10331), .A3(n10330), .A4(n10329), .ZN(
        n11933) );
  NAND2_X1 U13331 ( .A1(n9757), .A2(n11933), .ZN(n10334) );
  NAND2_X1 U13332 ( .A1(n12733), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n10333) );
  NAND4_X1 U13333 ( .A1(n10336), .A2(n10335), .A3(n10334), .A4(n10333), .ZN(
        n13773) );
  NAND2_X1 U13334 ( .A1(n13774), .A2(n13773), .ZN(n13775) );
  AOI22_X1 U13335 ( .A1(n12733), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n10267), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10361) );
  NAND2_X1 U13336 ( .A1(n10337), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n10360) );
  INV_X1 U13337 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10339) );
  INV_X1 U13338 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10338) );
  OAI22_X1 U13339 ( .A1(n10393), .A2(n10339), .B1(n10392), .B2(n10338), .ZN(
        n10344) );
  INV_X1 U13340 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10342) );
  NAND2_X1 U13341 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n10341) );
  NAND2_X1 U13342 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10340) );
  OAI211_X1 U13343 ( .C1(n12497), .C2(n10342), .A(n10341), .B(n10340), .ZN(
        n10343) );
  NOR2_X1 U13344 ( .A1(n10344), .A2(n10343), .ZN(n10358) );
  NAND2_X1 U13345 ( .A1(n10366), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10351) );
  NAND2_X1 U13346 ( .A1(n12523), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10350) );
  AOI22_X1 U13347 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10292), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10349) );
  INV_X1 U13348 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10346) );
  NAND2_X1 U13349 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12525), .ZN(
        n10345) );
  OAI21_X1 U13350 ( .B1(n12528), .B2(n10346), .A(n10345), .ZN(n10347) );
  AOI21_X1 U13351 ( .B1(n10322), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A(
        n10347), .ZN(n10348) );
  AOI22_X1 U13352 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10274), .B1(
        n12534), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10356) );
  INV_X1 U13353 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n20894) );
  INV_X1 U13354 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10353) );
  OAI22_X1 U13355 ( .A1(n12484), .A2(n20894), .B1(n12482), .B2(n10353), .ZN(
        n10354) );
  INV_X1 U13356 ( .A(n10354), .ZN(n10355) );
  NAND2_X1 U13357 ( .A1(n9757), .A2(n12306), .ZN(n10359) );
  AOI22_X1 U13358 ( .A1(n12733), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n10267), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10390) );
  NAND2_X1 U13359 ( .A1(n10337), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n10389) );
  NAND2_X1 U13360 ( .A1(n12523), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10365) );
  NAND2_X1 U13361 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n10364) );
  NAND2_X1 U13362 ( .A1(n10274), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n10363) );
  NAND2_X1 U13363 ( .A1(n10287), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n10362) );
  NAND4_X1 U13364 ( .A1(n10365), .A2(n10364), .A3(n10363), .A4(n10362), .ZN(
        n10379) );
  INV_X1 U13365 ( .A(n10366), .ZN(n10377) );
  INV_X1 U13366 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10376) );
  AOI22_X1 U13367 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10322), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10375) );
  INV_X1 U13368 ( .A(n10367), .ZN(n10372) );
  INV_X1 U13369 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10371) );
  NAND2_X1 U13370 ( .A1(n12524), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10370) );
  AOI22_X1 U13371 ( .A1(n10368), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12525), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10369) );
  OAI211_X1 U13372 ( .C1(n10372), .C2(n10371), .A(n10370), .B(n10369), .ZN(
        n10373) );
  INV_X1 U13373 ( .A(n10373), .ZN(n10374) );
  OAI211_X1 U13374 ( .C1(n10377), .C2(n10376), .A(n10375), .B(n10374), .ZN(
        n10378) );
  NOR2_X1 U13375 ( .A1(n10379), .A2(n10378), .ZN(n10386) );
  AOI22_X1 U13376 ( .A1(n12518), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12465), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10384) );
  INV_X1 U13377 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n20959) );
  NOR2_X1 U13378 ( .A1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n20959), .ZN(
        n20989) );
  NAND2_X1 U13379 ( .A1(n20989), .A2(n10380), .ZN(n10383) );
  NAND2_X1 U13380 ( .A1(n10352), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10382) );
  NAND2_X1 U13381 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10381) );
  INV_X1 U13382 ( .A(n12016), .ZN(n10387) );
  NAND2_X1 U13383 ( .A1(n9757), .A2(n10387), .ZN(n10388) );
  NAND3_X1 U13384 ( .A1(n10390), .A2(n10389), .A3(n10388), .ZN(n13973) );
  INV_X1 U13385 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12033) );
  INV_X1 U13386 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10391) );
  OAI22_X1 U13387 ( .A1(n10393), .A2(n12033), .B1(n10392), .B2(n10391), .ZN(
        n10398) );
  INV_X1 U13388 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10396) );
  NAND2_X1 U13389 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n10395) );
  NAND2_X1 U13390 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n10394) );
  OAI211_X1 U13391 ( .C1(n10396), .C2(n12497), .A(n10395), .B(n10394), .ZN(
        n10397) );
  NOR2_X1 U13392 ( .A1(n10398), .A2(n10397), .ZN(n10411) );
  NAND2_X1 U13393 ( .A1(n10366), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10404) );
  NAND2_X1 U13394 ( .A1(n12523), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n10403) );
  AOI22_X1 U13395 ( .A1(n10292), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10402) );
  INV_X1 U13396 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19249) );
  NAND2_X1 U13397 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n12525), .ZN(
        n10399) );
  OAI21_X1 U13398 ( .B1(n19249), .B2(n12528), .A(n10399), .ZN(n10400) );
  AOI21_X1 U13399 ( .B1(n10322), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A(
        n10400), .ZN(n10401) );
  AOI22_X1 U13400 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10274), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10409) );
  INV_X1 U13401 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10406) );
  INV_X1 U13402 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10405) );
  OAI22_X1 U13403 ( .A1(n12484), .A2(n10406), .B1(n12482), .B2(n10405), .ZN(
        n10407) );
  INV_X1 U13404 ( .A(n10407), .ZN(n10408) );
  NAND4_X1 U13405 ( .A1(n10411), .A2(n10410), .A3(n10409), .A4(n10408), .ZN(
        n12041) );
  NAND2_X1 U13406 ( .A1(n9757), .A2(n12041), .ZN(n10412) );
  AOI22_X1 U13407 ( .A1(n12733), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n10267), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10414) );
  NAND2_X1 U13408 ( .A1(n10337), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n10413) );
  NAND2_X1 U13409 ( .A1(n10414), .A2(n10413), .ZN(n15543) );
  NAND2_X1 U13410 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10418) );
  NAND2_X1 U13411 ( .A1(n10274), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10417) );
  NAND2_X1 U13412 ( .A1(n10352), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10416) );
  NAND2_X1 U13413 ( .A1(n10287), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10415) );
  NAND2_X1 U13414 ( .A1(n10366), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10425) );
  NAND2_X1 U13415 ( .A1(n12523), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10424) );
  AOI22_X1 U13416 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10292), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10423) );
  INV_X1 U13417 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10420) );
  INV_X1 U13418 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10419) );
  OAI22_X1 U13419 ( .A1(n12528), .A2(n10420), .B1(n10570), .B2(n10419), .ZN(
        n10421) );
  AOI21_X1 U13420 ( .B1(n10322), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A(
        n10421), .ZN(n10422) );
  NAND2_X1 U13421 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10429) );
  AOI22_X1 U13422 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10428) );
  NAND2_X1 U13423 ( .A1(n12518), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10427) );
  NAND2_X1 U13424 ( .A1(n12465), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10426) );
  AND3_X2 U13425 ( .A1(n10432), .A2(n10431), .A3(n10430), .ZN(n12158) );
  NAND2_X1 U13426 ( .A1(n9757), .A2(n12762), .ZN(n10433) );
  AOI22_X1 U13427 ( .A1(n12733), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n10267), .B2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10436) );
  NAND2_X1 U13428 ( .A1(n10337), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n10435) );
  NAND2_X1 U13429 ( .A1(n10436), .A2(n10435), .ZN(n15531) );
  AOI22_X1 U13430 ( .A1(n12733), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n10267), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10458) );
  NAND2_X1 U13431 ( .A1(n10337), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10457) );
  INV_X1 U13432 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10437) );
  OR2_X1 U13433 ( .A1(n12481), .A2(n10437), .ZN(n10441) );
  NAND2_X1 U13434 ( .A1(n10274), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n10440) );
  NAND2_X1 U13435 ( .A1(n10287), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n10439) );
  NAND2_X1 U13436 ( .A1(n10352), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n10438) );
  AND4_X1 U13437 ( .A1(n10441), .A2(n10440), .A3(n10439), .A4(n10438), .ZN(
        n10454) );
  NAND2_X1 U13438 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10446) );
  AOI22_X1 U13439 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10445) );
  NAND2_X1 U13440 ( .A1(n12518), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10444) );
  NAND2_X1 U13441 ( .A1(n12465), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n10443) );
  AND4_X1 U13442 ( .A1(n10446), .A2(n10445), .A3(n10444), .A4(n10443), .ZN(
        n10453) );
  NAND2_X1 U13443 ( .A1(n10366), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n10452) );
  NAND2_X1 U13444 ( .A1(n12523), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n10451) );
  AOI22_X1 U13445 ( .A1(n10292), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10450) );
  INV_X1 U13446 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n20792) );
  NAND2_X1 U13447 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n12525), .ZN(
        n10447) );
  OAI21_X1 U13448 ( .B1(n12528), .B2(n20792), .A(n10447), .ZN(n10448) );
  AOI21_X1 U13449 ( .B1(n10322), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n10448), .ZN(n10449) );
  INV_X1 U13450 ( .A(n13633), .ZN(n10455) );
  NAND2_X1 U13451 ( .A1(n9757), .A2(n10455), .ZN(n10456) );
  AOI22_X1 U13452 ( .A1(n12733), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n10267), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10475) );
  NAND2_X1 U13453 ( .A1(n10337), .A2(P2_REIP_REG_9__SCAN_IN), .ZN(n10474) );
  NAND2_X1 U13454 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10462) );
  AOI22_X1 U13455 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10461) );
  NAND2_X1 U13456 ( .A1(n12518), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n10460) );
  NAND2_X1 U13457 ( .A1(n12465), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n10459) );
  AND4_X1 U13458 ( .A1(n10462), .A2(n10461), .A3(n10460), .A4(n10459), .ZN(
        n10472) );
  NAND2_X1 U13459 ( .A1(n10366), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10468) );
  NAND2_X1 U13460 ( .A1(n10352), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n10467) );
  AOI22_X1 U13461 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10322), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10466) );
  INV_X1 U13462 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11941) );
  NAND2_X1 U13463 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n12525), .ZN(
        n10463) );
  OAI21_X1 U13464 ( .B1(n12528), .B2(n11941), .A(n10463), .ZN(n10464) );
  AOI21_X1 U13465 ( .B1(n10292), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A(
        n10464), .ZN(n10465) );
  AND4_X1 U13466 ( .A1(n10468), .A2(n10467), .A3(n10466), .A4(n10465), .ZN(
        n10471) );
  AOI22_X1 U13467 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10274), .B1(
        n12523), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10470) );
  AOI22_X1 U13468 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n10287), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10469) );
  NAND4_X1 U13469 ( .A1(n10472), .A2(n10471), .A3(n10470), .A4(n10469), .ZN(
        n12402) );
  NAND2_X1 U13470 ( .A1(n9757), .A2(n12402), .ZN(n10473) );
  NAND3_X1 U13471 ( .A1(n10475), .A2(n10474), .A3(n10473), .ZN(n15513) );
  AOI22_X1 U13472 ( .A1(n12733), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n10267), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n10493) );
  NAND2_X1 U13473 ( .A1(n10337), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n10492) );
  NAND2_X1 U13474 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n10479) );
  AOI22_X1 U13475 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10478) );
  NAND2_X1 U13476 ( .A1(n12518), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10477) );
  NAND2_X1 U13477 ( .A1(n12465), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10476) );
  AND4_X1 U13478 ( .A1(n10479), .A2(n10478), .A3(n10477), .A4(n10476), .ZN(
        n10490) );
  NAND2_X1 U13479 ( .A1(n10366), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10486) );
  NAND2_X1 U13480 ( .A1(n12523), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10485) );
  INV_X1 U13481 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n20910) );
  AOI22_X1 U13482 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n10292), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10484) );
  INV_X1 U13483 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10481) );
  NAND2_X1 U13484 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n12525), .ZN(
        n10480) );
  OAI21_X1 U13485 ( .B1(n12528), .B2(n10481), .A(n10480), .ZN(n10482) );
  AOI21_X1 U13486 ( .B1(n10322), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A(
        n10482), .ZN(n10483) );
  AND4_X1 U13487 ( .A1(n10486), .A2(n10485), .A3(n10484), .A4(n10483), .ZN(
        n10489) );
  AOI22_X1 U13488 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n10274), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10488) );
  AOI22_X1 U13489 ( .A1(n10352), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10287), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10487) );
  NAND4_X1 U13490 ( .A1(n10490), .A2(n10489), .A3(n10488), .A4(n10487), .ZN(
        n13681) );
  NAND2_X1 U13491 ( .A1(n9757), .A2(n13681), .ZN(n10491) );
  AOI22_X1 U13492 ( .A1(n12733), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n10267), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10511) );
  NAND2_X1 U13493 ( .A1(n10337), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n10510) );
  NAND2_X1 U13494 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n10497) );
  AOI22_X1 U13495 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10496) );
  NAND2_X1 U13496 ( .A1(n12518), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n10495) );
  NAND2_X1 U13497 ( .A1(n12465), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10494) );
  AND4_X1 U13498 ( .A1(n10497), .A2(n10496), .A3(n10495), .A4(n10494), .ZN(
        n10508) );
  NAND2_X1 U13499 ( .A1(n10352), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10504) );
  NAND2_X1 U13500 ( .A1(n10366), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n10503) );
  AOI22_X1 U13501 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10322), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10502) );
  INV_X1 U13502 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10499) );
  NAND2_X1 U13503 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n12525), .ZN(
        n10498) );
  OAI21_X1 U13504 ( .B1(n12528), .B2(n10499), .A(n10498), .ZN(n10500) );
  AOI21_X1 U13505 ( .B1(n10292), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n10500), .ZN(n10501) );
  AND4_X1 U13506 ( .A1(n10504), .A2(n10503), .A3(n10502), .A4(n10501), .ZN(
        n10507) );
  AOI22_X1 U13507 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12523), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10506) );
  AOI22_X1 U13508 ( .A1(n10274), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10287), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10505) );
  NAND4_X1 U13509 ( .A1(n10508), .A2(n10507), .A3(n10506), .A4(n10505), .ZN(
        n13684) );
  NAND2_X1 U13510 ( .A1(n9757), .A2(n13684), .ZN(n10509) );
  NAND3_X1 U13511 ( .A1(n10511), .A2(n10510), .A3(n10509), .ZN(n13117) );
  NAND2_X1 U13512 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10515) );
  AOI22_X1 U13513 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10514) );
  NAND2_X1 U13514 ( .A1(n12518), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n10513) );
  NAND2_X1 U13515 ( .A1(n12465), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10512) );
  AND4_X1 U13516 ( .A1(n10515), .A2(n10514), .A3(n10513), .A4(n10512), .ZN(
        n10526) );
  NAND2_X1 U13517 ( .A1(n10366), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n10522) );
  NAND2_X1 U13518 ( .A1(n12523), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10521) );
  AOI22_X1 U13519 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10292), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10520) );
  INV_X1 U13520 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10517) );
  NAND2_X1 U13521 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12525), .ZN(
        n10516) );
  OAI21_X1 U13522 ( .B1(n12528), .B2(n10517), .A(n10516), .ZN(n10518) );
  AOI21_X1 U13523 ( .B1(n10322), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A(
        n10518), .ZN(n10519) );
  AND4_X1 U13524 ( .A1(n10522), .A2(n10521), .A3(n10520), .A4(n10519), .ZN(
        n10525) );
  AOI22_X1 U13525 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10274), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10524) );
  AOI22_X1 U13526 ( .A1(n10352), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10287), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10523) );
  NAND4_X1 U13527 ( .A1(n10526), .A2(n10525), .A3(n10524), .A4(n10523), .ZN(
        n12404) );
  INV_X1 U13528 ( .A(n12404), .ZN(n13727) );
  AOI22_X1 U13529 ( .A1(n12733), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n10267), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n10527) );
  OAI21_X1 U13530 ( .B1(n10528), .B2(n13727), .A(n10527), .ZN(n10529) );
  AOI21_X1 U13531 ( .B1(P2_REIP_REG_12__SCAN_IN), .B2(n10337), .A(n10529), 
        .ZN(n16196) );
  NOR2_X2 U13532 ( .A1(n16195), .A2(n16196), .ZN(n15480) );
  INV_X1 U13533 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n15187) );
  AOI22_X1 U13534 ( .A1(n12733), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n10267), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10546) );
  AOI22_X1 U13535 ( .A1(n12518), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12465), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10533) );
  NAND2_X1 U13536 ( .A1(n20989), .A2(n12690), .ZN(n10532) );
  NAND2_X1 U13537 ( .A1(n10274), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n10531) );
  NAND2_X1 U13538 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10530) );
  AND4_X1 U13539 ( .A1(n10533), .A2(n10532), .A3(n10531), .A4(n10530), .ZN(
        n10544) );
  NAND2_X1 U13540 ( .A1(n10352), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10540) );
  AOI22_X1 U13541 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10322), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10539) );
  INV_X1 U13542 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10535) );
  NAND2_X1 U13543 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n12525), .ZN(
        n10534) );
  OAI21_X1 U13544 ( .B1(n12528), .B2(n10535), .A(n10534), .ZN(n10536) );
  AOI21_X1 U13545 ( .B1(n10292), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A(
        n10536), .ZN(n10538) );
  NAND2_X1 U13546 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n10537) );
  AND4_X1 U13547 ( .A1(n10540), .A2(n10539), .A3(n10538), .A4(n10537), .ZN(
        n10543) );
  AOI22_X1 U13548 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n10366), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10542) );
  AOI22_X1 U13549 ( .A1(n12523), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n10287), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10541) );
  NAND4_X1 U13550 ( .A1(n10544), .A2(n10543), .A3(n10542), .A4(n10541), .ZN(
        n13730) );
  NAND2_X1 U13551 ( .A1(n9757), .A2(n13730), .ZN(n10545) );
  OAI211_X1 U13552 ( .C1(n10547), .C2(n15187), .A(n10546), .B(n10545), .ZN(
        n15481) );
  NAND2_X1 U13553 ( .A1(n15480), .A2(n15481), .ZN(n15464) );
  AOI22_X1 U13554 ( .A1(n12733), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n10267), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n10565) );
  NAND2_X1 U13555 ( .A1(n10337), .A2(P2_REIP_REG_14__SCAN_IN), .ZN(n10564) );
  NAND2_X1 U13556 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n10551) );
  AOI22_X1 U13557 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10550) );
  NAND2_X1 U13558 ( .A1(n12518), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n10549) );
  NAND2_X1 U13559 ( .A1(n12465), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n10548) );
  AND4_X1 U13560 ( .A1(n10551), .A2(n10550), .A3(n10549), .A4(n10548), .ZN(
        n10562) );
  NAND2_X1 U13561 ( .A1(n10366), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n10558) );
  NAND2_X1 U13562 ( .A1(n12523), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10557) );
  AOI22_X1 U13563 ( .A1(n10292), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10556) );
  INV_X1 U13564 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10553) );
  NAND2_X1 U13565 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n12525), .ZN(
        n10552) );
  OAI21_X1 U13566 ( .B1(n12528), .B2(n10553), .A(n10552), .ZN(n10554) );
  AOI21_X1 U13567 ( .B1(n10322), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A(
        n10554), .ZN(n10555) );
  AND4_X1 U13568 ( .A1(n10558), .A2(n10557), .A3(n10556), .A4(n10555), .ZN(
        n10561) );
  AOI22_X1 U13569 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10274), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10560) );
  AOI22_X1 U13570 ( .A1(n10352), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10287), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10559) );
  NAND4_X1 U13571 ( .A1(n10562), .A2(n10561), .A3(n10560), .A4(n10559), .ZN(
        n13791) );
  NAND2_X1 U13572 ( .A1(n9757), .A2(n13791), .ZN(n10563) );
  NOR2_X2 U13573 ( .A1(n15464), .A2(n15465), .ZN(n13107) );
  AOI22_X1 U13574 ( .A1(n12733), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n10267), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n10584) );
  NAND2_X1 U13575 ( .A1(n10337), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n10583) );
  NAND2_X1 U13576 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10569) );
  AOI22_X1 U13577 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10568) );
  NAND2_X1 U13578 ( .A1(n12465), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10567) );
  NAND2_X1 U13579 ( .A1(n12518), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10566) );
  AND4_X1 U13580 ( .A1(n10569), .A2(n10568), .A3(n10567), .A4(n10566), .ZN(
        n10581) );
  NAND2_X1 U13581 ( .A1(n12523), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10577) );
  NAND2_X1 U13582 ( .A1(n10366), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10576) );
  AOI22_X1 U13583 ( .A1(n10442), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10322), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10575) );
  INV_X1 U13584 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n10572) );
  INV_X1 U13585 ( .A(n10570), .ZN(n12525) );
  NAND2_X1 U13586 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n12525), .ZN(
        n10571) );
  OAI21_X1 U13587 ( .B1(n12528), .B2(n10572), .A(n10571), .ZN(n10573) );
  AOI21_X1 U13588 ( .B1(n10292), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n10573), .ZN(n10574) );
  AND4_X1 U13589 ( .A1(n10577), .A2(n10576), .A3(n10575), .A4(n10574), .ZN(
        n10580) );
  AOI22_X1 U13590 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10274), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10579) );
  AOI22_X1 U13591 ( .A1(n10352), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10287), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10578) );
  NAND4_X1 U13592 ( .A1(n10581), .A2(n10580), .A3(n10579), .A4(n10578), .ZN(
        n13856) );
  NAND2_X1 U13593 ( .A1(n9757), .A2(n13856), .ZN(n10582) );
  INV_X1 U13594 ( .A(n13108), .ZN(n10585) );
  AOI22_X1 U13595 ( .A1(n12733), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n10267), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n10587) );
  NAND2_X1 U13596 ( .A1(n10337), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n10586) );
  AND2_X1 U13597 ( .A1(n10587), .A2(n10586), .ZN(n13984) );
  AOI22_X1 U13598 ( .A1(n12733), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n10267), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10589) );
  NAND2_X1 U13599 ( .A1(n10337), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n10588) );
  NAND2_X1 U13600 ( .A1(n10589), .A2(n10588), .ZN(n14002) );
  AOI22_X1 U13601 ( .A1(n12733), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n10267), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n10591) );
  NAND2_X1 U13602 ( .A1(n10337), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n10590) );
  AND2_X1 U13603 ( .A1(n10591), .A2(n10590), .ZN(n14797) );
  AOI22_X1 U13604 ( .A1(n12733), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n10267), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n10593) );
  NAND2_X1 U13605 ( .A1(n10337), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n10592) );
  NAND2_X1 U13606 ( .A1(n10593), .A2(n10592), .ZN(n15015) );
  AOI22_X1 U13607 ( .A1(n12733), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n10267), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n10595) );
  NAND2_X1 U13608 ( .A1(n10337), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n10594) );
  AND2_X1 U13609 ( .A1(n10595), .A2(n10594), .ZN(n14780) );
  AOI22_X1 U13610 ( .A1(n12733), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n10267), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10597) );
  NAND2_X1 U13611 ( .A1(n10337), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n10596) );
  NAND2_X1 U13612 ( .A1(n10597), .A2(n10596), .ZN(n14765) );
  NAND2_X1 U13613 ( .A1(n14764), .A2(n14765), .ZN(n14748) );
  AOI22_X1 U13614 ( .A1(n12733), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n10267), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10599) );
  NAND2_X1 U13615 ( .A1(n10337), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n10598) );
  AND2_X1 U13616 ( .A1(n10599), .A2(n10598), .ZN(n14746) );
  NOR2_X2 U13617 ( .A1(n14748), .A2(n14746), .ZN(n14733) );
  AOI22_X1 U13618 ( .A1(n12733), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n10267), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10601) );
  NAND2_X1 U13619 ( .A1(n10337), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n10600) );
  NAND2_X1 U13620 ( .A1(n10601), .A2(n10600), .ZN(n14734) );
  NAND2_X1 U13621 ( .A1(n14733), .A2(n14734), .ZN(n14735) );
  AOI22_X1 U13622 ( .A1(n12733), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n10267), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10603) );
  NAND2_X1 U13623 ( .A1(n10337), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n10602) );
  AND2_X1 U13624 ( .A1(n10603), .A2(n10602), .ZN(n15326) );
  AOI22_X1 U13625 ( .A1(n12733), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n10267), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10605) );
  NAND2_X1 U13626 ( .A1(n10337), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n10604) );
  AND2_X1 U13627 ( .A1(n10605), .A2(n10604), .ZN(n14991) );
  AOI22_X1 U13628 ( .A1(n12733), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n10267), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10607) );
  NAND2_X1 U13629 ( .A1(n10337), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n10606) );
  NAND2_X1 U13630 ( .A1(n10607), .A2(n10606), .ZN(n14986) );
  AOI22_X1 U13631 ( .A1(n12733), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n10267), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n10609) );
  NAND2_X1 U13632 ( .A1(n10337), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n10608) );
  AND2_X1 U13633 ( .A1(n10609), .A2(n10608), .ZN(n14979) );
  AOI22_X1 U13634 ( .A1(n12733), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n10267), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10611) );
  NAND2_X1 U13635 ( .A1(n10337), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n10610) );
  AND2_X1 U13636 ( .A1(n10611), .A2(n10610), .ZN(n12294) );
  AOI22_X1 U13637 ( .A1(n12733), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n10267), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10613) );
  NAND2_X1 U13638 ( .A1(n10337), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n10612) );
  NAND2_X1 U13639 ( .A1(n10613), .A2(n10612), .ZN(n14968) );
  AOI21_X1 U13640 ( .B1(n10615), .B2(n10614), .A(n12736), .ZN(n15260) );
  AOI22_X1 U13641 ( .A1(n12539), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12690), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10620) );
  NAND2_X1 U13642 ( .A1(n10662), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10616) );
  AOI22_X1 U13643 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12540), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10618) );
  NAND4_X1 U13644 ( .A1(n10621), .A2(n10620), .A3(n10619), .A4(n10618), .ZN(
        n10622) );
  NAND2_X1 U13645 ( .A1(n10622), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10629) );
  AOI22_X1 U13646 ( .A1(n10660), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9744), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10626) );
  AOI22_X1 U13647 ( .A1(n12539), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9746), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10625) );
  AOI22_X1 U13648 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12540), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10624) );
  AOI22_X1 U13649 ( .A1(n12550), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10623) );
  NAND4_X1 U13650 ( .A1(n10626), .A2(n10625), .A3(n10624), .A4(n10623), .ZN(
        n10627) );
  NAND2_X1 U13651 ( .A1(n10627), .A2(n10809), .ZN(n10628) );
  AOI22_X1 U13652 ( .A1(n12539), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n9761), .ZN(n10633) );
  AOI22_X1 U13653 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12540), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10632) );
  AOI22_X1 U13654 ( .A1(n12550), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10631) );
  NAND4_X1 U13655 ( .A1(n10634), .A2(n10633), .A3(n10632), .A4(n10631), .ZN(
        n10635) );
  NAND2_X1 U13656 ( .A1(n10635), .A2(n10809), .ZN(n10642) );
  AOI22_X1 U13657 ( .A1(n12539), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9746), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10638) );
  AOI22_X1 U13658 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9756), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10637) );
  NAND4_X1 U13659 ( .A1(n10639), .A2(n10638), .A3(n10637), .A4(n10636), .ZN(
        n10640) );
  NAND2_X1 U13660 ( .A1(n10640), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10641) );
  AOI22_X1 U13661 ( .A1(n12539), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9761), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10645) );
  AOI22_X1 U13662 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12540), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10644) );
  AOI22_X1 U13663 ( .A1(n12550), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10643) );
  NAND4_X1 U13664 ( .A1(n10646), .A2(n10645), .A3(n10644), .A4(n10643), .ZN(
        n10647) );
  NAND2_X1 U13665 ( .A1(n10647), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10654) );
  AOI22_X1 U13666 ( .A1(n12539), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12690), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10650) );
  AOI22_X1 U13667 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9756), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10649) );
  AOI22_X1 U13668 ( .A1(n12550), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10648) );
  NAND4_X1 U13669 ( .A1(n10651), .A2(n10650), .A3(n10649), .A4(n10648), .ZN(
        n10652) );
  NAND2_X1 U13670 ( .A1(n10652), .A2(n10809), .ZN(n10653) );
  AOI22_X1 U13671 ( .A1(n10660), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10661), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10658) );
  AOI22_X1 U13672 ( .A1(n12539), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n9761), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10657) );
  AOI22_X1 U13673 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(n9756), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10656) );
  AOI22_X1 U13674 ( .A1(n12550), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10655) );
  NAND4_X1 U13675 ( .A1(n10658), .A2(n10657), .A3(n10656), .A4(n10655), .ZN(
        n10659) );
  AOI22_X1 U13676 ( .A1(n12539), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10660), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10666) );
  AOI22_X1 U13677 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9761), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10665) );
  AOI22_X1 U13678 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9756), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10664) );
  AOI22_X1 U13679 ( .A1(n12550), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10662), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10663) );
  NAND4_X1 U13680 ( .A1(n10666), .A2(n10665), .A3(n10664), .A4(n10663), .ZN(
        n10667) );
  NAND2_X1 U13681 ( .A1(n10667), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10668) );
  NAND2_X1 U13682 ( .A1(n16287), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19741) );
  NOR2_X1 U13683 ( .A1(n10760), .A2(n18880), .ZN(n10688) );
  MUX2_X1 U13684 ( .A(n10670), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        n16229), .Z(n12204) );
  NAND2_X1 U13685 ( .A1(n12204), .A2(n11976), .ZN(n10672) );
  NAND2_X1 U13686 ( .A1(n10670), .A2(n16229), .ZN(n10671) );
  NAND2_X1 U13687 ( .A1(n10672), .A2(n10671), .ZN(n10681) );
  MUX2_X1 U13688 ( .A(n12371), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n10680) );
  NAND2_X1 U13689 ( .A1(n10681), .A2(n10680), .ZN(n10674) );
  NAND2_X1 U13690 ( .A1(n12371), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10673) );
  NAND2_X1 U13691 ( .A1(n10674), .A2(n10673), .ZN(n10679) );
  NOR2_X1 U13692 ( .A1(n10809), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n10675) );
  NOR2_X1 U13693 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15764), .ZN(
        n10676) );
  NAND2_X1 U13694 ( .A1(n10684), .A2(n10676), .ZN(n10705) );
  INV_X1 U13695 ( .A(n10677), .ZN(n10678) );
  XNOR2_X1 U13696 ( .A(n10679), .B(n10678), .ZN(n10703) );
  NAND2_X1 U13697 ( .A1(n10705), .A2(n10703), .ZN(n12230) );
  XNOR2_X1 U13698 ( .A(n10681), .B(n10680), .ZN(n12187) );
  XNOR2_X1 U13699 ( .A(n12204), .B(n11976), .ZN(n12183) );
  OR2_X1 U13700 ( .A1(n12187), .A2(n12183), .ZN(n10682) );
  OR2_X1 U13701 ( .A1(n12230), .A2(n10682), .ZN(n10687) );
  NAND2_X1 U13702 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15764), .ZN(
        n10683) );
  NAND2_X1 U13703 ( .A1(n10684), .A2(n10683), .ZN(n10686) );
  NAND2_X1 U13704 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16280), .ZN(
        n10685) );
  NAND2_X1 U13705 ( .A1(n10687), .A2(n12197), .ZN(n12232) );
  AND2_X2 U13706 ( .A1(n13134), .A2(n19869), .ZN(n13178) );
  INV_X1 U13707 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19747) );
  INV_X1 U13708 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19743) );
  NOR2_X1 U13709 ( .A1(n19743), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n18877) );
  INV_X1 U13710 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19760) );
  NAND2_X1 U13711 ( .A1(n19743), .A2(n19760), .ZN(n19754) );
  NAND2_X1 U13712 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19867) );
  NAND2_X1 U13713 ( .A1(n19871), .A2(n19867), .ZN(n12200) );
  NOR2_X1 U13714 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n12200), .ZN(n10696) );
  NAND2_X1 U13715 ( .A1(n13178), .A2(n10696), .ZN(n19026) );
  INV_X1 U13716 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n10699) );
  INV_X1 U13717 ( .A(n10728), .ZN(n19228) );
  AND2_X2 U13718 ( .A1(n10721), .A2(n10700), .ZN(n10737) );
  NAND2_X1 U13719 ( .A1(n9863), .A2(n16273), .ZN(n16265) );
  NOR2_X1 U13720 ( .A1(n19385), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19734) );
  INV_X1 U13721 ( .A(n19734), .ZN(n10691) );
  NOR2_X1 U13722 ( .A1(n19741), .A2(n10691), .ZN(n16285) );
  NAND2_X1 U13723 ( .A1(n10692), .A2(n19385), .ZN(n19636) );
  AND2_X2 U13724 ( .A1(n19820), .A2(n19861), .ZN(n19206) );
  NOR3_X1 U13725 ( .A1(n16285), .A2(n18915), .A3(n19206), .ZN(n10693) );
  AND2_X2 U13726 ( .A1(n19863), .A2(n10693), .ZN(n19028) );
  INV_X1 U13727 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19868) );
  NAND2_X1 U13728 ( .A1(n19868), .A2(n19867), .ZN(n10717) );
  INV_X1 U13729 ( .A(n10717), .ZN(n10914) );
  NOR2_X1 U13730 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n10914), .ZN(n10694) );
  AND2_X1 U13731 ( .A1(n13134), .A2(n10694), .ZN(n10695) );
  OR2_X1 U13732 ( .A1(n13178), .A2(n10695), .ZN(n10697) );
  INV_X1 U13733 ( .A(n10696), .ZN(n16288) );
  AOI22_X1 U13734 ( .A1(P2_EBX_REG_30__SCAN_IN), .A2(n18957), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19028), .ZN(n10698) );
  OAI21_X1 U13735 ( .B1(n10699), .B2(n19041), .A(n10698), .ZN(n10720) );
  INV_X1 U13736 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13259) );
  INV_X1 U13737 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n19032) );
  NAND2_X1 U13738 ( .A1(n13259), .A2(n19032), .ZN(n10702) );
  MUX2_X1 U13739 ( .A(n10702), .B(n12310), .S(n12150), .Z(n11983) );
  MUX2_X1 U13740 ( .A(n11933), .B(n10703), .S(n12247), .Z(n12179) );
  INV_X1 U13741 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10704) );
  MUX2_X1 U13742 ( .A(n12179), .B(n10704), .S(n19237), .Z(n11971) );
  MUX2_X1 U13743 ( .A(n12306), .B(n10705), .S(n12247), .Z(n12178) );
  INV_X1 U13744 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n10706) );
  MUX2_X1 U13745 ( .A(n12178), .B(n10706), .S(n19237), .Z(n11991) );
  NAND2_X1 U13746 ( .A1(n11993), .A2(n11991), .ZN(n12020) );
  MUX2_X1 U13747 ( .A(P2_EBX_REG_5__SCAN_IN), .B(n12016), .S(n12150), .Z(
        n12019) );
  INV_X1 U13748 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n18998) );
  MUX2_X1 U13749 ( .A(n18998), .B(n12041), .S(n12150), .Z(n12049) );
  MUX2_X1 U13750 ( .A(P2_EBX_REG_7__SCAN_IN), .B(n12158), .S(n12150), .Z(
        n12055) );
  INV_X1 U13751 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n10707) );
  INV_X1 U13752 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n14812) );
  NAND2_X1 U13753 ( .A1(n12067), .A2(n14812), .ZN(n12070) );
  NAND2_X1 U13754 ( .A1(n19237), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10708) );
  INV_X1 U13755 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10850) );
  NOR2_X1 U13756 ( .A1(n12150), .A2(n10850), .ZN(n12083) );
  OAI21_X1 U13757 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(P2_EBX_REG_14__SCAN_IN), 
        .A(n19237), .ZN(n10709) );
  NOR2_X1 U13758 ( .A1(P2_EBX_REG_17__SCAN_IN), .A2(P2_EBX_REG_16__SCAN_IN), 
        .ZN(n10710) );
  NOR2_X1 U13759 ( .A1(n12150), .A2(n10710), .ZN(n10711) );
  NOR2_X1 U13760 ( .A1(P2_EBX_REG_18__SCAN_IN), .A2(P2_EBX_REG_19__SCAN_IN), 
        .ZN(n10712) );
  INV_X1 U13761 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n14944) );
  NAND2_X1 U13762 ( .A1(n19237), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n12132) );
  NAND2_X1 U13763 ( .A1(n12090), .A2(n12132), .ZN(n12138) );
  INV_X1 U13764 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10713) );
  NOR2_X1 U13765 ( .A1(n12150), .A2(n10713), .ZN(n12137) );
  INV_X1 U13766 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n14915) );
  NAND2_X1 U13767 ( .A1(n19237), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n12166) );
  NAND2_X1 U13768 ( .A1(n19237), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n12174) );
  INV_X1 U13769 ( .A(n12174), .ZN(n10715) );
  NAND2_X1 U13770 ( .A1(n19237), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12757) );
  NAND2_X1 U13771 ( .A1(n19237), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10716) );
  NOR2_X1 U13772 ( .A1(n19863), .A2(n12247), .ZN(n10915) );
  AND2_X1 U13773 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n10717), .ZN(n10718) );
  NAND2_X1 U13774 ( .A1(n10915), .A2(n10718), .ZN(n19014) );
  NOR2_X1 U13775 ( .A1(n12760), .A2(n19014), .ZN(n10719) );
  AOI211_X1 U13776 ( .C1(n15260), .C2(n19029), .A(n10720), .B(n10719), .ZN(
        n10919) );
  INV_X1 U13777 ( .A(n10727), .ZN(n10738) );
  NAND2_X1 U13778 ( .A1(n10908), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10768) );
  INV_X1 U13779 ( .A(n10733), .ZN(n12211) );
  NAND2_X1 U13780 ( .A1(n10737), .A2(n10734), .ZN(n12248) );
  NAND2_X1 U13781 ( .A1(n12248), .A2(n10140), .ZN(n10736) );
  NAND2_X1 U13782 ( .A1(n12290), .A2(n16269), .ZN(n10756) );
  INV_X1 U13783 ( .A(n10737), .ZN(n10748) );
  NAND3_X1 U13784 ( .A1(n10738), .A2(n10742), .A3(n10748), .ZN(n12220) );
  NAND2_X1 U13785 ( .A1(n12251), .A2(n10729), .ZN(n10744) );
  NAND3_X1 U13786 ( .A1(n10744), .A2(n10743), .A3(n16269), .ZN(n10747) );
  NAND2_X1 U13787 ( .A1(n10739), .A2(n19869), .ZN(n12257) );
  NAND2_X1 U13788 ( .A1(n10747), .A2(n10746), .ZN(n10755) );
  MUX2_X1 U13789 ( .A(n10721), .B(n12707), .S(n12215), .Z(n10751) );
  AND2_X1 U13790 ( .A1(n10748), .A2(n19223), .ZN(n10750) );
  NAND2_X1 U13791 ( .A1(n10739), .A2(n10729), .ZN(n10749) );
  NAND3_X1 U13792 ( .A1(n10751), .A2(n10750), .A3(n10749), .ZN(n10754) );
  INV_X1 U13793 ( .A(n10752), .ZN(n10753) );
  NAND3_X1 U13794 ( .A1(n10754), .A2(n10753), .A3(n10690), .ZN(n12255) );
  NAND3_X1 U13795 ( .A1(n10756), .A2(n10755), .A3(n12255), .ZN(n10757) );
  AND2_X2 U13796 ( .A1(n12703), .A2(n12194), .ZN(n12263) );
  NAND2_X1 U13797 ( .A1(n10787), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10765) );
  INV_X1 U13798 ( .A(n10760), .ZN(n10762) );
  AND3_X2 U13799 ( .A1(n19245), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n11932), 
        .ZN(n12644) );
  AND2_X2 U13800 ( .A1(n10762), .A2(n12644), .ZN(n12742) );
  NAND2_X1 U13801 ( .A1(n12742), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10764) );
  INV_X1 U13802 ( .A(n19861), .ZN(n10808) );
  NAND2_X1 U13803 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10763) );
  NAND2_X1 U13804 ( .A1(n10768), .A2(n10767), .ZN(n11901) );
  NAND2_X1 U13805 ( .A1(n10795), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10774) );
  INV_X1 U13806 ( .A(n10769), .ZN(n14100) );
  NAND2_X1 U13807 ( .A1(n12258), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10771) );
  NAND2_X1 U13808 ( .A1(n19861), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10770) );
  OAI211_X1 U13809 ( .C1(n14100), .C2(n10771), .A(n10856), .B(n10770), .ZN(
        n10772) );
  INV_X1 U13810 ( .A(n10772), .ZN(n10773) );
  NAND2_X1 U13811 ( .A1(n10774), .A2(n10773), .ZN(n11900) );
  NAND2_X1 U13812 ( .A1(n10795), .A2(n16229), .ZN(n10777) );
  AOI22_X1 U13813 ( .A1(n10775), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19861), 
        .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10776) );
  INV_X1 U13814 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n14868) );
  NAND2_X1 U13815 ( .A1(n10787), .A2(P2_EBX_REG_1__SCAN_IN), .ZN(n10779) );
  NAND2_X1 U13816 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n10778) );
  NAND2_X1 U13817 ( .A1(n10779), .A2(n10778), .ZN(n10780) );
  NAND2_X1 U13818 ( .A1(n10782), .A2(n10783), .ZN(n11903) );
  NAND2_X1 U13819 ( .A1(n11899), .A2(n11903), .ZN(n10786) );
  INV_X1 U13820 ( .A(n10782), .ZN(n10785) );
  NAND2_X1 U13821 ( .A1(n10786), .A2(n11904), .ZN(n11898) );
  INV_X1 U13822 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10793) );
  INV_X1 U13823 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n10790) );
  NAND2_X1 U13824 ( .A1(n10787), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10789) );
  NAND2_X1 U13825 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10788) );
  OAI211_X1 U13826 ( .C1(n10790), .C2(n10800), .A(n10789), .B(n10788), .ZN(
        n10791) );
  INV_X1 U13827 ( .A(n10791), .ZN(n10792) );
  OAI21_X1 U13828 ( .B1(n12371), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16287), 
        .ZN(n10794) );
  AOI21_X2 U13829 ( .B1(n10795), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n10794), .ZN(n10797) );
  XNOR2_X2 U13830 ( .A(n10796), .B(n10797), .ZN(n11897) );
  INV_X1 U13831 ( .A(n10796), .ZN(n10798) );
  NAND2_X1 U13832 ( .A1(n10798), .A2(n10797), .ZN(n10799) );
  INV_X1 U13833 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13972) );
  INV_X1 U13834 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n10803) );
  NAND2_X1 U13835 ( .A1(n10787), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10802) );
  NAND2_X1 U13836 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n10801) );
  OAI211_X1 U13837 ( .C1(n10803), .C2(n10800), .A(n10802), .B(n10801), .ZN(
        n10804) );
  INV_X1 U13838 ( .A(n10804), .ZN(n10805) );
  INV_X1 U13839 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n10814) );
  INV_X1 U13840 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19209) );
  OR2_X1 U13841 ( .A1(n9719), .A2(n19209), .ZN(n10813) );
  AOI22_X1 U13842 ( .A1(n12741), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10812) );
  OAI211_X1 U13843 ( .C1(n10913), .C2(n10814), .A(n10813), .B(n10812), .ZN(
        n13420) );
  INV_X1 U13844 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n13974) );
  INV_X1 U13845 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13970) );
  OR2_X1 U13846 ( .A1(n9719), .A2(n13970), .ZN(n10816) );
  AOI22_X1 U13847 ( .A1(n12741), .A2(P2_EBX_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10815) );
  OAI211_X1 U13848 ( .C1(n13974), .C2(n10913), .A(n10816), .B(n10815), .ZN(
        n13485) );
  INV_X1 U13849 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n20868) );
  OR2_X1 U13850 ( .A1(n9719), .A2(n20868), .ZN(n10821) );
  NAND2_X1 U13851 ( .A1(n12742), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n10819) );
  NAND2_X1 U13852 ( .A1(n12741), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n10818) );
  NAND2_X1 U13853 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10817) );
  AND3_X1 U13854 ( .A1(n10819), .A2(n10818), .A3(n10817), .ZN(n10820) );
  INV_X1 U13855 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15539) );
  OR2_X1 U13856 ( .A1(n9719), .A2(n15539), .ZN(n10827) );
  INV_X1 U13857 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n10824) );
  NAND2_X1 U13858 ( .A1(n12741), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n10823) );
  NAND2_X1 U13859 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10822) );
  OAI211_X1 U13860 ( .C1(n10824), .C2(n10913), .A(n10823), .B(n10822), .ZN(
        n10825) );
  INV_X1 U13861 ( .A(n10825), .ZN(n10826) );
  NAND2_X1 U13862 ( .A1(n10827), .A2(n10826), .ZN(n13491) );
  INV_X1 U13863 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n10830) );
  NAND2_X1 U13864 ( .A1(n12741), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10829) );
  NAND2_X1 U13865 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10828) );
  OAI211_X1 U13866 ( .C1(n10830), .C2(n10913), .A(n10829), .B(n10828), .ZN(
        n10831) );
  AOI21_X1 U13867 ( .B1(n9751), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n10831), .ZN(n13539) );
  INV_X1 U13868 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n10836) );
  NAND2_X1 U13869 ( .A1(n12741), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10835) );
  NAND2_X1 U13870 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n10834) );
  OAI211_X1 U13871 ( .C1(n10836), .C2(n10913), .A(n10835), .B(n10834), .ZN(
        n10837) );
  AOI21_X1 U13872 ( .B1(n9751), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n10837), .ZN(n13630) );
  INV_X1 U13873 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n10840) );
  INV_X1 U13874 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16207) );
  OR2_X1 U13875 ( .A1(n9719), .A2(n16207), .ZN(n10839) );
  AOI22_X1 U13876 ( .A1(n12741), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n10838) );
  OAI211_X1 U13877 ( .C1(n10913), .C2(n10840), .A(n10839), .B(n10838), .ZN(
        n13675) );
  NAND2_X1 U13878 ( .A1(n13628), .A2(n13675), .ZN(n13676) );
  INV_X1 U13879 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n10843) );
  NAND2_X1 U13880 ( .A1(n12741), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10842) );
  NAND2_X1 U13881 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10841) );
  OAI211_X1 U13882 ( .C1(n10843), .C2(n10913), .A(n10842), .B(n10841), .ZN(
        n10844) );
  AOI21_X1 U13883 ( .B1(n9751), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n10844), .ZN(n13122) );
  INV_X1 U13884 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n10848) );
  NAND2_X1 U13885 ( .A1(n12741), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10847) );
  NAND2_X1 U13886 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10846) );
  OAI211_X1 U13887 ( .C1(n10848), .C2(n10913), .A(n10847), .B(n10846), .ZN(
        n10849) );
  AOI21_X1 U13888 ( .B1(n9751), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n10849), .ZN(n13697) );
  INV_X1 U13889 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15488) );
  OR2_X1 U13890 ( .A1(n9719), .A2(n15488), .ZN(n10854) );
  NOR2_X1 U13891 ( .A1(n10913), .A2(n15187), .ZN(n10852) );
  OAI22_X1 U13892 ( .A1(n10856), .A2(n10850), .B1(n16287), .B2(n15188), .ZN(
        n10851) );
  NOR2_X1 U13893 ( .A1(n10852), .A2(n10851), .ZN(n10853) );
  NAND2_X1 U13894 ( .A1(n10854), .A2(n10853), .ZN(n13724) );
  INV_X1 U13895 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n20881) );
  OR2_X1 U13896 ( .A1(n9719), .A2(n20881), .ZN(n10860) );
  INV_X1 U13897 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n10855) );
  NOR2_X1 U13898 ( .A1(n10913), .A2(n10855), .ZN(n10858) );
  INV_X1 U13899 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n12106) );
  OAI22_X1 U13900 ( .A1(n10856), .A2(n12106), .B1(n16287), .B2(n9997), .ZN(
        n10857) );
  NOR2_X1 U13901 ( .A1(n10858), .A2(n10857), .ZN(n10859) );
  NAND2_X1 U13902 ( .A1(n10860), .A2(n10859), .ZN(n13793) );
  INV_X1 U13903 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n10863) );
  NAND2_X1 U13904 ( .A1(n12741), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10862) );
  NAND2_X1 U13905 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10861) );
  OAI211_X1 U13906 ( .C1(n10863), .C2(n10913), .A(n10862), .B(n10861), .ZN(
        n10864) );
  AOI21_X1 U13907 ( .B1(n9751), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n10864), .ZN(n13105) );
  INV_X1 U13908 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n19775) );
  NAND2_X1 U13909 ( .A1(n12741), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10868) );
  NAND2_X1 U13910 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10867) );
  OAI211_X1 U13911 ( .C1(n19775), .C2(n10913), .A(n10868), .B(n10867), .ZN(
        n10869) );
  AOI21_X1 U13912 ( .B1(n9751), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n10869), .ZN(n13939) );
  INV_X1 U13913 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19777) );
  INV_X1 U13914 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21010) );
  OR2_X1 U13915 ( .A1(n9719), .A2(n21010), .ZN(n10871) );
  AOI22_X1 U13916 ( .A1(n12741), .A2(P2_EBX_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n10870) );
  OAI211_X1 U13917 ( .C1(n10913), .C2(n19777), .A(n10871), .B(n10870), .ZN(
        n14962) );
  INV_X1 U13918 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n10874) );
  INV_X1 U13919 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15410) );
  OR2_X1 U13920 ( .A1(n9719), .A2(n15410), .ZN(n10873) );
  AOI22_X1 U13921 ( .A1(n12741), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n10872) );
  OAI211_X1 U13922 ( .C1(n10913), .C2(n10874), .A(n10873), .B(n10872), .ZN(
        n14794) );
  INV_X1 U13923 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n10877) );
  NAND2_X1 U13924 ( .A1(n12741), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n10876) );
  NAND2_X1 U13925 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10875) );
  OAI211_X1 U13926 ( .C1(n10877), .C2(n10913), .A(n10876), .B(n10875), .ZN(
        n10878) );
  AOI21_X1 U13927 ( .B1(n9751), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n10878), .ZN(n14954) );
  INV_X1 U13928 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n10882) );
  NAND2_X1 U13929 ( .A1(n12741), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10881) );
  NAND2_X1 U13930 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10880) );
  OAI211_X1 U13931 ( .C1(n10882), .C2(n10913), .A(n10881), .B(n10880), .ZN(
        n10883) );
  AOI21_X1 U13932 ( .B1(n9751), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n10883), .ZN(n14777) );
  INV_X1 U13933 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n10886) );
  NAND2_X1 U13934 ( .A1(n12741), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10885) );
  NAND2_X1 U13935 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10884) );
  OAI211_X1 U13936 ( .C1(n10886), .C2(n10913), .A(n10885), .B(n10884), .ZN(
        n10887) );
  AOI21_X1 U13937 ( .B1(n9751), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n10887), .ZN(n14759) );
  INV_X1 U13938 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19783) );
  INV_X1 U13939 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15338) );
  OR2_X1 U13940 ( .A1(n9719), .A2(n15338), .ZN(n10889) );
  AOI22_X1 U13941 ( .A1(n12741), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n10888) );
  OAI211_X1 U13942 ( .C1(n10913), .C2(n19783), .A(n10889), .B(n10888), .ZN(
        n14744) );
  INV_X1 U13943 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n15102) );
  NAND2_X1 U13944 ( .A1(n12741), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10891) );
  NAND2_X1 U13945 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10890) );
  OAI211_X1 U13946 ( .C1(n15102), .C2(n10913), .A(n10891), .B(n10890), .ZN(
        n10892) );
  AOI21_X1 U13947 ( .B1(n9751), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n10892), .ZN(n14729) );
  INV_X1 U13948 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19786) );
  NAND2_X1 U13949 ( .A1(n12741), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10894) );
  NAND2_X1 U13950 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10893) );
  OAI211_X1 U13951 ( .C1(n19786), .C2(n10913), .A(n10894), .B(n10893), .ZN(
        n10895) );
  AOI21_X1 U13952 ( .B1(n9751), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n10895), .ZN(n14922) );
  INV_X1 U13953 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19788) );
  INV_X1 U13954 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15316) );
  OR2_X1 U13955 ( .A1(n9719), .A2(n15316), .ZN(n10897) );
  AOI22_X1 U13956 ( .A1(n12741), .A2(P2_EBX_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n10896) );
  OAI211_X1 U13957 ( .C1(n10913), .C2(n19788), .A(n10897), .B(n10896), .ZN(
        n14913) );
  INV_X1 U13958 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n10900) );
  INV_X1 U13959 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15307) );
  OR2_X1 U13960 ( .A1(n9719), .A2(n15307), .ZN(n10899) );
  AOI22_X1 U13961 ( .A1(n12741), .A2(P2_EBX_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n10898) );
  OAI211_X1 U13962 ( .C1(n10913), .C2(n10900), .A(n10899), .B(n10898), .ZN(
        n14908) );
  NAND2_X1 U13963 ( .A1(n14907), .A2(n14908), .ZN(n14897) );
  INV_X1 U13964 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19792) );
  NAND2_X1 U13965 ( .A1(n12741), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10902) );
  NAND2_X1 U13966 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10901) );
  OAI211_X1 U13967 ( .C1(n19792), .C2(n10913), .A(n10902), .B(n10901), .ZN(
        n10903) );
  AOI21_X1 U13968 ( .B1(n9751), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n10903), .ZN(n14898) );
  INV_X1 U13969 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19793) );
  NAND2_X1 U13970 ( .A1(n12741), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n10906) );
  NAND2_X1 U13971 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10905) );
  OAI211_X1 U13972 ( .C1(n19793), .C2(n10913), .A(n10906), .B(n10905), .ZN(
        n10907) );
  AOI21_X1 U13973 ( .B1(n9751), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n10907), .ZN(n12299) );
  INV_X1 U13974 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19795) );
  INV_X1 U13975 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15277) );
  OR2_X1 U13976 ( .A1(n9719), .A2(n15277), .ZN(n10910) );
  AOI22_X1 U13977 ( .A1(n12741), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n10909) );
  OAI211_X1 U13978 ( .C1(n10913), .C2(n19795), .A(n10910), .B(n10909), .ZN(
        n14882) );
  INV_X1 U13979 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n19798) );
  INV_X1 U13980 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15261) );
  OR2_X1 U13981 ( .A1(n9719), .A2(n15261), .ZN(n10912) );
  AOI22_X1 U13982 ( .A1(n12741), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n10911) );
  OAI211_X1 U13983 ( .C1(n10913), .C2(n19798), .A(n10912), .B(n10911), .ZN(
        n12740) );
  INV_X1 U13984 ( .A(n15270), .ZN(n10917) );
  NAND2_X1 U13985 ( .A1(n10915), .A2(n10914), .ZN(n19037) );
  NAND3_X1 U13986 ( .A1(n10920), .A2(n10919), .A3(n10918), .ZN(P2_U2825) );
  AND2_X2 U13987 ( .A1(n14149), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10927) );
  AOI22_X1 U13988 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11149), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n10925) );
  AOI22_X1 U13989 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n14118), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10924) );
  AND2_X2 U13990 ( .A1(n10926), .A2(n13459), .ZN(n11237) );
  AOI22_X1 U13991 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10923) );
  AOI22_X1 U13992 ( .A1(n14112), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10922) );
  NAND4_X1 U13993 ( .A1(n10925), .A2(n10924), .A3(n10923), .A4(n10922), .ZN(
        n10936) );
  AND2_X2 U13994 ( .A1(n13460), .A2(n10928), .ZN(n11597) );
  AOI22_X1 U13995 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10934) );
  AOI22_X1 U13996 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11070), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n10933) );
  AND2_X2 U13997 ( .A1(n13468), .A2(n10930), .ZN(n11297) );
  AOI22_X1 U13998 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11297), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10932) );
  AND2_X2 U13999 ( .A1(n10930), .A2(n10929), .ZN(n11254) );
  AOI22_X1 U14000 ( .A1(n11616), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10931) );
  NAND4_X1 U14001 ( .A1(n10934), .A2(n10933), .A3(n10932), .A4(n10931), .ZN(
        n10935) );
  NOR2_X1 U14002 ( .A1(n10936), .A2(n10935), .ZN(n11699) );
  AOI22_X1 U14003 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n14112), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10940) );
  AOI22_X1 U14004 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10939) );
  AOI22_X1 U14005 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10938) );
  AOI22_X1 U14006 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10937) );
  NAND4_X1 U14007 ( .A1(n10940), .A2(n10939), .A3(n10938), .A4(n10937), .ZN(
        n10946) );
  AOI22_X1 U14008 ( .A1(n14118), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11149), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n10944) );
  AOI22_X1 U14009 ( .A1(n11262), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10943) );
  AOI22_X1 U14010 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9725), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n10942) );
  AOI22_X1 U14011 ( .A1(n9721), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10941) );
  NAND4_X1 U14012 ( .A1(n10944), .A2(n10943), .A3(n10942), .A4(n10941), .ZN(
        n10945) );
  NOR2_X1 U14013 ( .A1(n10946), .A2(n10945), .ZN(n11677) );
  AOI22_X1 U14014 ( .A1(n10968), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11149), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n10950) );
  AOI22_X1 U14015 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10949) );
  AOI22_X1 U14016 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9725), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10948) );
  AOI22_X1 U14017 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11254), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10947) );
  NAND4_X1 U14018 ( .A1(n10950), .A2(n10949), .A3(n10948), .A4(n10947), .ZN(
        n10956) );
  AOI22_X1 U14019 ( .A1(n11262), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11597), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10954) );
  AOI22_X1 U14020 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10953) );
  AOI22_X1 U14021 ( .A1(n14112), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10952) );
  AOI22_X1 U14022 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10951) );
  NAND4_X1 U14023 ( .A1(n10954), .A2(n10953), .A3(n10952), .A4(n10951), .ZN(
        n10955) );
  NOR2_X1 U14024 ( .A1(n10956), .A2(n10955), .ZN(n11661) );
  AOI22_X1 U14025 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10961) );
  AOI22_X1 U14026 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10960) );
  AOI22_X1 U14027 ( .A1(n11262), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9725), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U14028 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10958) );
  NAND4_X1 U14029 ( .A1(n10961), .A2(n10960), .A3(n10959), .A4(n10958), .ZN(
        n10967) );
  AOI22_X1 U14030 ( .A1(n10968), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11149), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10965) );
  AOI22_X1 U14031 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10964) );
  AOI22_X1 U14032 ( .A1(n14112), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10963) );
  AOI22_X1 U14033 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10962) );
  NAND4_X1 U14034 ( .A1(n10965), .A2(n10964), .A3(n10963), .A4(n10962), .ZN(
        n10966) );
  NOR2_X1 U14035 ( .A1(n10967), .A2(n10966), .ZN(n11660) );
  OR2_X1 U14036 ( .A1(n11661), .A2(n11660), .ZN(n11672) );
  AOI22_X1 U14037 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n14112), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10972) );
  AOI22_X1 U14038 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n14118), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10971) );
  AOI22_X1 U14039 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10970) );
  AOI22_X1 U14040 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10969) );
  NAND4_X1 U14041 ( .A1(n10972), .A2(n10971), .A3(n10970), .A4(n10969), .ZN(
        n10978) );
  AOI22_X1 U14042 ( .A1(n11262), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10976) );
  INV_X1 U14043 ( .A(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n20992) );
  AOI22_X1 U14044 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10975) );
  AOI22_X1 U14045 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11149), .B1(
        n9725), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10974) );
  AOI22_X1 U14046 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11254), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10973) );
  NAND4_X1 U14047 ( .A1(n10976), .A2(n10975), .A3(n10974), .A4(n10973), .ZN(
        n10977) );
  NOR2_X1 U14048 ( .A1(n10978), .A2(n10977), .ZN(n11671) );
  NOR2_X1 U14049 ( .A1(n11677), .A2(n11678), .ZN(n11691) );
  AOI22_X1 U14050 ( .A1(n11262), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10982) );
  AOI22_X1 U14051 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10981) );
  AOI22_X1 U14052 ( .A1(n14112), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10980) );
  AOI22_X1 U14053 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10979) );
  NAND4_X1 U14054 ( .A1(n10982), .A2(n10981), .A3(n10980), .A4(n10979), .ZN(
        n10988) );
  AOI22_X1 U14055 ( .A1(n14118), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11149), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10986) );
  AOI22_X1 U14056 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10985) );
  AOI22_X1 U14057 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9725), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10984) );
  AOI22_X1 U14058 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10983) );
  NAND4_X1 U14059 ( .A1(n10986), .A2(n10985), .A3(n10984), .A4(n10983), .ZN(
        n10987) );
  OR2_X1 U14060 ( .A1(n10988), .A2(n10987), .ZN(n11689) );
  NAND2_X1 U14061 ( .A1(n11691), .A2(n11689), .ZN(n11700) );
  NOR2_X1 U14062 ( .A1(n11699), .A2(n11700), .ZN(n11711) );
  AOI22_X1 U14063 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10992) );
  INV_X1 U14064 ( .A(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n20942) );
  AOI22_X1 U14065 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10991) );
  AOI22_X1 U14066 ( .A1(n14112), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10990) );
  AOI22_X1 U14067 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11297), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10989) );
  NAND4_X1 U14068 ( .A1(n10992), .A2(n10991), .A3(n10990), .A4(n10989), .ZN(
        n10998) );
  AOI22_X1 U14069 ( .A1(n10968), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11149), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10996) );
  AOI22_X1 U14070 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10995) );
  AOI22_X1 U14071 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9749), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10994) );
  AOI22_X1 U14072 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10993) );
  NAND4_X1 U14073 ( .A1(n10996), .A2(n10995), .A3(n10994), .A4(n10993), .ZN(
        n10997) );
  OR2_X1 U14074 ( .A1(n10998), .A2(n10997), .ZN(n11709) );
  NAND2_X1 U14075 ( .A1(n11711), .A2(n11709), .ZN(n14126) );
  AOI22_X1 U14076 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11002) );
  AOI22_X1 U14077 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11262), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11001) );
  AOI22_X1 U14078 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11000) );
  AOI22_X1 U14079 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10999) );
  NAND4_X1 U14080 ( .A1(n11002), .A2(n11001), .A3(n11000), .A4(n10999), .ZN(
        n11008) );
  AOI22_X1 U14081 ( .A1(n14118), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11149), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11006) );
  AOI22_X1 U14082 ( .A1(n9721), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11070), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11005) );
  AOI22_X1 U14083 ( .A1(n14112), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11297), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11004) );
  AOI22_X1 U14084 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11003) );
  NAND4_X1 U14085 ( .A1(n11006), .A2(n11005), .A3(n11004), .A4(n11003), .ZN(
        n11007) );
  NOR2_X1 U14086 ( .A1(n11008), .A2(n11007), .ZN(n14127) );
  XOR2_X1 U14087 ( .A(n14126), .B(n14127), .Z(n11081) );
  NAND2_X1 U14088 ( .A1(n11095), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11012) );
  NAND2_X1 U14089 ( .A1(n10968), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11011) );
  NAND2_X1 U14090 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11010) );
  NAND2_X1 U14091 ( .A1(n11254), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11009) );
  AND4_X2 U14092 ( .A1(n11012), .A2(n11011), .A3(n11010), .A4(n11009), .ZN(
        n11028) );
  NAND2_X1 U14093 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11016) );
  NAND2_X1 U14094 ( .A1(n11597), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11015) );
  NAND2_X1 U14095 ( .A1(n11237), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11014) );
  NAND2_X1 U14096 ( .A1(n11090), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11013) );
  NAND2_X1 U14097 ( .A1(n11260), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11020) );
  NAND2_X1 U14098 ( .A1(n9760), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11019) );
  NAND2_X1 U14099 ( .A1(n9741), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11018) );
  NAND2_X1 U14100 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11017) );
  NAND2_X1 U14101 ( .A1(n11253), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11024) );
  NAND2_X1 U14102 ( .A1(n11252), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11023) );
  NAND2_X1 U14103 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11022) );
  NAND2_X1 U14104 ( .A1(n9750), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11021) );
  NAND4_X4 U14105 ( .A1(n11028), .A2(n11027), .A3(n11026), .A4(n11025), .ZN(
        n11167) );
  NAND2_X1 U14106 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n11032) );
  NAND2_X1 U14107 ( .A1(n11260), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11031) );
  NAND2_X1 U14108 ( .A1(n11597), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n11030) );
  NAND2_X1 U14109 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11029) );
  NAND2_X1 U14110 ( .A1(n11237), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11036) );
  NAND2_X1 U14111 ( .A1(n11090), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11035) );
  NAND2_X1 U14112 ( .A1(n9760), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11034) );
  NAND2_X1 U14113 ( .A1(n9742), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11033) );
  NAND2_X1 U14114 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n11040) );
  NAND2_X1 U14115 ( .A1(n11095), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n11039) );
  NAND2_X1 U14116 ( .A1(n11252), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n11038) );
  NAND2_X1 U14117 ( .A1(n9749), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11037) );
  NAND2_X1 U14118 ( .A1(n10968), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11045) );
  NAND2_X1 U14119 ( .A1(n11253), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n11044) );
  NAND2_X1 U14120 ( .A1(n11254), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11043) );
  NAND2_X1 U14121 ( .A1(n11107), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11042) );
  NAND2_X1 U14122 ( .A1(n11260), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11053) );
  NAND2_X1 U14123 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11052) );
  NAND2_X1 U14124 ( .A1(n9741), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11051) );
  NAND2_X1 U14125 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11050) );
  NAND2_X1 U14126 ( .A1(n10968), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11057) );
  NAND2_X1 U14127 ( .A1(n9755), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11056) );
  NAND2_X1 U14128 ( .A1(n11254), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11055) );
  NAND2_X1 U14129 ( .A1(n9759), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11054) );
  NAND2_X1 U14130 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11061) );
  NAND2_X1 U14131 ( .A1(n11597), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11060) );
  NAND2_X1 U14132 ( .A1(n11237), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11059) );
  NAND2_X1 U14133 ( .A1(n11090), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11058) );
  NAND2_X1 U14134 ( .A1(n11253), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11065) );
  NAND2_X1 U14135 ( .A1(n11252), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11064) );
  NAND2_X1 U14136 ( .A1(n11107), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11063) );
  NAND2_X1 U14137 ( .A1(n9750), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11062) );
  INV_X2 U14138 ( .A(n11165), .ZN(n11180) );
  AOI22_X1 U14139 ( .A1(n11237), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11090), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11074) );
  AOI22_X1 U14140 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11073) );
  AOI22_X1 U14141 ( .A1(n11597), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9749), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11072) );
  AOI22_X1 U14142 ( .A1(n10968), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11254), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11071) );
  AOI22_X1 U14143 ( .A1(n11260), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11297), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11078) );
  AOI22_X1 U14144 ( .A1(n11095), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9752), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11077) );
  AOI22_X1 U14145 ( .A1(n11253), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9748), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11076) );
  AOI22_X1 U14146 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11252), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11075) );
  INV_X1 U14147 ( .A(n11168), .ZN(n11080) );
  INV_X1 U14148 ( .A(n13196), .ZN(n14716) );
  NAND2_X1 U14149 ( .A1(n11081), .A2(n11714), .ZN(n11084) );
  NAND2_X1 U14150 ( .A1(n14137), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n11083) );
  INV_X1 U14151 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20579) );
  OAI21_X1 U14152 ( .B1(n20906), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n20579), .ZN(n11082) );
  NAND3_X1 U14153 ( .A1(n11084), .A2(n11083), .A3(n11082), .ZN(n11089) );
  INV_X1 U14154 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n20853) );
  INV_X1 U14155 ( .A(n11368), .ZN(n11085) );
  INV_X1 U14156 ( .A(n11685), .ZN(n11086) );
  NAND2_X1 U14157 ( .A1(n11086), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11695) );
  INV_X1 U14158 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14275) );
  INV_X1 U14159 ( .A(n11705), .ZN(n11087) );
  NAND2_X1 U14160 ( .A1(n11087), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n11717) );
  INV_X1 U14161 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11716) );
  XNOR2_X1 U14162 ( .A(n13739), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14437) );
  NOR2_X2 U14163 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n14135) );
  NAND2_X1 U14164 ( .A1(n14437), .A2(n14135), .ZN(n11088) );
  NAND2_X1 U14165 ( .A1(n11089), .A2(n11088), .ZN(n11723) );
  AOI22_X1 U14166 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11597), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11094) );
  AOI22_X1 U14167 ( .A1(n11237), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11090), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11093) );
  AOI22_X1 U14168 ( .A1(n11260), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9741), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11092) );
  AOI22_X1 U14169 ( .A1(n9760), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11297), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11091) );
  NAND4_X1 U14170 ( .A1(n11094), .A2(n11093), .A3(n11092), .A4(n11091), .ZN(
        n11101) );
  AOI22_X1 U14171 ( .A1(n11253), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9748), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11098) );
  AOI22_X1 U14172 ( .A1(n11252), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11070), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11097) );
  AOI22_X1 U14173 ( .A1(n11095), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11254), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11096) );
  NAND4_X1 U14174 ( .A1(n11099), .A2(n11098), .A3(n11097), .A4(n11096), .ZN(
        n11100) );
  AOI22_X1 U14175 ( .A1(n11253), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n10968), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11106) );
  AOI22_X1 U14176 ( .A1(n11090), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11597), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11105) );
  AOI22_X1 U14177 ( .A1(n11237), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11104) );
  AOI22_X1 U14178 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11254), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11103) );
  NAND4_X1 U14179 ( .A1(n11106), .A2(n11105), .A3(n11104), .A4(n11103), .ZN(
        n11113) );
  AOI22_X1 U14180 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11260), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11111) );
  AOI22_X1 U14181 ( .A1(n9754), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11107), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11110) );
  AOI22_X1 U14182 ( .A1(n11136), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11297), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11108) );
  NAND4_X1 U14183 ( .A1(n11111), .A2(n11110), .A3(n11109), .A4(n11108), .ZN(
        n11112) );
  NAND2_X1 U14184 ( .A1(n11095), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11118) );
  NAND2_X1 U14185 ( .A1(n10968), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11117) );
  NAND2_X1 U14186 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11116) );
  NAND2_X1 U14187 ( .A1(n11254), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11115) );
  NAND2_X1 U14188 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11122) );
  NAND2_X1 U14189 ( .A1(n11597), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11121) );
  NAND2_X1 U14190 ( .A1(n11237), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11120) );
  NAND2_X1 U14191 ( .A1(n11090), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11119) );
  NAND2_X1 U14192 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11125) );
  NAND2_X1 U14193 ( .A1(n11260), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11124) );
  NAND2_X1 U14194 ( .A1(n9741), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11123) );
  NAND2_X1 U14195 ( .A1(n11125), .A2(n10153), .ZN(n11126) );
  NAND2_X1 U14196 ( .A1(n11253), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11130) );
  NAND2_X1 U14197 ( .A1(n11252), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11129) );
  NAND2_X1 U14198 ( .A1(n9748), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11128) );
  NAND2_X1 U14199 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11127) );
  NAND4_X4 U14200 ( .A1(n11134), .A2(n11133), .A3(n11132), .A4(n11131), .ZN(
        n13748) );
  NOR2_X1 U14201 ( .A1(n11733), .A2(n13748), .ZN(n11135) );
  NAND2_X1 U14202 ( .A1(n11237), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11140) );
  NAND2_X1 U14203 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11139) );
  NAND2_X1 U14204 ( .A1(n9760), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11138) );
  NAND2_X1 U14205 ( .A1(n11297), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11137) );
  NAND2_X1 U14206 ( .A1(n11090), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11144) );
  NAND2_X1 U14207 ( .A1(n11597), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11143) );
  NAND2_X1 U14208 ( .A1(n11260), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11142) );
  NAND2_X1 U14209 ( .A1(n9741), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11141) );
  NAND2_X1 U14210 ( .A1(n9754), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11148) );
  NAND2_X1 U14211 ( .A1(n11252), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11147) );
  NAND2_X1 U14212 ( .A1(n11253), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11146) );
  NAND2_X1 U14213 ( .A1(n11254), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11145) );
  NAND2_X1 U14214 ( .A1(n10968), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11153) );
  NAND2_X1 U14215 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11152) );
  NAND2_X1 U14216 ( .A1(n11070), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11151) );
  NAND2_X1 U14217 ( .A1(n9747), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11150) );
  NAND2_X1 U14218 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20648) );
  OAI21_X1 U14219 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(P1_STATE_REG_2__SCAN_IN), 
        .A(n20648), .ZN(n13195) );
  NAND2_X1 U14220 ( .A1(n9722), .A2(n13195), .ZN(n11160) );
  NAND3_X1 U14221 ( .A1(n11183), .A2(n20139), .A3(n13470), .ZN(n13426) );
  AOI21_X1 U14222 ( .B1(n13153), .B2(n11160), .A(n13405), .ZN(n11161) );
  INV_X1 U14223 ( .A(n13470), .ZN(n13391) );
  NAND2_X1 U14224 ( .A1(n13391), .A2(n13746), .ZN(n11164) );
  NAND2_X1 U14225 ( .A1(n13386), .A2(n11787), .ZN(n11163) );
  NAND2_X1 U14226 ( .A1(n13445), .A2(n13748), .ZN(n11162) );
  NAND2_X1 U14227 ( .A1(n20139), .A2(n11782), .ZN(n11166) );
  NAND2_X1 U14228 ( .A1(n11166), .A2(n13568), .ZN(n13197) );
  NOR2_X2 U14229 ( .A1(n13197), .A2(n11167), .ZN(n11186) );
  NAND2_X1 U14230 ( .A1(n11186), .A2(n11168), .ZN(n11179) );
  NAND2_X1 U14231 ( .A1(n11168), .A2(n13748), .ZN(n11169) );
  NAND2_X1 U14232 ( .A1(n11169), .A2(n20721), .ZN(n11170) );
  NAND2_X1 U14233 ( .A1(n11179), .A2(n11170), .ZN(n13394) );
  NAND2_X1 U14234 ( .A1(n11179), .A2(n13196), .ZN(n11172) );
  NAND2_X1 U14235 ( .A1(n19883), .A2(n20639), .ZN(n13500) );
  NAND2_X1 U14236 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11200) );
  OAI21_X1 U14237 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n11200), .ZN(n20411) );
  OR2_X1 U14238 ( .A1(n15727), .A2(n20414), .ZN(n11194) );
  OAI21_X1 U14239 ( .B1(n13500), .B2(n20411), .A(n11194), .ZN(n11174) );
  INV_X1 U14240 ( .A(n11174), .ZN(n11175) );
  AND2_X2 U14241 ( .A1(n11176), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11195) );
  XNOR2_X2 U14242 ( .A(n11177), .B(n11195), .ZN(n20212) );
  INV_X2 U14243 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14149) );
  MUX2_X1 U14244 ( .A(n13500), .B(n15727), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n11178) );
  NAND3_X1 U14245 ( .A1(n11179), .A2(n13751), .A3(n13196), .ZN(n11191) );
  NAND2_X1 U14246 ( .A1(n13470), .A2(n11180), .ZN(n13399) );
  NAND4_X1 U14247 ( .A1(n13399), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n19883), 
        .A4(n13746), .ZN(n11181) );
  NOR2_X1 U14248 ( .A1(n11181), .A2(n13398), .ZN(n11190) );
  INV_X1 U14249 ( .A(n11182), .ZN(n13385) );
  INV_X1 U14250 ( .A(n11184), .ZN(n13562) );
  NAND3_X1 U14251 ( .A1(n11168), .A2(n13562), .A3(n13360), .ZN(n11185) );
  NAND2_X1 U14252 ( .A1(n13385), .A2(n11185), .ZN(n11189) );
  INV_X1 U14253 ( .A(n11186), .ZN(n11187) );
  NAND2_X1 U14254 ( .A1(n11187), .A2(n13955), .ZN(n11188) );
  INV_X1 U14255 ( .A(n11275), .ZN(n11192) );
  INV_X1 U14256 ( .A(n11194), .ZN(n11196) );
  OR2_X1 U14257 ( .A1(n11198), .A2(n10921), .ZN(n11205) );
  INV_X1 U14258 ( .A(n13500), .ZN(n11203) );
  INV_X1 U14259 ( .A(n11200), .ZN(n11199) );
  NAND2_X1 U14260 ( .A1(n11199), .A2(n20487), .ZN(n20455) );
  NAND2_X1 U14261 ( .A1(n11200), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11201) );
  NAND2_X1 U14262 ( .A1(n20455), .A2(n11201), .ZN(n20109) );
  INV_X1 U14263 ( .A(n15727), .ZN(n11202) );
  AOI22_X1 U14264 ( .A1(n11203), .A2(n20109), .B1(n11202), .B2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n11204) );
  INV_X1 U14265 ( .A(n11206), .ZN(n11207) );
  AOI22_X1 U14266 ( .A1(n11253), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n14118), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11212) );
  AOI22_X1 U14267 ( .A1(n11262), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11211) );
  AOI22_X1 U14268 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11210) );
  AOI22_X1 U14269 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11209) );
  NAND4_X1 U14270 ( .A1(n11212), .A2(n11211), .A3(n11210), .A4(n11209), .ZN(
        n11218) );
  AOI22_X1 U14271 ( .A1(n11260), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11216) );
  AOI22_X1 U14272 ( .A1(n9759), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11215) );
  AOI22_X1 U14273 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9725), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11214) );
  AOI22_X1 U14274 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11297), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11213) );
  NAND4_X1 U14275 ( .A1(n11216), .A2(n11215), .A3(n11214), .A4(n11213), .ZN(
        n11217) );
  AOI22_X1 U14276 ( .A1(n11775), .A2(n13522), .B1(n11770), .B2(
        P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11219) );
  AOI22_X1 U14277 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11253), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11226) );
  AOI22_X1 U14278 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11225) );
  AOI22_X1 U14279 ( .A1(n9754), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11224) );
  AOI22_X1 U14280 ( .A1(n10968), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11223) );
  NAND4_X1 U14281 ( .A1(n11226), .A2(n11225), .A3(n11224), .A4(n11223), .ZN(
        n11232) );
  AOI22_X1 U14282 ( .A1(n11237), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11230) );
  AOI22_X1 U14283 ( .A1(n11260), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11229) );
  AOI22_X1 U14284 ( .A1(n9759), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9725), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11228) );
  AOI22_X1 U14285 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11297), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11227) );
  NAND4_X1 U14286 ( .A1(n11230), .A2(n11229), .A3(n11228), .A4(n11227), .ZN(
        n11231) );
  NAND2_X1 U14287 ( .A1(n11222), .A2(n13954), .ZN(n13950) );
  AOI22_X1 U14288 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10968), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11236) );
  AOI22_X1 U14289 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11235) );
  AOI22_X1 U14290 ( .A1(n9755), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11234) );
  AOI22_X1 U14291 ( .A1(n11260), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11233) );
  NAND4_X1 U14292 ( .A1(n11236), .A2(n11235), .A3(n11234), .A4(n11233), .ZN(
        n11243) );
  AOI22_X1 U14293 ( .A1(n11237), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11241) );
  AOI22_X1 U14294 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11240) );
  AOI22_X1 U14295 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11239) );
  AOI22_X1 U14296 ( .A1(n11253), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9725), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11238) );
  NAND4_X1 U14297 ( .A1(n11241), .A2(n11240), .A3(n11239), .A4(n11238), .ZN(
        n11242) );
  INV_X1 U14298 ( .A(n11270), .ZN(n11277) );
  INV_X1 U14299 ( .A(n13954), .ZN(n11244) );
  NAND3_X1 U14300 ( .A1(n11277), .A2(n11244), .A3(n13520), .ZN(n11245) );
  INV_X1 U14301 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20883) );
  AOI21_X1 U14302 ( .B1(n11249), .B2(n13520), .A(n20639), .ZN(n11250) );
  OAI211_X1 U14303 ( .C1(n11764), .C2(n20883), .A(n11250), .B(n13950), .ZN(
        n11349) );
  INV_X1 U14304 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11272) );
  INV_X1 U14305 ( .A(n11251), .ZN(n11269) );
  AOI22_X1 U14306 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11253), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11259) );
  AOI22_X1 U14307 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n11597), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11258) );
  AOI22_X1 U14308 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11257) );
  BUF_X1 U14309 ( .A(n11254), .Z(n11255) );
  AOI22_X1 U14310 ( .A1(n9752), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11256) );
  NAND4_X1 U14311 ( .A1(n11259), .A2(n11258), .A3(n11257), .A4(n11256), .ZN(
        n11268) );
  AOI22_X1 U14313 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11260), .B1(
        n11261), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11266) );
  AOI22_X1 U14314 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n11095), .B1(
        n14118), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11265) );
  AOI22_X1 U14315 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n11616), .B1(
        n9725), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11264) );
  AOI22_X1 U14316 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11297), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11263) );
  NAND4_X1 U14317 ( .A1(n11266), .A2(n11265), .A3(n11264), .A4(n11263), .ZN(
        n11267) );
  NAND2_X1 U14318 ( .A1(n11269), .A2(n13521), .ZN(n11271) );
  OAI211_X1 U14319 ( .C1(n11272), .C2(n11764), .A(n11271), .B(n11270), .ZN(
        n11273) );
  INV_X1 U14320 ( .A(n11273), .ZN(n11274) );
  NAND2_X1 U14321 ( .A1(n11277), .A2(n13521), .ZN(n11278) );
  OR2_X1 U14322 ( .A1(n11198), .A2(n11280), .ZN(n11284) );
  NAND3_X1 U14323 ( .A1(n20486), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20323) );
  NOR3_X1 U14324 ( .A1(n20486), .A2(n20487), .A3(n20414), .ZN(n20589) );
  INV_X1 U14325 ( .A(n20589), .ZN(n20580) );
  INV_X1 U14326 ( .A(n20630), .ZN(n11281) );
  OAI21_X1 U14327 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20343), .A(
        n11281), .ZN(n20101) );
  OAI22_X1 U14328 ( .A1(n13500), .A2(n20101), .B1(n15727), .B2(n20486), .ZN(
        n11282) );
  INV_X1 U14329 ( .A(n11282), .ZN(n11283) );
  NAND2_X1 U14330 ( .A1(n20349), .A2(n20639), .ZN(n11296) );
  AOI22_X1 U14331 ( .A1(n11262), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11288) );
  AOI22_X1 U14332 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11287) );
  AOI22_X1 U14333 ( .A1(n11260), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11286) );
  AOI22_X1 U14334 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11297), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11285) );
  NAND4_X1 U14335 ( .A1(n11288), .A2(n11287), .A3(n11286), .A4(n11285), .ZN(
        n11294) );
  AOI22_X1 U14336 ( .A1(n10968), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9752), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11292) );
  AOI22_X1 U14337 ( .A1(n11253), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11291) );
  AOI22_X1 U14338 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9725), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11290) );
  AOI22_X1 U14339 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11289) );
  NAND4_X1 U14340 ( .A1(n11292), .A2(n11291), .A3(n11290), .A4(n11289), .ZN(
        n11293) );
  AOI22_X1 U14341 ( .A1(n11775), .A2(n13645), .B1(n11770), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11295) );
  AOI22_X1 U14342 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n10968), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11301) );
  AOI22_X1 U14343 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n14112), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11300) );
  AOI22_X1 U14344 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11299) );
  AOI22_X1 U14346 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11298) );
  NAND4_X1 U14347 ( .A1(n11301), .A2(n11300), .A3(n11299), .A4(n11298), .ZN(
        n11307) );
  AOI22_X1 U14348 ( .A1(n11262), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11305) );
  AOI22_X1 U14349 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11304) );
  AOI22_X1 U14350 ( .A1(n11597), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9725), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11303) );
  AOI22_X1 U14351 ( .A1(n9759), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11302) );
  NAND4_X1 U14352 ( .A1(n11305), .A2(n11304), .A3(n11303), .A4(n11302), .ZN(
        n11306) );
  NAND2_X1 U14353 ( .A1(n11775), .A2(n13805), .ZN(n11309) );
  NAND2_X1 U14354 ( .A1(n11770), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11308) );
  NAND2_X1 U14355 ( .A1(n11309), .A2(n11308), .ZN(n11376) );
  AOI22_X1 U14356 ( .A1(n11262), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11313) );
  AOI22_X1 U14357 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11312) );
  AOI22_X1 U14358 ( .A1(n14112), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11311) );
  AOI22_X1 U14359 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11310) );
  NAND4_X1 U14360 ( .A1(n11313), .A2(n11312), .A3(n11311), .A4(n11310), .ZN(
        n11319) );
  AOI22_X1 U14361 ( .A1(n14118), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n11149), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11317) );
  AOI22_X1 U14362 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11316) );
  INV_X1 U14363 ( .A(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n20991) );
  AOI22_X1 U14364 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9725), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11315) );
  AOI22_X1 U14365 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11314) );
  NAND4_X1 U14366 ( .A1(n11317), .A2(n11316), .A3(n11315), .A4(n11314), .ZN(
        n11318) );
  NAND2_X1 U14367 ( .A1(n11775), .A2(n13808), .ZN(n11321) );
  NAND2_X1 U14368 ( .A1(n11770), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11320) );
  NAND2_X1 U14369 ( .A1(n11321), .A2(n11320), .ZN(n11385) );
  AOI22_X1 U14370 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11149), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11326) );
  AOI22_X1 U14371 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n14112), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11325) );
  AOI22_X1 U14372 ( .A1(n11262), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11324) );
  AOI22_X1 U14373 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11323) );
  NAND4_X1 U14374 ( .A1(n11326), .A2(n11325), .A3(n11324), .A4(n11323), .ZN(
        n11332) );
  AOI22_X1 U14375 ( .A1(n9721), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(n9742), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11330) );
  AOI22_X1 U14376 ( .A1(n14118), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11329) );
  AOI22_X1 U14377 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9725), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11328) );
  AOI22_X1 U14378 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11327) );
  NAND4_X1 U14379 ( .A1(n11330), .A2(n11329), .A3(n11328), .A4(n11327), .ZN(
        n11331) );
  NAND2_X1 U14380 ( .A1(n11775), .A2(n13907), .ZN(n11334) );
  NAND2_X1 U14381 ( .A1(n11770), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11333) );
  NAND2_X1 U14382 ( .A1(n11775), .A2(n13954), .ZN(n11336) );
  NAND2_X1 U14383 ( .A1(n11770), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11335) );
  NAND2_X1 U14384 ( .A1(n11336), .A2(n11335), .ZN(n11337) );
  INV_X1 U14385 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n13822) );
  NOR2_X1 U14386 ( .A1(n11397), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11338) );
  OR2_X1 U14387 ( .A1(n11416), .A2(n11338), .ZN(n19920) );
  NAND2_X1 U14388 ( .A1(n19920), .A2(n14135), .ZN(n11340) );
  NAND2_X1 U14389 ( .A1(n14136), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11339) );
  OAI211_X1 U14390 ( .C1(n11354), .C2(n13822), .A(n11340), .B(n11339), .ZN(
        n11341) );
  AOI21_X1 U14391 ( .B1(n13905), .B2(n11413), .A(n11341), .ZN(n13820) );
  NAND2_X1 U14392 ( .A1(n13517), .A2(n11413), .ZN(n11346) );
  AND2_X1 U14393 ( .A1(n11159), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11379) );
  INV_X1 U14394 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n13580) );
  XNOR2_X1 U14395 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19992) );
  AOI21_X1 U14396 ( .B1(n14135), .B2(n19992), .A(n14136), .ZN(n11343) );
  OAI21_X1 U14397 ( .B1(n11354), .B2(n13580), .A(n11343), .ZN(n11344) );
  AOI21_X1 U14398 ( .B1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n11379), .A(
        n11344), .ZN(n11345) );
  NAND2_X1 U14399 ( .A1(n11346), .A2(n11345), .ZN(n11347) );
  NAND2_X1 U14400 ( .A1(n14136), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11367) );
  NAND2_X1 U14401 ( .A1(n11347), .A2(n11367), .ZN(n13532) );
  AOI21_X1 U14402 ( .B1(n13363), .B2(n11180), .A(n20640), .ZN(n13572) );
  INV_X1 U14403 ( .A(n11351), .ZN(n14145) );
  NAND2_X1 U14404 ( .A1(n14145), .A2(n11413), .ZN(n11357) );
  INV_X1 U14405 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n11353) );
  INV_X1 U14406 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n11352) );
  OAI22_X1 U14407 ( .A1(n11354), .A2(n11353), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n11352), .ZN(n11355) );
  AOI21_X1 U14408 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n11379), .A(
        n11355), .ZN(n11356) );
  NAND2_X1 U14409 ( .A1(n11357), .A2(n11356), .ZN(n13571) );
  NAND2_X1 U14410 ( .A1(n13572), .A2(n13571), .ZN(n13570) );
  INV_X1 U14411 ( .A(n14135), .ZN(n11423) );
  OR2_X1 U14412 ( .A1(n13571), .A2(n11423), .ZN(n11358) );
  NAND2_X1 U14413 ( .A1(n13570), .A2(n11358), .ZN(n13499) );
  INV_X1 U14414 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n11362) );
  INV_X1 U14415 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20930) );
  OAI22_X1 U14416 ( .A1(n11354), .A2(n11362), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20930), .ZN(n11363) );
  AOI21_X1 U14417 ( .B1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n11379), .A(
        n11363), .ZN(n11364) );
  NAND2_X1 U14418 ( .A1(n13499), .A2(n13498), .ZN(n13531) );
  NAND2_X1 U14419 ( .A1(n11366), .A2(n11365), .ZN(n13534) );
  INV_X1 U14420 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n11373) );
  INV_X1 U14421 ( .A(n11378), .ZN(n11371) );
  INV_X1 U14422 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11369) );
  NAND2_X1 U14423 ( .A1(n11369), .A2(n11368), .ZN(n11370) );
  NAND2_X1 U14424 ( .A1(n11371), .A2(n11370), .ZN(n19976) );
  AOI22_X1 U14425 ( .A1(n19976), .A2(n14135), .B1(n14136), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11372) );
  OAI21_X1 U14426 ( .B1(n11354), .B2(n11373), .A(n11372), .ZN(n11374) );
  AOI21_X1 U14427 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n11379), .A(
        n11374), .ZN(n11375) );
  NAND2_X1 U14428 ( .A1(n13575), .A2(n13574), .ZN(n13573) );
  XNOR2_X1 U14429 ( .A(n11377), .B(n11376), .ZN(n13715) );
  OAI21_X1 U14430 ( .B1(n11378), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n11387), .ZN(n19966) );
  INV_X1 U14431 ( .A(n11379), .ZN(n11382) );
  NAND2_X1 U14432 ( .A1(n20640), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11381) );
  NAND2_X1 U14433 ( .A1(n14137), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11380) );
  OAI211_X1 U14434 ( .C1(n11382), .C2(n13484), .A(n11381), .B(n11380), .ZN(
        n11383) );
  MUX2_X1 U14435 ( .A(n19966), .B(n11383), .S(n11423), .Z(n11384) );
  XNOR2_X1 U14436 ( .A(n11386), .B(n11385), .ZN(n13804) );
  NAND2_X1 U14437 ( .A1(n13804), .A2(n11413), .ZN(n11392) );
  AND2_X1 U14438 ( .A1(n11387), .A2(n20884), .ZN(n11388) );
  OR2_X1 U14439 ( .A1(n11388), .A2(n11395), .ZN(n19950) );
  NAND2_X1 U14440 ( .A1(n19950), .A2(n14135), .ZN(n11389) );
  OAI21_X1 U14441 ( .B1(n20884), .B2(n11559), .A(n11389), .ZN(n11390) );
  AOI21_X1 U14442 ( .B1(n14137), .B2(P1_EAX_REG_5__SCAN_IN), .A(n11390), .ZN(
        n11391) );
  NAND2_X1 U14443 ( .A1(n11392), .A2(n11391), .ZN(n13694) );
  NAND2_X1 U14444 ( .A1(n13672), .A2(n13694), .ZN(n13693) );
  NAND2_X1 U14445 ( .A1(n11394), .A2(n11393), .ZN(n13896) );
  INV_X1 U14446 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11399) );
  NOR2_X1 U14447 ( .A1(n11395), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11396) );
  OR2_X1 U14448 ( .A1(n11397), .A2(n11396), .ZN(n19935) );
  AOI22_X1 U14449 ( .A1(n19935), .A2(n14135), .B1(n14136), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11398) );
  OAI21_X1 U14450 ( .B1(n11354), .B2(n11399), .A(n11398), .ZN(n11400) );
  NAND2_X1 U14451 ( .A1(n11404), .A2(n11403), .ZN(n13819) );
  AOI22_X1 U14452 ( .A1(n14112), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11408) );
  AOI22_X1 U14453 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9725), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11407) );
  AOI22_X1 U14454 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11406) );
  AOI22_X1 U14455 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11405) );
  NAND4_X1 U14456 ( .A1(n11408), .A2(n11407), .A3(n11406), .A4(n11405), .ZN(
        n11415) );
  AOI22_X1 U14457 ( .A1(n14118), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11149), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11412) );
  AOI22_X1 U14458 ( .A1(n11262), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11411) );
  AOI22_X1 U14459 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11410) );
  AOI22_X1 U14460 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11409) );
  NAND4_X1 U14461 ( .A1(n11412), .A2(n11411), .A3(n11410), .A4(n11409), .ZN(
        n11414) );
  OAI21_X1 U14462 ( .B1(n11415), .B2(n11414), .A(n11413), .ZN(n11420) );
  NAND2_X1 U14463 ( .A1(n14137), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11419) );
  XNOR2_X1 U14464 ( .A(n11416), .B(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13959) );
  NAND2_X1 U14465 ( .A1(n13959), .A2(n14135), .ZN(n11418) );
  NAND2_X1 U14466 ( .A1(n14136), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11417) );
  NAND4_X1 U14467 ( .A1(n11420), .A2(n11419), .A3(n11418), .A4(n11417), .ZN(
        n13862) );
  XOR2_X1 U14468 ( .A(n13931), .B(n11422), .Z(n14039) );
  AOI22_X1 U14469 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n14118), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11427) );
  AOI22_X1 U14470 ( .A1(n11262), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n14112), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11426) );
  AOI22_X1 U14471 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11425) );
  AOI22_X1 U14472 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11424) );
  NAND4_X1 U14473 ( .A1(n11427), .A2(n11426), .A3(n11425), .A4(n11424), .ZN(
        n11433) );
  AOI22_X1 U14474 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11637), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11431) );
  AOI22_X1 U14475 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n11149), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11430) );
  AOI22_X1 U14476 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n9721), .B1(n9725), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11429) );
  AOI22_X1 U14477 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11428) );
  NAND4_X1 U14478 ( .A1(n11431), .A2(n11430), .A3(n11429), .A4(n11428), .ZN(
        n11432) );
  NOR2_X1 U14479 ( .A1(n11433), .A2(n11432), .ZN(n11434) );
  OAI22_X1 U14480 ( .A1(n11525), .A2(n11434), .B1(n11559), .B2(n13931), .ZN(
        n11436) );
  INV_X1 U14481 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n13937) );
  NOR2_X1 U14482 ( .A1(n11354), .A2(n13937), .ZN(n11435) );
  NOR2_X1 U14483 ( .A1(n11436), .A2(n11435), .ZN(n11437) );
  OAI21_X1 U14484 ( .B1(n14039), .B2(n11423), .A(n11437), .ZN(n13924) );
  XNOR2_X1 U14485 ( .A(n11438), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15908) );
  NAND2_X1 U14486 ( .A1(n15908), .A2(n14135), .ZN(n11454) );
  INV_X1 U14487 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n13998) );
  INV_X1 U14488 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n11439) );
  OAI22_X1 U14489 ( .A1(n11354), .A2(n13998), .B1(n11559), .B2(n11439), .ZN(
        n11452) );
  AOI22_X1 U14490 ( .A1(n14118), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11149), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11443) );
  AOI22_X1 U14491 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n14112), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11442) );
  AOI22_X1 U14492 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11441) );
  AOI22_X1 U14493 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9725), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11440) );
  NAND4_X1 U14494 ( .A1(n11443), .A2(n11442), .A3(n11441), .A4(n11440), .ZN(
        n11449) );
  AOI22_X1 U14495 ( .A1(n11262), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11447) );
  AOI22_X1 U14496 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11446) );
  AOI22_X1 U14497 ( .A1(n9742), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11445) );
  AOI22_X1 U14498 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11444) );
  NAND4_X1 U14499 ( .A1(n11447), .A2(n11446), .A3(n11445), .A4(n11444), .ZN(
        n11448) );
  NOR2_X1 U14500 ( .A1(n11449), .A2(n11448), .ZN(n11450) );
  NOR2_X1 U14501 ( .A1(n11525), .A2(n11450), .ZN(n11451) );
  NOR2_X1 U14502 ( .A1(n11452), .A2(n11451), .ZN(n11453) );
  NAND2_X1 U14503 ( .A1(n11454), .A2(n11453), .ZN(n13995) );
  INV_X1 U14504 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14047) );
  OAI21_X1 U14505 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11455), .A(
        n11478), .ZN(n15967) );
  AOI22_X1 U14506 ( .A1(n14135), .A2(n15967), .B1(n14136), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11456) );
  OAI21_X1 U14507 ( .B1(n11354), .B2(n14047), .A(n11456), .ZN(n14029) );
  AOI22_X1 U14508 ( .A1(n11262), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n14112), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U14509 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11459) );
  AOI22_X1 U14510 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11458) );
  AOI22_X1 U14511 ( .A1(n9742), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11457) );
  NAND4_X1 U14512 ( .A1(n11460), .A2(n11459), .A3(n11458), .A4(n11457), .ZN(
        n11466) );
  AOI22_X1 U14513 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11464) );
  AOI22_X1 U14514 ( .A1(n14118), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11149), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11463) );
  AOI22_X1 U14515 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11462) );
  AOI22_X1 U14516 ( .A1(n9721), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n9725), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11461) );
  NAND4_X1 U14517 ( .A1(n11464), .A2(n11463), .A3(n11462), .A4(n11461), .ZN(
        n11465) );
  NOR2_X1 U14518 ( .A1(n11466), .A2(n11465), .ZN(n11467) );
  NOR2_X1 U14519 ( .A1(n11525), .A2(n11467), .ZN(n14063) );
  AOI22_X1 U14520 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11149), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11471) );
  AOI22_X1 U14521 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n14118), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11470) );
  AOI22_X1 U14522 ( .A1(n14112), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11469) );
  AOI22_X1 U14523 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11468) );
  NAND4_X1 U14524 ( .A1(n11471), .A2(n11470), .A3(n11469), .A4(n11468), .ZN(
        n11477) );
  AOI22_X1 U14525 ( .A1(n11262), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11475) );
  AOI22_X1 U14526 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9725), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11474) );
  AOI22_X1 U14527 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11473) );
  AOI22_X1 U14528 ( .A1(n11616), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n11254), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11472) );
  NAND4_X1 U14529 ( .A1(n11475), .A2(n11474), .A3(n11473), .A4(n11472), .ZN(
        n11476) );
  NOR2_X1 U14530 ( .A1(n11477), .A2(n11476), .ZN(n11482) );
  NAND2_X1 U14531 ( .A1(n14137), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11481) );
  XNOR2_X1 U14532 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11478), .ZN(
        n15959) );
  OAI22_X1 U14533 ( .A1(n15959), .A2(n11423), .B1(n11559), .B2(n15885), .ZN(
        n11479) );
  INV_X1 U14534 ( .A(n11479), .ZN(n11480) );
  OAI211_X1 U14535 ( .C1(n11482), .C2(n11525), .A(n11481), .B(n11480), .ZN(
        n14067) );
  AOI22_X1 U14536 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n11635), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11486) );
  AOI22_X1 U14537 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11485) );
  AOI22_X1 U14538 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11484) );
  AOI22_X1 U14539 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11483) );
  NAND4_X1 U14540 ( .A1(n11486), .A2(n11485), .A3(n11484), .A4(n11483), .ZN(
        n11492) );
  AOI22_X1 U14541 ( .A1(n11262), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11490) );
  AOI22_X1 U14542 ( .A1(n14118), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9725), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11489) );
  AOI22_X1 U14543 ( .A1(n14112), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11488) );
  AOI22_X1 U14544 ( .A1(n11149), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11487) );
  NAND4_X1 U14545 ( .A1(n11490), .A2(n11489), .A3(n11488), .A4(n11487), .ZN(
        n11491) );
  NOR2_X1 U14546 ( .A1(n11492), .A2(n11491), .ZN(n11496) );
  NAND2_X1 U14547 ( .A1(n14137), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11495) );
  XNOR2_X1 U14548 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n11493), .ZN(
        n14554) );
  AOI22_X1 U14549 ( .A1(n14135), .A2(n14554), .B1(n14136), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11494) );
  OAI211_X1 U14550 ( .C1(n11496), .C2(n11525), .A(n11495), .B(n11494), .ZN(
        n14076) );
  XOR2_X1 U14551 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n11497), .Z(
        n15951) );
  AOI22_X1 U14552 ( .A1(n14118), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11149), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11501) );
  AOI22_X1 U14553 ( .A1(n9721), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(n9742), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11500) );
  AOI22_X1 U14554 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11499) );
  AOI22_X1 U14555 ( .A1(n11262), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9725), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11498) );
  NAND4_X1 U14556 ( .A1(n11501), .A2(n11500), .A3(n11499), .A4(n11498), .ZN(
        n11507) );
  AOI22_X1 U14557 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n14112), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11505) );
  AOI22_X1 U14558 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11504) );
  AOI22_X1 U14559 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11254), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11503) );
  AOI22_X1 U14560 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11502) );
  NAND4_X1 U14561 ( .A1(n11505), .A2(n11504), .A3(n11503), .A4(n11502), .ZN(
        n11506) );
  NOR2_X1 U14562 ( .A1(n11507), .A2(n11506), .ZN(n11509) );
  INV_X1 U14563 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n11508) );
  OAI22_X1 U14564 ( .A1(n11525), .A2(n11509), .B1(n11559), .B2(n11508), .ZN(
        n11511) );
  INV_X1 U14565 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n14056) );
  NOR2_X1 U14566 ( .A1(n11354), .A2(n14056), .ZN(n11510) );
  NOR2_X1 U14567 ( .A1(n11511), .A2(n11510), .ZN(n11512) );
  OAI21_X1 U14568 ( .B1(n15951), .B2(n11423), .A(n11512), .ZN(n14052) );
  XNOR2_X1 U14569 ( .A(n11513), .B(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15868) );
  AOI22_X1 U14570 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n14118), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11517) );
  AOI22_X1 U14571 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11516) );
  AOI22_X1 U14572 ( .A1(n11149), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11515) );
  AOI22_X1 U14573 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9725), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11514) );
  NAND4_X1 U14574 ( .A1(n11517), .A2(n11516), .A3(n11515), .A4(n11514), .ZN(
        n11523) );
  AOI22_X1 U14575 ( .A1(n11262), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11521) );
  AOI22_X1 U14576 ( .A1(n14112), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11520) );
  AOI22_X1 U14577 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11519) );
  AOI22_X1 U14578 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11518) );
  NAND4_X1 U14579 ( .A1(n11521), .A2(n11520), .A3(n11519), .A4(n11518), .ZN(
        n11522) );
  NOR2_X1 U14580 ( .A1(n11523), .A2(n11522), .ZN(n11524) );
  OAI22_X1 U14581 ( .A1(n11525), .A2(n11524), .B1(n11559), .B2(n15870), .ZN(
        n11528) );
  INV_X1 U14582 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n11526) );
  NOR2_X1 U14583 ( .A1(n11354), .A2(n11526), .ZN(n11527) );
  NOR2_X1 U14584 ( .A1(n11528), .A2(n11527), .ZN(n11529) );
  OAI21_X1 U14585 ( .B1(n15868), .B2(n11423), .A(n11529), .ZN(n14059) );
  AOI22_X1 U14586 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11635), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11533) );
  AOI22_X1 U14587 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11262), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11532) );
  AOI22_X1 U14588 ( .A1(n14112), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11531) );
  AOI22_X1 U14589 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11530) );
  NAND4_X1 U14590 ( .A1(n11533), .A2(n11532), .A3(n11531), .A4(n11530), .ZN(
        n11539) );
  AOI22_X1 U14591 ( .A1(n14118), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11149), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11537) );
  AOI22_X1 U14592 ( .A1(n9721), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11536) );
  AOI22_X1 U14593 ( .A1(n11616), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9725), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11535) );
  AOI22_X1 U14594 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11534) );
  NAND4_X1 U14595 ( .A1(n11537), .A2(n11536), .A3(n11535), .A4(n11534), .ZN(
        n11538) );
  NOR2_X1 U14596 ( .A1(n11539), .A2(n11538), .ZN(n11544) );
  INV_X1 U14597 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n11541) );
  NAND2_X1 U14598 ( .A1(n20640), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n11540) );
  OAI211_X1 U14599 ( .C1(n11354), .C2(n11541), .A(n11423), .B(n11540), .ZN(
        n11542) );
  INV_X1 U14600 ( .A(n11542), .ZN(n11543) );
  OAI21_X1 U14601 ( .B1(n14130), .B2(n11544), .A(n11543), .ZN(n11547) );
  OAI21_X1 U14602 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n11545), .A(
        n11558), .ZN(n15942) );
  OR2_X1 U14603 ( .A1(n11423), .A2(n15942), .ZN(n11546) );
  NAND2_X1 U14604 ( .A1(n11547), .A2(n11546), .ZN(n14357) );
  AOI22_X1 U14605 ( .A1(n11262), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U14606 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n9742), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11550) );
  AOI22_X1 U14607 ( .A1(n14118), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11254), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11549) );
  AOI22_X1 U14608 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9725), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11548) );
  NAND4_X1 U14609 ( .A1(n11551), .A2(n11550), .A3(n11549), .A4(n11548), .ZN(
        n11557) );
  AOI22_X1 U14610 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n14112), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11555) );
  AOI22_X1 U14611 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11149), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11554) );
  AOI22_X1 U14612 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11553) );
  AOI22_X1 U14613 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11552) );
  NAND4_X1 U14614 ( .A1(n11555), .A2(n11554), .A3(n11553), .A4(n11552), .ZN(
        n11556) );
  OAI21_X1 U14615 ( .B1(n11557), .B2(n11556), .A(n11714), .ZN(n11562) );
  XNOR2_X1 U14616 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n11558), .ZN(
        n15851) );
  OAI22_X1 U14617 ( .A1(n15851), .A2(n11423), .B1(n11559), .B2(n15849), .ZN(
        n11560) );
  AOI21_X1 U14618 ( .B1(n14137), .B2(P1_EAX_REG_17__SCAN_IN), .A(n11560), .ZN(
        n11561) );
  AOI22_X1 U14619 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10968), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11567) );
  AOI22_X1 U14620 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11566) );
  AOI22_X1 U14621 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11565) );
  AOI22_X1 U14622 ( .A1(n14112), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11564) );
  NAND4_X1 U14623 ( .A1(n11567), .A2(n11566), .A3(n11565), .A4(n11564), .ZN(
        n11573) );
  AOI22_X1 U14624 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11571) );
  AOI22_X1 U14625 ( .A1(n11262), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9725), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11570) );
  AOI22_X1 U14626 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11569) );
  AOI22_X1 U14627 ( .A1(n11149), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11254), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11568) );
  NAND4_X1 U14628 ( .A1(n11571), .A2(n11570), .A3(n11569), .A4(n11568), .ZN(
        n11572) );
  NOR2_X1 U14629 ( .A1(n11573), .A2(n11572), .ZN(n11577) );
  INV_X1 U14630 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n14410) );
  NAND2_X1 U14631 ( .A1(n20640), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11574) );
  OAI211_X1 U14632 ( .C1(n11354), .C2(n14410), .A(n11423), .B(n11574), .ZN(
        n11575) );
  INV_X1 U14633 ( .A(n11575), .ZN(n11576) );
  OAI21_X1 U14634 ( .B1(n14130), .B2(n11577), .A(n11576), .ZN(n11580) );
  OAI21_X1 U14635 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n11578), .A(
        n11594), .ZN(n15933) );
  OR2_X1 U14636 ( .A1(n11423), .A2(n15933), .ZN(n11579) );
  NAND2_X1 U14637 ( .A1(n11580), .A2(n11579), .ZN(n14408) );
  AOI22_X1 U14638 ( .A1(n11262), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11584) );
  AOI22_X1 U14639 ( .A1(n9721), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(n9742), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11583) );
  AOI22_X1 U14640 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11582) );
  AOI22_X1 U14641 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9725), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11581) );
  NAND4_X1 U14642 ( .A1(n11584), .A2(n11583), .A3(n11582), .A4(n11581), .ZN(
        n11590) );
  AOI22_X1 U14643 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n14112), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11588) );
  AOI22_X1 U14644 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n14118), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11587) );
  AOI22_X1 U14645 ( .A1(n11149), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11254), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11586) );
  AOI22_X1 U14646 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11585) );
  NAND4_X1 U14647 ( .A1(n11588), .A2(n11587), .A3(n11586), .A4(n11585), .ZN(
        n11589) );
  NOR2_X1 U14648 ( .A1(n11590), .A2(n11589), .ZN(n11593) );
  OAI21_X1 U14649 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15831), .A(n11423), 
        .ZN(n11591) );
  AOI21_X1 U14650 ( .B1(n14137), .B2(P1_EAX_REG_19__SCAN_IN), .A(n11591), .ZN(
        n11592) );
  OAI21_X1 U14651 ( .B1(n14130), .B2(n11593), .A(n11592), .ZN(n11596) );
  XNOR2_X1 U14652 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n11594), .ZN(
        n15837) );
  NAND2_X1 U14653 ( .A1(n15837), .A2(n14135), .ZN(n11595) );
  AOI22_X1 U14654 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11601) );
  AOI22_X1 U14655 ( .A1(n14112), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11600) );
  AOI22_X1 U14656 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11254), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11599) );
  AOI22_X1 U14657 ( .A1(n11597), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9749), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11598) );
  NAND4_X1 U14658 ( .A1(n11601), .A2(n11600), .A3(n11599), .A4(n11598), .ZN(
        n11607) );
  AOI22_X1 U14659 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11149), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11605) );
  AOI22_X1 U14660 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n14119), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U14661 ( .A1(n14118), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11603) );
  AOI22_X1 U14662 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11602) );
  NAND4_X1 U14663 ( .A1(n11605), .A2(n11604), .A3(n11603), .A4(n11602), .ZN(
        n11606) );
  NOR2_X1 U14664 ( .A1(n11607), .A2(n11606), .ZN(n11612) );
  INV_X1 U14665 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n11609) );
  NAND2_X1 U14666 ( .A1(n20640), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11608) );
  OAI211_X1 U14667 ( .C1(n11354), .C2(n11609), .A(n11423), .B(n11608), .ZN(
        n11610) );
  INV_X1 U14668 ( .A(n11610), .ZN(n11611) );
  OAI21_X1 U14669 ( .B1(n14130), .B2(n11612), .A(n11611), .ZN(n11615) );
  OAI21_X1 U14670 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n11613), .A(
        n11630), .ZN(n15921) );
  OR2_X1 U14671 ( .A1(n11423), .A2(n15921), .ZN(n11614) );
  AOI22_X1 U14672 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11149), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11620) );
  AOI22_X1 U14673 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n14112), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11619) );
  AOI22_X1 U14674 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U14675 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11616), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11617) );
  NAND4_X1 U14676 ( .A1(n11620), .A2(n11619), .A3(n11618), .A4(n11617), .ZN(
        n11626) );
  AOI22_X1 U14677 ( .A1(n9721), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11624) );
  AOI22_X1 U14678 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9750), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11623) );
  AOI22_X1 U14679 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11622) );
  AOI22_X1 U14680 ( .A1(n14118), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11621) );
  NAND4_X1 U14681 ( .A1(n11624), .A2(n11623), .A3(n11622), .A4(n11621), .ZN(
        n11625) );
  NOR2_X1 U14682 ( .A1(n11626), .A2(n11625), .ZN(n11629) );
  OAI21_X1 U14683 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20853), .A(n11423), 
        .ZN(n11627) );
  AOI21_X1 U14684 ( .B1(n14137), .B2(P1_EAX_REG_21__SCAN_IN), .A(n11627), .ZN(
        n11628) );
  OAI21_X1 U14685 ( .B1(n14130), .B2(n11629), .A(n11628), .ZN(n11634) );
  INV_X1 U14686 ( .A(n11630), .ZN(n11632) );
  INV_X1 U14687 ( .A(n11631), .ZN(n11654) );
  OAI21_X1 U14688 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n11632), .A(
        n11654), .ZN(n15812) );
  OR2_X1 U14689 ( .A1(n11423), .A2(n15812), .ZN(n11633) );
  NAND2_X1 U14690 ( .A1(n11634), .A2(n11633), .ZN(n14324) );
  AOI22_X1 U14691 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11641) );
  AOI22_X1 U14692 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11636), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11640) );
  AOI22_X1 U14693 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9721), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11639) );
  AOI22_X1 U14694 ( .A1(n11616), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11638) );
  NAND4_X1 U14695 ( .A1(n11641), .A2(n11640), .A3(n11639), .A4(n11638), .ZN(
        n11649) );
  AOI22_X1 U14696 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11149), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11647) );
  AOI22_X1 U14697 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n14118), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11646) );
  AOI22_X1 U14698 ( .A1(n14112), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9749), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11645) );
  AOI22_X1 U14699 ( .A1(n9742), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11642), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11644) );
  NAND4_X1 U14700 ( .A1(n11647), .A2(n11646), .A3(n11645), .A4(n11644), .ZN(
        n11648) );
  NOR2_X1 U14701 ( .A1(n11649), .A2(n11648), .ZN(n11653) );
  INV_X1 U14702 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n14394) );
  NAND2_X1 U14703 ( .A1(n20640), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11650) );
  OAI211_X1 U14704 ( .C1(n11354), .C2(n14394), .A(n11423), .B(n11650), .ZN(
        n11651) );
  INV_X1 U14705 ( .A(n11651), .ZN(n11652) );
  OAI21_X1 U14706 ( .B1(n14130), .B2(n11653), .A(n11652), .ZN(n11658) );
  INV_X1 U14707 ( .A(n11664), .ZN(n11656) );
  INV_X1 U14708 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15799) );
  NAND2_X1 U14709 ( .A1(n15799), .A2(n11654), .ZN(n11655) );
  NAND2_X1 U14710 ( .A1(n11656), .A2(n11655), .ZN(n15807) );
  NAND2_X1 U14711 ( .A1(n11658), .A2(n11657), .ZN(n14391) );
  XOR2_X1 U14712 ( .A(n11661), .B(n11660), .Z(n11662) );
  NAND2_X1 U14713 ( .A1(n11662), .A2(n11714), .ZN(n11667) );
  INV_X1 U14714 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15795) );
  OAI21_X1 U14715 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15795), .A(n11423), 
        .ZN(n11663) );
  AOI21_X1 U14716 ( .B1(n14137), .B2(P1_EAX_REG_23__SCAN_IN), .A(n11663), .ZN(
        n11666) );
  XNOR2_X1 U14717 ( .A(n11664), .B(n15795), .ZN(n15792) );
  AND2_X1 U14718 ( .A1(n15792), .A2(n14135), .ZN(n11665) );
  AOI21_X1 U14719 ( .B1(n11667), .B2(n11666), .A(n11665), .ZN(n14318) );
  INV_X1 U14720 ( .A(n11668), .ZN(n11669) );
  NAND2_X1 U14721 ( .A1(n11669), .A2(n20793), .ZN(n11670) );
  NAND2_X1 U14722 ( .A1(n11685), .A2(n11670), .ZN(n15782) );
  XNOR2_X1 U14723 ( .A(n11672), .B(n11671), .ZN(n11675) );
  INV_X1 U14724 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n14381) );
  NOR2_X1 U14725 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n20906), .ZN(
        n20988) );
  OAI22_X1 U14726 ( .A1(n11354), .A2(n14381), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20988), .ZN(n11673) );
  INV_X1 U14727 ( .A(n11673), .ZN(n11674) );
  OAI21_X1 U14728 ( .B1(n11675), .B2(n14130), .A(n11674), .ZN(n11676) );
  OAI21_X1 U14729 ( .B1(n11423), .B2(n15782), .A(n11676), .ZN(n14313) );
  XOR2_X1 U14730 ( .A(n11678), .B(n11677), .Z(n11679) );
  NAND2_X1 U14731 ( .A1(n11679), .A2(n11714), .ZN(n11684) );
  INV_X1 U14732 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n11681) );
  OAI21_X1 U14733 ( .B1(n20906), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n20579), .ZN(n11680) );
  OAI21_X1 U14734 ( .B1(n11354), .B2(n11681), .A(n11680), .ZN(n11682) );
  INV_X1 U14735 ( .A(n11682), .ZN(n11683) );
  NAND2_X1 U14736 ( .A1(n11684), .A2(n11683), .ZN(n11687) );
  XNOR2_X1 U14737 ( .A(n11685), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14487) );
  NAND2_X1 U14738 ( .A1(n14487), .A2(n14135), .ZN(n11686) );
  NAND2_X1 U14739 ( .A1(n11687), .A2(n11686), .ZN(n14284) );
  INV_X1 U14740 ( .A(n11689), .ZN(n11690) );
  XNOR2_X1 U14741 ( .A(n11691), .B(n11690), .ZN(n11694) );
  INV_X1 U14742 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14374) );
  NAND2_X1 U14743 ( .A1(n20640), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11692) );
  OAI211_X1 U14744 ( .C1(n11354), .C2(n14374), .A(n11423), .B(n11692), .ZN(
        n11693) );
  AOI21_X1 U14745 ( .B1(n11694), .B2(n11714), .A(n11693), .ZN(n11698) );
  NAND2_X1 U14746 ( .A1(n11695), .A2(n14275), .ZN(n11696) );
  NAND2_X1 U14747 ( .A1(n11705), .A2(n11696), .ZN(n14474) );
  NOR2_X1 U14748 ( .A1(n14474), .A2(n11423), .ZN(n11697) );
  XOR2_X1 U14749 ( .A(n11700), .B(n11699), .Z(n11701) );
  NAND2_X1 U14750 ( .A1(n11701), .A2(n11714), .ZN(n11708) );
  INV_X1 U14751 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n11703) );
  OAI21_X1 U14752 ( .B1(n20906), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n20579), .ZN(n11702) );
  OAI21_X1 U14753 ( .B1(n11354), .B2(n11703), .A(n11702), .ZN(n11704) );
  INV_X1 U14754 ( .A(n11704), .ZN(n11707) );
  XNOR2_X1 U14755 ( .A(n11705), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14468) );
  AOI21_X1 U14756 ( .B1(n11708), .B2(n11707), .A(n11706), .ZN(n14258) );
  NAND2_X1 U14757 ( .A1(n14255), .A2(n14258), .ZN(n14240) );
  INV_X1 U14758 ( .A(n11709), .ZN(n11710) );
  XNOR2_X1 U14759 ( .A(n11711), .B(n11710), .ZN(n11715) );
  INV_X1 U14760 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n14366) );
  NAND2_X1 U14761 ( .A1(n20640), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11712) );
  OAI211_X1 U14762 ( .C1(n11354), .C2(n14366), .A(n11423), .B(n11712), .ZN(
        n11713) );
  AOI21_X1 U14763 ( .B1(n11715), .B2(n11714), .A(n11713), .ZN(n11720) );
  NAND2_X1 U14764 ( .A1(n11717), .A2(n11716), .ZN(n11718) );
  NAND2_X1 U14765 ( .A1(n13739), .A2(n11718), .ZN(n14455) );
  NOR2_X1 U14766 ( .A1(n14455), .A2(n11423), .ZN(n11719) );
  INV_X1 U14767 ( .A(n11722), .ZN(n14241) );
  INV_X1 U14768 ( .A(n11723), .ZN(n11721) );
  INV_X1 U14769 ( .A(n14441), .ZN(n14365) );
  NAND2_X1 U14770 ( .A1(n20414), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11725) );
  NAND2_X1 U14771 ( .A1(n14718), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11724) );
  NAND2_X1 U14772 ( .A1(n11725), .A2(n11724), .ZN(n11740) );
  NAND2_X1 U14773 ( .A1(n20487), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11729) );
  NAND2_X1 U14774 ( .A1(n10921), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11726) );
  NAND2_X1 U14775 ( .A1(n11729), .A2(n11726), .ZN(n11748) );
  INV_X1 U14776 ( .A(n11748), .ZN(n11727) );
  AOI222_X1 U14777 ( .A1(n11767), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .B1(n11767), .B2(n13484), .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .C2(n13484), .ZN(n13160) );
  INV_X1 U14778 ( .A(n11775), .ZN(n11737) );
  OAI21_X1 U14779 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20517), .A(
        n11739), .ZN(n11731) );
  NOR2_X1 U14780 ( .A1(n11737), .A2(n11731), .ZN(n11735) );
  NAND2_X1 U14781 ( .A1(n14185), .A2(n13751), .ZN(n13643) );
  NOR2_X1 U14782 ( .A1(n11764), .A2(n13643), .ZN(n11776) );
  INV_X1 U14783 ( .A(n11731), .ZN(n11732) );
  OAI21_X1 U14784 ( .B1(n11733), .B2(n11249), .A(n11732), .ZN(n11734) );
  AND2_X1 U14785 ( .A1(n20120), .A2(n14185), .ZN(n11738) );
  OR2_X1 U14786 ( .A1(n11738), .A2(n11184), .ZN(n11762) );
  OAI22_X1 U14787 ( .A1(n11735), .A2(n11776), .B1(n11734), .B2(n11762), .ZN(
        n11746) );
  NAND2_X1 U14788 ( .A1(n20139), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11736) );
  NAND2_X1 U14789 ( .A1(n11737), .A2(n11736), .ZN(n11744) );
  INV_X1 U14790 ( .A(n11738), .ZN(n11743) );
  NAND2_X1 U14791 ( .A1(n11740), .A2(n11739), .ZN(n11741) );
  NAND2_X1 U14792 ( .A1(n11742), .A2(n11741), .ZN(n13156) );
  AOI22_X1 U14793 ( .A1(n11744), .A2(n11743), .B1(n11770), .B2(n13156), .ZN(
        n11747) );
  INV_X1 U14794 ( .A(n11744), .ZN(n11745) );
  NAND2_X1 U14795 ( .A1(n11745), .A2(n13751), .ZN(n11769) );
  OAI211_X1 U14796 ( .C1(n11746), .C2(n11747), .A(n11769), .B(n13156), .ZN(
        n11756) );
  NAND2_X1 U14797 ( .A1(n11747), .A2(n11746), .ZN(n11755) );
  NAND2_X1 U14798 ( .A1(n11749), .A2(n11748), .ZN(n11751) );
  NAND2_X1 U14799 ( .A1(n11751), .A2(n11750), .ZN(n13157) );
  INV_X1 U14800 ( .A(n13157), .ZN(n11753) );
  INV_X1 U14801 ( .A(n11762), .ZN(n11752) );
  NAND2_X1 U14802 ( .A1(n11775), .A2(n11753), .ZN(n11761) );
  OAI211_X1 U14803 ( .C1(n11753), .C2(n11764), .A(n11752), .B(n11761), .ZN(
        n11754) );
  NAND3_X1 U14804 ( .A1(n11756), .A2(n11755), .A3(n11754), .ZN(n11766) );
  AOI21_X1 U14805 ( .B1(n11759), .B2(n11758), .A(n11757), .ZN(n11760) );
  INV_X1 U14806 ( .A(n11760), .ZN(n13158) );
  INV_X1 U14807 ( .A(n11761), .ZN(n11763) );
  AOI22_X1 U14808 ( .A1(n13158), .A2(n13904), .B1(n11763), .B2(n11762), .ZN(
        n11765) );
  AOI22_X1 U14809 ( .A1(n11766), .A2(n11765), .B1(n11764), .B2(n13158), .ZN(
        n11772) );
  AND2_X1 U14810 ( .A1(n13484), .A2(n11767), .ZN(n11768) );
  NAND2_X1 U14811 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n11768), .ZN(
        n13159) );
  NOR2_X1 U14812 ( .A1(n13159), .A2(n11769), .ZN(n11771) );
  OAI22_X1 U14813 ( .A1(n11772), .A2(n11771), .B1(n11770), .B2(n13159), .ZN(
        n11773) );
  OAI21_X1 U14814 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n13484), .A(n11773), 
        .ZN(n11774) );
  AOI21_X1 U14815 ( .B1(n11775), .B2(n13160), .A(n11774), .ZN(n11778) );
  AND2_X1 U14816 ( .A1(n13160), .A2(n11776), .ZN(n11777) );
  NOR2_X1 U14817 ( .A1(n13196), .A2(n20120), .ZN(n11779) );
  NAND2_X1 U14818 ( .A1(n13436), .A2(n11779), .ZN(n13376) );
  NOR2_X1 U14819 ( .A1(n11780), .A2(n11249), .ZN(n13400) );
  INV_X1 U14820 ( .A(n13400), .ZN(n11781) );
  NAND2_X1 U14821 ( .A1(n15727), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19884) );
  NOR2_X1 U14822 ( .A1(n14185), .A2(n19884), .ZN(n11784) );
  NOR2_X1 U14823 ( .A1(n13568), .A2(n11167), .ZN(n11783) );
  NAND4_X1 U14824 ( .A1(n13470), .A2(n11784), .A3(n11783), .A4(n11782), .ZN(
        n13563) );
  OR2_X1 U14825 ( .A1(n13563), .A2(n14206), .ZN(n11785) );
  OAI21_X4 U14826 ( .B1(n13453), .B2(n19884), .A(n11785), .ZN(n14350) );
  NAND2_X2 U14827 ( .A1(n14350), .A2(n13568), .ZN(n14359) );
  MUX2_X1 U14828 ( .A(n11823), .B(n11879), .S(P1_EBX_REG_1__SCAN_IN), .Z(
        n11789) );
  INV_X1 U14829 ( .A(n13360), .ZN(n20130) );
  NAND2_X1 U14830 ( .A1(n20130), .A2(n13748), .ZN(n11803) );
  INV_X1 U14831 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13553) );
  NAND2_X1 U14832 ( .A1(n13702), .A2(n13553), .ZN(n11788) );
  NAND2_X1 U14833 ( .A1(n11789), .A2(n11788), .ZN(n11793) );
  INV_X1 U14834 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n11790) );
  OR2_X1 U14835 ( .A1(n11803), .A2(n11790), .ZN(n11792) );
  NAND2_X1 U14836 ( .A1(n14191), .A2(n11790), .ZN(n11791) );
  NAND2_X1 U14837 ( .A1(n11792), .A2(n11791), .ZN(n13703) );
  XNOR2_X1 U14838 ( .A(n11793), .B(n13703), .ZN(n13407) );
  NAND2_X1 U14839 ( .A1(n13407), .A2(n13381), .ZN(n11795) );
  INV_X1 U14840 ( .A(n11793), .ZN(n11794) );
  MUX2_X1 U14841 ( .A(n11883), .B(n14191), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n11797) );
  NOR2_X1 U14842 ( .A1(n14207), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11796) );
  NOR2_X1 U14843 ( .A1(n11797), .A2(n11796), .ZN(n13550) );
  INV_X1 U14844 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13871) );
  NAND2_X1 U14845 ( .A1(n11878), .A2(n13871), .ZN(n11801) );
  INV_X1 U14846 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13660) );
  NAND2_X1 U14847 ( .A1(n11803), .A2(n13660), .ZN(n11799) );
  NAND2_X1 U14848 ( .A1(n13381), .A2(n13871), .ZN(n11798) );
  NAND3_X1 U14849 ( .A1(n11799), .A2(n11879), .A3(n11798), .ZN(n11800) );
  AND2_X1 U14850 ( .A1(n11801), .A2(n11800), .ZN(n13652) );
  INV_X1 U14851 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n11802) );
  NAND2_X1 U14852 ( .A1(n11883), .A2(n11802), .ZN(n11806) );
  INV_X1 U14853 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20073) );
  NAND2_X1 U14854 ( .A1(n13381), .A2(n11802), .ZN(n11804) );
  OAI211_X1 U14855 ( .C1(n14191), .C2(n20073), .A(n11804), .B(n11803), .ZN(
        n11805) );
  NAND2_X1 U14856 ( .A1(n11806), .A2(n11805), .ZN(n13849) );
  INV_X1 U14857 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13812) );
  OAI21_X1 U14858 ( .B1(n14191), .B2(n13812), .A(n11803), .ZN(n11808) );
  INV_X1 U14859 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n19940) );
  NAND2_X1 U14860 ( .A1(n13381), .A2(n19940), .ZN(n11807) );
  NAND2_X1 U14861 ( .A1(n11808), .A2(n11807), .ZN(n11809) );
  OAI21_X1 U14862 ( .B1(P1_EBX_REG_5__SCAN_IN), .B2(n11888), .A(n11809), .ZN(
        n13814) );
  INV_X1 U14863 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n20007) );
  NAND2_X1 U14864 ( .A1(n11883), .A2(n20007), .ZN(n11812) );
  INV_X1 U14865 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16059) );
  NAND2_X1 U14866 ( .A1(n13381), .A2(n20007), .ZN(n11810) );
  OAI211_X1 U14867 ( .C1(n14191), .C2(n16059), .A(n11810), .B(n11803), .ZN(
        n11811) );
  INV_X1 U14868 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16044) );
  OAI21_X1 U14869 ( .B1(n14191), .B2(n16044), .A(n11803), .ZN(n11813) );
  OAI21_X1 U14870 ( .B1(P1_EBX_REG_7__SCAN_IN), .B2(n14206), .A(n11813), .ZN(
        n11815) );
  INV_X1 U14871 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n19912) );
  NAND2_X1 U14872 ( .A1(n11878), .A2(n19912), .ZN(n11814) );
  INV_X1 U14873 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13876) );
  NAND2_X1 U14874 ( .A1(n11883), .A2(n13876), .ZN(n11818) );
  INV_X1 U14875 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16045) );
  NAND2_X1 U14876 ( .A1(n13381), .A2(n13876), .ZN(n11816) );
  OAI211_X1 U14877 ( .C1(n14191), .C2(n16045), .A(n11816), .B(n11803), .ZN(
        n11817) );
  NAND2_X1 U14878 ( .A1(n11818), .A2(n11817), .ZN(n13865) );
  INV_X1 U14879 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n14158) );
  OAI21_X1 U14880 ( .B1(n14191), .B2(n14158), .A(n11803), .ZN(n11821) );
  INV_X1 U14881 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n11819) );
  NAND2_X1 U14882 ( .A1(n13381), .A2(n11819), .ZN(n11820) );
  NAND2_X1 U14883 ( .A1(n11821), .A2(n11820), .ZN(n11822) );
  OAI21_X1 U14884 ( .B1(P1_EBX_REG_9__SCAN_IN), .B2(n11888), .A(n11822), .ZN(
        n13926) );
  MUX2_X1 U14885 ( .A(n11823), .B(n11879), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n11825) );
  INV_X1 U14886 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16038) );
  NAND2_X1 U14887 ( .A1(n13702), .A2(n16038), .ZN(n11824) );
  NAND2_X1 U14888 ( .A1(n11825), .A2(n11824), .ZN(n14012) );
  INV_X1 U14889 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14034) );
  NAND2_X1 U14890 ( .A1(n11878), .A2(n14034), .ZN(n11829) );
  NAND2_X1 U14891 ( .A1(n11803), .A2(n14711), .ZN(n11827) );
  NAND2_X1 U14892 ( .A1(n13381), .A2(n14034), .ZN(n11826) );
  NAND3_X1 U14893 ( .A1(n11827), .A2(n11879), .A3(n11826), .ZN(n11828) );
  INV_X1 U14894 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15884) );
  NAND2_X1 U14895 ( .A1(n11883), .A2(n15884), .ZN(n11832) );
  INV_X1 U14896 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16022) );
  NAND2_X1 U14897 ( .A1(n13381), .A2(n15884), .ZN(n11830) );
  OAI211_X1 U14898 ( .C1(n14191), .C2(n16022), .A(n11830), .B(n11803), .ZN(
        n11831) );
  NAND2_X1 U14899 ( .A1(n11832), .A2(n11831), .ZN(n14072) );
  INV_X1 U14900 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14563) );
  NAND2_X1 U14901 ( .A1(n11803), .A2(n14563), .ZN(n11834) );
  INV_X1 U14902 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14083) );
  NAND2_X1 U14903 ( .A1(n13381), .A2(n14083), .ZN(n11833) );
  NAND3_X1 U14904 ( .A1(n11834), .A2(n11879), .A3(n11833), .ZN(n11835) );
  OAI21_X1 U14905 ( .B1(n11888), .B2(P1_EBX_REG_13__SCAN_IN), .A(n11835), .ZN(
        n14079) );
  INV_X1 U14906 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16009) );
  NAND2_X1 U14907 ( .A1(n16009), .A2(n13702), .ZN(n11837) );
  MUX2_X1 U14908 ( .A(n11823), .B(n11879), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n11836) );
  NAND2_X1 U14909 ( .A1(n11837), .A2(n11836), .ZN(n14054) );
  MUX2_X1 U14910 ( .A(n11823), .B(n11879), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n11839) );
  INV_X1 U14911 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14521) );
  NAND2_X1 U14912 ( .A1(n14521), .A2(n13702), .ZN(n11838) );
  AND2_X1 U14913 ( .A1(n11839), .A2(n11838), .ZN(n14353) );
  INV_X1 U14914 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14165) );
  OAI21_X1 U14915 ( .B1(n14191), .B2(n14165), .A(n11803), .ZN(n11841) );
  INV_X1 U14916 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n11842) );
  NAND2_X1 U14917 ( .A1(n13381), .A2(n11842), .ZN(n11840) );
  NAND2_X1 U14918 ( .A1(n11841), .A2(n11840), .ZN(n11844) );
  NAND2_X1 U14919 ( .A1(n11878), .A2(n11842), .ZN(n11843) );
  NAND2_X1 U14920 ( .A1(n11844), .A2(n11843), .ZN(n14354) );
  INV_X1 U14921 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n14688) );
  NAND2_X1 U14922 ( .A1(n11803), .A2(n14688), .ZN(n11846) );
  INV_X1 U14923 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n15848) );
  NAND2_X1 U14924 ( .A1(n13381), .A2(n15848), .ZN(n11845) );
  NAND3_X1 U14925 ( .A1(n11846), .A2(n11879), .A3(n11845), .ZN(n11847) );
  OAI21_X1 U14926 ( .B1(n11888), .B2(P1_EBX_REG_17__SCAN_IN), .A(n11847), .ZN(
        n14348) );
  INV_X1 U14927 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n15920) );
  NAND2_X1 U14928 ( .A1(n11883), .A2(n15920), .ZN(n11850) );
  NAND2_X1 U14929 ( .A1(n13381), .A2(n15920), .ZN(n11848) );
  OAI211_X1 U14930 ( .C1(n14191), .C2(n14175), .A(n11848), .B(n11803), .ZN(
        n11849) );
  INV_X1 U14931 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15749) );
  OAI21_X1 U14932 ( .B1(n14191), .B2(n15749), .A(n11803), .ZN(n11851) );
  OAI21_X1 U14933 ( .B1(P1_EBX_REG_19__SCAN_IN), .B2(n14206), .A(n11851), .ZN(
        n11854) );
  INV_X1 U14934 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n11852) );
  NAND2_X1 U14935 ( .A1(n11878), .A2(n11852), .ZN(n11853) );
  AND2_X1 U14936 ( .A1(n11854), .A2(n11853), .ZN(n14342) );
  INV_X1 U14937 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n11855) );
  NAND2_X1 U14938 ( .A1(n11883), .A2(n11855), .ZN(n11858) );
  INV_X1 U14939 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15753) );
  NAND2_X1 U14940 ( .A1(n11786), .A2(n11855), .ZN(n11856) );
  OAI211_X1 U14941 ( .C1(n14191), .C2(n15753), .A(n11856), .B(n11803), .ZN(
        n11857) );
  NAND2_X1 U14942 ( .A1(n11858), .A2(n11857), .ZN(n14336) );
  INV_X1 U14943 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15809) );
  NAND2_X1 U14944 ( .A1(n11878), .A2(n15809), .ZN(n11862) );
  INV_X1 U14945 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n14675) );
  NAND2_X1 U14946 ( .A1(n11803), .A2(n14675), .ZN(n11860) );
  NAND2_X1 U14947 ( .A1(n13381), .A2(n15809), .ZN(n11859) );
  NAND3_X1 U14948 ( .A1(n11860), .A2(n11879), .A3(n11859), .ZN(n11861) );
  AND2_X1 U14949 ( .A1(n11862), .A2(n11861), .ZN(n14326) );
  INV_X1 U14950 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15918) );
  NAND2_X1 U14951 ( .A1(n11883), .A2(n15918), .ZN(n11865) );
  INV_X1 U14952 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14667) );
  NAND2_X1 U14953 ( .A1(n13381), .A2(n15918), .ZN(n11863) );
  OAI211_X1 U14954 ( .C1(n14191), .C2(n14667), .A(n11863), .B(n11803), .ZN(
        n11864) );
  AND2_X1 U14955 ( .A1(n11865), .A2(n11864), .ZN(n14659) );
  INV_X1 U14956 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n11866) );
  NAND2_X1 U14957 ( .A1(n11878), .A2(n11866), .ZN(n11870) );
  INV_X1 U14958 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n20956) );
  NAND2_X1 U14959 ( .A1(n11803), .A2(n20956), .ZN(n11868) );
  NAND2_X1 U14960 ( .A1(n13381), .A2(n11866), .ZN(n11867) );
  NAND3_X1 U14961 ( .A1(n11868), .A2(n11879), .A3(n11867), .ZN(n11869) );
  AND2_X1 U14962 ( .A1(n11870), .A2(n11869), .ZN(n14320) );
  MUX2_X1 U14963 ( .A(n11823), .B(n11879), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n11871) );
  OAI21_X1 U14964 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14207), .A(
        n11871), .ZN(n14315) );
  INV_X1 U14965 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14635) );
  NAND2_X1 U14966 ( .A1(n11803), .A2(n14635), .ZN(n11874) );
  INV_X1 U14967 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n11872) );
  NAND2_X1 U14968 ( .A1(n13381), .A2(n11872), .ZN(n11873) );
  NAND3_X1 U14969 ( .A1(n11874), .A2(n11879), .A3(n11873), .ZN(n11875) );
  OAI21_X1 U14970 ( .B1(n11888), .B2(P1_EBX_REG_25__SCAN_IN), .A(n11875), .ZN(
        n14291) );
  MUX2_X1 U14971 ( .A(n11823), .B(n11879), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n11876) );
  OAI21_X1 U14972 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n14207), .A(
        n11876), .ZN(n14273) );
  INV_X1 U14973 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n11877) );
  NAND2_X1 U14974 ( .A1(n11878), .A2(n11877), .ZN(n11882) );
  INV_X1 U14975 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14462) );
  NAND2_X1 U14976 ( .A1(n11803), .A2(n14462), .ZN(n11880) );
  OAI211_X1 U14977 ( .C1(P1_EBX_REG_27__SCAN_IN), .C2(n14206), .A(n11880), .B(
        n11879), .ZN(n11881) );
  AND2_X1 U14978 ( .A1(n11882), .A2(n11881), .ZN(n14266) );
  MUX2_X1 U14979 ( .A(n11883), .B(n14191), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n11885) );
  NOR2_X1 U14980 ( .A1(n14207), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n11884) );
  NOR2_X1 U14981 ( .A1(n11885), .A2(n11884), .ZN(n14250) );
  OR2_X1 U14982 ( .A1(n14207), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11887) );
  INV_X1 U14983 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n20969) );
  NAND2_X1 U14984 ( .A1(n13381), .A2(n20969), .ZN(n11886) );
  NAND2_X1 U14985 ( .A1(n11887), .A2(n11886), .ZN(n14189) );
  OAI22_X1 U14986 ( .A1(n14189), .A2(n14191), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n11888), .ZN(n11889) );
  OR2_X1 U14987 ( .A1(n14248), .A2(n11889), .ZN(n11890) );
  NAND2_X1 U14988 ( .A1(n14204), .A2(n11890), .ZN(n14599) );
  NOR2_X1 U14989 ( .A1(n14350), .A2(n20969), .ZN(n11891) );
  AOI21_X1 U14990 ( .B1(n11893), .B2(n11892), .A(n11891), .ZN(n11894) );
  XNOR2_X2 U14991 ( .A(n11898), .B(n11897), .ZN(n11916) );
  NOR2_X2 U14992 ( .A1(n13777), .A2(n11916), .ZN(n11922) );
  INV_X1 U14993 ( .A(n11899), .ZN(n11905) );
  XNOR2_X2 U14994 ( .A(n11908), .B(n11905), .ZN(n15568) );
  INV_X1 U14995 ( .A(n15568), .ZN(n13258) );
  INV_X1 U14996 ( .A(n11918), .ZN(n11906) );
  INV_X2 U14997 ( .A(n11960), .ZN(n12011) );
  AOI22_X1 U14998 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12002), .B1(
        n12011), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11914) );
  INV_X1 U14999 ( .A(n11916), .ZN(n11907) );
  NOR2_X2 U15000 ( .A1(n13777), .A2(n11907), .ZN(n11920) );
  INV_X1 U15001 ( .A(n11908), .ZN(n11909) );
  NAND2_X1 U15003 ( .A1(n13777), .A2(n11907), .ZN(n11927) );
  NAND2_X1 U15004 ( .A1(n11919), .A2(n11917), .ZN(n11957) );
  AOI22_X1 U15005 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n11999), .B1(
        n12000), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11925) );
  AOI22_X1 U15006 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19353), .B1(
        n15614), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11924) );
  INV_X1 U15007 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11930) );
  INV_X1 U15008 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n20813) );
  OAI22_X1 U15009 ( .A1(n11930), .A2(n19494), .B1(n19601), .B2(n20813), .ZN(
        n11931) );
  NAND2_X1 U15010 ( .A1(n11933), .A2(n19869), .ZN(n11934) );
  INV_X1 U15011 ( .A(n12010), .ZN(n12031) );
  INV_X1 U15012 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13839) );
  NAND2_X1 U15013 ( .A1(n12000), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11938) );
  OAI211_X1 U15014 ( .C1(n12031), .C2(n13839), .A(n11938), .B(n9743), .ZN(
        n11939) );
  NOR2_X1 U15015 ( .A1(n11940), .A2(n11939), .ZN(n11967) );
  INV_X1 U15016 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11943) );
  INV_X1 U15017 ( .A(n12008), .ZN(n12032) );
  INV_X1 U15018 ( .A(n19262), .ZN(n11942) );
  OAI22_X1 U15019 ( .A1(n11943), .A2(n12032), .B1(n11942), .B2(n11941), .ZN(
        n11947) );
  INV_X1 U15020 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11945) );
  INV_X1 U15021 ( .A(n19353), .ZN(n11944) );
  INV_X1 U15022 ( .A(n12002), .ZN(n19295) );
  INV_X1 U15023 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12439) );
  OAI22_X1 U15024 ( .A1(n11945), .A2(n11944), .B1(n19295), .B2(n12439), .ZN(
        n11946) );
  NOR2_X1 U15025 ( .A1(n11947), .A2(n11946), .ZN(n11966) );
  INV_X1 U15026 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11949) );
  INV_X1 U15027 ( .A(n12007), .ZN(n11948) );
  INV_X1 U15028 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n19524) );
  OAI22_X1 U15029 ( .A1(n11949), .A2(n11948), .B1(n12001), .B2(n19524), .ZN(
        n11955) );
  INV_X1 U15030 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11953) );
  INV_X1 U15031 ( .A(n19433), .ZN(n11952) );
  INV_X1 U15032 ( .A(n12030), .ZN(n11951) );
  INV_X1 U15033 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11950) );
  OAI22_X1 U15034 ( .A1(n11953), .A2(n11952), .B1(n11951), .B2(n11950), .ZN(
        n11954) );
  NOR2_X1 U15035 ( .A1(n11955), .A2(n11954), .ZN(n11965) );
  INV_X1 U15036 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11958) );
  INV_X1 U15037 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11956) );
  OAI22_X1 U15038 ( .A1(n11958), .A2(n11957), .B1(n19601), .B2(n11956), .ZN(
        n11963) );
  INV_X1 U15039 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11961) );
  INV_X1 U15040 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11959) );
  OAI22_X1 U15041 ( .A1(n11961), .A2(n19494), .B1(n11960), .B2(n11959), .ZN(
        n11962) );
  NOR2_X1 U15042 ( .A1(n11963), .A2(n11962), .ZN(n11964) );
  NAND4_X1 U15043 ( .A1(n11967), .A2(n11966), .A3(n11965), .A4(n11964), .ZN(
        n11970) );
  NOR2_X1 U15044 ( .A1(n12308), .A2(n12310), .ZN(n11968) );
  NAND2_X1 U15045 ( .A1(n19869), .A2(n11968), .ZN(n12314) );
  NAND2_X1 U15046 ( .A1(n12314), .A2(n12313), .ZN(n11969) );
  INV_X1 U15047 ( .A(n11993), .ZN(n11973) );
  OR2_X1 U15048 ( .A1(n11982), .A2(n11971), .ZN(n11972) );
  NAND2_X1 U15049 ( .A1(n11973), .A2(n11972), .ZN(n14849) );
  AND2_X1 U15050 ( .A1(n14108), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11975) );
  NOR2_X1 U15051 ( .A1(n11976), .A2(n11975), .ZN(n12227) );
  INV_X1 U15052 ( .A(n12227), .ZN(n11977) );
  MUX2_X1 U15053 ( .A(n12308), .B(n11977), .S(n12247), .Z(n12207) );
  MUX2_X1 U15054 ( .A(n12207), .B(n19032), .S(n19237), .Z(n19027) );
  NOR2_X1 U15055 ( .A1(n19027), .A2(n15557), .ZN(n13212) );
  AND2_X1 U15056 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(P2_EBX_REG_0__SCAN_IN), 
        .ZN(n11978) );
  NAND2_X1 U15057 ( .A1(n19237), .A2(n11978), .ZN(n11979) );
  NAND2_X1 U15058 ( .A1(n11983), .A2(n11979), .ZN(n14873) );
  NOR2_X1 U15059 ( .A1(n14873), .A2(n15558), .ZN(n11981) );
  INV_X1 U15060 ( .A(n14873), .ZN(n11980) );
  OAI22_X1 U15061 ( .A1(n13212), .A2(n11981), .B1(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n11980), .ZN(n13262) );
  INV_X1 U15062 ( .A(n13262), .ZN(n11987) );
  INV_X1 U15063 ( .A(n11982), .ZN(n11986) );
  NAND2_X1 U15064 ( .A1(n11984), .A2(n11983), .ZN(n11985) );
  NAND2_X1 U15065 ( .A1(n11986), .A2(n11985), .ZN(n14858) );
  XNOR2_X1 U15066 ( .A(n14858), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13261) );
  NAND2_X1 U15067 ( .A1(n11987), .A2(n13261), .ZN(n13289) );
  INV_X1 U15068 ( .A(n14858), .ZN(n11988) );
  NAND2_X1 U15069 ( .A1(n11988), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11989) );
  AND2_X1 U15070 ( .A1(n13289), .A2(n11989), .ZN(n13763) );
  INV_X1 U15071 ( .A(n11991), .ZN(n11992) );
  XNOR2_X1 U15072 ( .A(n11993), .B(n11992), .ZN(n14833) );
  XNOR2_X1 U15073 ( .A(n14833), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19192) );
  INV_X1 U15074 ( .A(n19192), .ZN(n11994) );
  NAND2_X1 U15075 ( .A1(n14833), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11995) );
  INV_X1 U15076 ( .A(n11996), .ZN(n11998) );
  AOI22_X1 U15077 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n11999), .B1(
        n12000), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12006) );
  AOI22_X1 U15078 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19353), .B1(
        n15614), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12005) );
  AOI22_X1 U15079 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19433), .B1(
        n21051), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12004) );
  AOI22_X1 U15080 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n12002), .B1(
        n19262), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12003) );
  INV_X1 U15081 ( .A(n19601), .ZN(n12025) );
  AOI22_X1 U15082 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19497), .B1(
        n12025), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12015) );
  AOI22_X1 U15083 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n12007), .B1(
        n12030), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12014) );
  AOI22_X1 U15084 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n12008), .B1(
        n12009), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U15085 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n12010), .B1(
        n12011), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12012) );
  NAND2_X1 U15086 ( .A1(n12016), .A2(n19869), .ZN(n12017) );
  XNOR2_X1 U15087 ( .A(n12020), .B(n12019), .ZN(n19015) );
  INV_X1 U15088 ( .A(n12047), .ZN(n12046) );
  AOI22_X1 U15089 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19353), .B1(
        n15614), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12029) );
  AOI22_X1 U15090 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12007), .B1(
        n12025), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12028) );
  AOI22_X1 U15091 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n12011), .B1(
        n21051), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12027) );
  AOI22_X1 U15092 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12002), .B1(
        n19262), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12026) );
  NAND4_X1 U15093 ( .A1(n12029), .A2(n12028), .A3(n12027), .A4(n12026), .ZN(
        n12040) );
  AOI22_X1 U15094 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n11999), .B1(
        n12000), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12038) );
  AOI22_X1 U15095 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19433), .B1(
        n19497), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12037) );
  AOI22_X1 U15096 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12030), .B1(
        n12009), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12036) );
  OAI22_X1 U15097 ( .A1(n12033), .A2(n12032), .B1(n12031), .B2(n19249), .ZN(
        n12034) );
  INV_X1 U15098 ( .A(n12034), .ZN(n12035) );
  NAND4_X1 U15099 ( .A1(n12038), .A2(n12037), .A3(n12036), .A4(n12035), .ZN(
        n12039) );
  INV_X1 U15100 ( .A(n12041), .ZN(n12042) );
  NAND2_X1 U15101 ( .A1(n19869), .A2(n12042), .ZN(n12043) );
  NAND2_X1 U15102 ( .A1(n12047), .A2(n12329), .ZN(n12336) );
  OR2_X1 U15103 ( .A1(n12050), .A2(n12049), .ZN(n12051) );
  NAND2_X1 U15104 ( .A1(n12056), .A2(n12051), .ZN(n19000) );
  INV_X1 U15105 ( .A(n12054), .ZN(n15237) );
  NAND2_X1 U15106 ( .A1(n15237), .A2(n20868), .ZN(n12053) );
  NAND2_X1 U15107 ( .A1(n15233), .A2(n12053), .ZN(n12060) );
  AND2_X1 U15108 ( .A1(n12052), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15234) );
  NAND2_X1 U15109 ( .A1(n12053), .A2(n15234), .ZN(n12059) );
  NAND2_X1 U15110 ( .A1(n12054), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15238) );
  XNOR2_X1 U15111 ( .A(n12056), .B(n9913), .ZN(n18990) );
  NAND2_X1 U15112 ( .A1(n18990), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15528) );
  XNOR2_X1 U15113 ( .A(n9802), .B(n10148), .ZN(n14821) );
  INV_X1 U15114 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16216) );
  NOR2_X1 U15115 ( .A1(n12158), .A2(n16216), .ZN(n12057) );
  NAND2_X1 U15116 ( .A1(n14821), .A2(n12057), .ZN(n15241) );
  NAND2_X1 U15117 ( .A1(n14821), .A2(n12762), .ZN(n12061) );
  NAND2_X1 U15118 ( .A1(n12061), .A2(n16216), .ZN(n15242) );
  INV_X1 U15119 ( .A(n18990), .ZN(n12062) );
  NAND2_X1 U15120 ( .A1(n12062), .A2(n15539), .ZN(n15527) );
  AND2_X1 U15121 ( .A1(n15242), .A2(n15527), .ZN(n12063) );
  NAND2_X1 U15122 ( .A1(n19237), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n12064) );
  XNOR2_X1 U15123 ( .A(n12065), .B(n12064), .ZN(n18979) );
  NAND2_X1 U15124 ( .A1(n18979), .A2(n12762), .ZN(n12076) );
  INV_X1 U15125 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12075) );
  AND2_X1 U15126 ( .A1(n12076), .A2(n12075), .ZN(n15508) );
  INV_X1 U15127 ( .A(n15508), .ZN(n12066) );
  NAND2_X1 U15128 ( .A1(n19237), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n12068) );
  MUX2_X1 U15129 ( .A(n12068), .B(P2_EBX_REG_10__SCAN_IN), .S(n12067), .Z(
        n12069) );
  AND2_X1 U15130 ( .A1(n12069), .A2(n12155), .ZN(n14810) );
  NAND2_X1 U15131 ( .A1(n14810), .A2(n12762), .ZN(n12077) );
  NAND2_X1 U15132 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n12070), .ZN(n12071) );
  NOR2_X1 U15133 ( .A1(n12150), .A2(n12071), .ZN(n12072) );
  NOR2_X1 U15134 ( .A1(n12073), .A2(n12072), .ZN(n13120) );
  NAND2_X1 U15135 ( .A1(n13120), .A2(n12762), .ZN(n12074) );
  INV_X1 U15136 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15500) );
  NAND2_X1 U15137 ( .A1(n12074), .A2(n15500), .ZN(n15207) );
  OR2_X1 U15138 ( .A1(n12074), .A2(n15500), .ZN(n15208) );
  NOR2_X1 U15139 ( .A1(n12076), .A2(n12075), .ZN(n15509) );
  NOR2_X1 U15140 ( .A1(n16207), .A2(n12077), .ZN(n15219) );
  NOR2_X1 U15141 ( .A1(n15509), .A2(n15219), .ZN(n15205) );
  AND2_X1 U15142 ( .A1(n15208), .A2(n15205), .ZN(n15121) );
  NAND3_X1 U15143 ( .A1(n19237), .A2(n12078), .A3(P2_EBX_REG_12__SCAN_IN), 
        .ZN(n12079) );
  AND2_X1 U15144 ( .A1(n12085), .A2(n12079), .ZN(n18968) );
  INV_X1 U15145 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15194) );
  NOR2_X1 U15146 ( .A1(n12158), .A2(n15194), .ZN(n12080) );
  INV_X1 U15147 ( .A(n18968), .ZN(n12081) );
  OAI21_X1 U15148 ( .B1(n12081), .B2(n12158), .A(n15194), .ZN(n15196) );
  INV_X1 U15149 ( .A(n15196), .ZN(n12082) );
  INV_X1 U15150 ( .A(n12083), .ZN(n12084) );
  XNOR2_X1 U15151 ( .A(n12085), .B(n12084), .ZN(n18954) );
  NAND2_X1 U15152 ( .A1(n18954), .A2(n12762), .ZN(n12086) );
  NAND2_X1 U15153 ( .A1(n12086), .A2(n15488), .ZN(n15185) );
  NAND2_X1 U15154 ( .A1(n15183), .A2(n15185), .ZN(n15174) );
  NAND2_X1 U15155 ( .A1(n19237), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n12087) );
  NOR2_X1 U15156 ( .A1(n12088), .A2(n12087), .ZN(n12089) );
  NOR2_X1 U15157 ( .A1(n12090), .A2(n12089), .ZN(n14770) );
  INV_X1 U15158 ( .A(n14770), .ZN(n12091) );
  INV_X1 U15159 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15367) );
  OAI21_X1 U15160 ( .B1(n12091), .B2(n12158), .A(n15367), .ZN(n15119) );
  OR2_X1 U15161 ( .A1(n12113), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12115) );
  INV_X1 U15162 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n12092) );
  NOR2_X1 U15163 ( .A1(n12150), .A2(n12092), .ZN(n12093) );
  NAND2_X1 U15164 ( .A1(n12115), .A2(n12093), .ZN(n12094) );
  AND2_X1 U15165 ( .A1(n12094), .A2(n12111), .ZN(n12125) );
  INV_X1 U15166 ( .A(n12125), .ZN(n18905) );
  INV_X1 U15167 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15393) );
  OAI21_X1 U15168 ( .B1(n18905), .B2(n12158), .A(n15393), .ZN(n15389) );
  OR2_X1 U15169 ( .A1(n12104), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n12099) );
  NAND3_X1 U15170 ( .A1(n12104), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n19237), 
        .ZN(n12095) );
  NAND3_X1 U15171 ( .A1(n12099), .A2(n12155), .A3(n12095), .ZN(n18935) );
  OR2_X1 U15172 ( .A1(n18935), .A2(n12158), .ZN(n12096) );
  XNOR2_X1 U15173 ( .A(n12096), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15164) );
  INV_X1 U15174 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n12097) );
  NOR2_X1 U15175 ( .A1(n12150), .A2(n12097), .ZN(n12098) );
  NAND2_X1 U15176 ( .A1(n12099), .A2(n12098), .ZN(n12100) );
  NAND2_X1 U15177 ( .A1(n12100), .A2(n12113), .ZN(n18920) );
  OR2_X1 U15178 ( .A1(n18920), .A2(n12158), .ZN(n12101) );
  NAND2_X1 U15179 ( .A1(n12101), .A2(n21010), .ZN(n15152) );
  NAND2_X1 U15180 ( .A1(n12102), .A2(n12106), .ZN(n12103) );
  NAND3_X1 U15181 ( .A1(n12103), .A2(P2_EBX_REG_15__SCAN_IN), .A3(n19237), 
        .ZN(n12105) );
  NAND2_X1 U15182 ( .A1(n12105), .A2(n12104), .ZN(n13103) );
  INV_X1 U15183 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n20957) );
  NAND2_X1 U15184 ( .A1(n12122), .A2(n20957), .ZN(n15449) );
  AND2_X1 U15185 ( .A1(n15152), .A2(n15449), .ZN(n12109) );
  NOR2_X1 U15186 ( .A1(n12150), .A2(n12106), .ZN(n12107) );
  XNOR2_X1 U15187 ( .A(n12102), .B(n12107), .ZN(n18946) );
  NAND2_X1 U15188 ( .A1(n18946), .A2(n12762), .ZN(n12108) );
  NAND2_X1 U15189 ( .A1(n12108), .A2(n20881), .ZN(n15447) );
  AND4_X1 U15190 ( .A1(n15389), .A2(n15164), .A3(n12109), .A4(n15447), .ZN(
        n12118) );
  NAND2_X1 U15191 ( .A1(n19237), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n12110) );
  XNOR2_X1 U15192 ( .A(n12111), .B(n12110), .ZN(n14784) );
  INV_X1 U15193 ( .A(n12127), .ZN(n12112) );
  INV_X1 U15194 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12349) );
  NAND2_X1 U15195 ( .A1(n12112), .A2(n12349), .ZN(n15130) );
  NAND2_X1 U15196 ( .A1(n12113), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n12114) );
  MUX2_X1 U15197 ( .A(n12114), .B(n12113), .S(n12150), .Z(n12116) );
  NAND2_X1 U15198 ( .A1(n14790), .A2(n12762), .ZN(n12117) );
  NAND2_X1 U15199 ( .A1(n12117), .A2(n15410), .ZN(n15404) );
  NAND4_X1 U15200 ( .A1(n15119), .A2(n12118), .A3(n15130), .A4(n15404), .ZN(
        n12131) );
  NOR2_X1 U15201 ( .A1(n12158), .A2(n15367), .ZN(n12119) );
  NAND2_X1 U15202 ( .A1(n14770), .A2(n12119), .ZN(n15118) );
  OR2_X1 U15203 ( .A1(n12158), .A2(n21010), .ZN(n12120) );
  OR2_X1 U15204 ( .A1(n18920), .A2(n12120), .ZN(n15151) );
  INV_X1 U15205 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15427) );
  OR2_X1 U15206 ( .A1(n12158), .A2(n15427), .ZN(n12121) );
  OR2_X1 U15207 ( .A1(n18935), .A2(n12121), .ZN(n15149) );
  AND2_X1 U15208 ( .A1(n15151), .A2(n15149), .ZN(n15128) );
  OR2_X1 U15209 ( .A1(n12122), .A2(n20957), .ZN(n15450) );
  NOR2_X1 U15210 ( .A1(n12158), .A2(n20881), .ZN(n12123) );
  NAND2_X1 U15211 ( .A1(n18946), .A2(n12123), .ZN(n15175) );
  AND2_X1 U15212 ( .A1(n15450), .A2(n15175), .ZN(n15124) );
  NOR2_X1 U15213 ( .A1(n12158), .A2(n15393), .ZN(n12124) );
  NAND2_X1 U15214 ( .A1(n12125), .A2(n12124), .ZN(n15388) );
  NOR2_X1 U15215 ( .A1(n12158), .A2(n15488), .ZN(n12126) );
  NAND2_X1 U15216 ( .A1(n18954), .A2(n12126), .ZN(n15184) );
  AND4_X1 U15217 ( .A1(n15128), .A2(n15124), .A3(n15388), .A4(n15184), .ZN(
        n12129) );
  NAND2_X1 U15218 ( .A1(n12127), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15131) );
  NOR2_X1 U15219 ( .A1(n12158), .A2(n15410), .ZN(n12128) );
  NAND2_X1 U15220 ( .A1(n14790), .A2(n12128), .ZN(n15403) );
  AND4_X1 U15221 ( .A1(n15118), .A2(n12129), .A3(n15131), .A4(n15403), .ZN(
        n12130) );
  INV_X1 U15222 ( .A(n12132), .ZN(n12133) );
  NAND2_X1 U15223 ( .A1(n12134), .A2(n12133), .ZN(n12135) );
  NAND2_X1 U15224 ( .A1(n12138), .A2(n12135), .ZN(n14750) );
  OR2_X1 U15225 ( .A1(n14750), .A2(n12158), .ZN(n12136) );
  NAND2_X1 U15226 ( .A1(n12136), .A2(n15338), .ZN(n15111) );
  NAND2_X1 U15227 ( .A1(n12138), .A2(n12137), .ZN(n12139) );
  NAND2_X1 U15228 ( .A1(n12152), .A2(n12139), .ZN(n12140) );
  INV_X1 U15229 ( .A(n12140), .ZN(n14741) );
  NAND3_X1 U15230 ( .A1(n14741), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n12762), .ZN(n12145) );
  XNOR2_X1 U15231 ( .A(n12141), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15101) );
  INV_X1 U15232 ( .A(n15101), .ZN(n12142) );
  NAND2_X1 U15233 ( .A1(n12145), .A2(n12142), .ZN(n12144) );
  AND2_X1 U15234 ( .A1(n15111), .A2(n12144), .ZN(n12143) );
  NAND2_X1 U15235 ( .A1(n15098), .A2(n12143), .ZN(n12149) );
  INV_X1 U15236 ( .A(n12144), .ZN(n12147) );
  AND2_X1 U15237 ( .A1(n15110), .A2(n12145), .ZN(n12146) );
  INV_X1 U15238 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n14927) );
  NOR2_X1 U15239 ( .A1(n12150), .A2(n14927), .ZN(n12151) );
  NAND2_X1 U15240 ( .A1(n12152), .A2(n12151), .ZN(n12153) );
  NAND2_X1 U15241 ( .A1(n12153), .A2(n12155), .ZN(n12154) );
  NAND2_X1 U15242 ( .A1(n19237), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n12156) );
  OAI211_X1 U15243 ( .C1(n12157), .C2(n12156), .A(n12160), .B(n12155), .ZN(
        n16118) );
  OR2_X1 U15244 ( .A1(n16118), .A2(n12158), .ZN(n12159) );
  INV_X1 U15245 ( .A(n15069), .ZN(n12163) );
  NAND3_X1 U15246 ( .A1(n12160), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n19237), 
        .ZN(n12161) );
  NAND2_X1 U15247 ( .A1(n12161), .A2(n12768), .ZN(n16106) );
  XNOR2_X1 U15248 ( .A(n12164), .B(n15307), .ZN(n15070) );
  INV_X1 U15249 ( .A(n15070), .ZN(n12162) );
  NAND2_X1 U15250 ( .A1(n12163), .A2(n12162), .ZN(n12169) );
  OR2_X1 U15251 ( .A1(n12164), .A2(n15307), .ZN(n12165) );
  OR3_X1 U15252 ( .A1(n16118), .A2(n12158), .A3(n15316), .ZN(n15080) );
  NAND2_X1 U15253 ( .A1(n12165), .A2(n15080), .ZN(n12755) );
  NOR2_X1 U15254 ( .A1(n12756), .A2(n12755), .ZN(n12173) );
  INV_X1 U15255 ( .A(n12166), .ZN(n12167) );
  NAND2_X1 U15256 ( .A1(n12167), .A2(n10151), .ZN(n12168) );
  NAND2_X1 U15257 ( .A1(n12175), .A2(n12168), .ZN(n16094) );
  NAND2_X1 U15258 ( .A1(n12169), .A2(n12172), .ZN(n12170) );
  NAND3_X1 U15259 ( .A1(n12170), .A2(n10122), .A3(n9807), .ZN(n12171) );
  INV_X1 U15260 ( .A(n12171), .ZN(n15057) );
  OAI21_X1 U15261 ( .B1(n12173), .B2(n12172), .A(n15058), .ZN(n12177) );
  XNOR2_X1 U15262 ( .A(n12175), .B(n12174), .ZN(n16084) );
  NAND2_X1 U15263 ( .A1(n16084), .A2(n12762), .ZN(n12752) );
  XNOR2_X1 U15264 ( .A(n12752), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12176) );
  XNOR2_X1 U15265 ( .A(n12177), .B(n12176), .ZN(n12369) );
  AND2_X1 U15266 ( .A1(n12204), .A2(n12227), .ZN(n12181) );
  OAI21_X1 U15267 ( .B1(n12247), .B2(n12181), .A(n12187), .ZN(n12182) );
  NAND2_X1 U15268 ( .A1(n12180), .A2(n12182), .ZN(n12186) );
  INV_X1 U15269 ( .A(n12183), .ZN(n12184) );
  OAI211_X1 U15270 ( .C1(n9743), .C2(n12227), .A(n10690), .B(n12184), .ZN(
        n12185) );
  NAND2_X1 U15271 ( .A1(n12186), .A2(n12185), .ZN(n12190) );
  NAND2_X1 U15272 ( .A1(n16269), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19121) );
  NAND2_X1 U15273 ( .A1(n19121), .A2(n9743), .ZN(n12188) );
  INV_X1 U15274 ( .A(n12187), .ZN(n12228) );
  MUX2_X1 U15275 ( .A(n12188), .B(n12247), .S(n12228), .Z(n12189) );
  NAND2_X1 U15276 ( .A1(n12190), .A2(n12189), .ZN(n12192) );
  INV_X1 U15277 ( .A(n12230), .ZN(n12191) );
  NAND2_X1 U15278 ( .A1(n12192), .A2(n12191), .ZN(n12193) );
  NAND2_X1 U15279 ( .A1(n12195), .A2(n12197), .ZN(n12196) );
  MUX2_X1 U15280 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n12196), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n12202) );
  INV_X1 U15281 ( .A(n12197), .ZN(n12208) );
  INV_X1 U15282 ( .A(n19121), .ZN(n12198) );
  NAND2_X1 U15283 ( .A1(n12208), .A2(n12198), .ZN(n12199) );
  NAND2_X1 U15284 ( .A1(n16276), .A2(n9743), .ZN(n19118) );
  INV_X1 U15285 ( .A(n12200), .ZN(n16263) );
  NAND2_X1 U15286 ( .A1(n12201), .A2(n16263), .ZN(n12245) );
  AOI21_X1 U15287 ( .B1(n12202), .B2(n10690), .A(n10742), .ZN(n12203) );
  NAND2_X1 U15288 ( .A1(n19118), .A2(n12203), .ZN(n12244) );
  INV_X1 U15289 ( .A(n12204), .ZN(n12206) );
  OAI21_X1 U15290 ( .B1(n12207), .B2(n12206), .A(n12205), .ZN(n12210) );
  AOI21_X1 U15291 ( .B1(n12210), .B2(n12209), .A(n12208), .ZN(n19855) );
  NAND2_X1 U15292 ( .A1(n19869), .A2(n16269), .ZN(n12212) );
  NOR2_X1 U15293 ( .A1(n12248), .A2(n12212), .ZN(n12351) );
  NAND2_X1 U15294 ( .A1(n19855), .A2(n12351), .ZN(n12358) );
  MUX2_X1 U15295 ( .A(n12211), .B(n19223), .S(n19869), .Z(n12240) );
  NAND2_X1 U15296 ( .A1(n16273), .A2(n19867), .ZN(n12239) );
  OAI21_X1 U15297 ( .B1(n10727), .B2(n10737), .A(n12707), .ZN(n12214) );
  INV_X1 U15298 ( .A(n12212), .ZN(n12213) );
  NAND2_X1 U15299 ( .A1(n12214), .A2(n12213), .ZN(n12252) );
  NAND2_X1 U15300 ( .A1(n19869), .A2(n12215), .ZN(n12265) );
  NAND2_X1 U15301 ( .A1(n12265), .A2(n10690), .ZN(n12217) );
  NAND2_X1 U15302 ( .A1(n12217), .A2(n12216), .ZN(n12218) );
  NAND2_X1 U15303 ( .A1(n12218), .A2(n19223), .ZN(n12219) );
  AND3_X1 U15304 ( .A1(n12220), .A2(n12252), .A3(n12219), .ZN(n12225) );
  NAND2_X1 U15305 ( .A1(n12222), .A2(n19223), .ZN(n12223) );
  NAND2_X1 U15306 ( .A1(n12221), .A2(n12223), .ZN(n12224) );
  NAND3_X1 U15307 ( .A1(n10733), .A2(n16273), .A3(n16263), .ZN(n12226) );
  AND2_X1 U15308 ( .A1(n12267), .A2(n12226), .ZN(n14091) );
  NAND2_X1 U15309 ( .A1(n12228), .A2(n12227), .ZN(n12229) );
  NOR2_X1 U15310 ( .A1(n12230), .A2(n12229), .ZN(n12231) );
  OAI21_X1 U15311 ( .B1(n12232), .B2(n12231), .A(n16287), .ZN(n12237) );
  NAND2_X1 U15312 ( .A1(n16280), .A2(n12233), .ZN(n16259) );
  INV_X1 U15313 ( .A(n16259), .ZN(n12234) );
  NAND2_X1 U15314 ( .A1(n12481), .A2(n12234), .ZN(n12236) );
  INV_X1 U15315 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n18883) );
  AND2_X1 U15316 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n18883), .ZN(n12235) );
  NAND2_X1 U15317 ( .A1(n12236), .A2(n12235), .ZN(n19842) );
  INV_X1 U15318 ( .A(n12248), .ZN(n16270) );
  NAND3_X1 U15319 ( .A1(n19853), .A2(n16270), .A3(n9743), .ZN(n12238) );
  OAI211_X1 U15320 ( .C1(n12240), .C2(n12239), .A(n14091), .B(n12238), .ZN(
        n12241) );
  INV_X1 U15321 ( .A(n12241), .ZN(n12242) );
  AND2_X1 U15322 ( .A1(n12358), .A2(n12242), .ZN(n12243) );
  OAI211_X1 U15323 ( .C1(n19118), .C2(n12245), .A(n12244), .B(n12243), .ZN(
        n12246) );
  NOR2_X1 U15324 ( .A1(n12248), .A2(n12247), .ZN(n12356) );
  INV_X1 U15325 ( .A(n12356), .ZN(n19852) );
  AND2_X1 U15326 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15499) );
  AND3_X1 U15327 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12249) );
  AND2_X1 U15328 ( .A1(n15499), .A2(n12249), .ZN(n15432) );
  AND2_X1 U15329 ( .A1(n15432), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15420) );
  AND3_X1 U15330 ( .A1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12250) );
  NAND2_X1 U15331 ( .A1(n15420), .A2(n12250), .ZN(n15407) );
  NOR2_X1 U15332 ( .A1(n15407), .A2(n15410), .ZN(n12348) );
  NOR2_X1 U15333 ( .A1(n15558), .A2(n15557), .ZN(n15555) );
  NAND2_X1 U15334 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n15555), .ZN(
        n13292) );
  NAND2_X1 U15335 ( .A1(n12251), .A2(n9743), .ZN(n14099) );
  NAND2_X1 U15336 ( .A1(n14099), .A2(n12252), .ZN(n12253) );
  NAND2_X1 U15337 ( .A1(n12253), .A2(n10729), .ZN(n12262) );
  OAI22_X1 U15338 ( .A1(n12180), .A2(n10742), .B1(n10690), .B2(n19223), .ZN(
        n12254) );
  INV_X1 U15339 ( .A(n12254), .ZN(n12256) );
  AND2_X1 U15340 ( .A1(n12256), .A2(n12255), .ZN(n12261) );
  MUX2_X1 U15341 ( .A(n10723), .B(n12257), .S(n10759), .Z(n12259) );
  INV_X1 U15342 ( .A(n12180), .ZN(n19873) );
  OAI21_X1 U15343 ( .B1(n12259), .B2(n19873), .A(n12258), .ZN(n12260) );
  NAND3_X1 U15344 ( .A1(n12262), .A2(n12261), .A3(n12260), .ZN(n16241) );
  NOR2_X1 U15345 ( .A1(n16241), .A2(n12263), .ZN(n12264) );
  INV_X1 U15346 ( .A(n12265), .ZN(n12266) );
  NAND2_X1 U15347 ( .A1(n12267), .A2(n12266), .ZN(n15582) );
  NOR2_X1 U15348 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n15555), .ZN(
        n13294) );
  OAI22_X1 U15349 ( .A1(n13292), .A2(n15425), .B1(n12274), .B2(n13294), .ZN(
        n13772) );
  NAND2_X1 U15350 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13772), .ZN(
        n19222) );
  NOR2_X1 U15351 ( .A1(n19209), .A2(n13970), .ZN(n15549) );
  NAND2_X1 U15352 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15549), .ZN(
        n12271) );
  NOR2_X1 U15353 ( .A1(n19222), .A2(n12271), .ZN(n16215) );
  NOR2_X1 U15354 ( .A1(n15539), .A2(n16216), .ZN(n16219) );
  NAND2_X1 U15355 ( .A1(n16215), .A2(n16219), .ZN(n15469) );
  NAND2_X1 U15356 ( .A1(n12348), .A2(n15498), .ZN(n15394) );
  AND2_X1 U15357 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12283) );
  INV_X1 U15358 ( .A(n12283), .ZN(n12268) );
  NAND2_X1 U15359 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15328) );
  INV_X1 U15360 ( .A(n15328), .ZN(n15337) );
  NAND2_X1 U15361 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15337), .ZN(
        n12269) );
  NOR2_X1 U15362 ( .A1(n15349), .A2(n12269), .ZN(n15313) );
  NAND2_X1 U15363 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12287) );
  INV_X1 U15364 ( .A(n12287), .ZN(n12270) );
  NAND2_X1 U15365 ( .A1(n15313), .A2(n12270), .ZN(n15292) );
  INV_X1 U15366 ( .A(n15292), .ZN(n15279) );
  AND2_X1 U15367 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15278) );
  INV_X1 U15368 ( .A(n12271), .ZN(n12272) );
  NAND2_X1 U15369 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n12272), .ZN(
        n12273) );
  NAND2_X1 U15370 ( .A1(n15426), .A2(n12273), .ZN(n12278) );
  INV_X1 U15371 ( .A(n15425), .ZN(n12275) );
  INV_X1 U15372 ( .A(n12274), .ZN(n15419) );
  AOI22_X1 U15373 ( .A1(n12275), .A2(n13292), .B1(n15419), .B2(n13294), .ZN(
        n12276) );
  INV_X2 U15374 ( .A(n19206), .ZN(n19012) );
  NAND2_X1 U15375 ( .A1(n12352), .A2(n19012), .ZN(n13273) );
  NAND2_X1 U15376 ( .A1(n12276), .A2(n13273), .ZN(n13971) );
  INV_X1 U15377 ( .A(n13971), .ZN(n12277) );
  INV_X1 U15378 ( .A(n16219), .ZN(n12279) );
  NAND2_X1 U15379 ( .A1(n15426), .A2(n12279), .ZN(n12280) );
  AND2_X1 U15380 ( .A1(n16217), .A2(n12280), .ZN(n15468) );
  NAND2_X1 U15381 ( .A1(n15426), .A2(n15407), .ZN(n12281) );
  AND2_X1 U15382 ( .A1(n15468), .A2(n12281), .ZN(n15409) );
  NAND2_X1 U15383 ( .A1(n15426), .A2(n15410), .ZN(n12282) );
  NAND2_X1 U15384 ( .A1(n15409), .A2(n12282), .ZN(n15396) );
  NOR2_X1 U15385 ( .A1(n15556), .A2(n12283), .ZN(n12284) );
  NOR2_X1 U15386 ( .A1(n15396), .A2(n12284), .ZN(n15368) );
  NAND2_X1 U15387 ( .A1(n15426), .A2(n15367), .ZN(n12285) );
  NAND2_X1 U15388 ( .A1(n15368), .A2(n12285), .ZN(n15353) );
  NOR2_X1 U15389 ( .A1(n15556), .A2(n15337), .ZN(n12286) );
  INV_X1 U15390 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15092) );
  OR3_X1 U15391 ( .A1(n15353), .A2(n12286), .A3(n15092), .ZN(n15329) );
  NAND2_X1 U15392 ( .A1(n15368), .A2(n15556), .ZN(n12288) );
  NAND2_X1 U15393 ( .A1(n15329), .A2(n12288), .ZN(n15317) );
  NAND2_X1 U15394 ( .A1(n12288), .A2(n12287), .ZN(n12289) );
  NAND2_X1 U15395 ( .A1(n15317), .A2(n12289), .ZN(n15294) );
  AOI21_X1 U15396 ( .B1(n15279), .B2(n10123), .A(n15294), .ZN(n15276) );
  INV_X1 U15397 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12298) );
  INV_X1 U15398 ( .A(n12290), .ZN(n12291) );
  NAND2_X1 U15399 ( .A1(n12291), .A2(n10769), .ZN(n15581) );
  OAI21_X1 U15400 ( .B1(n19869), .B2(n10722), .A(n15581), .ZN(n12292) );
  INV_X1 U15401 ( .A(n12292), .ZN(n12293) );
  AND2_X1 U15402 ( .A1(n9813), .A2(n12294), .ZN(n12295) );
  NOR2_X1 U15403 ( .A1(n9769), .A2(n12295), .ZN(n16085) );
  NOR2_X1 U15404 ( .A1(n19012), .A2(n19793), .ZN(n12362) );
  INV_X1 U15405 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15056) );
  NOR3_X1 U15406 ( .A1(n15292), .A2(n15278), .A3(n15056), .ZN(n12296) );
  AOI211_X1 U15407 ( .C1(n19208), .C2(n16085), .A(n12362), .B(n12296), .ZN(
        n12297) );
  OAI21_X1 U15408 ( .B1(n15276), .B2(n12298), .A(n12297), .ZN(n12305) );
  AND2_X1 U15409 ( .A1(n14900), .A2(n12299), .ZN(n12301) );
  OR2_X1 U15410 ( .A1(n12301), .A2(n12300), .ZN(n14890) );
  INV_X1 U15411 ( .A(n12302), .ZN(n12303) );
  INV_X1 U15412 ( .A(n12308), .ZN(n13187) );
  NOR2_X1 U15413 ( .A1(n15557), .A2(n13187), .ZN(n13186) );
  INV_X1 U15414 ( .A(n12310), .ZN(n12309) );
  NAND2_X1 U15415 ( .A1(n13186), .A2(n12309), .ZN(n12312) );
  NOR2_X1 U15416 ( .A1(n13187), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12311) );
  XOR2_X1 U15417 ( .A(n12311), .B(n12310), .Z(n13214) );
  NAND2_X1 U15418 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13214), .ZN(
        n13213) );
  NAND2_X1 U15419 ( .A1(n12312), .A2(n13213), .ZN(n12315) );
  XOR2_X1 U15420 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n12315), .Z(
        n13267) );
  XNOR2_X1 U15421 ( .A(n12314), .B(n12313), .ZN(n13266) );
  NAND2_X1 U15422 ( .A1(n13267), .A2(n13266), .ZN(n12317) );
  NAND2_X1 U15423 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12315), .ZN(
        n12316) );
  NAND2_X1 U15424 ( .A1(n12317), .A2(n12316), .ZN(n12318) );
  XNOR2_X1 U15425 ( .A(n12318), .B(n13972), .ZN(n13766) );
  NAND2_X1 U15426 ( .A1(n13765), .A2(n13766), .ZN(n12320) );
  NAND2_X1 U15427 ( .A1(n12318), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12319) );
  INV_X1 U15428 ( .A(n12321), .ZN(n12323) );
  NAND2_X1 U15429 ( .A1(n12323), .A2(n12322), .ZN(n12324) );
  INV_X1 U15430 ( .A(n12325), .ZN(n12326) );
  INV_X1 U15431 ( .A(n12327), .ZN(n12333) );
  NAND2_X1 U15432 ( .A1(n12325), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12331) );
  NAND2_X1 U15433 ( .A1(n12333), .A2(n12331), .ZN(n12328) );
  INV_X1 U15434 ( .A(n12331), .ZN(n13965) );
  NAND2_X1 U15435 ( .A1(n13965), .A2(n12045), .ZN(n12330) );
  NAND2_X1 U15436 ( .A1(n12332), .A2(n12331), .ZN(n12334) );
  NAND2_X1 U15437 ( .A1(n12334), .A2(n12333), .ZN(n12335) );
  INV_X1 U15438 ( .A(n12343), .ZN(n12338) );
  NAND2_X1 U15439 ( .A1(n12336), .A2(n12158), .ZN(n12337) );
  NAND2_X1 U15440 ( .A1(n12345), .A2(n12337), .ZN(n12339) );
  INV_X1 U15441 ( .A(n12339), .ZN(n12342) );
  NAND2_X1 U15442 ( .A1(n12338), .A2(n12342), .ZN(n12341) );
  NAND2_X1 U15443 ( .A1(n12343), .A2(n12339), .ZN(n12340) );
  NAND2_X1 U15444 ( .A1(n15525), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15526) );
  NAND2_X1 U15445 ( .A1(n12343), .A2(n12342), .ZN(n12344) );
  NAND2_X1 U15446 ( .A1(n15229), .A2(n15231), .ZN(n15230) );
  INV_X1 U15447 ( .A(n12345), .ZN(n12346) );
  NOR2_X2 U15448 ( .A1(n15137), .A2(n15367), .ZN(n15108) );
  AND2_X1 U15449 ( .A1(n15278), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12350) );
  OAI21_X1 U15450 ( .B1(n15301), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12728), .ZN(n12365) );
  INV_X1 U15451 ( .A(n12351), .ZN(n19854) );
  NOR2_X1 U15452 ( .A1(n12365), .A2(n19215), .ZN(n12353) );
  INV_X1 U15453 ( .A(n12353), .ZN(n12354) );
  OAI211_X1 U15454 ( .C1(n12369), .C2(n16227), .A(n12355), .B(n12354), .ZN(
        P2_U3018) );
  NAND2_X1 U15455 ( .A1(n19853), .A2(n12356), .ZN(n12357) );
  NAND2_X1 U15456 ( .A1(n12358), .A2(n12357), .ZN(n12359) );
  NAND2_X1 U15457 ( .A1(n12359), .A2(n13249), .ZN(n18882) );
  NAND2_X1 U15458 ( .A1(n16287), .A2(n19385), .ZN(n19816) );
  NAND2_X1 U15459 ( .A1(n19636), .A2(n19816), .ZN(n19841) );
  NAND2_X1 U15460 ( .A1(n19841), .A2(n18874), .ZN(n12360) );
  AND2_X1 U15461 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19831) );
  NAND2_X1 U15462 ( .A1(n18874), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12396) );
  NAND2_X1 U15463 ( .A1(n19868), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n12361) );
  NAND2_X1 U15464 ( .A1(n12396), .A2(n12361), .ZN(n13191) );
  AOI21_X1 U15465 ( .B1(n19190), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n12362), .ZN(n12363) );
  OAI21_X1 U15466 ( .B1(n16089), .B2(n19205), .A(n12363), .ZN(n12364) );
  NOR2_X1 U15467 ( .A1(n12365), .A2(n19197), .ZN(n12366) );
  INV_X1 U15468 ( .A(n12366), .ZN(n12367) );
  OAI211_X1 U15469 ( .C1(n12369), .C2(n19198), .A(n12368), .B(n12367), .ZN(
        P2_U2986) );
  INV_X1 U15470 ( .A(n12396), .ZN(n12379) );
  NAND2_X1 U15471 ( .A1(n10721), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12370) );
  NAND2_X1 U15472 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19545) );
  NAND2_X1 U15473 ( .A1(n19545), .A2(n12371), .ZN(n12372) );
  NOR2_X1 U15474 ( .A1(n12371), .A2(n10670), .ZN(n19671) );
  NAND2_X1 U15475 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19671), .ZN(
        n12390) );
  NAND2_X1 U15476 ( .A1(n12372), .A2(n12390), .ZN(n15623) );
  NOR2_X1 U15477 ( .A1(n15623), .A2(n19636), .ZN(n12373) );
  AOI21_X1 U15478 ( .B1(n12394), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12373), .ZN(n12374) );
  NAND2_X1 U15479 ( .A1(n12644), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n12385) );
  AOI22_X1 U15480 ( .A1(n12394), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19820), .B2(n12376), .ZN(n12377) );
  AND2_X1 U15481 ( .A1(n12644), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12383) );
  XNOR2_X1 U15482 ( .A(n14104), .B(n12383), .ZN(n13254) );
  NAND2_X1 U15483 ( .A1(n15568), .A2(n12379), .ZN(n12382) );
  NAND2_X1 U15484 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n10670), .ZN(
        n19261) );
  NAND2_X1 U15485 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n12376), .ZN(
        n19290) );
  NAND2_X1 U15486 ( .A1(n19261), .A2(n19290), .ZN(n15622) );
  INV_X1 U15487 ( .A(n15622), .ZN(n12380) );
  NOR2_X1 U15488 ( .A1(n19636), .A2(n12380), .ZN(n19292) );
  AOI21_X1 U15489 ( .B1(n12394), .B2(n16229), .A(n19292), .ZN(n12381) );
  NAND2_X1 U15490 ( .A1(n12382), .A2(n12381), .ZN(n13253) );
  NAND2_X1 U15491 ( .A1(n13301), .A2(n13302), .ZN(n12389) );
  INV_X1 U15492 ( .A(n12385), .ZN(n12386) );
  NAND2_X1 U15493 ( .A1(n12387), .A2(n12386), .ZN(n12388) );
  INV_X1 U15494 ( .A(n12390), .ZN(n12391) );
  OAI21_X1 U15495 ( .B1(n12391), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n19820), .ZN(n12392) );
  NOR2_X1 U15496 ( .A1(n12392), .A2(n19724), .ZN(n12393) );
  AOI21_X1 U15497 ( .B1(n12394), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n12393), .ZN(n12395) );
  NAND2_X1 U15498 ( .A1(n12644), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12398) );
  XNOR2_X1 U15499 ( .A(n12397), .B(n12398), .ZN(n13476) );
  NAND2_X1 U15500 ( .A1(n13477), .A2(n13476), .ZN(n12401) );
  INV_X1 U15501 ( .A(n12398), .ZN(n12399) );
  AOI22_X1 U15502 ( .A1(n12397), .A2(n12399), .B1(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n10721), .ZN(n12400) );
  AND2_X1 U15503 ( .A1(n12644), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13416) );
  INV_X1 U15504 ( .A(n12402), .ZN(n13632) );
  NAND2_X1 U15505 ( .A1(n13728), .A2(n13791), .ZN(n13854) );
  NAND2_X1 U15506 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n12408) );
  AOI22_X1 U15507 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12407) );
  NAND2_X1 U15508 ( .A1(n12518), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n12406) );
  NAND2_X1 U15509 ( .A1(n12465), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12405) );
  AND4_X1 U15510 ( .A1(n12408), .A2(n12407), .A3(n12406), .A4(n12405), .ZN(
        n12418) );
  NAND2_X1 U15511 ( .A1(n10366), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12414) );
  NAND2_X1 U15512 ( .A1(n12523), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12413) );
  AOI22_X1 U15513 ( .A1(n10292), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12412) );
  INV_X1 U15514 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n20924) );
  NAND2_X1 U15515 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n12525), .ZN(
        n12409) );
  OAI21_X1 U15516 ( .B1(n12528), .B2(n20924), .A(n12409), .ZN(n12410) );
  AOI21_X1 U15517 ( .B1(n10322), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n12410), .ZN(n12411) );
  AND4_X1 U15518 ( .A1(n12414), .A2(n12413), .A3(n12412), .A4(n12411), .ZN(
        n12417) );
  AOI22_X1 U15519 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10274), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12416) );
  AOI22_X1 U15520 ( .A1(n10352), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10287), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12415) );
  NAND2_X1 U15521 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n12422) );
  AOI22_X1 U15522 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12421) );
  NAND2_X1 U15523 ( .A1(n12518), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n12420) );
  NAND2_X1 U15524 ( .A1(n12465), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12419) );
  AND4_X1 U15525 ( .A1(n12422), .A2(n12421), .A3(n12420), .A4(n12419), .ZN(
        n12433) );
  NAND2_X1 U15526 ( .A1(n10366), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12429) );
  NAND2_X1 U15527 ( .A1(n12523), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n12428) );
  AOI22_X1 U15528 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n10292), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12427) );
  INV_X1 U15529 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12424) );
  NAND2_X1 U15530 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n12525), .ZN(
        n12423) );
  OAI21_X1 U15531 ( .B1(n12528), .B2(n12424), .A(n12423), .ZN(n12425) );
  AOI21_X1 U15532 ( .B1(n10322), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n12425), .ZN(n12426) );
  AND4_X1 U15533 ( .A1(n12429), .A2(n12428), .A3(n12427), .A4(n12426), .ZN(
        n12432) );
  AOI22_X1 U15534 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n10274), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12431) );
  AOI22_X1 U15535 ( .A1(n10352), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10287), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12430) );
  NAND4_X1 U15536 ( .A1(n12433), .A2(n12432), .A3(n12431), .A4(n12430), .ZN(
        n14958) );
  NAND2_X1 U15537 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n12437) );
  AOI22_X1 U15538 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12436) );
  NAND2_X1 U15539 ( .A1(n12518), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n12435) );
  NAND2_X1 U15540 ( .A1(n12465), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12434) );
  AND4_X1 U15541 ( .A1(n12437), .A2(n12436), .A3(n12435), .A4(n12434), .ZN(
        n12448) );
  NAND2_X1 U15542 ( .A1(n10366), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12444) );
  NAND2_X1 U15543 ( .A1(n12523), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n12443) );
  AOI22_X1 U15544 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n10292), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12442) );
  NAND2_X1 U15545 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n12525), .ZN(
        n12438) );
  OAI21_X1 U15546 ( .B1(n12528), .B2(n12439), .A(n12438), .ZN(n12440) );
  AOI21_X1 U15547 ( .B1(n10322), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n12440), .ZN(n12441) );
  AND4_X1 U15548 ( .A1(n12444), .A2(n12443), .A3(n12442), .A4(n12441), .ZN(
        n12447) );
  AOI22_X1 U15549 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10274), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12446) );
  AOI22_X1 U15550 ( .A1(n10352), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n10287), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12445) );
  NAND4_X1 U15551 ( .A1(n12448), .A2(n12447), .A3(n12446), .A4(n12445), .ZN(
        n14001) );
  NAND2_X1 U15552 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n12452) );
  AOI22_X1 U15553 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12451) );
  NAND2_X1 U15554 ( .A1(n12518), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n12450) );
  NAND2_X1 U15555 ( .A1(n12465), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12449) );
  AND4_X1 U15556 ( .A1(n12452), .A2(n12451), .A3(n12450), .A4(n12449), .ZN(
        n12463) );
  NAND2_X1 U15557 ( .A1(n10366), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12459) );
  NAND2_X1 U15558 ( .A1(n12523), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n12458) );
  AOI22_X1 U15559 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n10292), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12457) );
  INV_X1 U15560 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12454) );
  NAND2_X1 U15561 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n12525), .ZN(
        n12453) );
  OAI21_X1 U15562 ( .B1(n12528), .B2(n12454), .A(n12453), .ZN(n12455) );
  AOI21_X1 U15563 ( .B1(n10322), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n12455), .ZN(n12456) );
  AND4_X1 U15564 ( .A1(n12459), .A2(n12458), .A3(n12457), .A4(n12456), .ZN(
        n12462) );
  AOI22_X1 U15565 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n10274), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12461) );
  AOI22_X1 U15566 ( .A1(n10352), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10287), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12460) );
  NAND4_X1 U15567 ( .A1(n12463), .A2(n12462), .A3(n12461), .A4(n12460), .ZN(
        n14953) );
  NAND2_X1 U15568 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n12469) );
  AOI22_X1 U15569 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12468) );
  NAND2_X1 U15570 ( .A1(n12518), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n12467) );
  NAND2_X1 U15571 ( .A1(n12465), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12466) );
  AND4_X1 U15572 ( .A1(n12469), .A2(n12468), .A3(n12467), .A4(n12466), .ZN(
        n12479) );
  NAND2_X1 U15573 ( .A1(n10366), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12475) );
  NAND2_X1 U15574 ( .A1(n12523), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n12474) );
  AOI22_X1 U15575 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10292), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12473) );
  INV_X1 U15576 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n20927) );
  NAND2_X1 U15577 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n12525), .ZN(
        n12470) );
  OAI21_X1 U15578 ( .B1(n12528), .B2(n20927), .A(n12470), .ZN(n12471) );
  AOI21_X1 U15579 ( .B1(n10322), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n12471), .ZN(n12472) );
  AND4_X1 U15580 ( .A1(n12475), .A2(n12474), .A3(n12473), .A4(n12472), .ZN(
        n12478) );
  AOI22_X1 U15581 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n10274), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12477) );
  AOI22_X1 U15582 ( .A1(n10352), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10287), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12476) );
  NAND4_X1 U15583 ( .A1(n12479), .A2(n12478), .A3(n12477), .A4(n12476), .ZN(
        n14948) );
  INV_X1 U15584 ( .A(n14948), .ZN(n12480) );
  NOR2_X1 U15585 ( .A1(n12481), .A2(n19249), .ZN(n12486) );
  INV_X1 U15586 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12483) );
  OAI22_X1 U15587 ( .A1(n12484), .A2(n12483), .B1(n12482), .B2(n10406), .ZN(
        n12485) );
  AOI211_X1 U15588 ( .C1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .C2(n10274), .A(
        n12486), .B(n12485), .ZN(n12493) );
  INV_X1 U15589 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12488) );
  NAND2_X1 U15590 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n12525), .ZN(
        n12487) );
  OAI21_X1 U15591 ( .B1(n12528), .B2(n12488), .A(n12487), .ZN(n12489) );
  AOI21_X1 U15592 ( .B1(n10322), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A(
        n12489), .ZN(n12492) );
  AOI22_X1 U15593 ( .A1(n10292), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12491) );
  AOI22_X1 U15594 ( .A1(n10366), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12523), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12490) );
  NAND4_X1 U15595 ( .A1(n12493), .A2(n12492), .A3(n12491), .A4(n12490), .ZN(
        n12499) );
  INV_X1 U15596 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12496) );
  AOI22_X1 U15597 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12518), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12495) );
  AOI22_X1 U15598 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12494) );
  OAI211_X1 U15599 ( .C1(n12497), .C2(n12496), .A(n12495), .B(n12494), .ZN(
        n12498) );
  NOR2_X1 U15600 ( .A1(n12499), .A2(n12498), .ZN(n14935) );
  INV_X1 U15601 ( .A(n14935), .ZN(n12515) );
  NAND2_X1 U15602 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n12503) );
  AOI22_X1 U15603 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12502) );
  NAND2_X1 U15604 ( .A1(n12518), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n12501) );
  NAND2_X1 U15605 ( .A1(n12465), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12500) );
  AND4_X1 U15606 ( .A1(n12503), .A2(n12502), .A3(n12501), .A4(n12500), .ZN(
        n12514) );
  NAND2_X1 U15607 ( .A1(n10366), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12510) );
  NAND2_X1 U15608 ( .A1(n12523), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n12509) );
  AOI22_X1 U15609 ( .A1(n10292), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12508) );
  INV_X1 U15610 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12505) );
  NAND2_X1 U15611 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n12525), .ZN(
        n12504) );
  OAI21_X1 U15612 ( .B1(n12528), .B2(n12505), .A(n12504), .ZN(n12506) );
  AOI21_X1 U15613 ( .B1(n10322), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n12506), .ZN(n12507) );
  AND4_X1 U15614 ( .A1(n12510), .A2(n12509), .A3(n12508), .A4(n12507), .ZN(
        n12513) );
  AOI22_X1 U15615 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n10274), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12512) );
  AOI22_X1 U15616 ( .A1(n10352), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10287), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12511) );
  NAND4_X1 U15617 ( .A1(n12514), .A2(n12513), .A3(n12512), .A4(n12511), .ZN(
        n14938) );
  AND2_X1 U15618 ( .A1(n12515), .A2(n14938), .ZN(n12516) );
  NAND2_X1 U15619 ( .A1(n12517), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n12522) );
  AOI22_X1 U15620 ( .A1(n10367), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10442), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12521) );
  NAND2_X1 U15621 ( .A1(n12518), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n12520) );
  NAND2_X1 U15622 ( .A1(n12465), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12519) );
  AND4_X1 U15623 ( .A1(n12522), .A2(n12521), .A3(n12520), .A4(n12519), .ZN(
        n12538) );
  NAND2_X1 U15624 ( .A1(n10366), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n12533) );
  NAND2_X1 U15625 ( .A1(n12523), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n12532) );
  AOI22_X1 U15626 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n10292), .B1(
        n12524), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12531) );
  INV_X1 U15627 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12527) );
  NAND2_X1 U15628 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n12525), .ZN(
        n12526) );
  OAI21_X1 U15629 ( .B1(n12528), .B2(n12527), .A(n12526), .ZN(n12529) );
  AOI21_X1 U15630 ( .B1(n10322), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n12529), .ZN(n12530) );
  AND4_X1 U15631 ( .A1(n12533), .A2(n12532), .A3(n12531), .A4(n12530), .ZN(
        n12537) );
  AOI22_X1 U15632 ( .A1(n12534), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n10274), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12536) );
  AOI22_X1 U15633 ( .A1(n10352), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10287), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12535) );
  NAND4_X1 U15634 ( .A1(n12538), .A2(n12537), .A3(n12536), .A4(n12535), .ZN(
        n12559) );
  AOI22_X1 U15635 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10660), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12549) );
  AOI22_X1 U15636 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12686), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12548) );
  AOI22_X1 U15637 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12689), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12547) );
  INV_X1 U15638 ( .A(n12541), .ZN(n15583) );
  NAND2_X1 U15639 ( .A1(n15583), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n12545) );
  NAND2_X1 U15640 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n12544) );
  AND2_X1 U15641 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12543) );
  OR2_X1 U15642 ( .A1(n12543), .A2(n12542), .ZN(n12693) );
  AND3_X1 U15643 ( .A1(n12545), .A2(n12544), .A3(n12693), .ZN(n12546) );
  NAND4_X1 U15644 ( .A1(n12549), .A2(n12548), .A3(n12547), .A4(n12546), .ZN(
        n12558) );
  AOI22_X1 U15645 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10660), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12556) );
  AOI22_X1 U15646 ( .A1(n9745), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12686), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12555) );
  AOI22_X1 U15647 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12689), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12554) );
  INV_X1 U15648 ( .A(n12693), .ZN(n12657) );
  NAND2_X1 U15649 ( .A1(n15583), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n12552) );
  NAND2_X1 U15650 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n12551) );
  AND3_X1 U15651 ( .A1(n12657), .A2(n12552), .A3(n12551), .ZN(n12553) );
  NAND4_X1 U15652 ( .A1(n12556), .A2(n12555), .A3(n12554), .A4(n12553), .ZN(
        n12557) );
  AND2_X1 U15653 ( .A1(n12558), .A2(n12557), .ZN(n12564) );
  NAND2_X1 U15654 ( .A1(n12582), .A2(n9743), .ZN(n12563) );
  INV_X1 U15655 ( .A(n12559), .ZN(n12561) );
  NAND2_X1 U15656 ( .A1(n9743), .A2(n12564), .ZN(n12560) );
  NAND2_X1 U15657 ( .A1(n12561), .A2(n12560), .ZN(n12562) );
  NAND2_X1 U15658 ( .A1(n12563), .A2(n12562), .ZN(n12586) );
  INV_X1 U15659 ( .A(n12564), .ZN(n12565) );
  NOR2_X1 U15660 ( .A1(n9743), .A2(n12565), .ZN(n14930) );
  INV_X1 U15661 ( .A(n14934), .ZN(n12566) );
  AOI22_X1 U15662 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n10661), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12572) );
  AOI22_X1 U15663 ( .A1(n10660), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9744), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12571) );
  AOI22_X1 U15664 ( .A1(n12686), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n15583), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12570) );
  NAND2_X1 U15665 ( .A1(n12689), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12568) );
  NAND2_X1 U15666 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n12567) );
  AND3_X1 U15667 ( .A1(n12657), .A2(n12568), .A3(n12567), .ZN(n12569) );
  NAND4_X1 U15668 ( .A1(n12572), .A2(n12571), .A3(n12570), .A4(n12569), .ZN(
        n12580) );
  AOI22_X1 U15669 ( .A1(n9745), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10661), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12578) );
  AOI22_X1 U15670 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12686), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12577) );
  AOI22_X1 U15671 ( .A1(n10660), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12689), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12576) );
  NAND2_X1 U15672 ( .A1(n15583), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12574) );
  NAND2_X1 U15673 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n12573) );
  AND3_X1 U15674 ( .A1(n12574), .A2(n12573), .A3(n12693), .ZN(n12575) );
  NAND4_X1 U15675 ( .A1(n12578), .A2(n12577), .A3(n12576), .A4(n12575), .ZN(
        n12579) );
  AND2_X1 U15676 ( .A1(n12580), .A2(n12579), .ZN(n12581) );
  INV_X1 U15677 ( .A(n12581), .ZN(n14918) );
  INV_X1 U15678 ( .A(n12582), .ZN(n12584) );
  AND2_X1 U15679 ( .A1(n12582), .A2(n12581), .ZN(n12588) );
  INV_X1 U15680 ( .A(n12644), .ZN(n12583) );
  AOI211_X1 U15681 ( .C1(n14918), .C2(n12584), .A(n12588), .B(n12583), .ZN(
        n14920) );
  INV_X1 U15682 ( .A(n14930), .ZN(n12585) );
  NOR3_X1 U15683 ( .A1(n12586), .A2(n14918), .A3(n12585), .ZN(n12587) );
  INV_X1 U15684 ( .A(n12588), .ZN(n12603) );
  AOI22_X1 U15685 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10660), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12594) );
  AOI22_X1 U15686 ( .A1(n9745), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12686), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12593) );
  AOI22_X1 U15687 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12689), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12592) );
  NAND2_X1 U15688 ( .A1(n15583), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n12590) );
  NAND2_X1 U15689 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n12589) );
  AND3_X1 U15690 ( .A1(n12590), .A2(n12589), .A3(n12693), .ZN(n12591) );
  NAND4_X1 U15691 ( .A1(n12594), .A2(n12593), .A3(n12592), .A4(n12591), .ZN(
        n12602) );
  AOI22_X1 U15692 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10660), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12600) );
  AOI22_X1 U15693 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12686), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12599) );
  AOI22_X1 U15694 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12689), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12598) );
  NAND2_X1 U15695 ( .A1(n15583), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12596) );
  NAND2_X1 U15696 ( .A1(n9746), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n12595) );
  AND3_X1 U15697 ( .A1(n12657), .A2(n12596), .A3(n12595), .ZN(n12597) );
  NAND4_X1 U15698 ( .A1(n12600), .A2(n12599), .A3(n12598), .A4(n12597), .ZN(
        n12601) );
  NAND2_X1 U15699 ( .A1(n12602), .A2(n12601), .ZN(n12605) );
  NAND2_X1 U15700 ( .A1(n12603), .A2(n12605), .ZN(n12604) );
  NAND3_X1 U15701 ( .A1(n12609), .A2(n12644), .A3(n12604), .ZN(n12607) );
  INV_X1 U15702 ( .A(n12605), .ZN(n12606) );
  NAND2_X1 U15703 ( .A1(n19869), .A2(n12606), .ZN(n14912) );
  OAI21_X2 U15704 ( .B1(n14911), .B2(n14912), .A(n9810), .ZN(n12627) );
  INV_X1 U15705 ( .A(n12609), .ZN(n12624) );
  AOI22_X1 U15706 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10661), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12615) );
  AOI22_X1 U15707 ( .A1(n10660), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9744), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12614) );
  AOI22_X1 U15708 ( .A1(n12686), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12689), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12613) );
  NAND2_X1 U15709 ( .A1(n15583), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n12611) );
  NAND2_X1 U15710 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n12610) );
  AND3_X1 U15711 ( .A1(n12611), .A2(n12610), .A3(n12693), .ZN(n12612) );
  NAND4_X1 U15712 ( .A1(n12615), .A2(n12614), .A3(n12613), .A4(n12612), .ZN(
        n12623) );
  AOI22_X1 U15713 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n10660), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12621) );
  AOI22_X1 U15714 ( .A1(n9745), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12686), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12620) );
  AOI22_X1 U15715 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n15583), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12619) );
  NAND2_X1 U15716 ( .A1(n12689), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12617) );
  NAND2_X1 U15717 ( .A1(n9746), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n12616) );
  AND3_X1 U15718 ( .A1(n12657), .A2(n12617), .A3(n12616), .ZN(n12618) );
  NAND4_X1 U15719 ( .A1(n12621), .A2(n12620), .A3(n12619), .A4(n12618), .ZN(
        n12622) );
  AND2_X1 U15720 ( .A1(n12623), .A2(n12622), .ZN(n12626) );
  NAND2_X1 U15721 ( .A1(n12624), .A2(n12626), .ZN(n12629) );
  OAI211_X1 U15722 ( .C1(n12624), .C2(n12626), .A(n12644), .B(n12629), .ZN(
        n12628) );
  INV_X1 U15723 ( .A(n12628), .ZN(n12625) );
  NAND2_X1 U15724 ( .A1(n19869), .A2(n12626), .ZN(n14904) );
  INV_X1 U15725 ( .A(n12629), .ZN(n12645) );
  AOI22_X1 U15726 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10660), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12635) );
  AOI22_X1 U15727 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12686), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12634) );
  AOI22_X1 U15728 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12689), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12633) );
  NAND2_X1 U15729 ( .A1(n15583), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n12631) );
  NAND2_X1 U15730 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n12630) );
  AND3_X1 U15731 ( .A1(n12631), .A2(n12630), .A3(n12693), .ZN(n12632) );
  NAND4_X1 U15732 ( .A1(n12635), .A2(n12634), .A3(n12633), .A4(n12632), .ZN(
        n12643) );
  AOI22_X1 U15733 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n10660), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12641) );
  AOI22_X1 U15734 ( .A1(n9745), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12686), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12640) );
  AOI22_X1 U15735 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12689), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12639) );
  NAND2_X1 U15736 ( .A1(n15583), .A2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n12637) );
  NAND2_X1 U15737 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n12636) );
  AND3_X1 U15738 ( .A1(n12657), .A2(n12637), .A3(n12636), .ZN(n12638) );
  NAND4_X1 U15739 ( .A1(n12641), .A2(n12640), .A3(n12639), .A4(n12638), .ZN(
        n12642) );
  AND2_X1 U15740 ( .A1(n12643), .A2(n12642), .ZN(n12646) );
  NAND2_X1 U15741 ( .A1(n12645), .A2(n12646), .ZN(n14885) );
  OAI211_X1 U15742 ( .C1(n12645), .C2(n12646), .A(n12644), .B(n14885), .ZN(
        n12648) );
  XNOR2_X1 U15743 ( .A(n12647), .B(n12648), .ZN(n14893) );
  NAND2_X1 U15744 ( .A1(n19869), .A2(n12646), .ZN(n14895) );
  NOR2_X1 U15745 ( .A1(n12647), .A2(n12648), .ZN(n14887) );
  AOI22_X1 U15746 ( .A1(n10660), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9745), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12654) );
  AOI22_X1 U15747 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12686), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12653) );
  AOI22_X1 U15748 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12689), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12652) );
  NAND2_X1 U15749 ( .A1(n15583), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n12650) );
  NAND2_X1 U15750 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n12649) );
  AND3_X1 U15751 ( .A1(n12650), .A2(n12649), .A3(n12693), .ZN(n12651) );
  NAND4_X1 U15752 ( .A1(n12654), .A2(n12653), .A3(n12652), .A4(n12651), .ZN(
        n12663) );
  AOI22_X1 U15753 ( .A1(n10660), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9744), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12661) );
  AOI22_X1 U15754 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12686), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12660) );
  AOI22_X1 U15755 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12689), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12659) );
  NAND2_X1 U15756 ( .A1(n15583), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n12656) );
  NAND2_X1 U15757 ( .A1(n9746), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n12655) );
  AND3_X1 U15758 ( .A1(n12657), .A2(n12656), .A3(n12655), .ZN(n12658) );
  NAND4_X1 U15759 ( .A1(n12661), .A2(n12660), .A3(n12659), .A4(n12658), .ZN(
        n12662) );
  AND2_X1 U15760 ( .A1(n12663), .A2(n12662), .ZN(n12677) );
  AOI22_X1 U15761 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10660), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12665) );
  AOI22_X1 U15762 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12686), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12664) );
  NAND2_X1 U15763 ( .A1(n12665), .A2(n12664), .ZN(n12676) );
  AOI22_X1 U15764 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12689), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12667) );
  AOI21_X1 U15765 ( .B1(n9746), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A(
        n12693), .ZN(n12666) );
  OAI211_X1 U15766 ( .C1(n12541), .C2(n10406), .A(n12667), .B(n12666), .ZN(
        n12675) );
  AOI22_X1 U15767 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10660), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12669) );
  AOI22_X1 U15768 ( .A1(n9745), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12686), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12668) );
  NAND2_X1 U15769 ( .A1(n12669), .A2(n12668), .ZN(n12674) );
  AOI22_X1 U15770 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12689), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12672) );
  NAND2_X1 U15771 ( .A1(n15583), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n12671) );
  NAND2_X1 U15772 ( .A1(n12690), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n12670) );
  NAND4_X1 U15773 ( .A1(n12672), .A2(n12693), .A3(n12671), .A4(n12670), .ZN(
        n12673) );
  OAI22_X1 U15774 ( .A1(n12676), .A2(n12675), .B1(n12674), .B2(n12673), .ZN(
        n12679) );
  INV_X1 U15775 ( .A(n12677), .ZN(n14888) );
  NOR3_X1 U15776 ( .A1(n14885), .A2(n19869), .A3(n14888), .ZN(n12678) );
  XOR2_X1 U15777 ( .A(n12679), .B(n12678), .Z(n14879) );
  INV_X1 U15778 ( .A(n12678), .ZN(n12680) );
  AOI22_X1 U15779 ( .A1(n10660), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9745), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12682) );
  AOI22_X1 U15780 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12686), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12681) );
  NAND2_X1 U15781 ( .A1(n12682), .A2(n12681), .ZN(n12698) );
  INV_X1 U15782 ( .A(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12685) );
  AOI22_X1 U15783 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12689), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12684) );
  AOI21_X1 U15784 ( .B1(n9746), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n12693), .ZN(n12683) );
  OAI211_X1 U15785 ( .C1(n12541), .C2(n12685), .A(n12684), .B(n12683), .ZN(
        n12697) );
  AOI22_X1 U15786 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10660), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12688) );
  AOI22_X1 U15787 ( .A1(n9744), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12686), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12687) );
  NAND2_X1 U15788 ( .A1(n12688), .A2(n12687), .ZN(n12696) );
  AOI22_X1 U15789 ( .A1(n10661), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12689), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12694) );
  NAND2_X1 U15790 ( .A1(n15583), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n12692) );
  NAND2_X1 U15791 ( .A1(n9761), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n12691) );
  NAND4_X1 U15792 ( .A1(n12694), .A2(n12693), .A3(n12692), .A4(n12691), .ZN(
        n12695) );
  OAI22_X1 U15793 ( .A1(n12698), .A2(n12697), .B1(n12696), .B2(n12695), .ZN(
        n12699) );
  INV_X1 U15794 ( .A(n15582), .ZN(n16271) );
  NAND2_X1 U15795 ( .A1(n12180), .A2(n19867), .ZN(n16262) );
  NOR2_X1 U15796 ( .A1(n16265), .A2(n16262), .ZN(n12702) );
  AOI21_X1 U15797 ( .B1(n16276), .B2(n16271), .A(n12702), .ZN(n14093) );
  NAND2_X1 U15798 ( .A1(n12703), .A2(n10723), .ZN(n12704) );
  NAND2_X1 U15799 ( .A1(n14093), .A2(n12704), .ZN(n12705) );
  AND2_X1 U15800 ( .A1(n19237), .A2(n12707), .ZN(n12708) );
  NOR4_X1 U15801 ( .A1(P2_ADDRESS_REG_16__SCAN_IN), .A2(
        P2_ADDRESS_REG_15__SCAN_IN), .A3(P2_ADDRESS_REG_14__SCAN_IN), .A4(
        P2_ADDRESS_REG_13__SCAN_IN), .ZN(n12712) );
  NOR4_X1 U15802 ( .A1(P2_ADDRESS_REG_20__SCAN_IN), .A2(
        P2_ADDRESS_REG_19__SCAN_IN), .A3(P2_ADDRESS_REG_18__SCAN_IN), .A4(
        P2_ADDRESS_REG_17__SCAN_IN), .ZN(n12711) );
  NOR4_X1 U15803 ( .A1(P2_ADDRESS_REG_7__SCAN_IN), .A2(
        P2_ADDRESS_REG_6__SCAN_IN), .A3(P2_ADDRESS_REG_5__SCAN_IN), .A4(
        P2_ADDRESS_REG_4__SCAN_IN), .ZN(n12710) );
  NOR4_X1 U15804 ( .A1(P2_ADDRESS_REG_12__SCAN_IN), .A2(
        P2_ADDRESS_REG_11__SCAN_IN), .A3(P2_ADDRESS_REG_10__SCAN_IN), .A4(
        P2_ADDRESS_REG_9__SCAN_IN), .ZN(n12709) );
  NAND4_X1 U15805 ( .A1(n12712), .A2(n12711), .A3(n12710), .A4(n12709), .ZN(
        n12717) );
  NOR4_X1 U15806 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_1__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n12715) );
  NOR4_X1 U15807 ( .A1(P2_ADDRESS_REG_24__SCAN_IN), .A2(
        P2_ADDRESS_REG_23__SCAN_IN), .A3(P2_ADDRESS_REG_22__SCAN_IN), .A4(
        P2_ADDRESS_REG_21__SCAN_IN), .ZN(n12714) );
  NOR4_X1 U15808 ( .A1(P2_ADDRESS_REG_28__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P2_ADDRESS_REG_26__SCAN_IN), .A4(
        P2_ADDRESS_REG_25__SCAN_IN), .ZN(n12713) );
  INV_X1 U15809 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19763) );
  NAND4_X1 U15810 ( .A1(n12715), .A2(n12714), .A3(n12713), .A4(n19763), .ZN(
        n12716) );
  NAND2_X1 U15811 ( .A1(n13830), .A2(BUF2_REG_14__SCAN_IN), .ZN(n12720) );
  INV_X1 U15812 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n12718) );
  OR2_X1 U15813 ( .A1(n13830), .A2(n12718), .ZN(n12719) );
  NAND2_X1 U15814 ( .A1(n12720), .A2(n12719), .ZN(n19184) );
  INV_X1 U15815 ( .A(n19184), .ZN(n12722) );
  INV_X1 U15816 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n12721) );
  OAI22_X1 U15817 ( .A1(n16141), .A2(n12722), .B1(n19072), .B2(n12721), .ZN(
        n12723) );
  AOI21_X1 U15818 ( .B1(n15260), .B2(n19106), .A(n12723), .ZN(n12726) );
  NAND2_X1 U15819 ( .A1(n19072), .A2(n12724), .ZN(n13339) );
  AOI22_X1 U15820 ( .A1(n19047), .A2(BUF2_REG_30__SCAN_IN), .B1(n19049), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n12725) );
  AND2_X1 U15821 ( .A1(n12726), .A2(n12725), .ZN(n12727) );
  OAI21_X1 U15822 ( .B1(n14203), .B2(n19082), .A(n12727), .ZN(P2_U2889) );
  NAND2_X1 U15823 ( .A1(n15032), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12729) );
  INV_X1 U15824 ( .A(n12782), .ZN(n12730) );
  NAND2_X1 U15825 ( .A1(n12730), .A2(n16223), .ZN(n12773) );
  NAND2_X1 U15826 ( .A1(n15278), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12737) );
  AOI21_X1 U15827 ( .B1(n15426), .B2(n12737), .A(n15294), .ZN(n15262) );
  OAI21_X1 U15828 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15556), .A(
        n15262), .ZN(n12731) );
  INV_X1 U15829 ( .A(n12731), .ZN(n12750) );
  AOI222_X1 U15830 ( .A1(n10337), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n12733), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n10267), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12734) );
  INV_X1 U15831 ( .A(n12734), .ZN(n12735) );
  NAND2_X1 U15832 ( .A1(n19206), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n12776) );
  NOR2_X1 U15833 ( .A1(n15292), .A2(n12737), .ZN(n15263) );
  NAND3_X1 U15834 ( .A1(n15263), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n12745), .ZN(n12738) );
  OAI211_X1 U15835 ( .C1(n16069), .C2(n16197), .A(n12776), .B(n12738), .ZN(
        n12739) );
  INV_X1 U15836 ( .A(n12739), .ZN(n12749) );
  NAND2_X1 U15837 ( .A1(n14880), .A2(n12740), .ZN(n12747) );
  AOI22_X1 U15838 ( .A1(n12741), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n12744) );
  NAND2_X1 U15839 ( .A1(n12742), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n12743) );
  OAI211_X1 U15840 ( .C1(n9719), .C2(n12745), .A(n12744), .B(n12743), .ZN(
        n12746) );
  OAI211_X1 U15841 ( .C1(n12745), .C2(n12750), .A(n12749), .B(n12748), .ZN(
        n12751) );
  INV_X1 U15842 ( .A(n12751), .ZN(n12772) );
  NAND2_X1 U15843 ( .A1(n15056), .A2(n12298), .ZN(n12754) );
  XNOR2_X1 U15844 ( .A(n12758), .B(n12757), .ZN(n12761) );
  AOI21_X1 U15845 ( .B1(n12759), .B2(n12762), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15034) );
  INV_X1 U15846 ( .A(n12761), .ZN(n16074) );
  NAND3_X1 U15847 ( .A1(n16074), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n12762), .ZN(n15046) );
  NOR2_X1 U15848 ( .A1(n12766), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12767) );
  MUX2_X1 U15849 ( .A(n12768), .B(n12767), .S(n19237), .Z(n16066) );
  NAND2_X1 U15850 ( .A1(n16066), .A2(n12762), .ZN(n12769) );
  XNOR2_X1 U15851 ( .A(n12770), .B(n9801), .ZN(n12779) );
  NAND2_X1 U15852 ( .A1(n12779), .A2(n19219), .ZN(n12771) );
  NAND3_X1 U15853 ( .A1(n12773), .A2(n12772), .A3(n12771), .ZN(P2_U3015) );
  NAND2_X1 U15854 ( .A1(n19190), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12775) );
  OAI211_X1 U15855 ( .C1(n12777), .C2(n19205), .A(n12776), .B(n12775), .ZN(
        n12778) );
  NAND2_X1 U15856 ( .A1(n12779), .A2(n16190), .ZN(n12780) );
  OAI211_X1 U15857 ( .C1(n12782), .C2(n19197), .A(n12781), .B(n12780), .ZN(
        P2_U2983) );
  AOI22_X1 U15858 ( .A1(n12834), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12787) );
  INV_X2 U15859 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18827) );
  INV_X2 U15860 ( .A(n17083), .ZN(n12832) );
  AOI22_X1 U15861 ( .A1(n12832), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12786) );
  NOR2_X2 U15862 ( .A1(n12789), .A2(n12791), .ZN(n17185) );
  AOI22_X1 U15863 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12785) );
  AOI22_X1 U15864 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12784) );
  NAND4_X1 U15865 ( .A1(n12787), .A2(n12786), .A3(n12785), .A4(n12784), .ZN(
        n12800) );
  INV_X2 U15866 ( .A(n12868), .ZN(n17188) );
  AOI22_X1 U15867 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12798) );
  INV_X2 U15868 ( .A(n16791), .ZN(n16876) );
  AOI22_X1 U15869 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n16876), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12797) );
  INV_X2 U15870 ( .A(n9767), .ZN(n17172) );
  AOI22_X1 U15871 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17172), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12796) );
  AOI22_X1 U15872 ( .A1(n17165), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n16869), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12795) );
  NAND4_X1 U15873 ( .A1(n12798), .A2(n12797), .A3(n12796), .A4(n12795), .ZN(
        n12799) );
  INV_X2 U15874 ( .A(n14086), .ZN(n17084) );
  AOI22_X1 U15875 ( .A1(n17084), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12804) );
  AOI22_X1 U15876 ( .A1(n16891), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12803) );
  AOI22_X1 U15877 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12802) );
  INV_X1 U15878 ( .A(n12835), .ZN(n17117) );
  INV_X2 U15879 ( .A(n17117), .ZN(n17166) );
  AOI22_X1 U15880 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n16876), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12801) );
  NAND4_X1 U15881 ( .A1(n12804), .A2(n12803), .A3(n12802), .A4(n12801), .ZN(
        n12810) );
  AOI22_X1 U15882 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12808) );
  AOI22_X1 U15883 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17172), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12807) );
  AOI22_X1 U15884 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12806) );
  AOI22_X1 U15885 ( .A1(n17165), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12805) );
  NAND4_X1 U15886 ( .A1(n12808), .A2(n12807), .A3(n12806), .A4(n12805), .ZN(
        n12809) );
  AOI22_X1 U15887 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n16876), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12814) );
  AOI22_X1 U15888 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12813) );
  AOI22_X1 U15889 ( .A1(n17084), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12812) );
  AOI22_X1 U15890 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12811) );
  NAND4_X1 U15891 ( .A1(n12814), .A2(n12813), .A3(n12812), .A4(n12811), .ZN(
        n12820) );
  AOI22_X1 U15892 ( .A1(n12834), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12818) );
  AOI22_X1 U15893 ( .A1(n17165), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12817) );
  INV_X2 U15894 ( .A(n9767), .ZN(n17193) );
  AOI22_X1 U15895 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n16869), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12816) );
  AOI22_X1 U15896 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12815) );
  NAND4_X1 U15897 ( .A1(n12818), .A2(n12817), .A3(n12816), .A4(n12815), .ZN(
        n12819) );
  AOI22_X1 U15898 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n12790), .B1(
        P3_INSTQUEUE_REG_6__1__SCAN_IN), .B2(n16864), .ZN(n12824) );
  AOI22_X1 U15899 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12823) );
  INV_X2 U15900 ( .A(n17083), .ZN(n17174) );
  AOI22_X1 U15901 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17174), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n16876), .ZN(n12822) );
  AOI22_X1 U15902 ( .A1(n16910), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17167), .ZN(n12821) );
  AOI22_X1 U15903 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17189), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n17173), .ZN(n12827) );
  AOI22_X1 U15904 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n16891), .B1(
        n17172), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12826) );
  NAND2_X1 U15905 ( .A1(n12834), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n12825) );
  INV_X1 U15906 ( .A(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n21028) );
  AOI22_X1 U15907 ( .A1(n12788), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12828) );
  OAI21_X1 U15908 ( .B1(n21028), .B2(n17117), .A(n12828), .ZN(n12829) );
  INV_X1 U15909 ( .A(n12829), .ZN(n12830) );
  AOI22_X1 U15910 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12843) );
  AOI22_X1 U15911 ( .A1(n16910), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17172), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12842) );
  AOI22_X1 U15912 ( .A1(n16876), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n16864), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12831) );
  OAI21_X1 U15913 ( .B1(n10128), .B2(n17232), .A(n12831), .ZN(n12841) );
  AOI22_X1 U15914 ( .A1(n12832), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12840) );
  AOI22_X1 U15915 ( .A1(n12834), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12833), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12839) );
  AOI22_X1 U15916 ( .A1(n16992), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12835), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12838) );
  AOI22_X1 U15917 ( .A1(n12790), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17167), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12837) );
  NAND2_X1 U15918 ( .A1(n17391), .A2(n13046), .ZN(n12865) );
  AOI22_X1 U15919 ( .A1(n16910), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12853) );
  INV_X2 U15920 ( .A(n10128), .ZN(n17184) );
  AOI22_X1 U15921 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12852) );
  AOI22_X1 U15922 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12844) );
  OAI21_X1 U15923 ( .B1(n12868), .B2(n21022), .A(n12844), .ZN(n12850) );
  AOI22_X1 U15924 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12848) );
  AOI22_X1 U15925 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n16876), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12847) );
  AOI22_X1 U15926 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12846) );
  AOI22_X1 U15927 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n16869), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12845) );
  NAND4_X1 U15928 ( .A1(n12848), .A2(n12847), .A3(n12846), .A4(n12845), .ZN(
        n12849) );
  AOI211_X1 U15929 ( .C1(n17164), .C2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n12850), .B(n12849), .ZN(n12851) );
  NAND3_X1 U15930 ( .A1(n12853), .A2(n12852), .A3(n12851), .ZN(n17375) );
  NAND2_X1 U15931 ( .A1(n12886), .A2(n17375), .ZN(n12864) );
  AOI22_X1 U15932 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17193), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12863) );
  AOI22_X1 U15933 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12862) );
  INV_X1 U15934 ( .A(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n20865) );
  AOI22_X1 U15935 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12854) );
  OAI21_X1 U15936 ( .B1(n16909), .B2(n20865), .A(n12854), .ZN(n12860) );
  AOI22_X1 U15937 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n16876), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12858) );
  AOI22_X1 U15938 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12857) );
  AOI22_X1 U15939 ( .A1(n16910), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12856) );
  AOI22_X1 U15940 ( .A1(n17084), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12855) );
  NAND4_X1 U15941 ( .A1(n12858), .A2(n12857), .A3(n12856), .A4(n12855), .ZN(
        n12859) );
  AOI211_X1 U15942 ( .C1(n17183), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n12860), .B(n12859), .ZN(n12861) );
  NAND3_X1 U15943 ( .A1(n12863), .A2(n12862), .A3(n12861), .ZN(n17367) );
  NAND2_X1 U15944 ( .A1(n12889), .A2(n17367), .ZN(n12892) );
  NOR2_X1 U15945 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17782), .ZN(
        n12907) );
  AOI21_X1 U15946 ( .B1(n17782), .B2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A(
        n12907), .ZN(n12913) );
  INV_X1 U15947 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17886) );
  INV_X1 U15948 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18011) );
  NAND2_X1 U15949 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18076) );
  INV_X1 U15950 ( .A(n18076), .ZN(n17747) );
  NAND2_X1 U15951 ( .A1(n17747), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18059) );
  INV_X1 U15952 ( .A(n18059), .ZN(n18046) );
  NAND2_X1 U15953 ( .A1(n18046), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17710) );
  INV_X1 U15954 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n20828) );
  NOR2_X1 U15955 ( .A1(n17710), .A2(n20828), .ZN(n18029) );
  NAND2_X1 U15956 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18029), .ZN(
        n18017) );
  INV_X1 U15957 ( .A(n18017), .ZN(n18009) );
  NAND2_X1 U15958 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18009), .ZN(
        n17994) );
  XOR2_X1 U15959 ( .A(n17372), .B(n12864), .Z(n17816) );
  XOR2_X1 U15960 ( .A(n17380), .B(n12865), .Z(n12882) );
  NAND2_X1 U15961 ( .A1(n13041), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12879) );
  XNOR2_X1 U15962 ( .A(n17391), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17867) );
  AOI22_X1 U15963 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12872) );
  INV_X1 U15964 ( .A(n12868), .ZN(n17152) );
  AOI22_X1 U15965 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12871) );
  AOI22_X1 U15966 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n16876), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12870) );
  AOI22_X1 U15967 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n16864), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12869) );
  NAND4_X1 U15968 ( .A1(n12872), .A2(n12871), .A3(n12870), .A4(n12869), .ZN(
        n12878) );
  AOI22_X1 U15969 ( .A1(n16891), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12876) );
  AOI22_X1 U15970 ( .A1(n16910), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17193), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12875) );
  AOI22_X1 U15971 ( .A1(n12834), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n16869), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12874) );
  AOI22_X1 U15972 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12832), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12873) );
  NAND4_X1 U15973 ( .A1(n12876), .A2(n12875), .A3(n12874), .A4(n12873), .ZN(
        n12877) );
  INV_X1 U15974 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n21021) );
  NOR2_X1 U15975 ( .A1(n17876), .A2(n21021), .ZN(n17875) );
  NAND2_X1 U15976 ( .A1(n17867), .A2(n17875), .ZN(n17866) );
  NAND2_X1 U15977 ( .A1(n12879), .A2(n17866), .ZN(n17858) );
  NAND2_X1 U15978 ( .A1(n17859), .A2(n17858), .ZN(n17857) );
  NAND2_X1 U15979 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12880), .ZN(
        n12881) );
  NAND2_X1 U15980 ( .A1(n17857), .A2(n12881), .ZN(n12884) );
  NAND2_X1 U15981 ( .A1(n12882), .A2(n12884), .ZN(n12885) );
  XNOR2_X1 U15982 ( .A(n12884), .B(n12883), .ZN(n17847) );
  NAND2_X1 U15983 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n17847), .ZN(
        n17846) );
  XOR2_X1 U15984 ( .A(n17375), .B(n12886), .Z(n12887) );
  NAND2_X1 U15985 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12887), .ZN(
        n12888) );
  INV_X1 U15986 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n20760) );
  XOR2_X1 U15987 ( .A(n17367), .B(n12889), .Z(n12890) );
  XOR2_X1 U15988 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n12890), .Z(
        n17802) );
  NAND2_X1 U15989 ( .A1(n17803), .A2(n17802), .ZN(n17801) );
  NAND2_X1 U15990 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12890), .ZN(
        n12891) );
  AOI21_X1 U15991 ( .B1(n16337), .B2(n12892), .A(n17782), .ZN(n12895) );
  NAND2_X1 U15992 ( .A1(n12895), .A2(n12894), .ZN(n12896) );
  INV_X1 U15993 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18100) );
  INV_X1 U15994 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18084) );
  NAND2_X1 U15995 ( .A1(n18100), .A2(n18084), .ZN(n17756) );
  INV_X1 U15996 ( .A(n17756), .ZN(n17693) );
  NOR4_X1 U15997 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12897) );
  INV_X1 U15998 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18016) );
  NAND4_X1 U15999 ( .A1(n12898), .A2(n17693), .A3(n12897), .A4(n18016), .ZN(
        n12899) );
  NAND2_X1 U16000 ( .A1(n12900), .A2(n12899), .ZN(n17674) );
  INV_X1 U16001 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n21020) );
  NOR2_X1 U16002 ( .A1(n21020), .A2(n18011), .ZN(n17989) );
  NAND2_X1 U16003 ( .A1(n17989), .A2(n17675), .ZN(n17619) );
  INV_X1 U16004 ( .A(n17989), .ZN(n17657) );
  NAND2_X1 U16005 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17947) );
  INV_X1 U16006 ( .A(n17947), .ZN(n17961) );
  NAND3_X1 U16007 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n17961), .ZN(n17601) );
  INV_X1 U16008 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17954) );
  NOR2_X1 U16009 ( .A1(n17601), .A2(n17954), .ZN(n17580) );
  NAND2_X1 U16010 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n17580), .ZN(
        n17921) );
  NOR2_X1 U16011 ( .A1(n17657), .A2(n17921), .ZN(n17539) );
  NAND2_X1 U16012 ( .A1(n17675), .A2(n17539), .ZN(n12901) );
  NOR2_X1 U16013 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17782), .ZN(
        n17649) );
  INV_X1 U16014 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17980) );
  NAND2_X1 U16015 ( .A1(n17649), .A2(n17980), .ZN(n17627) );
  NOR2_X1 U16016 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17627), .ZN(
        n17620) );
  INV_X1 U16017 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17946) );
  NAND2_X1 U16018 ( .A1(n17620), .A2(n17946), .ZN(n17600) );
  NAND2_X1 U16019 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17885) );
  NAND2_X1 U16020 ( .A1(n17782), .A2(n17885), .ZN(n12903) );
  INV_X1 U16021 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16317) );
  NAND2_X1 U16022 ( .A1(n10129), .A2(n16317), .ZN(n12911) );
  INV_X1 U16023 ( .A(n12911), .ZN(n12909) );
  INV_X1 U16024 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17892) );
  NOR3_X1 U16025 ( .A1(n17892), .A2(n12905), .A3(n16317), .ZN(n13072) );
  NAND2_X1 U16026 ( .A1(n16338), .A2(n13072), .ZN(n12910) );
  NAND2_X1 U16027 ( .A1(n17782), .A2(n12910), .ZN(n12912) );
  OAI21_X1 U16028 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n12907), .A(
        n12912), .ZN(n12908) );
  INV_X1 U16029 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n21009) );
  NAND2_X1 U16030 ( .A1(n21009), .A2(n15740), .ZN(n15739) );
  INV_X1 U16031 ( .A(n16337), .ZN(n17362) );
  AOI22_X1 U16032 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12917) );
  AOI22_X1 U16033 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17193), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12916) );
  AOI22_X1 U16034 ( .A1(n17190), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12915) );
  AOI22_X1 U16035 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n17167), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12914) );
  NAND4_X1 U16036 ( .A1(n12917), .A2(n12916), .A3(n12915), .A4(n12914), .ZN(
        n12923) );
  AOI22_X1 U16037 ( .A1(n17165), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12921) );
  AOI22_X1 U16038 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17164), .B1(
        n9720), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12920) );
  AOI22_X1 U16039 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n17188), .B1(
        n12832), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12919) );
  AOI22_X1 U16040 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12918) );
  NAND4_X1 U16041 ( .A1(n12921), .A2(n12920), .A3(n12919), .A4(n12918), .ZN(
        n12922) );
  NOR2_X1 U16042 ( .A1(n20757), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n16456) );
  NAND2_X1 U16043 ( .A1(n16456), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18708) );
  OAI22_X1 U16044 ( .A1(n18827), .A2(n18659), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13036) );
  INV_X1 U16045 ( .A(n13036), .ZN(n12936) );
  INV_X1 U16046 ( .A(n12935), .ZN(n12924) );
  NOR2_X1 U16047 ( .A1(n12936), .A2(n12924), .ZN(n12925) );
  AOI22_X1 U16048 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(n18663), .B2(n18820), .ZN(
        n12930) );
  OAI21_X1 U16049 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18820), .A(
        n12926), .ZN(n12927) );
  OAI22_X1 U16050 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18207), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n12927), .ZN(n12933) );
  NOR2_X1 U16051 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18207), .ZN(
        n12928) );
  NAND2_X1 U16052 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n12927), .ZN(
        n12932) );
  AOI22_X1 U16053 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n12933), .B1(
        n12928), .B2(n12932), .ZN(n13038) );
  OAI21_X1 U16054 ( .B1(n12931), .B2(n12930), .A(n13038), .ZN(n12929) );
  AOI21_X1 U16055 ( .B1(n12931), .B2(n12930), .A(n12929), .ZN(n12938) );
  INV_X1 U16056 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16785) );
  AND2_X1 U16057 ( .A1(n12932), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12934) );
  OAI22_X1 U16058 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n16785), .B1(
        n12934), .B2(n12933), .ZN(n12937) );
  NOR2_X1 U16059 ( .A1(n12938), .A2(n12937), .ZN(n13039) );
  AOI21_X1 U16060 ( .B1(n21023), .B2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(
        n12935), .ZN(n13037) );
  INV_X1 U16061 ( .A(n13037), .ZN(n12940) );
  XNOR2_X1 U16062 ( .A(n12936), .B(n12935), .ZN(n12939) );
  OAI21_X1 U16063 ( .B1(n13039), .B2(n12940), .A(n18682), .ZN(n18688) );
  AOI22_X1 U16064 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12944) );
  AOI22_X1 U16065 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17172), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12943) );
  AOI22_X1 U16066 ( .A1(n16891), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12942) );
  AOI22_X1 U16067 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12941) );
  NAND4_X1 U16068 ( .A1(n12944), .A2(n12943), .A3(n12942), .A4(n12941), .ZN(
        n12950) );
  AOI22_X1 U16069 ( .A1(n17165), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12832), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12948) );
  AOI22_X1 U16070 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n16869), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12947) );
  AOI22_X1 U16071 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n16876), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12946) );
  AOI22_X1 U16072 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12945) );
  NAND4_X1 U16073 ( .A1(n12948), .A2(n12947), .A3(n12946), .A4(n12945), .ZN(
        n12949) );
  AOI22_X1 U16074 ( .A1(n16891), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12954) );
  AOI22_X1 U16075 ( .A1(n17165), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12867), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12953) );
  INV_X2 U16076 ( .A(n16791), .ZN(n17190) );
  AOI22_X1 U16077 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12952) );
  AOI22_X1 U16078 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12951) );
  NAND4_X1 U16079 ( .A1(n12954), .A2(n12953), .A3(n12952), .A4(n12951), .ZN(
        n12961) );
  AOI22_X1 U16080 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12955) );
  OAI21_X1 U16081 ( .B1(n9767), .B2(n20743), .A(n12955), .ZN(n12960) );
  AOI22_X1 U16082 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12958) );
  AOI22_X1 U16083 ( .A1(n12834), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12832), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12957) );
  NAND3_X1 U16084 ( .A1(n12958), .A2(n12957), .A3(n12956), .ZN(n12959) );
  AOI22_X1 U16085 ( .A1(n16891), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17172), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12971) );
  AOI22_X1 U16086 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12970) );
  AOI22_X1 U16087 ( .A1(n17084), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12962) );
  OAI21_X1 U16088 ( .B1(n16909), .B2(n21022), .A(n12962), .ZN(n12968) );
  AOI22_X1 U16089 ( .A1(n12834), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12832), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12966) );
  AOI22_X1 U16090 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17189), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12965) );
  AOI22_X1 U16091 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n16869), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12964) );
  AOI22_X1 U16092 ( .A1(n16910), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12963) );
  NAND4_X1 U16093 ( .A1(n12966), .A2(n12965), .A3(n12964), .A4(n12963), .ZN(
        n12967) );
  AOI211_X1 U16094 ( .C1(n17188), .C2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n12968), .B(n12967), .ZN(n12969) );
  NAND3_X1 U16095 ( .A1(n12971), .A2(n12970), .A3(n12969), .ZN(n15641) );
  NOR2_X1 U16096 ( .A1(n18853), .A2(n15641), .ZN(n15666) );
  AOI22_X1 U16097 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12975) );
  AOI22_X1 U16098 ( .A1(n16910), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12974) );
  AOI22_X1 U16099 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17172), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12973) );
  AOI22_X1 U16100 ( .A1(n17084), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12972) );
  NAND4_X1 U16101 ( .A1(n12975), .A2(n12974), .A3(n12973), .A4(n12972), .ZN(
        n12981) );
  AOI22_X1 U16102 ( .A1(n12834), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12979) );
  AOI22_X1 U16103 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12832), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12978) );
  AOI22_X1 U16104 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n16869), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12977) );
  AOI22_X1 U16105 ( .A1(n16891), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12976) );
  NAND4_X1 U16106 ( .A1(n12979), .A2(n12978), .A3(n12977), .A4(n12976), .ZN(
        n12980) );
  AOI22_X1 U16107 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12985) );
  AOI22_X1 U16108 ( .A1(n16891), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12984) );
  AOI22_X1 U16109 ( .A1(n12834), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12983) );
  AOI22_X1 U16110 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12982) );
  NAND4_X1 U16111 ( .A1(n12985), .A2(n12984), .A3(n12983), .A4(n12982), .ZN(
        n12991) );
  AOI22_X1 U16112 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12989) );
  AOI22_X1 U16113 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n16869), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12988) );
  AOI22_X1 U16114 ( .A1(n9753), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12987) );
  AOI22_X1 U16115 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17172), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12986) );
  NAND4_X1 U16116 ( .A1(n12989), .A2(n12988), .A3(n12987), .A4(n12986), .ZN(
        n12990) );
  NOR2_X1 U16117 ( .A1(n18238), .A2(n18234), .ZN(n13024) );
  AOI22_X1 U16118 ( .A1(n16891), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13003) );
  INV_X2 U16119 ( .A(n17132), .ZN(n17164) );
  AOI22_X1 U16120 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n13002) );
  INV_X1 U16121 ( .A(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n20938) );
  AOI22_X1 U16122 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12993) );
  OAI21_X1 U16123 ( .B1(n9767), .B2(n20938), .A(n12993), .ZN(n13000) );
  AOI22_X1 U16124 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12998) );
  AOI22_X1 U16125 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12997) );
  AOI22_X1 U16126 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12996) );
  AOI22_X1 U16127 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12995) );
  NAND4_X1 U16128 ( .A1(n12998), .A2(n12997), .A3(n12996), .A4(n12995), .ZN(
        n12999) );
  NAND4_X1 U16129 ( .A1(n18225), .A2(n15666), .A3(n13024), .A4(n17330), .ZN(
        n13027) );
  INV_X1 U16130 ( .A(n15641), .ZN(n18229) );
  NAND2_X1 U16131 ( .A1(n17248), .A2(n18238), .ZN(n15769) );
  INV_X1 U16132 ( .A(n15769), .ZN(n18655) );
  INV_X1 U16133 ( .A(n13029), .ZN(n13015) );
  AOI22_X1 U16134 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13013) );
  AOI22_X1 U16135 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n16876), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13012) );
  AOI22_X1 U16136 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13004) );
  OAI21_X1 U16137 ( .B1(n17083), .B2(n17232), .A(n13004), .ZN(n13010) );
  AOI22_X1 U16138 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n16910), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n13008) );
  AOI22_X1 U16139 ( .A1(n16891), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13007) );
  AOI22_X1 U16140 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n16869), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13006) );
  AOI22_X1 U16141 ( .A1(n17057), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n13005) );
  NAND4_X1 U16142 ( .A1(n13008), .A2(n13007), .A3(n13006), .A4(n13005), .ZN(
        n13009) );
  AOI211_X1 U16143 ( .C1(n9720), .C2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A(
        n13010), .B(n13009), .ZN(n13011) );
  NAND3_X1 U16144 ( .A1(n13013), .A2(n13012), .A3(n13011), .ZN(n15678) );
  AOI211_X1 U16145 ( .C1(n18229), .C2(n18655), .A(n13015), .B(n15678), .ZN(
        n15669) );
  NOR3_X1 U16146 ( .A1(n18648), .A2(n15667), .A3(n15678), .ZN(n13017) );
  NOR2_X1 U16147 ( .A1(n18234), .A2(n15678), .ZN(n15684) );
  NOR2_X1 U16148 ( .A1(n13017), .A2(n15684), .ZN(n13026) );
  NAND2_X1 U16149 ( .A1(n18217), .A2(n18853), .ZN(n15663) );
  AOI21_X1 U16150 ( .B1(n17330), .B2(n15769), .A(n15663), .ZN(n15670) );
  NOR2_X1 U16151 ( .A1(n13026), .A2(n15670), .ZN(n13014) );
  OR2_X1 U16152 ( .A1(n13014), .A2(n18225), .ZN(n13022) );
  NOR2_X1 U16153 ( .A1(n13015), .A2(n13025), .ZN(n13016) );
  NAND2_X1 U16154 ( .A1(n18225), .A2(n13016), .ZN(n13021) );
  NAND2_X1 U16155 ( .A1(n13017), .A2(n18213), .ZN(n13019) );
  OAI21_X1 U16156 ( .B1(n18245), .B2(n13024), .A(n15641), .ZN(n13018) );
  NAND2_X1 U16157 ( .A1(n18234), .A2(n13030), .ZN(n15662) );
  NAND2_X1 U16158 ( .A1(n13029), .A2(n15663), .ZN(n18867) );
  NOR2_X1 U16159 ( .A1(n18217), .A2(n13031), .ZN(n13033) );
  XNOR2_X1 U16160 ( .A(n17448), .B(n18221), .ZN(n15679) );
  NAND3_X1 U16161 ( .A1(n13038), .A2(n13037), .A3(n13036), .ZN(n13040) );
  NAND2_X1 U16162 ( .A1(n13040), .A2(n13039), .ZN(n15639) );
  NOR2_X1 U16163 ( .A1(n13044), .A2(n17380), .ZN(n13053) );
  NAND2_X1 U16164 ( .A1(n13053), .A2(n17375), .ZN(n13043) );
  NOR2_X1 U16165 ( .A1(n17372), .A2(n13043), .ZN(n13056) );
  NAND2_X1 U16166 ( .A1(n13056), .A2(n17367), .ZN(n13042) );
  NOR2_X1 U16167 ( .A1(n16337), .A2(n13042), .ZN(n13063) );
  XOR2_X1 U16168 ( .A(n13042), .B(n16337), .Z(n17795) );
  XOR2_X1 U16169 ( .A(n13043), .B(n17372), .Z(n17821) );
  XOR2_X1 U16170 ( .A(n17380), .B(n13044), .Z(n13045) );
  NAND2_X1 U16171 ( .A1(n13045), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13052) );
  XOR2_X1 U16172 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n13045), .Z(
        n17844) );
  INV_X1 U16173 ( .A(n13046), .ZN(n17383) );
  NAND2_X1 U16174 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13048), .ZN(
        n13051) );
  INV_X1 U16175 ( .A(n17876), .ZN(n15770) );
  AOI21_X1 U16176 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n17391), .A(
        n15770), .ZN(n13050) );
  NOR2_X1 U16177 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n17391), .ZN(
        n13049) );
  AOI221_X1 U16178 ( .B1(n15770), .B2(n17391), .C1(n13050), .C2(n21021), .A(
        n13049), .ZN(n17855) );
  NAND2_X1 U16179 ( .A1(n13051), .A2(n17854), .ZN(n17843) );
  NAND2_X1 U16180 ( .A1(n17844), .A2(n17843), .ZN(n17842) );
  NAND2_X1 U16181 ( .A1(n13052), .A2(n17842), .ZN(n13054) );
  NAND2_X1 U16182 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13054), .ZN(
        n13055) );
  XOR2_X1 U16183 ( .A(n13053), .B(n17375), .Z(n17832) );
  INV_X1 U16184 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18152) );
  XNOR2_X1 U16185 ( .A(n18152), .B(n13054), .ZN(n17831) );
  NAND2_X1 U16186 ( .A1(n17832), .A2(n17831), .ZN(n17830) );
  XOR2_X1 U16187 ( .A(n13056), .B(n17367), .Z(n13058) );
  NAND2_X1 U16188 ( .A1(n13057), .A2(n13058), .ZN(n13059) );
  NAND2_X1 U16189 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n17805), .ZN(
        n17804) );
  INV_X1 U16190 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18106) );
  NAND2_X1 U16191 ( .A1(n13063), .A2(n13060), .ZN(n13064) );
  NAND2_X1 U16192 ( .A1(n13063), .A2(n13062), .ZN(n13061) );
  NAND2_X1 U16193 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17775), .ZN(
        n17774) );
  INV_X1 U16194 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18034) );
  INV_X1 U16195 ( .A(n17539), .ZN(n17575) );
  NAND2_X1 U16196 ( .A1(n17926), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17555) );
  NAND3_X1 U16197 ( .A1(n17521), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16340) );
  INV_X1 U16198 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18815) );
  NAND3_X1 U16199 ( .A1(n18815), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n13074) );
  NAND2_X1 U16200 ( .A1(n17521), .A2(n13072), .ZN(n16301) );
  OAI21_X1 U16201 ( .B1(n21009), .B2(n16301), .A(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13065) );
  OAI21_X1 U16202 ( .B1(n16340), .B2(n13074), .A(n13065), .ZN(n16333) );
  INV_X1 U16203 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18813) );
  NOR2_X1 U16204 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18866) );
  INV_X1 U16205 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18865) );
  NAND2_X1 U16206 ( .A1(n18865), .A2(n18808), .ZN(n16433) );
  INV_X1 U16207 ( .A(n16433), .ZN(n13066) );
  NOR2_X1 U16208 ( .A1(n18866), .A2(n13066), .ZN(n18848) );
  INV_X1 U16209 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18852) );
  NOR2_X1 U16210 ( .A1(n18813), .A2(n18852), .ZN(n17829) );
  INV_X1 U16211 ( .A(n17829), .ZN(n17845) );
  INV_X1 U16212 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16485) );
  NAND2_X1 U16213 ( .A1(n17812), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17800) );
  NAND4_X1 U16214 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A4(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17741) );
  NOR2_X1 U16215 ( .A1(n17741), .A2(n16702), .ZN(n16672) );
  NAND2_X1 U16216 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17715) );
  NAND2_X1 U16217 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17680) );
  NAND2_X1 U16218 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17641) );
  NAND2_X1 U16219 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17629), .ZN(
        n17606) );
  NAND2_X1 U16220 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17607) );
  NAND2_X1 U16221 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17562) );
  INV_X1 U16222 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17532) );
  INV_X1 U16223 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17512) );
  INV_X1 U16224 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17870) );
  NAND2_X1 U16225 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16321), .ZN(
        n13067) );
  XOR2_X2 U16226 ( .A(n16485), .B(n13067), .Z(n16758) );
  INV_X1 U16227 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18792) );
  NOR2_X1 U16228 ( .A1(n18792), .A2(n18193), .ZN(n16330) );
  NAND2_X1 U16229 ( .A1(n20757), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18721) );
  NOR2_X1 U16230 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18857) );
  AOI21_X1 U16231 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n18857), .ZN(n18718) );
  OR2_X1 U16232 ( .A1(n18828), .A2(n18718), .ZN(n18211) );
  NAND3_X1 U16233 ( .A1(n18865), .A2(n18808), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18359) );
  OR2_X1 U16234 ( .A1(n13069), .A2(n17714), .ZN(n16308) );
  XNOR2_X1 U16235 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13070) );
  NOR2_X1 U16236 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17665), .ZN(
        n16323) );
  NOR2_X1 U16237 ( .A1(n17870), .A2(n17511), .ZN(n16471) );
  NAND2_X1 U16238 ( .A1(n16471), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16475) );
  NOR2_X1 U16239 ( .A1(n16475), .A2(n17512), .ZN(n16474) );
  NAND2_X1 U16240 ( .A1(n18593), .A2(n13069), .ZN(n16311) );
  OAI211_X1 U16241 ( .C1(n16474), .C2(n18721), .A(n17877), .B(n16311), .ZN(
        n16313) );
  NOR2_X1 U16242 ( .A1(n16323), .A2(n16313), .ZN(n16307) );
  OAI22_X1 U16243 ( .A1(n16308), .A2(n13070), .B1(n16307), .B2(n16485), .ZN(
        n13071) );
  AOI211_X1 U16244 ( .C1(n9758), .C2(n16758), .A(n16330), .B(n13071), .ZN(
        n13079) );
  INV_X1 U16245 ( .A(n13072), .ZN(n16304) );
  INV_X1 U16246 ( .A(n17885), .ZN(n17895) );
  INV_X1 U16247 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17576) );
  NAND2_X1 U16248 ( .A1(n17539), .A2(n17940), .ZN(n17924) );
  NOR2_X1 U16249 ( .A1(n17576), .A2(n17924), .ZN(n17556) );
  NAND2_X1 U16250 ( .A1(n17895), .A2(n17556), .ZN(n17887) );
  NOR2_X1 U16251 ( .A1(n16304), .A2(n17887), .ZN(n15693) );
  NAND2_X1 U16252 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15693), .ZN(
        n13076) );
  INV_X1 U16253 ( .A(n13074), .ZN(n16332) );
  NAND2_X1 U16254 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n13075) );
  NOR2_X1 U16255 ( .A1(n13075), .A2(n17887), .ZN(n16341) );
  AOI22_X1 U16256 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n13076), .B1(
        n16332), .B2(n16341), .ZN(n16336) );
  INV_X1 U16257 ( .A(n16336), .ZN(n13077) );
  NAND2_X1 U16258 ( .A1(n13077), .A2(n17784), .ZN(n13078) );
  NOR4_X1 U16259 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13087) );
  NOR4_X1 U16260 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(
        P1_ADDRESS_REG_17__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n13086) );
  NOR4_X1 U16261 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13085) );
  NOR4_X1 U16262 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_8__SCAN_IN), .ZN(n13084) );
  AND4_X1 U16263 ( .A1(n13087), .A2(n13086), .A3(n13085), .A4(n13084), .ZN(
        n13093) );
  NOR4_X1 U16264 ( .A1(P1_ADDRESS_REG_2__SCAN_IN), .A2(
        P1_ADDRESS_REG_1__SCAN_IN), .A3(P1_ADDRESS_REG_28__SCAN_IN), .A4(
        P1_ADDRESS_REG_27__SCAN_IN), .ZN(n13091) );
  NOR4_X1 U16265 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(
        P1_ADDRESS_REG_21__SCAN_IN), .A3(P1_ADDRESS_REG_20__SCAN_IN), .A4(
        P1_ADDRESS_REG_19__SCAN_IN), .ZN(n13090) );
  NOR4_X1 U16266 ( .A1(P1_ADDRESS_REG_26__SCAN_IN), .A2(
        P1_ADDRESS_REG_25__SCAN_IN), .A3(P1_ADDRESS_REG_24__SCAN_IN), .A4(
        P1_ADDRESS_REG_23__SCAN_IN), .ZN(n13089) );
  INV_X1 U16267 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n13088) );
  AND4_X1 U16268 ( .A1(n13091), .A2(n13090), .A3(n13089), .A4(n13088), .ZN(
        n13092) );
  NAND2_X1 U16269 ( .A1(n13093), .A2(n13092), .ZN(n13094) );
  AND2_X2 U16270 ( .A1(n13094), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20107)
         );
  INV_X1 U16271 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20714) );
  NOR3_X1 U16272 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20714), .ZN(n13096) );
  NOR4_X1 U16273 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13095) );
  NAND4_X1 U16274 ( .A1(n20107), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13096), .A4(
        n13095), .ZN(U214) );
  NOR2_X1 U16275 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13098) );
  NOR4_X1 U16276 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13097) );
  NAND4_X1 U16277 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13098), .A4(n13097), .ZN(n13099) );
  NOR2_X1 U16278 ( .A1(n13225), .A2(n13099), .ZN(n16353) );
  NAND2_X1 U16279 ( .A1(n16353), .A2(U214), .ZN(U212) );
  NOR2_X1 U16280 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13099), .ZN(n16423)
         );
  NAND2_X1 U16281 ( .A1(n18915), .A2(n19019), .ZN(n16073) );
  AOI211_X1 U16282 ( .C1(n16166), .C2(n13100), .A(n18931), .B(n16073), .ZN(
        n13115) );
  INV_X1 U16283 ( .A(n16166), .ZN(n13102) );
  NAND2_X1 U16284 ( .A1(n19005), .A2(n18915), .ZN(n19040) );
  AOI22_X1 U16285 ( .A1(P2_EBX_REG_15__SCAN_IN), .A2(n18957), .B1(
        P2_REIP_REG_15__SCAN_IN), .B2(n19028), .ZN(n13101) );
  OAI211_X1 U16286 ( .C1(n13102), .C2(n19040), .A(n13101), .B(n19012), .ZN(
        n13114) );
  OAI22_X1 U16287 ( .A1(n13103), .A2(n19014), .B1(n19041), .B2(n20775), .ZN(
        n13113) );
  NAND2_X1 U16288 ( .A1(n13104), .A2(n13105), .ZN(n13106) );
  AND2_X1 U16289 ( .A1(n13940), .A2(n13106), .ZN(n16167) );
  INV_X1 U16290 ( .A(n16167), .ZN(n13111) );
  INV_X1 U16291 ( .A(n13107), .ZN(n15466) );
  NAND2_X1 U16292 ( .A1(n13108), .A2(n15466), .ZN(n13110) );
  NAND2_X1 U16293 ( .A1(n13110), .A2(n13109), .ZN(n19053) );
  OAI22_X1 U16294 ( .A1(n13111), .A2(n19037), .B1(n19053), .B2(n19026), .ZN(
        n13112) );
  AOI211_X1 U16295 ( .C1(n15213), .C2(n13116), .A(n18965), .B(n16073), .ZN(
        n13128) );
  OR2_X1 U16296 ( .A1(n13117), .A2(n9841), .ZN(n13118) );
  NAND2_X1 U16297 ( .A1(n13118), .A2(n16195), .ZN(n19061) );
  AOI22_X1 U16298 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n18957), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(n19028), .ZN(n13119) );
  OAI211_X1 U16299 ( .C1(n19061), .C2(n19026), .A(n13119), .B(n19012), .ZN(
        n13127) );
  INV_X1 U16300 ( .A(n13120), .ZN(n13121) );
  OAI22_X1 U16301 ( .A1(n13121), .A2(n19014), .B1(n19041), .B2(n15211), .ZN(
        n13126) );
  NAND2_X1 U16302 ( .A1(n13676), .A2(n13122), .ZN(n13123) );
  NAND2_X1 U16303 ( .A1(n9782), .A2(n13123), .ZN(n15497) );
  INV_X1 U16304 ( .A(n15213), .ZN(n13124) );
  OAI22_X1 U16305 ( .A1(n15497), .A2(n19037), .B1(n19040), .B2(n13124), .ZN(
        n13125) );
  OR4_X1 U16306 ( .A1(n13128), .A2(n13127), .A3(n13126), .A4(n13125), .ZN(
        P2_U2844) );
  NOR2_X1 U16307 ( .A1(n12221), .A2(n18880), .ZN(n19115) );
  NAND2_X1 U16308 ( .A1(n19115), .A2(n16273), .ZN(n14877) );
  INV_X1 U16309 ( .A(n14877), .ZN(n19044) );
  INV_X1 U16310 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13131) );
  INV_X1 U16311 ( .A(n13134), .ZN(n13130) );
  NOR2_X1 U16312 ( .A1(n19636), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n13132) );
  INV_X1 U16313 ( .A(n13132), .ZN(n13129) );
  OAI211_X1 U16314 ( .C1(n19044), .C2(n13131), .A(n13130), .B(n13129), .ZN(
        P2_U2814) );
  OAI21_X1 U16315 ( .B1(n13132), .B2(P2_READREQUEST_REG_SCAN_IN), .A(n19863), 
        .ZN(n13133) );
  OAI21_X1 U16316 ( .B1(n19873), .B2(n19863), .A(n13133), .ZN(P2_U3612) );
  OAI21_X1 U16317 ( .B1(n19869), .B2(n19867), .A(n13134), .ZN(n13244) );
  AOI22_X1 U16318 ( .A1(n13178), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n13244), 
        .B2(P2_UWORD_REG_5__SCAN_IN), .ZN(n13135) );
  NAND3_X1 U16319 ( .A1(n13134), .A2(n9743), .A3(n19867), .ZN(n13145) );
  OAI22_X1 U16320 ( .A1(n13225), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13828), .ZN(n19239) );
  INV_X1 U16321 ( .A(n19239), .ZN(n19075) );
  NAND2_X1 U16322 ( .A1(n19185), .A2(n19075), .ZN(n13242) );
  NAND2_X1 U16323 ( .A1(n13135), .A2(n13242), .ZN(P2_U2957) );
  AOI22_X1 U16324 ( .A1(P2_EAX_REG_27__SCAN_IN), .A2(n13178), .B1(n13244), 
        .B2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13137) );
  AOI22_X1 U16325 ( .A1(n13828), .A2(BUF1_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n13225), .ZN(n19060) );
  INV_X1 U16326 ( .A(n19060), .ZN(n13136) );
  NAND2_X1 U16327 ( .A1(n19185), .A2(n13136), .ZN(n13234) );
  NAND2_X1 U16328 ( .A1(n13137), .A2(n13234), .ZN(P2_U2963) );
  AOI22_X1 U16329 ( .A1(P2_EAX_REG_13__SCAN_IN), .A2(n13178), .B1(n13244), 
        .B2(P2_LWORD_REG_13__SCAN_IN), .ZN(n13139) );
  AOI22_X1 U16330 ( .A1(n13828), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n13830), .ZN(n19056) );
  INV_X1 U16331 ( .A(n19056), .ZN(n13138) );
  NAND2_X1 U16332 ( .A1(n19185), .A2(n13138), .ZN(n13140) );
  NAND2_X1 U16333 ( .A1(n13139), .A2(n13140), .ZN(P2_U2980) );
  AOI22_X1 U16334 ( .A1(P2_EAX_REG_29__SCAN_IN), .A2(n13178), .B1(n13244), 
        .B2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13141) );
  NAND2_X1 U16335 ( .A1(n13141), .A2(n13140), .ZN(P2_U2965) );
  INV_X1 U16336 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19165) );
  INV_X1 U16337 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16383) );
  INV_X1 U16338 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17489) );
  AOI22_X1 U16339 ( .A1(n13828), .A2(n16383), .B1(n17489), .B2(n13830), .ZN(
        n19068) );
  NAND2_X1 U16340 ( .A1(n19185), .A2(n19068), .ZN(n13144) );
  INV_X1 U16341 ( .A(n13244), .ZN(n13146) );
  NAND2_X1 U16342 ( .A1(n19187), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13142) );
  OAI211_X1 U16343 ( .C1(n19116), .C2(n19165), .A(n13144), .B(n13142), .ZN(
        P2_U2975) );
  INV_X1 U16344 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n19133) );
  NAND2_X1 U16345 ( .A1(n19187), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13143) );
  OAI211_X1 U16346 ( .C1(n19116), .C2(n19133), .A(n13144), .B(n13143), .ZN(
        P2_U2960) );
  INV_X1 U16347 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13148) );
  INV_X1 U16348 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13147) );
  AOI22_X1 U16349 ( .A1(n13828), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13830), .ZN(n19052) );
  OAI222_X1 U16350 ( .A1(n19116), .A2(n13148), .B1(n13147), .B2(n13146), .C1(
        n13145), .C2(n19052), .ZN(P2_U2982) );
  AOI22_X1 U16351 ( .A1(P2_EAX_REG_22__SCAN_IN), .A2(n13178), .B1(n19187), 
        .B2(P2_UWORD_REG_6__SCAN_IN), .ZN(n13150) );
  AOI22_X1 U16352 ( .A1(n13828), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n13225), .ZN(n19246) );
  INV_X1 U16353 ( .A(n19246), .ZN(n13149) );
  NAND2_X1 U16354 ( .A1(n19185), .A2(n13149), .ZN(n13168) );
  NAND2_X1 U16355 ( .A1(n13150), .A2(n13168), .ZN(P2_U2958) );
  AOI22_X1 U16356 ( .A1(P2_EAX_REG_26__SCAN_IN), .A2(n13178), .B1(n19187), 
        .B2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13152) );
  AOI22_X1 U16357 ( .A1(n13828), .A2(BUF1_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n13225), .ZN(n19063) );
  INV_X1 U16358 ( .A(n19063), .ZN(n13151) );
  NAND2_X1 U16359 ( .A1(n19185), .A2(n13151), .ZN(n13166) );
  NAND2_X1 U16360 ( .A1(n13152), .A2(n13166), .ZN(P2_U2962) );
  NOR3_X1 U16361 ( .A1(n13158), .A2(n13157), .A3(n13156), .ZN(n13161) );
  OAI21_X1 U16362 ( .B1(n13161), .B2(n13160), .A(n13159), .ZN(n13448) );
  AND2_X1 U16363 ( .A1(n13448), .A2(n13162), .ZN(n13194) );
  INV_X1 U16364 ( .A(n19884), .ZN(n13560) );
  NAND2_X1 U16365 ( .A1(n13194), .A2(n13560), .ZN(n13181) );
  NOR2_X2 U16366 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20547) );
  AND2_X1 U16367 ( .A1(n20547), .A2(n14146), .ZN(n13879) );
  AOI21_X1 U16368 ( .B1(n13181), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n13879), 
        .ZN(n13163) );
  NAND2_X1 U16369 ( .A1(n13567), .A2(n13163), .ZN(P1_U2801) );
  AOI22_X1 U16370 ( .A1(n13178), .A2(P2_EAX_REG_7__SCAN_IN), .B1(n19187), .B2(
        P2_LWORD_REG_7__SCAN_IN), .ZN(n13165) );
  AOI22_X1 U16371 ( .A1(n13828), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13830), .ZN(n19256) );
  INV_X1 U16372 ( .A(n19256), .ZN(n13164) );
  NAND2_X1 U16373 ( .A1(n19185), .A2(n13164), .ZN(n13230) );
  NAND2_X1 U16374 ( .A1(n13165), .A2(n13230), .ZN(P2_U2974) );
  AOI22_X1 U16375 ( .A1(n13178), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n19187), 
        .B2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13167) );
  NAND2_X1 U16376 ( .A1(n13167), .A2(n13166), .ZN(P2_U2977) );
  AOI22_X1 U16377 ( .A1(n13178), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n19187), .B2(
        P2_LWORD_REG_6__SCAN_IN), .ZN(n13169) );
  NAND2_X1 U16378 ( .A1(n13169), .A2(n13168), .ZN(P2_U2973) );
  AOI22_X1 U16379 ( .A1(n13178), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n19187), 
        .B2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13171) );
  AOI22_X1 U16380 ( .A1(n13828), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n13830), .ZN(n19058) );
  INV_X1 U16381 ( .A(n19058), .ZN(n13170) );
  NAND2_X1 U16382 ( .A1(n19185), .A2(n13170), .ZN(n13245) );
  NAND2_X1 U16383 ( .A1(n13171), .A2(n13245), .ZN(P2_U2979) );
  AOI22_X1 U16384 ( .A1(n13178), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n19187), .B2(
        P2_LWORD_REG_4__SCAN_IN), .ZN(n13173) );
  AOI22_X1 U16385 ( .A1(n13828), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n13225), .ZN(n19234) );
  INV_X1 U16386 ( .A(n19234), .ZN(n13172) );
  NAND2_X1 U16387 ( .A1(n19185), .A2(n13172), .ZN(n13238) );
  NAND2_X1 U16388 ( .A1(n13173), .A2(n13238), .ZN(P2_U2971) );
  AOI22_X1 U16389 ( .A1(n13178), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n19187), 
        .B2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13175) );
  AOI22_X1 U16390 ( .A1(n13828), .A2(BUF1_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n13830), .ZN(n19065) );
  INV_X1 U16391 ( .A(n19065), .ZN(n13174) );
  NAND2_X1 U16392 ( .A1(n19185), .A2(n13174), .ZN(n13240) );
  NAND2_X1 U16393 ( .A1(n13175), .A2(n13240), .ZN(P2_U2961) );
  AOI22_X1 U16394 ( .A1(n13178), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n19187), .B2(
        P2_LWORD_REG_1__SCAN_IN), .ZN(n13177) );
  AOI22_X1 U16395 ( .A1(n13828), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13830), .ZN(n14005) );
  INV_X1 U16396 ( .A(n14005), .ZN(n13176) );
  NAND2_X1 U16397 ( .A1(n19185), .A2(n13176), .ZN(n13179) );
  NAND2_X1 U16398 ( .A1(n13177), .A2(n13179), .ZN(P2_U2968) );
  AOI22_X1 U16399 ( .A1(n13178), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n19187), 
        .B2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13180) );
  NAND2_X1 U16400 ( .A1(n13180), .A2(n13179), .ZN(P2_U2953) );
  OAI21_X1 U16401 ( .B1(n13879), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n13734), 
        .ZN(n13183) );
  OAI21_X1 U16402 ( .B1(n11184), .B2(n14191), .A(n20716), .ZN(n13182) );
  NAND2_X1 U16403 ( .A1(n13183), .A2(n13182), .ZN(P1_U3487) );
  INV_X1 U16404 ( .A(n13212), .ZN(n13185) );
  NAND2_X1 U16405 ( .A1(n19027), .A2(n15557), .ZN(n13184) );
  NAND2_X1 U16406 ( .A1(n13185), .A2(n13184), .ZN(n13271) );
  INV_X1 U16407 ( .A(n13271), .ZN(n13190) );
  AOI21_X1 U16408 ( .B1(n15557), .B2(n13187), .A(n13186), .ZN(n13188) );
  INV_X1 U16409 ( .A(n13188), .ZN(n13272) );
  NAND2_X1 U16410 ( .A1(n19206), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13278) );
  OAI21_X1 U16411 ( .B1(n19197), .B2(n13272), .A(n13278), .ZN(n13189) );
  AOI21_X1 U16412 ( .B1(n16190), .B2(n13190), .A(n13189), .ZN(n13193) );
  OAI21_X1 U16413 ( .B1(n19190), .B2(n13191), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13192) );
  OAI211_X1 U16414 ( .C1(n16186), .C2(n19038), .A(n13193), .B(n13192), .ZN(
        P2_U3014) );
  OAI22_X1 U16415 ( .A1(n13496), .A2(n11184), .B1(n13153), .B2(n13194), .ZN(
        n19885) );
  NOR2_X1 U16416 ( .A1(n11184), .A2(n13381), .ZN(n13462) );
  OR2_X1 U16417 ( .A1(n13195), .A2(P1_STATE_REG_0__SCAN_IN), .ZN(n15746) );
  NAND2_X1 U16418 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20718) );
  INV_X1 U16419 ( .A(n20718), .ZN(n15745) );
  AOI21_X1 U16420 ( .B1(n13462), .B2(n15746), .A(n15745), .ZN(n20720) );
  NOR2_X1 U16421 ( .A1(n19885), .A2(n20720), .ZN(n15716) );
  OR2_X1 U16422 ( .A1(n15716), .A2(n19884), .ZN(n19891) );
  INV_X1 U16423 ( .A(n19891), .ZN(n13210) );
  INV_X1 U16424 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13209) );
  NOR2_X1 U16425 ( .A1(n13196), .A2(n11780), .ZN(n13466) );
  OR2_X1 U16426 ( .A1(n13466), .A2(n13400), .ZN(n13200) );
  INV_X1 U16427 ( .A(n13197), .ZN(n13199) );
  OR2_X1 U16428 ( .A1(n11168), .A2(n11167), .ZN(n13198) );
  AND2_X1 U16429 ( .A1(n13199), .A2(n13198), .ZN(n13389) );
  NAND2_X1 U16430 ( .A1(n13373), .A2(n13386), .ZN(n15713) );
  AND2_X1 U16431 ( .A1(n13466), .A2(n11184), .ZN(n13446) );
  INV_X1 U16432 ( .A(n13446), .ZN(n13203) );
  NAND2_X1 U16433 ( .A1(n13400), .A2(n13201), .ZN(n13202) );
  NAND3_X1 U16434 ( .A1(n15713), .A2(n13203), .A3(n13202), .ZN(n13205) );
  INV_X1 U16435 ( .A(n13448), .ZN(n13204) );
  AOI22_X1 U16436 ( .A1(n13436), .A2(n13205), .B1(n13162), .B2(n13204), .ZN(
        n13207) );
  AND2_X1 U16437 ( .A1(n13466), .A2(n13381), .ZN(n13384) );
  NAND2_X1 U16438 ( .A1(n13496), .A2(n13384), .ZN(n13206) );
  AOI21_X1 U16439 ( .B1(n13207), .B2(n13206), .A(n20148), .ZN(n15715) );
  NAND2_X1 U16440 ( .A1(n13210), .A2(n15715), .ZN(n13208) );
  OAI21_X1 U16441 ( .B1(n13210), .B2(n13209), .A(n13208), .ZN(P1_U3484) );
  INV_X1 U16442 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13219) );
  XNOR2_X1 U16443 ( .A(n14873), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13211) );
  XNOR2_X1 U16444 ( .A(n13212), .B(n13211), .ZN(n15560) );
  NOR2_X1 U16445 ( .A1(n19198), .A2(n15560), .ZN(n13218) );
  OAI21_X1 U16446 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13214), .A(
        n13213), .ZN(n15561) );
  INV_X1 U16447 ( .A(n15561), .ZN(n13215) );
  NOR2_X1 U16448 ( .A1(n19012), .A2(n14868), .ZN(n15562) );
  AOI21_X1 U16449 ( .B1(n16188), .B2(n13215), .A(n15562), .ZN(n13216) );
  OAI21_X1 U16450 ( .B1(n13219), .B2(n16194), .A(n13216), .ZN(n13217) );
  AOI211_X1 U16451 ( .C1(n16187), .C2(n13219), .A(n13218), .B(n13217), .ZN(
        n13220) );
  OAI21_X1 U16452 ( .B1(n13258), .B2(n16186), .A(n13220), .ZN(P2_U3013) );
  AOI22_X1 U16453 ( .A1(n13178), .A2(P2_EAX_REG_0__SCAN_IN), .B1(n19187), .B2(
        P2_LWORD_REG_0__SCAN_IN), .ZN(n13222) );
  AOI22_X1 U16454 ( .A1(n13828), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13225), .ZN(n19114) );
  INV_X1 U16455 ( .A(n19114), .ZN(n13221) );
  NAND2_X1 U16456 ( .A1(n19185), .A2(n13221), .ZN(n13232) );
  NAND2_X1 U16457 ( .A1(n13222), .A2(n13232), .ZN(P2_U2967) );
  AOI22_X1 U16458 ( .A1(n13178), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n19187), .B2(
        P2_LWORD_REG_2__SCAN_IN), .ZN(n13224) );
  AOI22_X1 U16459 ( .A1(n13828), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13225), .ZN(n19224) );
  INV_X1 U16460 ( .A(n19224), .ZN(n13223) );
  NAND2_X1 U16461 ( .A1(n19185), .A2(n13223), .ZN(n13236) );
  NAND2_X1 U16462 ( .A1(n13224), .A2(n13236), .ZN(P2_U2969) );
  AOI22_X1 U16463 ( .A1(n13178), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n19187), 
        .B2(P2_UWORD_REG_3__SCAN_IN), .ZN(n13227) );
  AOI22_X1 U16464 ( .A1(n13828), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13225), .ZN(n19229) );
  INV_X1 U16465 ( .A(n19229), .ZN(n13226) );
  NAND2_X1 U16466 ( .A1(n19185), .A2(n13226), .ZN(n13228) );
  NAND2_X1 U16467 ( .A1(n13227), .A2(n13228), .ZN(P2_U2955) );
  AOI22_X1 U16468 ( .A1(n13178), .A2(P2_EAX_REG_3__SCAN_IN), .B1(n19187), .B2(
        P2_LWORD_REG_3__SCAN_IN), .ZN(n13229) );
  NAND2_X1 U16469 ( .A1(n13229), .A2(n13228), .ZN(P2_U2970) );
  AOI22_X1 U16470 ( .A1(n13178), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n13244), 
        .B2(P2_UWORD_REG_7__SCAN_IN), .ZN(n13231) );
  NAND2_X1 U16471 ( .A1(n13231), .A2(n13230), .ZN(P2_U2959) );
  AOI22_X1 U16472 ( .A1(P2_EAX_REG_16__SCAN_IN), .A2(n13178), .B1(n19187), 
        .B2(P2_UWORD_REG_0__SCAN_IN), .ZN(n13233) );
  NAND2_X1 U16473 ( .A1(n13233), .A2(n13232), .ZN(P2_U2952) );
  AOI22_X1 U16474 ( .A1(P2_EAX_REG_11__SCAN_IN), .A2(n13178), .B1(n19187), 
        .B2(P2_LWORD_REG_11__SCAN_IN), .ZN(n13235) );
  NAND2_X1 U16475 ( .A1(n13235), .A2(n13234), .ZN(P2_U2978) );
  AOI22_X1 U16476 ( .A1(P2_EAX_REG_18__SCAN_IN), .A2(n13178), .B1(n19187), 
        .B2(P2_UWORD_REG_2__SCAN_IN), .ZN(n13237) );
  NAND2_X1 U16477 ( .A1(n13237), .A2(n13236), .ZN(P2_U2954) );
  AOI22_X1 U16478 ( .A1(P2_EAX_REG_20__SCAN_IN), .A2(n13178), .B1(n19187), 
        .B2(P2_UWORD_REG_4__SCAN_IN), .ZN(n13239) );
  NAND2_X1 U16479 ( .A1(n13239), .A2(n13238), .ZN(P2_U2956) );
  AOI22_X1 U16480 ( .A1(P2_EAX_REG_9__SCAN_IN), .A2(n13178), .B1(n19187), .B2(
        P2_LWORD_REG_9__SCAN_IN), .ZN(n13241) );
  NAND2_X1 U16481 ( .A1(n13241), .A2(n13240), .ZN(P2_U2976) );
  AOI22_X1 U16482 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n13178), .B1(n19187), .B2(
        P2_LWORD_REG_5__SCAN_IN), .ZN(n13243) );
  NAND2_X1 U16483 ( .A1(n13243), .A2(n13242), .ZN(P2_U2972) );
  AOI22_X1 U16484 ( .A1(P2_EAX_REG_28__SCAN_IN), .A2(n13178), .B1(n13244), 
        .B2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13246) );
  NAND2_X1 U16485 ( .A1(n13246), .A2(n13245), .ZN(P2_U2964) );
  NAND2_X1 U16486 ( .A1(n9743), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13247) );
  AND4_X1 U16487 ( .A1(n19245), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13247), 
        .A4(n19385), .ZN(n13248) );
  INV_X1 U16488 ( .A(n16276), .ZN(n16272) );
  INV_X1 U16489 ( .A(n15581), .ZN(n16275) );
  NAND2_X1 U16490 ( .A1(n16272), .A2(n16275), .ZN(n14092) );
  INV_X1 U16491 ( .A(n12263), .ZN(n15584) );
  NAND2_X1 U16492 ( .A1(n14092), .A2(n15584), .ZN(n13250) );
  MUX2_X1 U16493 ( .A(n19038), .B(n19032), .S(n13257), .Z(n13252) );
  OAI21_X1 U16494 ( .B1(n19846), .B2(n14966), .A(n13252), .ZN(P2_U2887) );
  NAND2_X1 U16495 ( .A1(n13254), .A2(n13253), .ZN(n13255) );
  MUX2_X1 U16496 ( .A(n13259), .B(n13258), .S(n13251), .Z(n13260) );
  OAI21_X1 U16497 ( .B1(n19838), .B2(n14966), .A(n13260), .ZN(P2_U2886) );
  INV_X1 U16498 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13265) );
  INV_X1 U16499 ( .A(n13261), .ZN(n13263) );
  NAND2_X1 U16500 ( .A1(n13263), .A2(n13262), .ZN(n13288) );
  NAND3_X1 U16501 ( .A1(n16190), .A2(n13289), .A3(n13288), .ZN(n13264) );
  NAND2_X1 U16502 ( .A1(n19206), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n13295) );
  OAI211_X1 U16503 ( .C1(n13265), .C2(n16194), .A(n13264), .B(n13295), .ZN(
        n13269) );
  XNOR2_X1 U16504 ( .A(n13267), .B(n13266), .ZN(n13291) );
  OAI22_X1 U16505 ( .A1(n19205), .A2(n14854), .B1(n19197), .B2(n13291), .ZN(
        n13268) );
  AOI211_X1 U16506 ( .C1(n15591), .C2(n19201), .A(n13269), .B(n13268), .ZN(
        n13270) );
  INV_X1 U16507 ( .A(n13270), .ZN(P2_U3012) );
  OAI22_X1 U16508 ( .A1(n19215), .A2(n13272), .B1(n16227), .B2(n13271), .ZN(
        n13281) );
  INV_X1 U16509 ( .A(n13273), .ZN(n15564) );
  NOR2_X1 U16510 ( .A1(n13275), .A2(n13274), .ZN(n13276) );
  NOR2_X1 U16511 ( .A1(n13277), .A2(n13276), .ZN(n19109) );
  AOI22_X1 U16512 ( .A1(n15564), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19208), .B2(n19109), .ZN(n13279) );
  OAI211_X1 U16513 ( .C1(n15520), .C2(n19038), .A(n13279), .B(n13278), .ZN(
        n13280) );
  AOI211_X1 U16514 ( .C1(n15557), .C2(n15426), .A(n13281), .B(n13280), .ZN(
        n13282) );
  INV_X1 U16515 ( .A(n13282), .ZN(P2_U3046) );
  NAND2_X1 U16516 ( .A1(n13284), .A2(n13283), .ZN(n13287) );
  INV_X1 U16517 ( .A(n13285), .ZN(n13286) );
  NAND2_X1 U16518 ( .A1(n13287), .A2(n13286), .ZN(n19829) );
  INV_X1 U16519 ( .A(n19829), .ZN(n19076) );
  NAND3_X1 U16520 ( .A1(n19219), .A2(n13289), .A3(n13288), .ZN(n13290) );
  OAI21_X1 U16521 ( .B1(n19215), .B2(n13291), .A(n13290), .ZN(n13299) );
  INV_X1 U16522 ( .A(n13292), .ZN(n13293) );
  OR2_X1 U16523 ( .A1(n13294), .A2(n13293), .ZN(n13297) );
  AOI22_X1 U16524 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n15564), .B1(
        n15419), .B2(n13297), .ZN(n13296) );
  OAI211_X1 U16525 ( .C1(n15425), .C2(n13297), .A(n13296), .B(n13295), .ZN(
        n13298) );
  AOI211_X1 U16526 ( .C1(n15591), .C2(n19212), .A(n13299), .B(n13298), .ZN(
        n13300) );
  OAI21_X1 U16527 ( .B1(n19076), .B2(n16197), .A(n13300), .ZN(P2_U3044) );
  INV_X1 U16528 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n14857) );
  MUX2_X1 U16529 ( .A(n14857), .B(n11907), .S(n13251), .Z(n13303) );
  OAI21_X1 U16530 ( .B1(n19825), .B2(n14966), .A(n13303), .ZN(P2_U2885) );
  INV_X1 U16531 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n20752) );
  AND2_X1 U16532 ( .A1(n13162), .A2(n13751), .ZN(n15704) );
  NAND3_X1 U16533 ( .A1(n13496), .A2(n13560), .A3(n15704), .ZN(n13304) );
  OAI21_X1 U16534 ( .B1(n13567), .B2(n13751), .A(n13304), .ZN(n13305) );
  INV_X1 U16535 ( .A(n15746), .ZN(n15723) );
  NAND2_X1 U16536 ( .A1(n20023), .A2(n13748), .ZN(n20008) );
  NAND2_X1 U16537 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16064) );
  OR2_X1 U16538 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16064), .ZN(n20013) );
  INV_X2 U16539 ( .A(n20013), .ZN(n20719) );
  AOI22_X1 U16540 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13306) );
  OAI21_X1 U16541 ( .B1(n20752), .B2(n20008), .A(n13306), .ZN(P1_U2906) );
  AOI22_X1 U16542 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13307) );
  OAI21_X1 U16543 ( .B1(n14381), .B2(n20008), .A(n13307), .ZN(P1_U2912) );
  AOI22_X1 U16544 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13308) );
  OAI21_X1 U16545 ( .B1(n11681), .B2(n20008), .A(n13308), .ZN(P1_U2911) );
  AOI22_X1 U16546 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13309) );
  OAI21_X1 U16547 ( .B1(n14410), .B2(n20008), .A(n13309), .ZN(P1_U2918) );
  AOI22_X1 U16548 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13310) );
  OAI21_X1 U16549 ( .B1(n14394), .B2(n20008), .A(n13310), .ZN(P1_U2914) );
  INV_X1 U16550 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13312) );
  AOI22_X1 U16551 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13311) );
  OAI21_X1 U16552 ( .B1(n13312), .B2(n20008), .A(n13311), .ZN(P1_U2915) );
  INV_X1 U16553 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13314) );
  AOI22_X1 U16554 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13313) );
  OAI21_X1 U16555 ( .B1(n13314), .B2(n20008), .A(n13313), .ZN(P1_U2913) );
  INV_X1 U16556 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n13316) );
  AOI22_X1 U16557 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13315) );
  OAI21_X1 U16558 ( .B1(n13316), .B2(n20008), .A(n13315), .ZN(P1_U2907) );
  AOI22_X1 U16559 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13317) );
  OAI21_X1 U16560 ( .B1(n14366), .B2(n20008), .A(n13317), .ZN(P1_U2908) );
  AOI22_X1 U16561 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13318) );
  OAI21_X1 U16562 ( .B1(n11703), .B2(n20008), .A(n13318), .ZN(P1_U2909) );
  AOI22_X1 U16563 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13319) );
  OAI21_X1 U16564 ( .B1(n14374), .B2(n20008), .A(n13319), .ZN(P1_U2910) );
  INV_X1 U16565 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13321) );
  AOI22_X1 U16566 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13320) );
  OAI21_X1 U16567 ( .B1(n13321), .B2(n20008), .A(n13320), .ZN(P1_U2917) );
  AOI22_X1 U16568 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13322) );
  OAI21_X1 U16569 ( .B1(n11609), .B2(n20008), .A(n13322), .ZN(P1_U2916) );
  AND2_X1 U16570 ( .A1(n20721), .A2(n15745), .ZN(n13323) );
  AND2_X2 U16571 ( .A1(n13357), .A2(n20120), .ZN(n20056) );
  INV_X2 U16572 ( .A(n13357), .ZN(n20055) );
  AOI22_X1 U16573 ( .A1(n20056), .A2(P1_EAX_REG_21__SCAN_IN), .B1(n20055), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13326) );
  NAND2_X1 U16574 ( .A1(n13357), .A2(n13751), .ZN(n13358) );
  INV_X1 U16575 ( .A(n20107), .ZN(n20105) );
  NAND2_X1 U16576 ( .A1(n20105), .A2(DATAI_5_), .ZN(n13325) );
  NAND2_X1 U16577 ( .A1(n20107), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13324) );
  AND2_X1 U16578 ( .A1(n13325), .A2(n13324), .ZN(n20138) );
  INV_X1 U16579 ( .A(n20138), .ZN(n14398) );
  NAND2_X1 U16580 ( .A1(n20043), .A2(n14398), .ZN(n13620) );
  NAND2_X1 U16581 ( .A1(n13326), .A2(n13620), .ZN(P1_U2942) );
  AOI22_X1 U16582 ( .A1(n20056), .A2(P1_EAX_REG_16__SCAN_IN), .B1(n20055), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13329) );
  NAND2_X1 U16583 ( .A1(n20105), .A2(DATAI_0_), .ZN(n13328) );
  NAND2_X1 U16584 ( .A1(n20107), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13327) );
  AND2_X1 U16585 ( .A1(n13328), .A2(n13327), .ZN(n20103) );
  INV_X1 U16586 ( .A(n20103), .ZN(n14423) );
  NAND2_X1 U16587 ( .A1(n20043), .A2(n14423), .ZN(n13626) );
  NAND2_X1 U16588 ( .A1(n13329), .A2(n13626), .ZN(P1_U2937) );
  AOI22_X1 U16589 ( .A1(n20056), .A2(P1_EAX_REG_24__SCAN_IN), .B1(n20055), 
        .B2(P1_UWORD_REG_8__SCAN_IN), .ZN(n13332) );
  INV_X1 U16590 ( .A(DATAI_8_), .ZN(n13331) );
  NAND2_X1 U16591 ( .A1(n20107), .A2(BUF1_REG_8__SCAN_IN), .ZN(n13330) );
  OAI21_X1 U16592 ( .B1(n20107), .B2(n13331), .A(n13330), .ZN(n14384) );
  NAND2_X1 U16593 ( .A1(n20043), .A2(n14384), .ZN(n13349) );
  NAND2_X1 U16594 ( .A1(n13332), .A2(n13349), .ZN(P1_U2945) );
  AOI22_X1 U16595 ( .A1(n20056), .A2(P1_EAX_REG_4__SCAN_IN), .B1(n20055), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13335) );
  NAND2_X1 U16596 ( .A1(n20105), .A2(DATAI_4_), .ZN(n13334) );
  NAND2_X1 U16597 ( .A1(n20107), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13333) );
  AND2_X1 U16598 ( .A1(n13334), .A2(n13333), .ZN(n20134) );
  INV_X1 U16599 ( .A(n20134), .ZN(n14402) );
  NAND2_X1 U16600 ( .A1(n20043), .A2(n14402), .ZN(n13607) );
  NAND2_X1 U16601 ( .A1(n13335), .A2(n13607), .ZN(P1_U2956) );
  AOI22_X1 U16602 ( .A1(n20056), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n20055), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13338) );
  NAND2_X1 U16603 ( .A1(n20105), .A2(DATAI_1_), .ZN(n13337) );
  NAND2_X1 U16604 ( .A1(n20107), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13336) );
  AND2_X1 U16605 ( .A1(n13337), .A2(n13336), .ZN(n20119) );
  INV_X1 U16606 ( .A(n20119), .ZN(n14417) );
  NAND2_X1 U16607 ( .A1(n20043), .A2(n14417), .ZN(n13624) );
  NAND2_X1 U16608 ( .A1(n13338), .A2(n13624), .ZN(P1_U2938) );
  NAND2_X1 U16609 ( .A1(n16141), .A2(n13339), .ZN(n19074) );
  XNOR2_X1 U16610 ( .A(n13341), .B(n13340), .ZN(n19833) );
  XNOR2_X1 U16611 ( .A(n19838), .B(n19833), .ZN(n13342) );
  NAND2_X1 U16612 ( .A1(n19110), .A2(n19109), .ZN(n19108) );
  NAND2_X1 U16613 ( .A1(n13342), .A2(n19108), .ZN(n19078) );
  OAI21_X1 U16614 ( .B1(n13342), .B2(n19108), .A(n19078), .ZN(n13343) );
  NAND2_X1 U16615 ( .A1(n13343), .A2(n19107), .ZN(n13345) );
  INV_X1 U16616 ( .A(n19072), .ZN(n19105) );
  AOI22_X1 U16617 ( .A1(n19106), .A2(n19833), .B1(n19105), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n13344) );
  OAI211_X1 U16618 ( .C1(n14005), .C2(n19113), .A(n13345), .B(n13344), .ZN(
        P2_U2918) );
  INV_X1 U16619 ( .A(n20056), .ZN(n13359) );
  INV_X1 U16620 ( .A(DATAI_14_), .ZN(n13347) );
  NAND2_X1 U16621 ( .A1(n20107), .A2(BUF1_REG_14__SCAN_IN), .ZN(n13346) );
  OAI21_X1 U16622 ( .B1(n20107), .B2(n13347), .A(n13346), .ZN(n14186) );
  NAND2_X1 U16623 ( .A1(n20043), .A2(n14186), .ZN(n20057) );
  NAND2_X1 U16624 ( .A1(n20055), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13348) );
  OAI211_X1 U16625 ( .C1(n13359), .C2(n20752), .A(n20057), .B(n13348), .ZN(
        P1_U2951) );
  INV_X1 U16626 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n13351) );
  NAND2_X1 U16627 ( .A1(n20055), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n13350) );
  OAI211_X1 U16628 ( .C1(n13359), .C2(n13351), .A(n13350), .B(n13349), .ZN(
        P1_U2960) );
  INV_X1 U16629 ( .A(DATAI_12_), .ZN(n13353) );
  NAND2_X1 U16630 ( .A1(n20107), .A2(BUF1_REG_12__SCAN_IN), .ZN(n13352) );
  OAI21_X1 U16631 ( .B1(n20107), .B2(n13353), .A(n13352), .ZN(n14368) );
  NAND2_X1 U16632 ( .A1(n20043), .A2(n14368), .ZN(n20051) );
  NAND2_X1 U16633 ( .A1(n20055), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n13354) );
  OAI211_X1 U16634 ( .C1(n13359), .C2(n14366), .A(n20051), .B(n13354), .ZN(
        P1_U2949) );
  INV_X1 U16635 ( .A(DATAI_15_), .ZN(n13356) );
  INV_X1 U16636 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13355) );
  MUX2_X1 U16637 ( .A(n13356), .B(n13355), .S(n20107), .Z(n14074) );
  INV_X1 U16638 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n20014) );
  OAI222_X1 U16639 ( .A1(n13359), .A2(n11526), .B1(n13358), .B2(n14074), .C1(
        n13357), .C2(n20014), .ZN(P1_U2967) );
  NAND2_X1 U16640 ( .A1(n11249), .A2(n13360), .ZN(n13524) );
  OAI21_X1 U16641 ( .B1(n20721), .B2(n13520), .A(n13524), .ZN(n13361) );
  INV_X1 U16642 ( .A(n13361), .ZN(n13362) );
  NAND2_X1 U16643 ( .A1(n20061), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n20063) );
  XNOR2_X1 U16644 ( .A(n13521), .B(n13520), .ZN(n13364) );
  INV_X1 U16645 ( .A(n11780), .ZN(n13387) );
  OAI211_X1 U16646 ( .C1(n13364), .C2(n20721), .A(n13387), .B(n14185), .ZN(
        n13365) );
  INV_X1 U16647 ( .A(n13365), .ZN(n13366) );
  OAI21_X1 U16648 ( .B1(n13367), .B2(n20120), .A(n13366), .ZN(n13530) );
  XNOR2_X1 U16649 ( .A(n13529), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13508) );
  NAND2_X1 U16650 ( .A1(n13439), .A2(n20718), .ZN(n13368) );
  AOI22_X1 U16651 ( .A1(n13368), .A2(n13748), .B1(n13955), .B2(n15746), .ZN(
        n13369) );
  OAI21_X1 U16652 ( .B1(n11159), .B2(n13369), .A(n13496), .ZN(n13372) );
  AOI21_X1 U16653 ( .B1(n13751), .B2(n15746), .A(n15745), .ZN(n13370) );
  NAND2_X1 U16654 ( .A1(n13448), .A2(n13370), .ZN(n13371) );
  MUX2_X1 U16655 ( .A(n13372), .B(n13371), .S(n13445), .Z(n13378) );
  INV_X1 U16656 ( .A(n13162), .ZN(n13375) );
  NAND2_X1 U16657 ( .A1(n13373), .A2(n13394), .ZN(n13374) );
  NAND2_X1 U16658 ( .A1(n13375), .A2(n13374), .ZN(n13443) );
  AND2_X1 U16659 ( .A1(n13376), .A2(n13443), .ZN(n13377) );
  NAND2_X1 U16660 ( .A1(n13378), .A2(n13377), .ZN(n13379) );
  AND2_X1 U16661 ( .A1(n13405), .A2(n11167), .ZN(n13380) );
  NOR2_X1 U16662 ( .A1(n13380), .A2(n13446), .ZN(n13382) );
  NAND2_X1 U16663 ( .A1(n13439), .A2(n13381), .ZN(n13440) );
  AND4_X1 U16664 ( .A1(n15713), .A2(n13447), .A3(n13382), .A4(n13440), .ZN(
        n13383) );
  NOR2_X2 U16665 ( .A1(n13408), .A2(n13383), .ZN(n20082) );
  NAND2_X1 U16666 ( .A1(n13385), .A2(n11184), .ZN(n13397) );
  OAI22_X1 U16667 ( .A1(n13702), .A2(n13387), .B1(n13386), .B2(n13746), .ZN(
        n13388) );
  INV_X1 U16668 ( .A(n13388), .ZN(n13396) );
  INV_X1 U16669 ( .A(n13389), .ZN(n13393) );
  AOI21_X1 U16670 ( .B1(n11180), .B2(n13445), .A(n20148), .ZN(n13390) );
  AOI21_X1 U16671 ( .B1(n13391), .B2(n13390), .A(n20120), .ZN(n13392) );
  AOI21_X1 U16672 ( .B1(n13393), .B2(n14191), .A(n13392), .ZN(n13395) );
  NAND4_X1 U16673 ( .A1(n13397), .A2(n13396), .A3(n13395), .A4(n13394), .ZN(
        n13430) );
  INV_X1 U16674 ( .A(n13398), .ZN(n13427) );
  OAI21_X1 U16675 ( .B1(n13427), .B2(n13400), .A(n13399), .ZN(n13401) );
  OR2_X1 U16676 ( .A1(n13430), .A2(n13401), .ZN(n13402) );
  NAND2_X1 U16677 ( .A1(n13403), .A2(n13402), .ZN(n13545) );
  NAND2_X1 U16678 ( .A1(n15755), .A2(n13545), .ZN(n13409) );
  NAND2_X1 U16679 ( .A1(n13403), .A2(n15704), .ZN(n20092) );
  INV_X1 U16680 ( .A(n20092), .ZN(n13404) );
  INV_X1 U16681 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20093) );
  NAND2_X1 U16682 ( .A1(n20093), .A2(n20092), .ZN(n13552) );
  NAND3_X1 U16683 ( .A1(n14580), .A2(n13553), .A3(n13552), .ZN(n13414) );
  AOI22_X1 U16684 ( .A1(n13153), .A2(n20120), .B1(n13405), .B2(n11222), .ZN(
        n13406) );
  XNOR2_X1 U16685 ( .A(n13407), .B(n14206), .ZN(n13888) );
  INV_X1 U16686 ( .A(n13888), .ZN(n13412) );
  NAND2_X1 U16687 ( .A1(n20066), .A2(n13408), .ZN(n20091) );
  NAND2_X1 U16688 ( .A1(n20093), .A2(n13409), .ZN(n20088) );
  AOI21_X1 U16689 ( .B1(n20091), .B2(n20088), .A(n13553), .ZN(n13411) );
  INV_X1 U16690 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20705) );
  NOR2_X1 U16691 ( .A1(n20066), .A2(n20705), .ZN(n13410) );
  AOI211_X1 U16692 ( .C1(n20085), .C2(n13412), .A(n13411), .B(n13410), .ZN(
        n13413) );
  OAI211_X1 U16693 ( .C1(n13508), .C2(n16025), .A(n13414), .B(n13413), .ZN(
        P1_U3030) );
  OR2_X1 U16694 ( .A1(n13417), .A2(n13416), .ZN(n13418) );
  NAND2_X1 U16695 ( .A1(n13415), .A2(n13418), .ZN(n19088) );
  NOR2_X1 U16696 ( .A1(n13421), .A2(n13420), .ZN(n13422) );
  OR2_X1 U16697 ( .A1(n13419), .A2(n13422), .ZN(n14837) );
  NOR2_X1 U16698 ( .A1(n14837), .A2(n13257), .ZN(n13423) );
  AOI21_X1 U16699 ( .B1(P2_EBX_REG_4__SCAN_IN), .B2(n13257), .A(n13423), .ZN(
        n13424) );
  OAI21_X1 U16700 ( .B1(n19088), .B2(n14966), .A(n13424), .ZN(P2_U2883) );
  NAND2_X1 U16701 ( .A1(n13427), .A2(n13426), .ZN(n13428) );
  NOR2_X1 U16702 ( .A1(n13428), .A2(n13439), .ZN(n13429) );
  NAND2_X1 U16703 ( .A1(n13447), .A2(n13429), .ZN(n13431) );
  OR2_X1 U16704 ( .A1(n13431), .A2(n13430), .ZN(n14144) );
  INV_X1 U16705 ( .A(n14144), .ZN(n14720) );
  XNOR2_X1 U16706 ( .A(n14718), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13433) );
  XNOR2_X1 U16707 ( .A(n10930), .B(n10921), .ZN(n13437) );
  NOR2_X1 U16708 ( .A1(n13462), .A2(n13437), .ZN(n13432) );
  AOI22_X1 U16709 ( .A1(n15704), .A2(n13433), .B1(n13466), .B2(n13432), .ZN(
        n13435) );
  NAND3_X1 U16710 ( .A1(n14720), .A2(n13470), .A3(n13437), .ZN(n13434) );
  OAI211_X1 U16711 ( .C1(n13425), .C2(n14720), .A(n13435), .B(n13434), .ZN(
        n13581) );
  NOR2_X1 U16712 ( .A1(n14146), .A2(n20093), .ZN(n14722) );
  INV_X1 U16713 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14572) );
  OAI22_X1 U16714 ( .A1(n14572), .A2(n13553), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14721) );
  INV_X1 U16715 ( .A(n14721), .ZN(n13438) );
  INV_X1 U16716 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20492) );
  AOI222_X1 U16717 ( .A1(n13581), .A2(n19883), .B1(n14722), .B2(n13438), .C1(
        n15731), .C2(n13437), .ZN(n13456) );
  OAI21_X1 U16718 ( .B1(n15704), .B2(n13439), .A(n15723), .ZN(n13441) );
  AOI21_X1 U16719 ( .B1(n13441), .B2(n13440), .A(n15745), .ZN(n13442) );
  NAND2_X1 U16720 ( .A1(n13496), .A2(n13442), .ZN(n13444) );
  OAI211_X1 U16721 ( .C1(n13746), .C2(n13445), .A(n13444), .B(n13443), .ZN(
        n13451) );
  NAND2_X1 U16722 ( .A1(n13496), .A2(n13446), .ZN(n13450) );
  INV_X1 U16723 ( .A(n13447), .ZN(n13590) );
  NAND3_X1 U16724 ( .A1(n13448), .A2(n13590), .A3(n20718), .ZN(n13449) );
  NAND2_X1 U16725 ( .A1(n13450), .A2(n13449), .ZN(n13561) );
  NOR2_X1 U16726 ( .A1(n13451), .A2(n13561), .ZN(n13452) );
  NOR2_X1 U16727 ( .A1(n20639), .A2(n16064), .ZN(n13595) );
  NAND2_X1 U16728 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n13595), .ZN(n13454) );
  OAI21_X1 U16729 ( .B1(n15699), .B2(n19884), .A(n13454), .ZN(n13482) );
  AOI21_X1 U16730 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20639), .A(n13482), 
        .ZN(n14151) );
  NAND2_X1 U16731 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n14151), .ZN(
        n13455) );
  OAI21_X1 U16732 ( .B1(n13456), .B2(n14151), .A(n13455), .ZN(P1_U3472) );
  INV_X1 U16733 ( .A(n20349), .ZN(n13668) );
  NAND2_X1 U16734 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13457) );
  INV_X1 U16735 ( .A(n13457), .ZN(n13458) );
  MUX2_X1 U16736 ( .A(n13458), .B(n13457), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13467) );
  INV_X1 U16737 ( .A(n13459), .ZN(n13464) );
  INV_X1 U16738 ( .A(n13460), .ZN(n13461) );
  MUX2_X1 U16739 ( .A(n13461), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n10930), .Z(n13463) );
  AOI21_X1 U16740 ( .B1(n13464), .B2(n13463), .A(n13462), .ZN(n13465) );
  AOI22_X1 U16741 ( .A1(n15704), .A2(n13467), .B1(n13466), .B2(n13465), .ZN(
        n13472) );
  INV_X1 U16742 ( .A(n10930), .ZN(n13469) );
  AOI211_X1 U16743 ( .C1(n13469), .C2(n11280), .A(n13468), .B(n11254), .ZN(
        n13473) );
  NAND3_X1 U16744 ( .A1(n14720), .A2(n13470), .A3(n13473), .ZN(n13471) );
  OAI211_X1 U16745 ( .C1(n13668), .C2(n14720), .A(n13472), .B(n13471), .ZN(
        n13582) );
  AOI22_X1 U16746 ( .A1(n19883), .A2(n13582), .B1(n15731), .B2(n13473), .ZN(
        n13475) );
  NAND2_X1 U16747 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n14151), .ZN(
        n13474) );
  OAI21_X1 U16748 ( .B1(n13475), .B2(n14151), .A(n13474), .ZN(P1_U3469) );
  MUX2_X1 U16749 ( .A(n10704), .B(n13478), .S(n13251), .Z(n13479) );
  OAI21_X1 U16750 ( .B1(n19818), .B2(n14966), .A(n13479), .ZN(P2_U2884) );
  INV_X1 U16751 ( .A(n14151), .ZN(n14726) );
  INV_X1 U16752 ( .A(n20244), .ZN(n20490) );
  OR2_X1 U16753 ( .A1(n13480), .A2(n20490), .ZN(n13481) );
  XNOR2_X1 U16754 ( .A(n13481), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n19952) );
  NAND4_X1 U16755 ( .A1(n13482), .A2(n19883), .A3(n13590), .A4(n19952), .ZN(
        n13483) );
  OAI21_X1 U16756 ( .B1(n13484), .B2(n14726), .A(n13483), .ZN(P1_U3468) );
  XOR2_X1 U16757 ( .A(n13415), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n13489)
         );
  OR2_X1 U16758 ( .A1(n13419), .A2(n13485), .ZN(n13486) );
  AND2_X1 U16759 ( .A1(n13486), .A2(n13513), .ZN(n19022) );
  INV_X1 U16760 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n19013) );
  NOR2_X1 U16761 ( .A1(n13251), .A2(n19013), .ZN(n13487) );
  AOI21_X1 U16762 ( .B1(n19022), .B2(n13251), .A(n13487), .ZN(n13488) );
  OAI21_X1 U16763 ( .B1(n13489), .B2(n14966), .A(n13488), .ZN(P2_U2882) );
  XNOR2_X1 U16764 ( .A(n13490), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13494) );
  OR2_X1 U16765 ( .A1(n13491), .A2(n13512), .ZN(n13492) );
  NAND2_X1 U16766 ( .A1(n13492), .A2(n13540), .ZN(n18993) );
  INV_X1 U16767 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n18992) );
  MUX2_X1 U16768 ( .A(n18993), .B(n18992), .S(n13257), .Z(n13493) );
  OAI21_X1 U16769 ( .B1(n13494), .B2(n14966), .A(n13493), .ZN(P2_U2880) );
  NOR2_X1 U16770 ( .A1(n15713), .A2(n19884), .ZN(n13495) );
  AND3_X1 U16771 ( .A1(n20639), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n13497) );
  OAI21_X1 U16772 ( .B1(n13499), .B2(n13498), .A(n13531), .ZN(n13886) );
  INV_X1 U16773 ( .A(n13886), .ZN(n13506) );
  NAND2_X1 U16774 ( .A1(n20581), .A2(n13500), .ZN(n20717) );
  NAND2_X1 U16775 ( .A1(n20717), .A2(n20639), .ZN(n13501) );
  NAND2_X1 U16776 ( .A1(n20639), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13503) );
  NAND2_X1 U16777 ( .A1(n20906), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13502) );
  NAND2_X1 U16778 ( .A1(n13503), .A2(n13502), .ZN(n20059) );
  INV_X2 U16779 ( .A(n20066), .ZN(n16053) );
  AOI22_X1 U16780 ( .A1(n20060), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n16053), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n13504) );
  OAI21_X1 U16781 ( .B1(n15978), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13504), .ZN(n13505) );
  AOI21_X1 U16782 ( .B1(n15975), .B2(n13506), .A(n13505), .ZN(n13507) );
  OAI21_X1 U16783 ( .B1(n13508), .B2(n15962), .A(n13507), .ZN(P1_U2998) );
  INV_X1 U16784 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13509) );
  NOR2_X1 U16785 ( .A1(n13415), .A2(n13509), .ZN(n13511) );
  INV_X1 U16786 ( .A(n13490), .ZN(n13510) );
  OAI211_X1 U16787 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n13511), .A(
        n13510), .B(n14941), .ZN(n13516) );
  AOI21_X1 U16788 ( .B1(n13514), .B2(n13513), .A(n13512), .ZN(n19008) );
  NAND2_X1 U16789 ( .A1(n13251), .A2(n19008), .ZN(n13515) );
  OAI211_X1 U16790 ( .C1(n13251), .C2(n18998), .A(n13516), .B(n13515), .ZN(
        P2_U2881) );
  NAND2_X1 U16791 ( .A1(n13664), .A2(n13904), .ZN(n13528) );
  INV_X1 U16792 ( .A(n13522), .ZN(n13519) );
  NAND2_X1 U16793 ( .A1(n13521), .A2(n13520), .ZN(n13518) );
  NAND2_X1 U16794 ( .A1(n13519), .A2(n13518), .ZN(n13644) );
  NAND3_X1 U16795 ( .A1(n13522), .A2(n13521), .A3(n13520), .ZN(n13523) );
  NAND2_X1 U16796 ( .A1(n13644), .A2(n13523), .ZN(n13526) );
  INV_X1 U16797 ( .A(n13524), .ZN(n13525) );
  AOI21_X1 U16798 ( .B1(n13955), .B2(n13526), .A(n13525), .ZN(n13527) );
  NAND2_X1 U16799 ( .A1(n13528), .A2(n13527), .ZN(n13638) );
  INV_X1 U16800 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13549) );
  XNOR2_X1 U16801 ( .A(n13638), .B(n13639), .ZN(n13559) );
  NAND2_X1 U16802 ( .A1(n13532), .A2(n13531), .ZN(n13533) );
  AND2_X1 U16803 ( .A1(n13534), .A2(n13533), .ZN(n19995) );
  NAND2_X1 U16804 ( .A1(n16053), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n13554) );
  NAND2_X1 U16805 ( .A1(n20060), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13535) );
  OAI211_X1 U16806 ( .C1(n15978), .C2(n19992), .A(n13554), .B(n13535), .ZN(
        n13536) );
  AOI21_X1 U16807 ( .B1(n15975), .B2(n19995), .A(n13536), .ZN(n13537) );
  OAI21_X1 U16808 ( .B1(n13559), .B2(n15962), .A(n13537), .ZN(P1_U2997) );
  XNOR2_X1 U16809 ( .A(n13538), .B(n13633), .ZN(n13544) );
  NAND2_X1 U16810 ( .A1(n13540), .A2(n13539), .ZN(n13541) );
  AND2_X1 U16811 ( .A1(n13629), .A2(n13541), .ZN(n16222) );
  NOR2_X1 U16812 ( .A1(n13251), .A2(n10707), .ZN(n13542) );
  AOI21_X1 U16813 ( .B1(n16222), .B2(n13251), .A(n13542), .ZN(n13543) );
  OAI21_X1 U16814 ( .B1(n13544), .B2(n14966), .A(n13543), .ZN(P2_U2879) );
  NAND2_X1 U16815 ( .A1(n13545), .A2(n20092), .ZN(n14574) );
  INV_X1 U16816 ( .A(n14574), .ZN(n14705) );
  OR2_X1 U16817 ( .A1(n13545), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13546) );
  NAND2_X1 U16818 ( .A1(n13546), .A2(n20091), .ZN(n13656) );
  OAI21_X1 U16819 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n14705), .A(
        n14577), .ZN(n13548) );
  INV_X1 U16820 ( .A(n15755), .ZN(n14709) );
  AND3_X1 U16821 ( .A1(n14709), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13547) );
  OAI21_X1 U16822 ( .B1(n13548), .B2(n13547), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13558) );
  OAI21_X1 U16823 ( .B1(n20093), .B2(n13553), .A(n13549), .ZN(n13797) );
  NOR2_X1 U16824 ( .A1(n15755), .A2(n13797), .ZN(n13657) );
  XNOR2_X1 U16825 ( .A(n13551), .B(n13550), .ZN(n19988) );
  NAND2_X1 U16826 ( .A1(n14574), .A2(n13552), .ZN(n16018) );
  OR3_X1 U16827 ( .A1(n13553), .A2(n16018), .A3(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13555) );
  OAI211_X1 U16828 ( .C1(n14712), .C2(n19988), .A(n13555), .B(n13554), .ZN(
        n13556) );
  NOR2_X1 U16829 ( .A1(n13657), .A2(n13556), .ZN(n13557) );
  OAI211_X1 U16830 ( .C1(n13559), .C2(n16025), .A(n13558), .B(n13557), .ZN(
        P1_U3029) );
  NAND2_X1 U16831 ( .A1(n13751), .A2(n20718), .ZN(n13566) );
  NAND2_X1 U16832 ( .A1(n13561), .A2(n13560), .ZN(n13565) );
  OR2_X1 U16833 ( .A1(n13563), .A2(n13562), .ZN(n13564) );
  OAI211_X4 U16834 ( .C1(n13567), .C2(n13566), .A(n13565), .B(n13564), .ZN(
        n14409) );
  NAND2_X1 U16835 ( .A1(n11168), .A2(n13568), .ZN(n13569) );
  OAI222_X1 U16836 ( .A1(n13886), .A2(n14431), .B1(n14075), .B2(n20119), .C1(
        n14409), .C2(n11362), .ZN(P1_U2903) );
  OAI21_X1 U16837 ( .B1(n13572), .B2(n13571), .A(n13570), .ZN(n20068) );
  OAI222_X1 U16838 ( .A1(n20068), .A2(n14431), .B1(n14075), .B2(n20103), .C1(
        n14409), .C2(n11353), .ZN(P1_U2904) );
  OAI21_X1 U16839 ( .B1(n13575), .B2(n13574), .A(n13573), .ZN(n13648) );
  NAND2_X1 U16840 ( .A1(n20105), .A2(DATAI_3_), .ZN(n13577) );
  NAND2_X1 U16841 ( .A1(n20107), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13576) );
  AND2_X1 U16842 ( .A1(n13577), .A2(n13576), .ZN(n20129) );
  OAI222_X1 U16843 ( .A1(n13648), .A2(n14431), .B1(n14075), .B2(n20129), .C1(
        n14409), .C2(n11373), .ZN(P1_U2901) );
  INV_X1 U16844 ( .A(n19995), .ZN(n13885) );
  NAND2_X1 U16845 ( .A1(n20105), .A2(DATAI_2_), .ZN(n13579) );
  NAND2_X1 U16846 ( .A1(n20107), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13578) );
  AND2_X1 U16847 ( .A1(n13579), .A2(n13578), .ZN(n20124) );
  OAI222_X1 U16848 ( .A1(n13885), .A2(n14431), .B1(n14075), .B2(n20124), .C1(
        n13580), .C2(n14409), .ZN(P1_U2902) );
  NOR2_X1 U16849 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n14146), .ZN(n13586) );
  MUX2_X1 U16850 ( .A(n13581), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15699), .Z(n15698) );
  AOI22_X1 U16851 ( .A1(n13586), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n14146), .B2(n15698), .ZN(n13584) );
  MUX2_X1 U16852 ( .A(n13582), .B(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15699), .Z(n15712) );
  AOI22_X1 U16853 ( .A1(n13586), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n14146), .B2(n15712), .ZN(n13583) );
  NOR2_X1 U16854 ( .A1(n13584), .A2(n13583), .ZN(n15722) );
  INV_X1 U16855 ( .A(n10928), .ZN(n13585) );
  NAND2_X1 U16856 ( .A1(n15722), .A2(n13585), .ZN(n13594) );
  NAND2_X1 U16857 ( .A1(n15699), .A2(n14146), .ZN(n13588) );
  INV_X1 U16858 ( .A(n13586), .ZN(n13587) );
  NAND2_X1 U16859 ( .A1(n13588), .A2(n13587), .ZN(n13589) );
  NAND2_X1 U16860 ( .A1(n13589), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n13592) );
  NAND3_X1 U16861 ( .A1(n19952), .A2(n13590), .A3(n14146), .ZN(n13591) );
  NAND2_X1 U16862 ( .A1(n13592), .A2(n13591), .ZN(n15721) );
  INV_X1 U16863 ( .A(n15721), .ZN(n13593) );
  NAND2_X1 U16864 ( .A1(n13594), .A2(n13593), .ZN(n13598) );
  OAI21_X1 U16865 ( .B1(n13598), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13595), .ZN(
        n13597) );
  NOR2_X1 U16866 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20722) );
  INV_X1 U16867 ( .A(n20722), .ZN(n13596) );
  NOR2_X1 U16868 ( .A1(n13598), .A2(n16064), .ZN(n15733) );
  NAND2_X1 U16869 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20492), .ZN(n13663) );
  INV_X1 U16870 ( .A(n13663), .ZN(n13599) );
  OAI22_X1 U16871 ( .A1(n13363), .A2(n20581), .B1(n11351), .B2(n13599), .ZN(
        n13600) );
  OAI21_X1 U16872 ( .B1(n15733), .B2(n13600), .A(n13689), .ZN(n13601) );
  OAI21_X1 U16873 ( .B1(n20517), .B2(n13689), .A(n13601), .ZN(P1_U3478) );
  AOI22_X1 U16874 ( .A1(n20056), .A2(P1_EAX_REG_7__SCAN_IN), .B1(n20055), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n13604) );
  NAND2_X1 U16875 ( .A1(n20105), .A2(DATAI_7_), .ZN(n13603) );
  NAND2_X1 U16876 ( .A1(n20107), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13602) );
  AND2_X1 U16877 ( .A1(n13603), .A2(n13602), .ZN(n20147) );
  INV_X1 U16878 ( .A(n20147), .ZN(n14388) );
  NAND2_X1 U16879 ( .A1(n20043), .A2(n14388), .ZN(n13613) );
  NAND2_X1 U16880 ( .A1(n13604), .A2(n13613), .ZN(P1_U2959) );
  AOI22_X1 U16881 ( .A1(n20056), .A2(P1_EAX_REG_18__SCAN_IN), .B1(n20055), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13606) );
  INV_X1 U16882 ( .A(n20124), .ZN(n13605) );
  NAND2_X1 U16883 ( .A1(n20043), .A2(n13605), .ZN(n13616) );
  NAND2_X1 U16884 ( .A1(n13606), .A2(n13616), .ZN(P1_U2939) );
  AOI22_X1 U16885 ( .A1(n20056), .A2(P1_EAX_REG_20__SCAN_IN), .B1(n20055), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13608) );
  NAND2_X1 U16886 ( .A1(n13608), .A2(n13607), .ZN(P1_U2941) );
  AOI22_X1 U16887 ( .A1(n20056), .A2(P1_EAX_REG_22__SCAN_IN), .B1(n20055), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13612) );
  NAND2_X1 U16888 ( .A1(n20105), .A2(DATAI_6_), .ZN(n13610) );
  NAND2_X1 U16889 ( .A1(n20107), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13609) );
  AND2_X1 U16890 ( .A1(n13610), .A2(n13609), .ZN(n20143) );
  INV_X1 U16891 ( .A(n20143), .ZN(n13611) );
  NAND2_X1 U16892 ( .A1(n20043), .A2(n13611), .ZN(n13622) );
  NAND2_X1 U16893 ( .A1(n13612), .A2(n13622), .ZN(P1_U2943) );
  AOI22_X1 U16894 ( .A1(n20056), .A2(P1_EAX_REG_23__SCAN_IN), .B1(n20055), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13614) );
  NAND2_X1 U16895 ( .A1(n13614), .A2(n13613), .ZN(P1_U2944) );
  AOI22_X1 U16896 ( .A1(n20056), .A2(P1_EAX_REG_19__SCAN_IN), .B1(n20055), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13615) );
  INV_X1 U16897 ( .A(n20129), .ZN(n14405) );
  NAND2_X1 U16898 ( .A1(n20043), .A2(n14405), .ZN(n13618) );
  NAND2_X1 U16899 ( .A1(n13615), .A2(n13618), .ZN(P1_U2940) );
  AOI22_X1 U16900 ( .A1(n20056), .A2(P1_EAX_REG_2__SCAN_IN), .B1(n20055), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n13617) );
  NAND2_X1 U16901 ( .A1(n13617), .A2(n13616), .ZN(P1_U2954) );
  AOI22_X1 U16902 ( .A1(n20056), .A2(P1_EAX_REG_3__SCAN_IN), .B1(n20055), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13619) );
  NAND2_X1 U16903 ( .A1(n13619), .A2(n13618), .ZN(P1_U2955) );
  AOI22_X1 U16904 ( .A1(n20056), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n20055), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n13621) );
  NAND2_X1 U16905 ( .A1(n13621), .A2(n13620), .ZN(P1_U2957) );
  AOI22_X1 U16906 ( .A1(n20056), .A2(P1_EAX_REG_6__SCAN_IN), .B1(n20055), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n13623) );
  NAND2_X1 U16907 ( .A1(n13623), .A2(n13622), .ZN(P1_U2958) );
  AOI22_X1 U16908 ( .A1(n20056), .A2(P1_EAX_REG_1__SCAN_IN), .B1(n20055), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13625) );
  NAND2_X1 U16909 ( .A1(n13625), .A2(n13624), .ZN(P1_U2953) );
  AOI22_X1 U16910 ( .A1(n20056), .A2(P1_EAX_REG_0__SCAN_IN), .B1(n20055), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13627) );
  NAND2_X1 U16911 ( .A1(n13627), .A2(n13626), .ZN(P1_U2952) );
  AOI21_X1 U16912 ( .B1(n13630), .B2(n13629), .A(n13628), .ZN(n13631) );
  INV_X1 U16913 ( .A(n13631), .ZN(n18982) );
  OAI21_X1 U16914 ( .B1(n13538), .B2(n13633), .A(n13632), .ZN(n13635) );
  NAND3_X1 U16915 ( .A1(n13635), .A2(n14941), .A3(n13634), .ZN(n13637) );
  NAND2_X1 U16916 ( .A1(n13257), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n13636) );
  OAI211_X1 U16917 ( .C1(n18982), .C2(n13257), .A(n13637), .B(n13636), .ZN(
        P2_U2878) );
  NAND2_X1 U16918 ( .A1(n13639), .A2(n13638), .ZN(n13642) );
  NAND2_X1 U16919 ( .A1(n13640), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13641) );
  OR2_X1 U16920 ( .A1(n20096), .A2(n13643), .ZN(n13647) );
  NAND2_X1 U16921 ( .A1(n13644), .A2(n13645), .ZN(n13807) );
  OAI211_X1 U16922 ( .C1(n13645), .C2(n13644), .A(n13807), .B(n13955), .ZN(
        n13646) );
  NAND2_X1 U16923 ( .A1(n13647), .A2(n13646), .ZN(n13710) );
  XNOR2_X1 U16924 ( .A(n13711), .B(n13710), .ZN(n13662) );
  INV_X1 U16925 ( .A(n13648), .ZN(n19978) );
  NAND2_X1 U16926 ( .A1(n16053), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n13655) );
  NAND2_X1 U16927 ( .A1(n20060), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13649) );
  OAI211_X1 U16928 ( .C1(n15978), .C2(n19976), .A(n13655), .B(n13649), .ZN(
        n13650) );
  AOI21_X1 U16929 ( .B1(n19978), .B2(n15975), .A(n13650), .ZN(n13651) );
  OAI21_X1 U16930 ( .B1(n13662), .B2(n15962), .A(n13651), .ZN(P1_U2996) );
  NAND2_X1 U16931 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n14022) );
  OAI21_X1 U16932 ( .B1(n14022), .B2(n16018), .A(n15755), .ZN(n14663) );
  NAND2_X1 U16933 ( .A1(n13653), .A2(n13652), .ZN(n13654) );
  NAND2_X1 U16934 ( .A1(n13850), .A2(n13654), .ZN(n19974) );
  OAI21_X1 U16935 ( .B1(n14712), .B2(n19974), .A(n13655), .ZN(n13659) );
  AOI211_X1 U16936 ( .C1(n14574), .C2(n14022), .A(n13657), .B(n13656), .ZN(
        n20074) );
  NOR2_X1 U16937 ( .A1(n20074), .A2(n13660), .ZN(n13658) );
  AOI211_X1 U16938 ( .C1(n20078), .C2(n13660), .A(n13659), .B(n13658), .ZN(
        n13661) );
  OAI21_X1 U16939 ( .B1(n16025), .B2(n13662), .A(n13661), .ZN(P1_U3028) );
  NAND2_X1 U16940 ( .A1(n13689), .A2(n13663), .ZN(n13692) );
  NOR2_X1 U16941 ( .A1(n20094), .A2(n20581), .ZN(n13688) );
  NOR2_X1 U16942 ( .A1(n20182), .A2(n20906), .ZN(n20459) );
  NAND2_X1 U16943 ( .A1(n20328), .A2(n20459), .ZN(n20325) );
  OAI211_X1 U16944 ( .C1(n20459), .C2(n20096), .A(n20460), .B(n20325), .ZN(
        n13666) );
  AOI22_X1 U16945 ( .A1(n13688), .A2(n13666), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20094), .ZN(n13667) );
  OAI21_X1 U16946 ( .B1(n13668), .B2(n13692), .A(n13667), .ZN(P1_U3475) );
  AOI21_X1 U16947 ( .B1(n20906), .B2(n20182), .A(n20459), .ZN(n13670) );
  AOI22_X1 U16948 ( .A1(n13688), .A2(n13670), .B1(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n20094), .ZN(n13671) );
  OAI21_X1 U16949 ( .B1(n13669), .B2(n13692), .A(n13671), .ZN(P1_U3477) );
  AOI21_X1 U16950 ( .B1(n13674), .B2(n13573), .A(n13673), .ZN(n19962) );
  INV_X1 U16951 ( .A(n19962), .ZN(n13853) );
  INV_X1 U16952 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20029) );
  OAI222_X1 U16953 ( .A1(n13853), .A2(n14431), .B1(n14075), .B2(n20134), .C1(
        n14409), .C2(n20029), .ZN(P1_U2900) );
  XOR2_X1 U16954 ( .A(n13634), .B(n13681), .Z(n13680) );
  OR2_X1 U16955 ( .A1(n13628), .A2(n13675), .ZN(n13677) );
  AND2_X1 U16956 ( .A1(n13677), .A2(n13676), .ZN(n16210) );
  NOR2_X1 U16957 ( .A1(n13251), .A2(n14812), .ZN(n13678) );
  AOI21_X1 U16958 ( .B1(n16210), .B2(n13251), .A(n13678), .ZN(n13679) );
  OAI21_X1 U16959 ( .B1(n13680), .B2(n14966), .A(n13679), .ZN(P2_U2877) );
  INV_X1 U16960 ( .A(n13681), .ZN(n13682) );
  NOR2_X1 U16961 ( .A1(n13634), .A2(n13682), .ZN(n13685) );
  OAI211_X1 U16962 ( .C1(n13685), .C2(n13684), .A(n14941), .B(n13683), .ZN(
        n13687) );
  NAND2_X1 U16963 ( .A1(n13257), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n13686) );
  OAI211_X1 U16964 ( .C1(n15497), .C2(n13257), .A(n13687), .B(n13686), .ZN(
        P2_U2876) );
  INV_X1 U16965 ( .A(n13688), .ZN(n13691) );
  XNOR2_X1 U16966 ( .A(n20459), .B(n13664), .ZN(n13690) );
  OAI222_X1 U16967 ( .A1(n13692), .A2(n13425), .B1(n13691), .B2(n13690), .C1(
        n20487), .C2(n13689), .ZN(P1_U3476) );
  OR2_X1 U16968 ( .A1(n13673), .A2(n13694), .ZN(n13695) );
  AND2_X1 U16969 ( .A1(n13693), .A2(n13695), .ZN(n19948) );
  INV_X1 U16970 ( .A(n19948), .ZN(n13889) );
  INV_X1 U16971 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13696) );
  OAI222_X1 U16972 ( .A1(n13889), .A2(n14431), .B1(n14075), .B2(n20138), .C1(
        n13696), .C2(n14409), .ZN(P1_U2899) );
  XNOR2_X1 U16973 ( .A(n13683), .B(n13727), .ZN(n13701) );
  AND2_X1 U16974 ( .A1(n9782), .A2(n13697), .ZN(n13698) );
  NOR2_X1 U16975 ( .A1(n13725), .A2(n13698), .ZN(n18970) );
  INV_X1 U16976 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n20941) );
  NOR2_X1 U16977 ( .A1(n13251), .A2(n20941), .ZN(n13699) );
  AOI21_X1 U16978 ( .B1(n18970), .B2(n13251), .A(n13699), .ZN(n13700) );
  OAI21_X1 U16979 ( .B1(n13701), .B2(n14966), .A(n13700), .ZN(P2_U2875) );
  NAND2_X1 U16980 ( .A1(n13702), .A2(n20093), .ZN(n13705) );
  INV_X1 U16981 ( .A(n13703), .ZN(n13704) );
  NAND2_X1 U16982 ( .A1(n13705), .A2(n13704), .ZN(n20083) );
  OAI222_X1 U16983 ( .A1(n20068), .A2(n14359), .B1(n14350), .B2(n11790), .C1(
        n20083), .C2(n20002), .ZN(P1_U2872) );
  NAND2_X1 U16984 ( .A1(n13693), .A2(n13707), .ZN(n13708) );
  AND2_X1 U16985 ( .A1(n13706), .A2(n13708), .ZN(n20005) );
  INV_X1 U16986 ( .A(n20005), .ZN(n13709) );
  OAI222_X1 U16987 ( .A1(n13709), .A2(n14431), .B1(n14075), .B2(n20143), .C1(
        n14409), .C2(n11399), .ZN(P1_U2898) );
  NAND2_X1 U16988 ( .A1(n13711), .A2(n13710), .ZN(n13714) );
  NAND2_X1 U16989 ( .A1(n13712), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13713) );
  NAND2_X1 U16990 ( .A1(n13715), .A2(n13904), .ZN(n13718) );
  XNOR2_X1 U16991 ( .A(n13807), .B(n13805), .ZN(n13716) );
  NAND2_X1 U16992 ( .A1(n13716), .A2(n13955), .ZN(n13717) );
  NAND2_X1 U16993 ( .A1(n13718), .A2(n13717), .ZN(n13801) );
  XNOR2_X1 U16994 ( .A(n13801), .B(n20073), .ZN(n13799) );
  XOR2_X1 U16995 ( .A(n9738), .B(n13799), .Z(n20076) );
  INV_X1 U16996 ( .A(n20076), .ZN(n13722) );
  NAND2_X1 U16997 ( .A1(n16053), .A2(P1_REIP_REG_4__SCAN_IN), .ZN(n20072) );
  NAND2_X1 U16998 ( .A1(n20060), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13719) );
  OAI211_X1 U16999 ( .C1(n15978), .C2(n19966), .A(n20072), .B(n13719), .ZN(
        n13720) );
  AOI21_X1 U17000 ( .B1(n19962), .B2(n15975), .A(n13720), .ZN(n13721) );
  OAI21_X1 U17001 ( .B1(n13722), .B2(n15962), .A(n13721), .ZN(P1_U2995) );
  NOR2_X1 U17002 ( .A1(n13725), .A2(n13724), .ZN(n13726) );
  OR2_X1 U17003 ( .A1(n13723), .A2(n13726), .ZN(n15482) );
  NOR2_X1 U17004 ( .A1(n13683), .A2(n13727), .ZN(n13731) );
  CLKBUF_X1 U17005 ( .A(n13728), .Z(n13792) );
  INV_X1 U17006 ( .A(n13792), .ZN(n13729) );
  OAI211_X1 U17007 ( .C1(n13731), .C2(n13730), .A(n13729), .B(n14941), .ZN(
        n13733) );
  NAND2_X1 U17008 ( .A1(n13257), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13732) );
  OAI211_X1 U17009 ( .C1(n15482), .C2(n13257), .A(n13733), .B(n13732), .ZN(
        P2_U2874) );
  NAND2_X1 U17010 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20722), .ZN(n15729) );
  OAI211_X1 U17011 ( .C1(n20639), .C2(n15729), .A(n20066), .B(n13734), .ZN(
        n13735) );
  INV_X1 U17012 ( .A(n13735), .ZN(n13738) );
  NOR2_X1 U17013 ( .A1(n14146), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n13736) );
  NAND2_X1 U17014 ( .A1(n14135), .A2(n13736), .ZN(n13737) );
  INV_X1 U17015 ( .A(n13739), .ZN(n13740) );
  NAND2_X1 U17016 ( .A1(n13740), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14110) );
  INV_X1 U17017 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14181) );
  INV_X1 U17018 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13741) );
  NOR2_X1 U17019 ( .A1(n14198), .A2(n14146), .ZN(n13743) );
  AND2_X1 U17020 ( .A1(n11184), .A2(n13747), .ZN(n13744) );
  INV_X1 U17021 ( .A(n19996), .ZN(n13790) );
  INV_X1 U17022 ( .A(n13747), .ZN(n13745) );
  NOR2_X1 U17023 ( .A1(n13746), .A2(n13745), .ZN(n19983) );
  AND2_X1 U17024 ( .A1(n13751), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13749) );
  NAND2_X1 U17025 ( .A1(n20718), .A2(n20906), .ZN(n15724) );
  INV_X1 U17026 ( .A(n13749), .ZN(n13752) );
  INV_X1 U17027 ( .A(n15724), .ZN(n13750) );
  OAI21_X1 U17028 ( .B1(n13751), .B2(n15723), .A(n13750), .ZN(n13754) );
  NAND3_X1 U17029 ( .A1(n13752), .A2(n13754), .A3(n13753), .ZN(n19986) );
  OAI22_X1 U17030 ( .A1(n20083), .A2(n19987), .B1(n11790), .B2(n19986), .ZN(
        n13757) );
  INV_X1 U17031 ( .A(n13753), .ZN(n13755) );
  AND2_X1 U17032 ( .A1(n19927), .A2(n19969), .ZN(n19929) );
  INV_X1 U17033 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n20711) );
  NOR2_X1 U17034 ( .A1(n19929), .A2(n20711), .ZN(n13756) );
  AOI211_X1 U17035 ( .C1(n14145), .C2(n19983), .A(n13757), .B(n13756), .ZN(
        n13760) );
  OAI21_X1 U17036 ( .B1(n19991), .B2(n19993), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13759) );
  OAI211_X1 U17037 ( .C1(n13790), .C2(n20068), .A(n13760), .B(n13759), .ZN(
        P1_U2840) );
  NAND2_X1 U17038 ( .A1(n13762), .A2(n13761), .ZN(n13764) );
  XNOR2_X1 U17039 ( .A(n13764), .B(n13763), .ZN(n13783) );
  XOR2_X1 U17040 ( .A(n13765), .B(n13766), .Z(n13781) );
  OAI22_X1 U17041 ( .A1(n16194), .A2(n13767), .B1(n10803), .B2(n19012), .ZN(
        n13768) );
  AOI21_X1 U17042 ( .B1(n16187), .B2(n14845), .A(n13768), .ZN(n13769) );
  OAI21_X1 U17043 ( .B1(n13478), .B2(n16186), .A(n13769), .ZN(n13770) );
  AOI21_X1 U17044 ( .B1(n13781), .B2(n16188), .A(n13770), .ZN(n13771) );
  OAI21_X1 U17045 ( .B1(n13783), .B2(n19198), .A(n13771), .ZN(P2_U3011) );
  MUX2_X1 U17046 ( .A(n13772), .B(n13971), .S(
        P2_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(n13780) );
  OR2_X1 U17047 ( .A1(n13774), .A2(n13773), .ZN(n13776) );
  NAND2_X1 U17048 ( .A1(n13776), .A2(n13775), .ZN(n19096) );
  AOI22_X1 U17049 ( .A1(n13777), .A2(n19212), .B1(P2_REIP_REG_3__SCAN_IN), 
        .B2(n19206), .ZN(n13778) );
  OAI21_X1 U17050 ( .B1(n19096), .B2(n16197), .A(n13778), .ZN(n13779) );
  AOI211_X1 U17051 ( .C1(n13781), .C2(n16223), .A(n13780), .B(n13779), .ZN(
        n13782) );
  OAI21_X1 U17052 ( .B1(n13783), .B2(n16227), .A(n13782), .ZN(P2_U3043) );
  INV_X1 U17053 ( .A(n13669), .ZN(n20553) );
  NAND2_X1 U17054 ( .A1(n20553), .A2(n19983), .ZN(n13785) );
  AOI22_X1 U17055 ( .A1(n19971), .A2(P1_EBX_REG_1__SCAN_IN), .B1(n19982), .B2(
        n20705), .ZN(n13784) );
  OAI211_X1 U17056 ( .C1(n13888), .C2(n19987), .A(n13785), .B(n13784), .ZN(
        n13786) );
  AOI21_X1 U17057 ( .B1(n19967), .B2(P1_REIP_REG_1__SCAN_IN), .A(n13786), .ZN(
        n13787) );
  OAI21_X1 U17058 ( .B1(n19965), .B2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13787), .ZN(n13788) );
  AOI21_X1 U17059 ( .B1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19991), .A(
        n13788), .ZN(n13789) );
  OAI21_X1 U17060 ( .B1(n13790), .B2(n13886), .A(n13789), .ZN(P1_U2839) );
  XNOR2_X1 U17061 ( .A(n13792), .B(n13791), .ZN(n13796) );
  OR2_X1 U17062 ( .A1(n13723), .A2(n13793), .ZN(n13794) );
  NAND2_X1 U17063 ( .A1(n13104), .A2(n13794), .ZN(n18949) );
  MUX2_X1 U17064 ( .A(n18949), .B(n12106), .S(n13257), .Z(n13795) );
  OAI21_X1 U17065 ( .B1(n13796), .B2(n14966), .A(n13795), .ZN(P2_U2873) );
  NAND2_X1 U17066 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20077) );
  OR2_X1 U17067 ( .A1(n20077), .A2(n14022), .ZN(n13798) );
  NOR2_X1 U17068 ( .A1(n13812), .A2(n20077), .ZN(n14021) );
  AND2_X1 U17069 ( .A1(n14021), .A2(n13797), .ZN(n14565) );
  OAI21_X1 U17070 ( .B1(n14565), .B2(n15755), .A(n14577), .ZN(n14707) );
  AOI21_X1 U17071 ( .B1(n13798), .B2(n14574), .A(n14707), .ZN(n13915) );
  NAND2_X1 U17072 ( .A1(n13800), .A2(n13799), .ZN(n13803) );
  NAND2_X1 U17073 ( .A1(n13801), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13802) );
  NAND2_X1 U17074 ( .A1(n13804), .A2(n13904), .ZN(n13811) );
  INV_X1 U17075 ( .A(n13805), .ZN(n13806) );
  NOR2_X1 U17076 ( .A1(n13807), .A2(n13806), .ZN(n13809) );
  NAND2_X1 U17077 ( .A1(n13809), .A2(n13808), .ZN(n13906) );
  OAI211_X1 U17078 ( .C1(n13809), .C2(n13808), .A(n13906), .B(n13955), .ZN(
        n13810) );
  NAND2_X1 U17079 ( .A1(n13811), .A2(n13810), .ZN(n13892) );
  XNOR2_X1 U17080 ( .A(n13892), .B(n13812), .ZN(n13890) );
  XOR2_X1 U17081 ( .A(n13891), .B(n13890), .Z(n15981) );
  NAND2_X1 U17082 ( .A1(n15981), .A2(n20082), .ZN(n13818) );
  NOR2_X1 U17083 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n20077), .ZN(
        n13917) );
  NOR2_X1 U17084 ( .A1(n13813), .A2(n13814), .ZN(n13815) );
  OR2_X1 U17085 ( .A1(n16050), .A2(n13815), .ZN(n19941) );
  NAND2_X1 U17086 ( .A1(n16053), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n15982) );
  OAI21_X1 U17087 ( .B1(n14712), .B2(n19941), .A(n15982), .ZN(n13816) );
  AOI21_X1 U17088 ( .B1(n20078), .B2(n13917), .A(n13816), .ZN(n13817) );
  OAI211_X1 U17089 ( .C1(n13915), .C2(n13812), .A(n13818), .B(n13817), .ZN(
        P1_U3026) );
  NAND2_X1 U17090 ( .A1(n13706), .A2(n13820), .ZN(n13821) );
  AND2_X1 U17091 ( .A1(n13819), .A2(n13821), .ZN(n19917) );
  INV_X1 U17092 ( .A(n19917), .ZN(n13848) );
  OAI222_X1 U17093 ( .A1(n13848), .A2(n14431), .B1(n14075), .B2(n20147), .C1(
        n13822), .C2(n14409), .ZN(P1_U2897) );
  NOR2_X2 U17094 ( .A1(n19610), .A2(n19815), .ZN(n19728) );
  OAI21_X1 U17095 ( .B1(n19728), .B2(n19281), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13823) );
  NAND2_X1 U17096 ( .A1(n13823), .A2(n19820), .ZN(n13836) );
  NAND2_X1 U17097 ( .A1(n19824), .A2(n12371), .ZN(n19324) );
  OR2_X1 U17098 ( .A1(n19324), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19265) );
  NOR2_X1 U17099 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19265), .ZN(
        n19255) );
  OR2_X1 U17100 ( .A1(n19724), .A2(n19255), .ZN(n13833) );
  INV_X1 U17101 ( .A(n19255), .ZN(n13840) );
  NAND2_X1 U17102 ( .A1(n19636), .A2(n13840), .ZN(n13824) );
  AOI21_X1 U17103 ( .B1(n12010), .B2(n19385), .A(n13824), .ZN(n13825) );
  NAND2_X1 U17104 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19843) );
  AOI21_X1 U17105 ( .B1(n10692), .B2(n16287), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n19866) );
  AOI22_X4 U17106 ( .A1(n18874), .A2(n14103), .B1(n19843), .B2(n19866), .ZN(
        n19436) );
  NOR2_X1 U17107 ( .A1(n13825), .A2(n19436), .ZN(n13826) );
  NOR2_X1 U17108 ( .A1(n19636), .A2(n19868), .ZN(n19834) );
  AOI22_X1 U17109 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19251), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n19252), .ZN(n19691) );
  AOI22_X1 U17110 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19252), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19251), .ZN(n19649) );
  INV_X1 U17111 ( .A(n19253), .ZN(n13831) );
  NAND2_X1 U17112 ( .A1(n9743), .A2(n13831), .ZN(n19270) );
  OAI22_X1 U17113 ( .A1(n19649), .A2(n19289), .B1(n19270), .B2(n13840), .ZN(
        n13832) );
  AOI21_X1 U17114 ( .B1(n19728), .B2(n19646), .A(n13832), .ZN(n13838) );
  INV_X1 U17115 ( .A(n13833), .ZN(n13835) );
  OAI21_X1 U17116 ( .B1(n12010), .B2(n19255), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13834) );
  NOR2_X2 U17117 ( .A1(n14005), .A2(n19436), .ZN(n19687) );
  NAND2_X1 U17118 ( .A1(n19257), .A2(n19687), .ZN(n13837) );
  OAI211_X1 U17119 ( .C1(n19250), .C2(n13839), .A(n13838), .B(n13837), .ZN(
        P2_U3049) );
  INV_X1 U17120 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13844) );
  AOI22_X1 U17121 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n19251), .B1(
        BUF1_REG_24__SCAN_IN), .B2(n19252), .ZN(n19685) );
  INV_X1 U17122 ( .A(n19685), .ZN(n19632) );
  AOI22_X1 U17123 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19252), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19251), .ZN(n19645) );
  NOR2_X2 U17124 ( .A1(n10690), .A2(n19253), .ZN(n19673) );
  INV_X1 U17125 ( .A(n19673), .ZN(n15634) );
  OAI22_X1 U17126 ( .A1(n19645), .A2(n19289), .B1(n15634), .B2(n13840), .ZN(
        n13841) );
  AOI21_X1 U17127 ( .B1(n19728), .B2(n19632), .A(n13841), .ZN(n13843) );
  NOR2_X2 U17128 ( .A1(n19114), .A2(n19436), .ZN(n19674) );
  NAND2_X1 U17129 ( .A1(n19257), .A2(n19674), .ZN(n13842) );
  OAI211_X1 U17130 ( .C1(n19250), .C2(n13844), .A(n13843), .B(n13842), .ZN(
        P2_U3048) );
  INV_X1 U17131 ( .A(n16052), .ZN(n13847) );
  INV_X1 U17132 ( .A(n13845), .ZN(n13846) );
  OAI21_X1 U17133 ( .B1(n13847), .B2(n13846), .A(n13866), .ZN(n19908) );
  OAI222_X1 U17134 ( .A1(n19908), .A2(n20002), .B1(n19912), .B2(n14350), .C1(
        n13848), .C2(n14359), .ZN(P1_U2865) );
  AND2_X1 U17135 ( .A1(n13850), .A2(n13849), .ZN(n13851) );
  NOR2_X1 U17136 ( .A1(n13813), .A2(n13851), .ZN(n20069) );
  AOI22_X1 U17137 ( .A1(n11892), .A2(n20069), .B1(n14337), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n13852) );
  OAI21_X1 U17138 ( .B1(n13853), .B2(n14359), .A(n13852), .ZN(P1_U2868) );
  INV_X1 U17139 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n13859) );
  OAI211_X1 U17140 ( .C1(n10020), .C2(n13856), .A(n14941), .B(n13855), .ZN(
        n13858) );
  NAND2_X1 U17141 ( .A1(n16167), .A2(n13251), .ZN(n13857) );
  OAI211_X1 U17142 ( .C1(n13251), .C2(n13859), .A(n13858), .B(n13857), .ZN(
        P2_U2872) );
  INV_X1 U17143 ( .A(n13819), .ZN(n13863) );
  INV_X1 U17144 ( .A(n13860), .ZN(n13861) );
  OAI21_X1 U17145 ( .B1(n13863), .B2(n13862), .A(n13861), .ZN(n13963) );
  AOI22_X1 U17146 ( .A1(n14429), .A2(n14384), .B1(P1_EAX_REG_8__SCAN_IN), .B2(
        n14428), .ZN(n13864) );
  OAI21_X1 U17147 ( .B1(n13963), .B2(n14431), .A(n13864), .ZN(P1_U2896) );
  AND2_X1 U17148 ( .A1(n13866), .A2(n13865), .ZN(n13867) );
  NOR2_X1 U17149 ( .A1(n13927), .A2(n13867), .ZN(n16040) );
  INV_X1 U17150 ( .A(n16040), .ZN(n13868) );
  OAI22_X1 U17151 ( .A1(n20002), .A2(n13868), .B1(n13876), .B2(n14350), .ZN(
        n13869) );
  INV_X1 U17152 ( .A(n13869), .ZN(n13870) );
  OAI21_X1 U17153 ( .B1(n13963), .B2(n14359), .A(n13870), .ZN(P1_U2864) );
  INV_X1 U17154 ( .A(n14359), .ZN(n20004) );
  OAI22_X1 U17155 ( .A1(n20002), .A2(n19974), .B1(n13871), .B2(n14350), .ZN(
        n13872) );
  AOI21_X1 U17156 ( .B1(n19978), .B2(n20004), .A(n13872), .ZN(n13873) );
  INV_X1 U17157 ( .A(n13873), .ZN(P1_U2869) );
  INV_X1 U17158 ( .A(n13959), .ZN(n13883) );
  INV_X1 U17159 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20908) );
  INV_X1 U17160 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n13874) );
  INV_X1 U17161 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n19936) );
  NAND4_X1 U17162 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n19937)
         );
  NOR3_X1 U17163 ( .A1(n13874), .A2(n19936), .A3(n19937), .ZN(n19915) );
  NAND2_X1 U17164 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19915), .ZN(n13877) );
  NOR2_X1 U17165 ( .A1(n20908), .A2(n13877), .ZN(n15826) );
  INV_X1 U17166 ( .A(n15826), .ZN(n13875) );
  NAND2_X1 U17167 ( .A1(n19982), .A2(n13875), .ZN(n13878) );
  OAI22_X1 U17168 ( .A1(n13878), .A2(n13877), .B1(n13876), .B2(n19986), .ZN(
        n13882) );
  NAND2_X1 U17169 ( .A1(n19927), .A2(n13878), .ZN(n14297) );
  INV_X1 U17170 ( .A(n14297), .ZN(n15828) );
  AOI22_X1 U17171 ( .A1(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19991), .B1(
        n19959), .B2(n16040), .ZN(n13880) );
  NAND2_X1 U17172 ( .A1(n19927), .A2(n13879), .ZN(n19953) );
  OAI211_X1 U17173 ( .C1(n15828), .C2(n20908), .A(n13880), .B(n19953), .ZN(
        n13881) );
  AOI211_X1 U17174 ( .C1(n19993), .C2(n13883), .A(n13882), .B(n13881), .ZN(
        n13884) );
  OAI21_X1 U17175 ( .B1(n15894), .B2(n13963), .A(n13884), .ZN(P1_U2832) );
  INV_X1 U17176 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n19985) );
  OAI222_X1 U17177 ( .A1(n19988), .A2(n20002), .B1(n19985), .B2(n14350), .C1(
        n13885), .C2(n14359), .ZN(P1_U2870) );
  INV_X1 U17178 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13887) );
  OAI222_X1 U17179 ( .A1(n13888), .A2(n20002), .B1(n13887), .B2(n14350), .C1(
        n13886), .C2(n14359), .ZN(P1_U2871) );
  OAI222_X1 U17180 ( .A1(n19941), .A2(n20002), .B1(n19940), .B2(n14350), .C1(
        n13889), .C2(n14359), .ZN(P1_U2867) );
  NAND2_X1 U17181 ( .A1(n14021), .A2(n20078), .ZN(n16030) );
  NOR2_X1 U17182 ( .A1(n16059), .A2(n16030), .ZN(n16043) );
  INV_X1 U17183 ( .A(n16043), .ZN(n13922) );
  NAND2_X1 U17184 ( .A1(n13891), .A2(n13890), .ZN(n13894) );
  NAND2_X1 U17185 ( .A1(n13892), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13893) );
  INV_X1 U17186 ( .A(n13896), .ZN(n13897) );
  OR2_X1 U17187 ( .A1(n13952), .A2(n13897), .ZN(n13900) );
  XNOR2_X1 U17188 ( .A(n13906), .B(n13907), .ZN(n13898) );
  NAND2_X1 U17189 ( .A1(n13898), .A2(n13955), .ZN(n13899) );
  NAND2_X1 U17190 ( .A1(n13901), .A2(n16059), .ZN(n15973) );
  INV_X1 U17191 ( .A(n13901), .ZN(n13902) );
  NAND2_X1 U17192 ( .A1(n13902), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15972) );
  NAND2_X1 U17193 ( .A1(n13905), .A2(n13904), .ZN(n13911) );
  INV_X1 U17194 ( .A(n13906), .ZN(n13908) );
  NAND2_X1 U17195 ( .A1(n13908), .A2(n13907), .ZN(n13953) );
  XNOR2_X1 U17196 ( .A(n13953), .B(n13954), .ZN(n13909) );
  NAND2_X1 U17197 ( .A1(n13909), .A2(n13955), .ZN(n13910) );
  NAND2_X1 U17198 ( .A1(n13911), .A2(n13910), .ZN(n13947) );
  XNOR2_X1 U17199 ( .A(n13947), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13912) );
  NAND2_X1 U17200 ( .A1(n13913), .A2(n13912), .ZN(n13914) );
  NAND2_X1 U17201 ( .A1(n13949), .A2(n13914), .ZN(n15968) );
  NAND2_X1 U17202 ( .A1(n15968), .A2(n20082), .ZN(n13921) );
  INV_X1 U17203 ( .A(n16018), .ZN(n13918) );
  INV_X1 U17204 ( .A(n13915), .ZN(n13916) );
  AOI21_X1 U17205 ( .B1(n13918), .B2(n13917), .A(n13916), .ZN(n16060) );
  OAI21_X1 U17206 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15995), .A(
        n16060), .ZN(n16041) );
  INV_X1 U17207 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n19909) );
  OAI22_X1 U17208 ( .A1(n14712), .A2(n19908), .B1(n19909), .B2(n20066), .ZN(
        n13919) );
  AOI21_X1 U17209 ( .B1(n16041), .B2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n13919), .ZN(n13920) );
  OAI211_X1 U17210 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n13922), .A(
        n13921), .B(n13920), .ZN(P1_U3024) );
  NOR2_X1 U17211 ( .A1(n13860), .A2(n13924), .ZN(n13925) );
  OR2_X1 U17212 ( .A1(n13923), .A2(n13925), .ZN(n14040) );
  NAND2_X1 U17213 ( .A1(n19982), .A2(n15826), .ZN(n13929) );
  OR2_X1 U17214 ( .A1(n13927), .A2(n13926), .ZN(n13928) );
  NAND2_X1 U17215 ( .A1(n14013), .A2(n13928), .ZN(n14020) );
  OAI22_X1 U17216 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n13929), .B1(n19987), 
        .B2(n14020), .ZN(n13933) );
  AOI22_X1 U17217 ( .A1(n19971), .A2(P1_EBX_REG_9__SCAN_IN), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n14297), .ZN(n13930) );
  OAI211_X1 U17218 ( .C1(n19956), .C2(n13931), .A(n13930), .B(n19953), .ZN(
        n13932) );
  AOI211_X1 U17219 ( .C1(n14039), .C2(n19993), .A(n13933), .B(n13932), .ZN(
        n13934) );
  OAI21_X1 U17220 ( .B1(n15894), .B2(n14040), .A(n13934), .ZN(P1_U2831) );
  INV_X1 U17221 ( .A(DATAI_9_), .ZN(n13936) );
  NAND2_X1 U17222 ( .A1(n20107), .A2(BUF1_REG_9__SCAN_IN), .ZN(n13935) );
  OAI21_X1 U17223 ( .B1(n20107), .B2(n13936), .A(n13935), .ZN(n20036) );
  INV_X1 U17224 ( .A(n20036), .ZN(n13938) );
  OAI222_X1 U17225 ( .A1(n14040), .A2(n14431), .B1(n14075), .B2(n13938), .C1(
        n13937), .C2(n14409), .ZN(P1_U2895) );
  AND2_X1 U17226 ( .A1(n13940), .A2(n13939), .ZN(n13942) );
  OR2_X1 U17227 ( .A1(n13942), .A2(n13941), .ZN(n18938) );
  AOI21_X1 U17228 ( .B1(n13944), .B2(n13855), .A(n13943), .ZN(n13983) );
  NAND2_X1 U17229 ( .A1(n13983), .A2(n14941), .ZN(n13946) );
  NAND2_X1 U17230 ( .A1(n13257), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n13945) );
  OAI211_X1 U17231 ( .C1(n18938), .C2(n13257), .A(n13946), .B(n13945), .ZN(
        P2_U2871) );
  OAI222_X1 U17232 ( .A1(n14020), .A2(n20002), .B1(n14350), .B2(n11819), .C1(
        n14359), .C2(n14040), .ZN(P1_U2863) );
  OR2_X1 U17233 ( .A1(n13947), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13948) );
  OR2_X1 U17234 ( .A1(n13950), .A2(n20639), .ZN(n13951) );
  OR2_X4 U17235 ( .A1(n13952), .A2(n13951), .ZN(n14160) );
  INV_X1 U17236 ( .A(n13953), .ZN(n13956) );
  NAND3_X1 U17237 ( .A1(n13956), .A2(n13955), .A3(n13954), .ZN(n13957) );
  NAND2_X1 U17238 ( .A1(n14160), .A2(n13957), .ZN(n14016) );
  XOR2_X1 U17239 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n14016), .Z(
        n13958) );
  XNOR2_X1 U17240 ( .A(n14015), .B(n13958), .ZN(n16042) );
  NAND2_X1 U17241 ( .A1(n16042), .A2(n20064), .ZN(n13962) );
  NOR2_X1 U17242 ( .A1(n20066), .A2(n20908), .ZN(n16039) );
  NOR2_X1 U17243 ( .A1(n15978), .A2(n13959), .ZN(n13960) );
  AOI211_X1 U17244 ( .C1(n20060), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16039), .B(n13960), .ZN(n13961) );
  OAI211_X1 U17245 ( .C1(n20106), .C2(n13963), .A(n13962), .B(n13961), .ZN(
        P1_U2991) );
  NOR2_X1 U17246 ( .A1(n13965), .A2(n13964), .ZN(n13966) );
  XNOR2_X1 U17247 ( .A(n13967), .B(n13966), .ZN(n16189) );
  INV_X1 U17248 ( .A(n16189), .ZN(n13982) );
  XOR2_X1 U17249 ( .A(n13968), .B(n13969), .Z(n16191) );
  AOI211_X1 U17250 ( .C1(n19209), .C2(n13970), .A(n15549), .B(n19222), .ZN(
        n13980) );
  NAND2_X1 U17251 ( .A1(n19022), .A2(n19212), .ZN(n13978) );
  AOI21_X1 U17252 ( .B1(n15426), .B2(n13972), .A(n13971), .ZN(n19210) );
  INV_X1 U17253 ( .A(n19210), .ZN(n13976) );
  XNOR2_X1 U17254 ( .A(n13973), .B(n9775), .ZN(n19085) );
  OAI22_X1 U17255 ( .A1(n16197), .A2(n19085), .B1(n19012), .B2(n13974), .ZN(
        n13975) );
  AOI21_X1 U17256 ( .B1(n13976), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n13975), .ZN(n13977) );
  NAND2_X1 U17257 ( .A1(n13978), .A2(n13977), .ZN(n13979) );
  AOI211_X1 U17258 ( .C1(n16191), .C2(n19219), .A(n13980), .B(n13979), .ZN(
        n13981) );
  OAI21_X1 U17259 ( .B1(n19215), .B2(n13982), .A(n13981), .ZN(P2_U3041) );
  INV_X1 U17260 ( .A(n13983), .ZN(n13992) );
  AND2_X1 U17261 ( .A1(n13109), .A2(n13984), .ZN(n13985) );
  OR2_X1 U17262 ( .A1(n14003), .A2(n13985), .ZN(n18937) );
  INV_X1 U17263 ( .A(n18937), .ZN(n13990) );
  INV_X1 U17264 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n19150) );
  OAI22_X1 U17265 ( .A1(n16141), .A2(n19114), .B1(n19072), .B2(n19150), .ZN(
        n13989) );
  INV_X1 U17266 ( .A(n19047), .ZN(n15026) );
  INV_X1 U17267 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n13987) );
  INV_X1 U17268 ( .A(n19049), .ZN(n15024) );
  INV_X1 U17269 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n13986) );
  OAI22_X1 U17270 ( .A1(n15026), .A2(n13987), .B1(n15024), .B2(n13986), .ZN(
        n13988) );
  AOI211_X1 U17271 ( .C1(n19106), .C2(n13990), .A(n13989), .B(n13988), .ZN(
        n13991) );
  OAI21_X1 U17272 ( .B1(n13992), .B2(n19082), .A(n13991), .ZN(P2_U2903) );
  INV_X1 U17273 ( .A(n13993), .ZN(n13994) );
  OAI21_X1 U17274 ( .B1(n13923), .B2(n13995), .A(n13994), .ZN(n15907) );
  INV_X1 U17275 ( .A(DATAI_10_), .ZN(n13997) );
  NAND2_X1 U17276 ( .A1(n20107), .A2(BUF1_REG_10__SCAN_IN), .ZN(n13996) );
  OAI21_X1 U17277 ( .B1(n20107), .B2(n13997), .A(n13996), .ZN(n20038) );
  INV_X1 U17278 ( .A(n20038), .ZN(n13999) );
  OAI222_X1 U17279 ( .A1(n15907), .A2(n14431), .B1(n14075), .B2(n13999), .C1(
        n13998), .C2(n14409), .ZN(P1_U2894) );
  AND2_X1 U17280 ( .A1(n13943), .A2(n14001), .ZN(n14959) );
  INV_X1 U17281 ( .A(n14959), .ZN(n14000) );
  OAI21_X1 U17282 ( .B1(n13943), .B2(n14001), .A(n14000), .ZN(n14967) );
  OR2_X1 U17283 ( .A1(n14003), .A2(n14002), .ZN(n14004) );
  NAND2_X1 U17284 ( .A1(n9827), .A2(n14004), .ZN(n18930) );
  INV_X1 U17285 ( .A(n18930), .ZN(n14010) );
  INV_X1 U17286 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n19147) );
  OAI22_X1 U17287 ( .A1(n16141), .A2(n14005), .B1(n19072), .B2(n19147), .ZN(
        n14009) );
  INV_X1 U17288 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n14007) );
  INV_X1 U17289 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n14006) );
  OAI22_X1 U17290 ( .A1(n15026), .A2(n14007), .B1(n15024), .B2(n14006), .ZN(
        n14008) );
  AOI211_X1 U17291 ( .C1(n19106), .C2(n14010), .A(n14009), .B(n14008), .ZN(
        n14011) );
  OAI21_X1 U17292 ( .B1(n14967), .B2(n19082), .A(n14011), .ZN(P2_U2902) );
  NAND2_X1 U17293 ( .A1(n14013), .A2(n14012), .ZN(n14014) );
  NAND2_X1 U17294 ( .A1(n14032), .A2(n14014), .ZN(n16027) );
  INV_X1 U17295 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n15902) );
  OAI222_X1 U17296 ( .A1(n16027), .A2(n20002), .B1(n15902), .B2(n14350), .C1(
        n14359), .C2(n15907), .ZN(P1_U2862) );
  MUX2_X1 U17297 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n14158), .S(
        n14160), .Z(n14018) );
  NAND2_X1 U17298 ( .A1(n14016), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14017) );
  XOR2_X1 U17299 ( .A(n14018), .B(n14156), .Z(n14044) );
  NAND3_X1 U17300 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16031) );
  NOR2_X1 U17301 ( .A1(n16031), .A2(n16030), .ZN(n14027) );
  INV_X1 U17302 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n14019) );
  OR2_X1 U17303 ( .A1(n20066), .A2(n14019), .ZN(n14037) );
  OAI21_X1 U17304 ( .B1(n14712), .B2(n14020), .A(n14037), .ZN(n14026) );
  INV_X1 U17305 ( .A(n14021), .ZN(n14023) );
  NOR2_X1 U17306 ( .A1(n14023), .A2(n14022), .ZN(n14706) );
  OAI211_X1 U17307 ( .C1(n14706), .C2(n14705), .A(n14565), .B(n14577), .ZN(
        n14024) );
  NAND2_X1 U17308 ( .A1(n15995), .A2(n14577), .ZN(n14582) );
  OAI21_X1 U17309 ( .B1(n14024), .B2(n16031), .A(n14582), .ZN(n16037) );
  NOR2_X1 U17310 ( .A1(n16037), .A2(n14158), .ZN(n14025) );
  AOI211_X1 U17311 ( .C1(n14027), .C2(n14158), .A(n14026), .B(n14025), .ZN(
        n14028) );
  OAI21_X1 U17312 ( .B1(n14044), .B2(n16025), .A(n14028), .ZN(P1_U3022) );
  OR2_X1 U17313 ( .A1(n13993), .A2(n14029), .ZN(n14030) );
  NAND2_X1 U17314 ( .A1(n14064), .A2(n14030), .ZN(n14066) );
  XNOR2_X1 U17315 ( .A(n14066), .B(n14063), .ZN(n15963) );
  NAND2_X1 U17316 ( .A1(n14032), .A2(n14031), .ZN(n14033) );
  NAND2_X1 U17317 ( .A1(n14071), .A2(n14033), .ZN(n15896) );
  OAI22_X1 U17318 ( .A1(n20002), .A2(n15896), .B1(n14034), .B2(n14350), .ZN(
        n14035) );
  AOI21_X1 U17319 ( .B1(n15963), .B2(n20004), .A(n14035), .ZN(n14036) );
  INV_X1 U17320 ( .A(n14036), .ZN(P1_U2861) );
  OAI21_X1 U17321 ( .B1(n15984), .B2(n13931), .A(n14037), .ZN(n14038) );
  AOI21_X1 U17322 ( .B1(n15979), .B2(n14039), .A(n14038), .ZN(n14043) );
  INV_X1 U17323 ( .A(n14040), .ZN(n14041) );
  NAND2_X1 U17324 ( .A1(n14041), .A2(n15975), .ZN(n14042) );
  OAI211_X1 U17325 ( .C1(n14044), .C2(n15962), .A(n14043), .B(n14042), .ZN(
        P1_U2990) );
  INV_X1 U17326 ( .A(n15963), .ZN(n14049) );
  INV_X1 U17327 ( .A(DATAI_11_), .ZN(n14046) );
  NAND2_X1 U17328 ( .A1(n20107), .A2(BUF1_REG_11__SCAN_IN), .ZN(n14045) );
  OAI21_X1 U17329 ( .B1(n20107), .B2(n14046), .A(n14045), .ZN(n20040) );
  INV_X1 U17330 ( .A(n20040), .ZN(n14048) );
  OAI222_X1 U17331 ( .A1(n14049), .A2(n14431), .B1(n14075), .B2(n14048), .C1(
        n14047), .C2(n14409), .ZN(P1_U2893) );
  NOR2_X1 U17332 ( .A1(n14051), .A2(n14052), .ZN(n14053) );
  OR2_X1 U17333 ( .A1(n14050), .A2(n14053), .ZN(n15877) );
  INV_X1 U17334 ( .A(n14061), .ZN(n14355) );
  AOI21_X1 U17335 ( .B1(n14054), .B2(n14082), .A(n14355), .ZN(n16011) );
  AOI22_X1 U17336 ( .A1(n16011), .A2(n11892), .B1(n14337), .B2(
        P1_EBX_REG_14__SCAN_IN), .ZN(n14055) );
  OAI21_X1 U17337 ( .B1(n15877), .B2(n14359), .A(n14055), .ZN(P1_U2858) );
  INV_X1 U17338 ( .A(n14186), .ZN(n14057) );
  OAI222_X1 U17339 ( .A1(n15877), .A2(n14431), .B1(n14075), .B2(n14057), .C1(
        n14056), .C2(n14409), .ZN(P1_U2890) );
  OR2_X1 U17340 ( .A1(n14050), .A2(n14059), .ZN(n14060) );
  NAND2_X1 U17341 ( .A1(n14058), .A2(n14060), .ZN(n15871) );
  XNOR2_X1 U17342 ( .A(n14061), .B(n14354), .ZN(n16002) );
  AOI22_X1 U17343 ( .A1(n16002), .A2(n11892), .B1(n14337), .B2(
        P1_EBX_REG_15__SCAN_IN), .ZN(n14062) );
  OAI21_X1 U17344 ( .B1(n15871), .B2(n14359), .A(n14062), .ZN(P1_U2857) );
  INV_X1 U17345 ( .A(n14063), .ZN(n14065) );
  OAI21_X1 U17346 ( .B1(n14066), .B2(n14065), .A(n14064), .ZN(n14068) );
  NAND2_X1 U17347 ( .A1(n14068), .A2(n14067), .ZN(n14078) );
  OR2_X1 U17348 ( .A1(n14068), .A2(n14067), .ZN(n14069) );
  AOI22_X1 U17349 ( .A1(n14429), .A2(n14368), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n14428), .ZN(n14070) );
  OAI21_X1 U17350 ( .B1(n15893), .B2(n14431), .A(n14070), .ZN(P1_U2892) );
  AOI21_X1 U17351 ( .B1(n14072), .B2(n14071), .A(n14080), .ZN(n16015) );
  AOI22_X1 U17352 ( .A1(n16015), .A2(n11892), .B1(n14337), .B2(
        P1_EBX_REG_12__SCAN_IN), .ZN(n14073) );
  OAI21_X1 U17353 ( .B1(n15893), .B2(n14359), .A(n14073), .ZN(P1_U2860) );
  OAI222_X1 U17354 ( .A1(n15871), .A2(n14431), .B1(n14075), .B2(n14074), .C1(
        n14409), .C2(n11526), .ZN(P1_U2889) );
  INV_X1 U17355 ( .A(n14076), .ZN(n14077) );
  AOI21_X1 U17356 ( .B1(n14078), .B2(n14077), .A(n14051), .ZN(n14556) );
  OR2_X1 U17357 ( .A1(n14080), .A2(n14079), .ZN(n14081) );
  NAND2_X1 U17358 ( .A1(n14082), .A2(n14081), .ZN(n14694) );
  OAI22_X1 U17359 ( .A1(n14694), .A2(n20002), .B1(n14083), .B2(n14350), .ZN(
        n14084) );
  AOI21_X1 U17360 ( .B1(n14556), .B2(n20004), .A(n14084), .ZN(n14085) );
  INV_X1 U17361 ( .A(n14085), .ZN(P1_U2859) );
  NAND3_X1 U17362 ( .A1(n14086), .A2(n15676), .A3(n16785), .ZN(n18200) );
  NOR2_X1 U17363 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18200), .ZN(n14087) );
  NAND3_X1 U17364 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18806)
         );
  OAI21_X1 U17365 ( .B1(n14087), .B2(n18806), .A(n18452), .ZN(n18206) );
  INV_X1 U17366 ( .A(n18206), .ZN(n14088) );
  NOR2_X1 U17367 ( .A1(n18848), .A2(n17829), .ZN(n15656) );
  AOI21_X1 U17368 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n15656), .ZN(n15657) );
  NOR2_X1 U17369 ( .A1(n14088), .A2(n15657), .ZN(n14090) );
  INV_X1 U17370 ( .A(n18359), .ZN(n18209) );
  NOR2_X1 U17371 ( .A1(n18808), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18250) );
  OR2_X1 U17372 ( .A1(n18250), .A2(n14088), .ZN(n15655) );
  OR2_X1 U17373 ( .A1(n18209), .A2(n15655), .ZN(n14089) );
  MUX2_X1 U17374 ( .A(n14090), .B(n14089), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  NOR2_X1 U17375 ( .A1(n18874), .A2(n19843), .ZN(n16298) );
  AND3_X1 U17376 ( .A1(n14093), .A2(n14092), .A3(n14091), .ZN(n14097) );
  INV_X1 U17377 ( .A(n19118), .ZN(n14095) );
  INV_X1 U17378 ( .A(n12221), .ZN(n14094) );
  NAND3_X1 U17379 ( .A1(n14095), .A2(n14094), .A3(n16263), .ZN(n14096) );
  OAI22_X1 U17380 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19385), .B1(n16242), 
        .B2(n18880), .ZN(n14098) );
  AOI21_X1 U17381 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16298), .A(n14098), .ZN(
        n19811) );
  INV_X1 U17382 ( .A(n19811), .ZN(n19813) );
  NAND2_X1 U17383 ( .A1(n19019), .A2(n14867), .ZN(n19046) );
  OAI21_X1 U17384 ( .B1(n19019), .B2(n15557), .A(n19046), .ZN(n15574) );
  NOR2_X1 U17385 ( .A1(n15574), .A2(n16287), .ZN(n14106) );
  NAND2_X1 U17386 ( .A1(n14100), .A2(n14099), .ZN(n15570) );
  MUX2_X1 U17387 ( .A(n10775), .B(n15570), .S(n14108), .Z(n14101) );
  AOI21_X1 U17388 ( .B1(n14102), .B2(n16241), .A(n14101), .ZN(n16246) );
  INV_X1 U17389 ( .A(n14103), .ZN(n19810) );
  OAI22_X1 U17390 ( .A1(n16246), .A2(n19816), .B1(n14104), .B2(n19810), .ZN(
        n14105) );
  OAI21_X1 U17391 ( .B1(n14106), .B2(n14105), .A(n19813), .ZN(n14107) );
  OAI21_X1 U17392 ( .B1(n19813), .B2(n14108), .A(n14107), .ZN(P2_U3601) );
  NOR2_X1 U17393 ( .A1(n14140), .A2(n20105), .ZN(n14109) );
  NAND2_X1 U17394 ( .A1(n14409), .A2(n14109), .ZN(n14411) );
  INV_X1 U17395 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16354) );
  XNOR2_X1 U17396 ( .A(n14110), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14224) );
  OAI21_X1 U17397 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n14181), .A(n11423), 
        .ZN(n14133) );
  AOI22_X1 U17398 ( .A1(n11635), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n14111), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14116) );
  AOI22_X1 U17399 ( .A1(n11261), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n14112), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14115) );
  AOI22_X1 U17400 ( .A1(n11636), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9742), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14114) );
  AOI22_X1 U17401 ( .A1(n11616), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11255), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n14113) );
  NAND4_X1 U17402 ( .A1(n14116), .A2(n14115), .A3(n14114), .A4(n14113), .ZN(
        n14125) );
  AOI22_X1 U17403 ( .A1(n14117), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11149), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14123) );
  AOI22_X1 U17404 ( .A1(n14119), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n14118), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14122) );
  AOI22_X1 U17405 ( .A1(n9721), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n9750), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n14121) );
  AOI22_X1 U17406 ( .A1(n11637), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11297), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n14120) );
  NAND4_X1 U17407 ( .A1(n14123), .A2(n14122), .A3(n14121), .A4(n14120), .ZN(
        n14124) );
  NOR2_X1 U17408 ( .A1(n14125), .A2(n14124), .ZN(n14129) );
  NOR2_X1 U17409 ( .A1(n14127), .A2(n14126), .ZN(n14128) );
  XOR2_X1 U17410 ( .A(n14129), .B(n14128), .Z(n14131) );
  NOR2_X1 U17411 ( .A1(n14131), .A2(n14130), .ZN(n14132) );
  AOI211_X1 U17412 ( .C1(n14137), .C2(P1_EAX_REG_30__SCAN_IN), .A(n14133), .B(
        n14132), .ZN(n14134) );
  AOI21_X1 U17413 ( .B1(n14135), .B2(n14224), .A(n14134), .ZN(n14154) );
  AOI22_X1 U17414 ( .A1(n14137), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n14136), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n14138) );
  INV_X1 U17415 ( .A(n14138), .ZN(n14139) );
  XNOR2_X2 U17416 ( .A(n14153), .B(n14139), .ZN(n14210) );
  NAND3_X1 U17417 ( .A1(n14210), .A2(n20148), .A3(n14409), .ZN(n14143) );
  NOR3_X1 U17418 ( .A1(n14428), .A2(n20107), .A3(n14140), .ZN(n14141) );
  AOI22_X1 U17419 ( .A1(n14422), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14428), .ZN(n14142) );
  OAI211_X1 U17420 ( .C1(n14411), .C2(n16354), .A(n14143), .B(n14142), .ZN(
        P1_U2873) );
  AOI22_X1 U17421 ( .A1(n14145), .A2(n14144), .B1(n14716), .B2(n14149), .ZN(
        n15702) );
  INV_X1 U17422 ( .A(n19883), .ZN(n14147) );
  OAI22_X1 U17423 ( .A1(n15702), .A2(n14147), .B1(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n14146), .ZN(n14148) );
  AOI21_X1 U17424 ( .B1(n15731), .B2(n14149), .A(n14148), .ZN(n14152) );
  AOI21_X1 U17425 ( .B1(n15704), .B2(n19883), .A(n14151), .ZN(n14150) );
  OAI22_X1 U17426 ( .A1(n14152), .A2(n14151), .B1(n14150), .B2(n14149), .ZN(
        P1_U3474) );
  INV_X1 U17427 ( .A(n14156), .ZN(n14157) );
  NAND2_X1 U17428 ( .A1(n14160), .A2(n14158), .ZN(n14159) );
  NAND2_X1 U17429 ( .A1(n14160), .A2(n14563), .ZN(n14161) );
  NAND2_X1 U17430 ( .A1(n15946), .A2(n14161), .ZN(n14552) );
  NOR2_X1 U17431 ( .A1(n14552), .A2(n14550), .ZN(n15945) );
  NAND3_X1 U17432 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14162) );
  NAND2_X1 U17433 ( .A1(n14160), .A2(n14162), .ZN(n14163) );
  NAND2_X1 U17434 ( .A1(n15945), .A2(n14163), .ZN(n14533) );
  NAND2_X1 U17435 ( .A1(n14545), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14164) );
  NOR2_X1 U17436 ( .A1(n14160), .A2(n14165), .ZN(n14536) );
  XNOR2_X1 U17437 ( .A(n14160), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15937) );
  NAND2_X1 U17438 ( .A1(n14160), .A2(n14165), .ZN(n15934) );
  AND2_X1 U17439 ( .A1(n15937), .A2(n15934), .ZN(n14166) );
  NAND2_X1 U17440 ( .A1(n14168), .A2(n14160), .ZN(n14169) );
  INV_X1 U17441 ( .A(n14170), .ZN(n15935) );
  NAND2_X1 U17442 ( .A1(n14711), .A2(n16038), .ZN(n14544) );
  OAI21_X1 U17443 ( .B1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n14544), .A(
        n14545), .ZN(n14532) );
  INV_X1 U17444 ( .A(n14532), .ZN(n14171) );
  XNOR2_X1 U17445 ( .A(n14160), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15927) );
  NAND2_X1 U17446 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14665) );
  INV_X1 U17447 ( .A(n14665), .ZN(n14172) );
  AND2_X2 U17448 ( .A1(n14500), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14176) );
  NOR2_X1 U17449 ( .A1(n14176), .A2(n14545), .ZN(n14478) );
  INV_X1 U17450 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14571) );
  AND3_X1 U17451 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14444) );
  NAND2_X1 U17452 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14581) );
  NOR2_X2 U17453 ( .A1(n14461), .A2(n14581), .ZN(n14433) );
  INV_X1 U17454 ( .A(n14176), .ZN(n14177) );
  INV_X1 U17455 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14643) );
  NAND3_X1 U17456 ( .A1(n20956), .A2(n14635), .A3(n14643), .ZN(n14448) );
  NOR2_X1 U17457 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14609) );
  INV_X1 U17458 ( .A(n14434), .ZN(n14180) );
  INV_X1 U17459 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14179) );
  INV_X1 U17460 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14591) );
  NAND2_X1 U17461 ( .A1(n14590), .A2(n20064), .ZN(n14184) );
  INV_X1 U17462 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14222) );
  NOR2_X1 U17463 ( .A1(n20066), .A2(n14222), .ZN(n14593) );
  NOR2_X1 U17464 ( .A1(n15984), .A2(n14181), .ZN(n14182) );
  AOI211_X1 U17465 ( .C1(n15979), .C2(n14224), .A(n14593), .B(n14182), .ZN(
        n14183) );
  OAI211_X1 U17466 ( .C1(n14220), .C2(n20106), .A(n14184), .B(n14183), .ZN(
        P1_U2969) );
  AOI22_X1 U17467 ( .A1(n14421), .A2(BUF1_REG_30__SCAN_IN), .B1(
        P1_EAX_REG_30__SCAN_IN), .B2(n14428), .ZN(n14188) );
  AOI22_X1 U17468 ( .A1(n14424), .A2(n14186), .B1(n14422), .B2(DATAI_30_), 
        .ZN(n14187) );
  OAI211_X1 U17469 ( .C1(n14220), .C2(n14431), .A(n14188), .B(n14187), .ZN(
        P1_U2874) );
  NAND2_X1 U17470 ( .A1(n14204), .A2(n14191), .ZN(n14190) );
  NAND2_X1 U17471 ( .A1(n14190), .A2(n14189), .ZN(n14193) );
  OR2_X1 U17472 ( .A1(n14248), .A2(n14191), .ZN(n14192) );
  NAND2_X1 U17473 ( .A1(n14193), .A2(n14192), .ZN(n14195) );
  AND2_X1 U17474 ( .A1(n14206), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14194) );
  AOI21_X1 U17475 ( .B1(n14207), .B2(P1_EBX_REG_30__SCAN_IN), .A(n14194), .ZN(
        n14205) );
  XNOR2_X1 U17476 ( .A(n14195), .B(n14205), .ZN(n14598) );
  INV_X1 U17477 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14227) );
  OAI222_X1 U17478 ( .A1(n14359), .A2(n14220), .B1(n20002), .B2(n14598), .C1(
        n14227), .C2(n14350), .ZN(P1_U2842) );
  NAND2_X1 U17479 ( .A1(n16053), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14583) );
  NAND2_X1 U17480 ( .A1(n20060), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14197) );
  OAI211_X1 U17481 ( .C1(n15978), .C2(n14198), .A(n14583), .B(n14197), .ZN(
        n14199) );
  AOI21_X1 U17482 ( .B1(n14210), .B2(n15975), .A(n14199), .ZN(n14200) );
  OAI21_X1 U17483 ( .B1(n14589), .B2(n15962), .A(n14200), .ZN(P1_U2968) );
  NOR2_X1 U17484 ( .A1(n15270), .A2(n13257), .ZN(n14201) );
  AOI21_X1 U17485 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n13257), .A(n14201), .ZN(
        n14202) );
  OAI21_X1 U17486 ( .B1(n14203), .B2(n14966), .A(n14202), .ZN(P2_U2857) );
  MUX2_X1 U17487 ( .A(n14205), .B(n11879), .S(n14204), .Z(n14209) );
  AOI22_X1 U17488 ( .A1(n14207), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n14206), .ZN(n14208) );
  NAND2_X1 U17489 ( .A1(n14210), .A2(n19932), .ZN(n14219) );
  AND2_X1 U17490 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n14212) );
  INV_X1 U17491 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n14472) );
  INV_X1 U17492 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n14294) );
  INV_X1 U17493 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20686) );
  INV_X1 U17494 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n20676) );
  NAND2_X1 U17495 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n14298) );
  NAND4_X1 U17496 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(P1_REIP_REG_12__SCAN_IN), 
        .A3(P1_REIP_REG_13__SCAN_IN), .A4(P1_REIP_REG_14__SCAN_IN), .ZN(n15859) );
  NAND2_X1 U17497 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n15858) );
  NOR4_X1 U17498 ( .A1(n20676), .A2(n14298), .A3(n15859), .A4(n15858), .ZN(
        n15829) );
  NAND4_X1 U17499 ( .A1(n15826), .A2(n15829), .A3(P1_REIP_REG_19__SCAN_IN), 
        .A4(P1_REIP_REG_18__SCAN_IN), .ZN(n15783) );
  NAND3_X1 U17500 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .A3(P1_REIP_REG_20__SCAN_IN), .ZN(n15784) );
  NOR3_X1 U17501 ( .A1(n20686), .A2(n15783), .A3(n15784), .ZN(n15773) );
  NAND2_X1 U17502 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n15773), .ZN(n14286) );
  OR2_X1 U17503 ( .A1(n14294), .A2(n14286), .ZN(n14274) );
  NOR3_X1 U17504 ( .A1(n14472), .A2(n14274), .A3(n19967), .ZN(n14259) );
  AND3_X1 U17505 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .A3(n14259), .ZN(n14211) );
  OR2_X1 U17506 ( .A1(n19929), .A2(n14211), .ZN(n14243) );
  OAI21_X1 U17507 ( .B1(n19929), .B2(n14212), .A(n14243), .ZN(n14230) );
  INV_X1 U17508 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14305) );
  NAND2_X1 U17509 ( .A1(n19991), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14216) );
  NAND2_X1 U17510 ( .A1(n19982), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14213) );
  NOR2_X1 U17511 ( .A1(n14274), .A2(n14213), .ZN(n14261) );
  AND3_X1 U17512 ( .A1(n14261), .A2(P1_REIP_REG_27__SCAN_IN), .A3(
        P1_REIP_REG_28__SCAN_IN), .ZN(n14234) );
  INV_X1 U17513 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n14214) );
  NAND4_X1 U17514 ( .A1(n14234), .A2(P1_REIP_REG_29__SCAN_IN), .A3(
        P1_REIP_REG_30__SCAN_IN), .A4(n14214), .ZN(n14215) );
  OAI211_X1 U17515 ( .C1(n14305), .C2(n19986), .A(n14216), .B(n14215), .ZN(
        n14217) );
  AOI21_X1 U17516 ( .B1(n14230), .B2(P1_REIP_REG_31__SCAN_IN), .A(n14217), 
        .ZN(n14218) );
  OAI211_X1 U17517 ( .C1(n14588), .C2(n19987), .A(n14219), .B(n14218), .ZN(
        P1_U2809) );
  INV_X1 U17518 ( .A(n14220), .ZN(n14221) );
  NAND2_X1 U17519 ( .A1(n14221), .A2(n19932), .ZN(n14232) );
  NAND2_X1 U17520 ( .A1(n14234), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14223) );
  NAND2_X1 U17521 ( .A1(n14223), .A2(n14222), .ZN(n14229) );
  NAND2_X1 U17522 ( .A1(n19993), .A2(n14224), .ZN(n14226) );
  NAND2_X1 U17523 ( .A1(n19991), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14225) );
  OAI211_X1 U17524 ( .C1(n19986), .C2(n14227), .A(n14226), .B(n14225), .ZN(
        n14228) );
  AOI21_X1 U17525 ( .B1(n14230), .B2(n14229), .A(n14228), .ZN(n14231) );
  OAI211_X1 U17526 ( .C1(n14598), .C2(n19987), .A(n14232), .B(n14231), .ZN(
        P1_U2810) );
  NAND2_X1 U17527 ( .A1(n14441), .A2(n19932), .ZN(n14239) );
  INV_X1 U17528 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n14233) );
  NOR2_X1 U17529 ( .A1(n14243), .A2(n14233), .ZN(n14237) );
  INV_X1 U17530 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14439) );
  AOI22_X1 U17531 ( .A1(n14234), .A2(n14233), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n19971), .ZN(n14235) );
  OAI21_X1 U17532 ( .B1(n19956), .B2(n14439), .A(n14235), .ZN(n14236) );
  AOI211_X1 U17533 ( .C1(n19993), .C2(n14437), .A(n14237), .B(n14236), .ZN(
        n14238) );
  OAI211_X1 U17534 ( .C1(n19987), .C2(n14599), .A(n14239), .B(n14238), .ZN(
        P1_U2811) );
  AOI21_X1 U17535 ( .B1(n14242), .B2(n14257), .A(n11722), .ZN(n14457) );
  INV_X1 U17536 ( .A(n14457), .ZN(n14371) );
  INV_X1 U17537 ( .A(n14243), .ZN(n14253) );
  INV_X1 U17538 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14306) );
  INV_X1 U17539 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14244) );
  NAND3_X1 U17540 ( .A1(n14261), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14244), 
        .ZN(n14245) );
  OAI21_X1 U17541 ( .B1(n14306), .B2(n19986), .A(n14245), .ZN(n14246) );
  AOI21_X1 U17542 ( .B1(n19991), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14246), .ZN(n14247) );
  OAI21_X1 U17543 ( .B1(n19965), .B2(n14455), .A(n14247), .ZN(n14252) );
  INV_X1 U17544 ( .A(n14248), .ZN(n14249) );
  OAI21_X1 U17545 ( .B1(n14250), .B2(n14265), .A(n14249), .ZN(n14612) );
  NOR2_X1 U17546 ( .A1(n14612), .A2(n19987), .ZN(n14251) );
  AOI211_X1 U17547 ( .C1(n14253), .C2(P1_REIP_REG_28__SCAN_IN), .A(n14252), 
        .B(n14251), .ZN(n14254) );
  OAI21_X1 U17548 ( .B1(n14371), .B2(n15894), .A(n14254), .ZN(P1_U2812) );
  NOR2_X1 U17549 ( .A1(n19929), .A2(n14259), .ZN(n14278) );
  INV_X1 U17550 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14464) );
  INV_X1 U17551 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n14260) );
  AOI22_X1 U17552 ( .A1(n14261), .A2(n14260), .B1(P1_EBX_REG_27__SCAN_IN), 
        .B2(n19971), .ZN(n14263) );
  NAND2_X1 U17553 ( .A1(n19993), .A2(n14468), .ZN(n14262) );
  OAI211_X1 U17554 ( .C1(n19956), .C2(n14464), .A(n14263), .B(n14262), .ZN(
        n14264) );
  AOI21_X1 U17555 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n14278), .A(n14264), 
        .ZN(n14268) );
  AOI21_X1 U17556 ( .B1(n14266), .B2(n14272), .A(n14265), .ZN(n14622) );
  NAND2_X1 U17557 ( .A1(n14622), .A2(n19959), .ZN(n14267) );
  OAI211_X1 U17558 ( .C1(n14465), .C2(n15894), .A(n14268), .B(n14267), .ZN(
        P1_U2813) );
  AOI21_X1 U17559 ( .B1(n14270), .B2(n14269), .A(n14256), .ZN(n14476) );
  INV_X1 U17560 ( .A(n14476), .ZN(n14378) );
  AOI21_X1 U17561 ( .B1(n14273), .B2(n14271), .A(n9953), .ZN(n14629) );
  NOR3_X1 U17562 ( .A1(n14274), .A2(P1_REIP_REG_26__SCAN_IN), .A3(n19969), 
        .ZN(n14277) );
  NOR2_X1 U17563 ( .A1(n19956), .A2(n14275), .ZN(n14276) );
  AOI211_X1 U17564 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n19971), .A(n14277), .B(
        n14276), .ZN(n14280) );
  NAND2_X1 U17565 ( .A1(n14278), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14279) );
  OAI211_X1 U17566 ( .C1(n19965), .C2(n14474), .A(n14280), .B(n14279), .ZN(
        n14281) );
  AOI21_X1 U17567 ( .B1(n14629), .B2(n19959), .A(n14281), .ZN(n14282) );
  OAI21_X1 U17568 ( .B1(n14378), .B2(n15894), .A(n14282), .ZN(P1_U2814) );
  NAND2_X1 U17569 ( .A1(n14312), .A2(n14284), .ZN(n14285) );
  NAND2_X1 U17570 ( .A1(n14269), .A2(n14285), .ZN(n14484) );
  NOR2_X1 U17571 ( .A1(n19969), .A2(n14286), .ZN(n14295) );
  INV_X1 U17572 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14483) );
  OR2_X1 U17573 ( .A1(n15773), .A2(n19969), .ZN(n14287) );
  AND2_X1 U17574 ( .A1(n19927), .A2(n14287), .ZN(n15785) );
  OAI21_X1 U17575 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n19969), .A(n15785), 
        .ZN(n14288) );
  AOI22_X1 U17576 ( .A1(n19971), .A2(P1_EBX_REG_25__SCAN_IN), .B1(n14288), 
        .B2(P1_REIP_REG_25__SCAN_IN), .ZN(n14290) );
  NAND2_X1 U17577 ( .A1(n19993), .A2(n14487), .ZN(n14289) );
  OAI211_X1 U17578 ( .C1(n19956), .C2(n14483), .A(n14290), .B(n14289), .ZN(
        n14293) );
  OAI21_X1 U17579 ( .B1(n14314), .B2(n14291), .A(n14271), .ZN(n14309) );
  NOR2_X1 U17580 ( .A1(n14309), .A2(n19987), .ZN(n14292) );
  AOI211_X1 U17581 ( .C1(n14295), .C2(n14294), .A(n14293), .B(n14292), .ZN(
        n14296) );
  OAI21_X1 U17582 ( .B1(n14484), .B2(n15894), .A(n14296), .ZN(P1_U2815) );
  INV_X1 U17583 ( .A(n14556), .ZN(n14432) );
  INV_X1 U17584 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n15888) );
  INV_X1 U17585 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n20668) );
  NAND3_X1 U17586 ( .A1(n19982), .A2(n15826), .A3(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n15905) );
  NOR2_X1 U17587 ( .A1(n20668), .A2(n15905), .ZN(n15899) );
  NAND2_X1 U17588 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n15899), .ZN(n15887) );
  NOR2_X1 U17589 ( .A1(n15888), .A2(n15887), .ZN(n15879) );
  INV_X1 U17590 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n20819) );
  INV_X1 U17591 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n20840) );
  NOR2_X1 U17592 ( .A1(n20840), .A2(n15888), .ZN(n14299) );
  AOI21_X1 U17593 ( .B1(n19982), .B2(n14298), .A(n14297), .ZN(n15913) );
  OAI21_X1 U17594 ( .B1(n14299), .B2(n19929), .A(n15913), .ZN(n15890) );
  AOI21_X1 U17595 ( .B1(n19991), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n19925), .ZN(n14302) );
  INV_X1 U17596 ( .A(n14554), .ZN(n14300) );
  AOI22_X1 U17597 ( .A1(n19993), .A2(n14300), .B1(n19971), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14301) );
  OAI211_X1 U17598 ( .C1(n19987), .C2(n14694), .A(n14302), .B(n14301), .ZN(
        n14303) );
  AOI221_X1 U17599 ( .B1(n15879), .B2(n20819), .C1(n15890), .C2(
        P1_REIP_REG_13__SCAN_IN), .A(n14303), .ZN(n14304) );
  OAI21_X1 U17600 ( .B1(n14432), .B2(n15894), .A(n14304), .ZN(P1_U2827) );
  OAI22_X1 U17601 ( .A1(n14588), .A2(n20002), .B1(n14305), .B2(n14350), .ZN(
        P1_U2841) );
  OAI222_X1 U17602 ( .A1(n14306), .A2(n14350), .B1(n20002), .B2(n14612), .C1(
        n14371), .C2(n14359), .ZN(P1_U2844) );
  AOI22_X1 U17603 ( .A1(n14622), .A2(n11892), .B1(n14337), .B2(
        P1_EBX_REG_27__SCAN_IN), .ZN(n14307) );
  OAI21_X1 U17604 ( .B1(n14465), .B2(n14359), .A(n14307), .ZN(P1_U2845) );
  AOI22_X1 U17605 ( .A1(n14629), .A2(n11892), .B1(n14337), .B2(
        P1_EBX_REG_26__SCAN_IN), .ZN(n14308) );
  OAI21_X1 U17606 ( .B1(n14378), .B2(n14359), .A(n14308), .ZN(P1_U2846) );
  INV_X1 U17607 ( .A(n14309), .ZN(n14638) );
  AOI22_X1 U17608 ( .A1(n14638), .A2(n11892), .B1(n14337), .B2(
        P1_EBX_REG_25__SCAN_IN), .ZN(n14310) );
  OAI21_X1 U17609 ( .B1(n14484), .B2(n14359), .A(n14310), .ZN(P1_U2847) );
  AOI21_X1 U17610 ( .B1(n14313), .B2(n14311), .A(n14283), .ZN(n15779) );
  INV_X1 U17611 ( .A(n15779), .ZN(n14387) );
  AOI21_X1 U17612 ( .B1(n14315), .B2(n14319), .A(n14314), .ZN(n15778) );
  AOI22_X1 U17613 ( .A1(n15778), .A2(n11892), .B1(n14337), .B2(
        P1_EBX_REG_24__SCAN_IN), .ZN(n14316) );
  OAI21_X1 U17614 ( .B1(n14387), .B2(n14359), .A(n14316), .ZN(P1_U2848) );
  OAI21_X1 U17615 ( .B1(n14317), .B2(n14318), .A(n14311), .ZN(n15790) );
  AOI21_X1 U17616 ( .B1(n14320), .B2(n9772), .A(n9959), .ZN(n15788) );
  AOI22_X1 U17617 ( .A1(n15788), .A2(n11892), .B1(n14337), .B2(
        P1_EBX_REG_23__SCAN_IN), .ZN(n14321) );
  OAI21_X1 U17618 ( .B1(n15790), .B2(n14359), .A(n14321), .ZN(P1_U2849) );
  INV_X1 U17619 ( .A(n14322), .ZN(n14392) );
  NAND2_X1 U17620 ( .A1(n14323), .A2(n14324), .ZN(n14325) );
  AND2_X1 U17621 ( .A1(n14392), .A2(n14325), .ZN(n15814) );
  INV_X1 U17622 ( .A(n15814), .ZN(n14401) );
  INV_X1 U17623 ( .A(n14660), .ZN(n14328) );
  NAND2_X1 U17624 ( .A1(n14334), .A2(n14326), .ZN(n14327) );
  NAND2_X1 U17625 ( .A1(n14328), .A2(n14327), .ZN(n15817) );
  OAI22_X1 U17626 ( .A1(n15817), .A2(n20002), .B1(n15809), .B2(n14350), .ZN(
        n14329) );
  INV_X1 U17627 ( .A(n14329), .ZN(n14330) );
  OAI21_X1 U17628 ( .B1(n14401), .B2(n14359), .A(n14330), .ZN(P1_U2851) );
  OAI21_X1 U17629 ( .B1(n14332), .B2(n14333), .A(n14323), .ZN(n15922) );
  INV_X1 U17630 ( .A(n14334), .ZN(n14335) );
  AOI21_X1 U17631 ( .B1(n14336), .B2(n14344), .A(n14335), .ZN(n15823) );
  AOI22_X1 U17632 ( .A1(n15823), .A2(n11892), .B1(n14337), .B2(
        P1_EBX_REG_20__SCAN_IN), .ZN(n14338) );
  OAI21_X1 U17633 ( .B1(n15922), .B2(n14359), .A(n14338), .ZN(P1_U2852) );
  INV_X1 U17634 ( .A(n14332), .ZN(n14340) );
  OAI21_X1 U17635 ( .B1(n14341), .B2(n14339), .A(n14340), .ZN(n15835) );
  NAND2_X1 U17636 ( .A1(n15843), .A2(n14342), .ZN(n14343) );
  NAND2_X1 U17637 ( .A1(n14344), .A2(n14343), .ZN(n15839) );
  OAI222_X1 U17638 ( .A1(n14359), .A2(n15835), .B1(n14350), .B2(n11852), .C1(
        n15839), .C2(n20002), .ZN(P1_U2853) );
  AOI21_X1 U17639 ( .B1(n14346), .B2(n9821), .A(n10039), .ZN(n15854) );
  NOR2_X1 U17640 ( .A1(n9839), .A2(n14348), .ZN(n14349) );
  OR2_X1 U17641 ( .A1(n14347), .A2(n14349), .ZN(n15857) );
  OAI22_X1 U17642 ( .A1(n15857), .A2(n20002), .B1(n15848), .B2(n14350), .ZN(
        n14351) );
  AOI21_X1 U17643 ( .B1(n15854), .B2(n20004), .A(n14351), .ZN(n14352) );
  INV_X1 U17644 ( .A(n14352), .ZN(P1_U2855) );
  AOI21_X1 U17645 ( .B1(n14355), .B2(n14354), .A(n14353), .ZN(n14356) );
  NOR2_X1 U17646 ( .A1(n14356), .A2(n9839), .ZN(n15996) );
  INV_X1 U17647 ( .A(n15996), .ZN(n14360) );
  INV_X1 U17648 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n15863) );
  NAND2_X1 U17649 ( .A1(n14058), .A2(n14357), .ZN(n14358) );
  AND2_X1 U17650 ( .A1(n9821), .A2(n14358), .ZN(n15939) );
  INV_X1 U17651 ( .A(n15939), .ZN(n14427) );
  OAI222_X1 U17652 ( .A1(n14360), .A2(n20002), .B1(n15863), .B2(n14350), .C1(
        n14427), .C2(n14359), .ZN(P1_U2856) );
  AOI22_X1 U17653 ( .A1(n14421), .A2(BUF1_REG_29__SCAN_IN), .B1(
        P1_EAX_REG_29__SCAN_IN), .B2(n14428), .ZN(n14364) );
  INV_X1 U17654 ( .A(DATAI_13_), .ZN(n14362) );
  NAND2_X1 U17655 ( .A1(n20107), .A2(BUF1_REG_13__SCAN_IN), .ZN(n14361) );
  OAI21_X1 U17656 ( .B1(n20107), .B2(n14362), .A(n14361), .ZN(n20042) );
  AOI22_X1 U17657 ( .A1(n14424), .A2(n20042), .B1(n14422), .B2(DATAI_29_), 
        .ZN(n14363) );
  OAI211_X1 U17658 ( .C1(n14365), .C2(n14431), .A(n14364), .B(n14363), .ZN(
        P1_U2875) );
  INV_X1 U17659 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n19233) );
  OAI22_X1 U17660 ( .A1(n14411), .A2(n19233), .B1(n14366), .B2(n14409), .ZN(
        n14367) );
  INV_X1 U17661 ( .A(n14367), .ZN(n14370) );
  AOI22_X1 U17662 ( .A1(n14424), .A2(n14368), .B1(n14422), .B2(DATAI_28_), 
        .ZN(n14369) );
  OAI211_X1 U17663 ( .C1(n14371), .C2(n14431), .A(n14370), .B(n14369), .ZN(
        P1_U2876) );
  AOI22_X1 U17664 ( .A1(n14421), .A2(BUF1_REG_27__SCAN_IN), .B1(
        P1_EAX_REG_27__SCAN_IN), .B2(n14428), .ZN(n14373) );
  AOI22_X1 U17665 ( .A1(n14424), .A2(n20040), .B1(n14422), .B2(DATAI_27_), 
        .ZN(n14372) );
  OAI211_X1 U17666 ( .C1(n14465), .C2(n14431), .A(n14373), .B(n14372), .ZN(
        P1_U2877) );
  INV_X1 U17667 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16360) );
  OAI22_X1 U17668 ( .A1(n14411), .A2(n16360), .B1(n14374), .B2(n14409), .ZN(
        n14375) );
  INV_X1 U17669 ( .A(n14375), .ZN(n14377) );
  AOI22_X1 U17670 ( .A1(n14424), .A2(n20038), .B1(n14422), .B2(DATAI_26_), 
        .ZN(n14376) );
  OAI211_X1 U17671 ( .C1(n14378), .C2(n14431), .A(n14377), .B(n14376), .ZN(
        P1_U2878) );
  AOI22_X1 U17672 ( .A1(n14421), .A2(BUF1_REG_25__SCAN_IN), .B1(
        P1_EAX_REG_25__SCAN_IN), .B2(n14428), .ZN(n14380) );
  AOI22_X1 U17673 ( .A1(n14424), .A2(n20036), .B1(n14422), .B2(DATAI_25_), 
        .ZN(n14379) );
  OAI211_X1 U17674 ( .C1(n14484), .C2(n14431), .A(n14380), .B(n14379), .ZN(
        P1_U2879) );
  INV_X1 U17675 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n14382) );
  OAI22_X1 U17676 ( .A1(n14411), .A2(n14382), .B1(n14381), .B2(n14409), .ZN(
        n14383) );
  INV_X1 U17677 ( .A(n14383), .ZN(n14386) );
  AOI22_X1 U17678 ( .A1(n14424), .A2(n14384), .B1(n14422), .B2(DATAI_24_), 
        .ZN(n14385) );
  OAI211_X1 U17679 ( .C1(n14387), .C2(n14431), .A(n14386), .B(n14385), .ZN(
        P1_U2880) );
  AOI22_X1 U17680 ( .A1(n14421), .A2(BUF1_REG_23__SCAN_IN), .B1(
        P1_EAX_REG_23__SCAN_IN), .B2(n14428), .ZN(n14390) );
  AOI22_X1 U17681 ( .A1(n14424), .A2(n14388), .B1(n14422), .B2(DATAI_23_), 
        .ZN(n14389) );
  OAI211_X1 U17682 ( .C1(n15790), .C2(n14431), .A(n14390), .B(n14389), .ZN(
        P1_U2881) );
  AND2_X1 U17683 ( .A1(n14392), .A2(n14391), .ZN(n14393) );
  OR2_X1 U17684 ( .A1(n14393), .A2(n14317), .ZN(n15915) );
  OAI22_X1 U17685 ( .A1(n14411), .A2(n15002), .B1(n14394), .B2(n14409), .ZN(
        n14396) );
  INV_X1 U17686 ( .A(n14424), .ZN(n14412) );
  NOR2_X1 U17687 ( .A1(n14412), .A2(n20143), .ZN(n14395) );
  AOI211_X1 U17688 ( .C1(n14422), .C2(DATAI_22_), .A(n14396), .B(n14395), .ZN(
        n14397) );
  OAI21_X1 U17689 ( .B1(n15915), .B2(n14431), .A(n14397), .ZN(P1_U2882) );
  AOI22_X1 U17690 ( .A1(n14421), .A2(BUF1_REG_21__SCAN_IN), .B1(
        P1_EAX_REG_21__SCAN_IN), .B2(n14428), .ZN(n14400) );
  AOI22_X1 U17691 ( .A1(n14424), .A2(n14398), .B1(n14422), .B2(DATAI_21_), 
        .ZN(n14399) );
  OAI211_X1 U17692 ( .C1(n14401), .C2(n14431), .A(n14400), .B(n14399), .ZN(
        P1_U2883) );
  AOI22_X1 U17693 ( .A1(n14421), .A2(BUF1_REG_20__SCAN_IN), .B1(
        P1_EAX_REG_20__SCAN_IN), .B2(n14428), .ZN(n14404) );
  AOI22_X1 U17694 ( .A1(n14424), .A2(n14402), .B1(n14422), .B2(DATAI_20_), 
        .ZN(n14403) );
  OAI211_X1 U17695 ( .C1(n15922), .C2(n14431), .A(n14404), .B(n14403), .ZN(
        P1_U2884) );
  AOI22_X1 U17696 ( .A1(n14421), .A2(BUF1_REG_19__SCAN_IN), .B1(
        P1_EAX_REG_19__SCAN_IN), .B2(n14428), .ZN(n14407) );
  AOI22_X1 U17697 ( .A1(n14424), .A2(n14405), .B1(n14422), .B2(DATAI_19_), 
        .ZN(n14406) );
  OAI211_X1 U17698 ( .C1(n15835), .C2(n14431), .A(n14407), .B(n14406), .ZN(
        P1_U2885) );
  AOI21_X1 U17699 ( .B1(n14408), .B2(n14345), .A(n14339), .ZN(n15930) );
  INV_X1 U17700 ( .A(n15930), .ZN(n14416) );
  INV_X1 U17701 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16371) );
  OAI22_X1 U17702 ( .A1(n14411), .A2(n16371), .B1(n14410), .B2(n14409), .ZN(
        n14414) );
  NOR2_X1 U17703 ( .A1(n14412), .A2(n20124), .ZN(n14413) );
  AOI211_X1 U17704 ( .C1(n14422), .C2(DATAI_18_), .A(n14414), .B(n14413), .ZN(
        n14415) );
  OAI21_X1 U17705 ( .B1(n14416), .B2(n14431), .A(n14415), .ZN(P1_U2886) );
  INV_X1 U17706 ( .A(n15854), .ZN(n14420) );
  AOI22_X1 U17707 ( .A1(n14421), .A2(BUF1_REG_17__SCAN_IN), .B1(
        P1_EAX_REG_17__SCAN_IN), .B2(n14428), .ZN(n14419) );
  AOI22_X1 U17708 ( .A1(n14424), .A2(n14417), .B1(n14422), .B2(DATAI_17_), 
        .ZN(n14418) );
  OAI211_X1 U17709 ( .C1(n14420), .C2(n14431), .A(n14419), .B(n14418), .ZN(
        P1_U2887) );
  AOI22_X1 U17710 ( .A1(n14421), .A2(BUF1_REG_16__SCAN_IN), .B1(
        P1_EAX_REG_16__SCAN_IN), .B2(n14428), .ZN(n14426) );
  AOI22_X1 U17711 ( .A1(n14424), .A2(n14423), .B1(n14422), .B2(DATAI_16_), 
        .ZN(n14425) );
  OAI211_X1 U17712 ( .C1(n14427), .C2(n14431), .A(n14426), .B(n14425), .ZN(
        P1_U2888) );
  AOI22_X1 U17713 ( .A1(n14429), .A2(n20042), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14428), .ZN(n14430) );
  OAI21_X1 U17714 ( .B1(n14432), .B2(n14431), .A(n14430), .ZN(P1_U2891) );
  INV_X1 U17715 ( .A(n14433), .ZN(n14435) );
  OAI21_X1 U17716 ( .B1(n14435), .B2(n14545), .A(n14434), .ZN(n14436) );
  XNOR2_X1 U17717 ( .A(n14436), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14605) );
  NAND2_X1 U17718 ( .A1(n15979), .A2(n14437), .ZN(n14438) );
  NAND2_X1 U17719 ( .A1(n16053), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14601) );
  OAI211_X1 U17720 ( .C1(n15984), .C2(n14439), .A(n14438), .B(n14601), .ZN(
        n14440) );
  AOI21_X1 U17721 ( .B1(n14441), .B2(n15975), .A(n14440), .ZN(n14442) );
  OAI21_X1 U17722 ( .B1(n14605), .B2(n15962), .A(n14442), .ZN(P1_U2970) );
  INV_X1 U17723 ( .A(n14444), .ZN(n14625) );
  NAND2_X1 U17724 ( .A1(n14160), .A2(n14625), .ZN(n14445) );
  NAND2_X1 U17725 ( .A1(n14443), .A2(n14445), .ZN(n14450) );
  NAND2_X1 U17726 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14446) );
  NOR2_X1 U17727 ( .A1(n14450), .A2(n14446), .ZN(n14452) );
  NAND2_X1 U17728 ( .A1(n14571), .A2(n14462), .ZN(n14447) );
  NOR2_X1 U17729 ( .A1(n14448), .A2(n14447), .ZN(n14449) );
  AND2_X1 U17730 ( .A1(n14450), .A2(n14449), .ZN(n14451) );
  MUX2_X1 U17731 ( .A(n14452), .B(n14451), .S(n14545), .Z(n14453) );
  XNOR2_X1 U17732 ( .A(n14453), .B(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14616) );
  NAND2_X1 U17733 ( .A1(n16053), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14606) );
  NAND2_X1 U17734 ( .A1(n20060), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14454) );
  OAI211_X1 U17735 ( .C1(n15978), .C2(n14455), .A(n14606), .B(n14454), .ZN(
        n14456) );
  AOI21_X1 U17736 ( .B1(n14457), .B2(n15975), .A(n14456), .ZN(n14458) );
  OAI21_X1 U17737 ( .B1(n15962), .B2(n14616), .A(n14458), .ZN(P1_U2971) );
  NAND2_X1 U17738 ( .A1(n14459), .A2(n9773), .ZN(n14460) );
  MUX2_X1 U17739 ( .A(n14461), .B(n14460), .S(n14545), .Z(n14463) );
  XNOR2_X1 U17740 ( .A(n14463), .B(n14462), .ZN(n14624) );
  NAND2_X1 U17741 ( .A1(n16053), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14618) );
  OAI21_X1 U17742 ( .B1(n15984), .B2(n14464), .A(n14618), .ZN(n14467) );
  NOR2_X1 U17743 ( .A1(n14465), .A2(n20106), .ZN(n14466) );
  AOI211_X1 U17744 ( .C1(n15979), .C2(n14468), .A(n14467), .B(n14466), .ZN(
        n14469) );
  OAI21_X1 U17745 ( .B1(n15962), .B2(n14624), .A(n14469), .ZN(P1_U2972) );
  INV_X1 U17746 ( .A(n14443), .ZN(n14489) );
  NOR2_X1 U17747 ( .A1(n14489), .A2(n14625), .ZN(n14470) );
  MUX2_X1 U17748 ( .A(n9773), .B(n14470), .S(n14160), .Z(n14471) );
  XNOR2_X1 U17749 ( .A(n14471), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14632) );
  NOR2_X1 U17750 ( .A1(n20066), .A2(n14472), .ZN(n14627) );
  AOI21_X1 U17751 ( .B1(n20060), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n14627), .ZN(n14473) );
  OAI21_X1 U17752 ( .B1(n15978), .B2(n14474), .A(n14473), .ZN(n14475) );
  AOI21_X1 U17753 ( .B1(n14476), .B2(n15975), .A(n14475), .ZN(n14477) );
  OAI21_X1 U17754 ( .B1(n15962), .B2(n14632), .A(n14477), .ZN(P1_U2973) );
  NAND3_X1 U17755 ( .A1(n14489), .A2(n20956), .A3(n14643), .ZN(n14481) );
  NAND2_X1 U17756 ( .A1(n14490), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14480) );
  MUX2_X1 U17757 ( .A(n14481), .B(n14480), .S(n14160), .Z(n14482) );
  XNOR2_X1 U17758 ( .A(n14482), .B(n14635), .ZN(n14640) );
  NAND2_X1 U17759 ( .A1(n16053), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14634) );
  OAI21_X1 U17760 ( .B1(n15984), .B2(n14483), .A(n14634), .ZN(n14486) );
  NOR2_X1 U17761 ( .A1(n14484), .A2(n20106), .ZN(n14485) );
  AOI211_X1 U17762 ( .C1(n15979), .C2(n14487), .A(n14486), .B(n14485), .ZN(
        n14488) );
  OAI21_X1 U17763 ( .B1(n14640), .B2(n15962), .A(n14488), .ZN(P1_U2974) );
  NAND2_X1 U17764 ( .A1(n14489), .A2(n14545), .ZN(n14491) );
  MUX2_X1 U17765 ( .A(n14491), .B(n14545), .S(n14490), .Z(n14492) );
  XNOR2_X1 U17766 ( .A(n14492), .B(n14643), .ZN(n14650) );
  NAND2_X1 U17767 ( .A1(n16053), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14645) );
  NAND2_X1 U17768 ( .A1(n20060), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14493) );
  OAI211_X1 U17769 ( .C1(n15978), .C2(n15782), .A(n14645), .B(n14493), .ZN(
        n14494) );
  AOI21_X1 U17770 ( .B1(n15779), .B2(n15975), .A(n14494), .ZN(n14495) );
  OAI21_X1 U17771 ( .B1(n14650), .B2(n15962), .A(n14495), .ZN(P1_U2975) );
  XNOR2_X1 U17772 ( .A(n14160), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14496) );
  XNOR2_X1 U17773 ( .A(n14443), .B(n14496), .ZN(n14657) );
  NAND2_X1 U17774 ( .A1(n16053), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14651) );
  OAI21_X1 U17775 ( .B1(n15984), .B2(n15795), .A(n14651), .ZN(n14498) );
  NOR2_X1 U17776 ( .A1(n15790), .A2(n20106), .ZN(n14497) );
  AOI211_X1 U17777 ( .C1(n15979), .C2(n15792), .A(n14498), .B(n14497), .ZN(
        n14499) );
  OAI21_X1 U17778 ( .B1(n14657), .B2(n15962), .A(n14499), .ZN(P1_U2976) );
  NAND2_X1 U17779 ( .A1(n14501), .A2(n14500), .ZN(n14502) );
  XNOR2_X1 U17780 ( .A(n14502), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14658) );
  NAND2_X1 U17781 ( .A1(n14658), .A2(n20064), .ZN(n14506) );
  INV_X1 U17782 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n14503) );
  NOR2_X1 U17783 ( .A1(n20066), .A2(n14503), .ZN(n14662) );
  NOR2_X1 U17784 ( .A1(n15978), .A2(n15807), .ZN(n14504) );
  AOI211_X1 U17785 ( .C1(n20060), .C2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n14662), .B(n14504), .ZN(n14505) );
  OAI211_X1 U17786 ( .C1(n20106), .C2(n15915), .A(n14506), .B(n14505), .ZN(
        P1_U2977) );
  NAND2_X1 U17787 ( .A1(n14507), .A2(n15749), .ZN(n14510) );
  OAI21_X1 U17788 ( .B1(n14508), .B2(n14545), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14509) );
  OAI211_X1 U17789 ( .C1(n14545), .C2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n14510), .B(n14509), .ZN(n14511) );
  XNOR2_X1 U17790 ( .A(n14511), .B(n14675), .ZN(n14678) );
  AOI22_X1 U17791 ( .A1(n20060), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n16053), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n14512) );
  OAI21_X1 U17792 ( .B1(n15978), .B2(n15812), .A(n14512), .ZN(n14513) );
  AOI21_X1 U17793 ( .B1(n15814), .B2(n15975), .A(n14513), .ZN(n14514) );
  OAI21_X1 U17794 ( .B1(n14678), .B2(n15962), .A(n14514), .ZN(P1_U2978) );
  NOR2_X1 U17795 ( .A1(n14160), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14515) );
  MUX2_X1 U17796 ( .A(n14160), .B(n14515), .S(n14508), .Z(n14516) );
  XNOR2_X1 U17797 ( .A(n14516), .B(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14684) );
  INV_X1 U17798 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n14517) );
  OR2_X1 U17799 ( .A1(n20066), .A2(n14517), .ZN(n14681) );
  OAI21_X1 U17800 ( .B1(n15984), .B2(n15831), .A(n14681), .ZN(n14519) );
  NOR2_X1 U17801 ( .A1(n15835), .A2(n20106), .ZN(n14518) );
  AOI211_X1 U17802 ( .C1(n15979), .C2(n15837), .A(n14519), .B(n14518), .ZN(
        n14520) );
  OAI21_X1 U17803 ( .B1(n15962), .B2(n14684), .A(n14520), .ZN(P1_U2980) );
  NAND2_X1 U17804 ( .A1(n14545), .A2(n14521), .ZN(n14526) );
  AOI21_X1 U17805 ( .B1(n14522), .B2(n14524), .A(n14523), .ZN(n14525) );
  MUX2_X1 U17806 ( .A(n14526), .B(n14545), .S(n14525), .Z(n14527) );
  XNOR2_X1 U17807 ( .A(n14527), .B(n14688), .ZN(n14693) );
  INV_X1 U17808 ( .A(n15851), .ZN(n14529) );
  AOI22_X1 U17809 ( .A1(n20060), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n16053), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n14528) );
  OAI21_X1 U17810 ( .B1(n15978), .B2(n14529), .A(n14528), .ZN(n14530) );
  AOI21_X1 U17811 ( .B1(n15854), .B2(n15975), .A(n14530), .ZN(n14531) );
  OAI21_X1 U17812 ( .B1(n14693), .B2(n15962), .A(n14531), .ZN(P1_U2982) );
  AND2_X1 U17813 ( .A1(n14522), .A2(n14532), .ZN(n15948) );
  NOR2_X1 U17814 ( .A1(n15948), .A2(n14533), .ZN(n15936) );
  NOR2_X1 U17815 ( .A1(n15936), .A2(n14534), .ZN(n14538) );
  INV_X1 U17816 ( .A(n15934), .ZN(n14535) );
  NOR2_X1 U17817 ( .A1(n14536), .A2(n14535), .ZN(n14537) );
  XNOR2_X1 U17818 ( .A(n14538), .B(n14537), .ZN(n16003) );
  NAND2_X1 U17819 ( .A1(n16003), .A2(n20064), .ZN(n14542) );
  INV_X1 U17820 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n14539) );
  OAI22_X1 U17821 ( .A1(n15984), .A2(n15870), .B1(n20066), .B2(n14539), .ZN(
        n14540) );
  AOI21_X1 U17822 ( .B1(n15979), .B2(n15868), .A(n14540), .ZN(n14541) );
  OAI211_X1 U17823 ( .C1(n20106), .C2(n15871), .A(n14542), .B(n14541), .ZN(
        P1_U2984) );
  NAND2_X1 U17824 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14543) );
  AND2_X1 U17825 ( .A1(n14160), .A2(n14543), .ZN(n15943) );
  OR2_X1 U17826 ( .A1(n14522), .A2(n15943), .ZN(n14547) );
  NAND2_X1 U17827 ( .A1(n14545), .A2(n14544), .ZN(n14546) );
  NAND2_X1 U17828 ( .A1(n14547), .A2(n14546), .ZN(n15957) );
  INV_X1 U17829 ( .A(n14550), .ZN(n14549) );
  NAND2_X1 U17830 ( .A1(n14545), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14548) );
  NAND2_X1 U17831 ( .A1(n14549), .A2(n14548), .ZN(n15956) );
  NOR2_X1 U17832 ( .A1(n15957), .A2(n15956), .ZN(n15955) );
  NOR2_X1 U17833 ( .A1(n15955), .A2(n14550), .ZN(n14551) );
  XOR2_X1 U17834 ( .A(n14552), .B(n14551), .Z(n14701) );
  NOR2_X1 U17835 ( .A1(n20066), .A2(n20819), .ZN(n14698) );
  AOI21_X1 U17836 ( .B1(n20060), .B2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n14698), .ZN(n14553) );
  OAI21_X1 U17837 ( .B1(n15978), .B2(n14554), .A(n14553), .ZN(n14555) );
  AOI21_X1 U17838 ( .B1(n14556), .B2(n15975), .A(n14555), .ZN(n14557) );
  OAI21_X1 U17839 ( .B1(n14701), .B2(n15962), .A(n14557), .ZN(P1_U2986) );
  MUX2_X1 U17840 ( .A(n14522), .B(n14558), .S(n14545), .Z(n14559) );
  XOR2_X1 U17841 ( .A(n16038), .B(n14559), .Z(n16034) );
  NAND2_X1 U17842 ( .A1(n16034), .A2(n20064), .ZN(n14562) );
  NOR2_X1 U17843 ( .A1(n20066), .A2(n20668), .ZN(n16028) );
  NOR2_X1 U17844 ( .A1(n15978), .A2(n15908), .ZN(n14560) );
  AOI211_X1 U17845 ( .C1(n20060), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16028), .B(n14560), .ZN(n14561) );
  OAI211_X1 U17846 ( .C1(n20106), .C2(n15907), .A(n14562), .B(n14561), .ZN(
        P1_U2989) );
  NOR3_X1 U17847 ( .A1(n16038), .A2(n14158), .A3(n16031), .ZN(n14710) );
  NAND2_X1 U17848 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14710), .ZN(
        n16019) );
  OR2_X1 U17849 ( .A1(n16022), .A2(n16019), .ZN(n14695) );
  NOR2_X1 U17850 ( .A1(n14563), .A2(n14695), .ZN(n16008) );
  NAND2_X1 U17851 ( .A1(n16008), .A2(n14706), .ZN(n14686) );
  INV_X1 U17852 ( .A(n14686), .ZN(n14564) );
  NAND2_X1 U17853 ( .A1(n13918), .A2(n14564), .ZN(n14641) );
  NAND2_X1 U17854 ( .A1(n14565), .A2(n16008), .ZN(n14573) );
  INV_X1 U17855 ( .A(n14573), .ZN(n14566) );
  NAND2_X1 U17856 ( .A1(n14709), .A2(n14566), .ZN(n14567) );
  NAND2_X1 U17857 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15993) );
  NOR3_X1 U17858 ( .A1(n16009), .A2(n14688), .A3(n15993), .ZN(n15987) );
  NAND2_X1 U17859 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15987), .ZN(
        n14575) );
  INV_X1 U17860 ( .A(n14575), .ZN(n14569) );
  AND2_X1 U17861 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14578) );
  INV_X1 U17862 ( .A(n14578), .ZN(n14666) );
  NOR2_X1 U17863 ( .A1(n14665), .A2(n14666), .ZN(n14568) );
  NAND2_X1 U17864 ( .A1(n14569), .A2(n14568), .ZN(n14570) );
  NOR3_X1 U17865 ( .A1(n14653), .A2(n14571), .A3(n14625), .ZN(n14607) );
  INV_X1 U17866 ( .A(n14581), .ZN(n14608) );
  NAND3_X1 U17867 ( .A1(n14607), .A2(n14608), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14592) );
  NAND2_X1 U17868 ( .A1(n14572), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14585) );
  INV_X1 U17869 ( .A(n14582), .ZN(n14579) );
  NOR2_X1 U17870 ( .A1(n14573), .A2(n14575), .ZN(n14664) );
  OAI21_X1 U17871 ( .B1(n14575), .B2(n14686), .A(n14574), .ZN(n14576) );
  OAI211_X1 U17872 ( .C1(n14664), .C2(n15755), .A(n14577), .B(n14576), .ZN(
        n15756) );
  OAI21_X1 U17873 ( .B1(n15756), .B2(n14665), .A(n14582), .ZN(n14672) );
  OAI21_X1 U17874 ( .B1(n14579), .B2(n14578), .A(n14672), .ZN(n14655) );
  AOI21_X1 U17875 ( .B1(n14625), .B2(n14580), .A(n14655), .ZN(n14636) );
  OAI21_X1 U17876 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n15995), .A(
        n14636), .ZN(n14617) );
  AOI21_X1 U17877 ( .B1(n14581), .B2(n14580), .A(n14617), .ZN(n14602) );
  OAI211_X1 U17878 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15995), .A(
        n14602), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14595) );
  NAND3_X1 U17879 ( .A1(n14595), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14582), .ZN(n14584) );
  OAI211_X1 U17880 ( .C1(n14592), .C2(n14585), .A(n14584), .B(n14583), .ZN(
        n14586) );
  INV_X1 U17881 ( .A(n14586), .ZN(n14587) );
  NAND2_X1 U17882 ( .A1(n14590), .A2(n20082), .ZN(n14597) );
  NAND2_X1 U17883 ( .A1(n14592), .A2(n14591), .ZN(n14594) );
  AOI21_X1 U17884 ( .B1(n14595), .B2(n14594), .A(n14593), .ZN(n14596) );
  OAI211_X1 U17885 ( .C1(n14598), .C2(n14712), .A(n14597), .B(n14596), .ZN(
        P1_U3001) );
  NAND3_X1 U17886 ( .A1(n14607), .A2(n14608), .A3(n14179), .ZN(n14600) );
  OAI211_X1 U17887 ( .C1(n14602), .C2(n14179), .A(n14601), .B(n14600), .ZN(
        n14603) );
  AOI21_X1 U17888 ( .B1(n11893), .B2(n20070), .A(n14603), .ZN(n14604) );
  OAI21_X1 U17889 ( .B1(n14605), .B2(n16025), .A(n14604), .ZN(P1_U3002) );
  INV_X1 U17890 ( .A(n14606), .ZN(n14611) );
  INV_X1 U17891 ( .A(n14607), .ZN(n14620) );
  NOR3_X1 U17892 ( .A1(n14620), .A2(n14609), .A3(n14608), .ZN(n14610) );
  AOI211_X1 U17893 ( .C1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .C2(n14617), .A(
        n14611), .B(n14610), .ZN(n14615) );
  INV_X1 U17894 ( .A(n14612), .ZN(n14613) );
  NAND2_X1 U17895 ( .A1(n14613), .A2(n20070), .ZN(n14614) );
  OAI211_X1 U17896 ( .C1(n14616), .C2(n16025), .A(n14615), .B(n14614), .ZN(
        P1_U3003) );
  NAND2_X1 U17897 ( .A1(n14617), .A2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14619) );
  OAI211_X1 U17898 ( .C1(n14620), .C2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14619), .B(n14618), .ZN(n14621) );
  AOI21_X1 U17899 ( .B1(n14622), .B2(n20070), .A(n14621), .ZN(n14623) );
  OAI21_X1 U17900 ( .B1(n14624), .B2(n16025), .A(n14623), .ZN(P1_U3004) );
  INV_X1 U17901 ( .A(n14636), .ZN(n14628) );
  NOR3_X1 U17902 ( .A1(n14653), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14625), .ZN(n14626) );
  AOI211_X1 U17903 ( .C1(n14628), .C2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n14627), .B(n14626), .ZN(n14631) );
  NAND2_X1 U17904 ( .A1(n14629), .A2(n20070), .ZN(n14630) );
  OAI211_X1 U17905 ( .C1(n14632), .C2(n16025), .A(n14631), .B(n14630), .ZN(
        P1_U3005) );
  INV_X1 U17906 ( .A(n14653), .ZN(n14644) );
  NAND4_X1 U17907 ( .A1(n14644), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A4(n14635), .ZN(n14633) );
  OAI211_X1 U17908 ( .C1(n14636), .C2(n14635), .A(n14634), .B(n14633), .ZN(
        n14637) );
  AOI21_X1 U17909 ( .B1(n14638), .B2(n20070), .A(n14637), .ZN(n14639) );
  OAI21_X1 U17910 ( .B1(n14640), .B2(n16025), .A(n14639), .ZN(P1_U3006) );
  AOI21_X1 U17911 ( .B1(n14641), .B2(n15755), .A(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n14642) );
  OAI21_X1 U17912 ( .B1(n14655), .B2(n14642), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14647) );
  NAND3_X1 U17913 ( .A1(n14644), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n14643), .ZN(n14646) );
  NAND3_X1 U17914 ( .A1(n14647), .A2(n14646), .A3(n14645), .ZN(n14648) );
  AOI21_X1 U17915 ( .B1(n15778), .B2(n20070), .A(n14648), .ZN(n14649) );
  OAI21_X1 U17916 ( .B1(n14650), .B2(n16025), .A(n14649), .ZN(P1_U3007) );
  NAND2_X1 U17917 ( .A1(n15788), .A2(n20070), .ZN(n14652) );
  OAI211_X1 U17918 ( .C1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n14653), .A(
        n14652), .B(n14651), .ZN(n14654) );
  AOI21_X1 U17919 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n14655), .A(
        n14654), .ZN(n14656) );
  OAI21_X1 U17920 ( .B1(n14657), .B2(n16025), .A(n14656), .ZN(P1_U3008) );
  NAND2_X1 U17921 ( .A1(n14658), .A2(n20082), .ZN(n14671) );
  OR2_X1 U17922 ( .A1(n14660), .A2(n14659), .ZN(n14661) );
  AND2_X1 U17923 ( .A1(n14661), .A2(n9772), .ZN(n15803) );
  AOI21_X1 U17924 ( .B1(n15803), .B2(n20070), .A(n14662), .ZN(n14670) );
  NAND2_X1 U17925 ( .A1(n14664), .A2(n14663), .ZN(n14679) );
  NOR2_X1 U17926 ( .A1(n14679), .A2(n14665), .ZN(n14676) );
  OAI211_X1 U17927 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n14676), .B(n14666), .ZN(
        n14669) );
  OR2_X1 U17928 ( .A1(n14672), .A2(n14667), .ZN(n14668) );
  NAND4_X1 U17929 ( .A1(n14671), .A2(n14670), .A3(n14669), .A4(n14668), .ZN(
        P1_U3009) );
  NOR2_X1 U17930 ( .A1(n14672), .A2(n14675), .ZN(n14674) );
  INV_X1 U17931 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20683) );
  OAI22_X1 U17932 ( .A1(n15817), .A2(n14712), .B1(n20683), .B2(n20066), .ZN(
        n14673) );
  AOI211_X1 U17933 ( .C1(n14676), .C2(n14675), .A(n14674), .B(n14673), .ZN(
        n14677) );
  OAI21_X1 U17934 ( .B1(n14678), .B2(n16025), .A(n14677), .ZN(P1_U3010) );
  INV_X1 U17935 ( .A(n14679), .ZN(n15754) );
  NAND2_X1 U17936 ( .A1(n15749), .A2(n15754), .ZN(n14680) );
  OAI211_X1 U17937 ( .C1(n15839), .C2(n14712), .A(n14681), .B(n14680), .ZN(
        n14682) );
  AOI21_X1 U17938 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15756), .A(
        n14682), .ZN(n14683) );
  OAI21_X1 U17939 ( .B1(n14684), .B2(n16025), .A(n14683), .ZN(P1_U3012) );
  INV_X1 U17940 ( .A(n15857), .ZN(n14691) );
  NOR2_X1 U17941 ( .A1(n20066), .A2(n20676), .ZN(n14690) );
  OAI21_X1 U17942 ( .B1(n15755), .B2(n16008), .A(n14705), .ZN(n14685) );
  AOI21_X1 U17943 ( .B1(n14686), .B2(n14685), .A(n14707), .ZN(n15994) );
  OAI21_X1 U17944 ( .B1(n15995), .B2(n15987), .A(n15994), .ZN(n14687) );
  INV_X1 U17945 ( .A(n14687), .ZN(n15992) );
  AOI221_X1 U17946 ( .B1(n15993), .B2(n14688), .C1(n16006), .C2(n14688), .A(
        n15992), .ZN(n14689) );
  AOI211_X1 U17947 ( .C1(n20085), .C2(n14691), .A(n14690), .B(n14689), .ZN(
        n14692) );
  OAI21_X1 U17948 ( .B1(n14693), .B2(n16025), .A(n14692), .ZN(P1_U3014) );
  INV_X1 U17949 ( .A(n14694), .ZN(n14699) );
  NOR2_X1 U17950 ( .A1(n14695), .A2(n16030), .ZN(n14696) );
  INV_X1 U17951 ( .A(n15994), .ZN(n16007) );
  MUX2_X1 U17952 ( .A(n14696), .B(n16007), .S(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(n14697) );
  AOI211_X1 U17953 ( .C1(n20085), .C2(n14699), .A(n14698), .B(n14697), .ZN(
        n14700) );
  OAI21_X1 U17954 ( .B1(n14701), .B2(n16025), .A(n14700), .ZN(P1_U3018) );
  NOR2_X1 U17955 ( .A1(n14558), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14703) );
  NOR2_X1 U17956 ( .A1(n14522), .A2(n16038), .ZN(n14702) );
  MUX2_X1 U17957 ( .A(n14703), .B(n14702), .S(n14160), .Z(n14704) );
  XNOR2_X1 U17958 ( .A(n14704), .B(n14711), .ZN(n15964) );
  AOI21_X1 U17959 ( .B1(n14710), .B2(n14706), .A(n14705), .ZN(n14708) );
  AOI211_X1 U17960 ( .C1(n14709), .C2(n16019), .A(n14708), .B(n14707), .ZN(
        n16016) );
  INV_X1 U17961 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14711) );
  NAND2_X1 U17962 ( .A1(n14710), .A2(n14711), .ZN(n16017) );
  OAI22_X1 U17963 ( .A1(n16016), .A2(n14711), .B1(n16030), .B2(n16017), .ZN(
        n14714) );
  OAI22_X1 U17964 ( .A1(n14712), .A2(n15896), .B1(n20066), .B2(n20840), .ZN(
        n14713) );
  AOI211_X1 U17965 ( .C1(n15964), .C2(n20082), .A(n14714), .B(n14713), .ZN(
        n14715) );
  INV_X1 U17966 ( .A(n14715), .ZN(P1_U3020) );
  INV_X1 U17967 ( .A(n15731), .ZN(n14725) );
  NOR2_X1 U17968 ( .A1(n10928), .A2(n10930), .ZN(n14717) );
  INV_X1 U17969 ( .A(n14717), .ZN(n14724) );
  AOI22_X1 U17970 ( .A1(n15704), .A2(n14718), .B1(n14717), .B2(n14716), .ZN(
        n14719) );
  OAI21_X1 U17971 ( .B1(n13669), .B2(n14720), .A(n14719), .ZN(n15700) );
  AOI22_X1 U17972 ( .A1(n15700), .A2(n19883), .B1(n14722), .B2(n14721), .ZN(
        n14723) );
  OAI21_X1 U17973 ( .B1(n14725), .B2(n14724), .A(n14723), .ZN(n14727) );
  MUX2_X1 U17974 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14727), .S(
        n14726), .Z(P1_U3473) );
  NAND2_X1 U17975 ( .A1(n14728), .A2(n14729), .ZN(n14730) );
  NAND2_X1 U17976 ( .A1(n14923), .A2(n14730), .ZN(n15344) );
  OAI211_X1 U17977 ( .C1(n14732), .C2(n15103), .A(n18915), .B(n14731), .ZN(
        n14743) );
  OAI22_X1 U17978 ( .A1(n10713), .A2(n19031), .B1(n15102), .B2(n18999), .ZN(
        n14740) );
  OR2_X1 U17979 ( .A1(n14734), .A2(n14733), .ZN(n14736) );
  AND2_X1 U17980 ( .A1(n14736), .A2(n14735), .ZN(n15341) );
  INV_X1 U17981 ( .A(n15341), .ZN(n14738) );
  OAI22_X1 U17982 ( .A1(n19026), .A2(n14738), .B1(n19041), .B2(n14737), .ZN(
        n14739) );
  AOI211_X1 U17983 ( .C1(n14741), .C2(n19035), .A(n14740), .B(n14739), .ZN(
        n14742) );
  OAI211_X1 U17984 ( .C1(n19037), .C2(n15344), .A(n14743), .B(n14742), .ZN(
        P2_U2832) );
  OR2_X1 U17985 ( .A1(n14760), .A2(n14744), .ZN(n14745) );
  NAND2_X1 U17986 ( .A1(n14728), .A2(n14745), .ZN(n15356) );
  INV_X1 U17987 ( .A(n15356), .ZN(n14757) );
  INV_X1 U17988 ( .A(n14746), .ZN(n14747) );
  XNOR2_X1 U17989 ( .A(n14748), .B(n14747), .ZN(n15352) );
  AOI22_X1 U17990 ( .A1(n18957), .A2(P2_EBX_REG_22__SCAN_IN), .B1(n19029), 
        .B2(n15352), .ZN(n14749) );
  OAI21_X1 U17991 ( .B1(n14750), .B2(n19014), .A(n14749), .ZN(n14756) );
  OAI211_X1 U17992 ( .C1(n15113), .C2(n14752), .A(n18915), .B(n14751), .ZN(
        n14754) );
  AOI22_X1 U17993 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n19003), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19028), .ZN(n14753) );
  NAND2_X1 U17994 ( .A1(n14754), .A2(n14753), .ZN(n14755) );
  AOI211_X1 U17995 ( .C1(n10916), .C2(n14757), .A(n14756), .B(n14755), .ZN(
        n14758) );
  INV_X1 U17996 ( .A(n14758), .ZN(P2_U2833) );
  NOR2_X1 U17997 ( .A1(n14760), .A2(n10150), .ZN(n15361) );
  INV_X1 U17998 ( .A(n15361), .ZN(n14773) );
  NOR2_X1 U17999 ( .A1(n19005), .A2(n14774), .ZN(n14763) );
  NAND2_X1 U18000 ( .A1(n14762), .A2(n14763), .ZN(n14761) );
  OAI211_X1 U18001 ( .C1(n14763), .C2(n14762), .A(n18915), .B(n14761), .ZN(
        n14772) );
  XNOR2_X1 U18002 ( .A(n14782), .B(n14765), .ZN(n16149) );
  NAND2_X1 U18003 ( .A1(n19029), .A2(n16149), .ZN(n14767) );
  AOI22_X1 U18004 ( .A1(P2_EBX_REG_21__SCAN_IN), .A2(n18957), .B1(
        P2_REIP_REG_21__SCAN_IN), .B2(n19028), .ZN(n14766) );
  OAI211_X1 U18005 ( .C1(n19041), .C2(n14768), .A(n14767), .B(n14766), .ZN(
        n14769) );
  AOI21_X1 U18006 ( .B1(n14770), .B2(n19035), .A(n14769), .ZN(n14771) );
  OAI211_X1 U18007 ( .C1(n19037), .C2(n14773), .A(n14772), .B(n14771), .ZN(
        P2_U2834) );
  AOI211_X1 U18008 ( .C1(n15144), .C2(n14775), .A(n14774), .B(n16073), .ZN(
        n14789) );
  OAI22_X1 U18009 ( .A1(n9999), .A2(n19041), .B1(n14776), .B2(n19040), .ZN(
        n14788) );
  INV_X1 U18010 ( .A(n14955), .ZN(n14779) );
  OAI21_X1 U18011 ( .B1(n14779), .B2(n10012), .A(n14778), .ZN(n15380) );
  NAND2_X1 U18012 ( .A1(n15016), .A2(n14780), .ZN(n14781) );
  AND2_X1 U18013 ( .A1(n14782), .A2(n14781), .ZN(n15376) );
  INV_X1 U18014 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n14950) );
  OAI22_X1 U18015 ( .A1(n14950), .A2(n19031), .B1(n10882), .B2(n18999), .ZN(
        n14783) );
  AOI21_X1 U18016 ( .B1(n19029), .B2(n15376), .A(n14783), .ZN(n14786) );
  NAND2_X1 U18017 ( .A1(n14784), .A2(n19035), .ZN(n14785) );
  OAI211_X1 U18018 ( .C1(n15380), .C2(n19037), .A(n14786), .B(n14785), .ZN(
        n14787) );
  OR3_X1 U18019 ( .A1(n14789), .A2(n14788), .A3(n14787), .ZN(P2_U2835) );
  INV_X1 U18020 ( .A(n14790), .ZN(n14806) );
  NOR2_X1 U18021 ( .A1(n19005), .A2(n14791), .ZN(n14792) );
  XNOR2_X1 U18022 ( .A(n14792), .B(n16165), .ZN(n14793) );
  NAND2_X1 U18023 ( .A1(n14793), .A2(n18915), .ZN(n14805) );
  INV_X1 U18024 ( .A(n14795), .ZN(n14796) );
  AOI21_X1 U18025 ( .B1(n10014), .B2(n14796), .A(n9819), .ZN(n16162) );
  NAND2_X1 U18026 ( .A1(n9827), .A2(n14797), .ZN(n14799) );
  INV_X1 U18027 ( .A(n15014), .ZN(n14798) );
  NAND2_X1 U18028 ( .A1(n14799), .A2(n14798), .ZN(n15412) );
  NOR2_X1 U18029 ( .A1(n15412), .A2(n19026), .ZN(n14803) );
  INV_X1 U18030 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n14801) );
  AOI22_X1 U18031 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19003), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n19028), .ZN(n14800) );
  OAI211_X1 U18032 ( .C1(n19031), .C2(n14801), .A(n14800), .B(n19012), .ZN(
        n14802) );
  AOI211_X1 U18033 ( .C1(n16162), .C2(n10916), .A(n14803), .B(n14802), .ZN(
        n14804) );
  OAI211_X1 U18034 ( .C1(n19014), .C2(n14806), .A(n14805), .B(n14804), .ZN(
        P2_U2837) );
  NOR2_X1 U18035 ( .A1(n19005), .A2(n14807), .ZN(n14808) );
  XNOR2_X1 U18036 ( .A(n14808), .B(n15224), .ZN(n14809) );
  NAND2_X1 U18037 ( .A1(n14809), .A2(n18915), .ZN(n14817) );
  AOI22_X1 U18038 ( .A1(n14810), .A2(n19035), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n19003), .ZN(n14811) );
  OAI211_X1 U18039 ( .C1(n14812), .C2(n19031), .A(n14811), .B(n19012), .ZN(
        n14813) );
  AOI21_X1 U18040 ( .B1(P2_REIP_REG_10__SCAN_IN), .B2(n19028), .A(n14813), 
        .ZN(n14816) );
  AOI21_X1 U18041 ( .B1(n14814), .B2(n15514), .A(n9841), .ZN(n19062) );
  AOI22_X1 U18042 ( .A1(n16210), .A2(n10916), .B1(n19029), .B2(n19062), .ZN(
        n14815) );
  NAND3_X1 U18043 ( .A1(n14817), .A2(n14816), .A3(n14815), .ZN(P2_U2845) );
  NOR2_X1 U18044 ( .A1(n19005), .A2(n14818), .ZN(n14819) );
  XNOR2_X1 U18045 ( .A(n14819), .B(n15245), .ZN(n14820) );
  NAND2_X1 U18046 ( .A1(n14820), .A2(n18915), .ZN(n14829) );
  AOI22_X1 U18047 ( .A1(n14821), .A2(n19035), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19003), .ZN(n14822) );
  OAI211_X1 U18048 ( .C1(n10707), .C2(n19031), .A(n14822), .B(n19012), .ZN(
        n14823) );
  AOI21_X1 U18049 ( .B1(P2_REIP_REG_8__SCAN_IN), .B2(n19028), .A(n14823), .ZN(
        n14828) );
  AOI21_X1 U18050 ( .B1(n14826), .B2(n14824), .A(n14825), .ZN(n19067) );
  AOI22_X1 U18051 ( .A1(n16222), .A2(n10916), .B1(n19029), .B2(n19067), .ZN(
        n14827) );
  NAND3_X1 U18052 ( .A1(n14829), .A2(n14828), .A3(n14827), .ZN(P2_U2847) );
  NOR2_X1 U18053 ( .A1(n19005), .A2(n14830), .ZN(n14831) );
  XNOR2_X1 U18054 ( .A(n14831), .B(n19204), .ZN(n14841) );
  AOI22_X1 U18055 ( .A1(P2_EBX_REG_4__SCAN_IN), .A2(n18957), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19028), .ZN(n14835) );
  AOI21_X1 U18056 ( .B1(n14832), .B2(n13775), .A(n9775), .ZN(n19207) );
  AOI22_X1 U18057 ( .A1(n19035), .A2(n14833), .B1(n19029), .B2(n19207), .ZN(
        n14834) );
  NAND3_X1 U18058 ( .A1(n14835), .A2(n14834), .A3(n19012), .ZN(n14836) );
  AOI21_X1 U18059 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n19003), .A(
        n14836), .ZN(n14839) );
  INV_X1 U18060 ( .A(n14837), .ZN(n19213) );
  NAND2_X1 U18061 ( .A1(n19213), .A2(n10916), .ZN(n14838) );
  OAI211_X1 U18062 ( .C1(n19088), .C2(n14877), .A(n14839), .B(n14838), .ZN(
        n14840) );
  AOI21_X1 U18063 ( .B1(n14841), .B2(n18915), .A(n14840), .ZN(n14842) );
  INV_X1 U18064 ( .A(n14842), .ZN(P2_U2851) );
  NAND2_X1 U18065 ( .A1(n19019), .A2(n14843), .ZN(n14844) );
  XNOR2_X1 U18066 ( .A(n14845), .B(n14844), .ZN(n14846) );
  NAND2_X1 U18067 ( .A1(n14846), .A2(n18915), .ZN(n14853) );
  OAI22_X1 U18068 ( .A1(n10704), .A2(n19031), .B1(n10803), .B2(n18999), .ZN(
        n14847) );
  AOI21_X1 U18069 ( .B1(n19003), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n14847), .ZN(n14848) );
  OAI21_X1 U18070 ( .B1(n19014), .B2(n14849), .A(n14848), .ZN(n14851) );
  NOR2_X1 U18071 ( .A1(n19096), .A2(n19026), .ZN(n14850) );
  AOI211_X1 U18072 ( .C1(n10916), .C2(n13777), .A(n14851), .B(n14850), .ZN(
        n14852) );
  OAI211_X1 U18073 ( .C1(n19818), .C2(n14877), .A(n14853), .B(n14852), .ZN(
        P2_U2852) );
  NOR2_X1 U18074 ( .A1(n19005), .A2(n14865), .ZN(n14855) );
  XNOR2_X1 U18075 ( .A(n14855), .B(n14854), .ZN(n14856) );
  NAND2_X1 U18076 ( .A1(n14856), .A2(n18915), .ZN(n14864) );
  OAI22_X1 U18077 ( .A1(n14857), .A2(n19031), .B1(n10790), .B2(n18999), .ZN(
        n14860) );
  NOR2_X1 U18078 ( .A1(n19014), .A2(n14858), .ZN(n14859) );
  AOI211_X1 U18079 ( .C1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .C2(n19003), .A(
        n14860), .B(n14859), .ZN(n14861) );
  OAI21_X1 U18080 ( .B1(n11907), .B2(n19037), .A(n14861), .ZN(n14862) );
  AOI21_X1 U18081 ( .B1(n19829), .B2(n19029), .A(n14862), .ZN(n14863) );
  OAI211_X1 U18082 ( .C1(n19825), .C2(n14877), .A(n14864), .B(n14863), .ZN(
        P2_U2853) );
  AOI211_X1 U18083 ( .C1(n14867), .C2(n14866), .A(n19005), .B(n14865), .ZN(
        n15576) );
  NAND2_X1 U18084 ( .A1(n15576), .A2(n18915), .ZN(n14876) );
  OAI22_X1 U18085 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19040), .B1(
        n19041), .B2(n13219), .ZN(n14870) );
  NOR2_X1 U18086 ( .A1(n18999), .A2(n14868), .ZN(n14869) );
  AOI211_X1 U18087 ( .C1(n18957), .C2(P2_EBX_REG_1__SCAN_IN), .A(n14870), .B(
        n14869), .ZN(n14872) );
  NAND2_X1 U18088 ( .A1(n19833), .A2(n19029), .ZN(n14871) );
  OAI211_X1 U18089 ( .C1(n19014), .C2(n14873), .A(n14872), .B(n14871), .ZN(
        n14874) );
  AOI21_X1 U18090 ( .B1(n15568), .B2(n10916), .A(n14874), .ZN(n14875) );
  OAI211_X1 U18091 ( .C1(n19838), .C2(n14877), .A(n14876), .B(n14875), .ZN(
        P2_U2854) );
  MUX2_X1 U18092 ( .A(n12774), .B(P2_EBX_REG_31__SCAN_IN), .S(n13257), .Z(
        P2_U2856) );
  NOR2_X1 U18093 ( .A1(n15275), .A2(n13257), .ZN(n14883) );
  AOI21_X1 U18094 ( .B1(P2_EBX_REG_29__SCAN_IN), .B2(n13257), .A(n14883), .ZN(
        n14884) );
  OAI21_X1 U18095 ( .B1(n14973), .B2(n14966), .A(n14884), .ZN(P2_U2858) );
  INV_X1 U18096 ( .A(n14885), .ZN(n14886) );
  NOR2_X1 U18097 ( .A1(n14887), .A2(n14886), .ZN(n14889) );
  XNOR2_X1 U18098 ( .A(n14889), .B(n14888), .ZN(n14977) );
  NOR2_X1 U18099 ( .A1(n14890), .A2(n13257), .ZN(n14891) );
  AOI21_X1 U18100 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n13257), .A(n14891), .ZN(
        n14892) );
  OAI21_X1 U18101 ( .B1(n14977), .B2(n14966), .A(n14892), .ZN(P2_U2859) );
  AOI21_X1 U18102 ( .B1(n14893), .B2(n14895), .A(n14894), .ZN(n14896) );
  INV_X1 U18103 ( .A(n14896), .ZN(n14984) );
  NAND2_X1 U18104 ( .A1(n14897), .A2(n14898), .ZN(n14899) );
  NAND2_X1 U18105 ( .A1(n14900), .A2(n14899), .ZN(n16096) );
  NOR2_X1 U18106 ( .A1(n16096), .A2(n13257), .ZN(n14901) );
  AOI21_X1 U18107 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n13257), .A(n14901), .ZN(
        n14902) );
  OAI21_X1 U18108 ( .B1(n14984), .B2(n14966), .A(n14902), .ZN(P2_U2860) );
  AOI21_X1 U18109 ( .B1(n14905), .B2(n14904), .A(n14903), .ZN(n14906) );
  INV_X1 U18110 ( .A(n14906), .ZN(n14990) );
  OAI21_X1 U18111 ( .B1(n14907), .B2(n14908), .A(n14897), .ZN(n16108) );
  NOR2_X1 U18112 ( .A1(n16108), .A2(n13257), .ZN(n14909) );
  AOI21_X1 U18113 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n13257), .A(n14909), .ZN(
        n14910) );
  OAI21_X1 U18114 ( .B1(n14990), .B2(n14966), .A(n14910), .ZN(P2_U2861) );
  XNOR2_X1 U18115 ( .A(n14911), .B(n14912), .ZN(n14996) );
  NOR2_X1 U18116 ( .A1(n9818), .A2(n14913), .ZN(n14914) );
  OR2_X1 U18117 ( .A1(n14907), .A2(n14914), .ZN(n16123) );
  MUX2_X1 U18118 ( .A(n16123), .B(n14915), .S(n13257), .Z(n14916) );
  OAI21_X1 U18119 ( .B1(n14996), .B2(n14966), .A(n14916), .ZN(P2_U2862) );
  NOR2_X1 U18120 ( .A1(n14918), .A2(n9743), .ZN(n14919) );
  XNOR2_X1 U18121 ( .A(n14920), .B(n14919), .ZN(n14921) );
  XNOR2_X1 U18122 ( .A(n14917), .B(n14921), .ZN(n16144) );
  NAND2_X1 U18123 ( .A1(n16144), .A2(n14941), .ZN(n14926) );
  AND2_X1 U18124 ( .A1(n14923), .A2(n14922), .ZN(n14924) );
  NOR2_X1 U18125 ( .A1(n9818), .A2(n14924), .ZN(n16133) );
  NAND2_X1 U18126 ( .A1(n16133), .A2(n13251), .ZN(n14925) );
  OAI211_X1 U18127 ( .C1(n13251), .C2(n14927), .A(n14926), .B(n14925), .ZN(
        P2_U2863) );
  OAI21_X1 U18128 ( .B1(n14928), .B2(n14930), .A(n14929), .ZN(n15000) );
  NOR2_X1 U18129 ( .A1(n15344), .A2(n13257), .ZN(n14931) );
  AOI21_X1 U18130 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n13257), .A(n14931), .ZN(
        n14932) );
  OAI21_X1 U18131 ( .B1(n15000), .B2(n14966), .A(n14932), .ZN(P2_U2864) );
  NAND2_X1 U18132 ( .A1(n14933), .A2(n14938), .ZN(n14940) );
  AOI21_X1 U18133 ( .B1(n14935), .B2(n14940), .A(n14934), .ZN(n15001) );
  NAND2_X1 U18134 ( .A1(n15001), .A2(n14941), .ZN(n14937) );
  NAND2_X1 U18135 ( .A1(n13257), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n14936) );
  OAI211_X1 U18136 ( .C1(n15356), .C2(n13257), .A(n14937), .B(n14936), .ZN(
        P2_U2865) );
  OR2_X1 U18137 ( .A1(n14933), .A2(n14938), .ZN(n14939) );
  NAND2_X1 U18138 ( .A1(n16150), .A2(n14941), .ZN(n14943) );
  NAND2_X1 U18139 ( .A1(n15361), .A2(n13251), .ZN(n14942) );
  OAI211_X1 U18140 ( .C1(n13251), .C2(n14944), .A(n14943), .B(n14942), .ZN(
        P2_U2866) );
  INV_X1 U18141 ( .A(n14946), .ZN(n14949) );
  INV_X1 U18142 ( .A(n14933), .ZN(n14947) );
  OAI21_X1 U18143 ( .B1(n14949), .B2(n14948), .A(n14947), .ZN(n15013) );
  MUX2_X1 U18144 ( .A(n15380), .B(n14950), .S(n13257), .Z(n14951) );
  OAI21_X1 U18145 ( .B1(n15013), .B2(n14966), .A(n14951), .ZN(P2_U2867) );
  OAI21_X1 U18146 ( .B1(n12464), .B2(n14953), .A(n14946), .ZN(n15023) );
  OAI21_X1 U18147 ( .B1(n9819), .B2(n10879), .A(n14955), .ZN(n18912) );
  NOR2_X1 U18148 ( .A1(n18912), .A2(n13257), .ZN(n14956) );
  AOI21_X1 U18149 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n13257), .A(n14956), .ZN(
        n14957) );
  OAI21_X1 U18150 ( .B1(n15023), .B2(n14966), .A(n14957), .ZN(P2_U2868) );
  OAI21_X1 U18151 ( .B1(n14959), .B2(n14958), .A(n14952), .ZN(n15031) );
  INV_X1 U18152 ( .A(n16162), .ZN(n15413) );
  NOR2_X1 U18153 ( .A1(n15413), .A2(n13257), .ZN(n14960) );
  AOI21_X1 U18154 ( .B1(P2_EBX_REG_18__SCAN_IN), .B2(n13257), .A(n14960), .ZN(
        n14961) );
  OAI21_X1 U18155 ( .B1(n15031), .B2(n14966), .A(n14961), .ZN(P2_U2869) );
  NOR2_X1 U18156 ( .A1(n13941), .A2(n14962), .ZN(n14963) );
  OR2_X1 U18157 ( .A1(n14795), .A2(n14963), .ZN(n18925) );
  NOR2_X1 U18158 ( .A1(n18925), .A2(n13257), .ZN(n14964) );
  AOI21_X1 U18159 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n13257), .A(n14964), .ZN(
        n14965) );
  OAI21_X1 U18160 ( .B1(n14967), .B2(n14966), .A(n14965), .ZN(P2_U2870) );
  XOR2_X1 U18161 ( .A(n14968), .B(n9769), .Z(n16075) );
  INV_X1 U18162 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14969) );
  OAI22_X1 U18163 ( .A1(n16141), .A2(n19056), .B1(n19072), .B2(n14969), .ZN(
        n14970) );
  AOI21_X1 U18164 ( .B1(n19106), .B2(n16075), .A(n14970), .ZN(n14972) );
  AOI22_X1 U18165 ( .A1(n19047), .A2(BUF2_REG_29__SCAN_IN), .B1(n19049), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n14971) );
  OAI211_X1 U18166 ( .C1(n14973), .C2(n19082), .A(n14972), .B(n14971), .ZN(
        P2_U2890) );
  INV_X1 U18167 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n19127) );
  OAI22_X1 U18168 ( .A1(n16141), .A2(n19058), .B1(n19072), .B2(n19127), .ZN(
        n14974) );
  AOI21_X1 U18169 ( .B1(n19106), .B2(n16085), .A(n14974), .ZN(n14976) );
  AOI22_X1 U18170 ( .A1(n19047), .A2(BUF2_REG_28__SCAN_IN), .B1(n19049), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n14975) );
  OAI211_X1 U18171 ( .C1(n14977), .C2(n19082), .A(n14976), .B(n14975), .ZN(
        P2_U2891) );
  NAND2_X1 U18172 ( .A1(n14978), .A2(n14979), .ZN(n14980) );
  INV_X1 U18173 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n19129) );
  OAI22_X1 U18174 ( .A1(n16141), .A2(n19060), .B1(n19072), .B2(n19129), .ZN(
        n14981) );
  AOI21_X1 U18175 ( .B1(n19106), .B2(n16097), .A(n14981), .ZN(n14983) );
  AOI22_X1 U18176 ( .A1(n19047), .A2(BUF2_REG_27__SCAN_IN), .B1(n19049), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n14982) );
  OAI211_X1 U18177 ( .C1(n14984), .C2(n19082), .A(n14983), .B(n14982), .ZN(
        P2_U2892) );
  OAI21_X1 U18178 ( .B1(n14985), .B2(n14986), .A(n14978), .ZN(n15302) );
  INV_X1 U18179 ( .A(n15302), .ZN(n16109) );
  INV_X1 U18180 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n19131) );
  OAI22_X1 U18181 ( .A1(n16141), .A2(n19063), .B1(n19072), .B2(n19131), .ZN(
        n14987) );
  AOI21_X1 U18182 ( .B1(n19106), .B2(n16109), .A(n14987), .ZN(n14989) );
  AOI22_X1 U18183 ( .A1(n19047), .A2(BUF2_REG_26__SCAN_IN), .B1(n19049), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n14988) );
  OAI211_X1 U18184 ( .C1(n14990), .C2(n19082), .A(n14989), .B(n14988), .ZN(
        P2_U2893) );
  AND2_X1 U18185 ( .A1(n9792), .A2(n14991), .ZN(n14992) );
  NOR2_X1 U18186 ( .A1(n14985), .A2(n14992), .ZN(n16121) );
  INV_X1 U18187 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n20748) );
  OAI22_X1 U18188 ( .A1(n16141), .A2(n19065), .B1(n19072), .B2(n20748), .ZN(
        n14993) );
  AOI21_X1 U18189 ( .B1(n19106), .B2(n16121), .A(n14993), .ZN(n14995) );
  AOI22_X1 U18190 ( .A1(n19047), .A2(BUF2_REG_25__SCAN_IN), .B1(n19049), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n14994) );
  OAI211_X1 U18191 ( .C1(n14996), .C2(n19082), .A(n14995), .B(n14994), .ZN(
        P2_U2894) );
  INV_X1 U18192 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n19135) );
  OAI22_X1 U18193 ( .A1(n16141), .A2(n19256), .B1(n19072), .B2(n19135), .ZN(
        n14997) );
  AOI21_X1 U18194 ( .B1(n19106), .B2(n15341), .A(n14997), .ZN(n14999) );
  AOI22_X1 U18195 ( .A1(n19047), .A2(BUF2_REG_23__SCAN_IN), .B1(n19049), .B2(
        BUF1_REG_23__SCAN_IN), .ZN(n14998) );
  OAI211_X1 U18196 ( .C1(n15000), .C2(n19082), .A(n14999), .B(n14998), .ZN(
        P2_U2896) );
  INV_X1 U18197 ( .A(n15001), .ZN(n15007) );
  INV_X1 U18198 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n19137) );
  OAI22_X1 U18199 ( .A1(n16141), .A2(n19246), .B1(n19072), .B2(n19137), .ZN(
        n15005) );
  INV_X1 U18200 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n15003) );
  INV_X1 U18201 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n15002) );
  OAI22_X1 U18202 ( .A1(n15026), .A2(n15003), .B1(n15024), .B2(n15002), .ZN(
        n15004) );
  AOI211_X1 U18203 ( .C1(n19106), .C2(n15352), .A(n15005), .B(n15004), .ZN(
        n15006) );
  OAI21_X1 U18204 ( .B1(n15007), .B2(n19082), .A(n15006), .ZN(P2_U2897) );
  INV_X1 U18205 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n19141) );
  OAI22_X1 U18206 ( .A1(n16141), .A2(n19234), .B1(n19072), .B2(n19141), .ZN(
        n15011) );
  INV_X1 U18207 ( .A(BUF2_REG_20__SCAN_IN), .ZN(n15009) );
  INV_X1 U18208 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n15008) );
  OAI22_X1 U18209 ( .A1(n15026), .A2(n15009), .B1(n15024), .B2(n15008), .ZN(
        n15010) );
  AOI211_X1 U18210 ( .C1(n19106), .C2(n15376), .A(n15011), .B(n15010), .ZN(
        n15012) );
  OAI21_X1 U18211 ( .B1(n15013), .B2(n19082), .A(n15012), .ZN(P2_U2899) );
  OR2_X1 U18212 ( .A1(n15015), .A2(n15014), .ZN(n15017) );
  AND2_X1 U18213 ( .A1(n15017), .A2(n15016), .ZN(n18910) );
  INV_X1 U18214 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n19143) );
  OAI22_X1 U18215 ( .A1(n16141), .A2(n19229), .B1(n19072), .B2(n19143), .ZN(
        n15021) );
  INV_X1 U18216 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n15019) );
  INV_X1 U18217 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n15018) );
  OAI22_X1 U18218 ( .A1(n15026), .A2(n15019), .B1(n15024), .B2(n15018), .ZN(
        n15020) );
  AOI211_X1 U18219 ( .C1(n19106), .C2(n18910), .A(n15021), .B(n15020), .ZN(
        n15022) );
  OAI21_X1 U18220 ( .B1(n15023), .B2(n19082), .A(n15022), .ZN(P2_U2900) );
  INV_X1 U18221 ( .A(n15412), .ZN(n15029) );
  INV_X1 U18222 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n19145) );
  OAI22_X1 U18223 ( .A1(n16141), .A2(n19224), .B1(n19072), .B2(n19145), .ZN(
        n15028) );
  INV_X1 U18224 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n15025) );
  OAI22_X1 U18225 ( .A1(n15026), .A2(n15025), .B1(n15024), .B2(n16371), .ZN(
        n15027) );
  AOI211_X1 U18226 ( .C1(n19106), .C2(n15029), .A(n15028), .B(n15027), .ZN(
        n15030) );
  OAI21_X1 U18227 ( .B1(n15031), .B2(n19082), .A(n15030), .ZN(P2_U2901) );
  XNOR2_X1 U18228 ( .A(n15053), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n15274) );
  NAND2_X1 U18229 ( .A1(n15033), .A2(n15046), .ZN(n15038) );
  INV_X1 U18230 ( .A(n15034), .ZN(n15036) );
  NAND2_X1 U18231 ( .A1(n15036), .A2(n15035), .ZN(n15037) );
  XNOR2_X1 U18232 ( .A(n15038), .B(n15037), .ZN(n15272) );
  INV_X1 U18233 ( .A(n15039), .ZN(n15041) );
  NAND2_X1 U18234 ( .A1(n19206), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n15264) );
  OAI21_X1 U18235 ( .B1(n16194), .B2(n10699), .A(n15264), .ZN(n15040) );
  AOI21_X1 U18236 ( .B1(n15041), .B2(n16187), .A(n15040), .ZN(n15042) );
  OAI21_X1 U18237 ( .B1(n15270), .B2(n16186), .A(n15042), .ZN(n15043) );
  AOI21_X1 U18238 ( .B1(n15272), .B2(n16190), .A(n15043), .ZN(n15044) );
  OAI21_X1 U18239 ( .B1(n19197), .B2(n15274), .A(n15044), .ZN(P2_U2984) );
  NAND2_X1 U18240 ( .A1(n15046), .A2(n15045), .ZN(n15048) );
  XOR2_X1 U18241 ( .A(n15048), .B(n15047), .Z(n15288) );
  NAND2_X1 U18242 ( .A1(n19206), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n15280) );
  OAI21_X1 U18243 ( .B1(n16194), .B2(n15049), .A(n15280), .ZN(n15051) );
  NOR2_X1 U18244 ( .A1(n15275), .A2(n16186), .ZN(n15050) );
  AOI211_X1 U18245 ( .C1(n16187), .C2(n15052), .A(n15051), .B(n15050), .ZN(
        n15055) );
  NAND2_X1 U18246 ( .A1(n15285), .A2(n16188), .ZN(n15054) );
  OAI211_X1 U18247 ( .C1(n15288), .C2(n19198), .A(n15055), .B(n15054), .ZN(
        P2_U2985) );
  NAND2_X1 U18248 ( .A1(n15068), .A2(n15056), .ZN(n15289) );
  NAND2_X1 U18249 ( .A1(n15289), .A2(n16188), .ZN(n15065) );
  OR2_X1 U18250 ( .A1(n15057), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15290) );
  NAND3_X1 U18251 ( .A1(n15290), .A2(n16190), .A3(n15058), .ZN(n15064) );
  NAND2_X1 U18252 ( .A1(n19206), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15291) );
  OAI21_X1 U18253 ( .B1(n16194), .B2(n15059), .A(n15291), .ZN(n15061) );
  NOR2_X1 U18254 ( .A1(n16096), .A2(n16186), .ZN(n15060) );
  AOI211_X1 U18255 ( .C1(n16187), .C2(n15062), .A(n15061), .B(n15060), .ZN(
        n15063) );
  OAI211_X1 U18256 ( .C1(n15301), .C2(n15065), .A(n15064), .B(n15063), .ZN(
        P2_U2987) );
  BUF_X1 U18257 ( .A(n15066), .Z(n15067) );
  OAI21_X1 U18258 ( .B1(n15067), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15068), .ZN(n15312) );
  NAND2_X1 U18259 ( .A1(n15069), .A2(n15080), .ZN(n15071) );
  MUX2_X1 U18260 ( .A(n15080), .B(n15071), .S(n15070), .Z(n15072) );
  AND2_X1 U18261 ( .A1(n12169), .A2(n15072), .ZN(n15310) );
  AND2_X1 U18262 ( .A1(n19206), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15304) );
  NOR2_X1 U18263 ( .A1(n16113), .A2(n19205), .ZN(n15073) );
  AOI211_X1 U18264 ( .C1(n19190), .C2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n15304), .B(n15073), .ZN(n15074) );
  OAI21_X1 U18265 ( .B1(n16108), .B2(n16186), .A(n15074), .ZN(n15075) );
  AOI21_X1 U18266 ( .B1(n15310), .B2(n16190), .A(n15075), .ZN(n15076) );
  OAI21_X1 U18267 ( .B1(n15312), .B2(n19197), .A(n15076), .ZN(P2_U2988) );
  INV_X1 U18268 ( .A(n15067), .ZN(n15078) );
  OAI21_X1 U18269 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n15077), .A(
        n15078), .ZN(n15324) );
  INV_X1 U18270 ( .A(n15080), .ZN(n15081) );
  NOR2_X1 U18271 ( .A1(n15082), .A2(n15081), .ZN(n15083) );
  XNOR2_X1 U18272 ( .A(n15079), .B(n15083), .ZN(n15322) );
  NOR2_X1 U18273 ( .A1(n16123), .A2(n16186), .ZN(n15086) );
  NAND2_X1 U18274 ( .A1(n19206), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15314) );
  NAND2_X1 U18275 ( .A1(n19190), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15084) );
  OAI211_X1 U18276 ( .C1(n16127), .C2(n19205), .A(n15314), .B(n15084), .ZN(
        n15085) );
  AOI211_X1 U18277 ( .C1(n15322), .C2(n16190), .A(n15086), .B(n15085), .ZN(
        n15087) );
  OAI21_X1 U18278 ( .B1(n15324), .B2(n19197), .A(n15087), .ZN(P2_U2989) );
  XNOR2_X1 U18279 ( .A(n15089), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15090) );
  XNOR2_X1 U18280 ( .A(n15088), .B(n15090), .ZN(n15336) );
  AOI21_X1 U18281 ( .B1(n15092), .B2(n15091), .A(n15077), .ZN(n15325) );
  NAND2_X1 U18282 ( .A1(n15325), .A2(n16188), .ZN(n15096) );
  NAND2_X1 U18283 ( .A1(n19206), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n15331) );
  NAND2_X1 U18284 ( .A1(n19190), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15093) );
  OAI211_X1 U18285 ( .C1(n16136), .C2(n19205), .A(n15331), .B(n15093), .ZN(
        n15094) );
  AOI21_X1 U18286 ( .B1(n16133), .B2(n19201), .A(n15094), .ZN(n15095) );
  OAI211_X1 U18287 ( .C1(n15336), .C2(n19198), .A(n15096), .B(n15095), .ZN(
        P2_U2990) );
  OAI21_X1 U18288 ( .B1(n9739), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15091), .ZN(n15348) );
  NAND2_X1 U18289 ( .A1(n15098), .A2(n15111), .ZN(n15099) );
  NAND2_X1 U18290 ( .A1(n15099), .A2(n15110), .ZN(n15100) );
  XOR2_X1 U18291 ( .A(n15101), .B(n15100), .Z(n15346) );
  NOR2_X1 U18292 ( .A1(n19012), .A2(n15102), .ZN(n15340) );
  NOR2_X1 U18293 ( .A1(n15103), .A2(n19205), .ZN(n15104) );
  AOI211_X1 U18294 ( .C1(n19190), .C2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n15340), .B(n15104), .ZN(n15105) );
  OAI21_X1 U18295 ( .B1(n15344), .B2(n16186), .A(n15105), .ZN(n15106) );
  AOI21_X1 U18296 ( .B1(n15346), .B2(n16190), .A(n15106), .ZN(n15107) );
  OAI21_X1 U18297 ( .B1(n15348), .B2(n19197), .A(n15107), .ZN(P2_U2991) );
  BUF_X1 U18298 ( .A(n15108), .Z(n15109) );
  OAI21_X1 U18299 ( .B1(n15109), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n15097), .ZN(n15360) );
  NAND2_X1 U18300 ( .A1(n15111), .A2(n15110), .ZN(n15112) );
  XNOR2_X1 U18301 ( .A(n15098), .B(n15112), .ZN(n15358) );
  NOR2_X1 U18302 ( .A1(n19012), .A2(n19783), .ZN(n15351) );
  NOR2_X1 U18303 ( .A1(n15113), .A2(n19205), .ZN(n15114) );
  AOI211_X1 U18304 ( .C1(n19190), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15351), .B(n15114), .ZN(n15115) );
  OAI21_X1 U18305 ( .B1(n15356), .B2(n16186), .A(n15115), .ZN(n15116) );
  AOI21_X1 U18306 ( .B1(n15358), .B2(n16190), .A(n15116), .ZN(n15117) );
  OAI21_X1 U18307 ( .B1(n15360), .B2(n19197), .A(n15117), .ZN(P2_U2992) );
  NAND2_X1 U18308 ( .A1(n15119), .A2(n15118), .ZN(n15133) );
  AND3_X1 U18309 ( .A1(n15121), .A2(n9825), .A3(n15184), .ZN(n15122) );
  NAND3_X1 U18310 ( .A1(n15123), .A2(n15185), .A3(n15447), .ZN(n15125) );
  NAND2_X1 U18311 ( .A1(n15125), .A2(n15124), .ZN(n15126) );
  NAND2_X1 U18312 ( .A1(n15126), .A2(n15449), .ZN(n15165) );
  INV_X1 U18313 ( .A(n15164), .ZN(n15127) );
  NAND2_X1 U18314 ( .A1(n15404), .A2(n15389), .ZN(n15129) );
  AND2_X1 U18315 ( .A1(n15131), .A2(n15130), .ZN(n15142) );
  NAND2_X1 U18316 ( .A1(n15143), .A2(n15142), .ZN(n15374) );
  NAND2_X1 U18317 ( .A1(n15374), .A2(n15131), .ZN(n15132) );
  NAND2_X1 U18318 ( .A1(n19206), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15362) );
  NAND2_X1 U18319 ( .A1(n19190), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15134) );
  OAI211_X1 U18320 ( .C1(n15135), .C2(n19205), .A(n15362), .B(n15134), .ZN(
        n15136) );
  AOI21_X1 U18321 ( .B1(n15361), .B2(n19201), .A(n15136), .ZN(n15140) );
  AOI21_X1 U18323 ( .B1(n15367), .B2(n15138), .A(n15109), .ZN(n15370) );
  NAND2_X1 U18324 ( .A1(n15370), .A2(n16188), .ZN(n15139) );
  OAI211_X1 U18325 ( .C1(n15372), .C2(n19198), .A(n15140), .B(n15139), .ZN(
        P2_U2993) );
  OAI21_X1 U18326 ( .B1(n15141), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15138), .ZN(n15385) );
  NOR2_X1 U18327 ( .A1(n15143), .A2(n15142), .ZN(n15373) );
  NOR2_X1 U18328 ( .A1(n15373), .A2(n19198), .ZN(n15147) );
  AOI22_X1 U18329 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n19190), .B1(
        n16187), .B2(n15144), .ZN(n15145) );
  NAND2_X1 U18330 ( .A1(n19206), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n15377) );
  OAI211_X1 U18331 ( .C1(n15380), .C2(n16186), .A(n15145), .B(n15377), .ZN(
        n15146) );
  AOI21_X1 U18332 ( .B1(n15147), .B2(n15374), .A(n15146), .ZN(n15148) );
  OAI21_X1 U18333 ( .B1(n19197), .B2(n15385), .A(n15148), .ZN(P2_U2994) );
  NAND2_X1 U18334 ( .A1(n15150), .A2(n15149), .ZN(n15154) );
  NAND2_X1 U18335 ( .A1(n15152), .A2(n15151), .ZN(n15153) );
  XNOR2_X1 U18336 ( .A(n15154), .B(n15153), .ZN(n15431) );
  NAND2_X1 U18337 ( .A1(n19206), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15428) );
  INV_X1 U18338 ( .A(n15155), .ZN(n18924) );
  OAI22_X1 U18339 ( .A1(n15156), .A2(n16194), .B1(n19205), .B2(n18924), .ZN(
        n15157) );
  INV_X1 U18340 ( .A(n15157), .ZN(n15158) );
  OAI211_X1 U18341 ( .C1(n18925), .C2(n16186), .A(n15428), .B(n15158), .ZN(
        n15162) );
  AND2_X2 U18342 ( .A1(n15172), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15457) );
  NAND2_X1 U18343 ( .A1(n15457), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15418) );
  INV_X1 U18344 ( .A(n15159), .ZN(n15160) );
  NOR2_X1 U18345 ( .A1(n15160), .A2(n15407), .ZN(n15402) );
  AOI211_X1 U18346 ( .C1(n21010), .C2(n15418), .A(n19197), .B(n15402), .ZN(
        n15161) );
  AOI211_X1 U18347 ( .C1(n16190), .C2(n15431), .A(n15162), .B(n15161), .ZN(
        n15163) );
  INV_X1 U18348 ( .A(n15163), .ZN(P2_U2997) );
  XNOR2_X1 U18349 ( .A(n15165), .B(n15164), .ZN(n15443) );
  INV_X1 U18350 ( .A(n15443), .ZN(n15171) );
  OAI211_X1 U18351 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15457), .A(
        n15418), .B(n16188), .ZN(n15170) );
  INV_X1 U18352 ( .A(n18938), .ZN(n15168) );
  NAND2_X1 U18353 ( .A1(n19206), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n15440) );
  NAND2_X1 U18354 ( .A1(n19190), .A2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15166) );
  OAI211_X1 U18355 ( .C1(n19205), .C2(n18932), .A(n15440), .B(n15166), .ZN(
        n15167) );
  AOI21_X1 U18356 ( .B1(n15168), .B2(n19201), .A(n15167), .ZN(n15169) );
  OAI211_X1 U18357 ( .C1(n15171), .C2(n19198), .A(n15170), .B(n15169), .ZN(
        P2_U2998) );
  NAND2_X1 U18358 ( .A1(n15159), .A2(n15432), .ZN(n15182) );
  INV_X1 U18359 ( .A(n15182), .ZN(n15173) );
  INV_X1 U18360 ( .A(n15172), .ZN(n15458) );
  OAI21_X1 U18361 ( .B1(n15173), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15458), .ZN(n15479) );
  NAND2_X1 U18362 ( .A1(n15174), .A2(n15184), .ZN(n15177) );
  NAND2_X1 U18363 ( .A1(n15447), .A2(n15175), .ZN(n15176) );
  NAND2_X1 U18364 ( .A1(n15177), .A2(n15176), .ZN(n15178) );
  NAND2_X1 U18365 ( .A1(n15448), .A2(n15178), .ZN(n15476) );
  OAI22_X1 U18366 ( .A1(n10855), .A2(n19012), .B1(n19205), .B2(n18944), .ZN(
        n15180) );
  OAI22_X1 U18367 ( .A1(n18949), .A2(n16186), .B1(n9997), .B2(n16194), .ZN(
        n15179) );
  AOI211_X1 U18368 ( .C1(n15476), .C2(n16190), .A(n15180), .B(n15179), .ZN(
        n15181) );
  OAI21_X1 U18369 ( .B1(n19197), .B2(n15479), .A(n15181), .ZN(P2_U3000) );
  NOR2_X2 U18370 ( .A1(n16175), .A2(n16207), .ZN(n15223) );
  NAND2_X1 U18371 ( .A1(n15223), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15203) );
  NOR2_X1 U18372 ( .A1(n15203), .A2(n15194), .ZN(n15193) );
  OAI21_X1 U18373 ( .B1(n15193), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15182), .ZN(n15493) );
  NAND2_X1 U18374 ( .A1(n15185), .A2(n15184), .ZN(n15186) );
  XNOR2_X1 U18375 ( .A(n15183), .B(n15186), .ZN(n15491) );
  OAI22_X1 U18376 ( .A1(n16194), .A2(n15188), .B1(n15187), .B2(n19012), .ZN(
        n15189) );
  AOI21_X1 U18377 ( .B1(n16187), .B2(n18959), .A(n15189), .ZN(n15190) );
  OAI21_X1 U18378 ( .B1(n15482), .B2(n16186), .A(n15190), .ZN(n15191) );
  AOI21_X1 U18379 ( .B1(n15491), .B2(n16190), .A(n15191), .ZN(n15192) );
  OAI21_X1 U18380 ( .B1(n15493), .B2(n19197), .A(n15192), .ZN(P2_U3001) );
  AOI21_X1 U18381 ( .B1(n15194), .B2(n15203), .A(n15193), .ZN(n16201) );
  AND2_X1 U18382 ( .A1(n9825), .A2(n15196), .ZN(n15197) );
  XNOR2_X1 U18383 ( .A(n15195), .B(n15197), .ZN(n16204) );
  AOI22_X1 U18384 ( .A1(n18970), .A2(n19201), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19190), .ZN(n15200) );
  OAI22_X1 U18385 ( .A1(n10848), .A2(n19012), .B1(n19205), .B2(n18967), .ZN(
        n15198) );
  INV_X1 U18386 ( .A(n15198), .ZN(n15199) );
  OAI211_X1 U18387 ( .C1(n16204), .C2(n19198), .A(n15200), .B(n15199), .ZN(
        n15201) );
  AOI21_X1 U18388 ( .B1(n16201), .B2(n16188), .A(n15201), .ZN(n15202) );
  INV_X1 U18389 ( .A(n15202), .ZN(P2_U3002) );
  OAI21_X1 U18390 ( .B1(n15223), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15203), .ZN(n15507) );
  INV_X1 U18391 ( .A(n15204), .ZN(n15206) );
  NAND2_X1 U18392 ( .A1(n15206), .A2(n15205), .ZN(n15210) );
  NAND2_X1 U18393 ( .A1(n15208), .A2(n15207), .ZN(n15209) );
  XNOR2_X1 U18394 ( .A(n15210), .B(n15209), .ZN(n15504) );
  NAND2_X1 U18395 ( .A1(n19206), .A2(P2_REIP_REG_11__SCAN_IN), .ZN(n15496) );
  OAI21_X1 U18396 ( .B1(n16194), .B2(n15211), .A(n15496), .ZN(n15212) );
  AOI21_X1 U18397 ( .B1(n16187), .B2(n15213), .A(n15212), .ZN(n15214) );
  OAI21_X1 U18398 ( .B1(n15497), .B2(n16186), .A(n15214), .ZN(n15215) );
  AOI21_X1 U18399 ( .B1(n15504), .B2(n16190), .A(n15215), .ZN(n15216) );
  OAI21_X1 U18400 ( .B1(n15507), .B2(n19197), .A(n15216), .ZN(P2_U3003) );
  INV_X1 U18401 ( .A(n15509), .ZN(n15218) );
  NAND2_X1 U18402 ( .A1(n15217), .A2(n15218), .ZN(n15222) );
  NOR2_X1 U18403 ( .A1(n15220), .A2(n15219), .ZN(n15221) );
  XNOR2_X1 U18404 ( .A(n15222), .B(n15221), .ZN(n16214) );
  AOI21_X1 U18405 ( .B1(n16207), .B2(n16175), .A(n15223), .ZN(n16211) );
  NAND2_X1 U18406 ( .A1(n16211), .A2(n16188), .ZN(n15228) );
  NAND2_X1 U18407 ( .A1(P2_REIP_REG_10__SCAN_IN), .A2(n19206), .ZN(n16205) );
  INV_X1 U18408 ( .A(n16205), .ZN(n15226) );
  INV_X1 U18409 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n20784) );
  OAI22_X1 U18410 ( .A1(n20784), .A2(n16194), .B1(n19205), .B2(n15224), .ZN(
        n15225) );
  AOI211_X1 U18411 ( .C1(n16210), .C2(n19201), .A(n15226), .B(n15225), .ZN(
        n15227) );
  OAI211_X1 U18412 ( .C1(n16214), .C2(n19198), .A(n15228), .B(n15227), .ZN(
        P2_U3004) );
  OAI21_X1 U18413 ( .B1(n15229), .B2(n15231), .A(n15230), .ZN(n15232) );
  INV_X1 U18414 ( .A(n15232), .ZN(n16224) );
  INV_X1 U18415 ( .A(n15233), .ZN(n15236) );
  INV_X1 U18416 ( .A(n15234), .ZN(n15235) );
  NAND2_X1 U18417 ( .A1(n15236), .A2(n15235), .ZN(n15254) );
  XNOR2_X1 U18418 ( .A(n15237), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15253) );
  NAND2_X1 U18419 ( .A1(n15254), .A2(n15253), .ZN(n15239) );
  NAND2_X1 U18420 ( .A1(n15239), .A2(n15238), .ZN(n15530) );
  NAND2_X1 U18421 ( .A1(n15530), .A2(n15527), .ZN(n15240) );
  NAND2_X1 U18422 ( .A1(n15240), .A2(n15528), .ZN(n15244) );
  AND2_X1 U18423 ( .A1(n15242), .A2(n15241), .ZN(n15243) );
  XNOR2_X1 U18424 ( .A(n15244), .B(n15243), .ZN(n16228) );
  AOI22_X1 U18425 ( .A1(n16222), .A2(n19201), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n19190), .ZN(n15248) );
  OAI22_X1 U18426 ( .A1(n10830), .A2(n19012), .B1(n19205), .B2(n15245), .ZN(
        n15246) );
  INV_X1 U18427 ( .A(n15246), .ZN(n15247) );
  OAI211_X1 U18428 ( .C1(n16228), .C2(n19198), .A(n15248), .B(n15247), .ZN(
        n15249) );
  AOI21_X1 U18429 ( .B1(n16224), .B2(n16188), .A(n15249), .ZN(n15250) );
  INV_X1 U18430 ( .A(n15250), .ZN(P2_U3006) );
  OAI21_X1 U18431 ( .B1(n15252), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15251), .ZN(n15554) );
  NOR2_X1 U18432 ( .A1(n15554), .A2(n19197), .ZN(n15259) );
  XNOR2_X1 U18433 ( .A(n15254), .B(n15253), .ZN(n15551) );
  AOI22_X1 U18434 ( .A1(n19201), .A2(n19008), .B1(n19190), .B2(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n15257) );
  INV_X1 U18435 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19765) );
  OAI22_X1 U18436 ( .A1(n19765), .A2(n19012), .B1(n19205), .B2(n19006), .ZN(
        n15255) );
  INV_X1 U18437 ( .A(n15255), .ZN(n15256) );
  OAI211_X1 U18438 ( .C1(n15551), .C2(n19198), .A(n15257), .B(n15256), .ZN(
        n15258) );
  OR2_X1 U18439 ( .A1(n15259), .A2(n15258), .ZN(P2_U3008) );
  NOR2_X1 U18440 ( .A1(n15262), .A2(n15261), .ZN(n15267) );
  INV_X1 U18441 ( .A(n15263), .ZN(n15265) );
  OAI21_X1 U18442 ( .B1(n15265), .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n15264), .ZN(n15266) );
  NOR2_X1 U18443 ( .A1(n15267), .A2(n15266), .ZN(n15268) );
  OAI211_X1 U18444 ( .C1(n15270), .C2(n15520), .A(n15269), .B(n15268), .ZN(
        n15271) );
  AOI21_X1 U18445 ( .B1(n15272), .B2(n19219), .A(n15271), .ZN(n15273) );
  OAI21_X1 U18446 ( .B1(n19215), .B2(n15274), .A(n15273), .ZN(P2_U3016) );
  INV_X1 U18447 ( .A(n15275), .ZN(n16076) );
  NOR2_X1 U18448 ( .A1(n15276), .A2(n15277), .ZN(n15284) );
  INV_X1 U18449 ( .A(n16075), .ZN(n15282) );
  NAND3_X1 U18450 ( .A1(n15279), .A2(n15278), .A3(n15277), .ZN(n15281) );
  OAI211_X1 U18451 ( .C1(n15282), .C2(n16197), .A(n15281), .B(n15280), .ZN(
        n15283) );
  AOI211_X1 U18452 ( .C1(n16076), .C2(n19212), .A(n15284), .B(n15283), .ZN(
        n15287) );
  NAND2_X1 U18453 ( .A1(n15285), .A2(n16223), .ZN(n15286) );
  OAI211_X1 U18454 ( .C1(n15288), .C2(n16227), .A(n15287), .B(n15286), .ZN(
        P2_U3017) );
  NAND2_X1 U18455 ( .A1(n15289), .A2(n16223), .ZN(n15300) );
  NAND3_X1 U18456 ( .A1(n15290), .A2(n19219), .A3(n15058), .ZN(n15299) );
  OAI21_X1 U18457 ( .B1(n15292), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15291), .ZN(n15293) );
  AOI21_X1 U18458 ( .B1(n19208), .B2(n16097), .A(n15293), .ZN(n15296) );
  NAND2_X1 U18459 ( .A1(n15294), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15295) );
  OAI211_X1 U18460 ( .C1(n16096), .C2(n15520), .A(n15296), .B(n15295), .ZN(
        n15297) );
  INV_X1 U18461 ( .A(n15297), .ZN(n15298) );
  OAI211_X1 U18462 ( .C1(n15301), .C2(n15300), .A(n15299), .B(n15298), .ZN(
        P2_U3019) );
  NOR2_X1 U18463 ( .A1(n16108), .A2(n15520), .ZN(n15309) );
  XNOR2_X1 U18464 ( .A(n15307), .B(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15305) );
  NOR2_X1 U18465 ( .A1(n16197), .A2(n15302), .ZN(n15303) );
  AOI211_X1 U18466 ( .C1(n15313), .C2(n15305), .A(n15304), .B(n15303), .ZN(
        n15306) );
  OAI21_X1 U18467 ( .B1(n15317), .B2(n15307), .A(n15306), .ZN(n15308) );
  AOI211_X1 U18468 ( .C1(n15310), .C2(n19219), .A(n15309), .B(n15308), .ZN(
        n15311) );
  OAI21_X1 U18469 ( .B1(n19215), .B2(n15312), .A(n15311), .ZN(P2_U3020) );
  INV_X1 U18470 ( .A(n15313), .ZN(n15315) );
  OAI21_X1 U18471 ( .B1(n15315), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n15314), .ZN(n15319) );
  NOR2_X1 U18472 ( .A1(n15317), .A2(n15316), .ZN(n15318) );
  AOI211_X1 U18473 ( .C1(n19208), .C2(n16121), .A(n15319), .B(n15318), .ZN(
        n15320) );
  OAI21_X1 U18474 ( .B1(n16123), .B2(n15520), .A(n15320), .ZN(n15321) );
  AOI21_X1 U18475 ( .B1(n15322), .B2(n19219), .A(n15321), .ZN(n15323) );
  OAI21_X1 U18476 ( .B1(n15324), .B2(n19215), .A(n15323), .ZN(P2_U3021) );
  NAND2_X1 U18477 ( .A1(n15325), .A2(n16223), .ZN(n15335) );
  NAND2_X1 U18478 ( .A1(n14735), .A2(n15326), .ZN(n15327) );
  NAND2_X1 U18479 ( .A1(n9792), .A2(n15327), .ZN(n16142) );
  NOR2_X1 U18480 ( .A1(n15349), .A2(n15328), .ZN(n15330) );
  OAI21_X1 U18481 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15330), .A(
        n15329), .ZN(n15332) );
  OAI211_X1 U18482 ( .C1(n16197), .C2(n16142), .A(n15332), .B(n15331), .ZN(
        n15333) );
  AOI21_X1 U18483 ( .B1(n16133), .B2(n19212), .A(n15333), .ZN(n15334) );
  OAI211_X1 U18484 ( .C1(n15336), .C2(n16227), .A(n15335), .B(n15334), .ZN(
        P2_U3022) );
  AOI211_X1 U18485 ( .C1(n10098), .C2(n15338), .A(n15337), .B(n15349), .ZN(
        n15339) );
  AOI211_X1 U18486 ( .C1(n19208), .C2(n15341), .A(n15340), .B(n15339), .ZN(
        n15343) );
  NAND2_X1 U18487 ( .A1(n15353), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15342) );
  OAI211_X1 U18488 ( .C1(n15344), .C2(n15520), .A(n15343), .B(n15342), .ZN(
        n15345) );
  AOI21_X1 U18489 ( .B1(n15346), .B2(n19219), .A(n15345), .ZN(n15347) );
  OAI21_X1 U18490 ( .B1(n15348), .B2(n19215), .A(n15347), .ZN(P2_U3023) );
  NOR2_X1 U18491 ( .A1(n15349), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15350) );
  AOI211_X1 U18492 ( .C1(n19208), .C2(n15352), .A(n15351), .B(n15350), .ZN(
        n15355) );
  NAND2_X1 U18493 ( .A1(n15353), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15354) );
  OAI211_X1 U18494 ( .C1(n15356), .C2(n15520), .A(n15355), .B(n15354), .ZN(
        n15357) );
  AOI21_X1 U18495 ( .B1(n15358), .B2(n19219), .A(n15357), .ZN(n15359) );
  OAI21_X1 U18496 ( .B1(n15360), .B2(n19215), .A(n15359), .ZN(P2_U3024) );
  NAND2_X1 U18497 ( .A1(n15361), .A2(n19212), .ZN(n15366) );
  OAI21_X1 U18498 ( .B1(n15363), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15362), .ZN(n15364) );
  AOI21_X1 U18499 ( .B1(n19208), .B2(n16149), .A(n15364), .ZN(n15365) );
  OAI211_X1 U18500 ( .C1(n15368), .C2(n15367), .A(n15366), .B(n15365), .ZN(
        n15369) );
  AOI21_X1 U18501 ( .B1(n15370), .B2(n16223), .A(n15369), .ZN(n15371) );
  OAI21_X1 U18502 ( .B1(n15372), .B2(n16227), .A(n15371), .ZN(P2_U3025) );
  INV_X1 U18503 ( .A(n15373), .ZN(n15375) );
  NAND3_X1 U18504 ( .A1(n15375), .A2(n19219), .A3(n15374), .ZN(n15384) );
  XNOR2_X1 U18505 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15379) );
  NAND2_X1 U18506 ( .A1(n19208), .A2(n15376), .ZN(n15378) );
  OAI211_X1 U18507 ( .C1(n15394), .C2(n15379), .A(n15378), .B(n15377), .ZN(
        n15382) );
  NOR2_X1 U18508 ( .A1(n15380), .A2(n15520), .ZN(n15381) );
  AOI211_X1 U18509 ( .C1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n15396), .A(
        n15382), .B(n15381), .ZN(n15383) );
  OAI211_X1 U18510 ( .C1(n15385), .C2(n19215), .A(n15384), .B(n15383), .ZN(
        P2_U3026) );
  INV_X1 U18511 ( .A(n15404), .ZN(n15386) );
  NOR2_X1 U18512 ( .A1(n15387), .A2(n15386), .ZN(n15391) );
  NAND2_X1 U18513 ( .A1(n15389), .A2(n15388), .ZN(n15390) );
  XNOR2_X1 U18514 ( .A(n15391), .B(n15390), .ZN(n16156) );
  INV_X1 U18515 ( .A(n16156), .ZN(n15401) );
  AOI21_X1 U18516 ( .B1(n15393), .B2(n15392), .A(n15141), .ZN(n16155) );
  OAI22_X1 U18517 ( .A1(n15394), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B1(
        n10877), .B2(n19012), .ZN(n15395) );
  AOI21_X1 U18518 ( .B1(n19208), .B2(n18910), .A(n15395), .ZN(n15398) );
  NAND2_X1 U18519 ( .A1(n15396), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15397) );
  OAI211_X1 U18520 ( .C1(n18912), .C2(n15520), .A(n15398), .B(n15397), .ZN(
        n15399) );
  AOI21_X1 U18521 ( .B1(n16155), .B2(n16223), .A(n15399), .ZN(n15400) );
  OAI21_X1 U18522 ( .B1(n15401), .B2(n16227), .A(n15400), .ZN(P2_U3027) );
  OAI21_X1 U18523 ( .B1(n15402), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15392), .ZN(n16160) );
  NAND2_X1 U18524 ( .A1(n15404), .A2(n15403), .ZN(n15405) );
  XNOR2_X1 U18525 ( .A(n15406), .B(n15405), .ZN(n16159) );
  INV_X1 U18526 ( .A(n16159), .ZN(n15416) );
  OR2_X1 U18527 ( .A1(n15407), .A2(n15469), .ZN(n15411) );
  NAND2_X1 U18528 ( .A1(P2_REIP_REG_18__SCAN_IN), .A2(n19206), .ZN(n15408) );
  OAI221_X1 U18529 ( .B1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15411), 
        .C1(n15410), .C2(n15409), .A(n15408), .ZN(n15415) );
  OAI22_X1 U18530 ( .A1(n15413), .A2(n15520), .B1(n16197), .B2(n15412), .ZN(
        n15414) );
  AOI211_X1 U18531 ( .C1(n15416), .C2(n19219), .A(n15415), .B(n15414), .ZN(
        n15417) );
  OAI21_X1 U18532 ( .B1(n19215), .B2(n16160), .A(n15417), .ZN(P2_U3028) );
  OAI21_X1 U18533 ( .B1(n16223), .B2(n15419), .A(n15418), .ZN(n15424) );
  INV_X1 U18534 ( .A(n15420), .ZN(n15421) );
  NAND2_X1 U18535 ( .A1(n15426), .A2(n15421), .ZN(n15422) );
  NAND2_X1 U18536 ( .A1(n15468), .A2(n15422), .ZN(n15459) );
  INV_X1 U18537 ( .A(n15459), .ZN(n15423) );
  OAI211_X1 U18538 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15425), .A(
        n15424), .B(n15423), .ZN(n15439) );
  AOI21_X1 U18539 ( .B1(n15427), .B2(n15426), .A(n15439), .ZN(n15437) );
  NOR2_X1 U18540 ( .A1(n18925), .A2(n15520), .ZN(n15430) );
  OAI21_X1 U18541 ( .B1(n16197), .B2(n18930), .A(n15428), .ZN(n15429) );
  AOI211_X1 U18542 ( .C1(n15431), .C2(n19219), .A(n15430), .B(n15429), .ZN(
        n15436) );
  NAND2_X1 U18543 ( .A1(n15457), .A2(n16223), .ZN(n15434) );
  NAND2_X1 U18544 ( .A1(n15432), .A2(n15498), .ZN(n15472) );
  INV_X1 U18545 ( .A(n15472), .ZN(n15453) );
  NAND3_X1 U18546 ( .A1(n15453), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15433) );
  NAND2_X1 U18547 ( .A1(n15434), .A2(n15433), .ZN(n15438) );
  NAND3_X1 U18548 ( .A1(n15438), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n21010), .ZN(n15435) );
  OAI211_X1 U18549 ( .C1(n15437), .C2(n21010), .A(n15436), .B(n15435), .ZN(
        P2_U3029) );
  INV_X1 U18550 ( .A(n15438), .ZN(n15446) );
  NAND2_X1 U18551 ( .A1(n15439), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15445) );
  NOR2_X1 U18552 ( .A1(n18938), .A2(n15520), .ZN(n15442) );
  OAI21_X1 U18553 ( .B1(n16197), .B2(n18937), .A(n15440), .ZN(n15441) );
  AOI211_X1 U18554 ( .C1(n15443), .C2(n19219), .A(n15442), .B(n15441), .ZN(
        n15444) );
  OAI211_X1 U18555 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15446), .A(
        n15445), .B(n15444), .ZN(P2_U3030) );
  NAND2_X1 U18556 ( .A1(n15448), .A2(n15447), .ZN(n15452) );
  NAND2_X1 U18557 ( .A1(n15450), .A2(n15449), .ZN(n15451) );
  XOR2_X1 U18558 ( .A(n15452), .B(n15451), .Z(n16169) );
  NAND2_X1 U18559 ( .A1(n16169), .A2(n19219), .ZN(n15463) );
  OR2_X1 U18560 ( .A1(n10863), .A2(n19012), .ZN(n15455) );
  NAND3_X1 U18561 ( .A1(n15453), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n20957), .ZN(n15454) );
  OAI211_X1 U18562 ( .C1(n16197), .C2(n19053), .A(n15455), .B(n15454), .ZN(
        n15456) );
  AOI21_X1 U18563 ( .B1(n16167), .B2(n19212), .A(n15456), .ZN(n15462) );
  AOI21_X1 U18564 ( .B1(n20957), .B2(n15458), .A(n15457), .ZN(n16168) );
  NAND2_X1 U18565 ( .A1(n16168), .A2(n16223), .ZN(n15461) );
  NAND2_X1 U18566 ( .A1(n15459), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15460) );
  NAND4_X1 U18567 ( .A1(n15463), .A2(n15462), .A3(n15461), .A4(n15460), .ZN(
        P2_U3031) );
  INV_X1 U18568 ( .A(n18949), .ZN(n15475) );
  NAND2_X1 U18569 ( .A1(n15465), .A2(n15464), .ZN(n15467) );
  NAND2_X1 U18570 ( .A1(n15467), .A2(n15466), .ZN(n19055) );
  OAI22_X1 U18571 ( .A1(n16197), .A2(n19055), .B1(n10855), .B2(n19012), .ZN(
        n15474) );
  NAND3_X1 U18572 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15499), .A3(
        n15498), .ZN(n15470) );
  NOR2_X1 U18573 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15470), .ZN(
        n16199) );
  INV_X1 U18574 ( .A(n15468), .ZN(n15522) );
  NOR2_X1 U18575 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15469), .ZN(
        n15517) );
  NOR2_X1 U18576 ( .A1(n15522), .A2(n15517), .ZN(n16206) );
  OAI21_X1 U18577 ( .B1(n15499), .B2(n15556), .A(n16206), .ZN(n16200) );
  NOR2_X1 U18578 ( .A1(n16199), .A2(n16200), .ZN(n15489) );
  NOR2_X1 U18579 ( .A1(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15470), .ZN(
        n15486) );
  NOR2_X1 U18580 ( .A1(n20881), .A2(n15486), .ZN(n15471) );
  AOI22_X1 U18581 ( .A1(n15472), .A2(n20881), .B1(n15489), .B2(n15471), .ZN(
        n15473) );
  AOI211_X1 U18582 ( .C1(n15475), .C2(n19212), .A(n15474), .B(n15473), .ZN(
        n15478) );
  NAND2_X1 U18583 ( .A1(n15476), .A2(n19219), .ZN(n15477) );
  OAI211_X1 U18584 ( .C1(n15479), .C2(n19215), .A(n15478), .B(n15477), .ZN(
        P2_U3032) );
  OAI21_X1 U18585 ( .B1(n15481), .B2(n15480), .A(n15464), .ZN(n19057) );
  INV_X1 U18586 ( .A(n15482), .ZN(n18961) );
  NOR2_X1 U18587 ( .A1(n15187), .A2(n19012), .ZN(n15483) );
  AOI21_X1 U18588 ( .B1(n18961), .B2(n19212), .A(n15483), .ZN(n15484) );
  OAI21_X1 U18589 ( .B1(n16197), .B2(n19057), .A(n15484), .ZN(n15485) );
  AOI21_X1 U18590 ( .B1(n15486), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15485), .ZN(n15487) );
  OAI21_X1 U18591 ( .B1(n15489), .B2(n15488), .A(n15487), .ZN(n15490) );
  AOI21_X1 U18592 ( .B1(n15491), .B2(n19219), .A(n15490), .ZN(n15492) );
  OAI21_X1 U18593 ( .B1(n15493), .B2(n19215), .A(n15492), .ZN(P2_U3033) );
  INV_X1 U18594 ( .A(n16206), .ZN(n15503) );
  INV_X1 U18595 ( .A(n19061), .ZN(n15494) );
  NAND2_X1 U18596 ( .A1(n19208), .A2(n15494), .ZN(n15495) );
  OAI211_X1 U18597 ( .C1(n15497), .C2(n15520), .A(n15496), .B(n15495), .ZN(
        n15502) );
  NAND2_X1 U18598 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15498), .ZN(
        n16208) );
  AOI211_X1 U18599 ( .C1(n16207), .C2(n15500), .A(n15499), .B(n16208), .ZN(
        n15501) );
  AOI211_X1 U18600 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15503), .A(
        n15502), .B(n15501), .ZN(n15506) );
  NAND2_X1 U18601 ( .A1(n15504), .A2(n19219), .ZN(n15505) );
  OAI211_X1 U18602 ( .C1(n15507), .C2(n19215), .A(n15506), .B(n15505), .ZN(
        P2_U3035) );
  NOR2_X1 U18603 ( .A1(n15509), .A2(n15508), .ZN(n15511) );
  XOR2_X1 U18604 ( .A(n15511), .B(n15510), .Z(n16173) );
  NOR2_X1 U18605 ( .A1(n15159), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n16172) );
  INV_X1 U18606 ( .A(n16172), .ZN(n15512) );
  NAND3_X1 U18607 ( .A1(n15512), .A2(n16223), .A3(n16175), .ZN(n15524) );
  OR2_X1 U18608 ( .A1(n15513), .A2(n14825), .ZN(n15515) );
  NAND2_X1 U18609 ( .A1(n15515), .A2(n15514), .ZN(n19066) );
  INV_X1 U18610 ( .A(n19066), .ZN(n15518) );
  NOR2_X1 U18611 ( .A1(n10836), .A2(n19012), .ZN(n15516) );
  AOI211_X1 U18612 ( .C1(n19208), .C2(n15518), .A(n15517), .B(n15516), .ZN(
        n15519) );
  OAI21_X1 U18613 ( .B1(n18982), .B2(n15520), .A(n15519), .ZN(n15521) );
  AOI21_X1 U18614 ( .B1(n15522), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15521), .ZN(n15523) );
  OAI211_X1 U18615 ( .C1(n16173), .C2(n16227), .A(n15524), .B(n15523), .ZN(
        P2_U3037) );
  OAI21_X1 U18616 ( .B1(n15525), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n15526), .ZN(n16181) );
  NAND2_X1 U18617 ( .A1(n15528), .A2(n15527), .ZN(n15529) );
  XNOR2_X1 U18618 ( .A(n15530), .B(n15529), .ZN(n16182) );
  NAND2_X1 U18619 ( .A1(n16215), .A2(n15539), .ZN(n15538) );
  INV_X1 U18620 ( .A(n18993), .ZN(n15536) );
  NOR2_X1 U18621 ( .A1(n10824), .A2(n19012), .ZN(n15535) );
  OR2_X1 U18622 ( .A1(n15532), .A2(n15531), .ZN(n15533) );
  NAND2_X1 U18623 ( .A1(n15533), .A2(n14824), .ZN(n19071) );
  NOR2_X1 U18624 ( .A1(n16197), .A2(n19071), .ZN(n15534) );
  AOI211_X1 U18625 ( .C1(n15536), .C2(n19212), .A(n15535), .B(n15534), .ZN(
        n15537) );
  OAI211_X1 U18626 ( .C1(n16217), .C2(n15539), .A(n15538), .B(n15537), .ZN(
        n15540) );
  AOI21_X1 U18627 ( .B1(n16182), .B2(n19219), .A(n15540), .ZN(n15541) );
  OAI21_X1 U18628 ( .B1(n16181), .B2(n19215), .A(n15541), .ZN(P2_U3039) );
  NOR2_X1 U18629 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n19222), .ZN(
        n15550) );
  NOR2_X1 U18630 ( .A1(n19765), .A2(n19012), .ZN(n15542) );
  AOI21_X1 U18631 ( .B1(n19212), .B2(n19008), .A(n15542), .ZN(n15547) );
  XNOR2_X1 U18632 ( .A(n15544), .B(n15543), .ZN(n19073) );
  INV_X1 U18633 ( .A(n19073), .ZN(n15545) );
  NAND2_X1 U18634 ( .A1(n19208), .A2(n15545), .ZN(n15546) );
  OAI211_X1 U18635 ( .C1(n16217), .C2(n20868), .A(n15547), .B(n15546), .ZN(
        n15548) );
  AOI21_X1 U18636 ( .B1(n15550), .B2(n15549), .A(n15548), .ZN(n15553) );
  OR2_X1 U18637 ( .A1(n15551), .A2(n16227), .ZN(n15552) );
  OAI211_X1 U18638 ( .C1(n15554), .C2(n19215), .A(n15553), .B(n15552), .ZN(
        P2_U3040) );
  AOI211_X1 U18639 ( .C1(n15558), .C2(n15557), .A(n15556), .B(n15555), .ZN(
        n15559) );
  INV_X1 U18640 ( .A(n15559), .ZN(n15567) );
  OAI22_X1 U18641 ( .A1(n19215), .A2(n15561), .B1(n16227), .B2(n15560), .ZN(
        n15563) );
  AOI211_X1 U18642 ( .C1(n19208), .C2(n19833), .A(n15563), .B(n15562), .ZN(
        n15566) );
  AOI22_X1 U18643 ( .A1(n19212), .A2(n15568), .B1(n15564), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15565) );
  NAND3_X1 U18644 ( .A1(n15567), .A2(n15566), .A3(n15565), .ZN(P2_U3045) );
  NAND2_X1 U18645 ( .A1(n15568), .A2(n16241), .ZN(n15573) );
  NOR2_X1 U18646 ( .A1(n15569), .A2(n15580), .ZN(n15571) );
  AOI22_X1 U18647 ( .A1(n15571), .A2(n15570), .B1(n10775), .B2(n10198), .ZN(
        n15572) );
  NAND2_X1 U18648 ( .A1(n15573), .A2(n15572), .ZN(n16248) );
  INV_X1 U18649 ( .A(n19816), .ZN(n18875) );
  INV_X1 U18650 ( .A(n15574), .ZN(n15575) );
  NOR2_X1 U18651 ( .A1(n16287), .A2(n15575), .ZN(n15592) );
  AOI21_X1 U18652 ( .B1(n19005), .B2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n15576), .ZN(n15594) );
  AOI22_X1 U18653 ( .A1(n16248), .A2(n18875), .B1(n15592), .B2(n15594), .ZN(
        n15577) );
  OAI21_X1 U18654 ( .B1(n19838), .B2(n19810), .A(n15577), .ZN(n15578) );
  MUX2_X1 U18655 ( .A(n15578), .B(n16229), .S(n19811), .Z(P2_U3600) );
  NOR2_X1 U18656 ( .A1(n19825), .A2(n19810), .ZN(n15596) );
  INV_X1 U18657 ( .A(n10775), .ZN(n16237) );
  AOI21_X1 U18658 ( .B1(n16229), .B2(n10197), .A(n15579), .ZN(n15589) );
  NOR2_X1 U18659 ( .A1(n15580), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n15586) );
  NAND2_X1 U18660 ( .A1(n15582), .A2(n15581), .ZN(n16234) );
  OAI21_X1 U18661 ( .B1(n15583), .B2(n15586), .A(n16234), .ZN(n15588) );
  AOI21_X1 U18662 ( .B1(n15585), .B2(n15584), .A(n15583), .ZN(n16230) );
  INV_X1 U18663 ( .A(n15586), .ZN(n16233) );
  NAND2_X1 U18664 ( .A1(n16230), .A2(n16233), .ZN(n15587) );
  OAI211_X1 U18665 ( .C1(n16237), .C2(n15589), .A(n15588), .B(n15587), .ZN(
        n15590) );
  AOI21_X1 U18666 ( .B1(n15591), .B2(n16241), .A(n15590), .ZN(n16245) );
  INV_X1 U18667 ( .A(n15592), .ZN(n15593) );
  OAI22_X1 U18668 ( .A1(n16245), .A2(n19816), .B1(n15594), .B2(n15593), .ZN(
        n15595) );
  OAI21_X1 U18669 ( .B1(n15596), .B2(n15595), .A(n19813), .ZN(n15597) );
  OAI21_X1 U18670 ( .B1(n19813), .B2(n10197), .A(n15597), .ZN(P2_U3599) );
  AND4_X1 U18671 ( .A1(n10752), .A2(n10723), .A3(n16259), .A4(n18875), .ZN(
        n15598) );
  MUX2_X1 U18672 ( .A(n15598), .B(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n19811), .Z(P2_U3595) );
  NOR3_X1 U18673 ( .A1(n12371), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19389) );
  INV_X1 U18674 ( .A(n19389), .ZN(n19391) );
  NOR2_X1 U18675 ( .A1(n12376), .A2(n19391), .ZN(n19408) );
  AOI21_X1 U18676 ( .B1(n19432), .B2(n19459), .A(n19868), .ZN(n15599) );
  NAND2_X1 U18677 ( .A1(n19824), .A2(n19671), .ZN(n19434) );
  NOR2_X1 U18678 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19434), .ZN(
        n19427) );
  AOI221_X1 U18679 ( .B1(n19408), .B2(n19385), .C1(n15599), .C2(n19385), .A(
        n19427), .ZN(n15600) );
  NOR3_X1 U18680 ( .A1(n12008), .A2(n19427), .A3(n10692), .ZN(n15602) );
  OR3_X1 U18681 ( .A1(n15600), .A2(n19436), .A3(n15602), .ZN(n19429) );
  INV_X1 U18682 ( .A(n19429), .ZN(n15607) );
  INV_X1 U18683 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15606) );
  AOI22_X1 U18684 ( .A1(n19448), .A2(n19682), .B1(n19424), .B2(n19632), .ZN(
        n15605) );
  NOR2_X1 U18685 ( .A1(n19408), .A2(n19427), .ZN(n15601) );
  OR2_X1 U18686 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n15601), .ZN(n15603) );
  AOI21_X1 U18687 ( .B1(n10692), .B2(n15603), .A(n15602), .ZN(n19428) );
  AOI22_X1 U18688 ( .A1(n19428), .A2(n19674), .B1(n19673), .B2(n19427), .ZN(
        n15604) );
  OAI211_X1 U18689 ( .C1(n15607), .C2(n15606), .A(n15605), .B(n15604), .ZN(
        P2_U3096) );
  NAND2_X1 U18690 ( .A1(n12371), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19544) );
  NOR2_X1 U18691 ( .A1(n19261), .A2(n19544), .ZN(n19516) );
  AOI21_X1 U18692 ( .B1(n19577), .B2(n19537), .A(n19868), .ZN(n15609) );
  NOR2_X1 U18693 ( .A1(n19516), .A2(n15609), .ZN(n15610) );
  NOR2_X1 U18694 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n15610), .ZN(n15611) );
  OAI21_X1 U18695 ( .B1(n15614), .B2(n10692), .A(n15611), .ZN(n15612) );
  NOR2_X1 U18696 ( .A1(n19290), .A2(n19544), .ZN(n19538) );
  INV_X1 U18697 ( .A(n19538), .ZN(n15618) );
  NAND2_X1 U18698 ( .A1(n15612), .A2(n15618), .ZN(n15613) );
  NAND2_X1 U18699 ( .A1(n15613), .A2(n19680), .ZN(n19541) );
  INV_X1 U18700 ( .A(n19541), .ZN(n19525) );
  INV_X1 U18701 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15621) );
  INV_X1 U18702 ( .A(n19292), .ZN(n15616) );
  OAI21_X1 U18703 ( .B1(n15614), .B2(n19538), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15615) );
  OAI21_X1 U18704 ( .B1(n19544), .B2(n15616), .A(n15615), .ZN(n19539) );
  AOI22_X1 U18705 ( .A1(n19560), .A2(n19682), .B1(n19540), .B2(n19632), .ZN(
        n15617) );
  OAI21_X1 U18706 ( .B1(n15634), .B2(n15618), .A(n15617), .ZN(n15619) );
  AOI21_X1 U18707 ( .B1(n19539), .B2(n19674), .A(n15619), .ZN(n15620) );
  OAI21_X1 U18708 ( .B1(n19525), .B2(n15621), .A(n15620), .ZN(P2_U3128) );
  NAND3_X1 U18709 ( .A1(n10670), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19605) );
  NOR2_X1 U18710 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19605), .ZN(
        n19594) );
  NOR2_X1 U18711 ( .A1(n15623), .A2(n15622), .ZN(n19354) );
  NAND2_X1 U18712 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19354), .ZN(
        n15629) );
  INV_X1 U18713 ( .A(n19610), .ZN(n15624) );
  NAND2_X1 U18714 ( .A1(n15624), .A2(n19547), .ZN(n19563) );
  INV_X1 U18715 ( .A(n19609), .ZN(n19604) );
  OAI21_X1 U18716 ( .B1(n19596), .B2(n19623), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n15625) );
  NAND2_X1 U18717 ( .A1(n15629), .A2(n15625), .ZN(n15626) );
  OAI21_X1 U18718 ( .B1(n19594), .B2(n19385), .A(n15626), .ZN(n15627) );
  NOR2_X1 U18719 ( .A1(n19436), .A2(n15627), .ZN(n15628) );
  NAND2_X1 U18720 ( .A1(n15628), .A2(n15631), .ZN(n19597) );
  INV_X1 U18721 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15637) );
  OAI21_X1 U18722 ( .B1(n15629), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n10692), 
        .ZN(n15630) );
  AND2_X1 U18723 ( .A1(n15631), .A2(n15630), .ZN(n19595) );
  INV_X1 U18724 ( .A(n19594), .ZN(n15633) );
  AOI22_X1 U18725 ( .A1(n19623), .A2(n19682), .B1(n19596), .B2(n19632), .ZN(
        n15632) );
  OAI21_X1 U18726 ( .B1(n15634), .B2(n15633), .A(n15632), .ZN(n15635) );
  AOI21_X1 U18727 ( .B1(n19595), .B2(n19674), .A(n15635), .ZN(n15636) );
  OAI21_X1 U18728 ( .B1(n19587), .B2(n15637), .A(n15636), .ZN(P2_U3144) );
  INV_X1 U18729 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n17110) );
  INV_X1 U18730 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n16779) );
  NAND3_X1 U18731 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17221) );
  NOR3_X1 U18732 ( .A1(n16779), .A2(n16801), .A3(n17221), .ZN(n17142) );
  INV_X1 U18733 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16707) );
  INV_X1 U18734 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17143) );
  INV_X1 U18735 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n17204) );
  NAND2_X1 U18736 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .ZN(n17208) );
  NOR4_X1 U18737 ( .A1(n16707), .A2(n17143), .A3(n17204), .A4(n17208), .ZN(
        n15638) );
  NAND4_X1 U18738 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .A3(n17142), .A4(n15638), .ZN(n16842) );
  NOR2_X1 U18739 ( .A1(n17110), .A2(n16842), .ZN(n15653) );
  NOR3_X1 U18740 ( .A1(n15641), .A2(n17330), .A3(n15640), .ZN(n15642) );
  OAI21_X1 U18741 ( .B1(n15653), .B2(n17330), .A(n17235), .ZN(n17108) );
  NAND2_X1 U18742 ( .A1(n18245), .A2(n17235), .ZN(n17240) );
  NOR2_X1 U18743 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(n17240), .ZN(n17109) );
  AOI22_X1 U18744 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n15652) );
  AOI22_X1 U18745 ( .A1(n12834), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15651) );
  INV_X1 U18746 ( .A(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n20825) );
  AOI22_X1 U18747 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n16869), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15643) );
  OAI21_X1 U18748 ( .B1(n9767), .B2(n20825), .A(n15643), .ZN(n15649) );
  AOI22_X1 U18749 ( .A1(n12832), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n16876), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15647) );
  AOI22_X1 U18750 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15646) );
  AOI22_X1 U18751 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15645) );
  AOI22_X1 U18752 ( .A1(n17084), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15644) );
  NAND4_X1 U18753 ( .A1(n15647), .A2(n15646), .A3(n15645), .A4(n15644), .ZN(
        n15648) );
  AOI211_X1 U18754 ( .C1(n9753), .C2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        n15649), .B(n15648), .ZN(n15650) );
  NAND3_X1 U18755 ( .A1(n15652), .A2(n15651), .A3(n15650), .ZN(n17335) );
  NOR2_X2 U18756 ( .A1(n17237), .A2(n18245), .ZN(n17238) );
  AOI222_X1 U18757 ( .A1(n17108), .A2(P3_EBX_REG_13__SCAN_IN), .B1(n17109), 
        .B2(n15653), .C1(n17335), .C2(n17238), .ZN(n15654) );
  INV_X1 U18758 ( .A(n15654), .ZN(P3_U2690) );
  NAND2_X1 U18759 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18427) );
  AOI221_X1 U18760 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18427), .C1(n15656), 
        .C2(n18427), .A(n15655), .ZN(n18205) );
  NOR2_X1 U18761 ( .A1(n15657), .A2(n18659), .ZN(n15658) );
  OAI21_X1 U18762 ( .B1(n15658), .B2(n18209), .A(n18206), .ZN(n18203) );
  AOI22_X1 U18763 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18205), .B1(
        n18203), .B2(n18663), .ZN(P3_U2865) );
  NAND2_X1 U18764 ( .A1(n15660), .A2(n15659), .ZN(n18680) );
  INV_X1 U18765 ( .A(n15661), .ZN(n17446) );
  NAND2_X1 U18766 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18854) );
  NAND2_X1 U18767 ( .A1(n18682), .A2(n18854), .ZN(n15672) );
  NOR2_X1 U18768 ( .A1(n15663), .A2(n15662), .ZN(n18700) );
  INV_X1 U18769 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n20922) );
  NAND2_X2 U18770 ( .A1(n18842), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18796) );
  INV_X1 U18771 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18737) );
  NAND2_X1 U18772 ( .A1(n18728), .A2(n18737), .ZN(n16436) );
  NAND3_X1 U18773 ( .A1(n20922), .A2(n18796), .A3(n16436), .ZN(n18851) );
  INV_X1 U18774 ( .A(n18851), .ZN(n15680) );
  OAI21_X1 U18775 ( .B1(n15664), .B2(n18700), .A(n15680), .ZN(n17397) );
  NOR3_X1 U18776 ( .A1(n15667), .A2(n15666), .A3(n15665), .ZN(n15668) );
  OAI211_X1 U18777 ( .C1(n18229), .C2(n18655), .A(n15669), .B(n15668), .ZN(
        n15671) );
  AOI21_X1 U18778 ( .B1(n16430), .B2(n15671), .A(n15670), .ZN(n15686) );
  OAI21_X1 U18779 ( .B1(n15672), .B2(n17397), .A(n15686), .ZN(n15673) );
  AOI211_X1 U18780 ( .C1(n18683), .C2(n15674), .A(n15768), .B(n15673), .ZN(
        n18691) );
  INV_X1 U18781 ( .A(n18691), .ZN(n18677) );
  NOR2_X1 U18782 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18808), .ZN(n18212) );
  INV_X1 U18783 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18201) );
  NOR2_X1 U18784 ( .A1(n18201), .A2(n18806), .ZN(n15675) );
  AOI21_X1 U18785 ( .B1(n15676), .B2(n16785), .A(n18680), .ZN(n18690) );
  NAND3_X1 U18786 ( .A1(n18830), .A2(n18866), .A3(n18690), .ZN(n15677) );
  OAI21_X1 U18787 ( .B1(n18830), .B2(n16785), .A(n15677), .ZN(P3_U3284) );
  NOR4_X1 U18788 ( .A1(n18217), .A2(n18238), .A3(n18688), .A4(n15678), .ZN(
        n15683) );
  INV_X1 U18789 ( .A(n18682), .ZN(n15681) );
  OAI21_X1 U18790 ( .B1(n15680), .B2(n15679), .A(n18854), .ZN(n16438) );
  NOR3_X1 U18791 ( .A1(n15684), .A2(n15681), .A3(n16438), .ZN(n15682) );
  AOI211_X1 U18792 ( .C1(n18683), .C2(n15684), .A(n15683), .B(n15682), .ZN(
        n15685) );
  AOI21_X2 U18793 ( .B1(n15686), .B2(n15685), .A(n18708), .ZN(n18191) );
  NOR2_X1 U18794 ( .A1(n18185), .A2(n18072), .ZN(n18113) );
  NOR2_X1 U18795 ( .A1(n17657), .A2(n17994), .ZN(n16347) );
  AOI21_X1 U18796 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18144) );
  INV_X1 U18797 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18131) );
  NAND3_X1 U18798 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18118) );
  NOR3_X1 U18799 ( .A1(n18106), .A2(n18131), .A3(n18118), .ZN(n18102) );
  NAND2_X1 U18800 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18102), .ZN(
        n17993) );
  NOR2_X1 U18801 ( .A1(n18144), .A2(n17993), .ZN(n18005) );
  NAND2_X1 U18802 ( .A1(n16347), .A2(n18005), .ZN(n17941) );
  OAI21_X1 U18803 ( .B1(n18094), .B2(n21021), .A(n18656), .ZN(n18171) );
  NAND2_X1 U18804 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18103) );
  NOR2_X1 U18805 ( .A1(n18103), .A2(n17993), .ZN(n15689) );
  NAND3_X1 U18806 ( .A1(n18171), .A2(n15689), .A3(n16347), .ZN(n15687) );
  OAI21_X1 U18807 ( .B1(n18685), .B2(n17941), .A(n15687), .ZN(n16346) );
  NAND2_X1 U18808 ( .A1(n17580), .A2(n16346), .ZN(n17906) );
  NAND2_X1 U18809 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17909) );
  NOR2_X1 U18810 ( .A1(n17885), .A2(n17909), .ZN(n16303) );
  NAND2_X1 U18811 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n16303), .ZN(
        n17518) );
  OR2_X1 U18812 ( .A1(n18185), .A2(n17518), .ZN(n16348) );
  NOR3_X1 U18813 ( .A1(n12905), .A2(n17906), .A3(n16348), .ZN(n16331) );
  NAND2_X1 U18814 ( .A1(n18069), .A2(n18191), .ZN(n18198) );
  NOR2_X1 U18815 ( .A1(n16340), .A2(n18198), .ZN(n15688) );
  AOI211_X1 U18816 ( .C1(n18113), .C2(n16341), .A(n16331), .B(n15688), .ZN(
        n15741) );
  INV_X1 U18817 ( .A(n15689), .ZN(n18006) );
  NOR2_X1 U18818 ( .A1(n17994), .A2(n18006), .ZN(n17986) );
  NOR2_X1 U18819 ( .A1(n17657), .A2(n17601), .ZN(n17944) );
  NAND2_X1 U18820 ( .A1(n17986), .A2(n17944), .ZN(n17882) );
  NOR2_X1 U18821 ( .A1(n17954), .A2(n17882), .ZN(n15691) );
  NAND2_X1 U18822 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15691), .ZN(
        n17883) );
  INV_X1 U18823 ( .A(n16303), .ZN(n15690) );
  INV_X1 U18824 ( .A(n17941), .ZN(n17987) );
  NAND2_X1 U18825 ( .A1(n17580), .A2(n17987), .ZN(n17927) );
  OAI21_X1 U18826 ( .B1(n15690), .B2(n17927), .A(n18145), .ZN(n17889) );
  OAI221_X1 U18827 ( .B1(n18656), .B2(n16303), .C1(n18656), .C2(n15691), .A(
        n17889), .ZN(n15692) );
  AOI221_X1 U18828 ( .B1(n17518), .B2(n18654), .C1(n17883), .C2(n18654), .A(
        n15692), .ZN(n15736) );
  OAI211_X1 U18829 ( .C1(n18052), .C2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n18191), .B(n15736), .ZN(n16339) );
  NAND2_X1 U18830 ( .A1(n18107), .A2(n18191), .ZN(n18180) );
  INV_X1 U18831 ( .A(n15693), .ZN(n16300) );
  AOI22_X1 U18832 ( .A1(n18113), .A2(n16300), .B1(n18184), .B2(n16301), .ZN(
        n15744) );
  OAI21_X1 U18833 ( .B1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n18180), .A(
        n15744), .ZN(n15694) );
  AOI21_X1 U18834 ( .B1(n18193), .B2(n16339), .A(n15694), .ZN(n15697) );
  OAI22_X1 U18835 ( .A1(n16338), .A2(n10129), .B1(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n12900), .ZN(n15695) );
  XOR2_X1 U18836 ( .A(n16317), .B(n15695), .Z(n16320) );
  AOI22_X1 U18837 ( .A1(n9726), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n9717), .B2(
        n16320), .ZN(n15696) );
  OAI221_X1 U18838 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15741), 
        .C1(n16317), .C2(n15697), .A(n15696), .ZN(P3_U2833) );
  INV_X1 U18839 ( .A(n15698), .ZN(n15710) );
  INV_X1 U18840 ( .A(n15699), .ZN(n15701) );
  NAND2_X1 U18841 ( .A1(n15701), .A2(n15700), .ZN(n15706) );
  INV_X1 U18842 ( .A(n15702), .ZN(n15703) );
  AOI21_X1 U18843 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n15704), .A(
        n15703), .ZN(n15705) );
  OAI211_X1 U18844 ( .C1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n15706), .A(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n15705), .ZN(n15708) );
  NAND2_X1 U18845 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n15706), .ZN(
        n15707) );
  NAND2_X1 U18846 ( .A1(n15708), .A2(n15707), .ZN(n15709) );
  AOI222_X1 U18847 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n15710), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15709), .C1(n15710), 
        .C2(n15709), .ZN(n15711) );
  AOI222_X1 U18848 ( .A1(n20486), .A2(n15712), .B1(n20486), .B2(n15711), .C1(
        n15712), .C2(n15711), .ZN(n15719) );
  INV_X1 U18849 ( .A(n15713), .ZN(n15714) );
  NOR2_X1 U18850 ( .A1(n15715), .A2(n15714), .ZN(n15718) );
  OAI21_X1 U18851 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15716), .ZN(n15717) );
  OAI211_X1 U18852 ( .C1(n15719), .C2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n15718), .B(n15717), .ZN(n15720) );
  NOR3_X1 U18853 ( .A1(n15722), .A2(n15721), .A3(n15720), .ZN(n15735) );
  INV_X1 U18854 ( .A(n15735), .ZN(n15728) );
  NOR3_X1 U18855 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20640), .A3(n20718), 
        .ZN(n15726) );
  NAND3_X1 U18856 ( .A1(n13153), .A2(n20120), .A3(n15723), .ZN(n15725) );
  OAI22_X1 U18857 ( .A1(n15727), .A2(n15726), .B1(n15725), .B2(n15724), .ZN(
        n16062) );
  AOI221_X1 U18858 ( .B1(n20639), .B2(n14146), .C1(n15728), .C2(n14146), .A(
        n16062), .ZN(n15730) );
  NOR2_X1 U18859 ( .A1(n15730), .A2(n20639), .ZN(n16065) );
  OAI211_X1 U18860 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n20718), .A(n16065), 
        .B(n15729), .ZN(n16063) );
  AOI21_X1 U18861 ( .B1(n20722), .B2(n15731), .A(n15730), .ZN(n15732) );
  OAI22_X1 U18862 ( .A1(n15733), .A2(n16063), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n15732), .ZN(n15734) );
  OAI21_X1 U18863 ( .B1(n15735), .B2(n19884), .A(n15734), .ZN(P1_U3161) );
  INV_X1 U18864 ( .A(n18180), .ZN(n15738) );
  OAI21_X1 U18865 ( .B1(n15736), .B2(n18185), .A(n18165), .ZN(n15737) );
  AOI21_X1 U18866 ( .B1(n15738), .B2(n16304), .A(n15737), .ZN(n16328) );
  OAI21_X1 U18867 ( .B1(n15740), .B2(n21009), .A(n15739), .ZN(n16310) );
  INV_X1 U18868 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18795) );
  NOR2_X1 U18869 ( .A1(n18193), .A2(n18795), .ZN(n16305) );
  NOR3_X1 U18870 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n15741), .A3(
        n16317), .ZN(n15742) );
  AOI211_X1 U18871 ( .C1(n9717), .C2(n16310), .A(n16305), .B(n15742), .ZN(
        n15743) );
  OAI221_X1 U18872 ( .B1(n21009), .B2(n16328), .C1(n21009), .C2(n15744), .A(
        n15743), .ZN(P3_U2832) );
  INV_X1 U18873 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20658) );
  INV_X1 U18874 ( .A(HOLD), .ZN(n19750) );
  NOR2_X1 U18875 ( .A1(n20658), .A2(n19750), .ZN(n20646) );
  AOI22_X1 U18876 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n15747) );
  NAND2_X1 U18877 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n15745), .ZN(n20644) );
  OAI211_X1 U18878 ( .C1(n20646), .C2(n15747), .A(n15746), .B(n20644), .ZN(
        P1_U3195) );
  INV_X1 U18879 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16425) );
  NOR2_X1 U18880 ( .A1(n20017), .A2(n16425), .ZN(P1_U2905) );
  NOR2_X1 U18881 ( .A1(n15748), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15751) );
  NOR2_X1 U18882 ( .A1(n14508), .A2(n15749), .ZN(n15750) );
  MUX2_X1 U18883 ( .A(n15751), .B(n15750), .S(n14160), .Z(n15752) );
  XOR2_X1 U18884 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n15752), .Z(
        n15924) );
  AOI22_X1 U18885 ( .A1(n15924), .A2(n20082), .B1(n20085), .B2(n15823), .ZN(
        n15760) );
  NAND3_X1 U18886 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15754), .A3(
        n15753), .ZN(n15759) );
  NAND2_X1 U18887 ( .A1(n16053), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15925) );
  AOI21_X1 U18888 ( .B1(n15755), .B2(n16018), .A(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15757) );
  OAI21_X1 U18889 ( .B1(n15757), .B2(n15756), .A(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15758) );
  NAND4_X1 U18890 ( .A1(n15760), .A2(n15759), .A3(n15925), .A4(n15758), .ZN(
        P1_U3011) );
  NOR2_X1 U18891 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n15761) );
  NOR3_X1 U18892 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n18874), .A3(n19867), 
        .ZN(n16286) );
  NOR4_X1 U18893 ( .A1(n15762), .A2(n15761), .A3(n16286), .A4(n16298), .ZN(
        P2_U3178) );
  INV_X1 U18894 ( .A(n19853), .ZN(n15763) );
  AOI221_X1 U18895 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16298), .C1(n15763), .C2(
        n16298), .A(n19680), .ZN(n19849) );
  INV_X1 U18896 ( .A(n19849), .ZN(n19850) );
  NOR2_X1 U18897 ( .A1(n15764), .A2(n19850), .ZN(P2_U3047) );
  NOR2_X1 U18898 ( .A1(n15766), .A2(n15765), .ZN(n15767) );
  NOR2_X1 U18899 ( .A1(n17330), .A2(n17388), .ZN(n17364) );
  INV_X1 U18900 ( .A(n17364), .ZN(n17359) );
  INV_X1 U18901 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n20971) );
  NAND2_X1 U18902 ( .A1(n17330), .A2(n17242), .ZN(n17389) );
  NOR2_X2 U18903 ( .A1(n15769), .A2(n17388), .ZN(n17392) );
  AOI22_X1 U18904 ( .A1(n17393), .A2(BUF2_REG_0__SCAN_IN), .B1(n17392), .B2(
        n15770), .ZN(n15771) );
  OAI221_X1 U18905 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17359), .C1(n20971), 
        .C2(n17242), .A(n15771), .ZN(P3_U2735) );
  INV_X1 U18906 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n15776) );
  NOR2_X1 U18907 ( .A1(n19969), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n15772) );
  AOI22_X1 U18908 ( .A1(n15773), .A2(n15772), .B1(n19971), .B2(
        P1_EBX_REG_24__SCAN_IN), .ZN(n15775) );
  NAND2_X1 U18909 ( .A1(n19991), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15774) );
  OAI211_X1 U18910 ( .C1(n15785), .C2(n15776), .A(n15775), .B(n15774), .ZN(
        n15777) );
  INV_X1 U18911 ( .A(n15777), .ZN(n15781) );
  AOI22_X1 U18912 ( .A1(n15779), .A2(n19932), .B1(n15778), .B2(n19959), .ZN(
        n15780) );
  OAI211_X1 U18913 ( .C1(n15782), .C2(n19965), .A(n15781), .B(n15780), .ZN(
        P1_U2816) );
  INV_X1 U18914 ( .A(n15783), .ZN(n15796) );
  NAND2_X1 U18915 ( .A1(n19982), .A2(n15796), .ZN(n15819) );
  OAI21_X1 U18916 ( .B1(n15784), .B2(n15819), .A(n20686), .ZN(n15787) );
  INV_X1 U18917 ( .A(n15785), .ZN(n15786) );
  AOI22_X1 U18918 ( .A1(n15787), .A2(n15786), .B1(n19971), .B2(
        P1_EBX_REG_23__SCAN_IN), .ZN(n15794) );
  INV_X1 U18919 ( .A(n15788), .ZN(n15789) );
  OAI22_X1 U18920 ( .A1(n15790), .A2(n15894), .B1(n15789), .B2(n19987), .ZN(
        n15791) );
  AOI21_X1 U18921 ( .B1(n15792), .B2(n19993), .A(n15791), .ZN(n15793) );
  OAI211_X1 U18922 ( .C1(n15795), .C2(n19956), .A(n15794), .B(n15793), .ZN(
        P1_U2817) );
  NAND2_X1 U18923 ( .A1(n15796), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15808) );
  INV_X1 U18924 ( .A(n19929), .ZN(n15797) );
  OAI21_X1 U18925 ( .B1(n19967), .B2(n15808), .A(n15797), .ZN(n15818) );
  OAI21_X1 U18926 ( .B1(P1_REIP_REG_21__SCAN_IN), .B2(n19969), .A(n15818), 
        .ZN(n15802) );
  NAND2_X1 U18927 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n15798) );
  NOR3_X1 U18928 ( .A1(P1_REIP_REG_22__SCAN_IN), .A2(n15798), .A3(n15819), 
        .ZN(n15801) );
  OAI22_X1 U18929 ( .A1(n19956), .A2(n15799), .B1(n19986), .B2(n15918), .ZN(
        n15800) );
  AOI211_X1 U18930 ( .C1(P1_REIP_REG_22__SCAN_IN), .C2(n15802), .A(n15801), 
        .B(n15800), .ZN(n15806) );
  INV_X1 U18931 ( .A(n15803), .ZN(n15914) );
  OAI22_X1 U18932 ( .A1(n15915), .A2(n15894), .B1(n15914), .B2(n19987), .ZN(
        n15804) );
  INV_X1 U18933 ( .A(n15804), .ZN(n15805) );
  OAI211_X1 U18934 ( .C1(n15807), .C2(n19965), .A(n15806), .B(n15805), .ZN(
        P1_U2818) );
  NOR3_X1 U18935 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n19969), .A3(n15808), 
        .ZN(n15811) );
  OAI22_X1 U18936 ( .A1(n15818), .A2(n20683), .B1(n15809), .B2(n19986), .ZN(
        n15810) );
  AOI211_X1 U18937 ( .C1(n19991), .C2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n15811), .B(n15810), .ZN(n15816) );
  INV_X1 U18938 ( .A(n15812), .ZN(n15813) );
  AOI22_X1 U18939 ( .A1(n15814), .A2(n19932), .B1(n15813), .B2(n19993), .ZN(
        n15815) );
  OAI211_X1 U18940 ( .C1(n15817), .C2(n19987), .A(n15816), .B(n15815), .ZN(
        P1_U2819) );
  INV_X1 U18941 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n21011) );
  INV_X1 U18942 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n15820) );
  AOI21_X1 U18943 ( .B1(n15820), .B2(n15819), .A(n15818), .ZN(n15821) );
  AOI21_X1 U18944 ( .B1(n19971), .B2(P1_EBX_REG_20__SCAN_IN), .A(n15821), .ZN(
        n15825) );
  OAI22_X1 U18945 ( .A1(n15922), .A2(n15894), .B1(n15921), .B2(n19965), .ZN(
        n15822) );
  AOI21_X1 U18946 ( .B1(n19959), .B2(n15823), .A(n15822), .ZN(n15824) );
  OAI211_X1 U18947 ( .C1(n21011), .C2(n19956), .A(n15825), .B(n15824), .ZN(
        P1_U2820) );
  INV_X1 U18948 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n15827) );
  NAND3_X1 U18949 ( .A1(n19982), .A2(n15826), .A3(n15829), .ZN(n15841) );
  AOI221_X1 U18950 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(P1_REIP_REG_18__SCAN_IN), .C1(n14517), .C2(n15827), .A(n15841), .ZN(n15833) );
  OAI21_X1 U18951 ( .B1(n15829), .B2(n19969), .A(n15828), .ZN(n15852) );
  AOI22_X1 U18952 ( .A1(n15852), .A2(P1_REIP_REG_19__SCAN_IN), .B1(
        P1_EBX_REG_19__SCAN_IN), .B2(n19971), .ZN(n15830) );
  OAI211_X1 U18953 ( .C1(n19956), .C2(n15831), .A(n15830), .B(n19953), .ZN(
        n15832) );
  NOR2_X1 U18954 ( .A1(n15833), .A2(n15832), .ZN(n15834) );
  OAI21_X1 U18955 ( .B1(n15835), .B2(n15894), .A(n15834), .ZN(n15836) );
  AOI21_X1 U18956 ( .B1(n15837), .B2(n19993), .A(n15836), .ZN(n15838) );
  OAI21_X1 U18957 ( .B1(n19987), .B2(n15839), .A(n15838), .ZN(P1_U2821) );
  AOI22_X1 U18958 ( .A1(n15852), .A2(P1_REIP_REG_18__SCAN_IN), .B1(n19971), 
        .B2(P1_EBX_REG_18__SCAN_IN), .ZN(n15840) );
  OAI21_X1 U18959 ( .B1(P1_REIP_REG_18__SCAN_IN), .B2(n15841), .A(n15840), 
        .ZN(n15842) );
  AOI211_X1 U18960 ( .C1(n19991), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n19925), .B(n15842), .ZN(n15847) );
  OAI21_X1 U18961 ( .B1(n14347), .B2(n15844), .A(n15843), .ZN(n15845) );
  INV_X1 U18962 ( .A(n15845), .ZN(n15988) );
  AOI22_X1 U18963 ( .A1(n15930), .A2(n19932), .B1(n19959), .B2(n15988), .ZN(
        n15846) );
  OAI211_X1 U18964 ( .C1(n15933), .C2(n19965), .A(n15847), .B(n15846), .ZN(
        P1_U2822) );
  OAI22_X1 U18965 ( .A1(n19956), .A2(n15849), .B1(n15848), .B2(n19986), .ZN(
        n15850) );
  AOI211_X1 U18966 ( .C1(n19993), .C2(n15851), .A(n19925), .B(n15850), .ZN(
        n15856) );
  NAND3_X1 U18967 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_14__SCAN_IN), 
        .A3(n15879), .ZN(n15876) );
  OAI21_X1 U18968 ( .B1(n15858), .B2(n15876), .A(n20676), .ZN(n15853) );
  AOI22_X1 U18969 ( .A1(n15854), .A2(n19932), .B1(n15853), .B2(n15852), .ZN(
        n15855) );
  OAI211_X1 U18970 ( .C1(n19987), .C2(n15857), .A(n15856), .B(n15855), .ZN(
        P1_U2823) );
  OAI21_X1 U18971 ( .B1(P1_REIP_REG_16__SCAN_IN), .B2(P1_REIP_REG_15__SCAN_IN), 
        .A(n15858), .ZN(n15867) );
  INV_X1 U18972 ( .A(n15859), .ZN(n15860) );
  OAI21_X1 U18973 ( .B1(n15860), .B2(n19929), .A(n15913), .ZN(n15878) );
  AOI22_X1 U18974 ( .A1(n19959), .A2(n15996), .B1(P1_REIP_REG_16__SCAN_IN), 
        .B2(n15878), .ZN(n15866) );
  INV_X1 U18975 ( .A(n15942), .ZN(n15861) );
  AOI22_X1 U18976 ( .A1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n19991), .B1(
        n19993), .B2(n15861), .ZN(n15862) );
  OAI211_X1 U18977 ( .C1(n19986), .C2(n15863), .A(n15862), .B(n19953), .ZN(
        n15864) );
  AOI21_X1 U18978 ( .B1(n15939), .B2(n19932), .A(n15864), .ZN(n15865) );
  OAI211_X1 U18979 ( .C1(n15876), .C2(n15867), .A(n15866), .B(n15865), .ZN(
        P1_U2824) );
  AOI22_X1 U18980 ( .A1(n15868), .A2(n19993), .B1(P1_REIP_REG_15__SCAN_IN), 
        .B2(n15878), .ZN(n15875) );
  AOI21_X1 U18981 ( .B1(n19971), .B2(P1_EBX_REG_15__SCAN_IN), .A(n19925), .ZN(
        n15869) );
  OAI21_X1 U18982 ( .B1(n15870), .B2(n19956), .A(n15869), .ZN(n15873) );
  NOR2_X1 U18983 ( .A1(n15871), .A2(n15894), .ZN(n15872) );
  AOI211_X1 U18984 ( .C1(n19959), .C2(n16002), .A(n15873), .B(n15872), .ZN(
        n15874) );
  OAI211_X1 U18985 ( .C1(P1_REIP_REG_15__SCAN_IN), .C2(n15876), .A(n15875), 
        .B(n15874), .ZN(P1_U2825) );
  AOI22_X1 U18986 ( .A1(n19991), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n19971), .B2(P1_EBX_REG_14__SCAN_IN), .ZN(n15883) );
  AOI21_X1 U18987 ( .B1(n16011), .B2(n19959), .A(n19925), .ZN(n15882) );
  INV_X1 U18988 ( .A(n15877), .ZN(n15952) );
  AOI22_X1 U18989 ( .A1(n15952), .A2(n19932), .B1(n19993), .B2(n15951), .ZN(
        n15881) );
  OAI221_X1 U18990 ( .B1(P1_REIP_REG_14__SCAN_IN), .B2(P1_REIP_REG_13__SCAN_IN), .C1(P1_REIP_REG_14__SCAN_IN), .C2(n15879), .A(n15878), .ZN(n15880) );
  NAND4_X1 U18991 ( .A1(n15883), .A2(n15882), .A3(n15881), .A4(n15880), .ZN(
        P1_U2826) );
  OAI22_X1 U18992 ( .A1(n19956), .A2(n15885), .B1(n15884), .B2(n19986), .ZN(
        n15886) );
  AOI211_X1 U18993 ( .C1(n16015), .C2(n19959), .A(n19925), .B(n15886), .ZN(
        n15892) );
  NAND2_X1 U18994 ( .A1(n15888), .A2(n15887), .ZN(n15889) );
  AOI22_X1 U18995 ( .A1(n15959), .A2(n19993), .B1(n15890), .B2(n15889), .ZN(
        n15891) );
  OAI211_X1 U18996 ( .C1(n15894), .C2(n15893), .A(n15892), .B(n15891), .ZN(
        P1_U2828) );
  NAND2_X1 U18997 ( .A1(n19971), .A2(P1_EBX_REG_11__SCAN_IN), .ZN(n15895) );
  OAI211_X1 U18998 ( .C1(n15896), .C2(n19987), .A(n19953), .B(n15895), .ZN(
        n15898) );
  NOR2_X1 U18999 ( .A1(n15913), .A2(n20840), .ZN(n15897) );
  AOI211_X1 U19000 ( .C1(n19991), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n15898), .B(n15897), .ZN(n15901) );
  AOI22_X1 U19001 ( .A1(n15963), .A2(n19932), .B1(n15899), .B2(n20840), .ZN(
        n15900) );
  OAI211_X1 U19002 ( .C1(n15967), .C2(n19965), .A(n15901), .B(n15900), .ZN(
        P1_U2829) );
  OAI22_X1 U19003 ( .A1(n16027), .A2(n19987), .B1(n19986), .B2(n15902), .ZN(
        n15903) );
  INV_X1 U19004 ( .A(n15903), .ZN(n15904) );
  OAI21_X1 U19005 ( .B1(P1_REIP_REG_10__SCAN_IN), .B2(n15905), .A(n15904), 
        .ZN(n15906) );
  AOI211_X1 U19006 ( .C1(n19991), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n19925), .B(n15906), .ZN(n15912) );
  INV_X1 U19007 ( .A(n15907), .ZN(n15910) );
  INV_X1 U19008 ( .A(n15908), .ZN(n15909) );
  AOI22_X1 U19009 ( .A1(n15910), .A2(n19932), .B1(n15909), .B2(n19993), .ZN(
        n15911) );
  OAI211_X1 U19010 ( .C1(n15913), .C2(n20668), .A(n15912), .B(n15911), .ZN(
        P1_U2830) );
  OAI22_X1 U19011 ( .A1(n15915), .A2(n14359), .B1(n15914), .B2(n20002), .ZN(
        n15916) );
  INV_X1 U19012 ( .A(n15916), .ZN(n15917) );
  OAI21_X1 U19013 ( .B1(n14350), .B2(n15918), .A(n15917), .ZN(P1_U2850) );
  AOI22_X1 U19014 ( .A1(n15930), .A2(n20004), .B1(n11892), .B2(n15988), .ZN(
        n15919) );
  OAI21_X1 U19015 ( .B1(n14350), .B2(n15920), .A(n15919), .ZN(P1_U2854) );
  OAI22_X1 U19016 ( .A1(n15922), .A2(n20106), .B1(n15921), .B2(n15978), .ZN(
        n15923) );
  AOI21_X1 U19017 ( .B1(n20064), .B2(n15924), .A(n15923), .ZN(n15926) );
  OAI211_X1 U19018 ( .C1(n21011), .C2(n15984), .A(n15926), .B(n15925), .ZN(
        P1_U2979) );
  AOI22_X1 U19019 ( .A1(n20060), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B1(
        n16053), .B2(P1_REIP_REG_18__SCAN_IN), .ZN(n15932) );
  OAI21_X1 U19020 ( .B1(n15928), .B2(n15927), .A(n14508), .ZN(n15929) );
  INV_X1 U19021 ( .A(n15929), .ZN(n15989) );
  AOI22_X1 U19022 ( .A1(n15989), .A2(n20064), .B1(n15975), .B2(n15930), .ZN(
        n15931) );
  OAI211_X1 U19023 ( .C1(n15978), .C2(n15933), .A(n15932), .B(n15931), .ZN(
        P1_U2981) );
  AOI22_X1 U19024 ( .A1(n20060), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n16053), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15941) );
  OAI21_X1 U19025 ( .B1(n15936), .B2(n15935), .A(n15934), .ZN(n15938) );
  XNOR2_X1 U19026 ( .A(n15938), .B(n15937), .ZN(n15997) );
  AOI22_X1 U19027 ( .A1(n15997), .A2(n20064), .B1(n15975), .B2(n15939), .ZN(
        n15940) );
  OAI211_X1 U19028 ( .C1(n15978), .C2(n15942), .A(n15941), .B(n15940), .ZN(
        P1_U2983) );
  INV_X1 U19029 ( .A(n15943), .ZN(n15944) );
  NAND2_X1 U19030 ( .A1(n15945), .A2(n15944), .ZN(n15947) );
  OAI21_X1 U19031 ( .B1(n15948), .B2(n15947), .A(n15946), .ZN(n15950) );
  XNOR2_X1 U19032 ( .A(n14160), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15949) );
  XNOR2_X1 U19033 ( .A(n15950), .B(n15949), .ZN(n16014) );
  AOI22_X1 U19034 ( .A1(n20060), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n16053), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15954) );
  AOI22_X1 U19035 ( .A1(n15952), .A2(n15975), .B1(n15979), .B2(n15951), .ZN(
        n15953) );
  OAI211_X1 U19036 ( .C1(n16014), .C2(n15962), .A(n15954), .B(n15953), .ZN(
        P1_U2985) );
  AOI21_X1 U19037 ( .B1(n15957), .B2(n15956), .A(n15955), .ZN(n16026) );
  AOI22_X1 U19038 ( .A1(n20060), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n16053), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15961) );
  AOI22_X1 U19039 ( .A1(n15979), .A2(n15959), .B1(n15975), .B2(n15958), .ZN(
        n15960) );
  OAI211_X1 U19040 ( .C1(n16026), .C2(n15962), .A(n15961), .B(n15960), .ZN(
        P1_U2987) );
  AOI22_X1 U19041 ( .A1(n20060), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n16053), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15966) );
  AOI22_X1 U19042 ( .A1(n20064), .A2(n15964), .B1(n15975), .B2(n15963), .ZN(
        n15965) );
  OAI211_X1 U19043 ( .C1(n15978), .C2(n15967), .A(n15966), .B(n15965), .ZN(
        P1_U2988) );
  AOI22_X1 U19044 ( .A1(n20060), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n16053), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15970) );
  AOI22_X1 U19045 ( .A1(n15968), .A2(n20064), .B1(n15975), .B2(n19917), .ZN(
        n15969) );
  OAI211_X1 U19046 ( .C1(n15978), .C2(n19920), .A(n15970), .B(n15969), .ZN(
        P1_U2992) );
  AOI22_X1 U19047 ( .A1(n20060), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n16053), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15977) );
  NAND2_X1 U19048 ( .A1(n15973), .A2(n15972), .ZN(n15974) );
  XNOR2_X1 U19049 ( .A(n15971), .B(n15974), .ZN(n16056) );
  AOI22_X1 U19050 ( .A1(n16056), .A2(n20064), .B1(n15975), .B2(n20005), .ZN(
        n15976) );
  OAI211_X1 U19051 ( .C1(n15978), .C2(n19935), .A(n15977), .B(n15976), .ZN(
        P1_U2993) );
  INV_X1 U19052 ( .A(n19950), .ZN(n15980) );
  AOI222_X1 U19053 ( .A1(n15981), .A2(n20064), .B1(n15975), .B2(n19948), .C1(
        n15980), .C2(n15979), .ZN(n15983) );
  OAI211_X1 U19054 ( .C1(n20884), .C2(n15984), .A(n15983), .B(n15982), .ZN(
        P1_U2994) );
  NOR2_X1 U19055 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15985), .ZN(
        n15986) );
  AOI22_X1 U19056 ( .A1(n16053), .A2(P1_REIP_REG_18__SCAN_IN), .B1(n15987), 
        .B2(n15986), .ZN(n15991) );
  AOI22_X1 U19057 ( .A1(n15989), .A2(n20082), .B1(n20085), .B2(n15988), .ZN(
        n15990) );
  OAI211_X1 U19058 ( .C1(n15992), .C2(n14175), .A(n15991), .B(n15990), .ZN(
        P1_U3013) );
  OAI21_X1 U19059 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n15993), .ZN(n16000) );
  OAI21_X1 U19060 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15995), .A(
        n15994), .ZN(n16001) );
  AOI22_X1 U19061 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n16001), .B1(
        n16053), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15999) );
  AOI22_X1 U19062 ( .A1(n15997), .A2(n20082), .B1(n20085), .B2(n15996), .ZN(
        n15998) );
  OAI211_X1 U19063 ( .C1(n16006), .C2(n16000), .A(n15999), .B(n15998), .ZN(
        P1_U3015) );
  AOI22_X1 U19064 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n16001), .B1(
        n16053), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n16005) );
  AOI22_X1 U19065 ( .A1(n16003), .A2(n20082), .B1(n20085), .B2(n16002), .ZN(
        n16004) );
  OAI211_X1 U19066 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16006), .A(
        n16005), .B(n16004), .ZN(P1_U3016) );
  AOI22_X1 U19067 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n16007), .B1(
        n16053), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n16013) );
  INV_X1 U19068 ( .A(n16030), .ZN(n16055) );
  AND3_X1 U19069 ( .A1(n16009), .A2(n16008), .A3(n16055), .ZN(n16010) );
  AOI21_X1 U19070 ( .B1(n16011), .B2(n20070), .A(n16010), .ZN(n16012) );
  OAI211_X1 U19071 ( .C1(n16014), .C2(n16025), .A(n16013), .B(n16012), .ZN(
        P1_U3017) );
  AOI22_X1 U19072 ( .A1(n16015), .A2(n20070), .B1(n16053), .B2(
        P1_REIP_REG_12__SCAN_IN), .ZN(n16024) );
  OAI21_X1 U19073 ( .B1(n16018), .B2(n16017), .A(n16016), .ZN(n16021) );
  OAI21_X1 U19074 ( .B1(n16019), .B2(n16030), .A(n16022), .ZN(n16020) );
  OAI21_X1 U19075 ( .B1(n16022), .B2(n16021), .A(n16020), .ZN(n16023) );
  OAI211_X1 U19076 ( .C1(n16026), .C2(n16025), .A(n16024), .B(n16023), .ZN(
        P1_U3019) );
  INV_X1 U19077 ( .A(n16027), .ZN(n16029) );
  AOI21_X1 U19078 ( .B1(n20085), .B2(n16029), .A(n16028), .ZN(n16036) );
  AOI211_X1 U19079 ( .C1(n16038), .C2(n14158), .A(n16031), .B(n16030), .ZN(
        n16033) );
  NAND2_X1 U19080 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16032) );
  AOI22_X1 U19081 ( .A1(n16034), .A2(n20082), .B1(n16033), .B2(n16032), .ZN(
        n16035) );
  OAI211_X1 U19082 ( .C1(n16038), .C2(n16037), .A(n16036), .B(n16035), .ZN(
        P1_U3021) );
  AOI21_X1 U19083 ( .B1(n20085), .B2(n16040), .A(n16039), .ZN(n16048) );
  AOI22_X1 U19084 ( .A1(n16042), .A2(n20082), .B1(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n16041), .ZN(n16047) );
  OAI221_X1 U19085 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(n16045), .C2(n16044), .A(
        n16043), .ZN(n16046) );
  NAND3_X1 U19086 ( .A1(n16048), .A2(n16047), .A3(n16046), .ZN(P1_U3023) );
  OR2_X1 U19087 ( .A1(n16050), .A2(n16049), .ZN(n16051) );
  NAND2_X1 U19088 ( .A1(n16052), .A2(n16051), .ZN(n20001) );
  INV_X1 U19089 ( .A(n20001), .ZN(n16054) );
  AOI22_X1 U19090 ( .A1(n20070), .A2(n16054), .B1(n16053), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n16058) );
  AOI22_X1 U19091 ( .A1(n16056), .A2(n20082), .B1(n16055), .B2(n16059), .ZN(
        n16057) );
  OAI211_X1 U19092 ( .C1(n16060), .C2(n16059), .A(n16058), .B(n16057), .ZN(
        P1_U3025) );
  OAI221_X1 U19093 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(
        P1_STATEBS16_REG_SCAN_IN), .C1(n20639), .C2(n20718), .A(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n20641) );
  NAND2_X1 U19094 ( .A1(n20641), .A2(n16064), .ZN(n16061) );
  AOI22_X1 U19095 ( .A1(n14146), .A2(n16063), .B1(n16062), .B2(n16061), .ZN(
        P1_U3162) );
  OAI22_X1 U19096 ( .A1(n16065), .A2(n20492), .B1(n20639), .B2(n16064), .ZN(
        P1_U3466) );
  AOI222_X1 U19097 ( .A1(n16066), .A2(n19035), .B1(P2_REIP_REG_31__SCAN_IN), 
        .B2(n19028), .C1(P2_EBX_REG_31__SCAN_IN), .C2(n18957), .ZN(n16067) );
  INV_X1 U19098 ( .A(n16067), .ZN(n16068) );
  AOI21_X1 U19099 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19003), .A(
        n16068), .ZN(n16071) );
  INV_X1 U19100 ( .A(n16069), .ZN(n19048) );
  AOI22_X1 U19101 ( .A1(n12774), .A2(n10916), .B1(n19029), .B2(n19048), .ZN(
        n16070) );
  OAI211_X1 U19102 ( .C1(n16073), .C2(n16072), .A(n16071), .B(n16070), .ZN(
        P2_U2824) );
  AOI22_X1 U19103 ( .A1(P2_EBX_REG_29__SCAN_IN), .A2(n18957), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n19028), .ZN(n16083) );
  AOI22_X1 U19104 ( .A1(n16074), .A2(n19035), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19003), .ZN(n16082) );
  AOI22_X1 U19105 ( .A1(n16076), .A2(n10916), .B1(n19029), .B2(n16075), .ZN(
        n16081) );
  OAI211_X1 U19106 ( .C1(n16079), .C2(n16078), .A(n18915), .B(n16077), .ZN(
        n16080) );
  NAND4_X1 U19107 ( .A1(n16083), .A2(n16082), .A3(n16081), .A4(n16080), .ZN(
        P2_U2826) );
  AOI22_X1 U19108 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(n18957), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19028), .ZN(n16093) );
  AOI22_X1 U19109 ( .A1(n16084), .A2(n19035), .B1(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n19003), .ZN(n16092) );
  AOI22_X1 U19110 ( .A1(n16086), .A2(n10916), .B1(n16085), .B2(n19029), .ZN(
        n16091) );
  OAI211_X1 U19111 ( .C1(n16089), .C2(n16088), .A(n18915), .B(n16087), .ZN(
        n16090) );
  NAND4_X1 U19112 ( .A1(n16093), .A2(n16092), .A3(n16091), .A4(n16090), .ZN(
        P2_U2827) );
  AOI22_X1 U19113 ( .A1(P2_EBX_REG_27__SCAN_IN), .A2(n18957), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n19028), .ZN(n16105) );
  INV_X1 U19114 ( .A(n16094), .ZN(n16095) );
  AOI22_X1 U19115 ( .A1(n16095), .A2(n19035), .B1(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n19003), .ZN(n16104) );
  INV_X1 U19116 ( .A(n16096), .ZN(n16098) );
  AOI22_X1 U19117 ( .A1(n16098), .A2(n10916), .B1(n16097), .B2(n19029), .ZN(
        n16103) );
  OAI211_X1 U19118 ( .C1(n16101), .C2(n16100), .A(n18915), .B(n16099), .ZN(
        n16102) );
  NAND4_X1 U19119 ( .A1(n16105), .A2(n16104), .A3(n16103), .A4(n16102), .ZN(
        P2_U2828) );
  AOI22_X1 U19120 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n18957), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n19028), .ZN(n16117) );
  OAI22_X1 U19121 ( .A1(n16106), .A2(n19014), .B1(n19041), .B2(n10005), .ZN(
        n16107) );
  INV_X1 U19122 ( .A(n16107), .ZN(n16116) );
  INV_X1 U19123 ( .A(n16108), .ZN(n16110) );
  AOI22_X1 U19124 ( .A1(n16110), .A2(n10916), .B1(n16109), .B2(n19029), .ZN(
        n16115) );
  OAI211_X1 U19125 ( .C1(n16113), .C2(n16112), .A(n18915), .B(n16111), .ZN(
        n16114) );
  NAND4_X1 U19126 ( .A1(n16117), .A2(n16116), .A3(n16115), .A4(n16114), .ZN(
        P2_U2829) );
  AOI22_X1 U19127 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n18957), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19028), .ZN(n16131) );
  OR2_X1 U19128 ( .A1(n16118), .A2(n19014), .ZN(n16120) );
  NAND2_X1 U19129 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19003), .ZN(
        n16119) );
  AND2_X1 U19130 ( .A1(n16120), .A2(n16119), .ZN(n16130) );
  INV_X1 U19131 ( .A(n16121), .ZN(n16122) );
  OAI22_X1 U19132 ( .A1(n16123), .A2(n19037), .B1(n16122), .B2(n19026), .ZN(
        n16124) );
  INV_X1 U19133 ( .A(n16124), .ZN(n16129) );
  OAI211_X1 U19134 ( .C1(n16127), .C2(n16126), .A(n18915), .B(n16125), .ZN(
        n16128) );
  NAND4_X1 U19135 ( .A1(n16131), .A2(n16130), .A3(n16129), .A4(n16128), .ZN(
        P2_U2830) );
  AOI22_X1 U19136 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n18957), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n19028), .ZN(n16140) );
  AOI22_X1 U19137 ( .A1(n9794), .A2(n19035), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n19003), .ZN(n16139) );
  NOR2_X1 U19138 ( .A1(n19026), .A2(n16142), .ZN(n16132) );
  AOI21_X1 U19139 ( .B1(n16133), .B2(n10916), .A(n16132), .ZN(n16138) );
  OAI211_X1 U19140 ( .C1(n16136), .C2(n16135), .A(n18915), .B(n16134), .ZN(
        n16137) );
  NAND4_X1 U19141 ( .A1(n16140), .A2(n16139), .A3(n16138), .A4(n16137), .ZN(
        P2_U2831) );
  INV_X1 U19142 ( .A(n16141), .ZN(n16148) );
  AOI22_X1 U19143 ( .A1(n16148), .A2(n19068), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n19105), .ZN(n16147) );
  AOI22_X1 U19144 ( .A1(n19047), .A2(BUF2_REG_24__SCAN_IN), .B1(n19049), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n16146) );
  INV_X1 U19145 ( .A(n16142), .ZN(n16143) );
  AOI22_X1 U19146 ( .A1(n16144), .A2(n19107), .B1(n19106), .B2(n16143), .ZN(
        n16145) );
  NAND3_X1 U19147 ( .A1(n16147), .A2(n16146), .A3(n16145), .ZN(P2_U2895) );
  AOI22_X1 U19148 ( .A1(n16148), .A2(n19075), .B1(P2_EAX_REG_21__SCAN_IN), 
        .B2(n19105), .ZN(n16153) );
  AOI22_X1 U19149 ( .A1(n19047), .A2(BUF2_REG_21__SCAN_IN), .B1(n19049), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n16152) );
  AOI22_X1 U19150 ( .A1(n16150), .A2(n19107), .B1(n19106), .B2(n16149), .ZN(
        n16151) );
  NAND3_X1 U19151 ( .A1(n16153), .A2(n16152), .A3(n16151), .ZN(P2_U2898) );
  OAI22_X1 U19152 ( .A1(n18918), .A2(n16194), .B1(n10877), .B2(n19012), .ZN(
        n16154) );
  AOI21_X1 U19153 ( .B1(n16187), .B2(n18909), .A(n16154), .ZN(n16158) );
  AOI22_X1 U19154 ( .A1(n16156), .A2(n16190), .B1(n16188), .B2(n16155), .ZN(
        n16157) );
  OAI211_X1 U19155 ( .C1(n16186), .C2(n18912), .A(n16158), .B(n16157), .ZN(
        P2_U2995) );
  AOI22_X1 U19156 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19190), .B1(
        P2_REIP_REG_18__SCAN_IN), .B2(n19206), .ZN(n16164) );
  OAI22_X1 U19157 ( .A1(n16160), .A2(n19197), .B1(n16159), .B2(n19198), .ZN(
        n16161) );
  AOI21_X1 U19158 ( .B1(n19201), .B2(n16162), .A(n16161), .ZN(n16163) );
  OAI211_X1 U19159 ( .C1(n19205), .C2(n16165), .A(n16164), .B(n16163), .ZN(
        P2_U2996) );
  AOI22_X1 U19160 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n19206), .B1(n16187), 
        .B2(n16166), .ZN(n16171) );
  AOI222_X1 U19161 ( .A1(n16169), .A2(n16190), .B1(n16188), .B2(n16168), .C1(
        n19201), .C2(n16167), .ZN(n16170) );
  OAI211_X1 U19162 ( .C1(n20775), .C2(n16194), .A(n16171), .B(n16170), .ZN(
        P2_U2999) );
  AOI22_X1 U19163 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19206), .B1(n16187), 
        .B2(n18977), .ZN(n16178) );
  NOR2_X1 U19164 ( .A1(n16172), .A2(n19197), .ZN(n16176) );
  OAI22_X1 U19165 ( .A1(n16173), .A2(n19198), .B1(n16186), .B2(n18982), .ZN(
        n16174) );
  AOI21_X1 U19166 ( .B1(n16176), .B2(n16175), .A(n16174), .ZN(n16177) );
  OAI211_X1 U19167 ( .C1(n16179), .C2(n16194), .A(n16178), .B(n16177), .ZN(
        P2_U3005) );
  OAI22_X1 U19168 ( .A1(n20789), .A2(n16194), .B1(n10824), .B2(n19012), .ZN(
        n16180) );
  AOI21_X1 U19169 ( .B1(n16187), .B2(n18988), .A(n16180), .ZN(n16185) );
  INV_X1 U19170 ( .A(n16181), .ZN(n16183) );
  AOI22_X1 U19171 ( .A1(n16183), .A2(n16188), .B1(n16190), .B2(n16182), .ZN(
        n16184) );
  OAI211_X1 U19172 ( .C1(n16186), .C2(n18993), .A(n16185), .B(n16184), .ZN(
        P2_U3007) );
  AOI22_X1 U19173 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19206), .B1(n16187), 
        .B2(n19021), .ZN(n16193) );
  AOI222_X1 U19174 ( .A1(n16191), .A2(n16190), .B1(n16189), .B2(n16188), .C1(
        n19201), .C2(n19022), .ZN(n16192) );
  OAI211_X1 U19175 ( .C1(n20749), .C2(n16194), .A(n16193), .B(n16192), .ZN(
        P2_U3009) );
  XNOR2_X1 U19176 ( .A(n16196), .B(n16195), .ZN(n19059) );
  OAI22_X1 U19177 ( .A1(n16197), .A2(n19059), .B1(n10848), .B2(n19012), .ZN(
        n16198) );
  AOI211_X1 U19178 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n16200), .A(
        n16199), .B(n16198), .ZN(n16203) );
  AOI22_X1 U19179 ( .A1(n16201), .A2(n16223), .B1(n19212), .B2(n18970), .ZN(
        n16202) );
  OAI211_X1 U19180 ( .C1(n16204), .C2(n16227), .A(n16203), .B(n16202), .ZN(
        P2_U3034) );
  OAI221_X1 U19181 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n16208), 
        .C1(n16207), .C2(n16206), .A(n16205), .ZN(n16209) );
  AOI21_X1 U19182 ( .B1(n19062), .B2(n19208), .A(n16209), .ZN(n16213) );
  AOI22_X1 U19183 ( .A1(n16211), .A2(n16223), .B1(n19212), .B2(n16210), .ZN(
        n16212) );
  OAI211_X1 U19184 ( .C1(n16214), .C2(n16227), .A(n16213), .B(n16212), .ZN(
        P2_U3036) );
  NOR2_X1 U19185 ( .A1(n19012), .A2(n10830), .ZN(n16221) );
  OAI21_X1 U19186 ( .B1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n16215), .ZN(n16218) );
  OAI22_X1 U19187 ( .A1(n16219), .A2(n16218), .B1(n16217), .B2(n16216), .ZN(
        n16220) );
  AOI211_X1 U19188 ( .C1(n19067), .C2(n19208), .A(n16221), .B(n16220), .ZN(
        n16226) );
  AOI22_X1 U19189 ( .A1(n16224), .A2(n16223), .B1(n19212), .B2(n16222), .ZN(
        n16225) );
  OAI211_X1 U19190 ( .C1(n16228), .C2(n16227), .A(n16226), .B(n16225), .ZN(
        P2_U3038) );
  NAND2_X1 U19191 ( .A1(n16229), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16236) );
  INV_X1 U19192 ( .A(n16236), .ZN(n16232) );
  INV_X1 U19193 ( .A(n16230), .ZN(n16231) );
  OAI211_X1 U19194 ( .C1(n16237), .C2(n16232), .A(n16231), .B(n16233), .ZN(
        n16239) );
  NAND2_X1 U19195 ( .A1(n16234), .A2(n16233), .ZN(n16235) );
  OAI211_X1 U19196 ( .C1(n16237), .C2(n16236), .A(n16235), .B(n12541), .ZN(
        n16238) );
  MUX2_X1 U19197 ( .A(n16239), .B(n16238), .S(n10809), .Z(n16240) );
  AOI21_X1 U19198 ( .B1(n13777), .B2(n16241), .A(n16240), .ZN(n19809) );
  NOR2_X1 U19199 ( .A1(n16281), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n16243) );
  AOI21_X1 U19200 ( .B1(n19809), .B2(n16281), .A(n16243), .ZN(n16284) );
  NOR2_X1 U19201 ( .A1(n16281), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n16244) );
  AOI21_X1 U19202 ( .B1(n16245), .B2(n16281), .A(n16244), .ZN(n16283) );
  INV_X1 U19203 ( .A(n16246), .ZN(n16247) );
  NOR2_X1 U19204 ( .A1(n12376), .A2(n16247), .ZN(n16251) );
  INV_X1 U19205 ( .A(n16248), .ZN(n16250) );
  OR2_X1 U19206 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n16251), .ZN(
        n16249) );
  AOI22_X1 U19207 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n16251), .B1(
        n16250), .B2(n16249), .ZN(n16253) );
  INV_X1 U19208 ( .A(n16283), .ZN(n16256) );
  NAND2_X1 U19209 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n16256), .ZN(
        n16252) );
  OAI211_X1 U19210 ( .C1(n16284), .C2(n19824), .A(n16253), .B(n16252), .ZN(
        n16254) );
  INV_X1 U19211 ( .A(n16254), .ZN(n16258) );
  INV_X1 U19212 ( .A(n16284), .ZN(n16255) );
  OAI21_X1 U19213 ( .B1(n16256), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n16255), .ZN(n16257) );
  AOI22_X1 U19214 ( .A1(n16258), .A2(n16281), .B1(n19824), .B2(n16257), .ZN(
        n16261) );
  NAND3_X1 U19215 ( .A1(n10752), .A2(n10723), .A3(n16259), .ZN(n16260) );
  OAI21_X1 U19216 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n16261), .A(
        n16260), .ZN(n16268) );
  INV_X1 U19217 ( .A(n16262), .ZN(n16264) );
  NOR3_X1 U19218 ( .A1(n16265), .A2(n16264), .A3(n16263), .ZN(n18881) );
  OAI21_X1 U19219 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n18881), .ZN(n16266) );
  INV_X1 U19220 ( .A(n16266), .ZN(n16267) );
  AOI211_X1 U19221 ( .C1(n16270), .C2(n16269), .A(n16268), .B(n16267), .ZN(
        n16279) );
  NAND2_X1 U19222 ( .A1(n16272), .A2(n16271), .ZN(n16278) );
  NOR2_X1 U19223 ( .A1(n10722), .A2(n16273), .ZN(n16274) );
  AOI21_X1 U19224 ( .B1(n16276), .B2(n16275), .A(n16274), .ZN(n16277) );
  AND2_X1 U19225 ( .A1(n16278), .A2(n16277), .ZN(n19858) );
  OAI211_X1 U19226 ( .C1(n16281), .C2(n16280), .A(n16279), .B(n19858), .ZN(
        n16282) );
  AOI21_X1 U19227 ( .B1(n16284), .B2(n16283), .A(n16282), .ZN(n16297) );
  AOI211_X1 U19228 ( .C1(n19853), .C2(n16298), .A(n16286), .B(n16285), .ZN(
        n16296) );
  AOI21_X1 U19229 ( .B1(n16297), .B2(n16287), .A(n18874), .ZN(n16290) );
  NOR3_X1 U19230 ( .A1(n10760), .A2(n9743), .A3(n16288), .ZN(n16289) );
  AOI21_X1 U19231 ( .B1(n18874), .B2(n19810), .A(n19866), .ZN(n16292) );
  INV_X1 U19232 ( .A(n16292), .ZN(n16294) );
  INV_X1 U19233 ( .A(n19867), .ZN(n19865) );
  NAND2_X1 U19234 ( .A1(n19737), .A2(n19865), .ZN(n16293) );
  AOI22_X1 U19235 ( .A1(n19737), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n16294), 
        .B2(n16293), .ZN(n16295) );
  OAI211_X1 U19236 ( .C1(n16297), .C2(n18880), .A(n16296), .B(n16295), .ZN(
        P2_U3176) );
  AOI221_X1 U19237 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n18874), .C1(
        P2_STATE2_REG_3__SCAN_IN), .C2(n19737), .A(n16298), .ZN(n16299) );
  INV_X1 U19238 ( .A(n16299), .ZN(P2_U3593) );
  NAND2_X1 U19239 ( .A1(n17784), .A2(n16300), .ZN(n16314) );
  NAND2_X1 U19240 ( .A1(n17869), .A2(n16301), .ZN(n16316) );
  NAND2_X1 U19241 ( .A1(n17944), .A2(n17658), .ZN(n17612) );
  NOR2_X1 U19242 ( .A1(n17954), .A2(n17612), .ZN(n17595) );
  INV_X1 U19243 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16489) );
  XNOR2_X1 U19244 ( .A(n16489), .B(n16321), .ZN(n16488) );
  AOI21_X1 U19245 ( .B1(n9758), .B2(n16488), .A(n16305), .ZN(n16306) );
  OAI221_X1 U19246 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16308), .C1(
        n16489), .C2(n16307), .A(n16306), .ZN(n16309) );
  INV_X1 U19247 ( .A(n16311), .ZN(n16312) );
  AOI22_X1 U19248 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n16313), .B1(
        n9849), .B2(n16312), .ZN(n16327) );
  INV_X1 U19249 ( .A(n16341), .ZN(n16315) );
  AOI21_X1 U19250 ( .B1(n16317), .B2(n16315), .A(n16314), .ZN(n16319) );
  AOI21_X1 U19251 ( .B1(n16317), .B2(n16340), .A(n16316), .ZN(n16318) );
  AOI211_X1 U19252 ( .C1(n16320), .C2(n17783), .A(n16319), .B(n16318), .ZN(
        n16326) );
  NAND2_X1 U19253 ( .A1(n9726), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16325) );
  INV_X1 U19254 ( .A(n16474), .ZN(n16322) );
  AOI21_X1 U19255 ( .B1(n9981), .B2(n16322), .A(n16321), .ZN(n16498) );
  OAI21_X1 U19256 ( .B1(n16323), .B2(n9758), .A(n16498), .ZN(n16324) );
  NAND4_X1 U19257 ( .A1(n16327), .A2(n16326), .A3(n16325), .A4(n16324), .ZN(
        P3_U2801) );
  INV_X1 U19258 ( .A(n18113), .ZN(n18044) );
  AOI221_X1 U19259 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16328), 
        .C1(n18180), .C2(n16328), .A(n18815), .ZN(n16329) );
  AOI211_X1 U19260 ( .C1(n16332), .C2(n16331), .A(n16330), .B(n16329), .ZN(
        n16335) );
  INV_X1 U19261 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18789) );
  AOI22_X1 U19262 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n12900), .B1(
        n17782), .B2(n12905), .ZN(n17516) );
  AOI21_X1 U19263 ( .B1(n17527), .B2(n17782), .A(n17526), .ZN(n17517) );
  NOR2_X1 U19264 ( .A1(n17516), .A2(n17517), .ZN(n17515) );
  OR2_X1 U19265 ( .A1(n16341), .A2(n18072), .ZN(n16342) );
  NOR2_X1 U19266 ( .A1(n18679), .A2(n18185), .ZN(n18136) );
  NAND2_X1 U19267 ( .A1(n17782), .A2(n18136), .ZN(n16349) );
  OAI22_X1 U19268 ( .A1(n18070), .A2(n18684), .B1(n13073), .B2(n18072), .ZN(
        n18057) );
  AOI21_X1 U19269 ( .B1(n16347), .B2(n18057), .A(n16346), .ZN(n17964) );
  NOR2_X1 U19270 ( .A1(n17964), .A2(n17601), .ZN(n17951) );
  NAND2_X1 U19271 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17951), .ZN(
        n17934) );
  OAI22_X1 U19272 ( .A1(n17515), .A2(n16349), .B1(n16348), .B2(n17934), .ZN(
        n16350) );
  NOR3_X1 U19273 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16352) );
  NOR4_X1 U19274 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16351) );
  NAND4_X1 U19275 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16352), .A3(n16351), .A4(
        U215), .ZN(U213) );
  INV_X1 U19276 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19120) );
  INV_X2 U19277 ( .A(U214), .ZN(n16394) );
  NOR2_X2 U19278 ( .A1(n16394), .A2(n16353), .ZN(n16392) );
  OAI222_X1 U19279 ( .A1(U212), .A2(n19120), .B1(n16397), .B2(n16354), .C1(
        U214), .C2(n16425), .ZN(U216) );
  INV_X1 U19280 ( .A(U212), .ZN(n16395) );
  AOI222_X1 U19281 ( .A1(n16394), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16392), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n16395), .C2(P2_DATAO_REG_30__SCAN_IN), 
        .ZN(n16355) );
  INV_X1 U19282 ( .A(n16355), .ZN(U217) );
  AOI222_X1 U19283 ( .A1(n16394), .A2(P1_DATAO_REG_29__SCAN_IN), .B1(n16392), 
        .B2(BUF1_REG_29__SCAN_IN), .C1(n16395), .C2(P2_DATAO_REG_29__SCAN_IN), 
        .ZN(n16356) );
  INV_X1 U19284 ( .A(n16356), .ZN(U218) );
  AOI22_X1 U19285 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n16395), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n16394), .ZN(n16357) );
  OAI21_X1 U19286 ( .B1(n19233), .B2(n16397), .A(n16357), .ZN(U219) );
  INV_X1 U19287 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n19227) );
  AOI22_X1 U19288 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(n16395), .B1(
        P1_DATAO_REG_27__SCAN_IN), .B2(n16394), .ZN(n16358) );
  OAI21_X1 U19289 ( .B1(n19227), .B2(n16397), .A(n16358), .ZN(U220) );
  AOI22_X1 U19290 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n16395), .B1(
        P1_DATAO_REG_26__SCAN_IN), .B2(n16394), .ZN(n16359) );
  OAI21_X1 U19291 ( .B1(n16360), .B2(n16397), .A(n16359), .ZN(U221) );
  AOI222_X1 U19292 ( .A1(n16394), .A2(P1_DATAO_REG_25__SCAN_IN), .B1(n16392), 
        .B2(BUF1_REG_25__SCAN_IN), .C1(n16395), .C2(P2_DATAO_REG_25__SCAN_IN), 
        .ZN(n16361) );
  INV_X1 U19293 ( .A(n16361), .ZN(U222) );
  AOI22_X1 U19294 ( .A1(P2_DATAO_REG_24__SCAN_IN), .A2(n16395), .B1(
        P1_DATAO_REG_24__SCAN_IN), .B2(n16394), .ZN(n16362) );
  OAI21_X1 U19295 ( .B1(n14382), .B2(n16397), .A(n16362), .ZN(U223) );
  INV_X1 U19296 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n16364) );
  AOI22_X1 U19297 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(n16395), .B1(
        P1_DATAO_REG_23__SCAN_IN), .B2(n16394), .ZN(n16363) );
  OAI21_X1 U19298 ( .B1(n16364), .B2(n16397), .A(n16363), .ZN(U224) );
  AOI22_X1 U19299 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(n16395), .B1(
        P1_DATAO_REG_22__SCAN_IN), .B2(n16394), .ZN(n16365) );
  OAI21_X1 U19300 ( .B1(n15002), .B2(n16397), .A(n16365), .ZN(U225) );
  INV_X1 U19301 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n16367) );
  AOI22_X1 U19302 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n16395), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n16394), .ZN(n16366) );
  OAI21_X1 U19303 ( .B1(n16367), .B2(n16397), .A(n16366), .ZN(U226) );
  AOI22_X1 U19304 ( .A1(P2_DATAO_REG_20__SCAN_IN), .A2(n16395), .B1(
        P1_DATAO_REG_20__SCAN_IN), .B2(n16394), .ZN(n16368) );
  OAI21_X1 U19305 ( .B1(n15008), .B2(n16397), .A(n16368), .ZN(U227) );
  AOI22_X1 U19306 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n16395), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n16394), .ZN(n16369) );
  OAI21_X1 U19307 ( .B1(n15018), .B2(n16397), .A(n16369), .ZN(U228) );
  AOI22_X1 U19308 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n16395), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n16394), .ZN(n16370) );
  OAI21_X1 U19309 ( .B1(n16371), .B2(n16397), .A(n16370), .ZN(U229) );
  AOI22_X1 U19310 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n16395), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n16394), .ZN(n16372) );
  OAI21_X1 U19311 ( .B1(n14006), .B2(n16397), .A(n16372), .ZN(U230) );
  AOI222_X1 U19312 ( .A1(n16395), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n16392), 
        .B2(BUF1_REG_16__SCAN_IN), .C1(n16394), .C2(P1_DATAO_REG_16__SCAN_IN), 
        .ZN(n16373) );
  INV_X1 U19313 ( .A(n16373), .ZN(U231) );
  AOI22_X1 U19314 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n16395), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n16394), .ZN(n16374) );
  OAI21_X1 U19315 ( .B1(n13355), .B2(n16397), .A(n16374), .ZN(U232) );
  AOI22_X1 U19316 ( .A1(P2_DATAO_REG_14__SCAN_IN), .A2(n16395), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16394), .ZN(n16375) );
  OAI21_X1 U19317 ( .B1(n12718), .B2(n16397), .A(n16375), .ZN(U233) );
  INV_X1 U19318 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n20965) );
  AOI22_X1 U19319 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n16392), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16395), .ZN(n16376) );
  OAI21_X1 U19320 ( .B1(n20965), .B2(U214), .A(n16376), .ZN(U234) );
  INV_X1 U19321 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16378) );
  AOI22_X1 U19322 ( .A1(BUF1_REG_12__SCAN_IN), .A2(n16392), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n16394), .ZN(n16377) );
  OAI21_X1 U19323 ( .B1(n16378), .B2(U212), .A(n16377), .ZN(U235) );
  INV_X1 U19324 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16380) );
  AOI22_X1 U19325 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n16392), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16394), .ZN(n16379) );
  OAI21_X1 U19326 ( .B1(n16380), .B2(U212), .A(n16379), .ZN(U236) );
  INV_X1 U19327 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n19160) );
  AOI22_X1 U19328 ( .A1(BUF1_REG_10__SCAN_IN), .A2(n16392), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16394), .ZN(n16381) );
  OAI21_X1 U19329 ( .B1(n19160), .B2(U212), .A(n16381), .ZN(U237) );
  INV_X1 U19330 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n19162) );
  AOI22_X1 U19331 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n16392), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n16394), .ZN(n16382) );
  OAI21_X1 U19332 ( .B1(n19162), .B2(U212), .A(n16382), .ZN(U238) );
  INV_X1 U19333 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16405) );
  INV_X1 U19334 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n20950) );
  OAI222_X1 U19335 ( .A1(U212), .A2(n16405), .B1(n16397), .B2(n16383), .C1(
        U214), .C2(n20950), .ZN(U239) );
  INV_X1 U19336 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16404) );
  AOI22_X1 U19337 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16392), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16394), .ZN(n16384) );
  OAI21_X1 U19338 ( .B1(n16404), .B2(U212), .A(n16384), .ZN(U240) );
  INV_X1 U19339 ( .A(BUF1_REG_6__SCAN_IN), .ZN(n16386) );
  AOI22_X1 U19340 ( .A1(P2_DATAO_REG_6__SCAN_IN), .A2(n16395), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16394), .ZN(n16385) );
  OAI21_X1 U19341 ( .B1(n16386), .B2(n16397), .A(n16385), .ZN(U241) );
  INV_X1 U19342 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16388) );
  AOI22_X1 U19343 ( .A1(P2_DATAO_REG_5__SCAN_IN), .A2(n16395), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n16394), .ZN(n16387) );
  OAI21_X1 U19344 ( .B1(n16388), .B2(n16397), .A(n16387), .ZN(U242) );
  AOI222_X1 U19345 ( .A1(n16394), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n16392), 
        .B2(BUF1_REG_4__SCAN_IN), .C1(n16395), .C2(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n16389) );
  INV_X1 U19346 ( .A(n16389), .ZN(U243) );
  INV_X1 U19347 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16401) );
  AOI22_X1 U19348 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16392), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16394), .ZN(n16390) );
  OAI21_X1 U19349 ( .B1(n16401), .B2(U212), .A(n16390), .ZN(U244) );
  INV_X1 U19350 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n16400) );
  AOI22_X1 U19351 ( .A1(BUF1_REG_2__SCAN_IN), .A2(n16392), .B1(
        P1_DATAO_REG_2__SCAN_IN), .B2(n16394), .ZN(n16391) );
  OAI21_X1 U19352 ( .B1(n16400), .B2(U212), .A(n16391), .ZN(U245) );
  INV_X1 U19353 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n16399) );
  AOI22_X1 U19354 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n16392), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n16394), .ZN(n16393) );
  OAI21_X1 U19355 ( .B1(n16399), .B2(U212), .A(n16393), .ZN(U246) );
  INV_X1 U19356 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n20871) );
  AOI22_X1 U19357 ( .A1(P2_DATAO_REG_0__SCAN_IN), .A2(n16395), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16394), .ZN(n16396) );
  OAI21_X1 U19358 ( .B1(n20871), .B2(n16397), .A(n16396), .ZN(U247) );
  OAI22_X1 U19359 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16424), .ZN(n16398) );
  INV_X1 U19360 ( .A(n16398), .ZN(U251) );
  INV_X1 U19361 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n20954) );
  AOI22_X1 U19362 ( .A1(n16424), .A2(n16399), .B1(n20954), .B2(U215), .ZN(U252) );
  INV_X1 U19363 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n20804) );
  AOI22_X1 U19364 ( .A1(n16424), .A2(n16400), .B1(n20804), .B2(U215), .ZN(U253) );
  INV_X1 U19365 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18224) );
  AOI22_X1 U19366 ( .A1(n16424), .A2(n16401), .B1(n18224), .B2(U215), .ZN(U254) );
  INV_X1 U19367 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n19172) );
  INV_X1 U19368 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18228) );
  AOI22_X1 U19369 ( .A1(n16424), .A2(n19172), .B1(n18228), .B2(U215), .ZN(U255) );
  OAI22_X1 U19370 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16424), .ZN(n16402) );
  INV_X1 U19371 ( .A(n16402), .ZN(U256) );
  OAI22_X1 U19372 ( .A1(U215), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n16424), .ZN(n16403) );
  INV_X1 U19373 ( .A(n16403), .ZN(U257) );
  INV_X1 U19374 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18242) );
  AOI22_X1 U19375 ( .A1(n16424), .A2(n16404), .B1(n18242), .B2(U215), .ZN(U258) );
  AOI22_X1 U19376 ( .A1(n16423), .A2(n16405), .B1(n17489), .B2(U215), .ZN(U259) );
  INV_X1 U19377 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17492) );
  AOI22_X1 U19378 ( .A1(n16424), .A2(n19162), .B1(n17492), .B2(U215), .ZN(U260) );
  INV_X1 U19379 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17496) );
  AOI22_X1 U19380 ( .A1(n16423), .A2(n19160), .B1(n17496), .B2(U215), .ZN(U261) );
  OAI22_X1 U19381 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16423), .ZN(n16406) );
  INV_X1 U19382 ( .A(n16406), .ZN(U262) );
  OAI22_X1 U19383 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16423), .ZN(n16407) );
  INV_X1 U19384 ( .A(n16407), .ZN(U263) );
  OAI22_X1 U19385 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16423), .ZN(n16408) );
  INV_X1 U19386 ( .A(n16408), .ZN(U264) );
  OAI22_X1 U19387 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16423), .ZN(n16409) );
  INV_X1 U19388 ( .A(n16409), .ZN(U265) );
  OAI22_X1 U19389 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16423), .ZN(n16410) );
  INV_X1 U19390 ( .A(n16410), .ZN(U266) );
  OAI22_X1 U19391 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16424), .ZN(n16411) );
  INV_X1 U19392 ( .A(n16411), .ZN(U267) );
  OAI22_X1 U19393 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16423), .ZN(n16412) );
  INV_X1 U19394 ( .A(n16412), .ZN(U268) );
  OAI22_X1 U19395 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16424), .ZN(n16413) );
  INV_X1 U19396 ( .A(n16413), .ZN(U269) );
  OAI22_X1 U19397 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16424), .ZN(n16414) );
  INV_X1 U19398 ( .A(n16414), .ZN(U270) );
  OAI22_X1 U19399 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16424), .ZN(n16415) );
  INV_X1 U19400 ( .A(n16415), .ZN(U271) );
  OAI22_X1 U19401 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16424), .ZN(n16416) );
  INV_X1 U19402 ( .A(n16416), .ZN(U272) );
  OAI22_X1 U19403 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16424), .ZN(n16417) );
  INV_X1 U19404 ( .A(n16417), .ZN(U273) );
  OAI22_X1 U19405 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16424), .ZN(n16418) );
  INV_X1 U19406 ( .A(n16418), .ZN(U274) );
  OAI22_X1 U19407 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16424), .ZN(n16419) );
  INV_X1 U19408 ( .A(n16419), .ZN(U275) );
  INV_X1 U19409 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n20850) );
  INV_X1 U19410 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18216) );
  AOI22_X1 U19411 ( .A1(n16423), .A2(n20850), .B1(n18216), .B2(U215), .ZN(U276) );
  OAI22_X1 U19412 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16424), .ZN(n16420) );
  INV_X1 U19413 ( .A(n16420), .ZN(U277) );
  OAI22_X1 U19414 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16424), .ZN(n16421) );
  INV_X1 U19415 ( .A(n16421), .ZN(U278) );
  OAI22_X1 U19416 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16424), .ZN(n16422) );
  INV_X1 U19417 ( .A(n16422), .ZN(U279) );
  INV_X1 U19418 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n20773) );
  INV_X1 U19419 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18232) );
  AOI22_X1 U19420 ( .A1(n16424), .A2(n20773), .B1(n18232), .B2(U215), .ZN(U280) );
  INV_X1 U19421 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19123) );
  INV_X1 U19422 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n19244) );
  AOI22_X1 U19423 ( .A1(n16423), .A2(n19123), .B1(n19244), .B2(U215), .ZN(U281) );
  INV_X1 U19424 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18241) );
  AOI22_X1 U19425 ( .A1(n16424), .A2(n19120), .B1(n18241), .B2(U215), .ZN(U282) );
  INV_X1 U19426 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n17398) );
  AOI222_X1 U19427 ( .A1(n19120), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16425), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .C1(n17398), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16426) );
  INV_X2 U19428 ( .A(n16428), .ZN(n16427) );
  INV_X1 U19429 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n21025) );
  INV_X1 U19430 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19769) );
  AOI22_X1 U19431 ( .A1(n16427), .A2(n21025), .B1(n19769), .B2(n16428), .ZN(
        U347) );
  INV_X1 U19432 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n20812) );
  INV_X1 U19433 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n20905) );
  AOI22_X1 U19434 ( .A1(n16427), .A2(n20812), .B1(n20905), .B2(n16428), .ZN(
        U348) );
  INV_X1 U19435 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18750) );
  INV_X1 U19436 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19768) );
  AOI22_X1 U19437 ( .A1(n16427), .A2(n18750), .B1(n19768), .B2(n16428), .ZN(
        U349) );
  INV_X1 U19438 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n20770) );
  INV_X1 U19439 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19767) );
  AOI22_X1 U19440 ( .A1(n16427), .A2(n20770), .B1(n19767), .B2(n16428), .ZN(
        U350) );
  INV_X1 U19441 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18748) );
  INV_X1 U19442 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19766) );
  AOI22_X1 U19443 ( .A1(n16427), .A2(n18748), .B1(n19766), .B2(n16428), .ZN(
        U351) );
  INV_X1 U19444 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18746) );
  INV_X1 U19445 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19764) );
  AOI22_X1 U19446 ( .A1(n16427), .A2(n18746), .B1(n19764), .B2(n16428), .ZN(
        U352) );
  INV_X1 U19447 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18745) );
  AOI22_X1 U19448 ( .A1(n16427), .A2(n18745), .B1(n19763), .B2(n16428), .ZN(
        U353) );
  INV_X1 U19449 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18743) );
  INV_X1 U19450 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19762) );
  AOI22_X1 U19451 ( .A1(n16427), .A2(n18743), .B1(n19762), .B2(n16428), .ZN(
        U354) );
  INV_X1 U19452 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18794) );
  INV_X1 U19453 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19799) );
  AOI22_X1 U19454 ( .A1(n16427), .A2(n18794), .B1(n19799), .B2(n16428), .ZN(
        U355) );
  INV_X1 U19455 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18791) );
  INV_X1 U19456 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19796) );
  AOI22_X1 U19457 ( .A1(n16427), .A2(n18791), .B1(n19796), .B2(n16428), .ZN(
        U356) );
  INV_X1 U19458 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18788) );
  INV_X1 U19459 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19794) );
  AOI22_X1 U19460 ( .A1(n16427), .A2(n18788), .B1(n19794), .B2(n16428), .ZN(
        U357) );
  INV_X1 U19461 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18787) );
  INV_X1 U19462 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19791) );
  AOI22_X1 U19463 ( .A1(n16427), .A2(n18787), .B1(n19791), .B2(n16428), .ZN(
        U358) );
  INV_X1 U19464 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18785) );
  INV_X1 U19465 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19790) );
  AOI22_X1 U19466 ( .A1(n16427), .A2(n18785), .B1(n19790), .B2(n16428), .ZN(
        U359) );
  INV_X1 U19467 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18783) );
  INV_X1 U19468 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19789) );
  AOI22_X1 U19469 ( .A1(n16427), .A2(n18783), .B1(n19789), .B2(n16428), .ZN(
        U360) );
  INV_X1 U19470 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18780) );
  INV_X1 U19471 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19787) );
  AOI22_X1 U19472 ( .A1(n16427), .A2(n18780), .B1(n19787), .B2(n16428), .ZN(
        U361) );
  INV_X1 U19473 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18778) );
  INV_X1 U19474 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19785) );
  AOI22_X1 U19475 ( .A1(n16427), .A2(n18778), .B1(n19785), .B2(n16428), .ZN(
        U362) );
  INV_X1 U19476 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18776) );
  INV_X1 U19477 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19784) );
  AOI22_X1 U19478 ( .A1(n16427), .A2(n18776), .B1(n19784), .B2(n16428), .ZN(
        U363) );
  INV_X1 U19479 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18774) );
  INV_X1 U19480 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19782) );
  AOI22_X1 U19481 ( .A1(n16427), .A2(n18774), .B1(n19782), .B2(n16428), .ZN(
        U364) );
  INV_X1 U19482 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18741) );
  INV_X1 U19483 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n20803) );
  AOI22_X1 U19484 ( .A1(n16427), .A2(n18741), .B1(n20803), .B2(n16428), .ZN(
        U365) );
  INV_X1 U19485 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18772) );
  INV_X1 U19486 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19781) );
  AOI22_X1 U19487 ( .A1(n16427), .A2(n18772), .B1(n19781), .B2(n16428), .ZN(
        U366) );
  INV_X1 U19488 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18770) );
  INV_X1 U19489 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19780) );
  AOI22_X1 U19490 ( .A1(n16427), .A2(n18770), .B1(n19780), .B2(n16428), .ZN(
        U367) );
  INV_X1 U19491 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18768) );
  INV_X1 U19492 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19779) );
  AOI22_X1 U19493 ( .A1(n16427), .A2(n18768), .B1(n19779), .B2(n16428), .ZN(
        U368) );
  INV_X1 U19494 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18766) );
  INV_X1 U19495 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19778) );
  AOI22_X1 U19496 ( .A1(n16427), .A2(n18766), .B1(n19778), .B2(n16428), .ZN(
        U369) );
  INV_X1 U19497 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18764) );
  INV_X1 U19498 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19776) );
  AOI22_X1 U19499 ( .A1(n16427), .A2(n18764), .B1(n19776), .B2(n16428), .ZN(
        U370) );
  INV_X1 U19500 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18762) );
  INV_X1 U19501 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19774) );
  AOI22_X1 U19502 ( .A1(n16427), .A2(n18762), .B1(n19774), .B2(n16428), .ZN(
        U371) );
  INV_X1 U19503 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18759) );
  INV_X1 U19504 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19773) );
  AOI22_X1 U19505 ( .A1(n16427), .A2(n18759), .B1(n19773), .B2(n16428), .ZN(
        U372) );
  INV_X1 U19506 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18758) );
  INV_X1 U19507 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19772) );
  AOI22_X1 U19508 ( .A1(n16427), .A2(n18758), .B1(n19772), .B2(n16428), .ZN(
        U373) );
  INV_X1 U19509 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18756) );
  INV_X1 U19510 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19771) );
  AOI22_X1 U19511 ( .A1(n16427), .A2(n18756), .B1(n19771), .B2(n16428), .ZN(
        U374) );
  INV_X1 U19512 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18754) );
  INV_X1 U19513 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19770) );
  AOI22_X1 U19514 ( .A1(n16427), .A2(n18754), .B1(n19770), .B2(n16428), .ZN(
        U375) );
  INV_X1 U19515 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18738) );
  INV_X1 U19516 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19761) );
  AOI22_X1 U19517 ( .A1(n16427), .A2(n18738), .B1(n19761), .B2(n16428), .ZN(
        U376) );
  NAND2_X1 U19518 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18737), .ZN(n18725) );
  AOI22_X1 U19519 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18725), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n20922), .ZN(n18805) );
  AOI21_X1 U19520 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18805), .ZN(n16429) );
  INV_X1 U19521 ( .A(n16429), .ZN(P3_U2633) );
  INV_X1 U19522 ( .A(n16456), .ZN(n18712) );
  NAND2_X1 U19523 ( .A1(n17446), .A2(n16430), .ZN(n16437) );
  INV_X1 U19524 ( .A(n16437), .ZN(n16431) );
  NAND2_X1 U19525 ( .A1(n18849), .A2(n18682), .ZN(n17445) );
  OAI21_X1 U19526 ( .B1(n16431), .B2(n17445), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16432) );
  OAI21_X1 U19527 ( .B1(n16433), .B2(n18712), .A(n16432), .ZN(P3_U2634) );
  AOI21_X1 U19528 ( .B1(n20922), .B2(n18737), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16434) );
  AOI22_X1 U19529 ( .A1(n18842), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16434), 
        .B2(n18863), .ZN(P3_U2635) );
  INV_X1 U19530 ( .A(BS16), .ZN(n16435) );
  AOI21_X1 U19531 ( .B1(n16436), .B2(n16435), .A(n18802), .ZN(n18801) );
  INV_X1 U19532 ( .A(n18801), .ZN(n18803) );
  OAI21_X1 U19533 ( .B1(n18805), .B2(n18852), .A(n18803), .ZN(P3_U2636) );
  NAND3_X1 U19534 ( .A1(n18682), .A2(n16438), .A3(n16437), .ZN(n18693) );
  NAND2_X1 U19535 ( .A1(n18849), .A2(n18693), .ZN(n18846) );
  INV_X1 U19536 ( .A(n18846), .ZN(n16440) );
  OAI21_X1 U19537 ( .B1(n16440), .B2(n18201), .A(n16439), .ZN(P3_U2637) );
  NOR4_X1 U19538 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16444) );
  NOR4_X1 U19539 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16443) );
  NOR4_X1 U19540 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16442) );
  NOR4_X1 U19541 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16441) );
  NAND4_X1 U19542 ( .A1(n16444), .A2(n16443), .A3(n16442), .A4(n16441), .ZN(
        n16450) );
  NOR4_X1 U19543 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16448) );
  AOI211_X1 U19544 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_12__SCAN_IN), .B(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16447) );
  NOR4_X1 U19545 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16446) );
  NOR4_X1 U19546 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16445) );
  NAND4_X1 U19547 ( .A1(n16448), .A2(n16447), .A3(n16446), .A4(n16445), .ZN(
        n16449) );
  NOR2_X1 U19548 ( .A1(n16450), .A2(n16449), .ZN(n18841) );
  INV_X1 U19549 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16452) );
  NOR3_X1 U19550 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16453) );
  OAI21_X1 U19551 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16453), .A(n18841), .ZN(
        n16451) );
  OAI21_X1 U19552 ( .B1(n18841), .B2(n16452), .A(n16451), .ZN(P3_U2638) );
  INV_X1 U19553 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16455) );
  NOR2_X1 U19554 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18835) );
  OAI21_X1 U19555 ( .B1(n16453), .B2(n18835), .A(n18841), .ZN(n16454) );
  OAI21_X1 U19556 ( .B1(n18841), .B2(n16455), .A(n16454), .ZN(P3_U2639) );
  INV_X1 U19557 ( .A(n18868), .ZN(n18847) );
  AND4_X1 U19558 ( .A1(n20757), .A2(n18865), .A3(n18852), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n16823) );
  NOR2_X2 U19559 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18808), .ZN(n18713) );
  NAND2_X1 U19560 ( .A1(n16456), .A2(n18713), .ZN(n18706) );
  INV_X1 U19561 ( .A(n18854), .ZN(n18710) );
  AOI211_X1 U19562 ( .C1(n18217), .C2(n18851), .A(n18710), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n16458) );
  NAND2_X1 U19563 ( .A1(n18868), .A2(n18853), .ZN(n16461) );
  AOI211_X1 U19564 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n17448), .A(n16458), .B(
        n16461), .ZN(n16457) );
  INV_X1 U19565 ( .A(n16458), .ZN(n18701) );
  INV_X1 U19566 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18782) );
  INV_X1 U19567 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18777) );
  INV_X1 U19568 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18773) );
  INV_X1 U19569 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18769) );
  INV_X1 U19570 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18765) );
  INV_X1 U19571 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18757) );
  INV_X1 U19572 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18753) );
  INV_X1 U19573 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18749) );
  NAND3_X1 U19574 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16782) );
  NOR2_X1 U19575 ( .A1(n18744), .A2(n16782), .ZN(n16766) );
  NAND2_X1 U19576 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16766), .ZN(n16748) );
  NOR3_X1 U19577 ( .A1(n18749), .A2(n18747), .A3(n16748), .ZN(n16735) );
  NAND2_X1 U19578 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16735), .ZN(n16731) );
  NAND2_X1 U19579 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16709) );
  NOR3_X1 U19580 ( .A1(n18753), .A2(n16731), .A3(n16709), .ZN(n16687) );
  NAND2_X1 U19581 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16687), .ZN(n16675) );
  NOR2_X1 U19582 ( .A1(n18757), .A2(n16675), .ZN(n16664) );
  NAND2_X1 U19583 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n16664), .ZN(n16641) );
  NAND2_X1 U19584 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .ZN(n16627) );
  NOR3_X1 U19585 ( .A1(n18765), .A2(n16641), .A3(n16627), .ZN(n16606) );
  NAND2_X1 U19586 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16606), .ZN(n16615) );
  NOR2_X1 U19587 ( .A1(n18769), .A2(n16615), .ZN(n16601) );
  NAND2_X1 U19588 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16601), .ZN(n16584) );
  NOR2_X1 U19589 ( .A1(n18773), .A2(n16584), .ZN(n16580) );
  NAND2_X1 U19590 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16580), .ZN(n16566) );
  NOR2_X1 U19591 ( .A1(n18777), .A2(n16566), .ZN(n16564) );
  NAND2_X1 U19592 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16564), .ZN(n16543) );
  NOR2_X1 U19593 ( .A1(n18782), .A2(n16543), .ZN(n16528) );
  NAND2_X1 U19594 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16528), .ZN(n16476) );
  NOR2_X1 U19595 ( .A1(n16825), .A2(n16476), .ZN(n16521) );
  NAND4_X1 U19596 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .A4(n16521), .ZN(n16479) );
  NOR3_X1 U19597 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18795), .A3(n16479), 
        .ZN(n16459) );
  AOI21_X1 U19598 ( .B1(n16838), .B2(P3_EBX_REG_31__SCAN_IN), .A(n16459), .ZN(
        n16484) );
  NAND2_X1 U19599 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n17448), .ZN(n16460) );
  AOI211_X4 U19600 ( .C1(n18852), .C2(n18854), .A(n16461), .B(n16460), .ZN(
        n16837) );
  NOR3_X1 U19601 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16808) );
  NAND2_X1 U19602 ( .A1(n16808), .A2(n16801), .ZN(n16800) );
  NOR2_X1 U19603 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16800), .ZN(n16784) );
  INV_X1 U19604 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16773) );
  NAND2_X1 U19605 ( .A1(n16784), .A2(n16773), .ZN(n16772) );
  INV_X1 U19606 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17210) );
  NAND2_X1 U19607 ( .A1(n16756), .A2(n17210), .ZN(n16746) );
  NAND2_X1 U19608 ( .A1(n16732), .A2(n17143), .ZN(n16720) );
  NAND2_X1 U19609 ( .A1(n16708), .A2(n16707), .ZN(n16699) );
  INV_X1 U19610 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n21008) );
  NAND2_X1 U19611 ( .A1(n16684), .A2(n21008), .ZN(n16679) );
  INV_X1 U19612 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n20783) );
  NAND2_X1 U19613 ( .A1(n16663), .A2(n20783), .ZN(n16655) );
  INV_X1 U19614 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n20806) );
  NAND2_X1 U19615 ( .A1(n16639), .A2(n20806), .ZN(n16635) );
  INV_X1 U19616 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n20786) );
  NAND2_X1 U19617 ( .A1(n16617), .A2(n20786), .ZN(n16612) );
  INV_X1 U19618 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17012) );
  NAND2_X1 U19619 ( .A1(n16598), .A2(n17012), .ZN(n16588) );
  INV_X1 U19620 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16570) );
  NAND2_X1 U19621 ( .A1(n16574), .A2(n16570), .ZN(n16569) );
  NOR2_X1 U19622 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16569), .ZN(n16540) );
  INV_X1 U19623 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16551) );
  NAND2_X1 U19624 ( .A1(n16540), .A2(n16551), .ZN(n16530) );
  NOR2_X1 U19625 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16530), .ZN(n16529) );
  INV_X1 U19626 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16960) );
  NAND2_X1 U19627 ( .A1(n16529), .A2(n16960), .ZN(n16522) );
  NOR2_X1 U19628 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16522), .ZN(n16507) );
  INV_X1 U19629 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16847) );
  NAND2_X1 U19630 ( .A1(n16507), .A2(n16847), .ZN(n16486) );
  NOR2_X1 U19631 ( .A1(n16827), .A2(n16486), .ZN(n16493) );
  INV_X1 U19632 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16852) );
  OAI21_X1 U19633 ( .B1(n16471), .B2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16475), .ZN(n17529) );
  INV_X1 U19634 ( .A(n17529), .ZN(n16519) );
  NOR2_X1 U19635 ( .A1(n17870), .A2(n17561), .ZN(n16470) );
  AND2_X1 U19636 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n16470), .ZN(
        n16462) );
  NAND2_X1 U19637 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17542), .ZN(
        n16472) );
  OAI21_X1 U19638 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16462), .A(
        n16472), .ZN(n16463) );
  INV_X1 U19639 ( .A(n16463), .ZN(n17554) );
  INV_X1 U19640 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17572) );
  XNOR2_X1 U19641 ( .A(n17572), .B(n16470), .ZN(n17568) );
  INV_X1 U19642 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n16465) );
  INV_X1 U19643 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n16466) );
  NOR2_X1 U19644 ( .A1(n17870), .A2(n17640), .ZN(n17639) );
  INV_X1 U19645 ( .A(n17639), .ZN(n16628) );
  NOR2_X1 U19646 ( .A1(n17641), .A2(n16628), .ZN(n17603) );
  INV_X1 U19647 ( .A(n17603), .ZN(n16607) );
  NOR2_X1 U19648 ( .A1(n16466), .A2(n16607), .ZN(n16468) );
  NAND2_X1 U19649 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16468), .ZN(
        n16464) );
  NAND2_X1 U19650 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17585), .ZN(
        n17552) );
  INV_X1 U19651 ( .A(n17552), .ZN(n17587) );
  AOI21_X1 U19652 ( .B1(n16465), .B2(n16464), .A(n17587), .ZN(n17605) );
  AOI21_X1 U19653 ( .B1(n16466), .B2(n16607), .A(n16468), .ZN(n17633) );
  NAND2_X1 U19654 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16467), .ZN(
        n16673) );
  NOR2_X1 U19655 ( .A1(n9987), .A2(n16673), .ZN(n17677) );
  NAND2_X1 U19656 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17677), .ZN(
        n16651) );
  OAI21_X1 U19657 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16651), .A(
        n16758), .ZN(n16645) );
  NOR2_X1 U19658 ( .A1(n17633), .A2(n16597), .ZN(n16596) );
  NOR2_X1 U19659 ( .A1(n16596), .A2(n16820), .ZN(n16587) );
  INV_X1 U19660 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17617) );
  XNOR2_X1 U19661 ( .A(n17617), .B(n16468), .ZN(n17613) );
  INV_X1 U19662 ( .A(n16820), .ZN(n16469) );
  INV_X1 U19663 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17591) );
  AOI21_X1 U19664 ( .B1(n17591), .B2(n17552), .A(n16470), .ZN(n17588) );
  NOR2_X1 U19665 ( .A1(n16554), .A2(n16820), .ZN(n16542) );
  INV_X1 U19666 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16473) );
  AOI21_X1 U19667 ( .B1(n16473), .B2(n16472), .A(n16471), .ZN(n17543) );
  NOR2_X1 U19668 ( .A1(n16517), .A2(n16820), .ZN(n16510) );
  AOI21_X1 U19669 ( .B1(n16475), .B2(n17512), .A(n16474), .ZN(n17514) );
  NOR4_X1 U19670 ( .A1(n16488), .A2(n16487), .A3(n16820), .A4(n18717), .ZN(
        n16482) );
  NAND3_X1 U19671 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(P3_REIP_REG_27__SCAN_IN), .ZN(n16478) );
  NAND2_X1 U19672 ( .A1(n16807), .A2(n16476), .ZN(n16477) );
  NAND2_X1 U19673 ( .A1(n16783), .A2(n16477), .ZN(n16527) );
  AOI21_X1 U19674 ( .B1(n16807), .B2(n16478), .A(n16527), .ZN(n16506) );
  NOR2_X1 U19675 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16479), .ZN(n16491) );
  INV_X1 U19676 ( .A(n16491), .ZN(n16480) );
  AOI21_X1 U19677 ( .B1(n16506), .B2(n16480), .A(n18792), .ZN(n16481) );
  OAI211_X1 U19678 ( .C1(n16485), .C2(n16804), .A(n16484), .B(n16483), .ZN(
        P3_U2640) );
  NAND2_X1 U19679 ( .A1(n16837), .A2(n16486), .ZN(n16502) );
  OAI22_X1 U19680 ( .A1(n16506), .A2(n18795), .B1(n16489), .B2(n16804), .ZN(
        n16490) );
  AOI211_X1 U19681 ( .C1(n16492), .C2(n16823), .A(n16491), .B(n16490), .ZN(
        n16495) );
  OAI21_X1 U19682 ( .B1(n16838), .B2(n16493), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16494) );
  INV_X1 U19683 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18790) );
  AOI211_X1 U19684 ( .C1(n16498), .C2(n16497), .A(n16496), .B(n18717), .ZN(
        n16501) );
  NAND3_X1 U19685 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_27__SCAN_IN), 
        .A3(n16521), .ZN(n16499) );
  OAI22_X1 U19686 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16499), .B1(n9981), 
        .B2(n16804), .ZN(n16500) );
  AOI211_X1 U19687 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16838), .A(n16501), .B(
        n16500), .ZN(n16505) );
  INV_X1 U19688 ( .A(n16502), .ZN(n16503) );
  OAI21_X1 U19689 ( .B1(n16507), .B2(n16847), .A(n16503), .ZN(n16504) );
  OAI211_X1 U19690 ( .C1(n16506), .C2(n18790), .A(n16505), .B(n16504), .ZN(
        P3_U2642) );
  AOI211_X1 U19691 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16522), .A(n16507), .B(
        n16827), .ZN(n16516) );
  INV_X1 U19692 ( .A(n16508), .ZN(n16509) );
  AOI211_X1 U19693 ( .C1(n17514), .C2(n16510), .A(n16509), .B(n18717), .ZN(
        n16515) );
  NAND2_X1 U19694 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16521), .ZN(n16513) );
  INV_X1 U19695 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18786) );
  AOI21_X1 U19696 ( .B1(n16521), .B2(n18786), .A(n16527), .ZN(n16512) );
  AOI22_X1 U19697 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n16821), .B1(
        n16838), .B2(P3_EBX_REG_28__SCAN_IN), .ZN(n16511) );
  OAI221_X1 U19698 ( .B1(P3_REIP_REG_28__SCAN_IN), .B2(n16513), .C1(n18789), 
        .C2(n16512), .A(n16511), .ZN(n16514) );
  OR3_X1 U19699 ( .A1(n16516), .A2(n16515), .A3(n16514), .ZN(P3_U2643) );
  AOI22_X1 U19700 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n16821), .B1(
        n16838), .B2(P3_EBX_REG_27__SCAN_IN), .ZN(n16526) );
  AOI211_X1 U19701 ( .C1(n16519), .C2(n16518), .A(n16517), .B(n18717), .ZN(
        n16520) );
  AOI21_X1 U19702 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n16527), .A(n16520), 
        .ZN(n16525) );
  NAND2_X1 U19703 ( .A1(n16521), .A2(n18786), .ZN(n16524) );
  OAI211_X1 U19704 ( .C1(n16529), .C2(n16960), .A(n16837), .B(n16522), .ZN(
        n16523) );
  NAND4_X1 U19705 ( .A1(n16526), .A2(n16525), .A3(n16524), .A4(n16523), .ZN(
        P3_U2644) );
  INV_X1 U19706 ( .A(n16527), .ZN(n16539) );
  AOI21_X1 U19707 ( .B1(n16807), .B2(n16528), .A(P3_REIP_REG_26__SCAN_IN), 
        .ZN(n16538) );
  AOI22_X1 U19708 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16821), .B1(
        n16838), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16537) );
  AOI211_X1 U19709 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16530), .A(n16529), .B(
        n16827), .ZN(n16535) );
  INV_X1 U19710 ( .A(n16531), .ZN(n16532) );
  AOI211_X1 U19711 ( .C1(n17543), .C2(n16533), .A(n16532), .B(n18717), .ZN(
        n16534) );
  NOR2_X1 U19712 ( .A1(n16535), .A2(n16534), .ZN(n16536) );
  OAI211_X1 U19713 ( .C1(n16539), .C2(n16538), .A(n16537), .B(n16536), .ZN(
        P3_U2645) );
  OR2_X1 U19714 ( .A1(n16827), .A2(n16540), .ZN(n16553) );
  AOI21_X1 U19715 ( .B1(n16837), .B2(n16540), .A(n16838), .ZN(n16550) );
  AOI211_X1 U19716 ( .C1(n17554), .C2(n16542), .A(n16541), .B(n18717), .ZN(
        n16548) );
  NOR2_X1 U19717 ( .A1(n16825), .A2(n16543), .ZN(n16546) );
  INV_X1 U19718 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18779) );
  OAI21_X1 U19719 ( .B1(n16564), .B2(n16825), .A(n16783), .ZN(n16560) );
  AOI21_X1 U19720 ( .B1(n16807), .B2(n18779), .A(n16560), .ZN(n16544) );
  INV_X1 U19721 ( .A(n16544), .ZN(n16545) );
  MUX2_X1 U19722 ( .A(n16546), .B(n16545), .S(P3_REIP_REG_25__SCAN_IN), .Z(
        n16547) );
  AOI211_X1 U19723 ( .C1(n16821), .C2(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n16548), .B(n16547), .ZN(n16549) );
  OAI221_X1 U19724 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n16553), .C1(n16551), 
        .C2(n16550), .A(n16549), .ZN(P3_U2646) );
  NOR2_X1 U19725 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16825), .ZN(n16552) );
  AOI22_X1 U19726 ( .A1(n16838), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16564), 
        .B2(n16552), .ZN(n16559) );
  AOI21_X1 U19727 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16569), .A(n16553), .ZN(
        n16557) );
  AOI211_X1 U19728 ( .C1(n17568), .C2(n16555), .A(n16554), .B(n18717), .ZN(
        n16556) );
  AOI211_X1 U19729 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16560), .A(n16557), 
        .B(n16556), .ZN(n16558) );
  OAI211_X1 U19730 ( .C1(n17572), .C2(n16804), .A(n16559), .B(n16558), .ZN(
        P3_U2647) );
  INV_X1 U19731 ( .A(n16560), .ZN(n16573) );
  INV_X1 U19732 ( .A(n16561), .ZN(n16562) );
  AOI211_X1 U19733 ( .C1(n17588), .C2(n16563), .A(n16562), .B(n18717), .ZN(
        n16568) );
  OR2_X1 U19734 ( .A1(n16825), .A2(n16564), .ZN(n16565) );
  OAI22_X1 U19735 ( .A1(n17591), .A2(n16804), .B1(n16566), .B2(n16565), .ZN(
        n16567) );
  AOI211_X1 U19736 ( .C1(P3_EBX_REG_23__SCAN_IN), .C2(n16838), .A(n16568), .B(
        n16567), .ZN(n16572) );
  OAI211_X1 U19737 ( .C1(n16574), .C2(n16570), .A(n16837), .B(n16569), .ZN(
        n16571) );
  OAI211_X1 U19738 ( .C1(n16573), .C2(n18777), .A(n16572), .B(n16571), .ZN(
        P3_U2648) );
  AOI221_X1 U19739 ( .B1(n18773), .B2(n16807), .C1(n16584), .C2(n16807), .A(
        n16834), .ZN(n16583) );
  INV_X1 U19740 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18775) );
  AOI22_X1 U19741 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n16821), .B1(
        n16838), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n16582) );
  NOR2_X1 U19742 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16825), .ZN(n16579) );
  AOI211_X1 U19743 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16588), .A(n16574), .B(
        n16827), .ZN(n16578) );
  AOI211_X1 U19744 ( .C1(n17605), .C2(n16576), .A(n16575), .B(n18717), .ZN(
        n16577) );
  AOI211_X1 U19745 ( .C1(n16580), .C2(n16579), .A(n16578), .B(n16577), .ZN(
        n16581) );
  OAI211_X1 U19746 ( .C1(n16583), .C2(n18775), .A(n16582), .B(n16581), .ZN(
        P3_U2649) );
  INV_X1 U19747 ( .A(n16584), .ZN(n16593) );
  NOR2_X1 U19748 ( .A1(n16825), .A2(n16593), .ZN(n16602) );
  NOR2_X1 U19749 ( .A1(n16834), .A2(n16602), .ZN(n16605) );
  INV_X1 U19750 ( .A(n16605), .ZN(n16592) );
  INV_X1 U19751 ( .A(n16585), .ZN(n16586) );
  AOI211_X1 U19752 ( .C1(n17613), .C2(n16587), .A(n16586), .B(n18717), .ZN(
        n16591) );
  OAI211_X1 U19753 ( .C1(n16598), .C2(n17012), .A(n16837), .B(n16588), .ZN(
        n16589) );
  OAI21_X1 U19754 ( .B1(n17012), .B2(n16824), .A(n16589), .ZN(n16590) );
  AOI211_X1 U19755 ( .C1(P3_REIP_REG_21__SCAN_IN), .C2(n16592), .A(n16591), 
        .B(n16590), .ZN(n16595) );
  NAND3_X1 U19756 ( .A1(n16807), .A2(n16593), .A3(n18773), .ZN(n16594) );
  OAI211_X1 U19757 ( .C1(n16804), .C2(n17617), .A(n16595), .B(n16594), .ZN(
        P3_U2650) );
  INV_X1 U19758 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18771) );
  AOI22_X1 U19759 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n16821), .B1(
        n16838), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n16604) );
  AOI211_X1 U19760 ( .C1(n17633), .C2(n16597), .A(n16596), .B(n18717), .ZN(
        n16600) );
  AOI211_X1 U19761 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16612), .A(n16598), .B(
        n16827), .ZN(n16599) );
  AOI211_X1 U19762 ( .C1(n16602), .C2(n16601), .A(n16600), .B(n16599), .ZN(
        n16603) );
  OAI211_X1 U19763 ( .C1(n16605), .C2(n18771), .A(n16604), .B(n16603), .ZN(
        P3_U2651) );
  NAND2_X1 U19764 ( .A1(n16807), .A2(n18769), .ZN(n16616) );
  INV_X1 U19765 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18767) );
  AND3_X1 U19766 ( .A1(n18767), .A2(n16807), .A3(n16606), .ZN(n16619) );
  OAI21_X1 U19767 ( .B1(n16606), .B2(n16825), .A(n16783), .ZN(n16633) );
  INV_X1 U19768 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17655) );
  NOR2_X1 U19769 ( .A1(n17655), .A2(n16628), .ZN(n16620) );
  OAI21_X1 U19770 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16620), .A(
        n16607), .ZN(n17644) );
  OAI21_X1 U19771 ( .B1(n16620), .B2(n16820), .A(n16645), .ZN(n16608) );
  XOR2_X1 U19772 ( .A(n17644), .B(n16608), .Z(n16610) );
  AOI22_X1 U19773 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n16821), .B1(
        n16838), .B2(P3_EBX_REG_19__SCAN_IN), .ZN(n16609) );
  OAI211_X1 U19774 ( .C1(n18717), .C2(n16610), .A(n16609), .B(n18193), .ZN(
        n16611) );
  AOI221_X1 U19775 ( .B1(n16619), .B2(P3_REIP_REG_19__SCAN_IN), .C1(n16633), 
        .C2(P3_REIP_REG_19__SCAN_IN), .A(n16611), .ZN(n16614) );
  OAI211_X1 U19776 ( .C1(n16617), .C2(n20786), .A(n16837), .B(n16612), .ZN(
        n16613) );
  OAI211_X1 U19777 ( .C1(n16616), .C2(n16615), .A(n16614), .B(n16613), .ZN(
        P3_U2652) );
  AOI211_X1 U19778 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16635), .A(n16617), .B(
        n16827), .ZN(n16618) );
  AOI21_X1 U19779 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n16838), .A(n16618), .ZN(
        n16626) );
  AOI211_X1 U19780 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(n16821), .A(
        n9726), .B(n16619), .ZN(n16625) );
  AOI21_X1 U19781 ( .B1(n17655), .B2(n16628), .A(n16620), .ZN(n16621) );
  INV_X1 U19782 ( .A(n16621), .ZN(n17652) );
  OAI21_X1 U19783 ( .B1(n17639), .B2(n16820), .A(n16645), .ZN(n16622) );
  XNOR2_X1 U19784 ( .A(n17652), .B(n16622), .ZN(n16623) );
  AOI22_X1 U19785 ( .A1(n16823), .A2(n16623), .B1(P3_REIP_REG_18__SCAN_IN), 
        .B2(n16633), .ZN(n16624) );
  NAND3_X1 U19786 ( .A1(n16626), .A2(n16625), .A3(n16624), .ZN(P3_U2653) );
  AOI22_X1 U19787 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16821), .B1(
        n16838), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n16638) );
  NAND3_X1 U19788 ( .A1(n16807), .A2(P3_REIP_REG_14__SCAN_IN), .A3(n16664), 
        .ZN(n16652) );
  NOR2_X1 U19789 ( .A1(n16627), .A2(n16652), .ZN(n16634) );
  AND2_X1 U19790 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17661), .ZN(
        n16643) );
  OAI21_X1 U19791 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16643), .A(
        n16628), .ZN(n17666) );
  NOR2_X1 U19792 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17870), .ZN(
        n16816) );
  AOI21_X1 U19793 ( .B1(n17661), .B2(n16816), .A(n16820), .ZN(n16629) );
  INV_X1 U19794 ( .A(n16629), .ZN(n16631) );
  OAI21_X1 U19795 ( .B1(n17666), .B2(n16631), .A(n16823), .ZN(n16630) );
  AOI21_X1 U19796 ( .B1(n17666), .B2(n16631), .A(n16630), .ZN(n16632) );
  AOI221_X1 U19797 ( .B1(n16634), .B2(n18765), .C1(n16633), .C2(
        P3_REIP_REG_17__SCAN_IN), .A(n16632), .ZN(n16637) );
  OAI211_X1 U19798 ( .C1(n16639), .C2(n20806), .A(n16837), .B(n16635), .ZN(
        n16636) );
  NAND4_X1 U19799 ( .A1(n16638), .A2(n16637), .A3(n18193), .A4(n16636), .ZN(
        P3_U2654) );
  INV_X1 U19800 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16650) );
  AOI211_X1 U19801 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16655), .A(n16639), .B(
        n16827), .ZN(n16640) );
  AOI211_X1 U19802 ( .C1(n16838), .C2(P3_EBX_REG_16__SCAN_IN), .A(n9726), .B(
        n16640), .ZN(n16649) );
  NOR2_X1 U19803 ( .A1(n16834), .A2(n16641), .ZN(n16667) );
  NAND2_X1 U19804 ( .A1(n16783), .A2(n16825), .ZN(n16836) );
  INV_X1 U19805 ( .A(n16836), .ZN(n16642) );
  AOI21_X1 U19806 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16667), .A(n16642), 
        .ZN(n16653) );
  INV_X1 U19807 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18761) );
  NOR2_X1 U19808 ( .A1(n18761), .A2(n16652), .ZN(n16647) );
  INV_X1 U19809 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18763) );
  INV_X1 U19810 ( .A(n16645), .ZN(n16660) );
  AOI21_X1 U19811 ( .B1(n16650), .B2(n16651), .A(n16643), .ZN(n17678) );
  INV_X1 U19812 ( .A(n17678), .ZN(n16644) );
  AOI221_X1 U19813 ( .B1(n16660), .B2(n17678), .C1(n16645), .C2(n16644), .A(
        n18717), .ZN(n16646) );
  AOI221_X1 U19814 ( .B1(n16653), .B2(P3_REIP_REG_16__SCAN_IN), .C1(n16647), 
        .C2(n18763), .A(n16646), .ZN(n16648) );
  OAI211_X1 U19815 ( .C1(n16650), .C2(n16804), .A(n16649), .B(n16648), .ZN(
        P3_U2655) );
  OAI21_X1 U19816 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17677), .A(
        n16651), .ZN(n17687) );
  INV_X1 U19817 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16833) );
  OAI21_X1 U19818 ( .B1(n16820), .B2(n16833), .A(n16823), .ZN(n16832) );
  AOI211_X1 U19819 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n16758), .A(
        n17687), .B(n16832), .ZN(n16659) );
  INV_X1 U19820 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17690) );
  INV_X1 U19821 ( .A(n16652), .ZN(n16654) );
  OAI21_X1 U19822 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16654), .A(n16653), 
        .ZN(n16657) );
  OAI211_X1 U19823 ( .C1(n16663), .C2(n20783), .A(n16837), .B(n16655), .ZN(
        n16656) );
  OAI211_X1 U19824 ( .C1(n16804), .C2(n17690), .A(n16657), .B(n16656), .ZN(
        n16658) );
  AOI211_X1 U19825 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n16838), .A(n16659), .B(
        n16658), .ZN(n16662) );
  NAND3_X1 U19826 ( .A1(n16660), .A2(n16823), .A3(n17687), .ZN(n16661) );
  NAND3_X1 U19827 ( .A1(n16662), .A2(n18193), .A3(n16661), .ZN(P3_U2656) );
  INV_X1 U19828 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n17111) );
  AOI211_X1 U19829 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16679), .A(n16663), .B(
        n16827), .ZN(n16669) );
  AOI22_X1 U19830 ( .A1(n16807), .A2(n16664), .B1(P3_REIP_REG_14__SCAN_IN), 
        .B2(n16836), .ZN(n16666) );
  AOI21_X1 U19831 ( .B1(n9987), .B2(n16673), .A(n17677), .ZN(n17704) );
  OAI21_X1 U19832 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16673), .A(
        n16758), .ZN(n16671) );
  XOR2_X1 U19833 ( .A(n17704), .B(n16671), .Z(n16665) );
  OAI22_X1 U19834 ( .A1(n16667), .A2(n16666), .B1(n18717), .B2(n16665), .ZN(
        n16668) );
  AOI211_X1 U19835 ( .C1(n16821), .C2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16669), .B(n16668), .ZN(n16670) );
  OAI211_X1 U19836 ( .C1(n16824), .C2(n17111), .A(n16670), .B(n18193), .ZN(
        P3_U2657) );
  AOI22_X1 U19837 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n16821), .B1(
        n16838), .B2(P3_EBX_REG_13__SCAN_IN), .ZN(n16683) );
  NOR2_X1 U19838 ( .A1(n18717), .A2(n16671), .ZN(n16677) );
  INV_X1 U19839 ( .A(n16672), .ZN(n16689) );
  INV_X1 U19840 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16776) );
  NAND2_X1 U19841 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17812), .ZN(
        n16777) );
  NOR2_X1 U19842 ( .A1(n16776), .A2(n16777), .ZN(n16767) );
  NAND2_X1 U19843 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16767), .ZN(
        n16754) );
  NOR2_X1 U19844 ( .A1(n16689), .A2(n16754), .ZN(n17712) );
  NAND2_X1 U19845 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17712), .ZN(
        n16688) );
  INV_X1 U19846 ( .A(n16688), .ZN(n16674) );
  OAI21_X1 U19847 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16674), .A(
        n16673), .ZN(n17718) );
  NOR3_X1 U19848 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16825), .A3(n16675), 
        .ZN(n16676) );
  AOI211_X1 U19849 ( .C1(n16677), .C2(n17718), .A(n9726), .B(n16676), .ZN(
        n16682) );
  NOR2_X1 U19850 ( .A1(P3_REIP_REG_12__SCAN_IN), .A2(n16825), .ZN(n16686) );
  OAI21_X1 U19851 ( .B1(n16687), .B2(n16825), .A(n16783), .ZN(n16705) );
  NAND2_X1 U19852 ( .A1(n16823), .A2(n16820), .ZN(n16819) );
  AOI211_X1 U19853 ( .C1(n16688), .C2(n16819), .A(n17718), .B(n16832), .ZN(
        n16678) );
  AOI221_X1 U19854 ( .B1(n16686), .B2(P3_REIP_REG_13__SCAN_IN), .C1(n16705), 
        .C2(P3_REIP_REG_13__SCAN_IN), .A(n16678), .ZN(n16681) );
  OAI211_X1 U19855 ( .C1(n16684), .C2(n21008), .A(n16837), .B(n16679), .ZN(
        n16680) );
  NAND4_X1 U19856 ( .A1(n16683), .A2(n16682), .A3(n16681), .A4(n16680), .ZN(
        P3_U2658) );
  AOI22_X1 U19857 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16821), .B1(
        n16838), .B2(P3_EBX_REG_12__SCAN_IN), .ZN(n16694) );
  AOI211_X1 U19858 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16699), .A(n16684), .B(
        n16827), .ZN(n16685) );
  AOI211_X1 U19859 ( .C1(n16687), .C2(n16686), .A(n9726), .B(n16685), .ZN(
        n16693) );
  OAI21_X1 U19860 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n17712), .A(
        n16688), .ZN(n17729) );
  NAND2_X1 U19861 ( .A1(n17777), .A2(n16816), .ZN(n16757) );
  OAI21_X1 U19862 ( .B1(n16689), .B2(n16757), .A(n16758), .ZN(n16690) );
  XOR2_X1 U19863 ( .A(n17729), .B(n16690), .Z(n16691) );
  AOI22_X1 U19864 ( .A1(n16823), .A2(n16691), .B1(P3_REIP_REG_12__SCAN_IN), 
        .B2(n16705), .ZN(n16692) );
  NAND3_X1 U19865 ( .A1(n16694), .A2(n16693), .A3(n16692), .ZN(P3_U2659) );
  NOR2_X1 U19866 ( .A1(n16825), .A2(n16731), .ZN(n16710) );
  INV_X1 U19867 ( .A(n16710), .ZN(n16726) );
  OAI21_X1 U19868 ( .B1(n16709), .B2(n16726), .A(n18753), .ZN(n16704) );
  NAND2_X1 U19869 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16695) );
  INV_X1 U19870 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17791) );
  NOR2_X1 U19871 ( .A1(n17791), .A2(n16754), .ZN(n16744) );
  NAND2_X1 U19872 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16744), .ZN(
        n16736) );
  OR2_X1 U19873 ( .A1(n16695), .A2(n16736), .ZN(n16714) );
  AOI21_X1 U19874 ( .B1(n16702), .B2(n16714), .A(n17712), .ZN(n16696) );
  INV_X1 U19875 ( .A(n16696), .ZN(n17745) );
  OAI21_X1 U19876 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16714), .A(
        n16758), .ZN(n16698) );
  AOI21_X1 U19877 ( .B1(n17745), .B2(n16698), .A(n18717), .ZN(n16697) );
  OAI21_X1 U19878 ( .B1(n17745), .B2(n16698), .A(n16697), .ZN(n16701) );
  OAI211_X1 U19879 ( .C1(n16708), .C2(n16707), .A(n16837), .B(n16699), .ZN(
        n16700) );
  OAI211_X1 U19880 ( .C1(n16804), .C2(n16702), .A(n16701), .B(n16700), .ZN(
        n16703) );
  AOI21_X1 U19881 ( .B1(n16705), .B2(n16704), .A(n16703), .ZN(n16706) );
  OAI211_X1 U19882 ( .C1(n16824), .C2(n16707), .A(n16706), .B(n18193), .ZN(
        P3_U2660) );
  AOI21_X1 U19883 ( .B1(n16807), .B2(n16731), .A(n16834), .ZN(n16743) );
  INV_X1 U19884 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18752) );
  AOI211_X1 U19885 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16720), .A(n16708), .B(
        n16827), .ZN(n16713) );
  INV_X1 U19886 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n17144) );
  OAI211_X1 U19887 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(P3_REIP_REG_9__SCAN_IN), 
        .A(n16710), .B(n16709), .ZN(n16711) );
  OAI211_X1 U19888 ( .C1(n16824), .C2(n17144), .A(n18193), .B(n16711), .ZN(
        n16712) );
  AOI211_X1 U19889 ( .C1(n16821), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n16713), .B(n16712), .ZN(n16719) );
  INV_X1 U19890 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n17751) );
  NOR2_X1 U19891 ( .A1(n17751), .A2(n16736), .ZN(n16715) );
  OAI21_X1 U19892 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16715), .A(
        n16714), .ZN(n17752) );
  INV_X1 U19893 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16738) );
  NOR3_X1 U19894 ( .A1(n17791), .A2(n16738), .A3(n16757), .ZN(n16724) );
  NAND2_X1 U19895 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16724), .ZN(
        n16723) );
  NAND2_X1 U19896 ( .A1(n16758), .A2(n16723), .ZN(n16717) );
  AOI21_X1 U19897 ( .B1(n17752), .B2(n16717), .A(n18717), .ZN(n16716) );
  OAI21_X1 U19898 ( .B1(n17752), .B2(n16717), .A(n16716), .ZN(n16718) );
  OAI211_X1 U19899 ( .C1(n16743), .C2(n18752), .A(n16719), .B(n16718), .ZN(
        P3_U2661) );
  INV_X1 U19900 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18751) );
  OAI211_X1 U19901 ( .C1(n16732), .C2(n17143), .A(n16837), .B(n16720), .ZN(
        n16721) );
  OAI21_X1 U19902 ( .B1(n17143), .B2(n16824), .A(n16721), .ZN(n16729) );
  INV_X1 U19903 ( .A(n16736), .ZN(n16722) );
  AOI22_X1 U19904 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16736), .B1(
        n16722), .B2(n17751), .ZN(n17766) );
  OAI211_X1 U19905 ( .C1(n16724), .C2(n17766), .A(n16758), .B(n16723), .ZN(
        n16725) );
  OAI22_X1 U19906 ( .A1(n17751), .A2(n16804), .B1(n18717), .B2(n16725), .ZN(
        n16728) );
  OAI22_X1 U19907 ( .A1(P3_REIP_REG_9__SCAN_IN), .A2(n16726), .B1(n16819), 
        .B2(n17766), .ZN(n16727) );
  NOR4_X1 U19908 ( .A1(n9726), .A2(n16729), .A3(n16728), .A4(n16727), .ZN(
        n16730) );
  OAI21_X1 U19909 ( .B1(n16743), .B2(n18751), .A(n16730), .ZN(P3_U2662) );
  INV_X1 U19910 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n20834) );
  AND2_X1 U19911 ( .A1(n16731), .A2(n16807), .ZN(n16734) );
  AOI211_X1 U19912 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16746), .A(n16732), .B(
        n16827), .ZN(n16733) );
  AOI211_X1 U19913 ( .C1(n16735), .C2(n16734), .A(n9726), .B(n16733), .ZN(
        n16742) );
  OAI21_X1 U19914 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16744), .A(
        n16736), .ZN(n17779) );
  OAI21_X1 U19915 ( .B1(n17791), .B2(n16757), .A(n16758), .ZN(n16737) );
  XOR2_X1 U19916 ( .A(n17779), .B(n16737), .Z(n16740) );
  OAI22_X1 U19917 ( .A1(n16738), .A2(n16804), .B1(n16824), .B2(n17204), .ZN(
        n16739) );
  AOI21_X1 U19918 ( .B1(n16823), .B2(n16740), .A(n16739), .ZN(n16741) );
  OAI211_X1 U19919 ( .C1(n16743), .C2(n20834), .A(n16742), .B(n16741), .ZN(
        P3_U2663) );
  NAND2_X1 U19920 ( .A1(n16758), .A2(n16757), .ZN(n16745) );
  AOI21_X1 U19921 ( .B1(n17791), .B2(n16754), .A(n16744), .ZN(n17797) );
  XOR2_X1 U19922 ( .A(n16745), .B(n17797), .Z(n16753) );
  OAI211_X1 U19923 ( .C1(n16756), .C2(n17210), .A(n16837), .B(n16746), .ZN(
        n16747) );
  OAI211_X1 U19924 ( .C1(n16824), .C2(n17210), .A(n18193), .B(n16747), .ZN(
        n16751) );
  NAND3_X1 U19925 ( .A1(n16807), .A2(P3_REIP_REG_5__SCAN_IN), .A3(n16766), 
        .ZN(n16765) );
  XOR2_X1 U19926 ( .A(P3_REIP_REG_7__SCAN_IN), .B(n18747), .Z(n16749) );
  AOI21_X1 U19927 ( .B1(n16807), .B2(n16748), .A(n16834), .ZN(n16770) );
  OAI22_X1 U19928 ( .A1(n16765), .A2(n16749), .B1(n18749), .B2(n16770), .ZN(
        n16750) );
  AOI211_X1 U19929 ( .C1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n16821), .A(
        n16751), .B(n16750), .ZN(n16752) );
  OAI21_X1 U19930 ( .B1(n16753), .B2(n18717), .A(n16752), .ZN(P3_U2664) );
  INV_X1 U19931 ( .A(n16767), .ZN(n16755) );
  OAI21_X1 U19932 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16767), .A(
        n16754), .ZN(n17806) );
  AOI211_X1 U19933 ( .C1(n16758), .C2(n16755), .A(n17806), .B(n16832), .ZN(
        n16763) );
  AOI211_X1 U19934 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16772), .A(n16756), .B(
        n16827), .ZN(n16762) );
  AOI22_X1 U19935 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16821), .B1(
        n16838), .B2(P3_EBX_REG_6__SCAN_IN), .ZN(n16760) );
  NAND4_X1 U19936 ( .A1(n16823), .A2(n16758), .A3(n17806), .A4(n16757), .ZN(
        n16759) );
  NAND3_X1 U19937 ( .A1(n16760), .A2(n18193), .A3(n16759), .ZN(n16761) );
  NOR3_X1 U19938 ( .A1(n16763), .A2(n16762), .A3(n16761), .ZN(n16764) );
  OAI221_X1 U19939 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n16765), .C1(n18747), 
        .C2(n16770), .A(n16764), .ZN(P3_U2665) );
  AOI21_X1 U19940 ( .B1(n16807), .B2(n16766), .A(P3_REIP_REG_5__SCAN_IN), .ZN(
        n16769) );
  AOI21_X1 U19941 ( .B1(n16776), .B2(n16777), .A(n16767), .ZN(n17823) );
  AOI21_X1 U19942 ( .B1(n17812), .B2(n16816), .A(n16820), .ZN(n16778) );
  XNOR2_X1 U19943 ( .A(n17823), .B(n16778), .ZN(n16768) );
  OAI22_X1 U19944 ( .A1(n16770), .A2(n16769), .B1(n18717), .B2(n16768), .ZN(
        n16771) );
  AOI211_X1 U19945 ( .C1(n16838), .C2(P3_EBX_REG_5__SCAN_IN), .A(n9726), .B(
        n16771), .ZN(n16775) );
  OAI211_X1 U19946 ( .C1(n16784), .C2(n16773), .A(n16837), .B(n16772), .ZN(
        n16774) );
  OAI211_X1 U19947 ( .C1(n16804), .C2(n16776), .A(n16775), .B(n16774), .ZN(
        P3_U2666) );
  NOR2_X1 U19948 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17828), .ZN(
        n17839) );
  NOR2_X1 U19949 ( .A1(n17870), .A2(n17828), .ZN(n16792) );
  OAI21_X1 U19950 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16792), .A(
        n16777), .ZN(n17836) );
  AOI22_X1 U19951 ( .A1(n16816), .A2(n17839), .B1(n16778), .B2(n17836), .ZN(
        n16790) );
  NOR3_X1 U19952 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16825), .A3(n16782), .ZN(
        n16781) );
  OAI22_X1 U19953 ( .A1(n16824), .A2(n16779), .B1(n17836), .B2(n16819), .ZN(
        n16780) );
  AOI211_X1 U19954 ( .C1(n16821), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n16781), .B(n16780), .ZN(n16789) );
  NAND2_X1 U19955 ( .A1(n16807), .A2(n16782), .ZN(n16797) );
  NAND2_X1 U19956 ( .A1(n16783), .A2(n16797), .ZN(n16799) );
  AOI211_X1 U19957 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16800), .A(n16784), .B(
        n16827), .ZN(n16787) );
  NOR2_X1 U19958 ( .A1(n18853), .A2(n18847), .ZN(n18870) );
  INV_X1 U19959 ( .A(n18870), .ZN(n16841) );
  OAI221_X1 U19960 ( .B1(n16841), .B2(n10128), .C1(n16841), .C2(n16785), .A(
        n18193), .ZN(n16786) );
  AOI211_X1 U19961 ( .C1(P3_REIP_REG_4__SCAN_IN), .C2(n16799), .A(n16787), .B(
        n16786), .ZN(n16788) );
  OAI211_X1 U19962 ( .C1(n16790), .C2(n18717), .A(n16789), .B(n16788), .ZN(
        P3_U2667) );
  INV_X1 U19963 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17848) );
  NAND2_X1 U19964 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16806) );
  NAND2_X1 U19965 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18666) );
  NOR2_X1 U19966 ( .A1(n21023), .A2(n18666), .ZN(n18649) );
  OAI21_X1 U19967 ( .B1(n18649), .B2(n18812), .A(n16791), .ZN(n18809) );
  AOI22_X1 U19968 ( .A1(n16838), .A2(P3_EBX_REG_3__SCAN_IN), .B1(n18870), .B2(
        n18809), .ZN(n16796) );
  INV_X1 U19969 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17863) );
  NOR2_X1 U19970 ( .A1(n17870), .A2(n17863), .ZN(n16793) );
  INV_X1 U19971 ( .A(n16793), .ZN(n16805) );
  AOI21_X1 U19972 ( .B1(n17848), .B2(n16805), .A(n16792), .ZN(n17852) );
  AOI21_X1 U19973 ( .B1(n16793), .B2(n16833), .A(n16820), .ZN(n16815) );
  AOI21_X1 U19974 ( .B1(n17852), .B2(n16815), .A(n18717), .ZN(n16794) );
  OAI21_X1 U19975 ( .B1(n17852), .B2(n16815), .A(n16794), .ZN(n16795) );
  OAI211_X1 U19976 ( .C1(n16797), .C2(n16806), .A(n16796), .B(n16795), .ZN(
        n16798) );
  AOI21_X1 U19977 ( .B1(P3_REIP_REG_3__SCAN_IN), .B2(n16799), .A(n16798), .ZN(
        n16803) );
  OAI211_X1 U19978 ( .C1(n16808), .C2(n16801), .A(n16837), .B(n16800), .ZN(
        n16802) );
  OAI211_X1 U19979 ( .C1(n16804), .C2(n17848), .A(n16803), .B(n16802), .ZN(
        P3_U2668) );
  OAI21_X1 U19980 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16805), .ZN(n17860) );
  AOI21_X1 U19981 ( .B1(n18820), .B2(n18665), .A(n18649), .ZN(n18816) );
  AOI22_X1 U19982 ( .A1(n16834), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n18816), 
        .B2(n18870), .ZN(n16814) );
  AOI22_X1 U19983 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n16821), .B1(
        n16838), .B2(P3_EBX_REG_2__SCAN_IN), .ZN(n16813) );
  OAI211_X1 U19984 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16807), .B(n16806), .ZN(n16812) );
  OR2_X1 U19985 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), .ZN(
        n16809) );
  AOI211_X1 U19986 ( .C1(n16809), .C2(P3_EBX_REG_2__SCAN_IN), .A(n16827), .B(
        n16808), .ZN(n16810) );
  INV_X1 U19987 ( .A(n16810), .ZN(n16811) );
  AND4_X1 U19988 ( .A1(n16814), .A2(n16813), .A3(n16812), .A4(n16811), .ZN(
        n16818) );
  OAI211_X1 U19989 ( .C1(n16816), .C2(n17860), .A(n16823), .B(n16815), .ZN(
        n16817) );
  OAI211_X1 U19990 ( .C1(n16819), .C2(n17860), .A(n16818), .B(n16817), .ZN(
        P3_U2669) );
  NOR2_X1 U19991 ( .A1(n16820), .A2(n16833), .ZN(n16822) );
  AOI21_X1 U19992 ( .B1(n16823), .B2(n16822), .A(n16821), .ZN(n16831) );
  INV_X1 U19993 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n20848) );
  OAI22_X1 U19994 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16825), .B1(n16824), 
        .B2(n20848), .ZN(n16829) );
  NAND2_X1 U19995 ( .A1(P3_EBX_REG_1__SCAN_IN), .A2(P3_EBX_REG_0__SCAN_IN), 
        .ZN(n17228) );
  OAI21_X1 U19996 ( .B1(P3_EBX_REG_1__SCAN_IN), .B2(P3_EBX_REG_0__SCAN_IN), 
        .A(n17228), .ZN(n17236) );
  NAND2_X1 U19997 ( .A1(n16826), .A2(n18665), .ZN(n18821) );
  OAI22_X1 U19998 ( .A1(n16827), .A2(n17236), .B1(n18821), .B2(n16841), .ZN(
        n16828) );
  AOI211_X1 U19999 ( .C1(n16834), .C2(P3_REIP_REG_1__SCAN_IN), .A(n16829), .B(
        n16828), .ZN(n16830) );
  OAI221_X1 U20000 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16832), .C1(
        n17870), .C2(n16831), .A(n16830), .ZN(P3_U2670) );
  NOR3_X1 U20001 ( .A1(n18866), .A2(n16834), .A3(n16833), .ZN(n16835) );
  AOI21_X1 U20002 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n16836), .A(n16835), .ZN(
        n16840) );
  OAI21_X1 U20003 ( .B1(n16838), .B2(n16837), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n16839) );
  OAI211_X1 U20004 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n16841), .A(
        n16840), .B(n16839), .ZN(P3_U2671) );
  INV_X1 U20005 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16843) );
  NAND4_X1 U20006 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(P3_EBX_REG_13__SCAN_IN), 
        .A3(P3_EBX_REG_12__SCAN_IN), .A4(n17115), .ZN(n17095) );
  NAND4_X1 U20007 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(P3_EBX_REG_17__SCAN_IN), 
        .A3(P3_EBX_REG_16__SCAN_IN), .A4(n17077), .ZN(n17051) );
  INV_X1 U20008 ( .A(n17051), .ZN(n17039) );
  NAND2_X1 U20009 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n17039), .ZN(n17038) );
  NOR2_X1 U20010 ( .A1(n16843), .A2(n17038), .ZN(n17011) );
  NAND2_X1 U20011 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .ZN(n16846) );
  NAND2_X1 U20012 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(P3_EBX_REG_24__SCAN_IN), 
        .ZN(n16845) );
  NAND2_X1 U20013 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n16844) );
  NOR4_X1 U20014 ( .A1(n16847), .A2(n16846), .A3(n16845), .A4(n16844), .ZN(
        n16848) );
  NAND4_X1 U20015 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_21__SCAN_IN), 
        .A3(n17011), .A4(n16848), .ZN(n16851) );
  NOR2_X1 U20016 ( .A1(n16852), .A2(n16851), .ZN(n16952) );
  NAND2_X1 U20017 ( .A1(n17233), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16850) );
  NAND2_X1 U20018 ( .A1(n16952), .A2(n18245), .ZN(n16849) );
  OAI22_X1 U20019 ( .A1(n16952), .A2(n16850), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16849), .ZN(P3_U2672) );
  NAND2_X1 U20020 ( .A1(n16852), .A2(n16851), .ZN(n16853) );
  NAND2_X1 U20021 ( .A1(n16853), .A2(n17233), .ZN(n16951) );
  AOI22_X1 U20022 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16857) );
  AOI22_X1 U20023 ( .A1(n17188), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12832), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16856) );
  AOI22_X1 U20024 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16855) );
  AOI22_X1 U20025 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16854) );
  NAND4_X1 U20026 ( .A1(n16857), .A2(n16856), .A3(n16855), .A4(n16854), .ZN(
        n16863) );
  AOI22_X1 U20027 ( .A1(n16910), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16861) );
  AOI22_X1 U20028 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16860) );
  AOI22_X1 U20029 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17193), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16859) );
  AOI22_X1 U20030 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n16876), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16858) );
  NAND4_X1 U20031 ( .A1(n16861), .A2(n16860), .A3(n16859), .A4(n16858), .ZN(
        n16862) );
  NOR2_X1 U20032 ( .A1(n16863), .A2(n16862), .ZN(n16954) );
  AOI22_X1 U20033 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12832), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16868) );
  AOI22_X1 U20034 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n16867) );
  AOI22_X1 U20035 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n16866) );
  AOI22_X1 U20036 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16865) );
  NAND4_X1 U20037 ( .A1(n16868), .A2(n16867), .A3(n16866), .A4(n16865), .ZN(
        n16875) );
  AOI22_X1 U20038 ( .A1(n16891), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n16873) );
  AOI22_X1 U20039 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16872) );
  AOI22_X1 U20040 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n16869), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16871) );
  AOI22_X1 U20041 ( .A1(n17084), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n16876), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n16870) );
  NAND4_X1 U20042 ( .A1(n16873), .A2(n16872), .A3(n16871), .A4(n16870), .ZN(
        n16874) );
  NOR2_X1 U20043 ( .A1(n16875), .A2(n16874), .ZN(n16964) );
  AOI22_X1 U20044 ( .A1(n17165), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16880) );
  AOI22_X1 U20045 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16879) );
  AOI22_X1 U20046 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17193), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n16878) );
  AOI22_X1 U20047 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n16876), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n16877) );
  NAND4_X1 U20048 ( .A1(n16880), .A2(n16879), .A3(n16878), .A4(n16877), .ZN(
        n16886) );
  AOI22_X1 U20049 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n16884) );
  AOI22_X1 U20050 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n16883) );
  AOI22_X1 U20051 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16882) );
  AOI22_X1 U20052 ( .A1(n16891), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n16881) );
  NAND4_X1 U20053 ( .A1(n16884), .A2(n16883), .A3(n16882), .A4(n16881), .ZN(
        n16885) );
  NOR2_X1 U20054 ( .A1(n16886), .A2(n16885), .ZN(n16973) );
  AOI22_X1 U20055 ( .A1(n17165), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17193), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n16890) );
  AOI22_X1 U20056 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n16889) );
  AOI22_X1 U20057 ( .A1(n17084), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16888) );
  AOI22_X1 U20058 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16887) );
  NAND4_X1 U20059 ( .A1(n16890), .A2(n16889), .A3(n16888), .A4(n16887), .ZN(
        n16897) );
  AOI22_X1 U20060 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n16895) );
  AOI22_X1 U20061 ( .A1(n17190), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n16894) );
  AOI22_X1 U20062 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17057), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n16893) );
  AOI22_X1 U20063 ( .A1(n16891), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n16892) );
  NAND4_X1 U20064 ( .A1(n16895), .A2(n16894), .A3(n16893), .A4(n16892), .ZN(
        n16896) );
  NOR2_X1 U20065 ( .A1(n16897), .A2(n16896), .ZN(n16982) );
  AOI22_X1 U20066 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12832), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16901) );
  AOI22_X1 U20067 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16900) );
  AOI22_X1 U20068 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16899) );
  AOI22_X1 U20069 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16898) );
  NAND4_X1 U20070 ( .A1(n16901), .A2(n16900), .A3(n16899), .A4(n16898), .ZN(
        n16907) );
  AOI22_X1 U20071 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n16905) );
  AOI22_X1 U20072 ( .A1(n17084), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16904) );
  AOI22_X1 U20073 ( .A1(n16910), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16903) );
  AOI22_X1 U20074 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9720), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16902) );
  NAND4_X1 U20075 ( .A1(n16905), .A2(n16904), .A3(n16903), .A4(n16902), .ZN(
        n16906) );
  NOR2_X1 U20076 ( .A1(n16907), .A2(n16906), .ZN(n16983) );
  NOR2_X1 U20077 ( .A1(n16982), .A2(n16983), .ZN(n16981) );
  AOI22_X1 U20078 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17057), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n17166), .ZN(n16919) );
  AOI22_X1 U20079 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17173), .ZN(n16918) );
  INV_X1 U20080 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n20864) );
  AOI22_X1 U20081 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17193), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n16908) );
  OAI21_X1 U20082 ( .B1(n16909), .B2(n20864), .A(n16908), .ZN(n16916) );
  AOI22_X1 U20083 ( .A1(n17165), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16914) );
  AOI22_X1 U20084 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17190), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17162), .ZN(n16913) );
  AOI22_X1 U20085 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n16912) );
  AOI22_X1 U20086 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n17174), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n12992), .ZN(n16911) );
  NAND4_X1 U20087 ( .A1(n16914), .A2(n16913), .A3(n16912), .A4(n16911), .ZN(
        n16915) );
  AOI211_X1 U20088 ( .C1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .C2(n17192), .A(
        n16916), .B(n16915), .ZN(n16917) );
  NAND3_X1 U20089 ( .A1(n16919), .A2(n16918), .A3(n16917), .ZN(n16978) );
  NAND2_X1 U20090 ( .A1(n16981), .A2(n16978), .ZN(n16977) );
  NOR2_X1 U20091 ( .A1(n16973), .A2(n16977), .ZN(n16972) );
  AOI22_X1 U20092 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16929) );
  AOI22_X1 U20093 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n16928) );
  INV_X1 U20094 ( .A(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17131) );
  AOI22_X1 U20095 ( .A1(n17188), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n16920) );
  OAI21_X1 U20096 ( .B1(n17083), .B2(n17131), .A(n16920), .ZN(n16926) );
  AOI22_X1 U20097 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17165), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n16924) );
  AOI22_X1 U20098 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16923) );
  AOI22_X1 U20099 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n16922) );
  AOI22_X1 U20100 ( .A1(n17162), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16921) );
  NAND4_X1 U20101 ( .A1(n16924), .A2(n16923), .A3(n16922), .A4(n16921), .ZN(
        n16925) );
  AOI211_X1 U20102 ( .C1(n17183), .C2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n16926), .B(n16925), .ZN(n16927) );
  NAND3_X1 U20103 ( .A1(n16929), .A2(n16928), .A3(n16927), .ZN(n16969) );
  NAND2_X1 U20104 ( .A1(n16972), .A2(n16969), .ZN(n16968) );
  NOR2_X1 U20105 ( .A1(n16964), .A2(n16968), .ZN(n16963) );
  AOI22_X1 U20106 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16939) );
  AOI22_X1 U20107 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16938) );
  AOI22_X1 U20108 ( .A1(n17190), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n16930) );
  OAI21_X1 U20109 ( .B1(n17187), .B2(n20825), .A(n16930), .ZN(n16936) );
  AOI22_X1 U20110 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16934) );
  AOI22_X1 U20111 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16933) );
  AOI22_X1 U20112 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12832), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16932) );
  AOI22_X1 U20113 ( .A1(n17188), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16931) );
  NAND4_X1 U20114 ( .A1(n16934), .A2(n16933), .A3(n16932), .A4(n16931), .ZN(
        n16935) );
  AOI211_X1 U20115 ( .C1(n17192), .C2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n16936), .B(n16935), .ZN(n16937) );
  NAND3_X1 U20116 ( .A1(n16939), .A2(n16938), .A3(n16937), .ZN(n16958) );
  NAND2_X1 U20117 ( .A1(n16963), .A2(n16958), .ZN(n16957) );
  NOR2_X1 U20118 ( .A1(n16954), .A2(n16957), .ZN(n16953) );
  AOI22_X1 U20119 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16943) );
  AOI22_X1 U20120 ( .A1(n17188), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16942) );
  AOI22_X1 U20121 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16941) );
  AOI22_X1 U20122 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16940) );
  NAND4_X1 U20123 ( .A1(n16943), .A2(n16942), .A3(n16941), .A4(n16940), .ZN(
        n16949) );
  AOI22_X1 U20124 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12832), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n16947) );
  AOI22_X1 U20125 ( .A1(n17165), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17193), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16946) );
  AOI22_X1 U20126 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16945) );
  AOI22_X1 U20127 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16944) );
  NAND4_X1 U20128 ( .A1(n16947), .A2(n16946), .A3(n16945), .A4(n16944), .ZN(
        n16948) );
  NOR2_X1 U20129 ( .A1(n16949), .A2(n16948), .ZN(n16950) );
  XOR2_X1 U20130 ( .A(n16953), .B(n16950), .Z(n17249) );
  OAI22_X1 U20131 ( .A1(n16952), .A2(n16951), .B1(n17249), .B2(n17233), .ZN(
        P3_U2673) );
  NOR2_X1 U20132 ( .A1(n17330), .A2(n17038), .ZN(n17026) );
  NAND3_X1 U20133 ( .A1(P3_EBX_REG_23__SCAN_IN), .A2(P3_EBX_REG_22__SCAN_IN), 
        .A3(n16987), .ZN(n16980) );
  NAND2_X1 U20134 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16976), .ZN(n16967) );
  INV_X1 U20135 ( .A(n16967), .ZN(n16971) );
  NAND3_X1 U20136 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .A3(n16971), .ZN(n16959) );
  AOI21_X1 U20137 ( .B1(n16954), .B2(n16957), .A(n16953), .ZN(n17253) );
  INV_X1 U20138 ( .A(n17253), .ZN(n16956) );
  NAND3_X1 U20139 ( .A1(n16959), .A2(P3_EBX_REG_29__SCAN_IN), .A3(n17233), 
        .ZN(n16955) );
  OAI221_X1 U20140 ( .B1(n16959), .B2(P3_EBX_REG_29__SCAN_IN), .C1(n17233), 
        .C2(n16956), .A(n16955), .ZN(P3_U2674) );
  OAI21_X1 U20141 ( .B1(n16963), .B2(n16958), .A(n16957), .ZN(n17261) );
  NAND3_X1 U20142 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n17233), .A3(n16959), 
        .ZN(n16962) );
  OR3_X1 U20143 ( .A1(n16960), .A2(n16967), .A3(P3_EBX_REG_28__SCAN_IN), .ZN(
        n16961) );
  OAI211_X1 U20144 ( .C1(n17233), .C2(n17261), .A(n16962), .B(n16961), .ZN(
        P3_U2675) );
  AOI21_X1 U20145 ( .B1(n16964), .B2(n16968), .A(n16963), .ZN(n17262) );
  INV_X1 U20146 ( .A(n17262), .ZN(n16966) );
  NAND3_X1 U20147 ( .A1(n16967), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17233), 
        .ZN(n16965) );
  OAI221_X1 U20148 ( .B1(n16967), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17233), 
        .C2(n16966), .A(n16965), .ZN(P3_U2676) );
  AOI21_X1 U20149 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17233), .A(n16976), .ZN(
        n16970) );
  OAI21_X1 U20150 ( .B1(n16972), .B2(n16969), .A(n16968), .ZN(n17270) );
  OAI22_X1 U20151 ( .A1(n16971), .A2(n16970), .B1(n17270), .B2(n17233), .ZN(
        P3_U2677) );
  AOI22_X1 U20152 ( .A1(P3_EBX_REG_25__SCAN_IN), .A2(n17233), .B1(
        P3_EBX_REG_24__SCAN_IN), .B2(n16986), .ZN(n16975) );
  AOI21_X1 U20153 ( .B1(n16973), .B2(n16977), .A(n16972), .ZN(n17271) );
  INV_X1 U20154 ( .A(n17271), .ZN(n16974) );
  OAI22_X1 U20155 ( .A1(n16976), .A2(n16975), .B1(n16974), .B2(n17233), .ZN(
        P3_U2678) );
  OAI21_X1 U20156 ( .B1(n16981), .B2(n16978), .A(n16977), .ZN(n17281) );
  NAND3_X1 U20157 ( .A1(n16980), .A2(P3_EBX_REG_24__SCAN_IN), .A3(n17233), 
        .ZN(n16979) );
  OAI221_X1 U20158 ( .B1(n16980), .B2(P3_EBX_REG_24__SCAN_IN), .C1(n17233), 
        .C2(n17281), .A(n16979), .ZN(P3_U2679) );
  AND2_X1 U20159 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16987), .ZN(n17000) );
  AOI21_X1 U20160 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17233), .A(n17000), .ZN(
        n16985) );
  AOI21_X1 U20161 ( .B1(n16983), .B2(n16982), .A(n16981), .ZN(n17285) );
  INV_X1 U20162 ( .A(n17285), .ZN(n16984) );
  OAI22_X1 U20163 ( .A1(n16986), .A2(n16985), .B1(n16984), .B2(n17233), .ZN(
        P3_U2680) );
  AOI21_X1 U20164 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17233), .A(n16987), .ZN(
        n16999) );
  AOI22_X1 U20165 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16991) );
  AOI22_X1 U20166 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17193), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16990) );
  AOI22_X1 U20167 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16989) );
  AOI22_X1 U20168 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16988) );
  NAND4_X1 U20169 ( .A1(n16991), .A2(n16990), .A3(n16989), .A4(n16988), .ZN(
        n16998) );
  AOI22_X1 U20170 ( .A1(n16910), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17163), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16996) );
  AOI22_X1 U20171 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16995) );
  AOI22_X1 U20172 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16994) );
  AOI22_X1 U20173 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16993) );
  NAND4_X1 U20174 ( .A1(n16996), .A2(n16995), .A3(n16994), .A4(n16993), .ZN(
        n16997) );
  NOR2_X1 U20175 ( .A1(n16998), .A2(n16997), .ZN(n17290) );
  OAI22_X1 U20176 ( .A1(n17000), .A2(n16999), .B1(n17290), .B2(n17233), .ZN(
        P3_U2681) );
  AOI22_X1 U20177 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17004) );
  AOI22_X1 U20178 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17003) );
  AOI22_X1 U20179 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12867), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17002) );
  AOI22_X1 U20180 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17001) );
  NAND4_X1 U20181 ( .A1(n17004), .A2(n17003), .A3(n17002), .A4(n17001), .ZN(
        n17010) );
  AOI22_X1 U20182 ( .A1(n16910), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n17008) );
  AOI22_X1 U20183 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17007) );
  AOI22_X1 U20184 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17006) );
  AOI22_X1 U20185 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n17005) );
  NAND4_X1 U20186 ( .A1(n17008), .A2(n17007), .A3(n17006), .A4(n17005), .ZN(
        n17009) );
  NOR2_X1 U20187 ( .A1(n17010), .A2(n17009), .ZN(n17297) );
  NOR2_X1 U20188 ( .A1(n17238), .A2(n17011), .ZN(n17025) );
  AOI22_X1 U20189 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17025), .B1(n17013), 
        .B2(n17012), .ZN(n17014) );
  OAI21_X1 U20190 ( .B1(n17297), .B2(n17233), .A(n17014), .ZN(P3_U2682) );
  AOI22_X1 U20191 ( .A1(n9753), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17018) );
  AOI22_X1 U20192 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17017) );
  AOI22_X1 U20193 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17016) );
  AOI22_X1 U20194 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17015) );
  NAND4_X1 U20195 ( .A1(n17018), .A2(n17017), .A3(n17016), .A4(n17015), .ZN(
        n17024) );
  AOI22_X1 U20196 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17022) );
  AOI22_X1 U20197 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17021) );
  AOI22_X1 U20198 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17020) );
  AOI22_X1 U20199 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17019) );
  NAND4_X1 U20200 ( .A1(n17022), .A2(n17021), .A3(n17020), .A4(n17019), .ZN(
        n17023) );
  NOR2_X1 U20201 ( .A1(n17024), .A2(n17023), .ZN(n17302) );
  OAI21_X1 U20202 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n17026), .A(n17025), .ZN(
        n17027) );
  OAI21_X1 U20203 ( .B1(n17302), .B2(n17233), .A(n17027), .ZN(P3_U2683) );
  AOI22_X1 U20204 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17031) );
  AOI22_X1 U20205 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17030) );
  AOI22_X1 U20206 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17029) );
  AOI22_X1 U20207 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17028) );
  NAND4_X1 U20208 ( .A1(n17031), .A2(n17030), .A3(n17029), .A4(n17028), .ZN(
        n17037) );
  AOI22_X1 U20209 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17035) );
  AOI22_X1 U20210 ( .A1(n9753), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17034) );
  AOI22_X1 U20211 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17172), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17033) );
  AOI22_X1 U20212 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17032) );
  NAND4_X1 U20213 ( .A1(n17035), .A2(n17034), .A3(n17033), .A4(n17032), .ZN(
        n17036) );
  NOR2_X1 U20214 ( .A1(n17037), .A2(n17036), .ZN(n17306) );
  OAI21_X1 U20215 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n17039), .A(n17038), .ZN(
        n17040) );
  AOI22_X1 U20216 ( .A1(n17238), .A2(n17306), .B1(n17040), .B2(n17233), .ZN(
        P3_U2684) );
  AOI22_X1 U20217 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17044) );
  AOI22_X1 U20218 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17152), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17043) );
  AOI22_X1 U20219 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17042) );
  AOI22_X1 U20220 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17041) );
  NAND4_X1 U20221 ( .A1(n17044), .A2(n17043), .A3(n17042), .A4(n17041), .ZN(
        n17050) );
  AOI22_X1 U20222 ( .A1(n9753), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12832), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17048) );
  AOI22_X1 U20223 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17047) );
  AOI22_X1 U20224 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17046) );
  AOI22_X1 U20225 ( .A1(n17084), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17045) );
  NAND4_X1 U20226 ( .A1(n17048), .A2(n17047), .A3(n17046), .A4(n17045), .ZN(
        n17049) );
  NOR2_X1 U20227 ( .A1(n17050), .A2(n17049), .ZN(n17311) );
  INV_X1 U20228 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n17078) );
  NAND2_X1 U20229 ( .A1(n18245), .A2(n17077), .ZN(n17064) );
  NOR3_X1 U20230 ( .A1(n20806), .A2(n17078), .A3(n17064), .ZN(n17066) );
  OAI21_X1 U20231 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17066), .A(n17051), .ZN(
        n17052) );
  AOI22_X1 U20232 ( .A1(n17238), .A2(n17311), .B1(n17052), .B2(n17233), .ZN(
        P3_U2685) );
  AOI22_X1 U20233 ( .A1(n9753), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17056) );
  AOI22_X1 U20234 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17173), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17055) );
  AOI22_X1 U20235 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n12992), .ZN(n17054) );
  AOI22_X1 U20236 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17190), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17167), .ZN(n17053) );
  NAND4_X1 U20237 ( .A1(n17056), .A2(n17055), .A3(n17054), .A4(n17053), .ZN(
        n17063) );
  AOI22_X1 U20238 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n17162), .ZN(n17061) );
  AOI22_X1 U20239 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n17163), .ZN(n17060) );
  AOI22_X1 U20240 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17174), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17057), .ZN(n17059) );
  AOI22_X1 U20241 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17166), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17193), .ZN(n17058) );
  NAND4_X1 U20242 ( .A1(n17061), .A2(n17060), .A3(n17059), .A4(n17058), .ZN(
        n17062) );
  NOR2_X1 U20243 ( .A1(n17063), .A2(n17062), .ZN(n17315) );
  INV_X1 U20244 ( .A(n17064), .ZN(n17079) );
  AOI22_X1 U20245 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n17233), .B1(
        P3_EBX_REG_16__SCAN_IN), .B2(n17079), .ZN(n17065) );
  OAI22_X1 U20246 ( .A1(n17315), .A2(n17233), .B1(n17066), .B2(n17065), .ZN(
        P3_U2686) );
  AOI22_X1 U20247 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17070) );
  AOI22_X1 U20248 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17069) );
  AOI22_X1 U20249 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17068) );
  AOI22_X1 U20250 ( .A1(n17084), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17067) );
  NAND4_X1 U20251 ( .A1(n17070), .A2(n17069), .A3(n17068), .A4(n17067), .ZN(
        n17076) );
  AOI22_X1 U20252 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17074) );
  AOI22_X1 U20253 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17073) );
  AOI22_X1 U20254 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17072) );
  AOI22_X1 U20255 ( .A1(n9753), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17071) );
  NAND4_X1 U20256 ( .A1(n17074), .A2(n17073), .A3(n17072), .A4(n17071), .ZN(
        n17075) );
  NOR2_X1 U20257 ( .A1(n17076), .A2(n17075), .ZN(n17322) );
  NOR2_X1 U20258 ( .A1(n17238), .A2(n17077), .ZN(n17081) );
  AOI22_X1 U20259 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17081), .B1(n17079), 
        .B2(n17078), .ZN(n17080) );
  OAI21_X1 U20260 ( .B1(n17322), .B2(n17233), .A(n17080), .ZN(P3_U2687) );
  INV_X1 U20261 ( .A(n17081), .ZN(n17096) );
  AOI22_X1 U20262 ( .A1(n9753), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12867), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17093) );
  AOI22_X1 U20263 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17092) );
  INV_X1 U20264 ( .A(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n20822) );
  AOI22_X1 U20265 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17082) );
  OAI21_X1 U20266 ( .B1(n17083), .B2(n20822), .A(n17082), .ZN(n17090) );
  AOI22_X1 U20267 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17172), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17088) );
  AOI22_X1 U20268 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17087) );
  AOI22_X1 U20269 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17086) );
  AOI22_X1 U20270 ( .A1(n17084), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17085) );
  NAND4_X1 U20271 ( .A1(n17088), .A2(n17087), .A3(n17086), .A4(n17085), .ZN(
        n17089) );
  AOI211_X1 U20272 ( .C1(n17097), .C2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n17090), .B(n17089), .ZN(n17091) );
  NAND3_X1 U20273 ( .A1(n17093), .A2(n17092), .A3(n17091), .ZN(n17323) );
  NAND2_X1 U20274 ( .A1(n17238), .A2(n17323), .ZN(n17094) );
  OAI221_X1 U20275 ( .B1(n17096), .B2(n20783), .C1(n17096), .C2(n17095), .A(
        n17094), .ZN(P3_U2688) );
  AOI22_X1 U20276 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17101) );
  AOI22_X1 U20277 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17100) );
  AOI22_X1 U20278 ( .A1(n9753), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17099) );
  AOI22_X1 U20279 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17098) );
  NAND4_X1 U20280 ( .A1(n17101), .A2(n17100), .A3(n17099), .A4(n17098), .ZN(
        n17107) );
  AOI22_X1 U20281 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17105) );
  AOI22_X1 U20282 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17104) );
  AOI22_X1 U20283 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n17103) );
  AOI22_X1 U20284 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n17102) );
  NAND4_X1 U20285 ( .A1(n17105), .A2(n17104), .A3(n17103), .A4(n17102), .ZN(
        n17106) );
  NOR2_X1 U20286 ( .A1(n17107), .A2(n17106), .ZN(n17333) );
  OAI21_X1 U20287 ( .B1(n17109), .B2(n17108), .A(P3_EBX_REG_14__SCAN_IN), .ZN(
        n17114) );
  NOR2_X1 U20288 ( .A1(n21008), .A2(n17110), .ZN(n17112) );
  NAND4_X1 U20289 ( .A1(n18245), .A2(n17115), .A3(n17112), .A4(n17111), .ZN(
        n17113) );
  OAI211_X1 U20290 ( .C1(n17333), .C2(n17233), .A(n17114), .B(n17113), .ZN(
        P3_U2689) );
  NAND2_X1 U20291 ( .A1(n18245), .A2(n17115), .ZN(n17129) );
  NOR2_X1 U20292 ( .A1(n17238), .A2(n17115), .ZN(n17145) );
  AOI22_X1 U20293 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17127) );
  AOI22_X1 U20294 ( .A1(n12832), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17172), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17126) );
  AOI22_X1 U20295 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17116) );
  OAI21_X1 U20296 ( .B1(n17117), .B2(n21022), .A(n17116), .ZN(n17124) );
  AOI22_X1 U20297 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17122) );
  AOI22_X1 U20298 ( .A1(n17165), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17121) );
  AOI22_X1 U20299 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n17120) );
  AOI22_X1 U20300 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17119) );
  NAND4_X1 U20301 ( .A1(n17122), .A2(n17121), .A3(n17120), .A4(n17119), .ZN(
        n17123) );
  AOI211_X1 U20302 ( .C1(n17164), .C2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n17124), .B(n17123), .ZN(n17125) );
  NAND3_X1 U20303 ( .A1(n17127), .A2(n17126), .A3(n17125), .ZN(n17338) );
  AOI22_X1 U20304 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n17145), .B1(n17238), 
        .B2(n17338), .ZN(n17128) );
  OAI21_X1 U20305 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17129), .A(n17128), .ZN(
        P3_U2691) );
  AOI22_X1 U20306 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17141) );
  AOI22_X1 U20307 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17140) );
  AOI22_X1 U20308 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17172), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17130) );
  OAI21_X1 U20309 ( .B1(n17132), .B2(n17131), .A(n17130), .ZN(n17138) );
  AOI22_X1 U20310 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17136) );
  AOI22_X1 U20311 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17135) );
  AOI22_X1 U20312 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17134) );
  AOI22_X1 U20313 ( .A1(n17167), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17133) );
  NAND4_X1 U20314 ( .A1(n17136), .A2(n17135), .A3(n17134), .A4(n17133), .ZN(
        n17137) );
  AOI211_X1 U20315 ( .C1(n9753), .C2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A(
        n17138), .B(n17137), .ZN(n17139) );
  NAND3_X1 U20316 ( .A1(n17141), .A2(n17140), .A3(n17139), .ZN(n17342) );
  INV_X1 U20317 ( .A(n17342), .ZN(n17147) );
  INV_X1 U20318 ( .A(n17208), .ZN(n17211) );
  NAND2_X1 U20319 ( .A1(n17235), .A2(n17142), .ZN(n17209) );
  INV_X1 U20320 ( .A(n17209), .ZN(n17218) );
  NAND3_X1 U20321 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17211), .A3(n17218), .ZN(
        n17205) );
  NOR3_X1 U20322 ( .A1(n17143), .A2(n17204), .A3(n17205), .ZN(n17159) );
  INV_X1 U20323 ( .A(n17159), .ZN(n17181) );
  NOR2_X1 U20324 ( .A1(n17144), .A2(n17181), .ZN(n17161) );
  OAI21_X1 U20325 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17161), .A(n17145), .ZN(
        n17146) );
  OAI21_X1 U20326 ( .B1(n17147), .B2(n17233), .A(n17146), .ZN(P3_U2692) );
  AOI22_X1 U20327 ( .A1(n17166), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17151) );
  AOI22_X1 U20328 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17150) );
  AOI22_X1 U20329 ( .A1(n17163), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17149) );
  AOI22_X1 U20330 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17167), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17148) );
  NAND4_X1 U20331 ( .A1(n17151), .A2(n17150), .A3(n17149), .A4(n17148), .ZN(
        n17158) );
  AOI22_X1 U20332 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17184), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17156) );
  AOI22_X1 U20333 ( .A1(n17152), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17162), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17155) );
  AOI22_X1 U20334 ( .A1(n9753), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17154) );
  AOI22_X1 U20335 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17097), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17153) );
  NAND4_X1 U20336 ( .A1(n17156), .A2(n17155), .A3(n17154), .A4(n17153), .ZN(
        n17157) );
  NOR2_X1 U20337 ( .A1(n17158), .A2(n17157), .ZN(n17345) );
  OAI21_X1 U20338 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17159), .A(n17233), .ZN(
        n17160) );
  OAI22_X1 U20339 ( .A1(n17345), .A2(n17233), .B1(n17161), .B2(n17160), .ZN(
        P3_U2693) );
  AOI22_X1 U20340 ( .A1(n17183), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17162), .ZN(n17171) );
  AOI22_X1 U20341 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n17163), .ZN(n17170) );
  AOI22_X1 U20342 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n17166), .B1(
        n16910), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17169) );
  AOI22_X1 U20343 ( .A1(n17097), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n17167), .ZN(n17168) );
  NAND4_X1 U20344 ( .A1(n17171), .A2(n17170), .A3(n17169), .A4(n17168), .ZN(
        n17180) );
  AOI22_X1 U20345 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17188), .B1(
        n17172), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17178) );
  AOI22_X1 U20346 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n17173), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n17190), .ZN(n17177) );
  AOI22_X1 U20347 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17174), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n12992), .ZN(n17176) );
  AOI22_X1 U20348 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17118), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17175) );
  NAND4_X1 U20349 ( .A1(n17178), .A2(n17177), .A3(n17176), .A4(n17175), .ZN(
        n17179) );
  NOR2_X1 U20350 ( .A1(n17180), .A2(n17179), .ZN(n17350) );
  INV_X1 U20351 ( .A(n17205), .ZN(n17203) );
  OAI221_X1 U20352 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(P3_EBX_REG_8__SCAN_IN), 
        .C1(P3_EBX_REG_9__SCAN_IN), .C2(n17203), .A(n17181), .ZN(n17182) );
  AOI22_X1 U20353 ( .A1(n17238), .A2(n17350), .B1(n17182), .B2(n17233), .ZN(
        P3_U2694) );
  AOI22_X1 U20354 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17183), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17202) );
  AOI22_X1 U20355 ( .A1(n17184), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17166), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17201) );
  AOI22_X1 U20356 ( .A1(n17118), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17185), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17186) );
  OAI21_X1 U20357 ( .B1(n17187), .B2(n20743), .A(n17186), .ZN(n17199) );
  AOI22_X1 U20358 ( .A1(n17189), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17188), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17197) );
  AOI22_X1 U20359 ( .A1(n17191), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17190), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17196) );
  AOI22_X1 U20360 ( .A1(n9720), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17192), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17195) );
  AOI22_X1 U20361 ( .A1(n17193), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12992), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17194) );
  NAND4_X1 U20362 ( .A1(n17197), .A2(n17196), .A3(n17195), .A4(n17194), .ZN(
        n17198) );
  AOI211_X1 U20363 ( .C1(n12832), .C2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A(
        n17199), .B(n17198), .ZN(n17200) );
  NAND3_X1 U20364 ( .A1(n17202), .A2(n17201), .A3(n17200), .ZN(n17357) );
  OAI33_X1 U20365 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17330), .A3(n17205), .B1(
        n17204), .B2(n17238), .B3(n17203), .ZN(n17206) );
  AOI21_X1 U20366 ( .B1(n17238), .B2(n17357), .A(n17206), .ZN(n17207) );
  INV_X1 U20367 ( .A(n17207), .ZN(P3_U2695) );
  OAI21_X1 U20368 ( .B1(n17208), .B2(n17209), .A(P3_EBX_REG_7__SCAN_IN), .ZN(
        n17214) );
  INV_X1 U20369 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17213) );
  NOR2_X1 U20370 ( .A1(n17330), .A2(n17209), .ZN(n17224) );
  NAND3_X1 U20371 ( .A1(n17211), .A2(n17224), .A3(n17210), .ZN(n17212) );
  OAI221_X1 U20372 ( .B1(n17238), .B2(n17214), .C1(n17233), .C2(n17213), .A(
        n17212), .ZN(P3_U2696) );
  NAND2_X1 U20373 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17224), .ZN(n17217) );
  INV_X1 U20374 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17216) );
  NAND3_X1 U20375 ( .A1(n17217), .A2(P3_EBX_REG_6__SCAN_IN), .A3(n17233), .ZN(
        n17215) );
  OAI221_X1 U20376 ( .B1(n17217), .B2(P3_EBX_REG_6__SCAN_IN), .C1(n17233), 
        .C2(n17216), .A(n17215), .ZN(P3_U2697) );
  INV_X1 U20377 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17220) );
  OAI211_X1 U20378 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n17218), .A(n17217), .B(
        n17233), .ZN(n17219) );
  OAI21_X1 U20379 ( .B1(n17233), .B2(n17220), .A(n17219), .ZN(P3_U2698) );
  NOR2_X1 U20380 ( .A1(n17221), .A2(n17240), .ZN(n17230) );
  AOI22_X1 U20381 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17233), .B1(
        P3_EBX_REG_3__SCAN_IN), .B2(n17230), .ZN(n17223) );
  INV_X1 U20382 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17222) );
  OAI22_X1 U20383 ( .A1(n17224), .A2(n17223), .B1(n17222), .B2(n17233), .ZN(
        P3_U2699) );
  INV_X1 U20384 ( .A(n17230), .ZN(n17227) );
  INV_X1 U20385 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17226) );
  NAND3_X1 U20386 ( .A1(n17227), .A2(P3_EBX_REG_3__SCAN_IN), .A3(n17233), .ZN(
        n17225) );
  OAI221_X1 U20387 ( .B1(n17227), .B2(P3_EBX_REG_3__SCAN_IN), .C1(n17233), 
        .C2(n17226), .A(n17225), .ZN(P3_U2700) );
  INV_X1 U20388 ( .A(n17228), .ZN(n17229) );
  AOI221_X1 U20389 ( .B1(n17229), .B2(n17235), .C1(n17330), .C2(n17235), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17231) );
  AOI211_X1 U20390 ( .C1(n17238), .C2(n17232), .A(n17231), .B(n17230), .ZN(
        P3_U2701) );
  INV_X1 U20391 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17234) );
  OAI222_X1 U20392 ( .A1(n17240), .A2(n17236), .B1(n20848), .B2(n17235), .C1(
        n17234), .C2(n17233), .ZN(P3_U2702) );
  AOI22_X1 U20393 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17238), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17237), .ZN(n17239) );
  OAI21_X1 U20394 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17240), .A(n17239), .ZN(
        P3_U2703) );
  INV_X1 U20395 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17472) );
  INV_X1 U20396 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17468) );
  INV_X1 U20397 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17466) );
  INV_X1 U20398 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17450) );
  INV_X1 U20399 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17427) );
  NAND2_X1 U20400 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(P3_EAX_REG_1__SCAN_IN), 
        .ZN(n17360) );
  NAND2_X1 U20401 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .ZN(n17361) );
  NAND4_X1 U20402 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17241) );
  NOR3_X1 U20403 ( .A1(n17360), .A2(n17361), .A3(n17241), .ZN(n17365) );
  INV_X1 U20404 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17500) );
  INV_X1 U20405 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17498) );
  INV_X1 U20406 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17423) );
  NOR3_X1 U20407 ( .A1(n17500), .A2(n17498), .A3(n17423), .ZN(n17334) );
  INV_X1 U20408 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17504) );
  INV_X1 U20409 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17458) );
  INV_X1 U20410 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17456) );
  INV_X1 U20411 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17454) );
  INV_X1 U20412 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17452) );
  NOR4_X1 U20413 ( .A1(n17458), .A2(n17456), .A3(n17454), .A4(n17452), .ZN(
        n17288) );
  AND2_X1 U20414 ( .A1(n17288), .A2(n10138), .ZN(n17244) );
  INV_X1 U20415 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17464) );
  NAND2_X1 U20416 ( .A1(n18245), .A2(n17282), .ZN(n17276) );
  NAND2_X1 U20417 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17263), .ZN(n17258) );
  NAND2_X1 U20418 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17255), .ZN(n17254) );
  NOR2_X1 U20419 ( .A1(P3_EAX_REG_31__SCAN_IN), .A2(n17254), .ZN(n17246) );
  NAND2_X1 U20420 ( .A1(n17389), .A2(n17254), .ZN(n17252) );
  OAI21_X1 U20421 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17359), .A(n17252), .ZN(
        n17245) );
  AOI22_X1 U20422 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17246), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17245), .ZN(n17247) );
  OAI21_X1 U20423 ( .B1(n18241), .B2(n17289), .A(n17247), .ZN(P3_U2704) );
  INV_X1 U20424 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17478) );
  NOR2_X2 U20425 ( .A1(n17248), .A2(n17389), .ZN(n17317) );
  OAI22_X1 U20426 ( .A1(n17249), .A2(n17384), .B1(n19244), .B2(n17289), .ZN(
        n17250) );
  AOI21_X1 U20427 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17317), .A(n17250), .ZN(
        n17251) );
  OAI221_X1 U20428 ( .B1(P3_EAX_REG_30__SCAN_IN), .B2(n17254), .C1(n17478), 
        .C2(n17252), .A(n17251), .ZN(P3_U2705) );
  AOI22_X1 U20429 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17317), .B1(n17392), .B2(
        n17253), .ZN(n17257) );
  OAI211_X1 U20430 ( .C1(n17255), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17389), .B(
        n17254), .ZN(n17256) );
  OAI211_X1 U20431 ( .C1(n17289), .C2(n18232), .A(n17257), .B(n17256), .ZN(
        P3_U2706) );
  AOI22_X1 U20432 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17317), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17316), .ZN(n17260) );
  OAI211_X1 U20433 ( .C1(n17263), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17389), .B(
        n17258), .ZN(n17259) );
  OAI211_X1 U20434 ( .C1(n17261), .C2(n17384), .A(n17260), .B(n17259), .ZN(
        P3_U2707) );
  INV_X1 U20435 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n20810) );
  AOI22_X1 U20436 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17317), .B1(n17392), .B2(
        n17262), .ZN(n17266) );
  AOI211_X1 U20437 ( .C1(n17472), .C2(n17267), .A(n17263), .B(n17354), .ZN(
        n17264) );
  INV_X1 U20438 ( .A(n17264), .ZN(n17265) );
  OAI211_X1 U20439 ( .C1(n17289), .C2(n20810), .A(n17266), .B(n17265), .ZN(
        P3_U2708) );
  AOI22_X1 U20440 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17317), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17316), .ZN(n17269) );
  OAI211_X1 U20441 ( .C1(n17272), .C2(P3_EAX_REG_26__SCAN_IN), .A(n17389), .B(
        n17267), .ZN(n17268) );
  OAI211_X1 U20442 ( .C1(n17270), .C2(n17384), .A(n17269), .B(n17268), .ZN(
        P3_U2709) );
  AOI22_X1 U20443 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17317), .B1(n17392), .B2(
        n17271), .ZN(n17275) );
  AOI211_X1 U20444 ( .C1(n17468), .C2(n17277), .A(n17272), .B(n17354), .ZN(
        n17273) );
  INV_X1 U20445 ( .A(n17273), .ZN(n17274) );
  OAI211_X1 U20446 ( .C1(n17289), .C2(n18216), .A(n17275), .B(n17274), .ZN(
        P3_U2710) );
  AOI22_X1 U20447 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17317), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17316), .ZN(n17280) );
  OAI21_X1 U20448 ( .B1(n17466), .B2(n17354), .A(n17276), .ZN(n17278) );
  NAND2_X1 U20449 ( .A1(n17278), .A2(n17277), .ZN(n17279) );
  OAI211_X1 U20450 ( .C1(n17281), .C2(n17384), .A(n17280), .B(n17279), .ZN(
        P3_U2711) );
  AOI22_X1 U20451 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17317), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17316), .ZN(n17287) );
  AOI211_X1 U20452 ( .C1(n17464), .C2(n17283), .A(n17354), .B(n17282), .ZN(
        n17284) );
  AOI21_X1 U20453 ( .B1(n17285), .B2(n17392), .A(n17284), .ZN(n17286) );
  NAND2_X1 U20454 ( .A1(n17287), .A2(n17286), .ZN(P3_U2712) );
  AND3_X1 U20455 ( .A1(n18245), .A2(n17318), .A3(n17288), .ZN(n17298) );
  NAND2_X1 U20456 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17298), .ZN(n17294) );
  NAND2_X1 U20457 ( .A1(n17294), .A2(P3_EAX_REG_22__SCAN_IN), .ZN(n17293) );
  OAI22_X1 U20458 ( .A1(n17290), .A2(n17384), .B1(n15003), .B2(n17289), .ZN(
        n17291) );
  AOI21_X1 U20459 ( .B1(BUF2_REG_6__SCAN_IN), .B2(n17317), .A(n17291), .ZN(
        n17292) );
  OAI221_X1 U20460 ( .B1(n17294), .B2(P3_EAX_REG_22__SCAN_IN), .C1(n17293), 
        .C2(n17354), .A(n17292), .ZN(P3_U2713) );
  AOI22_X1 U20461 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17317), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n17316), .ZN(n17296) );
  OAI211_X1 U20462 ( .C1(n17298), .C2(P3_EAX_REG_21__SCAN_IN), .A(n17389), .B(
        n17294), .ZN(n17295) );
  OAI211_X1 U20463 ( .C1(n17297), .C2(n17384), .A(n17296), .B(n17295), .ZN(
        P3_U2714) );
  AOI22_X1 U20464 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17317), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17316), .ZN(n17301) );
  NAND2_X1 U20465 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17318), .ZN(n17312) );
  NOR2_X1 U20466 ( .A1(n17454), .A2(n17312), .ZN(n17307) );
  NAND2_X1 U20467 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17307), .ZN(n17303) );
  AOI211_X1 U20468 ( .C1(n17458), .C2(n17303), .A(n17298), .B(n17354), .ZN(
        n17299) );
  INV_X1 U20469 ( .A(n17299), .ZN(n17300) );
  OAI211_X1 U20470 ( .C1(n17302), .C2(n17384), .A(n17301), .B(n17300), .ZN(
        P3_U2715) );
  AOI22_X1 U20471 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17317), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17316), .ZN(n17305) );
  OAI211_X1 U20472 ( .C1(n17307), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17389), .B(
        n17303), .ZN(n17304) );
  OAI211_X1 U20473 ( .C1(n17306), .C2(n17384), .A(n17305), .B(n17304), .ZN(
        P3_U2716) );
  AOI22_X1 U20474 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17317), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17316), .ZN(n17310) );
  AOI211_X1 U20475 ( .C1(n17454), .C2(n17312), .A(n17307), .B(n17354), .ZN(
        n17308) );
  INV_X1 U20476 ( .A(n17308), .ZN(n17309) );
  OAI211_X1 U20477 ( .C1(n17311), .C2(n17384), .A(n17310), .B(n17309), .ZN(
        P3_U2717) );
  AOI22_X1 U20478 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17317), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17316), .ZN(n17314) );
  OAI211_X1 U20479 ( .C1(n17318), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17389), .B(
        n17312), .ZN(n17313) );
  OAI211_X1 U20480 ( .C1(n17315), .C2(n17384), .A(n17314), .B(n17313), .ZN(
        P3_U2718) );
  AOI22_X1 U20481 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17317), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17316), .ZN(n17321) );
  AOI211_X1 U20482 ( .C1(n17450), .C2(n17324), .A(n17354), .B(n17318), .ZN(
        n17319) );
  INV_X1 U20483 ( .A(n17319), .ZN(n17320) );
  OAI211_X1 U20484 ( .C1(n17322), .C2(n17384), .A(n17321), .B(n17320), .ZN(
        P3_U2719) );
  AOI22_X1 U20485 ( .A1(n17392), .A2(n17323), .B1(BUF2_REG_15__SCAN_IN), .B2(
        n17393), .ZN(n17327) );
  OAI211_X1 U20486 ( .C1(P3_EAX_REG_15__SCAN_IN), .C2(n17325), .A(n17389), .B(
        n17324), .ZN(n17326) );
  NAND2_X1 U20487 ( .A1(n17327), .A2(n17326), .ZN(P3_U2720) );
  INV_X1 U20488 ( .A(n17329), .ZN(n17328) );
  OAI33_X1 U20489 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17330), .A3(n17329), 
        .B1(n17504), .B2(n17354), .B3(n17328), .ZN(n17331) );
  AOI21_X1 U20490 ( .B1(BUF2_REG_14__SCAN_IN), .B2(n17393), .A(n17331), .ZN(
        n17332) );
  OAI21_X1 U20491 ( .B1(n17333), .B2(n17384), .A(n17332), .ZN(P3_U2721) );
  INV_X1 U20492 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17425) );
  NAND2_X1 U20493 ( .A1(n18245), .A2(n17353), .ZN(n17348) );
  NAND2_X1 U20494 ( .A1(n17334), .A2(n17352), .ZN(n17337) );
  INV_X1 U20495 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17502) );
  NAND2_X1 U20496 ( .A1(n17389), .A2(n17337), .ZN(n17340) );
  AOI22_X1 U20497 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17393), .B1(n17392), .B2(
        n17335), .ZN(n17336) );
  OAI221_X1 U20498 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17337), .C1(n17502), 
        .C2(n17340), .A(n17336), .ZN(P3_U2722) );
  NAND3_X1 U20499 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(P3_EAX_REG_10__SCAN_IN), 
        .A3(n17352), .ZN(n17341) );
  AOI22_X1 U20500 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17393), .B1(n17392), .B2(
        n17338), .ZN(n17339) );
  OAI221_X1 U20501 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17341), .C1(n17500), 
        .C2(n17340), .A(n17339), .ZN(P3_U2723) );
  NAND2_X1 U20502 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17352), .ZN(n17344) );
  NAND2_X1 U20503 ( .A1(n17389), .A2(n17344), .ZN(n17347) );
  AOI22_X1 U20504 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17393), .B1(n17392), .B2(
        n17342), .ZN(n17343) );
  OAI221_X1 U20505 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17344), .C1(n17498), 
        .C2(n17347), .A(n17343), .ZN(P3_U2724) );
  NOR2_X1 U20506 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17352), .ZN(n17346) );
  OAI222_X1 U20507 ( .A1(n17387), .A2(n17496), .B1(n17347), .B2(n17346), .C1(
        n17384), .C2(n17345), .ZN(P3_U2725) );
  OAI21_X1 U20508 ( .B1(n17425), .B2(n17354), .A(n17348), .ZN(n17349) );
  INV_X1 U20509 ( .A(n17349), .ZN(n17351) );
  OAI222_X1 U20510 ( .A1(n17387), .A2(n17492), .B1(n17352), .B2(n17351), .C1(
        n17384), .C2(n17350), .ZN(P3_U2726) );
  AOI211_X1 U20511 ( .C1(n17427), .C2(n17355), .A(n17354), .B(n17353), .ZN(
        n17356) );
  AOI21_X1 U20512 ( .B1(n17392), .B2(n17357), .A(n17356), .ZN(n17358) );
  OAI21_X1 U20513 ( .B1(n17489), .B2(n17387), .A(n17358), .ZN(P3_U2727) );
  INV_X1 U20514 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17436) );
  NOR2_X1 U20515 ( .A1(n17360), .A2(n17359), .ZN(n17396) );
  NAND2_X1 U20516 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17396), .ZN(n17379) );
  NOR2_X1 U20517 ( .A1(n17436), .A2(n17379), .ZN(n17382) );
  NAND2_X1 U20518 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17382), .ZN(n17371) );
  NOR2_X1 U20519 ( .A1(n17361), .A2(n17371), .ZN(n17370) );
  AOI21_X1 U20520 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17389), .A(n17370), .ZN(
        n17366) );
  AOI22_X1 U20521 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17393), .B1(n17392), .B2(
        n17362), .ZN(n17363) );
  OAI221_X1 U20522 ( .B1(n17366), .B2(n17365), .C1(n17366), .C2(n17364), .A(
        n17363), .ZN(P3_U2728) );
  INV_X1 U20523 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18237) );
  INV_X1 U20524 ( .A(n17371), .ZN(n17378) );
  AOI22_X1 U20525 ( .A1(n17378), .A2(P3_EAX_REG_5__SCAN_IN), .B1(
        P3_EAX_REG_6__SCAN_IN), .B2(n17389), .ZN(n17369) );
  INV_X1 U20526 ( .A(n17367), .ZN(n17368) );
  OAI222_X1 U20527 ( .A1(n17387), .A2(n18237), .B1(n17370), .B2(n17369), .C1(
        n17384), .C2(n17368), .ZN(P3_U2729) );
  INV_X1 U20528 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18233) );
  INV_X1 U20529 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17432) );
  NOR2_X1 U20530 ( .A1(n17432), .A2(n17371), .ZN(n17374) );
  AOI21_X1 U20531 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17389), .A(n17378), .ZN(
        n17373) );
  OAI222_X1 U20532 ( .A1(n18233), .A2(n17387), .B1(n17374), .B2(n17373), .C1(
        n17384), .C2(n17372), .ZN(P3_U2730) );
  AOI21_X1 U20533 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17389), .A(n17382), .ZN(
        n17377) );
  INV_X1 U20534 ( .A(n17375), .ZN(n17376) );
  OAI222_X1 U20535 ( .A1(n18228), .A2(n17387), .B1(n17378), .B2(n17377), .C1(
        n17384), .C2(n17376), .ZN(P3_U2731) );
  INV_X1 U20536 ( .A(n17379), .ZN(n17386) );
  AOI21_X1 U20537 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17389), .A(n17386), .ZN(
        n17381) );
  OAI222_X1 U20538 ( .A1(n18224), .A2(n17387), .B1(n17382), .B2(n17381), .C1(
        n17384), .C2(n17380), .ZN(P3_U2732) );
  AOI21_X1 U20539 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17389), .A(n17396), .ZN(
        n17385) );
  OAI222_X1 U20540 ( .A1(n20804), .A2(n17387), .B1(n17386), .B2(n17385), .C1(
        n17384), .C2(n17383), .ZN(P3_U2733) );
  NOR2_X1 U20541 ( .A1(n17388), .A2(n20971), .ZN(n17390) );
  OAI21_X1 U20542 ( .B1(P3_EAX_REG_1__SCAN_IN), .B2(n17390), .A(n17389), .ZN(
        n17395) );
  AOI22_X1 U20543 ( .A1(n17393), .A2(BUF2_REG_1__SCAN_IN), .B1(n17392), .B2(
        n17391), .ZN(n17394) );
  OAI21_X1 U20544 ( .B1(n17396), .B2(n17395), .A(n17394), .ZN(P3_U2734) );
  INV_X1 U20545 ( .A(n18721), .ZN(n17553) );
  NAND2_X1 U20546 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17553), .ZN(n17410) );
  NOR2_X1 U20547 ( .A1(n17438), .A2(n17398), .ZN(P3_U2736) );
  NOR2_X1 U20548 ( .A1(n17442), .A2(n18213), .ZN(n17408) );
  INV_X2 U20549 ( .A(n17410), .ZN(n17440) );
  AOI22_X1 U20550 ( .A1(n17440), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17399) );
  OAI21_X1 U20551 ( .B1(n17478), .B2(n17416), .A(n17399), .ZN(P3_U2737) );
  INV_X1 U20552 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17476) );
  AOI22_X1 U20553 ( .A1(n17440), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17400) );
  OAI21_X1 U20554 ( .B1(n17476), .B2(n17416), .A(n17400), .ZN(P3_U2738) );
  INV_X1 U20555 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17474) );
  AOI22_X1 U20556 ( .A1(n17440), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17401) );
  OAI21_X1 U20557 ( .B1(n17474), .B2(n17416), .A(n17401), .ZN(P3_U2739) );
  AOI22_X1 U20558 ( .A1(n17440), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17402) );
  OAI21_X1 U20559 ( .B1(n17472), .B2(n17416), .A(n17402), .ZN(P3_U2740) );
  INV_X1 U20560 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17470) );
  AOI22_X1 U20561 ( .A1(n17440), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17403) );
  OAI21_X1 U20562 ( .B1(n17470), .B2(n17416), .A(n17403), .ZN(P3_U2741) );
  AOI22_X1 U20563 ( .A1(n17440), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17404) );
  OAI21_X1 U20564 ( .B1(n17468), .B2(n17416), .A(n17404), .ZN(P3_U2742) );
  AOI22_X1 U20565 ( .A1(n17440), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17405) );
  OAI21_X1 U20566 ( .B1(n17466), .B2(n17416), .A(n17405), .ZN(P3_U2743) );
  AOI22_X1 U20567 ( .A1(n17440), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17406) );
  OAI21_X1 U20568 ( .B1(n17464), .B2(n17416), .A(n17406), .ZN(P3_U2744) );
  INV_X1 U20569 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17462) );
  AOI22_X1 U20570 ( .A1(n17440), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17407) );
  OAI21_X1 U20571 ( .B1(n17462), .B2(n17416), .A(n17407), .ZN(P3_U2745) );
  INV_X1 U20572 ( .A(P3_UWORD_REG_5__SCAN_IN), .ZN(n20972) );
  AOI22_X1 U20573 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17408), .B1(n17439), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17409) );
  OAI21_X1 U20574 ( .B1(n20972), .B2(n17410), .A(n17409), .ZN(P3_U2746) );
  AOI22_X1 U20575 ( .A1(n17440), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17411) );
  OAI21_X1 U20576 ( .B1(n17458), .B2(n17416), .A(n17411), .ZN(P3_U2747) );
  AOI22_X1 U20577 ( .A1(n17440), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17412) );
  OAI21_X1 U20578 ( .B1(n17456), .B2(n17416), .A(n17412), .ZN(P3_U2748) );
  AOI22_X1 U20579 ( .A1(n17440), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17413) );
  OAI21_X1 U20580 ( .B1(n17454), .B2(n17416), .A(n17413), .ZN(P3_U2749) );
  AOI22_X1 U20581 ( .A1(n17440), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17414) );
  OAI21_X1 U20582 ( .B1(n17452), .B2(n17416), .A(n17414), .ZN(P3_U2750) );
  AOI22_X1 U20583 ( .A1(P3_DATAO_REG_16__SCAN_IN), .A2(n17439), .B1(n17440), 
        .B2(P3_UWORD_REG_0__SCAN_IN), .ZN(n17415) );
  OAI21_X1 U20584 ( .B1(n17450), .B2(n17416), .A(n17415), .ZN(P3_U2751) );
  INV_X1 U20585 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17509) );
  AOI22_X1 U20586 ( .A1(n17440), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17417) );
  OAI21_X1 U20587 ( .B1(n17509), .B2(n17442), .A(n17417), .ZN(P3_U2752) );
  AOI22_X1 U20588 ( .A1(n17440), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17418) );
  OAI21_X1 U20589 ( .B1(n17504), .B2(n17442), .A(n17418), .ZN(P3_U2753) );
  AOI22_X1 U20590 ( .A1(n17440), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17419) );
  OAI21_X1 U20591 ( .B1(n17502), .B2(n17442), .A(n17419), .ZN(P3_U2754) );
  AOI22_X1 U20592 ( .A1(n17440), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17420) );
  OAI21_X1 U20593 ( .B1(n17500), .B2(n17442), .A(n17420), .ZN(P3_U2755) );
  AOI22_X1 U20594 ( .A1(n17440), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17421) );
  OAI21_X1 U20595 ( .B1(n17498), .B2(n17442), .A(n17421), .ZN(P3_U2756) );
  AOI22_X1 U20596 ( .A1(n17440), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17422) );
  OAI21_X1 U20597 ( .B1(n17423), .B2(n17442), .A(n17422), .ZN(P3_U2757) );
  AOI22_X1 U20598 ( .A1(n17440), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17424) );
  OAI21_X1 U20599 ( .B1(n17425), .B2(n17442), .A(n17424), .ZN(P3_U2758) );
  AOI22_X1 U20600 ( .A1(n17440), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17426) );
  OAI21_X1 U20601 ( .B1(n17427), .B2(n17442), .A(n17426), .ZN(P3_U2759) );
  INV_X1 U20602 ( .A(P3_DATAO_REG_7__SCAN_IN), .ZN(n20823) );
  AOI22_X1 U20603 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17443), .B1(n17440), .B2(
        P3_LWORD_REG_7__SCAN_IN), .ZN(n17428) );
  OAI21_X1 U20604 ( .B1(n20823), .B2(n17438), .A(n17428), .ZN(P3_U2760) );
  INV_X1 U20605 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17430) );
  AOI22_X1 U20606 ( .A1(n17440), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17429) );
  OAI21_X1 U20607 ( .B1(n17430), .B2(n17442), .A(n17429), .ZN(P3_U2761) );
  AOI22_X1 U20608 ( .A1(n17440), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17431) );
  OAI21_X1 U20609 ( .B1(n17432), .B2(n17442), .A(n17431), .ZN(P3_U2762) );
  INV_X1 U20610 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17434) );
  AOI22_X1 U20611 ( .A1(n17440), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17433) );
  OAI21_X1 U20612 ( .B1(n17434), .B2(n17442), .A(n17433), .ZN(P3_U2763) );
  AOI22_X1 U20613 ( .A1(n17440), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17435) );
  OAI21_X1 U20614 ( .B1(n17436), .B2(n17442), .A(n17435), .ZN(P3_U2764) );
  INV_X1 U20615 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n20837) );
  AOI22_X1 U20616 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17443), .B1(n17440), .B2(
        P3_LWORD_REG_2__SCAN_IN), .ZN(n17437) );
  OAI21_X1 U20617 ( .B1(n20837), .B2(n17438), .A(n17437), .ZN(P3_U2765) );
  INV_X1 U20618 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17481) );
  AOI22_X1 U20619 ( .A1(n17440), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17439), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17441) );
  OAI21_X1 U20620 ( .B1(n17481), .B2(n17442), .A(n17441), .ZN(P3_U2766) );
  AOI222_X1 U20621 ( .A1(P3_LWORD_REG_0__SCAN_IN), .A2(n17440), .B1(n17443), 
        .B2(P3_EAX_REG_0__SCAN_IN), .C1(n17439), .C2(P3_DATAO_REG_0__SCAN_IN), 
        .ZN(n17444) );
  INV_X1 U20622 ( .A(n17444), .ZN(P3_U2767) );
  AOI22_X1 U20623 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17506), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17490), .ZN(n17449) );
  OAI21_X1 U20624 ( .B1(n17450), .B2(n17508), .A(n17449), .ZN(P3_U2768) );
  AOI22_X1 U20625 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17506), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17490), .ZN(n17451) );
  OAI21_X1 U20626 ( .B1(n17452), .B2(n17508), .A(n17451), .ZN(P3_U2769) );
  AOI22_X1 U20627 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17506), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17490), .ZN(n17453) );
  OAI21_X1 U20628 ( .B1(n17454), .B2(n17508), .A(n17453), .ZN(P3_U2770) );
  AOI22_X1 U20629 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17506), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17490), .ZN(n17455) );
  OAI21_X1 U20630 ( .B1(n17456), .B2(n17508), .A(n17455), .ZN(P3_U2771) );
  AOI22_X1 U20631 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17506), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17490), .ZN(n17457) );
  OAI21_X1 U20632 ( .B1(n17458), .B2(n17508), .A(n17457), .ZN(P3_U2772) );
  INV_X1 U20633 ( .A(n17508), .ZN(n17493) );
  AOI22_X1 U20634 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17506), .B1(
        P3_EAX_REG_21__SCAN_IN), .B2(n17493), .ZN(n17459) );
  OAI21_X1 U20635 ( .B1(n17460), .B2(n20972), .A(n17459), .ZN(P3_U2773) );
  AOI22_X1 U20636 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17506), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17490), .ZN(n17461) );
  OAI21_X1 U20637 ( .B1(n17462), .B2(n17508), .A(n17461), .ZN(P3_U2774) );
  AOI22_X1 U20638 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17506), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17490), .ZN(n17463) );
  OAI21_X1 U20639 ( .B1(n17464), .B2(n17508), .A(n17463), .ZN(P3_U2775) );
  AOI22_X1 U20640 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17506), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17490), .ZN(n17465) );
  OAI21_X1 U20641 ( .B1(n17466), .B2(n17508), .A(n17465), .ZN(P3_U2776) );
  AOI22_X1 U20642 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17506), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17490), .ZN(n17467) );
  OAI21_X1 U20643 ( .B1(n17468), .B2(n17508), .A(n17467), .ZN(P3_U2777) );
  AOI22_X1 U20644 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17506), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17490), .ZN(n17469) );
  OAI21_X1 U20645 ( .B1(n17470), .B2(n17508), .A(n17469), .ZN(P3_U2778) );
  AOI22_X1 U20646 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17506), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17490), .ZN(n17471) );
  OAI21_X1 U20647 ( .B1(n17472), .B2(n17508), .A(n17471), .ZN(P3_U2779) );
  AOI22_X1 U20648 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17506), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17490), .ZN(n17473) );
  OAI21_X1 U20649 ( .B1(n17474), .B2(n17508), .A(n17473), .ZN(P3_U2780) );
  AOI22_X1 U20650 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17506), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17505), .ZN(n17475) );
  OAI21_X1 U20651 ( .B1(n17476), .B2(n17508), .A(n17475), .ZN(P3_U2781) );
  AOI22_X1 U20652 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17506), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17490), .ZN(n17477) );
  OAI21_X1 U20653 ( .B1(n17478), .B2(n17508), .A(n17477), .ZN(P3_U2782) );
  AOI22_X1 U20654 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17506), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17490), .ZN(n17479) );
  OAI21_X1 U20655 ( .B1(n20971), .B2(n17508), .A(n17479), .ZN(P3_U2783) );
  AOI22_X1 U20656 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17506), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17490), .ZN(n17480) );
  OAI21_X1 U20657 ( .B1(n17481), .B2(n17508), .A(n17480), .ZN(P3_U2784) );
  AOI22_X1 U20658 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17493), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17490), .ZN(n17482) );
  OAI21_X1 U20659 ( .B1(n20804), .B2(n17495), .A(n17482), .ZN(P3_U2785) );
  AOI22_X1 U20660 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17493), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17490), .ZN(n17483) );
  OAI21_X1 U20661 ( .B1(n18224), .B2(n17495), .A(n17483), .ZN(P3_U2786) );
  AOI22_X1 U20662 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17493), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17490), .ZN(n17484) );
  OAI21_X1 U20663 ( .B1(n18228), .B2(n17495), .A(n17484), .ZN(P3_U2787) );
  AOI22_X1 U20664 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17493), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17490), .ZN(n17485) );
  OAI21_X1 U20665 ( .B1(n18233), .B2(n17495), .A(n17485), .ZN(P3_U2788) );
  AOI22_X1 U20666 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17493), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17490), .ZN(n17486) );
  OAI21_X1 U20667 ( .B1(n18237), .B2(n17495), .A(n17486), .ZN(P3_U2789) );
  AOI22_X1 U20668 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17493), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17490), .ZN(n17487) );
  OAI21_X1 U20669 ( .B1(n18242), .B2(n17495), .A(n17487), .ZN(P3_U2790) );
  AOI22_X1 U20670 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17493), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17490), .ZN(n17488) );
  OAI21_X1 U20671 ( .B1(n17489), .B2(n17495), .A(n17488), .ZN(P3_U2791) );
  AOI22_X1 U20672 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17493), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17490), .ZN(n17491) );
  OAI21_X1 U20673 ( .B1(n17492), .B2(n17495), .A(n17491), .ZN(P3_U2792) );
  AOI22_X1 U20674 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17493), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17505), .ZN(n17494) );
  OAI21_X1 U20675 ( .B1(n17496), .B2(n17495), .A(n17494), .ZN(P3_U2793) );
  AOI22_X1 U20676 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17506), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17505), .ZN(n17497) );
  OAI21_X1 U20677 ( .B1(n17498), .B2(n17508), .A(n17497), .ZN(P3_U2794) );
  AOI22_X1 U20678 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17506), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17505), .ZN(n17499) );
  OAI21_X1 U20679 ( .B1(n17500), .B2(n17508), .A(n17499), .ZN(P3_U2795) );
  AOI22_X1 U20680 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17506), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17505), .ZN(n17501) );
  OAI21_X1 U20681 ( .B1(n17502), .B2(n17508), .A(n17501), .ZN(P3_U2796) );
  AOI22_X1 U20682 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17506), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17505), .ZN(n17503) );
  OAI21_X1 U20683 ( .B1(n17504), .B2(n17508), .A(n17503), .ZN(P3_U2797) );
  AOI22_X1 U20684 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17506), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17505), .ZN(n17507) );
  OAI21_X1 U20685 ( .B1(n17509), .B2(n17508), .A(n17507), .ZN(P3_U2798) );
  AOI21_X1 U20686 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17542), .A(
        n18721), .ZN(n17510) );
  AOI211_X1 U20687 ( .C1(n17829), .C2(n17511), .A(n17864), .B(n17510), .ZN(
        n17546) );
  OAI21_X1 U20688 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17665), .A(
        n17546), .ZN(n17531) );
  NOR2_X1 U20689 ( .A1(n17714), .A2(n17511), .ZN(n17533) );
  XOR2_X1 U20690 ( .A(n17512), .B(n17532), .Z(n17513) );
  AOI22_X1 U20691 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17531), .B1(
        n17533), .B2(n17513), .ZN(n17525) );
  AOI22_X1 U20692 ( .A1(n9726), .A2(P3_REIP_REG_28__SCAN_IN), .B1(n9758), .B2(
        n17514), .ZN(n17524) );
  AOI21_X1 U20693 ( .B1(n17517), .B2(n17516), .A(n17515), .ZN(n17520) );
  NOR2_X1 U20694 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17518), .ZN(
        n17519) );
  AOI22_X1 U20695 ( .A1(n17783), .A2(n17520), .B1(n17595), .B2(n17519), .ZN(
        n17523) );
  INV_X1 U20696 ( .A(n17521), .ZN(n17888) );
  AOI22_X1 U20697 ( .A1(n17869), .A2(n17888), .B1(n17784), .B2(n17887), .ZN(
        n17550) );
  NAND2_X1 U20698 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17550), .ZN(
        n17535) );
  OAI211_X1 U20699 ( .C1(n17869), .C2(n17784), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n17535), .ZN(n17522) );
  NAND4_X1 U20700 ( .A1(n17525), .A2(n17524), .A3(n17523), .A4(n17522), .ZN(
        P3_U2802) );
  NAND2_X1 U20701 ( .A1(n10102), .A2(n17527), .ZN(n17528) );
  XOR2_X1 U20702 ( .A(n17528), .B(n12900), .Z(n17898) );
  OAI22_X1 U20703 ( .A1(n18193), .A2(n18786), .B1(n9718), .B2(n17529), .ZN(
        n17530) );
  AOI221_X1 U20704 ( .B1(n17533), .B2(n17532), .C1(n17531), .C2(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(n17530), .ZN(n17538) );
  INV_X1 U20705 ( .A(n17534), .ZN(n17536) );
  OAI21_X1 U20706 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17536), .A(
        n17535), .ZN(n17537) );
  OAI211_X1 U20707 ( .C1(n17898), .C2(n17761), .A(n17538), .B(n17537), .ZN(
        P3_U2803) );
  NAND4_X1 U20708 ( .A1(n17539), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A4(n17658), .ZN(n17551) );
  INV_X1 U20709 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17899) );
  AOI21_X1 U20710 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17541), .A(
        n17540), .ZN(n17905) );
  INV_X1 U20711 ( .A(n17905), .ZN(n17548) );
  AOI21_X1 U20712 ( .B1(n17542), .B2(n18593), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17545) );
  OAI21_X1 U20713 ( .B1(n9758), .B2(n13068), .A(n17543), .ZN(n17544) );
  NAND2_X1 U20714 ( .A1(n9726), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17903) );
  OAI211_X1 U20715 ( .C1(n17546), .C2(n17545), .A(n17544), .B(n17903), .ZN(
        n17547) );
  AOI21_X1 U20716 ( .B1(n17783), .B2(n17548), .A(n17547), .ZN(n17549) );
  OAI221_X1 U20717 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17551), 
        .C1(n17899), .C2(n17550), .A(n17549), .ZN(P3_U2804) );
  AND2_X1 U20718 ( .A1(n17561), .A2(n18593), .ZN(n17584) );
  AOI211_X1 U20719 ( .C1(n17553), .C2(n17552), .A(n17864), .B(n17584), .ZN(
        n17592) );
  OAI21_X1 U20720 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17665), .A(
        n17592), .ZN(n17571) );
  AOI22_X1 U20721 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17571), .B1(
        n9758), .B2(n17554), .ZN(n17565) );
  XOR2_X1 U20722 ( .A(n17886), .B(n17555), .Z(n17918) );
  XOR2_X1 U20723 ( .A(n17886), .B(n17556), .Z(n17920) );
  OAI21_X1 U20724 ( .B1(n12900), .B2(n17558), .A(n17557), .ZN(n17559) );
  XOR2_X1 U20725 ( .A(n17559), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17916) );
  OAI22_X1 U20726 ( .A1(n17720), .A2(n17920), .B1(n17761), .B2(n17916), .ZN(
        n17560) );
  AOI21_X1 U20727 ( .B1(n17869), .B2(n17918), .A(n17560), .ZN(n17564) );
  NAND2_X1 U20728 ( .A1(n9726), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17914) );
  NOR2_X1 U20729 ( .A1(n17714), .A2(n17561), .ZN(n17573) );
  OAI211_X1 U20730 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17573), .B(n17562), .ZN(n17563) );
  NAND4_X1 U20731 ( .A1(n17565), .A2(n17564), .A3(n17914), .A4(n17563), .ZN(
        P3_U2805) );
  AOI21_X1 U20732 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17567), .A(
        n17566), .ZN(n17932) );
  INV_X1 U20733 ( .A(n17568), .ZN(n17569) );
  OAI22_X1 U20734 ( .A1(n18193), .A2(n18779), .B1(n9718), .B2(n17569), .ZN(
        n17570) );
  AOI221_X1 U20735 ( .B1(n17573), .B2(n17572), .C1(n17571), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17570), .ZN(n17579) );
  INV_X1 U20736 ( .A(n17924), .ZN(n17574) );
  OAI22_X1 U20737 ( .A1(n17926), .A2(n17881), .B1(n17574), .B2(n17720), .ZN(
        n17594) );
  NOR2_X1 U20738 ( .A1(n17575), .A2(n17686), .ZN(n17577) );
  AOI22_X1 U20739 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17594), .B1(
        n17577), .B2(n17576), .ZN(n17578) );
  OAI211_X1 U20740 ( .C1(n17932), .C2(n17761), .A(n17579), .B(n17578), .ZN(
        P3_U2806) );
  INV_X1 U20741 ( .A(n17580), .ZN(n17581) );
  OAI21_X1 U20742 ( .B1(n17651), .B2(n17581), .A(n17600), .ZN(n17582) );
  OAI211_X1 U20743 ( .C1(n17782), .C2(n17954), .A(n17599), .B(n17582), .ZN(
        n17583) );
  XOR2_X1 U20744 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n17583), .Z(
        n17938) );
  INV_X1 U20745 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17933) );
  AOI22_X1 U20746 ( .A1(n9726), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n17585), 
        .B2(n17584), .ZN(n17590) );
  NOR2_X1 U20747 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17665), .ZN(
        n17586) );
  AOI22_X1 U20748 ( .A1(n9758), .A2(n17588), .B1(n17587), .B2(n17586), .ZN(
        n17589) );
  OAI211_X1 U20749 ( .C1(n17592), .C2(n17591), .A(n17590), .B(n17589), .ZN(
        n17593) );
  AOI221_X1 U20750 ( .B1(n17595), .B2(n17933), .C1(n17594), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n17593), .ZN(n17596) );
  OAI21_X1 U20751 ( .B1(n17761), .B2(n17938), .A(n17596), .ZN(P3_U2807) );
  NOR2_X1 U20752 ( .A1(n17869), .A2(n17784), .ZN(n17634) );
  NAND2_X1 U20753 ( .A1(n17869), .A2(n18023), .ZN(n17700) );
  OAI21_X1 U20754 ( .B1(n17940), .B2(n17720), .A(n17700), .ZN(n17597) );
  INV_X1 U20755 ( .A(n17597), .ZN(n17685) );
  OAI21_X1 U20756 ( .B1(n17944), .B2(n17634), .A(n17685), .ZN(n17598) );
  INV_X1 U20757 ( .A(n17598), .ZN(n17624) );
  AOI221_X1 U20758 ( .B1(n17601), .B2(n17600), .C1(n17619), .C2(n17600), .A(
        n17625), .ZN(n17602) );
  XOR2_X1 U20759 ( .A(n17602), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(
        n17939) );
  OAI21_X1 U20760 ( .B1(n17603), .B2(n18721), .A(n17877), .ZN(n17604) );
  AOI21_X1 U20761 ( .B1(n17829), .B2(n17606), .A(n17604), .ZN(n17631) );
  OAI21_X1 U20762 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17665), .A(
        n17631), .ZN(n17616) );
  AOI22_X1 U20763 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n17616), .B1(
        n9758), .B2(n17605), .ZN(n17609) );
  NOR2_X1 U20764 ( .A1(n17714), .A2(n17606), .ZN(n17618) );
  OAI211_X1 U20765 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17618), .B(n17607), .ZN(n17608) );
  OAI211_X1 U20766 ( .C1(n18775), .C2(n18193), .A(n17609), .B(n17608), .ZN(
        n17610) );
  AOI21_X1 U20767 ( .B1(n17783), .B2(n17939), .A(n17610), .ZN(n17611) );
  OAI221_X1 U20768 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17612), 
        .C1(n17954), .C2(n17624), .A(n17611), .ZN(P3_U2808) );
  INV_X1 U20769 ( .A(n17613), .ZN(n17614) );
  OAI22_X1 U20770 ( .A1(n18193), .A2(n18773), .B1(n9718), .B2(n17614), .ZN(
        n17615) );
  AOI221_X1 U20771 ( .B1(n17618), .B2(n17617), .C1(n17616), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17615), .ZN(n17623) );
  INV_X1 U20772 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17963) );
  NOR3_X1 U20773 ( .A1(n17963), .A2(n12900), .A3(n17619), .ZN(n17637) );
  AOI22_X1 U20774 ( .A1(n17961), .A2(n17637), .B1(n17651), .B2(n17620), .ZN(
        n17621) );
  XOR2_X1 U20775 ( .A(n17946), .B(n17621), .Z(n17966) );
  NOR2_X1 U20776 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17947), .ZN(
        n17965) );
  NAND2_X1 U20777 ( .A1(n17989), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17956) );
  NOR2_X1 U20778 ( .A1(n17686), .A2(n17956), .ZN(n17647) );
  AOI22_X1 U20779 ( .A1(n17783), .A2(n17966), .B1(n17965), .B2(n17647), .ZN(
        n17622) );
  OAI211_X1 U20780 ( .C1(n17624), .C2(n17946), .A(n17623), .B(n17622), .ZN(
        P3_U2809) );
  INV_X1 U20781 ( .A(n17637), .ZN(n17626) );
  AOI221_X1 U20782 ( .B1(n17980), .B2(n17627), .C1(n17626), .C2(n17627), .A(
        n17625), .ZN(n17628) );
  XNOR2_X1 U20783 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B(n17628), .ZN(
        n17978) );
  AOI21_X1 U20784 ( .B1(n17629), .B2(n18593), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17630) );
  OAI22_X1 U20785 ( .A1(n17631), .A2(n17630), .B1(n18193), .B2(n18771), .ZN(
        n17632) );
  AOI221_X1 U20786 ( .B1(n9758), .B2(n17633), .C1(n13068), .C2(n17633), .A(
        n17632), .ZN(n17636) );
  NOR2_X1 U20787 ( .A1(n17980), .A2(n17956), .ZN(n17970) );
  OAI21_X1 U20788 ( .B1(n17634), .B2(n17970), .A(n17685), .ZN(n17646) );
  NOR2_X1 U20789 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17980), .ZN(
        n17969) );
  AOI22_X1 U20790 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17646), .B1(
        n17969), .B2(n17647), .ZN(n17635) );
  OAI211_X1 U20791 ( .C1(n17761), .C2(n17978), .A(n17636), .B(n17635), .ZN(
        P3_U2810) );
  AOI21_X1 U20792 ( .B1(n17651), .B2(n17649), .A(n17637), .ZN(n17638) );
  XOR2_X1 U20793 ( .A(n17638), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Z(
        n17984) );
  AOI21_X1 U20794 ( .B1(n17829), .B2(n17640), .A(n17864), .ZN(n17672) );
  OAI21_X1 U20795 ( .B1(n17639), .B2(n18721), .A(n17672), .ZN(n17654) );
  NOR2_X1 U20796 ( .A1(n18193), .A2(n18769), .ZN(n17979) );
  AOI21_X1 U20797 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17654), .A(
        n17979), .ZN(n17643) );
  NOR2_X1 U20798 ( .A1(n17714), .A2(n17640), .ZN(n17656) );
  OAI211_X1 U20799 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17656), .B(n17641), .ZN(n17642) );
  OAI211_X1 U20800 ( .C1(n9718), .C2(n17644), .A(n17643), .B(n17642), .ZN(
        n17645) );
  AOI221_X1 U20801 ( .B1(n17647), .B2(n17980), .C1(n17646), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n17645), .ZN(n17648) );
  OAI21_X1 U20802 ( .B1(n17984), .B2(n17761), .A(n17648), .ZN(P3_U2811) );
  AOI21_X1 U20803 ( .B1(n17782), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17649), .ZN(n17650) );
  XNOR2_X1 U20804 ( .A(n17651), .B(n17650), .ZN(n17999) );
  NAND2_X1 U20805 ( .A1(n9726), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17997) );
  OAI21_X1 U20806 ( .B1(n9718), .B2(n17652), .A(n17997), .ZN(n17653) );
  AOI221_X1 U20807 ( .B1(n17656), .B2(n17655), .C1(n17654), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17653), .ZN(n17660) );
  OAI21_X1 U20808 ( .B1(n17989), .B2(n17686), .A(n17685), .ZN(n17669) );
  NOR2_X1 U20809 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17657), .ZN(
        n17995) );
  AOI22_X1 U20810 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17669), .B1(
        n17658), .B2(n17995), .ZN(n17659) );
  OAI211_X1 U20811 ( .C1(n17761), .C2(n17999), .A(n17660), .B(n17659), .ZN(
        P3_U2812) );
  AOI21_X1 U20812 ( .B1(n17661), .B2(n18593), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17673) );
  OAI21_X1 U20813 ( .B1(n18011), .B2(n17686), .A(n21020), .ZN(n17668) );
  INV_X1 U20814 ( .A(n17662), .ZN(n17663) );
  AOI21_X1 U20815 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17664), .A(
        n17663), .ZN(n18004) );
  OAI22_X1 U20816 ( .A1(n18004), .A2(n17761), .B1(n17861), .B2(n17666), .ZN(
        n17667) );
  AOI21_X1 U20817 ( .B1(n17669), .B2(n17668), .A(n17667), .ZN(n17671) );
  NAND2_X1 U20818 ( .A1(n9726), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n17670) );
  OAI211_X1 U20819 ( .C1(n17673), .C2(n17672), .A(n17671), .B(n17670), .ZN(
        P3_U2813) );
  OAI21_X1 U20820 ( .B1(n12900), .B2(n17675), .A(n17674), .ZN(n17676) );
  XOR2_X1 U20821 ( .A(n17676), .B(n18011), .Z(n18013) );
  AOI21_X1 U20822 ( .B1(n17829), .B2(n17679), .A(n17864), .ZN(n17702) );
  OAI21_X1 U20823 ( .B1(n17677), .B2(n18721), .A(n17702), .ZN(n17689) );
  AOI22_X1 U20824 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17689), .B1(
        n9758), .B2(n17678), .ZN(n17682) );
  NOR2_X1 U20825 ( .A1(n17714), .A2(n17679), .ZN(n17691) );
  OAI211_X1 U20826 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17691), .B(n17680), .ZN(n17681) );
  OAI211_X1 U20827 ( .C1(n18763), .C2(n18193), .A(n17682), .B(n17681), .ZN(
        n17683) );
  AOI21_X1 U20828 ( .B1(n17783), .B2(n18013), .A(n17683), .ZN(n17684) );
  OAI221_X1 U20829 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17686), 
        .C1(n18011), .C2(n17685), .A(n17684), .ZN(P3_U2814) );
  NOR2_X1 U20830 ( .A1(n17705), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n18022) );
  OAI22_X1 U20831 ( .A1(n18193), .A2(n18761), .B1(n9718), .B2(n17687), .ZN(
        n17688) );
  AOI221_X1 U20832 ( .B1(n17691), .B2(n17690), .C1(n17689), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17688), .ZN(n17699) );
  INV_X1 U20833 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18062) );
  NOR2_X1 U20834 ( .A1(n18059), .A2(n17692), .ZN(n17722) );
  NOR2_X1 U20835 ( .A1(n20828), .A2(n18034), .ZN(n17694) );
  NOR2_X1 U20836 ( .A1(n17782), .A2(n10104), .ZN(n17762) );
  NAND2_X1 U20837 ( .A1(n17693), .A2(n17762), .ZN(n17738) );
  NOR2_X1 U20838 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17738), .ZN(
        n17727) );
  AOI22_X1 U20839 ( .A1(n17722), .A2(n17694), .B1(n17727), .B2(n20828), .ZN(
        n17695) );
  AOI221_X1 U20840 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18062), 
        .C1(n12900), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(n17695), .ZN(
        n17696) );
  XOR2_X1 U20841 ( .A(n17696), .B(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .Z(
        n18025) );
  NOR2_X1 U20842 ( .A1(n17940), .A2(n17720), .ZN(n17697) );
  NAND2_X1 U20843 ( .A1(n18073), .A2(n18009), .ZN(n17701) );
  NAND2_X1 U20844 ( .A1(n18016), .A2(n17701), .ZN(n18020) );
  AOI22_X1 U20845 ( .A1(n17783), .A2(n18025), .B1(n17697), .B2(n18020), .ZN(
        n17698) );
  OAI211_X1 U20846 ( .C1(n18022), .C2(n17700), .A(n17699), .B(n17698), .ZN(
        P3_U2815) );
  NOR2_X1 U20847 ( .A1(n17710), .A2(n13073), .ZN(n18051) );
  OAI221_X1 U20848 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18051), .A(n17701), .ZN(
        n18043) );
  OR2_X1 U20849 ( .A1(n17713), .A2(n18454), .ZN(n17742) );
  AOI221_X1 U20850 ( .B1(n17715), .B2(n9987), .C1(n17742), .C2(n9987), .A(
        n17702), .ZN(n17703) );
  INV_X1 U20851 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18760) );
  NOR2_X1 U20852 ( .A1(n18193), .A2(n18760), .ZN(n18036) );
  AOI211_X1 U20853 ( .C1(n17704), .C2(n17871), .A(n17703), .B(n18036), .ZN(
        n17709) );
  AOI221_X1 U20854 ( .B1(n20828), .B2(n18034), .C1(n18047), .C2(n18034), .A(
        n17705), .ZN(n18040) );
  NAND2_X1 U20855 ( .A1(n17782), .A2(n18073), .ZN(n17739) );
  INV_X1 U20856 ( .A(n17739), .ZN(n17763) );
  NOR2_X1 U20857 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17706) );
  AOI22_X1 U20858 ( .A1(n18029), .A2(n17763), .B1(n17706), .B2(n17727), .ZN(
        n17707) );
  XOR2_X1 U20859 ( .A(n18034), .B(n17707), .Z(n18039) );
  AOI22_X1 U20860 ( .A1(n17869), .A2(n18040), .B1(n17783), .B2(n18039), .ZN(
        n17708) );
  OAI211_X1 U20861 ( .C1(n17720), .C2(n18043), .A(n17709), .B(n17708), .ZN(
        P3_U2816) );
  NAND2_X1 U20862 ( .A1(n9930), .A2(n20828), .ZN(n18056) );
  NAND2_X1 U20863 ( .A1(n17829), .A2(n17713), .ZN(n17711) );
  OAI211_X1 U20864 ( .C1(n17712), .C2(n18721), .A(n17711), .B(n17877), .ZN(
        n17733) );
  NOR2_X1 U20865 ( .A1(n17714), .A2(n17713), .ZN(n17732) );
  OAI211_X1 U20866 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17732), .B(n17715), .ZN(n17717) );
  NAND2_X1 U20867 ( .A1(n9726), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17716) );
  OAI211_X1 U20868 ( .C1(n9718), .C2(n17718), .A(n17717), .B(n17716), .ZN(
        n17719) );
  AOI21_X1 U20869 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17733), .A(
        n17719), .ZN(n17726) );
  OAI22_X1 U20870 ( .A1(n17721), .A2(n17881), .B1(n18051), .B2(n17720), .ZN(
        n17734) );
  NOR2_X1 U20871 ( .A1(n18062), .A2(n12900), .ZN(n17723) );
  OAI22_X1 U20872 ( .A1(n17727), .A2(n17723), .B1(n17722), .B2(n18062), .ZN(
        n17724) );
  XOR2_X1 U20873 ( .A(n20828), .B(n17724), .Z(n18045) );
  AOI22_X1 U20874 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17734), .B1(
        n17783), .B2(n18045), .ZN(n17725) );
  OAI211_X1 U20875 ( .C1(n17773), .C2(n18056), .A(n17726), .B(n17725), .ZN(
        P3_U2817) );
  AOI21_X1 U20876 ( .B1(n17763), .B2(n18046), .A(n17727), .ZN(n17728) );
  XOR2_X1 U20877 ( .A(n17728), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n18066) );
  INV_X1 U20878 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17731) );
  INV_X1 U20879 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18755) );
  OAI22_X1 U20880 ( .A1(n18193), .A2(n18755), .B1(n9718), .B2(n17729), .ZN(
        n17730) );
  AOI221_X1 U20881 ( .B1(n17733), .B2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C1(
        n17732), .C2(n17731), .A(n17730), .ZN(n17737) );
  OAI21_X1 U20882 ( .B1(n18059), .B2(n17773), .A(n18062), .ZN(n17735) );
  NAND2_X1 U20883 ( .A1(n17735), .A2(n17734), .ZN(n17736) );
  OAI211_X1 U20884 ( .C1(n18066), .C2(n17761), .A(n17737), .B(n17736), .ZN(
        P3_U2818) );
  OR2_X1 U20885 ( .A1(n18076), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18081) );
  OAI21_X1 U20886 ( .B1(n18076), .B2(n17739), .A(n17738), .ZN(n17740) );
  XOR2_X1 U20887 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n17740), .Z(
        n18067) );
  NAND2_X1 U20888 ( .A1(n17777), .A2(n18593), .ZN(n17789) );
  NOR2_X1 U20889 ( .A1(n17741), .A2(n17789), .ZN(n17754) );
  OAI211_X1 U20890 ( .C1(n17754), .C2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n17872), .B(n17742), .ZN(n17744) );
  NAND2_X1 U20891 ( .A1(n9726), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n17743) );
  OAI211_X1 U20892 ( .C1(n17861), .C2(n17745), .A(n17744), .B(n17743), .ZN(
        n17746) );
  AOI21_X1 U20893 ( .B1(n17783), .B2(n18067), .A(n17746), .ZN(n17749) );
  NOR2_X1 U20894 ( .A1(n17747), .A2(n17773), .ZN(n17757) );
  AOI22_X1 U20895 ( .A1(n13073), .A2(n17784), .B1(n17869), .B2(n18070), .ZN(
        n17772) );
  INV_X1 U20896 ( .A(n17772), .ZN(n17758) );
  OAI21_X1 U20897 ( .B1(n17757), .B2(n17758), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17748) );
  OAI211_X1 U20898 ( .C1(n17773), .C2(n18081), .A(n17749), .B(n17748), .ZN(
        P3_U2819) );
  AOI22_X1 U20899 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17763), .B1(
        n17762), .B2(n18100), .ZN(n17750) );
  XOR2_X1 U20900 ( .A(n17750), .B(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .Z(
        n18091) );
  NAND2_X1 U20901 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17776) );
  NOR3_X1 U20902 ( .A1(n17776), .A2(n17751), .A3(n17789), .ZN(n17768) );
  AOI21_X1 U20903 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n17872), .A(
        n17768), .ZN(n17753) );
  OAI22_X1 U20904 ( .A1(n17754), .A2(n17753), .B1(n17861), .B2(n17752), .ZN(
        n17755) );
  AOI21_X1 U20905 ( .B1(n9726), .B2(P3_REIP_REG_10__SCAN_IN), .A(n17755), .ZN(
        n17760) );
  AOI22_X1 U20906 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17758), .B1(
        n17757), .B2(n17756), .ZN(n17759) );
  OAI211_X1 U20907 ( .C1(n18091), .C2(n17761), .A(n17760), .B(n17759), .ZN(
        P3_U2820) );
  NOR2_X1 U20908 ( .A1(n17763), .A2(n17762), .ZN(n17764) );
  XOR2_X1 U20909 ( .A(n17764), .B(n18100), .Z(n18097) );
  NOR2_X1 U20910 ( .A1(n18193), .A2(n18751), .ZN(n17770) );
  NOR2_X1 U20911 ( .A1(n17776), .A2(n17789), .ZN(n17765) );
  AOI21_X1 U20912 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17872), .A(
        n17765), .ZN(n17767) );
  OAI22_X1 U20913 ( .A1(n17768), .A2(n17767), .B1(n17861), .B2(n17766), .ZN(
        n17769) );
  AOI211_X1 U20914 ( .C1(n17783), .C2(n18097), .A(n17770), .B(n17769), .ZN(
        n17771) );
  OAI221_X1 U20915 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17773), .C1(
        n18100), .C2(n17772), .A(n17771), .ZN(P3_U2821) );
  OAI21_X1 U20916 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17775), .A(
        n17774), .ZN(n18117) );
  OAI21_X1 U20917 ( .B1(n17777), .B2(n17845), .A(n17877), .ZN(n17790) );
  NOR2_X1 U20918 ( .A1(n18193), .A2(n20834), .ZN(n18108) );
  OAI211_X1 U20919 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n17777), .B(n17776), .ZN(n17778)
         );
  OAI22_X1 U20920 ( .A1(n17861), .A2(n17779), .B1(n18454), .B2(n17778), .ZN(
        n17780) );
  AOI211_X1 U20921 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17790), .A(
        n18108), .B(n17780), .ZN(n17786) );
  OAI21_X1 U20922 ( .B1(n17782), .B2(n18114), .A(n17781), .ZN(n18111) );
  AOI22_X1 U20923 ( .A1(n17784), .A2(n18114), .B1(n17783), .B2(n18111), .ZN(
        n17785) );
  OAI211_X1 U20924 ( .C1(n17881), .C2(n18117), .A(n17786), .B(n17785), .ZN(
        P3_U2822) );
  OAI21_X1 U20925 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17788), .A(
        n17787), .ZN(n18120) );
  INV_X1 U20926 ( .A(n17789), .ZN(n17792) );
  NOR2_X1 U20927 ( .A1(n18193), .A2(n18749), .ZN(n18119) );
  AOI221_X1 U20928 ( .B1(n17792), .B2(n17791), .C1(n17790), .C2(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(n18119), .ZN(n17799) );
  AOI21_X1 U20929 ( .B1(n17795), .B2(n17794), .A(n17793), .ZN(n17796) );
  XOR2_X1 U20930 ( .A(n17796), .B(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .Z(
        n18122) );
  AOI22_X1 U20931 ( .A1(n17869), .A2(n18122), .B1(n17797), .B2(n17871), .ZN(
        n17798) );
  OAI211_X1 U20932 ( .C1(n17880), .C2(n18120), .A(n17799), .B(n17798), .ZN(
        P3_U2823) );
  OAI21_X1 U20933 ( .B1(n18454), .B2(n17800), .A(n17872), .ZN(n17826) );
  NOR2_X1 U20934 ( .A1(n17800), .A2(n18454), .ZN(n17809) );
  OAI21_X1 U20935 ( .B1(n17803), .B2(n17802), .A(n17801), .ZN(n18129) );
  OAI22_X1 U20936 ( .A1(n17880), .A2(n18129), .B1(n18193), .B2(n18747), .ZN(
        n17808) );
  OAI21_X1 U20937 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n17805), .A(
        n17804), .ZN(n18134) );
  OAI22_X1 U20938 ( .A1(n17861), .A2(n17806), .B1(n17881), .B2(n18134), .ZN(
        n17807) );
  AOI211_X1 U20939 ( .C1(n17809), .C2(n17811), .A(n17808), .B(n17807), .ZN(
        n17810) );
  OAI21_X1 U20940 ( .B1(n17811), .B2(n17826), .A(n17810), .ZN(P3_U2824) );
  AOI21_X1 U20941 ( .B1(n17812), .B2(n17877), .A(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17827) );
  INV_X1 U20942 ( .A(n17813), .ZN(n17814) );
  AOI21_X1 U20943 ( .B1(n17816), .B2(n17815), .A(n17814), .ZN(n17817) );
  XOR2_X1 U20944 ( .A(n17817), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(
        n18135) );
  AOI22_X1 U20945 ( .A1(n17818), .A2(n18135), .B1(n9726), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17825) );
  AOI21_X1 U20946 ( .B1(n17821), .B2(n17820), .A(n17819), .ZN(n17822) );
  XOR2_X1 U20947 ( .A(n17822), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(
        n18137) );
  AOI22_X1 U20948 ( .A1(n17869), .A2(n18137), .B1(n17823), .B2(n17871), .ZN(
        n17824) );
  OAI211_X1 U20949 ( .C1(n17827), .C2(n17826), .A(n17825), .B(n17824), .ZN(
        P3_U2825) );
  AOI21_X1 U20950 ( .B1(n17829), .B2(n17828), .A(n17864), .ZN(n17849) );
  OAI21_X1 U20951 ( .B1(n17832), .B2(n17831), .A(n17830), .ZN(n18149) );
  OAI22_X1 U20952 ( .A1(n17881), .A2(n18149), .B1(n18193), .B2(n18744), .ZN(
        n17838) );
  OAI21_X1 U20953 ( .B1(n17835), .B2(n17834), .A(n17833), .ZN(n18155) );
  OAI22_X1 U20954 ( .A1(n17861), .A2(n17836), .B1(n17880), .B2(n18155), .ZN(
        n17837) );
  AOI211_X1 U20955 ( .C1(n18593), .C2(n17839), .A(n17838), .B(n17837), .ZN(
        n17840) );
  OAI21_X1 U20956 ( .B1(n17849), .B2(n17841), .A(n17840), .ZN(P3_U2826) );
  OAI21_X1 U20957 ( .B1(n17844), .B2(n17843), .A(n17842), .ZN(n18159) );
  NOR4_X1 U20958 ( .A1(n17864), .A2(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        n17863), .A4(n17845), .ZN(n17851) );
  OAI21_X1 U20959 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n17847), .A(
        n17846), .ZN(n18158) );
  OAI22_X1 U20960 ( .A1(n17849), .A2(n17848), .B1(n17880), .B2(n18158), .ZN(
        n17850) );
  AOI211_X1 U20961 ( .C1(n17852), .C2(n17871), .A(n17851), .B(n17850), .ZN(
        n17853) );
  NAND2_X1 U20962 ( .A1(n9726), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18162) );
  OAI211_X1 U20963 ( .C1(n17881), .C2(n18159), .A(n17853), .B(n18162), .ZN(
        P3_U2827) );
  OAI21_X1 U20964 ( .B1(n17856), .B2(n17855), .A(n17854), .ZN(n18179) );
  OAI21_X1 U20965 ( .B1(n17859), .B2(n17858), .A(n17857), .ZN(n18175) );
  OAI22_X1 U20966 ( .A1(n17861), .A2(n17860), .B1(n17880), .B2(n18175), .ZN(
        n17862) );
  AOI221_X1 U20967 ( .B1(n17864), .B2(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .C1(
        n18593), .C2(n17863), .A(n17862), .ZN(n17865) );
  NAND2_X1 U20968 ( .A1(n9726), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18177) );
  OAI211_X1 U20969 ( .C1(n17881), .C2(n18179), .A(n17865), .B(n18177), .ZN(
        P3_U2828) );
  OAI21_X1 U20970 ( .B1(n17867), .B2(n17875), .A(n17866), .ZN(n18190) );
  NAND2_X1 U20971 ( .A1(n21021), .A2(n17876), .ZN(n17868) );
  XNOR2_X1 U20972 ( .A(n17868), .B(n17867), .ZN(n18183) );
  AOI22_X1 U20973 ( .A1(n17869), .A2(n18183), .B1(n9726), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17874) );
  AOI22_X1 U20974 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17872), .B1(
        n17871), .B2(n17870), .ZN(n17873) );
  OAI211_X1 U20975 ( .C1(n17880), .C2(n18190), .A(n17874), .B(n17873), .ZN(
        P3_U2829) );
  AOI21_X1 U20976 ( .B1(n17876), .B2(n21021), .A(n17875), .ZN(n18199) );
  INV_X1 U20977 ( .A(n18199), .ZN(n18197) );
  NAND3_X1 U20978 ( .A1(n18813), .A2(n18721), .A3(n17877), .ZN(n17878) );
  AOI22_X1 U20979 ( .A1(n9726), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17878), .ZN(n17879) );
  OAI221_X1 U20980 ( .B1(n18199), .B2(n17881), .C1(n18197), .C2(n17880), .A(
        n17879), .ZN(P3_U2830) );
  NAND2_X1 U20981 ( .A1(n9726), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17897) );
  NOR2_X1 U20982 ( .A1(n17909), .A2(n17934), .ZN(n17902) );
  NOR2_X1 U20983 ( .A1(n18647), .A2(n18654), .ZN(n18147) );
  INV_X1 U20984 ( .A(n18147), .ZN(n18166) );
  INV_X1 U20985 ( .A(n17882), .ZN(n17884) );
  OAI21_X1 U20986 ( .B1(n17954), .B2(n18654), .A(n17883), .ZN(n17948) );
  AOI21_X1 U20987 ( .B1(n17884), .B2(n17948), .A(n18147), .ZN(n17923) );
  AOI21_X1 U20988 ( .B1(n18166), .B2(n17909), .A(n17923), .ZN(n17907) );
  AOI22_X1 U20989 ( .A1(n18647), .A2(n17886), .B1(n18654), .B2(n17885), .ZN(
        n17891) );
  AOI22_X1 U20990 ( .A1(n18069), .A2(n17888), .B1(n17943), .B2(n17887), .ZN(
        n17890) );
  OAI22_X1 U20991 ( .A1(n17893), .A2(n18185), .B1(n17892), .B2(n18165), .ZN(
        n17894) );
  OAI221_X1 U20992 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17895), 
        .C1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n17902), .A(n17894), .ZN(
        n17896) );
  OAI211_X1 U20993 ( .C1(n17898), .C2(n18090), .A(n17897), .B(n17896), .ZN(
        P3_U2835) );
  OAI22_X1 U20994 ( .A1(n18185), .A2(n17900), .B1(n18165), .B2(n17899), .ZN(
        n17901) );
  OAI221_X1 U20995 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n17902), .A(n17901), .ZN(
        n17904) );
  OAI211_X1 U20996 ( .C1(n17905), .C2(n18090), .A(n17904), .B(n17903), .ZN(
        P3_U2836) );
  NOR2_X1 U20997 ( .A1(n17906), .A2(n17909), .ZN(n17912) );
  INV_X1 U20998 ( .A(n17907), .ZN(n17908) );
  AOI221_X1 U20999 ( .B1(n17909), .B2(n18145), .C1(n17927), .C2(n18145), .A(
        n17908), .ZN(n17910) );
  INV_X1 U21000 ( .A(n17910), .ZN(n17911) );
  MUX2_X1 U21001 ( .A(n17912), .B(n17911), .S(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(n17913) );
  AOI22_X1 U21002 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n18187), .B1(
        n18191), .B2(n17913), .ZN(n17915) );
  OAI211_X1 U21003 ( .C1(n17916), .C2(n18090), .A(n17915), .B(n17914), .ZN(
        n17917) );
  AOI21_X1 U21004 ( .B1(n18184), .B2(n17918), .A(n17917), .ZN(n17919) );
  OAI21_X1 U21005 ( .B1(n18044), .B2(n17920), .A(n17919), .ZN(P3_U2837) );
  NOR4_X1 U21006 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17964), .A3(
        n17921), .A4(n18185), .ZN(n17922) );
  AOI21_X1 U21007 ( .B1(P3_REIP_REG_24__SCAN_IN), .B2(n9726), .A(n17922), .ZN(
        n17931) );
  AOI211_X1 U21008 ( .C1(n17943), .C2(n17924), .A(n17923), .B(n18187), .ZN(
        n17925) );
  OAI21_X1 U21009 ( .B1(n17926), .B2(n18684), .A(n17925), .ZN(n17929) );
  AOI211_X1 U21010 ( .C1(n18145), .C2(n17927), .A(n17933), .B(n17929), .ZN(
        n17928) );
  NOR2_X1 U21011 ( .A1(n9726), .A2(n17928), .ZN(n17936) );
  OAI211_X1 U21012 ( .C1(n18107), .C2(n17929), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17936), .ZN(n17930) );
  OAI211_X1 U21013 ( .C1(n17932), .C2(n18090), .A(n17931), .B(n17930), .ZN(
        P3_U2838) );
  OAI21_X1 U21014 ( .B1(n18187), .B2(n17934), .A(n17933), .ZN(n17935) );
  AOI22_X1 U21015 ( .A1(n9726), .A2(P3_REIP_REG_23__SCAN_IN), .B1(n17936), 
        .B2(n17935), .ZN(n17937) );
  OAI21_X1 U21016 ( .B1(n18090), .B2(n17938), .A(n17937), .ZN(P3_U2839) );
  AOI22_X1 U21017 ( .A1(n9726), .A2(P3_REIP_REG_22__SCAN_IN), .B1(n9717), .B2(
        n17939), .ZN(n17953) );
  NOR2_X1 U21018 ( .A1(n17940), .A2(n18072), .ZN(n18021) );
  AOI21_X1 U21019 ( .B1(n18069), .B2(n18023), .A(n18021), .ZN(n17958) );
  OAI21_X1 U21020 ( .B1(n17963), .B2(n17941), .A(n18145), .ZN(n17942) );
  OAI221_X1 U21021 ( .B1(n18656), .B2(n17986), .C1(n18656), .C2(n17970), .A(
        n17942), .ZN(n17971) );
  NOR2_X1 U21022 ( .A1(n18069), .A2(n17943), .ZN(n17988) );
  OAI22_X1 U21023 ( .A1(n18656), .A2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n17944), .B2(n17988), .ZN(n17945) );
  NOR2_X1 U21024 ( .A1(n17971), .A2(n17945), .ZN(n17960) );
  INV_X1 U21025 ( .A(n18052), .ZN(n18082) );
  AOI22_X1 U21026 ( .A1(n18145), .A2(n17947), .B1(n18082), .B2(n17946), .ZN(
        n17949) );
  NAND4_X1 U21027 ( .A1(n17958), .A2(n17960), .A3(n17949), .A4(n17948), .ZN(
        n17950) );
  OAI211_X1 U21028 ( .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17951), .A(
        n18191), .B(n17950), .ZN(n17952) );
  OAI211_X1 U21029 ( .C1(n18165), .C2(n17954), .A(n17953), .B(n17952), .ZN(
        P3_U2840) );
  NOR2_X1 U21030 ( .A1(n18145), .A2(n18654), .ZN(n18186) );
  INV_X1 U21031 ( .A(n17994), .ZN(n17955) );
  NOR2_X1 U21032 ( .A1(n21021), .A2(n18006), .ZN(n18093) );
  NAND2_X1 U21033 ( .A1(n17955), .A2(n18093), .ZN(n18007) );
  OAI21_X1 U21034 ( .B1(n17956), .B2(n18007), .A(n18654), .ZN(n17957) );
  INV_X1 U21035 ( .A(n17957), .ZN(n17959) );
  NAND2_X1 U21036 ( .A1(n18191), .A2(n17958), .ZN(n18010) );
  NOR2_X1 U21037 ( .A1(n17959), .A2(n18010), .ZN(n17973) );
  OAI211_X1 U21038 ( .C1(n17961), .C2(n18186), .A(n17973), .B(n17960), .ZN(
        n17962) );
  NAND2_X1 U21039 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17962), .ZN(
        n17968) );
  NOR3_X1 U21040 ( .A1(n17964), .A2(n18185), .A3(n17963), .ZN(n17981) );
  AOI22_X1 U21041 ( .A1(n9717), .A2(n17966), .B1(n17981), .B2(n17965), .ZN(
        n17967) );
  OAI221_X1 U21042 ( .B1(n9726), .B2(n17968), .C1(n18193), .C2(n18773), .A(
        n17967), .ZN(P3_U2841) );
  AOI22_X1 U21043 ( .A1(n9726), .A2(P3_REIP_REG_20__SCAN_IN), .B1(n17981), 
        .B2(n17969), .ZN(n17977) );
  INV_X1 U21044 ( .A(n17970), .ZN(n17972) );
  INV_X1 U21045 ( .A(n17988), .ZN(n18075) );
  AOI21_X1 U21046 ( .B1(n17972), .B2(n18075), .A(n17971), .ZN(n17974) );
  AOI21_X1 U21047 ( .B1(n17974), .B2(n17973), .A(n9726), .ZN(n17982) );
  NOR3_X1 U21048 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18186), .A3(
        n18865), .ZN(n17975) );
  OAI21_X1 U21049 ( .B1(n17982), .B2(n17975), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17976) );
  OAI211_X1 U21050 ( .C1(n17978), .C2(n18090), .A(n17977), .B(n17976), .ZN(
        P3_U2842) );
  AOI221_X1 U21051 ( .B1(n17982), .B2(P3_INSTADDRPOINTER_REG_19__SCAN_IN), 
        .C1(n17981), .C2(n17980), .A(n17979), .ZN(n17983) );
  OAI21_X1 U21052 ( .B1(n17984), .B2(n18090), .A(n17983), .ZN(P3_U2843) );
  NOR2_X1 U21053 ( .A1(n18094), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18167) );
  INV_X1 U21054 ( .A(n18167), .ZN(n17985) );
  NAND3_X1 U21055 ( .A1(n17986), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n17985), .ZN(n17991) );
  OAI22_X1 U21056 ( .A1(n17989), .A2(n17988), .B1(n17987), .B2(n18685), .ZN(
        n17990) );
  AOI211_X1 U21057 ( .C1(n18166), .C2(n17991), .A(n18010), .B(n17990), .ZN(
        n18000) );
  AOI221_X1 U21058 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n18000), 
        .C1(n18147), .C2(n18000), .A(n9726), .ZN(n17996) );
  INV_X1 U21059 ( .A(n18144), .ZN(n17992) );
  INV_X1 U21060 ( .A(n18103), .ZN(n18146) );
  AOI22_X1 U21061 ( .A1(n18145), .A2(n17992), .B1(n18171), .B2(n18146), .ZN(
        n18157) );
  NOR2_X1 U21062 ( .A1(n18157), .A2(n17993), .ZN(n18058) );
  OAI21_X1 U21063 ( .B1(n18058), .B2(n18057), .A(n18191), .ZN(n18101) );
  NOR2_X1 U21064 ( .A1(n17994), .A2(n18101), .ZN(n18012) );
  AOI22_X1 U21065 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17996), .B1(
        n18012), .B2(n17995), .ZN(n17998) );
  OAI211_X1 U21066 ( .C1(n18090), .C2(n17999), .A(n17998), .B(n17997), .ZN(
        P3_U2844) );
  NOR2_X1 U21067 ( .A1(n9726), .A2(n18000), .ZN(n18001) );
  AOI22_X1 U21068 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18001), .B1(
        n9726), .B2(P3_REIP_REG_17__SCAN_IN), .ZN(n18003) );
  NAND3_X1 U21069 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n18012), .A3(
        n21020), .ZN(n18002) );
  OAI211_X1 U21070 ( .C1(n18004), .C2(n18090), .A(n18003), .B(n18002), .ZN(
        P3_U2845) );
  NOR2_X1 U21071 ( .A1(n18005), .A2(n18685), .ZN(n18068) );
  NAND2_X1 U21072 ( .A1(n18647), .A2(n18006), .ZN(n18092) );
  INV_X1 U21073 ( .A(n18092), .ZN(n18083) );
  NOR2_X1 U21074 ( .A1(n18068), .A2(n18083), .ZN(n18031) );
  OAI21_X1 U21075 ( .B1(n18016), .B2(n18654), .A(n18007), .ZN(n18008) );
  OAI211_X1 U21076 ( .C1(n18052), .C2(n18009), .A(n18031), .B(n18008), .ZN(
        n18019) );
  OAI221_X1 U21077 ( .B1(n18010), .B2(n18107), .C1(n18010), .C2(n18019), .A(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18015) );
  AOI22_X1 U21078 ( .A1(n18013), .A2(n9717), .B1(n18012), .B2(n18011), .ZN(
        n18014) );
  OAI221_X1 U21079 ( .B1(n9726), .B2(n18015), .C1(n18193), .C2(n18763), .A(
        n18014), .ZN(P3_U2846) );
  INV_X1 U21080 ( .A(n18058), .ZN(n18030) );
  OAI21_X1 U21081 ( .B1(n18017), .B2(n18030), .A(n18016), .ZN(n18018) );
  AOI22_X1 U21082 ( .A1(n18021), .A2(n18020), .B1(n18019), .B2(n18018), .ZN(
        n18028) );
  AOI22_X1 U21083 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18187), .B1(
        n9726), .B2(P3_REIP_REG_15__SCAN_IN), .ZN(n18027) );
  NOR2_X1 U21084 ( .A1(n18022), .A2(n18198), .ZN(n18024) );
  AOI22_X1 U21085 ( .A1(n18025), .A2(n9717), .B1(n18024), .B2(n18023), .ZN(
        n18026) );
  OAI211_X1 U21086 ( .C1(n18028), .C2(n18185), .A(n18027), .B(n18026), .ZN(
        P3_U2847) );
  INV_X1 U21087 ( .A(n18029), .ZN(n18033) );
  OAI21_X1 U21088 ( .B1(n18033), .B2(n18030), .A(n18034), .ZN(n18038) );
  AOI21_X1 U21089 ( .B1(n9930), .B2(n18093), .A(n18094), .ZN(n18048) );
  OAI211_X1 U21090 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n18186), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B(n18031), .ZN(n18032) );
  AOI211_X1 U21091 ( .C1(n18082), .C2(n18033), .A(n18048), .B(n18032), .ZN(
        n18035) );
  OAI22_X1 U21092 ( .A1(n18035), .A2(n18185), .B1(n18034), .B2(n18165), .ZN(
        n18037) );
  AOI21_X1 U21093 ( .B1(n18038), .B2(n18037), .A(n18036), .ZN(n18042) );
  AOI22_X1 U21094 ( .A1(n18184), .A2(n18040), .B1(n9717), .B2(n18039), .ZN(
        n18041) );
  OAI211_X1 U21095 ( .C1(n18044), .C2(n18043), .A(n18042), .B(n18041), .ZN(
        P3_U2848) );
  AOI22_X1 U21096 ( .A1(n9726), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n9717), .B2(
        n18045), .ZN(n18055) );
  AOI21_X1 U21097 ( .B1(n18046), .B2(n18092), .A(n18052), .ZN(n18078) );
  AOI211_X1 U21098 ( .C1(n18069), .C2(n18047), .A(n18068), .B(n18078), .ZN(
        n18050) );
  INV_X1 U21099 ( .A(n18048), .ZN(n18049) );
  OAI211_X1 U21100 ( .C1(n18051), .C2(n18072), .A(n18050), .B(n18049), .ZN(
        n18061) );
  OAI21_X1 U21101 ( .B1(n18052), .B2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18191), .ZN(n18053) );
  OAI211_X1 U21102 ( .C1(n18061), .C2(n18053), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18193), .ZN(n18054) );
  OAI211_X1 U21103 ( .C1(n18101), .C2(n18056), .A(n18055), .B(n18054), .ZN(
        P3_U2849) );
  AOI22_X1 U21104 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18187), .B1(
        n9726), .B2(P3_REIP_REG_12__SCAN_IN), .ZN(n18065) );
  NOR2_X1 U21105 ( .A1(n18058), .A2(n18057), .ZN(n18060) );
  NOR2_X1 U21106 ( .A1(n18060), .A2(n18059), .ZN(n18063) );
  OAI221_X1 U21107 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18063), 
        .C1(n18062), .C2(n18061), .A(n18191), .ZN(n18064) );
  OAI211_X1 U21108 ( .C1(n18066), .C2(n18090), .A(n18065), .B(n18064), .ZN(
        P3_U2850) );
  AOI22_X1 U21109 ( .A1(n9726), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n9717), .B2(
        n18067), .ZN(n18080) );
  AOI21_X1 U21110 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18093), .A(
        n18094), .ZN(n18074) );
  AOI211_X1 U21111 ( .C1(n18070), .C2(n18069), .A(n18068), .B(n18185), .ZN(
        n18071) );
  OAI21_X1 U21112 ( .B1(n18073), .B2(n18072), .A(n18071), .ZN(n18096) );
  AOI211_X1 U21113 ( .C1(n18076), .C2(n18075), .A(n18074), .B(n18096), .ZN(
        n18086) );
  OAI21_X1 U21114 ( .B1(n18094), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18086), .ZN(n18077) );
  OAI211_X1 U21115 ( .C1(n18078), .C2(n18077), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18193), .ZN(n18079) );
  OAI211_X1 U21116 ( .C1(n18081), .C2(n18101), .A(n18080), .B(n18079), .ZN(
        P3_U2851) );
  OAI21_X1 U21117 ( .B1(n18083), .B2(n18100), .A(n18082), .ZN(n18085) );
  AOI21_X1 U21118 ( .B1(n18086), .B2(n18085), .A(n18084), .ZN(n18088) );
  NOR3_X1 U21119 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18100), .A3(
        n18101), .ZN(n18087) );
  AOI221_X1 U21120 ( .B1(P3_REIP_REG_10__SCAN_IN), .B2(n9726), .C1(n18088), 
        .C2(n18193), .A(n18087), .ZN(n18089) );
  OAI21_X1 U21121 ( .B1(n18091), .B2(n18090), .A(n18089), .ZN(P3_U2852) );
  OAI21_X1 U21122 ( .B1(n18094), .B2(n18093), .A(n18092), .ZN(n18095) );
  OAI21_X1 U21123 ( .B1(n18096), .B2(n18095), .A(n18193), .ZN(n18099) );
  AOI22_X1 U21124 ( .A1(n9726), .A2(P3_REIP_REG_9__SCAN_IN), .B1(n9717), .B2(
        n18097), .ZN(n18098) );
  OAI221_X1 U21125 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n18101), .C1(
        n18100), .C2(n18099), .A(n18098), .ZN(P3_U2853) );
  NOR2_X1 U21126 ( .A1(n18157), .A2(n18185), .ZN(n18139) );
  AND2_X1 U21127 ( .A1(n18102), .A2(n18139), .ZN(n18110) );
  NOR3_X1 U21128 ( .A1(n18167), .A2(n18118), .A3(n18103), .ZN(n18105) );
  OAI21_X1 U21129 ( .B1(n18144), .B2(n18118), .A(n18145), .ZN(n18104) );
  OAI21_X1 U21130 ( .B1(n18147), .B2(n18105), .A(n18104), .ZN(n18127) );
  AOI211_X1 U21131 ( .C1(n18107), .C2(n18131), .A(n18106), .B(n18127), .ZN(
        n18126) );
  OAI21_X1 U21132 ( .B1(n18126), .B2(n18180), .A(n18165), .ZN(n18109) );
  AOI221_X1 U21133 ( .B1(n18110), .B2(n9900), .C1(n18109), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18108), .ZN(n18116) );
  AOI22_X1 U21134 ( .A1(n18114), .A2(n18113), .B1(n9717), .B2(n18111), .ZN(
        n18115) );
  OAI211_X1 U21135 ( .C1(n18198), .C2(n18117), .A(n18116), .B(n18115), .ZN(
        P3_U2854) );
  INV_X1 U21136 ( .A(n18139), .ZN(n18143) );
  NOR2_X1 U21137 ( .A1(n18118), .A2(n18143), .ZN(n18132) );
  AOI22_X1 U21138 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18191), .B1(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18132), .ZN(n18125) );
  AOI21_X1 U21139 ( .B1(n18187), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n18119), .ZN(n18124) );
  INV_X1 U21140 ( .A(n18120), .ZN(n18121) );
  AOI22_X1 U21141 ( .A1(n18184), .A2(n18122), .B1(n18136), .B2(n18121), .ZN(
        n18123) );
  OAI211_X1 U21142 ( .C1(n18126), .C2(n18125), .A(n18124), .B(n18123), .ZN(
        P3_U2855) );
  AOI21_X1 U21143 ( .B1(n18127), .B2(n18191), .A(n18187), .ZN(n18128) );
  INV_X1 U21144 ( .A(n18128), .ZN(n18138) );
  INV_X1 U21145 ( .A(n18136), .ZN(n18196) );
  OAI22_X1 U21146 ( .A1(n18193), .A2(n18747), .B1(n18196), .B2(n18129), .ZN(
        n18130) );
  AOI221_X1 U21147 ( .B1(n18132), .B2(n18131), .C1(n18138), .C2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A(n18130), .ZN(n18133) );
  OAI21_X1 U21148 ( .B1(n18198), .B2(n18134), .A(n18133), .ZN(P3_U2856) );
  AOI22_X1 U21149 ( .A1(n9726), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18136), .B2(
        n18135), .ZN(n18142) );
  AOI22_X1 U21150 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18138), .B1(
        n18184), .B2(n18137), .ZN(n18141) );
  NAND4_X1 U21151 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n18139), .A4(n20760), .ZN(
        n18140) );
  NAND3_X1 U21152 ( .A1(n18142), .A2(n18141), .A3(n18140), .ZN(P3_U2857) );
  INV_X1 U21153 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18164) );
  NOR2_X1 U21154 ( .A1(n18164), .A2(n18143), .ZN(n18153) );
  NAND2_X1 U21155 ( .A1(n18145), .A2(n18144), .ZN(n18173) );
  OAI211_X1 U21156 ( .C1(n18147), .C2(n18146), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n18173), .ZN(n18148) );
  NOR2_X1 U21157 ( .A1(n18167), .A2(n18148), .ZN(n18156) );
  OAI21_X1 U21158 ( .B1(n18156), .B2(n18180), .A(n18165), .ZN(n18151) );
  OAI22_X1 U21159 ( .A1(n18193), .A2(n18744), .B1(n18198), .B2(n18149), .ZN(
        n18150) );
  AOI221_X1 U21160 ( .B1(n18153), .B2(n18152), .C1(n18151), .C2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A(n18150), .ZN(n18154) );
  OAI21_X1 U21161 ( .B1(n18196), .B2(n18155), .A(n18154), .ZN(P3_U2858) );
  AOI211_X1 U21162 ( .C1(n18157), .C2(n18164), .A(n18156), .B(n18185), .ZN(
        n18161) );
  OAI22_X1 U21163 ( .A1(n18198), .A2(n18159), .B1(n18196), .B2(n18158), .ZN(
        n18160) );
  NOR2_X1 U21164 ( .A1(n18161), .A2(n18160), .ZN(n18163) );
  OAI211_X1 U21165 ( .C1(n18165), .C2(n18164), .A(n18163), .B(n18162), .ZN(
        P3_U2859) );
  NAND2_X1 U21166 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18169) );
  INV_X1 U21167 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18814) );
  OAI21_X1 U21168 ( .B1(n18167), .B2(n18814), .A(n18166), .ZN(n18168) );
  OAI21_X1 U21169 ( .B1(n18169), .B2(n18685), .A(n18168), .ZN(n18172) );
  NOR2_X1 U21170 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18814), .ZN(
        n18170) );
  AOI22_X1 U21171 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18172), .B1(
        n18171), .B2(n18170), .ZN(n18174) );
  OAI211_X1 U21172 ( .C1(n18679), .C2(n18175), .A(n18174), .B(n18173), .ZN(
        n18176) );
  AOI22_X1 U21173 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18187), .B1(
        n18191), .B2(n18176), .ZN(n18178) );
  OAI211_X1 U21174 ( .C1(n18198), .C2(n18179), .A(n18178), .B(n18177), .ZN(
        P3_U2860) );
  INV_X1 U21175 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18739) );
  NOR2_X1 U21176 ( .A1(n18193), .A2(n18739), .ZN(n18182) );
  AOI211_X1 U21177 ( .C1(n18656), .C2(n21021), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18180), .ZN(n18181) );
  AOI211_X1 U21178 ( .C1(n18184), .C2(n18183), .A(n18182), .B(n18181), .ZN(
        n18189) );
  NOR3_X1 U21179 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18186), .A3(
        n18185), .ZN(n18192) );
  OAI21_X1 U21180 ( .B1(n18187), .B2(n18192), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18188) );
  OAI211_X1 U21181 ( .C1(n18190), .C2(n18196), .A(n18189), .B(n18188), .ZN(
        P3_U2861) );
  AOI21_X1 U21182 ( .B1(n18656), .B2(n18191), .A(n21021), .ZN(n18194) );
  AOI221_X1 U21183 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(n9726), .C1(n18194), 
        .C2(n18193), .A(n18192), .ZN(n18195) );
  OAI221_X1 U21184 ( .B1(n18199), .B2(n18198), .C1(n18197), .C2(n18196), .A(
        n18195), .ZN(P3_U2862) );
  AOI211_X1 U21185 ( .C1(n18201), .C2(n18200), .A(n18865), .B(n18813), .ZN(
        n18703) );
  OAI21_X1 U21186 ( .B1(n18703), .B2(n18250), .A(n18206), .ZN(n18202) );
  OAI221_X1 U21187 ( .B1(n21027), .B2(n18848), .C1(n21027), .C2(n18206), .A(
        n18202), .ZN(P3_U2863) );
  INV_X1 U21188 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18249) );
  NOR2_X1 U21189 ( .A1(n18663), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18383) );
  INV_X1 U21190 ( .A(n18383), .ZN(n18385) );
  NOR2_X1 U21191 ( .A1(n18249), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18478) );
  NAND2_X1 U21192 ( .A1(n18209), .A2(n18478), .ZN(n18500) );
  AND2_X1 U21193 ( .A1(n18385), .A2(n18500), .ZN(n18204) );
  OAI22_X1 U21194 ( .A1(n18205), .A2(n18249), .B1(n18204), .B2(n18203), .ZN(
        P3_U2866) );
  NOR2_X1 U21195 ( .A1(n18207), .A2(n18206), .ZN(P3_U2867) );
  NAND2_X1 U21196 ( .A1(n18593), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18597) );
  NAND2_X1 U21197 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18208) );
  NAND2_X1 U21198 ( .A1(n21027), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18451) );
  NOR2_X2 U21199 ( .A1(n18208), .A2(n18451), .ZN(n18581) );
  INV_X1 U21200 ( .A(n18581), .ZN(n18265) );
  NOR2_X1 U21201 ( .A1(n18208), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18592) );
  NAND2_X1 U21202 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18592), .ZN(
        n18646) );
  INV_X1 U21203 ( .A(n18646), .ZN(n18630) );
  NAND2_X1 U21204 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18593), .ZN(n18557) );
  INV_X1 U21205 ( .A(n18557), .ZN(n18589) );
  INV_X1 U21206 ( .A(n18452), .ZN(n18503) );
  AND2_X1 U21207 ( .A1(n18503), .A2(BUF2_REG_0__SCAN_IN), .ZN(n18588) );
  NAND2_X1 U21208 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18658) );
  NOR2_X2 U21209 ( .A1(n18658), .A2(n18208), .ZN(n18641) );
  NAND2_X1 U21210 ( .A1(n18659), .A2(n21027), .ZN(n18660) );
  NOR2_X1 U21211 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18292) );
  INV_X1 U21212 ( .A(n18292), .ZN(n18293) );
  NOR2_X2 U21213 ( .A1(n18660), .A2(n18293), .ZN(n18312) );
  NOR2_X1 U21214 ( .A1(n18641), .A2(n18312), .ZN(n18270) );
  NOR2_X1 U21215 ( .A1(n18713), .A2(n18270), .ZN(n18243) );
  AOI22_X1 U21216 ( .A1(n18630), .A2(n18589), .B1(n18588), .B2(n18243), .ZN(
        n18215) );
  AOI21_X1 U21217 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n18270), .ZN(n18210) );
  NAND2_X1 U21218 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18659), .ZN(
        n18430) );
  AND2_X1 U21219 ( .A1(n18451), .A2(n18430), .ZN(n18501) );
  OR2_X1 U21220 ( .A1(n18208), .A2(n18501), .ZN(n18550) );
  NOR2_X1 U21221 ( .A1(n18452), .A2(n18550), .ZN(n18554) );
  AOI22_X1 U21222 ( .A1(n18503), .A2(n18210), .B1(n18209), .B2(n18554), .ZN(
        n18246) );
  NAND2_X1 U21223 ( .A1(n18212), .A2(n18211), .ZN(n18244) );
  NOR2_X2 U21224 ( .A1(n18213), .A2(n18244), .ZN(n18594) );
  AOI22_X1 U21225 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18246), .B1(
        n18312), .B2(n18594), .ZN(n18214) );
  OAI211_X1 U21226 ( .C1(n18597), .C2(n18265), .A(n18215), .B(n18214), .ZN(
        P3_U2868) );
  NOR2_X1 U21227 ( .A1(n18216), .A2(n18454), .ZN(n18530) );
  AND2_X1 U21228 ( .A1(n18593), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18599) );
  NOR2_X2 U21229 ( .A1(n18452), .A2(n20954), .ZN(n18598) );
  AOI22_X1 U21230 ( .A1(n18581), .A2(n18599), .B1(n18243), .B2(n18598), .ZN(
        n18219) );
  NOR2_X2 U21231 ( .A1(n18217), .A2(n18244), .ZN(n18600) );
  AOI22_X1 U21232 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18246), .B1(
        n18312), .B2(n18600), .ZN(n18218) );
  OAI211_X1 U21233 ( .C1(n18646), .C2(n18603), .A(n18219), .B(n18218), .ZN(
        P3_U2869) );
  INV_X1 U21234 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n18220) );
  NOR2_X1 U21235 ( .A1(n18220), .A2(n18454), .ZN(n18560) );
  INV_X1 U21236 ( .A(n18560), .ZN(n18609) );
  NAND2_X1 U21237 ( .A1(n18593), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18563) );
  INV_X1 U21238 ( .A(n18563), .ZN(n18605) );
  NOR2_X2 U21239 ( .A1(n18452), .A2(n20804), .ZN(n18604) );
  AOI22_X1 U21240 ( .A1(n18581), .A2(n18605), .B1(n18243), .B2(n18604), .ZN(
        n18223) );
  NOR2_X2 U21241 ( .A1(n18221), .A2(n18244), .ZN(n18606) );
  AOI22_X1 U21242 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18246), .B1(
        n18312), .B2(n18606), .ZN(n18222) );
  OAI211_X1 U21243 ( .C1(n18646), .C2(n18609), .A(n18223), .B(n18222), .ZN(
        P3_U2870) );
  NOR2_X1 U21244 ( .A1(n20810), .A2(n18454), .ZN(n18611) );
  INV_X1 U21245 ( .A(n18611), .ZN(n18567) );
  NAND2_X1 U21246 ( .A1(n18593), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18615) );
  INV_X1 U21247 ( .A(n18615), .ZN(n18564) );
  NOR2_X2 U21248 ( .A1(n18452), .A2(n18224), .ZN(n18610) );
  AOI22_X1 U21249 ( .A1(n18581), .A2(n18564), .B1(n18243), .B2(n18610), .ZN(
        n18227) );
  NOR2_X2 U21250 ( .A1(n18225), .A2(n18244), .ZN(n18612) );
  AOI22_X1 U21251 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18246), .B1(
        n18312), .B2(n18612), .ZN(n18226) );
  OAI211_X1 U21252 ( .C1(n18646), .C2(n18567), .A(n18227), .B(n18226), .ZN(
        P3_U2871) );
  INV_X1 U21253 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n19232) );
  NOR2_X1 U21254 ( .A1(n19232), .A2(n18454), .ZN(n18617) );
  INV_X1 U21255 ( .A(n18617), .ZN(n18516) );
  NAND2_X1 U21256 ( .A1(n18593), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18621) );
  INV_X1 U21257 ( .A(n18621), .ZN(n18512) );
  NOR2_X2 U21258 ( .A1(n18452), .A2(n18228), .ZN(n18616) );
  AOI22_X1 U21259 ( .A1(n18581), .A2(n18512), .B1(n18243), .B2(n18616), .ZN(
        n18231) );
  NOR2_X2 U21260 ( .A1(n18229), .A2(n18244), .ZN(n18618) );
  AOI22_X1 U21261 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18246), .B1(
        n18312), .B2(n18618), .ZN(n18230) );
  OAI211_X1 U21262 ( .C1(n18646), .C2(n18516), .A(n18231), .B(n18230), .ZN(
        P3_U2872) );
  NOR2_X1 U21263 ( .A1(n18232), .A2(n18454), .ZN(n18623) );
  INV_X1 U21264 ( .A(n18623), .ZN(n18573) );
  NAND2_X1 U21265 ( .A1(n18593), .A2(BUF2_REG_21__SCAN_IN), .ZN(n18627) );
  INV_X1 U21266 ( .A(n18627), .ZN(n18570) );
  NOR2_X2 U21267 ( .A1(n18452), .A2(n18233), .ZN(n18622) );
  AOI22_X1 U21268 ( .A1(n18581), .A2(n18570), .B1(n18243), .B2(n18622), .ZN(
        n18236) );
  NOR2_X2 U21269 ( .A1(n18234), .A2(n18244), .ZN(n18624) );
  AOI22_X1 U21270 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18246), .B1(
        n18312), .B2(n18624), .ZN(n18235) );
  OAI211_X1 U21271 ( .C1(n18646), .C2(n18573), .A(n18236), .B(n18235), .ZN(
        P3_U2873) );
  NOR2_X1 U21272 ( .A1(n15003), .A2(n18454), .ZN(n18629) );
  INV_X1 U21273 ( .A(n18629), .ZN(n18578) );
  NAND2_X1 U21274 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18593), .ZN(n18635) );
  INV_X1 U21275 ( .A(n18635), .ZN(n18575) );
  NOR2_X2 U21276 ( .A1(n18237), .A2(n18452), .ZN(n18628) );
  AOI22_X1 U21277 ( .A1(n18630), .A2(n18575), .B1(n18243), .B2(n18628), .ZN(
        n18240) );
  NOR2_X2 U21278 ( .A1(n18238), .A2(n18244), .ZN(n18631) );
  AOI22_X1 U21279 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18246), .B1(
        n18312), .B2(n18631), .ZN(n18239) );
  OAI211_X1 U21280 ( .C1(n18265), .C2(n18578), .A(n18240), .B(n18239), .ZN(
        P3_U2874) );
  NOR2_X1 U21281 ( .A1(n18454), .A2(n18241), .ZN(n18639) );
  INV_X1 U21282 ( .A(n18639), .ZN(n18586) );
  NAND2_X1 U21283 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18593), .ZN(n18645) );
  INV_X1 U21284 ( .A(n18645), .ZN(n18580) );
  NOR2_X2 U21285 ( .A1(n18242), .A2(n18452), .ZN(n18637) );
  AOI22_X1 U21286 ( .A1(n18581), .A2(n18580), .B1(n18243), .B2(n18637), .ZN(
        n18248) );
  NOR2_X2 U21287 ( .A1(n18245), .A2(n18244), .ZN(n18640) );
  AOI22_X1 U21288 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18246), .B1(
        n18312), .B2(n18640), .ZN(n18247) );
  OAI211_X1 U21289 ( .C1(n18646), .C2(n18586), .A(n18248), .B(n18247), .ZN(
        P3_U2875) );
  INV_X1 U21290 ( .A(n18641), .ZN(n18290) );
  AOI22_X1 U21291 ( .A1(n18581), .A2(n18589), .B1(n18588), .B2(n18266), .ZN(
        n18252) );
  NOR2_X1 U21292 ( .A1(n18249), .A2(n18427), .ZN(n18590) );
  NOR2_X1 U21293 ( .A1(n18452), .A2(n18250), .ZN(n18591) );
  AND2_X1 U21294 ( .A1(n18659), .A2(n18591), .ZN(n18337) );
  AOI22_X1 U21295 ( .A1(n18593), .A2(n18590), .B1(n18292), .B2(n18337), .ZN(
        n18267) );
  NOR2_X2 U21296 ( .A1(n18430), .A2(n18293), .ZN(n18333) );
  AOI22_X1 U21297 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18267), .B1(
        n18594), .B2(n18333), .ZN(n18251) );
  OAI211_X1 U21298 ( .C1(n18597), .C2(n18290), .A(n18252), .B(n18251), .ZN(
        P3_U2876) );
  AOI22_X1 U21299 ( .A1(n18641), .A2(n18599), .B1(n18598), .B2(n18266), .ZN(
        n18254) );
  AOI22_X1 U21300 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18267), .B1(
        n18600), .B2(n18333), .ZN(n18253) );
  OAI211_X1 U21301 ( .C1(n18265), .C2(n18603), .A(n18254), .B(n18253), .ZN(
        P3_U2877) );
  AOI22_X1 U21302 ( .A1(n18581), .A2(n18560), .B1(n18604), .B2(n18266), .ZN(
        n18256) );
  AOI22_X1 U21303 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18267), .B1(
        n18606), .B2(n18333), .ZN(n18255) );
  OAI211_X1 U21304 ( .C1(n18290), .C2(n18563), .A(n18256), .B(n18255), .ZN(
        P3_U2878) );
  AOI22_X1 U21305 ( .A1(n18581), .A2(n18611), .B1(n18610), .B2(n18266), .ZN(
        n18258) );
  AOI22_X1 U21306 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18267), .B1(
        n18612), .B2(n18333), .ZN(n18257) );
  OAI211_X1 U21307 ( .C1(n18290), .C2(n18615), .A(n18258), .B(n18257), .ZN(
        P3_U2879) );
  AOI22_X1 U21308 ( .A1(n18581), .A2(n18617), .B1(n18616), .B2(n18266), .ZN(
        n18260) );
  AOI22_X1 U21309 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18267), .B1(
        n18618), .B2(n18333), .ZN(n18259) );
  OAI211_X1 U21310 ( .C1(n18290), .C2(n18621), .A(n18260), .B(n18259), .ZN(
        P3_U2880) );
  AOI22_X1 U21311 ( .A1(n18641), .A2(n18570), .B1(n18622), .B2(n18266), .ZN(
        n18262) );
  AOI22_X1 U21312 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18267), .B1(
        n18624), .B2(n18333), .ZN(n18261) );
  OAI211_X1 U21313 ( .C1(n18265), .C2(n18573), .A(n18262), .B(n18261), .ZN(
        P3_U2881) );
  AOI22_X1 U21314 ( .A1(n18641), .A2(n18629), .B1(n18628), .B2(n18266), .ZN(
        n18264) );
  AOI22_X1 U21315 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18267), .B1(
        n18631), .B2(n18333), .ZN(n18263) );
  OAI211_X1 U21316 ( .C1(n18265), .C2(n18635), .A(n18264), .B(n18263), .ZN(
        P3_U2882) );
  AOI22_X1 U21317 ( .A1(n18581), .A2(n18639), .B1(n18637), .B2(n18266), .ZN(
        n18269) );
  AOI22_X1 U21318 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18267), .B1(
        n18640), .B2(n18333), .ZN(n18268) );
  OAI211_X1 U21319 ( .C1(n18290), .C2(n18645), .A(n18269), .B(n18268), .ZN(
        P3_U2883) );
  INV_X1 U21320 ( .A(n18312), .ZN(n18309) );
  NOR2_X2 U21321 ( .A1(n18451), .A2(n18293), .ZN(n18355) );
  NOR2_X1 U21322 ( .A1(n18333), .A2(n18355), .ZN(n18315) );
  NOR2_X1 U21323 ( .A1(n18713), .A2(n18315), .ZN(n18286) );
  AOI22_X1 U21324 ( .A1(n18641), .A2(n18589), .B1(n18588), .B2(n18286), .ZN(
        n18273) );
  OAI22_X1 U21325 ( .A1(n18270), .A2(n18454), .B1(n18315), .B2(n18452), .ZN(
        n18271) );
  OAI21_X1 U21326 ( .B1(n18355), .B2(n18808), .A(n18271), .ZN(n18287) );
  AOI22_X1 U21327 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18287), .B1(
        n18594), .B2(n18355), .ZN(n18272) );
  OAI211_X1 U21328 ( .C1(n18597), .C2(n18309), .A(n18273), .B(n18272), .ZN(
        P3_U2884) );
  AOI22_X1 U21329 ( .A1(n18312), .A2(n18599), .B1(n18598), .B2(n18286), .ZN(
        n18275) );
  AOI22_X1 U21330 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18287), .B1(
        n18600), .B2(n18355), .ZN(n18274) );
  OAI211_X1 U21331 ( .C1(n18290), .C2(n18603), .A(n18275), .B(n18274), .ZN(
        P3_U2885) );
  AOI22_X1 U21332 ( .A1(n18641), .A2(n18560), .B1(n18604), .B2(n18286), .ZN(
        n18277) );
  AOI22_X1 U21333 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18287), .B1(
        n18606), .B2(n18355), .ZN(n18276) );
  OAI211_X1 U21334 ( .C1(n18309), .C2(n18563), .A(n18277), .B(n18276), .ZN(
        P3_U2886) );
  AOI22_X1 U21335 ( .A1(n18312), .A2(n18564), .B1(n18610), .B2(n18286), .ZN(
        n18279) );
  AOI22_X1 U21336 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18287), .B1(
        n18612), .B2(n18355), .ZN(n18278) );
  OAI211_X1 U21337 ( .C1(n18290), .C2(n18567), .A(n18279), .B(n18278), .ZN(
        P3_U2887) );
  AOI22_X1 U21338 ( .A1(n18641), .A2(n18617), .B1(n18616), .B2(n18286), .ZN(
        n18281) );
  AOI22_X1 U21339 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18287), .B1(
        n18618), .B2(n18355), .ZN(n18280) );
  OAI211_X1 U21340 ( .C1(n18309), .C2(n18621), .A(n18281), .B(n18280), .ZN(
        P3_U2888) );
  AOI22_X1 U21341 ( .A1(n18312), .A2(n18570), .B1(n18622), .B2(n18286), .ZN(
        n18283) );
  AOI22_X1 U21342 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18287), .B1(
        n18624), .B2(n18355), .ZN(n18282) );
  OAI211_X1 U21343 ( .C1(n18290), .C2(n18573), .A(n18283), .B(n18282), .ZN(
        P3_U2889) );
  AOI22_X1 U21344 ( .A1(n18312), .A2(n18629), .B1(n18628), .B2(n18286), .ZN(
        n18285) );
  AOI22_X1 U21345 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18287), .B1(
        n18631), .B2(n18355), .ZN(n18284) );
  OAI211_X1 U21346 ( .C1(n18290), .C2(n18635), .A(n18285), .B(n18284), .ZN(
        P3_U2890) );
  AOI22_X1 U21347 ( .A1(n18312), .A2(n18580), .B1(n18637), .B2(n18286), .ZN(
        n18289) );
  AOI22_X1 U21348 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18287), .B1(
        n18640), .B2(n18355), .ZN(n18288) );
  OAI211_X1 U21349 ( .C1(n18290), .C2(n18586), .A(n18289), .B(n18288), .ZN(
        P3_U2891) );
  INV_X1 U21350 ( .A(n18333), .ZN(n18329) );
  AOI22_X1 U21351 ( .A1(n18659), .A2(n18359), .B1(n18658), .B2(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18291) );
  AND2_X1 U21352 ( .A1(n18503), .A2(n18291), .ZN(n18384) );
  NAND2_X1 U21353 ( .A1(n18292), .A2(n18384), .ZN(n18311) );
  NOR2_X1 U21354 ( .A1(n18659), .A2(n18293), .ZN(n18338) );
  INV_X1 U21355 ( .A(n18338), .ZN(n18294) );
  NOR2_X1 U21356 ( .A1(n18713), .A2(n18294), .ZN(n18310) );
  AOI22_X1 U21357 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18311), .B1(
        n18588), .B2(n18310), .ZN(n18296) );
  NAND2_X1 U21358 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18338), .ZN(
        n18382) );
  INV_X1 U21359 ( .A(n18382), .ZN(n18374) );
  AOI22_X1 U21360 ( .A1(n18312), .A2(n18589), .B1(n18594), .B2(n18374), .ZN(
        n18295) );
  OAI211_X1 U21361 ( .C1(n18597), .C2(n18329), .A(n18296), .B(n18295), .ZN(
        P3_U2892) );
  AOI22_X1 U21362 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18311), .B1(
        n18598), .B2(n18310), .ZN(n18298) );
  AOI22_X1 U21363 ( .A1(n18600), .A2(n18374), .B1(n18599), .B2(n18333), .ZN(
        n18297) );
  OAI211_X1 U21364 ( .C1(n18309), .C2(n18603), .A(n18298), .B(n18297), .ZN(
        P3_U2893) );
  AOI22_X1 U21365 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18311), .B1(
        n18604), .B2(n18310), .ZN(n18300) );
  AOI22_X1 U21366 ( .A1(n18312), .A2(n18560), .B1(n18606), .B2(n18374), .ZN(
        n18299) );
  OAI211_X1 U21367 ( .C1(n18563), .C2(n18329), .A(n18300), .B(n18299), .ZN(
        P3_U2894) );
  AOI22_X1 U21368 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18311), .B1(
        n18610), .B2(n18310), .ZN(n18302) );
  AOI22_X1 U21369 ( .A1(n18312), .A2(n18611), .B1(n18612), .B2(n18374), .ZN(
        n18301) );
  OAI211_X1 U21370 ( .C1(n18615), .C2(n18329), .A(n18302), .B(n18301), .ZN(
        P3_U2895) );
  AOI22_X1 U21371 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18311), .B1(
        n18616), .B2(n18310), .ZN(n18304) );
  AOI22_X1 U21372 ( .A1(n18618), .A2(n18374), .B1(n18512), .B2(n18333), .ZN(
        n18303) );
  OAI211_X1 U21373 ( .C1(n18309), .C2(n18516), .A(n18304), .B(n18303), .ZN(
        P3_U2896) );
  AOI22_X1 U21374 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18311), .B1(
        n18622), .B2(n18310), .ZN(n18306) );
  AOI22_X1 U21375 ( .A1(n18624), .A2(n18374), .B1(n18570), .B2(n18333), .ZN(
        n18305) );
  OAI211_X1 U21376 ( .C1(n18309), .C2(n18573), .A(n18306), .B(n18305), .ZN(
        P3_U2897) );
  AOI22_X1 U21377 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18311), .B1(
        n18628), .B2(n18310), .ZN(n18308) );
  AOI22_X1 U21378 ( .A1(n18629), .A2(n18333), .B1(n18631), .B2(n18374), .ZN(
        n18307) );
  OAI211_X1 U21379 ( .C1(n18309), .C2(n18635), .A(n18308), .B(n18307), .ZN(
        P3_U2898) );
  AOI22_X1 U21380 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18311), .B1(
        n18637), .B2(n18310), .ZN(n18314) );
  AOI22_X1 U21381 ( .A1(n18312), .A2(n18639), .B1(n18640), .B2(n18374), .ZN(
        n18313) );
  OAI211_X1 U21382 ( .C1(n18645), .C2(n18329), .A(n18314), .B(n18313), .ZN(
        P3_U2899) );
  INV_X1 U21383 ( .A(n18597), .ZN(n18551) );
  NOR2_X2 U21384 ( .A1(n18660), .A2(n18385), .ZN(n18378) );
  NOR2_X1 U21385 ( .A1(n18374), .A2(n18378), .ZN(n18360) );
  NOR2_X1 U21386 ( .A1(n18713), .A2(n18360), .ZN(n18332) );
  AOI22_X1 U21387 ( .A1(n18551), .A2(n18355), .B1(n18588), .B2(n18332), .ZN(
        n18318) );
  OAI21_X1 U21388 ( .B1(n18315), .B2(n18359), .A(n18360), .ZN(n18316) );
  OAI211_X1 U21389 ( .C1(n18378), .C2(n18808), .A(n18503), .B(n18316), .ZN(
        n18334) );
  AOI22_X1 U21390 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18334), .B1(
        n18594), .B2(n18378), .ZN(n18317) );
  OAI211_X1 U21391 ( .C1(n18557), .C2(n18329), .A(n18318), .B(n18317), .ZN(
        P3_U2900) );
  AOI22_X1 U21392 ( .A1(n18599), .A2(n18355), .B1(n18598), .B2(n18332), .ZN(
        n18320) );
  AOI22_X1 U21393 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18334), .B1(
        n18600), .B2(n18378), .ZN(n18319) );
  OAI211_X1 U21394 ( .C1(n18603), .C2(n18329), .A(n18320), .B(n18319), .ZN(
        P3_U2901) );
  AOI22_X1 U21395 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18334), .B1(
        n18604), .B2(n18332), .ZN(n18322) );
  AOI22_X1 U21396 ( .A1(n18606), .A2(n18378), .B1(n18605), .B2(n18355), .ZN(
        n18321) );
  OAI211_X1 U21397 ( .C1(n18609), .C2(n18329), .A(n18322), .B(n18321), .ZN(
        P3_U2902) );
  AOI22_X1 U21398 ( .A1(n18610), .A2(n18332), .B1(n18564), .B2(n18355), .ZN(
        n18324) );
  AOI22_X1 U21399 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18334), .B1(
        n18612), .B2(n18378), .ZN(n18323) );
  OAI211_X1 U21400 ( .C1(n18567), .C2(n18329), .A(n18324), .B(n18323), .ZN(
        P3_U2903) );
  INV_X1 U21401 ( .A(n18355), .ZN(n18347) );
  AOI22_X1 U21402 ( .A1(n18617), .A2(n18333), .B1(n18616), .B2(n18332), .ZN(
        n18326) );
  AOI22_X1 U21403 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18334), .B1(
        n18618), .B2(n18378), .ZN(n18325) );
  OAI211_X1 U21404 ( .C1(n18621), .C2(n18347), .A(n18326), .B(n18325), .ZN(
        P3_U2904) );
  AOI22_X1 U21405 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18334), .B1(
        n18622), .B2(n18332), .ZN(n18328) );
  AOI22_X1 U21406 ( .A1(n18624), .A2(n18378), .B1(n18570), .B2(n18355), .ZN(
        n18327) );
  OAI211_X1 U21407 ( .C1(n18573), .C2(n18329), .A(n18328), .B(n18327), .ZN(
        P3_U2905) );
  AOI22_X1 U21408 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18334), .B1(
        n18628), .B2(n18332), .ZN(n18331) );
  AOI22_X1 U21409 ( .A1(n18631), .A2(n18378), .B1(n18575), .B2(n18333), .ZN(
        n18330) );
  OAI211_X1 U21410 ( .C1(n18578), .C2(n18347), .A(n18331), .B(n18330), .ZN(
        P3_U2906) );
  AOI22_X1 U21411 ( .A1(n18639), .A2(n18333), .B1(n18637), .B2(n18332), .ZN(
        n18336) );
  AOI22_X1 U21412 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18334), .B1(
        n18640), .B2(n18378), .ZN(n18335) );
  OAI211_X1 U21413 ( .C1(n18645), .C2(n18347), .A(n18336), .B(n18335), .ZN(
        P3_U2907) );
  AOI22_X1 U21414 ( .A1(n18551), .A2(n18374), .B1(n18588), .B2(n18354), .ZN(
        n18340) );
  AOI22_X1 U21415 ( .A1(n18593), .A2(n18338), .B1(n18337), .B2(n18383), .ZN(
        n18356) );
  NOR2_X2 U21416 ( .A1(n18430), .A2(n18385), .ZN(n18423) );
  AOI22_X1 U21417 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18356), .B1(
        n18594), .B2(n18423), .ZN(n18339) );
  OAI211_X1 U21418 ( .C1(n18557), .C2(n18347), .A(n18340), .B(n18339), .ZN(
        P3_U2908) );
  AOI22_X1 U21419 ( .A1(n18599), .A2(n18374), .B1(n18598), .B2(n18354), .ZN(
        n18342) );
  AOI22_X1 U21420 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18356), .B1(
        n18600), .B2(n18423), .ZN(n18341) );
  OAI211_X1 U21421 ( .C1(n18603), .C2(n18347), .A(n18342), .B(n18341), .ZN(
        P3_U2909) );
  AOI22_X1 U21422 ( .A1(n18605), .A2(n18374), .B1(n18604), .B2(n18354), .ZN(
        n18344) );
  AOI22_X1 U21423 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18356), .B1(
        n18606), .B2(n18423), .ZN(n18343) );
  OAI211_X1 U21424 ( .C1(n18609), .C2(n18347), .A(n18344), .B(n18343), .ZN(
        P3_U2910) );
  AOI22_X1 U21425 ( .A1(n18610), .A2(n18354), .B1(n18564), .B2(n18374), .ZN(
        n18346) );
  AOI22_X1 U21426 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18356), .B1(
        n18612), .B2(n18423), .ZN(n18345) );
  OAI211_X1 U21427 ( .C1(n18567), .C2(n18347), .A(n18346), .B(n18345), .ZN(
        P3_U2911) );
  AOI22_X1 U21428 ( .A1(n18617), .A2(n18355), .B1(n18616), .B2(n18354), .ZN(
        n18349) );
  AOI22_X1 U21429 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18356), .B1(
        n18618), .B2(n18423), .ZN(n18348) );
  OAI211_X1 U21430 ( .C1(n18621), .C2(n18382), .A(n18349), .B(n18348), .ZN(
        P3_U2912) );
  AOI22_X1 U21431 ( .A1(n18623), .A2(n18355), .B1(n18622), .B2(n18354), .ZN(
        n18351) );
  AOI22_X1 U21432 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18356), .B1(
        n18624), .B2(n18423), .ZN(n18350) );
  OAI211_X1 U21433 ( .C1(n18627), .C2(n18382), .A(n18351), .B(n18350), .ZN(
        P3_U2913) );
  AOI22_X1 U21434 ( .A1(n18628), .A2(n18354), .B1(n18575), .B2(n18355), .ZN(
        n18353) );
  AOI22_X1 U21435 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18356), .B1(
        n18631), .B2(n18423), .ZN(n18352) );
  OAI211_X1 U21436 ( .C1(n18578), .C2(n18382), .A(n18353), .B(n18352), .ZN(
        P3_U2914) );
  AOI22_X1 U21437 ( .A1(n18639), .A2(n18355), .B1(n18637), .B2(n18354), .ZN(
        n18358) );
  AOI22_X1 U21438 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18356), .B1(
        n18640), .B2(n18423), .ZN(n18357) );
  OAI211_X1 U21439 ( .C1(n18645), .C2(n18382), .A(n18358), .B(n18357), .ZN(
        P3_U2915) );
  INV_X1 U21440 ( .A(n18378), .ZN(n18404) );
  NOR2_X1 U21441 ( .A1(n18423), .A2(n18437), .ZN(n18405) );
  NOR2_X1 U21442 ( .A1(n18713), .A2(n18405), .ZN(n18377) );
  AOI22_X1 U21443 ( .A1(n18589), .A2(n18374), .B1(n18588), .B2(n18377), .ZN(
        n18363) );
  OAI21_X1 U21444 ( .B1(n18360), .B2(n18359), .A(n18405), .ZN(n18361) );
  OAI211_X1 U21445 ( .C1(n18437), .C2(n18808), .A(n18503), .B(n18361), .ZN(
        n18379) );
  AOI22_X1 U21446 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18379), .B1(
        n18594), .B2(n18437), .ZN(n18362) );
  OAI211_X1 U21447 ( .C1(n18597), .C2(n18404), .A(n18363), .B(n18362), .ZN(
        P3_U2916) );
  AOI22_X1 U21448 ( .A1(n18599), .A2(n18378), .B1(n18598), .B2(n18377), .ZN(
        n18365) );
  AOI22_X1 U21449 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18379), .B1(
        n18600), .B2(n18437), .ZN(n18364) );
  OAI211_X1 U21450 ( .C1(n18603), .C2(n18382), .A(n18365), .B(n18364), .ZN(
        P3_U2917) );
  AOI22_X1 U21451 ( .A1(n18605), .A2(n18378), .B1(n18604), .B2(n18377), .ZN(
        n18367) );
  AOI22_X1 U21452 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18379), .B1(
        n18606), .B2(n18437), .ZN(n18366) );
  OAI211_X1 U21453 ( .C1(n18609), .C2(n18382), .A(n18367), .B(n18366), .ZN(
        P3_U2918) );
  AOI22_X1 U21454 ( .A1(n18611), .A2(n18374), .B1(n18610), .B2(n18377), .ZN(
        n18369) );
  AOI22_X1 U21455 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18379), .B1(
        n18612), .B2(n18437), .ZN(n18368) );
  OAI211_X1 U21456 ( .C1(n18615), .C2(n18404), .A(n18369), .B(n18368), .ZN(
        P3_U2919) );
  AOI22_X1 U21457 ( .A1(n18512), .A2(n18378), .B1(n18616), .B2(n18377), .ZN(
        n18371) );
  AOI22_X1 U21458 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18379), .B1(
        n18618), .B2(n18437), .ZN(n18370) );
  OAI211_X1 U21459 ( .C1(n18516), .C2(n18382), .A(n18371), .B(n18370), .ZN(
        P3_U2920) );
  AOI22_X1 U21460 ( .A1(n18623), .A2(n18374), .B1(n18622), .B2(n18377), .ZN(
        n18373) );
  AOI22_X1 U21461 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18379), .B1(
        n18624), .B2(n18437), .ZN(n18372) );
  OAI211_X1 U21462 ( .C1(n18627), .C2(n18404), .A(n18373), .B(n18372), .ZN(
        P3_U2921) );
  AOI22_X1 U21463 ( .A1(n18628), .A2(n18377), .B1(n18575), .B2(n18374), .ZN(
        n18376) );
  AOI22_X1 U21464 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18379), .B1(
        n18631), .B2(n18437), .ZN(n18375) );
  OAI211_X1 U21465 ( .C1(n18578), .C2(n18404), .A(n18376), .B(n18375), .ZN(
        P3_U2922) );
  AOI22_X1 U21466 ( .A1(n18580), .A2(n18378), .B1(n18637), .B2(n18377), .ZN(
        n18381) );
  AOI22_X1 U21467 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18379), .B1(
        n18640), .B2(n18437), .ZN(n18380) );
  OAI211_X1 U21468 ( .C1(n18586), .C2(n18382), .A(n18381), .B(n18380), .ZN(
        P3_U2923) );
  NAND2_X1 U21469 ( .A1(n18384), .A2(n18383), .ZN(n18401) );
  AOI22_X1 U21470 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18401), .B1(
        n18588), .B2(n18400), .ZN(n18387) );
  NOR2_X2 U21471 ( .A1(n18658), .A2(n18385), .ZN(n18473) );
  AOI22_X1 U21472 ( .A1(n18551), .A2(n18423), .B1(n18594), .B2(n18473), .ZN(
        n18386) );
  OAI211_X1 U21473 ( .C1(n18557), .C2(n18404), .A(n18387), .B(n18386), .ZN(
        P3_U2924) );
  AOI22_X1 U21474 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18401), .B1(
        n18598), .B2(n18400), .ZN(n18389) );
  AOI22_X1 U21475 ( .A1(n18600), .A2(n18473), .B1(n18599), .B2(n18423), .ZN(
        n18388) );
  OAI211_X1 U21476 ( .C1(n18603), .C2(n18404), .A(n18389), .B(n18388), .ZN(
        P3_U2925) );
  AOI22_X1 U21477 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18401), .B1(
        n18604), .B2(n18400), .ZN(n18391) );
  AOI22_X1 U21478 ( .A1(n18606), .A2(n18473), .B1(n18605), .B2(n18423), .ZN(
        n18390) );
  OAI211_X1 U21479 ( .C1(n18609), .C2(n18404), .A(n18391), .B(n18390), .ZN(
        P3_U2926) );
  AOI22_X1 U21480 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18401), .B1(
        n18610), .B2(n18400), .ZN(n18393) );
  AOI22_X1 U21481 ( .A1(n18612), .A2(n18473), .B1(n18564), .B2(n18423), .ZN(
        n18392) );
  OAI211_X1 U21482 ( .C1(n18567), .C2(n18404), .A(n18393), .B(n18392), .ZN(
        P3_U2927) );
  AOI22_X1 U21483 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18401), .B1(
        n18616), .B2(n18400), .ZN(n18395) );
  AOI22_X1 U21484 ( .A1(n18618), .A2(n18473), .B1(n18512), .B2(n18423), .ZN(
        n18394) );
  OAI211_X1 U21485 ( .C1(n18516), .C2(n18404), .A(n18395), .B(n18394), .ZN(
        P3_U2928) );
  AOI22_X1 U21486 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18401), .B1(
        n18622), .B2(n18400), .ZN(n18397) );
  AOI22_X1 U21487 ( .A1(n18624), .A2(n18473), .B1(n18570), .B2(n18423), .ZN(
        n18396) );
  OAI211_X1 U21488 ( .C1(n18573), .C2(n18404), .A(n18397), .B(n18396), .ZN(
        P3_U2929) );
  AOI22_X1 U21489 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18401), .B1(
        n18628), .B2(n18400), .ZN(n18399) );
  AOI22_X1 U21490 ( .A1(n18629), .A2(n18423), .B1(n18631), .B2(n18473), .ZN(
        n18398) );
  OAI211_X1 U21491 ( .C1(n18635), .C2(n18404), .A(n18399), .B(n18398), .ZN(
        P3_U2930) );
  AOI22_X1 U21492 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18401), .B1(
        n18637), .B2(n18400), .ZN(n18403) );
  AOI22_X1 U21493 ( .A1(n18640), .A2(n18473), .B1(n18580), .B2(n18423), .ZN(
        n18402) );
  OAI211_X1 U21494 ( .C1(n18586), .C2(n18404), .A(n18403), .B(n18402), .ZN(
        P3_U2931) );
  INV_X1 U21495 ( .A(n18423), .ZN(n18421) );
  INV_X1 U21496 ( .A(n18478), .ZN(n18479) );
  NOR2_X2 U21497 ( .A1(n18660), .A2(n18479), .ZN(n18496) );
  NOR2_X1 U21498 ( .A1(n18473), .A2(n18496), .ZN(n18455) );
  NOR2_X1 U21499 ( .A1(n18713), .A2(n18455), .ZN(n18422) );
  AOI22_X1 U21500 ( .A1(n18551), .A2(n18437), .B1(n18588), .B2(n18422), .ZN(
        n18408) );
  OAI22_X1 U21501 ( .A1(n18405), .A2(n18454), .B1(n18455), .B2(n18452), .ZN(
        n18406) );
  OAI21_X1 U21502 ( .B1(n18496), .B2(n18808), .A(n18406), .ZN(n18424) );
  AOI22_X1 U21503 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18424), .B1(
        n18594), .B2(n18496), .ZN(n18407) );
  OAI211_X1 U21504 ( .C1(n18557), .C2(n18421), .A(n18408), .B(n18407), .ZN(
        P3_U2932) );
  AOI22_X1 U21505 ( .A1(n18599), .A2(n18437), .B1(n18598), .B2(n18422), .ZN(
        n18410) );
  AOI22_X1 U21506 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18424), .B1(
        n18600), .B2(n18496), .ZN(n18409) );
  OAI211_X1 U21507 ( .C1(n18603), .C2(n18421), .A(n18410), .B(n18409), .ZN(
        P3_U2933) );
  AOI22_X1 U21508 ( .A1(n18605), .A2(n18437), .B1(n18604), .B2(n18422), .ZN(
        n18412) );
  AOI22_X1 U21509 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18424), .B1(
        n18606), .B2(n18496), .ZN(n18411) );
  OAI211_X1 U21510 ( .C1(n18609), .C2(n18421), .A(n18412), .B(n18411), .ZN(
        P3_U2934) );
  AOI22_X1 U21511 ( .A1(n18610), .A2(n18422), .B1(n18564), .B2(n18437), .ZN(
        n18414) );
  AOI22_X1 U21512 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18424), .B1(
        n18612), .B2(n18496), .ZN(n18413) );
  OAI211_X1 U21513 ( .C1(n18567), .C2(n18421), .A(n18414), .B(n18413), .ZN(
        P3_U2935) );
  INV_X1 U21514 ( .A(n18437), .ZN(n18444) );
  AOI22_X1 U21515 ( .A1(n18617), .A2(n18423), .B1(n18616), .B2(n18422), .ZN(
        n18416) );
  AOI22_X1 U21516 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18424), .B1(
        n18618), .B2(n18496), .ZN(n18415) );
  OAI211_X1 U21517 ( .C1(n18621), .C2(n18444), .A(n18416), .B(n18415), .ZN(
        P3_U2936) );
  AOI22_X1 U21518 ( .A1(n18622), .A2(n18422), .B1(n18570), .B2(n18437), .ZN(
        n18418) );
  AOI22_X1 U21519 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18424), .B1(
        n18624), .B2(n18496), .ZN(n18417) );
  OAI211_X1 U21520 ( .C1(n18573), .C2(n18421), .A(n18418), .B(n18417), .ZN(
        P3_U2937) );
  AOI22_X1 U21521 ( .A1(n18629), .A2(n18437), .B1(n18628), .B2(n18422), .ZN(
        n18420) );
  AOI22_X1 U21522 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18424), .B1(
        n18631), .B2(n18496), .ZN(n18419) );
  OAI211_X1 U21523 ( .C1(n18635), .C2(n18421), .A(n18420), .B(n18419), .ZN(
        P3_U2938) );
  AOI22_X1 U21524 ( .A1(n18639), .A2(n18423), .B1(n18637), .B2(n18422), .ZN(
        n18426) );
  AOI22_X1 U21525 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18424), .B1(
        n18640), .B2(n18496), .ZN(n18425) );
  OAI211_X1 U21526 ( .C1(n18645), .C2(n18444), .A(n18426), .B(n18425), .ZN(
        P3_U2939) );
  INV_X1 U21527 ( .A(n18473), .ZN(n18471) );
  AOI22_X1 U21528 ( .A1(n18589), .A2(n18437), .B1(n18588), .B2(n18447), .ZN(
        n18432) );
  NOR2_X1 U21529 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18427), .ZN(
        n18429) );
  NOR2_X1 U21530 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18479), .ZN(
        n18428) );
  AOI22_X1 U21531 ( .A1(n18593), .A2(n18429), .B1(n18591), .B2(n18428), .ZN(
        n18448) );
  NOR2_X2 U21532 ( .A1(n18430), .A2(n18479), .ZN(n18523) );
  AOI22_X1 U21533 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18448), .B1(
        n18594), .B2(n18523), .ZN(n18431) );
  OAI211_X1 U21534 ( .C1(n18597), .C2(n18471), .A(n18432), .B(n18431), .ZN(
        P3_U2940) );
  AOI22_X1 U21535 ( .A1(n18599), .A2(n18473), .B1(n18598), .B2(n18447), .ZN(
        n18434) );
  AOI22_X1 U21536 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18448), .B1(
        n18600), .B2(n18523), .ZN(n18433) );
  OAI211_X1 U21537 ( .C1(n18603), .C2(n18444), .A(n18434), .B(n18433), .ZN(
        P3_U2941) );
  AOI22_X1 U21538 ( .A1(n18605), .A2(n18473), .B1(n18604), .B2(n18447), .ZN(
        n18436) );
  AOI22_X1 U21539 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18448), .B1(
        n18606), .B2(n18523), .ZN(n18435) );
  OAI211_X1 U21540 ( .C1(n18609), .C2(n18444), .A(n18436), .B(n18435), .ZN(
        P3_U2942) );
  AOI22_X1 U21541 ( .A1(n18611), .A2(n18437), .B1(n18610), .B2(n18447), .ZN(
        n18439) );
  AOI22_X1 U21542 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18448), .B1(
        n18612), .B2(n18523), .ZN(n18438) );
  OAI211_X1 U21543 ( .C1(n18615), .C2(n18471), .A(n18439), .B(n18438), .ZN(
        P3_U2943) );
  AOI22_X1 U21544 ( .A1(n18617), .A2(n18437), .B1(n18616), .B2(n18447), .ZN(
        n18441) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18448), .B1(
        n18618), .B2(n18523), .ZN(n18440) );
  OAI211_X1 U21546 ( .C1(n18621), .C2(n18471), .A(n18441), .B(n18440), .ZN(
        P3_U2944) );
  AOI22_X1 U21547 ( .A1(n18622), .A2(n18447), .B1(n18570), .B2(n18473), .ZN(
        n18443) );
  AOI22_X1 U21548 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18448), .B1(
        n18624), .B2(n18523), .ZN(n18442) );
  OAI211_X1 U21549 ( .C1(n18573), .C2(n18444), .A(n18443), .B(n18442), .ZN(
        P3_U2945) );
  AOI22_X1 U21550 ( .A1(n18628), .A2(n18447), .B1(n18575), .B2(n18437), .ZN(
        n18446) );
  AOI22_X1 U21551 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18448), .B1(
        n18631), .B2(n18523), .ZN(n18445) );
  OAI211_X1 U21552 ( .C1(n18578), .C2(n18471), .A(n18446), .B(n18445), .ZN(
        P3_U2946) );
  AOI22_X1 U21553 ( .A1(n18639), .A2(n18437), .B1(n18637), .B2(n18447), .ZN(
        n18450) );
  AOI22_X1 U21554 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18448), .B1(
        n18640), .B2(n18523), .ZN(n18449) );
  OAI211_X1 U21555 ( .C1(n18645), .C2(n18471), .A(n18450), .B(n18449), .ZN(
        P3_U2947) );
  INV_X1 U21556 ( .A(n18496), .ZN(n18494) );
  INV_X1 U21557 ( .A(n18523), .ZN(n18515) );
  NOR2_X2 U21558 ( .A1(n18451), .A2(n18479), .ZN(n18546) );
  INV_X1 U21559 ( .A(n18546), .ZN(n18544) );
  AOI21_X1 U21560 ( .B1(n18515), .B2(n18544), .A(n18713), .ZN(n18472) );
  AOI22_X1 U21561 ( .A1(n18589), .A2(n18473), .B1(n18588), .B2(n18472), .ZN(
        n18458) );
  NOR2_X1 U21562 ( .A1(n18523), .A2(n18546), .ZN(n18453) );
  OAI22_X1 U21563 ( .A1(n18455), .A2(n18454), .B1(n18453), .B2(n18452), .ZN(
        n18456) );
  OAI21_X1 U21564 ( .B1(n18546), .B2(n18808), .A(n18456), .ZN(n18474) );
  AOI22_X1 U21565 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18474), .B1(
        n18594), .B2(n18546), .ZN(n18457) );
  OAI211_X1 U21566 ( .C1(n18597), .C2(n18494), .A(n18458), .B(n18457), .ZN(
        P3_U2948) );
  AOI22_X1 U21567 ( .A1(n18599), .A2(n18496), .B1(n18598), .B2(n18472), .ZN(
        n18460) );
  AOI22_X1 U21568 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18474), .B1(
        n18600), .B2(n18546), .ZN(n18459) );
  OAI211_X1 U21569 ( .C1(n18603), .C2(n18471), .A(n18460), .B(n18459), .ZN(
        P3_U2949) );
  AOI22_X1 U21570 ( .A1(n18605), .A2(n18496), .B1(n18604), .B2(n18472), .ZN(
        n18462) );
  AOI22_X1 U21571 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18474), .B1(
        n18606), .B2(n18546), .ZN(n18461) );
  OAI211_X1 U21572 ( .C1(n18609), .C2(n18471), .A(n18462), .B(n18461), .ZN(
        P3_U2950) );
  AOI22_X1 U21573 ( .A1(n18611), .A2(n18473), .B1(n18610), .B2(n18472), .ZN(
        n18464) );
  AOI22_X1 U21574 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18474), .B1(
        n18612), .B2(n18546), .ZN(n18463) );
  OAI211_X1 U21575 ( .C1(n18615), .C2(n18494), .A(n18464), .B(n18463), .ZN(
        P3_U2951) );
  AOI22_X1 U21576 ( .A1(n18512), .A2(n18496), .B1(n18616), .B2(n18472), .ZN(
        n18466) );
  AOI22_X1 U21577 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18474), .B1(
        n18618), .B2(n18546), .ZN(n18465) );
  OAI211_X1 U21578 ( .C1(n18516), .C2(n18471), .A(n18466), .B(n18465), .ZN(
        P3_U2952) );
  AOI22_X1 U21579 ( .A1(n18623), .A2(n18473), .B1(n18622), .B2(n18472), .ZN(
        n18468) );
  AOI22_X1 U21580 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18474), .B1(
        n18624), .B2(n18546), .ZN(n18467) );
  OAI211_X1 U21581 ( .C1(n18627), .C2(n18494), .A(n18468), .B(n18467), .ZN(
        P3_U2953) );
  AOI22_X1 U21582 ( .A1(n18629), .A2(n18496), .B1(n18628), .B2(n18472), .ZN(
        n18470) );
  AOI22_X1 U21583 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18474), .B1(
        n18631), .B2(n18546), .ZN(n18469) );
  OAI211_X1 U21584 ( .C1(n18635), .C2(n18471), .A(n18470), .B(n18469), .ZN(
        P3_U2954) );
  AOI22_X1 U21585 ( .A1(n18639), .A2(n18473), .B1(n18637), .B2(n18472), .ZN(
        n18476) );
  AOI22_X1 U21586 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18474), .B1(
        n18640), .B2(n18546), .ZN(n18475) );
  OAI211_X1 U21587 ( .C1(n18645), .C2(n18494), .A(n18476), .B(n18475), .ZN(
        P3_U2955) );
  NOR2_X1 U21588 ( .A1(n18659), .A2(n18479), .ZN(n18527) );
  INV_X1 U21589 ( .A(n18527), .ZN(n18477) );
  NOR2_X1 U21590 ( .A1(n18713), .A2(n18477), .ZN(n18495) );
  AOI22_X1 U21591 ( .A1(n18551), .A2(n18523), .B1(n18588), .B2(n18495), .ZN(
        n18481) );
  OAI211_X1 U21592 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18593), .A(
        n18591), .B(n18478), .ZN(n18497) );
  NOR2_X2 U21593 ( .A1(n18658), .A2(n18479), .ZN(n18574) );
  AOI22_X1 U21594 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18497), .B1(
        n18594), .B2(n18574), .ZN(n18480) );
  OAI211_X1 U21595 ( .C1(n18557), .C2(n18494), .A(n18481), .B(n18480), .ZN(
        P3_U2956) );
  AOI22_X1 U21596 ( .A1(n18599), .A2(n18523), .B1(n18598), .B2(n18495), .ZN(
        n18483) );
  AOI22_X1 U21597 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18497), .B1(
        n18600), .B2(n18574), .ZN(n18482) );
  OAI211_X1 U21598 ( .C1(n18603), .C2(n18494), .A(n18483), .B(n18482), .ZN(
        P3_U2957) );
  AOI22_X1 U21599 ( .A1(n18560), .A2(n18496), .B1(n18604), .B2(n18495), .ZN(
        n18485) );
  AOI22_X1 U21600 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18497), .B1(
        n18606), .B2(n18574), .ZN(n18484) );
  OAI211_X1 U21601 ( .C1(n18563), .C2(n18515), .A(n18485), .B(n18484), .ZN(
        P3_U2958) );
  AOI22_X1 U21602 ( .A1(n18610), .A2(n18495), .B1(n18564), .B2(n18523), .ZN(
        n18487) );
  AOI22_X1 U21603 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18497), .B1(
        n18612), .B2(n18574), .ZN(n18486) );
  OAI211_X1 U21604 ( .C1(n18567), .C2(n18494), .A(n18487), .B(n18486), .ZN(
        P3_U2959) );
  AOI22_X1 U21605 ( .A1(n18617), .A2(n18496), .B1(n18616), .B2(n18495), .ZN(
        n18489) );
  AOI22_X1 U21606 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18497), .B1(
        n18618), .B2(n18574), .ZN(n18488) );
  OAI211_X1 U21607 ( .C1(n18621), .C2(n18515), .A(n18489), .B(n18488), .ZN(
        P3_U2960) );
  AOI22_X1 U21608 ( .A1(n18622), .A2(n18495), .B1(n18570), .B2(n18523), .ZN(
        n18491) );
  AOI22_X1 U21609 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18497), .B1(
        n18624), .B2(n18574), .ZN(n18490) );
  OAI211_X1 U21610 ( .C1(n18573), .C2(n18494), .A(n18491), .B(n18490), .ZN(
        P3_U2961) );
  AOI22_X1 U21611 ( .A1(n18629), .A2(n18523), .B1(n18628), .B2(n18495), .ZN(
        n18493) );
  AOI22_X1 U21612 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18497), .B1(
        n18631), .B2(n18574), .ZN(n18492) );
  OAI211_X1 U21613 ( .C1(n18635), .C2(n18494), .A(n18493), .B(n18492), .ZN(
        P3_U2962) );
  AOI22_X1 U21614 ( .A1(n18639), .A2(n18496), .B1(n18637), .B2(n18495), .ZN(
        n18499) );
  AOI22_X1 U21615 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18497), .B1(
        n18640), .B2(n18574), .ZN(n18498) );
  OAI211_X1 U21616 ( .C1(n18645), .C2(n18515), .A(n18499), .B(n18498), .ZN(
        P3_U2963) );
  NAND2_X1 U21617 ( .A1(n21027), .A2(n18592), .ZN(n18634) );
  INV_X1 U21618 ( .A(n18634), .ZN(n18638) );
  NOR2_X1 U21619 ( .A1(n18574), .A2(n18638), .ZN(n18552) );
  NOR2_X1 U21620 ( .A1(n18713), .A2(n18552), .ZN(n18521) );
  AOI22_X1 U21621 ( .A1(n18551), .A2(n18546), .B1(n18588), .B2(n18521), .ZN(
        n18505) );
  OAI21_X1 U21622 ( .B1(n18501), .B2(n18500), .A(n18552), .ZN(n18502) );
  OAI211_X1 U21623 ( .C1(n18638), .C2(n18808), .A(n18503), .B(n18502), .ZN(
        n18522) );
  AOI22_X1 U21624 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18522), .B1(
        n18594), .B2(n18638), .ZN(n18504) );
  OAI211_X1 U21625 ( .C1(n18557), .C2(n18515), .A(n18505), .B(n18504), .ZN(
        P3_U2964) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18522), .B1(
        n18598), .B2(n18521), .ZN(n18507) );
  AOI22_X1 U21627 ( .A1(n18600), .A2(n18638), .B1(n18599), .B2(n18546), .ZN(
        n18506) );
  OAI211_X1 U21628 ( .C1(n18603), .C2(n18515), .A(n18507), .B(n18506), .ZN(
        P3_U2965) );
  AOI22_X1 U21629 ( .A1(n18605), .A2(n18546), .B1(n18604), .B2(n18521), .ZN(
        n18509) );
  AOI22_X1 U21630 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18522), .B1(
        n18606), .B2(n18638), .ZN(n18508) );
  OAI211_X1 U21631 ( .C1(n18609), .C2(n18515), .A(n18509), .B(n18508), .ZN(
        P3_U2966) );
  AOI22_X1 U21632 ( .A1(n18611), .A2(n18523), .B1(n18610), .B2(n18521), .ZN(
        n18511) );
  AOI22_X1 U21633 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18522), .B1(
        n18612), .B2(n18638), .ZN(n18510) );
  OAI211_X1 U21634 ( .C1(n18615), .C2(n18544), .A(n18511), .B(n18510), .ZN(
        P3_U2967) );
  AOI22_X1 U21635 ( .A1(n18512), .A2(n18546), .B1(n18616), .B2(n18521), .ZN(
        n18514) );
  AOI22_X1 U21636 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18522), .B1(
        n18618), .B2(n18638), .ZN(n18513) );
  OAI211_X1 U21637 ( .C1(n18516), .C2(n18515), .A(n18514), .B(n18513), .ZN(
        P3_U2968) );
  AOI22_X1 U21638 ( .A1(n18623), .A2(n18523), .B1(n18622), .B2(n18521), .ZN(
        n18518) );
  AOI22_X1 U21639 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18522), .B1(
        n18624), .B2(n18638), .ZN(n18517) );
  OAI211_X1 U21640 ( .C1(n18627), .C2(n18544), .A(n18518), .B(n18517), .ZN(
        P3_U2969) );
  AOI22_X1 U21641 ( .A1(n18628), .A2(n18521), .B1(n18575), .B2(n18523), .ZN(
        n18520) );
  AOI22_X1 U21642 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18522), .B1(
        n18631), .B2(n18638), .ZN(n18519) );
  OAI211_X1 U21643 ( .C1(n18578), .C2(n18544), .A(n18520), .B(n18519), .ZN(
        P3_U2970) );
  AOI22_X1 U21644 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18522), .B1(
        n18637), .B2(n18521), .ZN(n18525) );
  AOI22_X1 U21645 ( .A1(n18639), .A2(n18523), .B1(n18640), .B2(n18638), .ZN(
        n18524) );
  OAI211_X1 U21646 ( .C1(n18645), .C2(n18544), .A(n18525), .B(n18524), .ZN(
        P3_U2971) );
  INV_X1 U21647 ( .A(n18592), .ZN(n18526) );
  NOR2_X1 U21648 ( .A1(n18713), .A2(n18526), .ZN(n18545) );
  AOI22_X1 U21649 ( .A1(n18551), .A2(n18574), .B1(n18588), .B2(n18545), .ZN(
        n18529) );
  AOI22_X1 U21650 ( .A1(n18593), .A2(n18527), .B1(n18592), .B2(n18591), .ZN(
        n18547) );
  AOI22_X1 U21651 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18547), .B1(
        n18594), .B2(n18630), .ZN(n18528) );
  OAI211_X1 U21652 ( .C1(n18557), .C2(n18544), .A(n18529), .B(n18528), .ZN(
        P3_U2972) );
  INV_X1 U21653 ( .A(n18600), .ZN(n18533) );
  AOI22_X1 U21654 ( .A1(n18530), .A2(n18546), .B1(n18598), .B2(n18545), .ZN(
        n18532) );
  AOI22_X1 U21655 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18547), .B1(
        n18599), .B2(n18574), .ZN(n18531) );
  OAI211_X1 U21656 ( .C1(n18646), .C2(n18533), .A(n18532), .B(n18531), .ZN(
        P3_U2973) );
  AOI22_X1 U21657 ( .A1(n18605), .A2(n18574), .B1(n18604), .B2(n18545), .ZN(
        n18535) );
  AOI22_X1 U21658 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18547), .B1(
        n18630), .B2(n18606), .ZN(n18534) );
  OAI211_X1 U21659 ( .C1(n18609), .C2(n18544), .A(n18535), .B(n18534), .ZN(
        P3_U2974) );
  INV_X1 U21660 ( .A(n18574), .ZN(n18585) );
  AOI22_X1 U21661 ( .A1(n18611), .A2(n18546), .B1(n18610), .B2(n18545), .ZN(
        n18537) );
  AOI22_X1 U21662 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18547), .B1(
        n18630), .B2(n18612), .ZN(n18536) );
  OAI211_X1 U21663 ( .C1(n18615), .C2(n18585), .A(n18537), .B(n18536), .ZN(
        P3_U2975) );
  AOI22_X1 U21664 ( .A1(n18617), .A2(n18546), .B1(n18616), .B2(n18545), .ZN(
        n18539) );
  AOI22_X1 U21665 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18547), .B1(
        n18630), .B2(n18618), .ZN(n18538) );
  OAI211_X1 U21666 ( .C1(n18621), .C2(n18585), .A(n18539), .B(n18538), .ZN(
        P3_U2976) );
  AOI22_X1 U21667 ( .A1(n18623), .A2(n18546), .B1(n18622), .B2(n18545), .ZN(
        n18541) );
  AOI22_X1 U21668 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18547), .B1(
        n18630), .B2(n18624), .ZN(n18540) );
  OAI211_X1 U21669 ( .C1(n18627), .C2(n18585), .A(n18541), .B(n18540), .ZN(
        P3_U2977) );
  AOI22_X1 U21670 ( .A1(n18629), .A2(n18574), .B1(n18628), .B2(n18545), .ZN(
        n18543) );
  AOI22_X1 U21671 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18547), .B1(
        n18630), .B2(n18631), .ZN(n18542) );
  OAI211_X1 U21672 ( .C1(n18635), .C2(n18544), .A(n18543), .B(n18542), .ZN(
        P3_U2978) );
  AOI22_X1 U21673 ( .A1(n18639), .A2(n18546), .B1(n18637), .B2(n18545), .ZN(
        n18549) );
  AOI22_X1 U21674 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18547), .B1(
        n18630), .B2(n18640), .ZN(n18548) );
  OAI211_X1 U21675 ( .C1(n18645), .C2(n18585), .A(n18549), .B(n18548), .ZN(
        P3_U2979) );
  NOR2_X1 U21676 ( .A1(n18713), .A2(n18550), .ZN(n18579) );
  AOI22_X1 U21677 ( .A1(n18551), .A2(n18638), .B1(n18588), .B2(n18579), .ZN(
        n18556) );
  NOR2_X1 U21678 ( .A1(n18552), .A2(n18454), .ZN(n18553) );
  OAI22_X1 U21679 ( .A1(n18581), .A2(n18808), .B1(n18554), .B2(n18553), .ZN(
        n18582) );
  AOI22_X1 U21680 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18582), .B1(
        n18581), .B2(n18594), .ZN(n18555) );
  OAI211_X1 U21681 ( .C1(n18557), .C2(n18585), .A(n18556), .B(n18555), .ZN(
        P3_U2980) );
  AOI22_X1 U21682 ( .A1(n18599), .A2(n18638), .B1(n18598), .B2(n18579), .ZN(
        n18559) );
  AOI22_X1 U21683 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18582), .B1(
        n18581), .B2(n18600), .ZN(n18558) );
  OAI211_X1 U21684 ( .C1(n18603), .C2(n18585), .A(n18559), .B(n18558), .ZN(
        P3_U2981) );
  AOI22_X1 U21685 ( .A1(n18560), .A2(n18574), .B1(n18604), .B2(n18579), .ZN(
        n18562) );
  AOI22_X1 U21686 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18582), .B1(
        n18581), .B2(n18606), .ZN(n18561) );
  OAI211_X1 U21687 ( .C1(n18563), .C2(n18634), .A(n18562), .B(n18561), .ZN(
        P3_U2982) );
  AOI22_X1 U21688 ( .A1(n18610), .A2(n18579), .B1(n18564), .B2(n18638), .ZN(
        n18566) );
  AOI22_X1 U21689 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18582), .B1(
        n18581), .B2(n18612), .ZN(n18565) );
  OAI211_X1 U21690 ( .C1(n18567), .C2(n18585), .A(n18566), .B(n18565), .ZN(
        P3_U2983) );
  AOI22_X1 U21691 ( .A1(n18617), .A2(n18574), .B1(n18616), .B2(n18579), .ZN(
        n18569) );
  AOI22_X1 U21692 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18582), .B1(
        n18581), .B2(n18618), .ZN(n18568) );
  OAI211_X1 U21693 ( .C1(n18621), .C2(n18634), .A(n18569), .B(n18568), .ZN(
        P3_U2984) );
  AOI22_X1 U21694 ( .A1(n18622), .A2(n18579), .B1(n18570), .B2(n18638), .ZN(
        n18572) );
  AOI22_X1 U21695 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18582), .B1(
        n18581), .B2(n18624), .ZN(n18571) );
  OAI211_X1 U21696 ( .C1(n18573), .C2(n18585), .A(n18572), .B(n18571), .ZN(
        P3_U2985) );
  AOI22_X1 U21697 ( .A1(n18628), .A2(n18579), .B1(n18575), .B2(n18574), .ZN(
        n18577) );
  AOI22_X1 U21698 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18582), .B1(
        n18581), .B2(n18631), .ZN(n18576) );
  OAI211_X1 U21699 ( .C1(n18578), .C2(n18634), .A(n18577), .B(n18576), .ZN(
        P3_U2986) );
  AOI22_X1 U21700 ( .A1(n18580), .A2(n18638), .B1(n18637), .B2(n18579), .ZN(
        n18584) );
  AOI22_X1 U21701 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18582), .B1(
        n18581), .B2(n18640), .ZN(n18583) );
  OAI211_X1 U21702 ( .C1(n18586), .C2(n18585), .A(n18584), .B(n18583), .ZN(
        P3_U2987) );
  INV_X1 U21703 ( .A(n18590), .ZN(n18587) );
  NOR2_X1 U21704 ( .A1(n18713), .A2(n18587), .ZN(n18636) );
  AOI22_X1 U21705 ( .A1(n18589), .A2(n18638), .B1(n18588), .B2(n18636), .ZN(
        n18596) );
  AOI22_X1 U21706 ( .A1(n18593), .A2(n18592), .B1(n18591), .B2(n18590), .ZN(
        n18642) );
  AOI22_X1 U21707 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18642), .B1(
        n18641), .B2(n18594), .ZN(n18595) );
  OAI211_X1 U21708 ( .C1(n18597), .C2(n18646), .A(n18596), .B(n18595), .ZN(
        P3_U2988) );
  AOI22_X1 U21709 ( .A1(n18630), .A2(n18599), .B1(n18598), .B2(n18636), .ZN(
        n18602) );
  AOI22_X1 U21710 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18642), .B1(
        n18641), .B2(n18600), .ZN(n18601) );
  OAI211_X1 U21711 ( .C1(n18603), .C2(n18634), .A(n18602), .B(n18601), .ZN(
        P3_U2989) );
  AOI22_X1 U21712 ( .A1(n18630), .A2(n18605), .B1(n18604), .B2(n18636), .ZN(
        n18608) );
  AOI22_X1 U21713 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18642), .B1(
        n18641), .B2(n18606), .ZN(n18607) );
  OAI211_X1 U21714 ( .C1(n18609), .C2(n18634), .A(n18608), .B(n18607), .ZN(
        P3_U2990) );
  AOI22_X1 U21715 ( .A1(n18611), .A2(n18638), .B1(n18610), .B2(n18636), .ZN(
        n18614) );
  AOI22_X1 U21716 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18642), .B1(
        n18641), .B2(n18612), .ZN(n18613) );
  OAI211_X1 U21717 ( .C1(n18646), .C2(n18615), .A(n18614), .B(n18613), .ZN(
        P3_U2991) );
  AOI22_X1 U21718 ( .A1(n18617), .A2(n18638), .B1(n18616), .B2(n18636), .ZN(
        n18620) );
  AOI22_X1 U21719 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18642), .B1(
        n18641), .B2(n18618), .ZN(n18619) );
  OAI211_X1 U21720 ( .C1(n18646), .C2(n18621), .A(n18620), .B(n18619), .ZN(
        P3_U2992) );
  AOI22_X1 U21721 ( .A1(n18623), .A2(n18638), .B1(n18622), .B2(n18636), .ZN(
        n18626) );
  AOI22_X1 U21722 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18642), .B1(
        n18641), .B2(n18624), .ZN(n18625) );
  OAI211_X1 U21723 ( .C1(n18646), .C2(n18627), .A(n18626), .B(n18625), .ZN(
        P3_U2993) );
  AOI22_X1 U21724 ( .A1(n18630), .A2(n18629), .B1(n18628), .B2(n18636), .ZN(
        n18633) );
  AOI22_X1 U21725 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18642), .B1(
        n18641), .B2(n18631), .ZN(n18632) );
  OAI211_X1 U21726 ( .C1(n18635), .C2(n18634), .A(n18633), .B(n18632), .ZN(
        P3_U2994) );
  AOI22_X1 U21727 ( .A1(n18639), .A2(n18638), .B1(n18637), .B2(n18636), .ZN(
        n18644) );
  AOI22_X1 U21728 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18642), .B1(
        n18641), .B2(n18640), .ZN(n18643) );
  OAI211_X1 U21729 ( .C1(n18646), .C2(n18645), .A(n18644), .B(n18643), .ZN(
        P3_U2995) );
  NOR2_X1 U21730 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18698) );
  NOR2_X1 U21731 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18647), .ZN(
        n18667) );
  OAI21_X1 U21732 ( .B1(n18827), .B2(n18667), .A(n18820), .ZN(n18652) );
  AOI22_X1 U21733 ( .A1(n18648), .A2(n9832), .B1(n18647), .B2(n18666), .ZN(
        n18650) );
  AOI21_X1 U21734 ( .B1(n18651), .B2(n18650), .A(n18649), .ZN(n18670) );
  NAND2_X1 U21735 ( .A1(n18652), .A2(n18670), .ZN(n18653) );
  OAI21_X1 U21736 ( .B1(n18816), .B2(n18685), .A(n18653), .ZN(n18818) );
  AOI22_X1 U21737 ( .A1(n18691), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n18818), .B2(n18677), .ZN(n18674) );
  INV_X1 U21738 ( .A(n18674), .ZN(n18664) );
  NOR2_X1 U21739 ( .A1(n18655), .A2(n18654), .ZN(n18657) );
  AOI22_X1 U21740 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18656), .B1(
        n18657), .B2(n21023), .ZN(n18829) );
  OAI22_X1 U21741 ( .A1(n18657), .A2(n18821), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18667), .ZN(n18825) );
  AOI222_X1 U21742 ( .A1(n18829), .A2(n18825), .B1(n18829), .B2(n18659), .C1(
        n18825), .C2(n18658), .ZN(n18661) );
  OAI21_X1 U21743 ( .B1(n18691), .B2(n18661), .A(n18660), .ZN(n18662) );
  OAI21_X1 U21744 ( .B1(n18664), .B2(n18663), .A(n18662), .ZN(n18675) );
  OAI21_X1 U21745 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18674), .A(
        n18675), .ZN(n18697) );
  AND2_X1 U21746 ( .A1(n18820), .A2(n18665), .ZN(n18669) );
  OAI22_X1 U21747 ( .A1(n18669), .A2(n18685), .B1(n18667), .B2(n18666), .ZN(
        n18668) );
  INV_X1 U21748 ( .A(n18668), .ZN(n18672) );
  NOR2_X1 U21749 ( .A1(n18670), .A2(n18669), .ZN(n18671) );
  MUX2_X1 U21750 ( .A(n18672), .B(n18671), .S(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n18673) );
  INV_X1 U21751 ( .A(n18673), .ZN(n18810) );
  OAI221_X1 U21752 ( .B1(n18675), .B2(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), 
        .C1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(n18674), .ZN(n18676) );
  OAI221_X1 U21753 ( .B1(n18677), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .C1(n18691), .C2(n18810), .A(n18676), .ZN(n18678) );
  INV_X1 U21754 ( .A(n18678), .ZN(n18696) );
  NOR2_X1 U21755 ( .A1(P3_MORE_REG_SCAN_IN), .A2(P3_FLUSH_REG_SCAN_IN), .ZN(
        n18694) );
  OAI221_X1 U21756 ( .B1(n18682), .B2(n18681), .C1(n18682), .C2(n18680), .A(
        n18679), .ZN(n18687) );
  AOI21_X1 U21757 ( .B1(n18685), .B2(n18684), .A(n18683), .ZN(n18686) );
  AOI21_X1 U21758 ( .B1(n18688), .B2(n18687), .A(n18686), .ZN(n18845) );
  AOI211_X1 U21759 ( .C1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(n18691), .A(
        n18690), .B(n18689), .ZN(n18692) );
  OAI211_X1 U21760 ( .C1(n18694), .C2(n18693), .A(n18845), .B(n18692), .ZN(
        n18695) );
  AOI211_X1 U21761 ( .C1(n18698), .C2(n18697), .A(n18696), .B(n18695), .ZN(
        n18709) );
  AOI22_X1 U21762 ( .A1(n18828), .A2(n18857), .B1(n18710), .B2(n17440), .ZN(
        n18699) );
  INV_X1 U21763 ( .A(n18699), .ZN(n18705) );
  INV_X1 U21764 ( .A(n18700), .ZN(n18702) );
  OAI211_X1 U21765 ( .C1(n18702), .C2(n18701), .A(n18849), .B(n18709), .ZN(
        n18807) );
  OAI21_X1 U21766 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18854), .A(n18807), 
        .ZN(n18711) );
  NOR2_X1 U21767 ( .A1(n18703), .A2(n18711), .ZN(n18704) );
  MUX2_X1 U21768 ( .A(n18705), .B(n18704), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18707) );
  OAI211_X1 U21769 ( .C1(n18709), .C2(n18708), .A(n18707), .B(n18706), .ZN(
        P3_U2996) );
  NAND2_X1 U21770 ( .A1(n18710), .A2(n17440), .ZN(n18716) );
  NOR4_X1 U21771 ( .A1(n18813), .A2(n20757), .A3(n18854), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18719) );
  INV_X1 U21772 ( .A(n18719), .ZN(n18715) );
  OR3_X1 U21773 ( .A1(n18713), .A2(n18712), .A3(n18711), .ZN(n18714) );
  NAND4_X1 U21774 ( .A1(n18717), .A2(n18716), .A3(n18715), .A4(n18714), .ZN(
        P3_U2997) );
  OAI21_X1 U21775 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18718), .ZN(n18720) );
  AOI21_X1 U21776 ( .B1(n18721), .B2(n18720), .A(n18719), .ZN(P3_U2998) );
  AND2_X1 U21777 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18802), .ZN(
        P3_U2999) );
  AND2_X1 U21778 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18802), .ZN(
        P3_U3000) );
  AND2_X1 U21779 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18802), .ZN(
        P3_U3001) );
  AND2_X1 U21780 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18802), .ZN(
        P3_U3002) );
  AND2_X1 U21781 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18802), .ZN(
        P3_U3003) );
  AND2_X1 U21782 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18802), .ZN(
        P3_U3004) );
  AND2_X1 U21783 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18802), .ZN(
        P3_U3005) );
  AND2_X1 U21784 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18802), .ZN(
        P3_U3006) );
  AND2_X1 U21785 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18802), .ZN(
        P3_U3007) );
  AND2_X1 U21786 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18802), .ZN(
        P3_U3008) );
  AND2_X1 U21787 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18802), .ZN(
        P3_U3009) );
  AND2_X1 U21788 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18802), .ZN(
        P3_U3010) );
  AND2_X1 U21789 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18802), .ZN(
        P3_U3011) );
  AND2_X1 U21790 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18802), .ZN(
        P3_U3012) );
  AND2_X1 U21791 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18802), .ZN(
        P3_U3013) );
  AND2_X1 U21792 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18802), .ZN(
        P3_U3014) );
  AND2_X1 U21793 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18802), .ZN(
        P3_U3015) );
  AND2_X1 U21794 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18802), .ZN(
        P3_U3016) );
  AND2_X1 U21795 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18802), .ZN(
        P3_U3017) );
  INV_X1 U21796 ( .A(P3_DATAWIDTH_REG_12__SCAN_IN), .ZN(n20835) );
  NOR2_X1 U21797 ( .A1(n20835), .A2(n18805), .ZN(P3_U3018) );
  AND2_X1 U21798 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18802), .ZN(
        P3_U3019) );
  AND2_X1 U21799 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18802), .ZN(
        P3_U3020) );
  AND2_X1 U21800 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18802), .ZN(P3_U3021) );
  AND2_X1 U21801 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18802), .ZN(P3_U3022) );
  AND2_X1 U21802 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18802), .ZN(P3_U3023) );
  AND2_X1 U21803 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18802), .ZN(P3_U3024) );
  AND2_X1 U21804 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18802), .ZN(P3_U3025) );
  AND2_X1 U21805 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18802), .ZN(P3_U3026) );
  AND2_X1 U21806 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18802), .ZN(P3_U3027) );
  AND2_X1 U21807 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18802), .ZN(P3_U3028) );
  NOR2_X1 U21808 ( .A1(n18737), .A2(n19750), .ZN(n18732) );
  INV_X1 U21809 ( .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18722) );
  NOR2_X1 U21810 ( .A1(n18732), .A2(n18722), .ZN(n18727) );
  OAI21_X1 U21811 ( .B1(n18728), .B2(n19750), .A(n18727), .ZN(n18723) );
  AOI22_X1 U21812 ( .A1(n20922), .A2(n18737), .B1(n18863), .B2(n18723), .ZN(
        n18724) );
  NAND3_X1 U21813 ( .A1(NA), .A2(n20922), .A3(n18728), .ZN(n18733) );
  OAI211_X1 U21814 ( .C1(n18854), .C2(n18725), .A(n18724), .B(n18733), .ZN(
        P3_U3029) );
  NOR2_X1 U21815 ( .A1(n18728), .A2(n19750), .ZN(n18726) );
  AOI22_X1 U21816 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18727), .B1(n18726), 
        .B2(n18737), .ZN(n18729) );
  NOR2_X1 U21817 ( .A1(n18854), .A2(n18728), .ZN(n18734) );
  INV_X1 U21818 ( .A(n18734), .ZN(n18730) );
  NAND3_X1 U21819 ( .A1(n18729), .A2(n18851), .A3(n18730), .ZN(P3_U3030) );
  OAI22_X1 U21820 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18730), .ZN(n18731) );
  OAI22_X1 U21821 ( .A1(n18732), .A2(n18731), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18736) );
  OAI211_X1 U21822 ( .C1(n18734), .C2(n20922), .A(n18733), .B(
        P3_STATE_REG_2__SCAN_IN), .ZN(n18735) );
  OAI21_X1 U21823 ( .B1(n20922), .B2(n18736), .A(n18735), .ZN(P3_U3031) );
  INV_X1 U21824 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18740) );
  OAI222_X1 U21825 ( .A1(n18739), .A2(n18796), .B1(n18738), .B2(n18793), .C1(
        n18740), .C2(n18781), .ZN(P3_U3032) );
  INV_X1 U21826 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18742) );
  INV_X1 U21827 ( .A(n18863), .ZN(n18862) );
  OAI222_X1 U21828 ( .A1(n18781), .A2(n18742), .B1(n18741), .B2(n18862), .C1(
        n18740), .C2(n18796), .ZN(P3_U3033) );
  OAI222_X1 U21829 ( .A1(n18781), .A2(n18744), .B1(n18743), .B2(n18793), .C1(
        n18742), .C2(n18796), .ZN(P3_U3034) );
  INV_X1 U21830 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n20851) );
  OAI222_X1 U21831 ( .A1(n18781), .A2(n20851), .B1(n18745), .B2(n18862), .C1(
        n18744), .C2(n18796), .ZN(P3_U3035) );
  OAI222_X1 U21832 ( .A1(n18781), .A2(n18747), .B1(n18746), .B2(n18793), .C1(
        n20851), .C2(n18796), .ZN(P3_U3036) );
  OAI222_X1 U21833 ( .A1(n18781), .A2(n18749), .B1(n18748), .B2(n18862), .C1(
        n18747), .C2(n18796), .ZN(P3_U3037) );
  OAI222_X1 U21834 ( .A1(n18781), .A2(n20834), .B1(n20770), .B2(n18862), .C1(
        n18749), .C2(n18796), .ZN(P3_U3038) );
  OAI222_X1 U21835 ( .A1(n20834), .A2(n18796), .B1(n18750), .B2(n18862), .C1(
        n18751), .C2(n18781), .ZN(P3_U3039) );
  OAI222_X1 U21836 ( .A1(n18781), .A2(n18752), .B1(n20812), .B2(n18862), .C1(
        n18751), .C2(n18796), .ZN(P3_U3040) );
  OAI222_X1 U21837 ( .A1(n18781), .A2(n18753), .B1(n21025), .B2(n18862), .C1(
        n18752), .C2(n18796), .ZN(P3_U3041) );
  OAI222_X1 U21838 ( .A1(n18781), .A2(n18755), .B1(n18754), .B2(n18862), .C1(
        n18753), .C2(n18796), .ZN(P3_U3042) );
  OAI222_X1 U21839 ( .A1(n18781), .A2(n18757), .B1(n18756), .B2(n18862), .C1(
        n18755), .C2(n18796), .ZN(P3_U3043) );
  OAI222_X1 U21840 ( .A1(n18781), .A2(n18760), .B1(n18758), .B2(n18862), .C1(
        n18757), .C2(n18796), .ZN(P3_U3044) );
  OAI222_X1 U21841 ( .A1(n18760), .A2(n18796), .B1(n18759), .B2(n18862), .C1(
        n18761), .C2(n18781), .ZN(P3_U3045) );
  OAI222_X1 U21842 ( .A1(n18781), .A2(n18763), .B1(n18762), .B2(n18862), .C1(
        n18761), .C2(n18796), .ZN(P3_U3046) );
  OAI222_X1 U21843 ( .A1(n18781), .A2(n18765), .B1(n18764), .B2(n18862), .C1(
        n18763), .C2(n18796), .ZN(P3_U3047) );
  OAI222_X1 U21844 ( .A1(n18781), .A2(n18767), .B1(n18766), .B2(n18862), .C1(
        n18765), .C2(n18796), .ZN(P3_U3048) );
  OAI222_X1 U21845 ( .A1(n18781), .A2(n18769), .B1(n18768), .B2(n18862), .C1(
        n18767), .C2(n18796), .ZN(P3_U3049) );
  OAI222_X1 U21846 ( .A1(n18781), .A2(n18771), .B1(n18770), .B2(n18862), .C1(
        n18769), .C2(n18796), .ZN(P3_U3050) );
  OAI222_X1 U21847 ( .A1(n18781), .A2(n18773), .B1(n18772), .B2(n18862), .C1(
        n18771), .C2(n18796), .ZN(P3_U3051) );
  OAI222_X1 U21848 ( .A1(n18781), .A2(n18775), .B1(n18774), .B2(n18862), .C1(
        n18773), .C2(n18796), .ZN(P3_U3052) );
  OAI222_X1 U21849 ( .A1(n18781), .A2(n18777), .B1(n18776), .B2(n18862), .C1(
        n18775), .C2(n18796), .ZN(P3_U3053) );
  OAI222_X1 U21850 ( .A1(n18781), .A2(n18779), .B1(n18778), .B2(n18842), .C1(
        n18777), .C2(n18796), .ZN(P3_U3054) );
  OAI222_X1 U21851 ( .A1(n18781), .A2(n18782), .B1(n18780), .B2(n18793), .C1(
        n18779), .C2(n18796), .ZN(P3_U3055) );
  INV_X1 U21852 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18784) );
  OAI222_X1 U21853 ( .A1(n18781), .A2(n18784), .B1(n18783), .B2(n18793), .C1(
        n18782), .C2(n18796), .ZN(P3_U3056) );
  OAI222_X1 U21854 ( .A1(n18781), .A2(n18786), .B1(n18785), .B2(n18793), .C1(
        n18784), .C2(n18796), .ZN(P3_U3057) );
  OAI222_X1 U21855 ( .A1(n18781), .A2(n18789), .B1(n18787), .B2(n18793), .C1(
        n18786), .C2(n18796), .ZN(P3_U3058) );
  OAI222_X1 U21856 ( .A1(n18789), .A2(n18796), .B1(n18788), .B2(n18793), .C1(
        n18790), .C2(n18781), .ZN(P3_U3059) );
  OAI222_X1 U21857 ( .A1(n18781), .A2(n18795), .B1(n18791), .B2(n18793), .C1(
        n18790), .C2(n18796), .ZN(P3_U3060) );
  OAI222_X1 U21858 ( .A1(n18796), .A2(n18795), .B1(n18794), .B2(n18793), .C1(
        n18792), .C2(n18781), .ZN(P3_U3061) );
  OAI22_X1 U21859 ( .A1(n18863), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18862), .ZN(n18797) );
  INV_X1 U21860 ( .A(n18797), .ZN(P3_U3274) );
  OAI22_X1 U21861 ( .A1(n18863), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18862), .ZN(n18798) );
  INV_X1 U21862 ( .A(n18798), .ZN(P3_U3275) );
  OAI22_X1 U21863 ( .A1(n18863), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18862), .ZN(n18799) );
  INV_X1 U21864 ( .A(n18799), .ZN(P3_U3276) );
  OAI22_X1 U21865 ( .A1(n18863), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18862), .ZN(n18800) );
  INV_X1 U21866 ( .A(n18800), .ZN(P3_U3277) );
  INV_X1 U21867 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18834) );
  AOI21_X1 U21868 ( .B1(n18802), .B2(n18834), .A(n18801), .ZN(P3_U3280) );
  INV_X1 U21869 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18804) );
  OAI21_X1 U21870 ( .B1(n18805), .B2(n18804), .A(n18803), .ZN(P3_U3281) );
  OAI221_X1 U21871 ( .B1(n18808), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18808), 
        .C2(n18807), .A(n18806), .ZN(P3_U3282) );
  AOI22_X1 U21872 ( .A1(n18866), .A2(n18810), .B1(n18828), .B2(n18809), .ZN(
        n18811) );
  AOI22_X1 U21873 ( .A1(n18832), .A2(n18812), .B1(n18811), .B2(n18830), .ZN(
        P3_U3285) );
  NOR2_X1 U21874 ( .A1(n18813), .A2(n21021), .ZN(n18822) );
  OAI22_X1 U21875 ( .A1(n18815), .A2(n18814), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18823) );
  INV_X1 U21876 ( .A(n18823), .ZN(n18817) );
  AOI222_X1 U21877 ( .A1(n18818), .A2(n18866), .B1(n18822), .B2(n18817), .C1(
        n18828), .C2(n18816), .ZN(n18819) );
  AOI22_X1 U21878 ( .A1(n18832), .A2(n18820), .B1(n18819), .B2(n18830), .ZN(
        P3_U3288) );
  INV_X1 U21879 ( .A(n18821), .ZN(n18824) );
  AOI222_X1 U21880 ( .A1(n18825), .A2(n18866), .B1(n18828), .B2(n18824), .C1(
        n18823), .C2(n18822), .ZN(n18826) );
  AOI22_X1 U21881 ( .A1(n18832), .A2(n18827), .B1(n18826), .B2(n18830), .ZN(
        P3_U3289) );
  AOI222_X1 U21882 ( .A1(n21021), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18866), 
        .B2(n18829), .C1(n21023), .C2(n18828), .ZN(n18831) );
  AOI22_X1 U21883 ( .A1(n18832), .A2(n21023), .B1(n18831), .B2(n18830), .ZN(
        P3_U3290) );
  NOR3_X1 U21884 ( .A1(n18834), .A2(P3_REIP_REG_0__SCAN_IN), .A3(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18833) );
  AOI221_X1 U21885 ( .B1(n18835), .B2(n18834), .C1(P3_REIP_REG_1__SCAN_IN), 
        .C2(P3_REIP_REG_0__SCAN_IN), .A(n18833), .ZN(n18837) );
  INV_X1 U21886 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18836) );
  INV_X1 U21887 ( .A(n18841), .ZN(n18838) );
  AOI22_X1 U21888 ( .A1(n18841), .A2(n18837), .B1(n18836), .B2(n18838), .ZN(
        P3_U3292) );
  NOR2_X1 U21889 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n18840) );
  INV_X1 U21890 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18839) );
  AOI22_X1 U21891 ( .A1(n18841), .A2(n18840), .B1(n18839), .B2(n18838), .ZN(
        P3_U3293) );
  INV_X1 U21892 ( .A(P3_READREQUEST_REG_SCAN_IN), .ZN(n18869) );
  OAI22_X1 U21893 ( .A1(n18863), .A2(n18869), .B1(P3_W_R_N_REG_SCAN_IN), .B2(
        n18842), .ZN(n18843) );
  INV_X1 U21894 ( .A(n18843), .ZN(P3_U3294) );
  NAND2_X1 U21895 ( .A1(n18846), .A2(P3_MORE_REG_SCAN_IN), .ZN(n18844) );
  OAI21_X1 U21896 ( .B1(n18846), .B2(n18845), .A(n18844), .ZN(P3_U3295) );
  OAI21_X1 U21897 ( .B1(n18849), .B2(n18848), .A(n18847), .ZN(n18850) );
  AOI21_X1 U21898 ( .B1(n17440), .B2(n18854), .A(n18850), .ZN(n18861) );
  AOI21_X1 U21899 ( .B1(n18853), .B2(n18852), .A(n18851), .ZN(n18855) );
  OAI211_X1 U21900 ( .C1(n18856), .C2(n18855), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18854), .ZN(n18858) );
  AOI21_X1 U21901 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18858), .A(n18857), 
        .ZN(n18860) );
  NAND2_X1 U21902 ( .A1(n18861), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18859) );
  OAI21_X1 U21903 ( .B1(n18861), .B2(n18860), .A(n18859), .ZN(P3_U3296) );
  OAI22_X1 U21904 ( .A1(n18863), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18862), .ZN(n18864) );
  INV_X1 U21905 ( .A(n18864), .ZN(P3_U3297) );
  AOI21_X1 U21906 ( .B1(n18866), .B2(n18865), .A(n18868), .ZN(n18872) );
  AOI22_X1 U21907 ( .A1(n18872), .A2(n18869), .B1(n18868), .B2(n18867), .ZN(
        P3_U3298) );
  INV_X1 U21908 ( .A(P3_MEMORYFETCH_REG_SCAN_IN), .ZN(n18871) );
  AOI21_X1 U21909 ( .B1(n18872), .B2(n18871), .A(n18870), .ZN(P3_U3299) );
  NAND2_X1 U21910 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19760), .ZN(n19749) );
  NAND2_X1 U21911 ( .A1(n19747), .A2(n19743), .ZN(n19748) );
  OAI21_X1 U21912 ( .B1(n19747), .B2(n19749), .A(n19748), .ZN(n19808) );
  AOI21_X1 U21913 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19808), .ZN(n18873) );
  INV_X1 U21914 ( .A(n18873), .ZN(P2_U2815) );
  NOR2_X1 U21915 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n18874), .ZN(n19736) );
  AOI22_X1 U21916 ( .A1(n18875), .A2(n19736), .B1(P2_CODEFETCH_REG_SCAN_IN), 
        .B2(n19863), .ZN(n18876) );
  INV_X1 U21917 ( .A(n18876), .ZN(P2_U2816) );
  INV_X1 U21918 ( .A(n18877), .ZN(n19880) );
  INV_X1 U21919 ( .A(n19754), .ZN(n18879) );
  AOI22_X1 U21920 ( .A1(P2_D_C_N_REG_SCAN_IN), .A2(n19880), .B1(n18879), .B2(
        n19747), .ZN(n18878) );
  OAI21_X1 U21921 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n19880), .A(n18878), 
        .ZN(P2_U2817) );
  OAI21_X1 U21922 ( .B1(n18879), .B2(BS16), .A(n19808), .ZN(n19806) );
  OAI21_X1 U21923 ( .B1(n19808), .B2(n19868), .A(n19806), .ZN(P2_U2818) );
  NOR2_X1 U21924 ( .A1(n18881), .A2(n18880), .ZN(n19859) );
  OAI21_X1 U21925 ( .B1(n19859), .B2(n18883), .A(n18882), .ZN(P2_U2819) );
  NOR4_X1 U21926 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_11__SCAN_IN), .A3(P2_DATAWIDTH_REG_12__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_13__SCAN_IN), .ZN(n18893) );
  NOR4_X1 U21927 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_7__SCAN_IN), .A3(P2_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_9__SCAN_IN), .ZN(n18892) );
  AOI211_X1 U21928 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_3__SCAN_IN), .B(
        P2_DATAWIDTH_REG_4__SCAN_IN), .ZN(n18884) );
  INV_X1 U21929 ( .A(P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n20925) );
  INV_X1 U21930 ( .A(P2_DATAWIDTH_REG_21__SCAN_IN), .ZN(n21026) );
  NAND3_X1 U21931 ( .A1(n18884), .A2(n20925), .A3(n21026), .ZN(n18890) );
  NOR4_X1 U21932 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_20__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18888) );
  NOR4_X1 U21933 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_16__SCAN_IN), .A3(P2_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n18887) );
  NOR4_X1 U21934 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18886) );
  NOR4_X1 U21935 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18885) );
  NAND4_X1 U21936 ( .A1(n18888), .A2(n18887), .A3(n18886), .A4(n18885), .ZN(
        n18889) );
  NOR4_X1 U21937 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_2__SCAN_IN), .A3(n18890), .A4(n18889), .ZN(n18891) );
  NAND3_X1 U21938 ( .A1(n18893), .A2(n18892), .A3(n18891), .ZN(n18902) );
  NOR2_X1 U21939 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18902), .ZN(n18896) );
  INV_X1 U21940 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18894) );
  AOI22_X1 U21941 ( .A1(n18896), .A2(n18897), .B1(n18902), .B2(n18894), .ZN(
        P2_U2820) );
  OR3_X1 U21942 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18901) );
  INV_X1 U21943 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18895) );
  AOI22_X1 U21944 ( .A1(n18896), .A2(n18901), .B1(n18902), .B2(n18895), .ZN(
        P2_U2821) );
  INV_X1 U21945 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19807) );
  NAND2_X1 U21946 ( .A1(n18896), .A2(n19807), .ZN(n18900) );
  INV_X1 U21947 ( .A(n18902), .ZN(n18904) );
  OAI21_X1 U21948 ( .B1(n18897), .B2(n14868), .A(n18904), .ZN(n18898) );
  OAI21_X1 U21949 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18904), .A(n18898), 
        .ZN(n18899) );
  OAI221_X1 U21950 ( .B1(n18900), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18900), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18899), .ZN(P2_U2822) );
  INV_X1 U21951 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18903) );
  OAI221_X1 U21952 ( .B1(n18904), .B2(n18903), .C1(n18902), .C2(n18901), .A(
        n18900), .ZN(P2_U2823) );
  OAI22_X1 U21953 ( .A1(n18905), .A2(n19014), .B1(n10877), .B2(n18999), .ZN(
        n18906) );
  AOI211_X1 U21954 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n18957), .A(n19206), .B(
        n18906), .ZN(n18917) );
  NAND2_X1 U21955 ( .A1(n19019), .A2(n18907), .ZN(n18908) );
  XNOR2_X1 U21956 ( .A(n18909), .B(n18908), .ZN(n18914) );
  INV_X1 U21957 ( .A(n18910), .ZN(n18911) );
  OAI22_X1 U21958 ( .A1(n18912), .A2(n19037), .B1(n18911), .B2(n19026), .ZN(
        n18913) );
  AOI21_X1 U21959 ( .B1(n18915), .B2(n18914), .A(n18913), .ZN(n18916) );
  OAI211_X1 U21960 ( .C1(n18918), .C2(n19041), .A(n18917), .B(n18916), .ZN(
        P2_U2836) );
  AOI22_X1 U21961 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19003), .B1(
        P2_REIP_REG_17__SCAN_IN), .B2(n19028), .ZN(n18919) );
  OAI21_X1 U21962 ( .B1(n18920), .B2(n19014), .A(n18919), .ZN(n18921) );
  AOI211_X1 U21963 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n18957), .A(n19206), .B(
        n18921), .ZN(n18929) );
  NAND2_X1 U21964 ( .A1(n19019), .A2(n18922), .ZN(n18923) );
  XOR2_X1 U21965 ( .A(n18924), .B(n18923), .Z(n18927) );
  INV_X1 U21966 ( .A(n18925), .ZN(n18926) );
  AOI22_X1 U21967 ( .A1(n18927), .A2(n18915), .B1(n18926), .B2(n10916), .ZN(
        n18928) );
  OAI211_X1 U21968 ( .C1(n18930), .C2(n19026), .A(n18929), .B(n18928), .ZN(
        P2_U2838) );
  NOR2_X1 U21969 ( .A1(n19005), .A2(n18931), .ZN(n18933) );
  XOR2_X1 U21970 ( .A(n18933), .B(n18932), .Z(n18942) );
  AOI22_X1 U21971 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n19003), .B1(
        P2_REIP_REG_16__SCAN_IN), .B2(n19028), .ZN(n18934) );
  OAI21_X1 U21972 ( .B1(n18935), .B2(n19014), .A(n18934), .ZN(n18936) );
  AOI211_X1 U21973 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n18957), .A(n19206), .B(
        n18936), .ZN(n18941) );
  OAI22_X1 U21974 ( .A1(n18938), .A2(n19037), .B1(n18937), .B2(n19026), .ZN(
        n18939) );
  INV_X1 U21975 ( .A(n18939), .ZN(n18940) );
  OAI211_X1 U21976 ( .C1(n19738), .C2(n18942), .A(n18941), .B(n18940), .ZN(
        P2_U2839) );
  NOR2_X1 U21977 ( .A1(n19005), .A2(n18943), .ZN(n18945) );
  XOR2_X1 U21978 ( .A(n18945), .B(n18944), .Z(n18953) );
  AOI22_X1 U21979 ( .A1(n18946), .A2(n19035), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19003), .ZN(n18947) );
  OAI211_X1 U21980 ( .C1(n12106), .C2(n19031), .A(n18947), .B(n19012), .ZN(
        n18948) );
  AOI21_X1 U21981 ( .B1(P2_REIP_REG_14__SCAN_IN), .B2(n19028), .A(n18948), 
        .ZN(n18952) );
  OAI22_X1 U21982 ( .A1(n18949), .A2(n19037), .B1(n19055), .B2(n19026), .ZN(
        n18950) );
  INV_X1 U21983 ( .A(n18950), .ZN(n18951) );
  OAI211_X1 U21984 ( .C1(n19738), .C2(n18953), .A(n18952), .B(n18951), .ZN(
        P2_U2841) );
  AOI22_X1 U21985 ( .A1(n18954), .A2(n19035), .B1(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n19003), .ZN(n18955) );
  OAI21_X1 U21986 ( .B1(n15187), .B2(n18999), .A(n18955), .ZN(n18956) );
  AOI211_X1 U21987 ( .C1(P2_EBX_REG_13__SCAN_IN), .C2(n18957), .A(n19206), .B(
        n18956), .ZN(n18964) );
  NAND2_X1 U21988 ( .A1(n19019), .A2(n18958), .ZN(n18960) );
  XNOR2_X1 U21989 ( .A(n18960), .B(n18959), .ZN(n18962) );
  AOI22_X1 U21990 ( .A1(n18962), .A2(n18915), .B1(n18961), .B2(n10916), .ZN(
        n18963) );
  OAI211_X1 U21991 ( .C1(n19057), .C2(n19026), .A(n18964), .B(n18963), .ZN(
        P2_U2842) );
  NOR2_X1 U21992 ( .A1(n19005), .A2(n18965), .ZN(n18966) );
  XOR2_X1 U21993 ( .A(n18967), .B(n18966), .Z(n18975) );
  AOI22_X1 U21994 ( .A1(n18968), .A2(n19035), .B1(P2_REIP_REG_12__SCAN_IN), 
        .B2(n19028), .ZN(n18969) );
  OAI211_X1 U21995 ( .C1(n20941), .C2(n19031), .A(n18969), .B(n19012), .ZN(
        n18973) );
  INV_X1 U21996 ( .A(n18970), .ZN(n18971) );
  OAI22_X1 U21997 ( .A1(n18971), .A2(n19037), .B1(n19026), .B2(n19059), .ZN(
        n18972) );
  AOI211_X1 U21998 ( .C1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(n19003), .A(
        n18973), .B(n18972), .ZN(n18974) );
  OAI21_X1 U21999 ( .B1(n19738), .B2(n18975), .A(n18974), .ZN(P2_U2843) );
  NAND2_X1 U22000 ( .A1(n19019), .A2(n18976), .ZN(n18978) );
  XOR2_X1 U22001 ( .A(n18978), .B(n18977), .Z(n18986) );
  INV_X1 U22002 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n18981) );
  AOI22_X1 U22003 ( .A1(n18979), .A2(n19035), .B1(P2_REIP_REG_9__SCAN_IN), 
        .B2(n19028), .ZN(n18980) );
  OAI211_X1 U22004 ( .C1(n18981), .C2(n19031), .A(n18980), .B(n19012), .ZN(
        n18984) );
  OAI22_X1 U22005 ( .A1(n18982), .A2(n19037), .B1(n19066), .B2(n19026), .ZN(
        n18983) );
  AOI211_X1 U22006 ( .C1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n19003), .A(
        n18984), .B(n18983), .ZN(n18985) );
  OAI21_X1 U22007 ( .B1(n18986), .B2(n19738), .A(n18985), .ZN(P2_U2846) );
  NAND2_X1 U22008 ( .A1(n19019), .A2(n18987), .ZN(n18989) );
  XOR2_X1 U22009 ( .A(n18989), .B(n18988), .Z(n18997) );
  AOI22_X1 U22010 ( .A1(n18990), .A2(n19035), .B1(P2_REIP_REG_7__SCAN_IN), 
        .B2(n19028), .ZN(n18991) );
  OAI211_X1 U22011 ( .C1(n18992), .C2(n19031), .A(n18991), .B(n19012), .ZN(
        n18995) );
  OAI22_X1 U22012 ( .A1(n18993), .A2(n19037), .B1(n19071), .B2(n19026), .ZN(
        n18994) );
  AOI211_X1 U22013 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n19003), .A(
        n18995), .B(n18994), .ZN(n18996) );
  OAI21_X1 U22014 ( .B1(n18997), .B2(n19738), .A(n18996), .ZN(P2_U2848) );
  OAI21_X1 U22015 ( .B1(n18998), .B2(n19031), .A(n19012), .ZN(n19002) );
  OAI22_X1 U22016 ( .A1(n19000), .A2(n19014), .B1(n19765), .B2(n18999), .ZN(
        n19001) );
  AOI211_X1 U22017 ( .C1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n19003), .A(
        n19002), .B(n19001), .ZN(n19011) );
  NOR2_X1 U22018 ( .A1(n19005), .A2(n19004), .ZN(n19007) );
  XNOR2_X1 U22019 ( .A(n19007), .B(n19006), .ZN(n19009) );
  AOI22_X1 U22020 ( .A1(n19009), .A2(n18915), .B1(n10916), .B2(n19008), .ZN(
        n19010) );
  OAI211_X1 U22021 ( .C1(n19026), .C2(n19073), .A(n19011), .B(n19010), .ZN(
        P2_U2849) );
  OAI21_X1 U22022 ( .B1(n19013), .B2(n19031), .A(n19012), .ZN(n19017) );
  OAI22_X1 U22023 ( .A1(n19015), .A2(n19014), .B1(n19041), .B2(n20749), .ZN(
        n19016) );
  AOI211_X1 U22024 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19028), .A(n19017), .B(
        n19016), .ZN(n19025) );
  NAND2_X1 U22025 ( .A1(n19019), .A2(n19018), .ZN(n19020) );
  XNOR2_X1 U22026 ( .A(n19021), .B(n19020), .ZN(n19023) );
  AOI22_X1 U22027 ( .A1(n19023), .A2(n18915), .B1(n10916), .B2(n19022), .ZN(
        n19024) );
  OAI211_X1 U22028 ( .C1(n19026), .C2(n19085), .A(n19025), .B(n19024), .ZN(
        P2_U2850) );
  INV_X1 U22029 ( .A(n19027), .ZN(n19034) );
  AOI22_X1 U22030 ( .A1(n19029), .A2(n19109), .B1(n19028), .B2(
        P2_REIP_REG_0__SCAN_IN), .ZN(n19030) );
  OAI21_X1 U22031 ( .B1(n19032), .B2(n19031), .A(n19030), .ZN(n19033) );
  AOI21_X1 U22032 ( .B1(n19035), .B2(n19034), .A(n19033), .ZN(n19036) );
  OAI21_X1 U22033 ( .B1(n19038), .B2(n19037), .A(n19036), .ZN(n19043) );
  AOI21_X1 U22034 ( .B1(n19041), .B2(n19040), .A(n19039), .ZN(n19042) );
  AOI211_X1 U22035 ( .C1(n19110), .C2(n19044), .A(n19043), .B(n19042), .ZN(
        n19045) );
  OAI21_X1 U22036 ( .B1(n19738), .B2(n19046), .A(n19045), .ZN(P2_U2855) );
  AOI22_X1 U22037 ( .A1(n19048), .A2(n19106), .B1(n19047), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19051) );
  AOI22_X1 U22038 ( .A1(P2_EAX_REG_31__SCAN_IN), .A2(n19105), .B1(n19049), 
        .B2(BUF1_REG_31__SCAN_IN), .ZN(n19050) );
  NAND2_X1 U22039 ( .A1(n19051), .A2(n19050), .ZN(P2_U2888) );
  OAI222_X1 U22040 ( .A1(n19053), .A2(n19086), .B1(n13148), .B2(n19072), .C1(
        n19052), .C2(n19113), .ZN(P2_U2904) );
  AOI22_X1 U22041 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19105), .B1(n19184), 
        .B2(n19074), .ZN(n19054) );
  OAI21_X1 U22042 ( .B1(n19086), .B2(n19055), .A(n19054), .ZN(P2_U2905) );
  INV_X1 U22043 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19155) );
  OAI222_X1 U22044 ( .A1(n19057), .A2(n19086), .B1(n19155), .B2(n19072), .C1(
        n19113), .C2(n19056), .ZN(P2_U2906) );
  INV_X1 U22045 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19157) );
  OAI222_X1 U22046 ( .A1(n19059), .A2(n19086), .B1(n19157), .B2(n19072), .C1(
        n19113), .C2(n19058), .ZN(P2_U2907) );
  INV_X1 U22047 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19159) );
  OAI222_X1 U22048 ( .A1(n19061), .A2(n19086), .B1(n19159), .B2(n19072), .C1(
        n19113), .C2(n19060), .ZN(P2_U2908) );
  INV_X1 U22049 ( .A(n19062), .ZN(n19064) );
  INV_X1 U22050 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n19161) );
  OAI222_X1 U22051 ( .A1(n19064), .A2(n19086), .B1(n19161), .B2(n19072), .C1(
        n19113), .C2(n19063), .ZN(P2_U2909) );
  INV_X1 U22052 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19163) );
  OAI222_X1 U22053 ( .A1(n19066), .A2(n19086), .B1(n19163), .B2(n19072), .C1(
        n19113), .C2(n19065), .ZN(P2_U2910) );
  INV_X1 U22054 ( .A(n19067), .ZN(n19070) );
  AOI22_X1 U22055 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19105), .B1(n19068), .B2(
        n19074), .ZN(n19069) );
  OAI21_X1 U22056 ( .B1(n19086), .B2(n19070), .A(n19069), .ZN(P2_U2911) );
  INV_X1 U22057 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19167) );
  OAI222_X1 U22058 ( .A1(n19071), .A2(n19086), .B1(n19167), .B2(n19072), .C1(
        n19113), .C2(n19256), .ZN(P2_U2912) );
  INV_X1 U22059 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19169) );
  OAI222_X1 U22060 ( .A1(n19073), .A2(n19086), .B1(n19169), .B2(n19072), .C1(
        n19113), .C2(n19246), .ZN(P2_U2913) );
  AOI22_X1 U22061 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19105), .B1(n19075), .B2(
        n19074), .ZN(n19084) );
  NAND2_X1 U22062 ( .A1(n19818), .A2(n19096), .ZN(n19081) );
  XOR2_X1 U22063 ( .A(n19096), .B(n19818), .Z(n19094) );
  NAND2_X1 U22064 ( .A1(n19825), .A2(n19076), .ZN(n19080) );
  XNOR2_X1 U22065 ( .A(n19825), .B(n19829), .ZN(n19101) );
  INV_X1 U22066 ( .A(n19833), .ZN(n19077) );
  NAND2_X1 U22067 ( .A1(n19838), .A2(n19077), .ZN(n19079) );
  NAND2_X1 U22068 ( .A1(n19079), .A2(n19078), .ZN(n19100) );
  NAND2_X1 U22069 ( .A1(n19101), .A2(n19100), .ZN(n19099) );
  NAND2_X1 U22070 ( .A1(n19080), .A2(n19099), .ZN(n19093) );
  NAND2_X1 U22071 ( .A1(n19094), .A2(n19093), .ZN(n19092) );
  AOI21_X1 U22072 ( .B1(n19081), .B2(n19092), .A(n19207), .ZN(n19087) );
  OR3_X1 U22073 ( .A1(n19088), .A2(n19087), .A3(n19082), .ZN(n19083) );
  OAI211_X1 U22074 ( .C1(n19086), .C2(n19085), .A(n19084), .B(n19083), .ZN(
        P2_U2914) );
  AOI22_X1 U22075 ( .A1(n19106), .A2(n19207), .B1(n19105), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n19091) );
  XOR2_X1 U22076 ( .A(n19088), .B(n19087), .Z(n19089) );
  NAND2_X1 U22077 ( .A1(n19089), .A2(n19107), .ZN(n19090) );
  OAI211_X1 U22078 ( .C1(n19234), .C2(n19113), .A(n19091), .B(n19090), .ZN(
        P2_U2915) );
  OAI21_X1 U22079 ( .B1(n19094), .B2(n19093), .A(n19092), .ZN(n19095) );
  NAND2_X1 U22080 ( .A1(n19095), .A2(n19107), .ZN(n19098) );
  INV_X1 U22081 ( .A(n19096), .ZN(n19821) );
  AOI22_X1 U22082 ( .A1(n19821), .A2(n19106), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19105), .ZN(n19097) );
  OAI211_X1 U22083 ( .C1(n19229), .C2(n19113), .A(n19098), .B(n19097), .ZN(
        P2_U2916) );
  AOI22_X1 U22084 ( .A1(n19829), .A2(n19106), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19105), .ZN(n19104) );
  OAI21_X1 U22085 ( .B1(n19101), .B2(n19100), .A(n19099), .ZN(n19102) );
  NAND2_X1 U22086 ( .A1(n19102), .A2(n19107), .ZN(n19103) );
  OAI211_X1 U22087 ( .C1(n19224), .C2(n19113), .A(n19104), .B(n19103), .ZN(
        P2_U2917) );
  AOI22_X1 U22088 ( .A1(n19106), .A2(n19109), .B1(n19105), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n19112) );
  OAI211_X1 U22089 ( .C1(n19110), .C2(n19109), .A(n19108), .B(n19107), .ZN(
        n19111) );
  OAI211_X1 U22090 ( .C1(n19114), .C2(n19113), .A(n19112), .B(n19111), .ZN(
        P2_U2919) );
  INV_X1 U22091 ( .A(n19115), .ZN(n19117) );
  OAI21_X1 U22092 ( .B1(n19118), .B2(n19117), .A(n19116), .ZN(n19119) );
  OR2_X1 U22093 ( .A1(n19843), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19864) );
  NOR2_X1 U22094 ( .A1(n19173), .A2(n19120), .ZN(P2_U2920) );
  INV_X1 U22095 ( .A(n19149), .ZN(n19124) );
  AOI22_X1 U22096 ( .A1(P2_EAX_REG_30__SCAN_IN), .A2(n19124), .B1(n9727), .B2(
        P2_UWORD_REG_14__SCAN_IN), .ZN(n19122) );
  OAI21_X1 U22097 ( .B1(n19173), .B2(n19123), .A(n19122), .ZN(P2_U2921) );
  AOI22_X1 U22098 ( .A1(P2_EAX_REG_29__SCAN_IN), .A2(n19124), .B1(n9727), .B2(
        P2_UWORD_REG_13__SCAN_IN), .ZN(n19125) );
  OAI21_X1 U22099 ( .B1(n20773), .B2(n19173), .A(n19125), .ZN(P2_U2922) );
  AOI22_X1 U22100 ( .A1(n9727), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n19126) );
  OAI21_X1 U22101 ( .B1(n19127), .B2(n19149), .A(n19126), .ZN(P2_U2923) );
  AOI22_X1 U22102 ( .A1(n9727), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n19128) );
  OAI21_X1 U22103 ( .B1(n19129), .B2(n19149), .A(n19128), .ZN(P2_U2924) );
  AOI22_X1 U22104 ( .A1(n9727), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n19130) );
  OAI21_X1 U22105 ( .B1(n19131), .B2(n19149), .A(n19130), .ZN(P2_U2925) );
  INV_X1 U22106 ( .A(P2_UWORD_REG_9__SCAN_IN), .ZN(n20826) );
  OAI222_X1 U22107 ( .A1(n19173), .A2(n20850), .B1(n19149), .B2(n20748), .C1(
        n19864), .C2(n20826), .ZN(P2_U2926) );
  AOI22_X1 U22108 ( .A1(n9727), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n19132) );
  OAI21_X1 U22109 ( .B1(n19133), .B2(n19149), .A(n19132), .ZN(P2_U2927) );
  AOI22_X1 U22110 ( .A1(n9727), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n19134) );
  OAI21_X1 U22111 ( .B1(n19135), .B2(n19149), .A(n19134), .ZN(P2_U2928) );
  AOI22_X1 U22112 ( .A1(n9727), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n19136) );
  OAI21_X1 U22113 ( .B1(n19137), .B2(n19149), .A(n19136), .ZN(P2_U2929) );
  INV_X1 U22114 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n19139) );
  AOI22_X1 U22115 ( .A1(n9727), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n19138) );
  OAI21_X1 U22116 ( .B1(n19139), .B2(n19149), .A(n19138), .ZN(P2_U2930) );
  AOI22_X1 U22117 ( .A1(n9727), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n19140) );
  OAI21_X1 U22118 ( .B1(n19141), .B2(n19149), .A(n19140), .ZN(P2_U2931) );
  AOI22_X1 U22119 ( .A1(n9727), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n19142) );
  OAI21_X1 U22120 ( .B1(n19143), .B2(n19149), .A(n19142), .ZN(P2_U2932) );
  AOI22_X1 U22121 ( .A1(n9727), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n19144) );
  OAI21_X1 U22122 ( .B1(n19145), .B2(n19149), .A(n19144), .ZN(P2_U2933) );
  AOI22_X1 U22123 ( .A1(n9727), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n19146) );
  OAI21_X1 U22124 ( .B1(n19147), .B2(n19149), .A(n19146), .ZN(P2_U2934) );
  AOI22_X1 U22125 ( .A1(n9727), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n19148) );
  OAI21_X1 U22126 ( .B1(n19150), .B2(n19149), .A(n19148), .ZN(P2_U2935) );
  AOI22_X1 U22127 ( .A1(n9727), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19151) );
  OAI21_X1 U22128 ( .B1(n13148), .B2(n19182), .A(n19151), .ZN(P2_U2936) );
  INV_X1 U22129 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19153) );
  AOI22_X1 U22130 ( .A1(n9727), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19152) );
  OAI21_X1 U22131 ( .B1(n19153), .B2(n19182), .A(n19152), .ZN(P2_U2937) );
  AOI22_X1 U22132 ( .A1(n9727), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19154) );
  OAI21_X1 U22133 ( .B1(n19155), .B2(n19182), .A(n19154), .ZN(P2_U2938) );
  AOI22_X1 U22134 ( .A1(n9727), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19156) );
  OAI21_X1 U22135 ( .B1(n19157), .B2(n19182), .A(n19156), .ZN(P2_U2939) );
  AOI22_X1 U22136 ( .A1(n9727), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19158) );
  OAI21_X1 U22137 ( .B1(n19159), .B2(n19182), .A(n19158), .ZN(P2_U2940) );
  INV_X1 U22138 ( .A(P2_LWORD_REG_10__SCAN_IN), .ZN(n20787) );
  OAI222_X1 U22139 ( .A1(n19864), .A2(n20787), .B1(n19182), .B2(n19161), .C1(
        n19173), .C2(n19160), .ZN(P2_U2941) );
  INV_X1 U22140 ( .A(P2_LWORD_REG_9__SCAN_IN), .ZN(n20759) );
  OAI222_X1 U22141 ( .A1(n19864), .A2(n20759), .B1(n19182), .B2(n19163), .C1(
        n19173), .C2(n19162), .ZN(P2_U2942) );
  AOI22_X1 U22142 ( .A1(n9727), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19164) );
  OAI21_X1 U22143 ( .B1(n19165), .B2(n19182), .A(n19164), .ZN(P2_U2943) );
  AOI22_X1 U22144 ( .A1(n9727), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19166) );
  OAI21_X1 U22145 ( .B1(n19167), .B2(n19182), .A(n19166), .ZN(P2_U2944) );
  AOI22_X1 U22146 ( .A1(n9727), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19168) );
  OAI21_X1 U22147 ( .B1(n19169), .B2(n19182), .A(n19168), .ZN(P2_U2945) );
  INV_X1 U22148 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19171) );
  AOI22_X1 U22149 ( .A1(n9727), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19170) );
  OAI21_X1 U22150 ( .B1(n19171), .B2(n19182), .A(n19170), .ZN(P2_U2946) );
  INV_X1 U22151 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n20939) );
  INV_X1 U22152 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n20870) );
  OAI222_X1 U22153 ( .A1(n19864), .A2(n20939), .B1(n19182), .B2(n20870), .C1(
        n19173), .C2(n19172), .ZN(P2_U2947) );
  INV_X1 U22154 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19175) );
  AOI22_X1 U22155 ( .A1(n9727), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19174) );
  OAI21_X1 U22156 ( .B1(n19175), .B2(n19182), .A(n19174), .ZN(P2_U2948) );
  INV_X1 U22157 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19177) );
  AOI22_X1 U22158 ( .A1(n9727), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19176) );
  OAI21_X1 U22159 ( .B1(n19177), .B2(n19182), .A(n19176), .ZN(P2_U2949) );
  INV_X1 U22160 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19179) );
  AOI22_X1 U22161 ( .A1(n9727), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19178) );
  OAI21_X1 U22162 ( .B1(n19179), .B2(n19182), .A(n19178), .ZN(P2_U2950) );
  INV_X1 U22163 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n19183) );
  AOI22_X1 U22164 ( .A1(n9727), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19180), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19181) );
  OAI21_X1 U22165 ( .B1(n19183), .B2(n19182), .A(n19181), .ZN(P2_U2951) );
  AOI22_X1 U22166 ( .A1(P2_EAX_REG_30__SCAN_IN), .A2(n13178), .B1(n19187), 
        .B2(P2_UWORD_REG_14__SCAN_IN), .ZN(n19186) );
  NAND2_X1 U22167 ( .A1(n19185), .A2(n19184), .ZN(n19188) );
  NAND2_X1 U22168 ( .A1(n19186), .A2(n19188), .ZN(P2_U2966) );
  AOI22_X1 U22169 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n13178), .B1(n19187), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n19189) );
  NAND2_X1 U22170 ( .A1(n19189), .A2(n19188), .ZN(P2_U2981) );
  AOI22_X1 U22171 ( .A1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n19190), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19206), .ZN(n19203) );
  XOR2_X1 U22172 ( .A(n19191), .B(n19192), .Z(n19218) );
  INV_X1 U22173 ( .A(n19218), .ZN(n19199) );
  INV_X1 U22174 ( .A(n19193), .ZN(n19196) );
  INV_X1 U22175 ( .A(n19194), .ZN(n19195) );
  AOI21_X1 U22176 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n19196), .A(
        n19195), .ZN(n19216) );
  OAI22_X1 U22177 ( .A1(n19199), .A2(n19198), .B1(n19216), .B2(n19197), .ZN(
        n19200) );
  AOI21_X1 U22178 ( .B1(n19201), .B2(n19213), .A(n19200), .ZN(n19202) );
  OAI211_X1 U22179 ( .C1(n19205), .C2(n19204), .A(n19203), .B(n19202), .ZN(
        P2_U3010) );
  AOI22_X1 U22180 ( .A1(n19208), .A2(n19207), .B1(n19206), .B2(
        P2_REIP_REG_4__SCAN_IN), .ZN(n19221) );
  NOR2_X1 U22181 ( .A1(n19210), .A2(n19209), .ZN(n19211) );
  AOI21_X1 U22182 ( .B1(n19213), .B2(n19212), .A(n19211), .ZN(n19214) );
  OAI21_X1 U22183 ( .B1(n19216), .B2(n19215), .A(n19214), .ZN(n19217) );
  AOI21_X1 U22184 ( .B1(n19219), .B2(n19218), .A(n19217), .ZN(n19220) );
  OAI211_X1 U22185 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n19222), .A(
        n19221), .B(n19220), .ZN(P2_U3042) );
  AOI22_X1 U22186 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19252), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19251), .ZN(n19528) );
  AOI22_X1 U22187 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n19251), .B1(
        BUF1_REG_26__SCAN_IN), .B2(n19252), .ZN(n19697) );
  NOR2_X2 U22188 ( .A1(n19223), .A2(n19253), .ZN(n19692) );
  AOI22_X1 U22189 ( .A1(n19581), .A2(n19728), .B1(n19255), .B2(n19692), .ZN(
        n19226) );
  NOR2_X2 U22190 ( .A1(n19224), .A2(n19436), .ZN(n19693) );
  AOI22_X1 U22191 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19258), .B1(
        n19693), .B2(n19257), .ZN(n19225) );
  OAI211_X1 U22192 ( .C1(n19528), .C2(n19289), .A(n19226), .B(n19225), .ZN(
        P2_U3050) );
  AOI22_X1 U22193 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19252), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19251), .ZN(n19656) );
  INV_X1 U22194 ( .A(n19251), .ZN(n19243) );
  NOR2_X2 U22195 ( .A1(n19228), .A2(n19253), .ZN(n19698) );
  AOI22_X1 U22196 ( .A1(n19653), .A2(n19728), .B1(n19255), .B2(n19698), .ZN(
        n19231) );
  NOR2_X2 U22197 ( .A1(n19229), .A2(n19436), .ZN(n19699) );
  AOI22_X1 U22198 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19258), .B1(
        n19699), .B2(n19257), .ZN(n19230) );
  OAI211_X1 U22199 ( .C1(n19656), .C2(n19289), .A(n19231), .B(n19230), .ZN(
        P2_U3051) );
  AOI22_X2 U22200 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19252), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19251), .ZN(n19709) );
  OAI22_X2 U22201 ( .A1(n19233), .A2(n19242), .B1(n19232), .B2(n19243), .ZN(
        n19706) );
  NOR2_X2 U22202 ( .A1(n10742), .A2(n19253), .ZN(n19704) );
  AOI22_X1 U22203 ( .A1(n19706), .A2(n19728), .B1(n19255), .B2(n19704), .ZN(
        n19236) );
  NOR2_X2 U22204 ( .A1(n19234), .A2(n19436), .ZN(n19705) );
  AOI22_X1 U22205 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19258), .B1(
        n19705), .B2(n19257), .ZN(n19235) );
  OAI211_X1 U22206 ( .C1(n19709), .C2(n19289), .A(n19236), .B(n19235), .ZN(
        P2_U3052) );
  AOI22_X1 U22207 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n19252), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n19251), .ZN(n19714) );
  AOI22_X1 U22208 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n19252), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n19251), .ZN(n19567) );
  AOI22_X1 U22209 ( .A1(n19711), .A2(n19728), .B1(n19255), .B2(n19238), .ZN(
        n19241) );
  NOR2_X2 U22210 ( .A1(n19239), .A2(n19436), .ZN(n19710) );
  AOI22_X1 U22211 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19258), .B1(
        n19710), .B2(n19257), .ZN(n19240) );
  OAI211_X1 U22212 ( .C1(n19714), .C2(n19289), .A(n19241), .B(n19240), .ZN(
        P2_U3053) );
  INV_X1 U22213 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n20790) );
  NOR2_X2 U22214 ( .A1(n19245), .A2(n19253), .ZN(n19715) );
  AOI22_X1 U22215 ( .A1(n19717), .A2(n19728), .B1(n19255), .B2(n19715), .ZN(
        n19248) );
  NOR2_X2 U22216 ( .A1(n19246), .A2(n19436), .ZN(n19716) );
  AOI22_X1 U22217 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n19252), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n19251), .ZN(n19722) );
  INV_X1 U22218 ( .A(n19722), .ZN(n19568) );
  AOI22_X1 U22219 ( .A1(n19716), .A2(n19257), .B1(n19281), .B2(n19568), .ZN(
        n19247) );
  OAI211_X1 U22220 ( .C1(n19250), .C2(n19249), .A(n19248), .B(n19247), .ZN(
        P2_U3054) );
  AOI22_X1 U22221 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19252), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19251), .ZN(n19670) );
  AOI22_X1 U22222 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19252), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19251), .ZN(n19733) );
  INV_X1 U22223 ( .A(n19733), .ZN(n19665) );
  NOR2_X2 U22224 ( .A1(n19254), .A2(n19253), .ZN(n19723) );
  AOI22_X1 U22225 ( .A1(n19665), .A2(n19728), .B1(n19255), .B2(n19723), .ZN(
        n19260) );
  NOR2_X2 U22226 ( .A1(n19256), .A2(n19436), .ZN(n19725) );
  AOI22_X1 U22227 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19258), .B1(
        n19725), .B2(n19257), .ZN(n19259) );
  OAI211_X1 U22228 ( .C1(n19670), .C2(n19289), .A(n19260), .B(n19259), .ZN(
        P2_U3055) );
  NOR2_X1 U22229 ( .A1(n19261), .A2(n19324), .ZN(n19284) );
  NOR3_X1 U22230 ( .A1(n19262), .A2(n19284), .A3(n10692), .ZN(n19263) );
  AOI211_X2 U22231 ( .C1(n19265), .C2(n10692), .A(n19734), .B(n19263), .ZN(
        n19285) );
  AOI22_X1 U22232 ( .A1(n19285), .A2(n19674), .B1(n19673), .B2(n19284), .ZN(
        n19269) );
  INV_X1 U22233 ( .A(n19284), .ZN(n19264) );
  AOI211_X1 U22234 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19264), .A(n19436), 
        .B(n19263), .ZN(n19267) );
  NAND2_X1 U22235 ( .A1(n19818), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19435) );
  OAI21_X1 U22236 ( .B1(n19435), .B2(n19491), .A(n19265), .ZN(n19266) );
  NAND2_X1 U22237 ( .A1(n19267), .A2(n19266), .ZN(n19286) );
  AOI22_X1 U22238 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19286), .B1(
        n19281), .B2(n19632), .ZN(n19268) );
  OAI211_X1 U22239 ( .C1(n19645), .C2(n19316), .A(n19269), .B(n19268), .ZN(
        P2_U3056) );
  AOI22_X1 U22240 ( .A1(n19285), .A2(n19687), .B1(n19686), .B2(n19284), .ZN(
        n19272) );
  AOI22_X1 U22241 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19286), .B1(
        n19281), .B2(n19646), .ZN(n19271) );
  OAI211_X1 U22242 ( .C1(n19649), .C2(n19316), .A(n19272), .B(n19271), .ZN(
        P2_U3057) );
  AOI22_X1 U22243 ( .A1(n19285), .A2(n19693), .B1(n19692), .B2(n19284), .ZN(
        n19274) );
  INV_X1 U22244 ( .A(n19528), .ZN(n19694) );
  AOI22_X1 U22245 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19286), .B1(
        n19319), .B2(n19694), .ZN(n19273) );
  OAI211_X1 U22246 ( .C1(n19697), .C2(n19289), .A(n19274), .B(n19273), .ZN(
        P2_U3058) );
  AOI22_X1 U22247 ( .A1(n19285), .A2(n19699), .B1(n19698), .B2(n19284), .ZN(
        n19276) );
  INV_X1 U22248 ( .A(n19656), .ZN(n19700) );
  AOI22_X1 U22249 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19286), .B1(
        n19319), .B2(n19700), .ZN(n19275) );
  OAI211_X1 U22250 ( .C1(n19703), .C2(n19289), .A(n19276), .B(n19275), .ZN(
        P2_U3059) );
  AOI22_X1 U22251 ( .A1(n19285), .A2(n19705), .B1(n19704), .B2(n19284), .ZN(
        n19278) );
  AOI22_X1 U22252 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19286), .B1(
        n19281), .B2(n19706), .ZN(n19277) );
  OAI211_X1 U22253 ( .C1(n19709), .C2(n19316), .A(n19278), .B(n19277), .ZN(
        P2_U3060) );
  AOI22_X1 U22254 ( .A1(n19285), .A2(n19710), .B1(n19238), .B2(n19284), .ZN(
        n19280) );
  INV_X1 U22255 ( .A(n19714), .ZN(n19564) );
  AOI22_X1 U22256 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19286), .B1(
        n19319), .B2(n19564), .ZN(n19279) );
  OAI211_X1 U22257 ( .C1(n19567), .C2(n19289), .A(n19280), .B(n19279), .ZN(
        P2_U3061) );
  AOI22_X1 U22258 ( .A1(n19285), .A2(n19716), .B1(n19715), .B2(n19284), .ZN(
        n19283) );
  AOI22_X1 U22259 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19286), .B1(
        n19281), .B2(n19717), .ZN(n19282) );
  OAI211_X1 U22260 ( .C1(n19722), .C2(n19316), .A(n19283), .B(n19282), .ZN(
        P2_U3062) );
  AOI22_X1 U22261 ( .A1(n19285), .A2(n19725), .B1(n19723), .B2(n19284), .ZN(
        n19288) );
  INV_X1 U22262 ( .A(n19670), .ZN(n19727) );
  AOI22_X1 U22263 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19286), .B1(
        n19319), .B2(n19727), .ZN(n19287) );
  OAI211_X1 U22264 ( .C1(n19733), .C2(n19289), .A(n19288), .B(n19287), .ZN(
        P2_U3063) );
  NOR2_X1 U22265 ( .A1(n19290), .A2(n19324), .ZN(n19317) );
  OAI21_X1 U22266 ( .B1(n12002), .B2(n19317), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19293) );
  INV_X1 U22267 ( .A(n19324), .ZN(n19291) );
  NAND2_X1 U22268 ( .A1(n19292), .A2(n19291), .ZN(n19297) );
  NAND2_X1 U22269 ( .A1(n19293), .A2(n19297), .ZN(n19318) );
  AOI22_X1 U22270 ( .A1(n19318), .A2(n19674), .B1(n19673), .B2(n19317), .ZN(
        n19303) );
  INV_X1 U22271 ( .A(n19317), .ZN(n19294) );
  OAI21_X1 U22272 ( .B1(n19295), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19294), 
        .ZN(n19300) );
  OAI21_X1 U22273 ( .B1(n19348), .B2(n19319), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19298) );
  NAND2_X1 U22274 ( .A1(n19298), .A2(n19297), .ZN(n19299) );
  MUX2_X1 U22275 ( .A(n19300), .B(n19299), .S(n19820), .Z(n19301) );
  NAND2_X1 U22276 ( .A1(n19301), .A2(n19680), .ZN(n19320) );
  AOI22_X1 U22277 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19320), .B1(
        n19348), .B2(n19682), .ZN(n19302) );
  OAI211_X1 U22278 ( .C1(n19685), .C2(n19316), .A(n19303), .B(n19302), .ZN(
        P2_U3064) );
  AOI22_X1 U22279 ( .A1(n19318), .A2(n19687), .B1(n19686), .B2(n19317), .ZN(
        n19305) );
  AOI22_X1 U22280 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19320), .B1(
        n19319), .B2(n19646), .ZN(n19304) );
  OAI211_X1 U22281 ( .C1(n19649), .C2(n19346), .A(n19305), .B(n19304), .ZN(
        P2_U3065) );
  AOI22_X1 U22282 ( .A1(n19318), .A2(n19693), .B1(n19692), .B2(n19317), .ZN(
        n19307) );
  AOI22_X1 U22283 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19320), .B1(
        n19319), .B2(n19581), .ZN(n19306) );
  OAI211_X1 U22284 ( .C1(n19528), .C2(n19346), .A(n19307), .B(n19306), .ZN(
        P2_U3066) );
  AOI22_X1 U22285 ( .A1(n19318), .A2(n19699), .B1(n19698), .B2(n19317), .ZN(
        n19309) );
  AOI22_X1 U22286 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19320), .B1(
        n19348), .B2(n19700), .ZN(n19308) );
  OAI211_X1 U22287 ( .C1(n19703), .C2(n19316), .A(n19309), .B(n19308), .ZN(
        P2_U3067) );
  AOI22_X1 U22288 ( .A1(n19318), .A2(n19705), .B1(n19704), .B2(n19317), .ZN(
        n19311) );
  AOI22_X1 U22289 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19320), .B1(
        n19319), .B2(n19706), .ZN(n19310) );
  OAI211_X1 U22290 ( .C1(n19709), .C2(n19346), .A(n19311), .B(n19310), .ZN(
        P2_U3068) );
  AOI22_X1 U22291 ( .A1(n19318), .A2(n19710), .B1(n19238), .B2(n19317), .ZN(
        n19313) );
  AOI22_X1 U22292 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19320), .B1(
        n19319), .B2(n19711), .ZN(n19312) );
  OAI211_X1 U22293 ( .C1(n19714), .C2(n19346), .A(n19313), .B(n19312), .ZN(
        P2_U3069) );
  AOI22_X1 U22294 ( .A1(n19318), .A2(n19716), .B1(n19715), .B2(n19317), .ZN(
        n19315) );
  AOI22_X1 U22295 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19320), .B1(
        n19348), .B2(n19568), .ZN(n19314) );
  OAI211_X1 U22296 ( .C1(n19571), .C2(n19316), .A(n19315), .B(n19314), .ZN(
        P2_U3070) );
  AOI22_X1 U22297 ( .A1(n19318), .A2(n19725), .B1(n19723), .B2(n19317), .ZN(
        n19322) );
  AOI22_X1 U22298 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19320), .B1(
        n19319), .B2(n19665), .ZN(n19321) );
  OAI211_X1 U22299 ( .C1(n19670), .C2(n19346), .A(n19322), .B(n19321), .ZN(
        P2_U3071) );
  NOR2_X1 U22300 ( .A1(n19545), .A2(n19324), .ZN(n19347) );
  AOI22_X1 U22301 ( .A1(n19632), .A2(n19348), .B1(n19673), .B2(n19347), .ZN(
        n19333) );
  OAI21_X1 U22302 ( .B1(n19435), .B2(n19323), .A(n19820), .ZN(n19331) );
  NOR2_X1 U22303 ( .A1(n10670), .A2(n19324), .ZN(n19328) );
  OAI21_X1 U22304 ( .B1(n12007), .B2(n10692), .A(n19385), .ZN(n19326) );
  INV_X1 U22305 ( .A(n19347), .ZN(n19325) );
  AOI21_X1 U22306 ( .B1(n19326), .B2(n19325), .A(n19436), .ZN(n19327) );
  OAI21_X1 U22307 ( .B1(n19331), .B2(n19328), .A(n19327), .ZN(n19350) );
  INV_X1 U22308 ( .A(n19328), .ZN(n19330) );
  OAI21_X1 U22309 ( .B1(n12007), .B2(n19347), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19329) );
  OAI21_X1 U22310 ( .B1(n19331), .B2(n19330), .A(n19329), .ZN(n19349) );
  AOI22_X1 U22311 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19350), .B1(
        n19674), .B2(n19349), .ZN(n19332) );
  OAI211_X1 U22312 ( .C1(n19645), .C2(n19366), .A(n19333), .B(n19332), .ZN(
        P2_U3072) );
  INV_X1 U22313 ( .A(n19649), .ZN(n19688) );
  AOI22_X1 U22314 ( .A1(n19688), .A2(n19381), .B1(n19686), .B2(n19347), .ZN(
        n19335) );
  AOI22_X1 U22315 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19350), .B1(
        n19687), .B2(n19349), .ZN(n19334) );
  OAI211_X1 U22316 ( .C1(n19691), .C2(n19346), .A(n19335), .B(n19334), .ZN(
        P2_U3073) );
  AOI22_X1 U22317 ( .A1(n19581), .A2(n19348), .B1(n19347), .B2(n19692), .ZN(
        n19337) );
  AOI22_X1 U22318 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19350), .B1(
        n19693), .B2(n19349), .ZN(n19336) );
  OAI211_X1 U22319 ( .C1(n19528), .C2(n19366), .A(n19337), .B(n19336), .ZN(
        P2_U3074) );
  AOI22_X1 U22320 ( .A1(n19653), .A2(n19348), .B1(n19347), .B2(n19698), .ZN(
        n19339) );
  AOI22_X1 U22321 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19350), .B1(
        n19699), .B2(n19349), .ZN(n19338) );
  OAI211_X1 U22322 ( .C1(n19656), .C2(n19366), .A(n19339), .B(n19338), .ZN(
        P2_U3075) );
  AOI22_X1 U22323 ( .A1(n19706), .A2(n19348), .B1(n19347), .B2(n19704), .ZN(
        n19341) );
  AOI22_X1 U22324 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19350), .B1(
        n19705), .B2(n19349), .ZN(n19340) );
  OAI211_X1 U22325 ( .C1(n19709), .C2(n19366), .A(n19341), .B(n19340), .ZN(
        P2_U3076) );
  AOI22_X1 U22326 ( .A1(n19711), .A2(n19348), .B1(n19347), .B2(n19238), .ZN(
        n19343) );
  AOI22_X1 U22327 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19350), .B1(
        n19710), .B2(n19349), .ZN(n19342) );
  OAI211_X1 U22328 ( .C1(n19714), .C2(n19366), .A(n19343), .B(n19342), .ZN(
        P2_U3077) );
  AOI22_X1 U22329 ( .A1(n19568), .A2(n19381), .B1(n19347), .B2(n19715), .ZN(
        n19345) );
  AOI22_X1 U22330 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19350), .B1(
        n19716), .B2(n19349), .ZN(n19344) );
  OAI211_X1 U22331 ( .C1(n19571), .C2(n19346), .A(n19345), .B(n19344), .ZN(
        P2_U3078) );
  AOI22_X1 U22332 ( .A1(n19665), .A2(n19348), .B1(n19347), .B2(n19723), .ZN(
        n19352) );
  AOI22_X1 U22333 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19350), .B1(
        n19725), .B2(n19349), .ZN(n19351) );
  OAI211_X1 U22334 ( .C1(n19670), .C2(n19366), .A(n19352), .B(n19351), .ZN(
        P2_U3079) );
  NAND2_X1 U22335 ( .A1(n12376), .A2(n19389), .ZN(n19360) );
  INV_X1 U22336 ( .A(n19360), .ZN(n19379) );
  NAND2_X1 U22337 ( .A1(n19354), .A2(n19824), .ZN(n19356) );
  OAI21_X1 U22338 ( .B1(n19356), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n10692), 
        .ZN(n19355) );
  AND2_X1 U22339 ( .A1(n19358), .A2(n19355), .ZN(n19380) );
  AOI22_X1 U22340 ( .A1(n19380), .A2(n19674), .B1(n19673), .B2(n19379), .ZN(
        n19365) );
  INV_X1 U22341 ( .A(n19356), .ZN(n19363) );
  AOI21_X1 U22342 ( .B1(n19366), .B2(n19413), .A(n19868), .ZN(n19362) );
  INV_X1 U22343 ( .A(n19358), .ZN(n19359) );
  AOI211_X1 U22344 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19360), .A(n19436), 
        .B(n19359), .ZN(n19361) );
  AOI22_X1 U22345 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19382), .B1(
        n19401), .B2(n19682), .ZN(n19364) );
  OAI211_X1 U22346 ( .C1(n19685), .C2(n19366), .A(n19365), .B(n19364), .ZN(
        P2_U3080) );
  AOI22_X1 U22347 ( .A1(n19380), .A2(n19687), .B1(n19686), .B2(n19379), .ZN(
        n19368) );
  AOI22_X1 U22348 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19382), .B1(
        n19381), .B2(n19646), .ZN(n19367) );
  OAI211_X1 U22349 ( .C1(n19649), .C2(n19413), .A(n19368), .B(n19367), .ZN(
        P2_U3081) );
  AOI22_X1 U22350 ( .A1(n19380), .A2(n19693), .B1(n19692), .B2(n19379), .ZN(
        n19370) );
  AOI22_X1 U22351 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19382), .B1(
        n19381), .B2(n19581), .ZN(n19369) );
  OAI211_X1 U22352 ( .C1(n19528), .C2(n19413), .A(n19370), .B(n19369), .ZN(
        P2_U3082) );
  AOI22_X1 U22353 ( .A1(n19380), .A2(n19699), .B1(n19698), .B2(n19379), .ZN(
        n19372) );
  AOI22_X1 U22354 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19382), .B1(
        n19381), .B2(n19653), .ZN(n19371) );
  OAI211_X1 U22355 ( .C1(n19656), .C2(n19413), .A(n19372), .B(n19371), .ZN(
        P2_U3083) );
  AOI22_X1 U22356 ( .A1(n19380), .A2(n19705), .B1(n19704), .B2(n19379), .ZN(
        n19374) );
  AOI22_X1 U22357 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19382), .B1(
        n19381), .B2(n19706), .ZN(n19373) );
  OAI211_X1 U22358 ( .C1(n19709), .C2(n19413), .A(n19374), .B(n19373), .ZN(
        P2_U3084) );
  AOI22_X1 U22359 ( .A1(n19380), .A2(n19710), .B1(n19238), .B2(n19379), .ZN(
        n19376) );
  AOI22_X1 U22360 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19382), .B1(
        n19381), .B2(n19711), .ZN(n19375) );
  OAI211_X1 U22361 ( .C1(n19714), .C2(n19413), .A(n19376), .B(n19375), .ZN(
        P2_U3085) );
  AOI22_X1 U22362 ( .A1(n19380), .A2(n19716), .B1(n19715), .B2(n19379), .ZN(
        n19378) );
  AOI22_X1 U22363 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19382), .B1(
        n19381), .B2(n19717), .ZN(n19377) );
  OAI211_X1 U22364 ( .C1(n19722), .C2(n19413), .A(n19378), .B(n19377), .ZN(
        P2_U3086) );
  AOI22_X1 U22365 ( .A1(n19380), .A2(n19725), .B1(n19723), .B2(n19379), .ZN(
        n19384) );
  AOI22_X1 U22366 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19382), .B1(
        n19381), .B2(n19665), .ZN(n19383) );
  OAI211_X1 U22367 ( .C1(n19670), .C2(n19413), .A(n19384), .B(n19383), .ZN(
        P2_U3087) );
  AOI22_X1 U22368 ( .A1(n19682), .A2(n19424), .B1(n19673), .B2(n19408), .ZN(
        n19394) );
  OAI21_X1 U22369 ( .B1(n19435), .B2(n19609), .A(n19820), .ZN(n19392) );
  NAND2_X1 U22370 ( .A1(n12030), .A2(n19385), .ZN(n19387) );
  INV_X1 U22371 ( .A(n19408), .ZN(n19386) );
  NAND3_X1 U22372 ( .A1(n19387), .A2(n19636), .A3(n19386), .ZN(n19388) );
  OAI211_X1 U22373 ( .C1(n19392), .C2(n19389), .A(n19680), .B(n19388), .ZN(
        n19410) );
  OAI21_X1 U22374 ( .B1(n12030), .B2(n19408), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19390) );
  OAI21_X1 U22375 ( .B1(n19392), .B2(n19391), .A(n19390), .ZN(n19409) );
  AOI22_X1 U22376 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19410), .B1(
        n19674), .B2(n19409), .ZN(n19393) );
  OAI211_X1 U22377 ( .C1(n19685), .C2(n19413), .A(n19394), .B(n19393), .ZN(
        P2_U3088) );
  AOI22_X1 U22378 ( .A1(n19688), .A2(n19424), .B1(n19686), .B2(n19408), .ZN(
        n19396) );
  AOI22_X1 U22379 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19410), .B1(
        n19687), .B2(n19409), .ZN(n19395) );
  OAI211_X1 U22380 ( .C1(n19691), .C2(n19413), .A(n19396), .B(n19395), .ZN(
        P2_U3089) );
  AOI22_X1 U22381 ( .A1(n19581), .A2(n19401), .B1(n19692), .B2(n19408), .ZN(
        n19398) );
  AOI22_X1 U22382 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19410), .B1(
        n19693), .B2(n19409), .ZN(n19397) );
  OAI211_X1 U22383 ( .C1(n19528), .C2(n19432), .A(n19398), .B(n19397), .ZN(
        P2_U3090) );
  AOI22_X1 U22384 ( .A1(n19653), .A2(n19401), .B1(n19408), .B2(n19698), .ZN(
        n19400) );
  AOI22_X1 U22385 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19410), .B1(
        n19699), .B2(n19409), .ZN(n19399) );
  OAI211_X1 U22386 ( .C1(n19656), .C2(n19432), .A(n19400), .B(n19399), .ZN(
        P2_U3091) );
  AOI22_X1 U22387 ( .A1(n19706), .A2(n19401), .B1(n19408), .B2(n19704), .ZN(
        n19403) );
  AOI22_X1 U22388 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19410), .B1(
        n19705), .B2(n19409), .ZN(n19402) );
  OAI211_X1 U22389 ( .C1(n19709), .C2(n19432), .A(n19403), .B(n19402), .ZN(
        P2_U3092) );
  AOI22_X1 U22390 ( .A1(n19564), .A2(n19424), .B1(n19408), .B2(n19238), .ZN(
        n19405) );
  AOI22_X1 U22391 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19410), .B1(
        n19710), .B2(n19409), .ZN(n19404) );
  OAI211_X1 U22392 ( .C1(n19567), .C2(n19413), .A(n19405), .B(n19404), .ZN(
        P2_U3093) );
  AOI22_X1 U22393 ( .A1(n19568), .A2(n19424), .B1(n19715), .B2(n19408), .ZN(
        n19407) );
  AOI22_X1 U22394 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19410), .B1(
        n19716), .B2(n19409), .ZN(n19406) );
  OAI211_X1 U22395 ( .C1(n19571), .C2(n19413), .A(n19407), .B(n19406), .ZN(
        P2_U3094) );
  AOI22_X1 U22396 ( .A1(n19727), .A2(n19424), .B1(n19408), .B2(n19723), .ZN(
        n19412) );
  AOI22_X1 U22397 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19410), .B1(
        n19725), .B2(n19409), .ZN(n19411) );
  OAI211_X1 U22398 ( .C1(n19733), .C2(n19413), .A(n19412), .B(n19411), .ZN(
        P2_U3095) );
  AOI22_X1 U22399 ( .A1(n19428), .A2(n19687), .B1(n19427), .B2(n19686), .ZN(
        n19415) );
  AOI22_X1 U22400 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19429), .B1(
        n19448), .B2(n19688), .ZN(n19414) );
  OAI211_X1 U22401 ( .C1(n19691), .C2(n19432), .A(n19415), .B(n19414), .ZN(
        P2_U3097) );
  AOI22_X1 U22402 ( .A1(n19428), .A2(n19693), .B1(n19427), .B2(n19692), .ZN(
        n19417) );
  AOI22_X1 U22403 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19429), .B1(
        n19448), .B2(n19694), .ZN(n19416) );
  OAI211_X1 U22404 ( .C1(n19697), .C2(n19432), .A(n19417), .B(n19416), .ZN(
        P2_U3098) );
  AOI22_X1 U22405 ( .A1(n19428), .A2(n19699), .B1(n19427), .B2(n19698), .ZN(
        n19419) );
  AOI22_X1 U22406 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19429), .B1(
        n19424), .B2(n19653), .ZN(n19418) );
  OAI211_X1 U22407 ( .C1(n19656), .C2(n19459), .A(n19419), .B(n19418), .ZN(
        P2_U3099) );
  AOI22_X1 U22408 ( .A1(n19428), .A2(n19705), .B1(n19427), .B2(n19704), .ZN(
        n19421) );
  AOI22_X1 U22409 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19429), .B1(
        n19424), .B2(n19706), .ZN(n19420) );
  OAI211_X1 U22410 ( .C1(n19709), .C2(n19459), .A(n19421), .B(n19420), .ZN(
        P2_U3100) );
  AOI22_X1 U22411 ( .A1(n19428), .A2(n19710), .B1(n19427), .B2(n19238), .ZN(
        n19423) );
  AOI22_X1 U22412 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19429), .B1(
        n19448), .B2(n19564), .ZN(n19422) );
  OAI211_X1 U22413 ( .C1(n19567), .C2(n19432), .A(n19423), .B(n19422), .ZN(
        P2_U3101) );
  AOI22_X1 U22414 ( .A1(n19428), .A2(n19716), .B1(n19427), .B2(n19715), .ZN(
        n19426) );
  AOI22_X1 U22415 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19429), .B1(
        n19424), .B2(n19717), .ZN(n19425) );
  OAI211_X1 U22416 ( .C1(n19722), .C2(n19459), .A(n19426), .B(n19425), .ZN(
        P2_U3102) );
  AOI22_X1 U22417 ( .A1(n19428), .A2(n19725), .B1(n19427), .B2(n19723), .ZN(
        n19431) );
  AOI22_X1 U22418 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19429), .B1(
        n19448), .B2(n19727), .ZN(n19430) );
  OAI211_X1 U22419 ( .C1(n19733), .C2(n19432), .A(n19431), .B(n19430), .ZN(
        P2_U3103) );
  NOR2_X1 U22420 ( .A1(n12376), .A2(n19434), .ZN(n19467) );
  AOI22_X1 U22421 ( .A1(n19455), .A2(n19674), .B1(n19673), .B2(n19467), .ZN(
        n19441) );
  INV_X1 U22422 ( .A(n19434), .ZN(n19438) );
  NOR2_X1 U22423 ( .A1(n19435), .A2(n19815), .ZN(n19819) );
  INV_X1 U22424 ( .A(n19467), .ZN(n19464) );
  AOI211_X1 U22425 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19464), .A(n19436), 
        .B(n9838), .ZN(n19437) );
  OAI21_X1 U22426 ( .B1(n19438), .B2(n19819), .A(n19437), .ZN(n19456) );
  AOI22_X1 U22427 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19456), .B1(
        n19486), .B2(n19682), .ZN(n19440) );
  OAI211_X1 U22428 ( .C1(n19685), .C2(n19459), .A(n19441), .B(n19440), .ZN(
        P2_U3104) );
  AOI22_X1 U22429 ( .A1(n19455), .A2(n19687), .B1(n19686), .B2(n19467), .ZN(
        n19443) );
  AOI22_X1 U22430 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19456), .B1(
        n19448), .B2(n19646), .ZN(n19442) );
  OAI211_X1 U22431 ( .C1(n19649), .C2(n19484), .A(n19443), .B(n19442), .ZN(
        P2_U3105) );
  AOI22_X1 U22432 ( .A1(n19455), .A2(n19693), .B1(n19692), .B2(n19467), .ZN(
        n19445) );
  AOI22_X1 U22433 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19456), .B1(
        n19448), .B2(n19581), .ZN(n19444) );
  OAI211_X1 U22434 ( .C1(n19528), .C2(n19484), .A(n19445), .B(n19444), .ZN(
        P2_U3106) );
  AOI22_X1 U22435 ( .A1(n19455), .A2(n19699), .B1(n19698), .B2(n19467), .ZN(
        n19447) );
  AOI22_X1 U22436 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19456), .B1(
        n19448), .B2(n19653), .ZN(n19446) );
  OAI211_X1 U22437 ( .C1(n19656), .C2(n19484), .A(n19447), .B(n19446), .ZN(
        P2_U3107) );
  AOI22_X1 U22438 ( .A1(n19455), .A2(n19705), .B1(n19704), .B2(n19467), .ZN(
        n19450) );
  AOI22_X1 U22439 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19456), .B1(
        n19448), .B2(n19706), .ZN(n19449) );
  OAI211_X1 U22440 ( .C1(n19709), .C2(n19484), .A(n19450), .B(n19449), .ZN(
        P2_U3108) );
  AOI22_X1 U22441 ( .A1(n19455), .A2(n19710), .B1(n19238), .B2(n19467), .ZN(
        n19452) );
  AOI22_X1 U22442 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19456), .B1(
        n19486), .B2(n19564), .ZN(n19451) );
  OAI211_X1 U22443 ( .C1(n19567), .C2(n19459), .A(n19452), .B(n19451), .ZN(
        P2_U3109) );
  AOI22_X1 U22444 ( .A1(n19455), .A2(n19716), .B1(n19715), .B2(n19467), .ZN(
        n19454) );
  AOI22_X1 U22445 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19456), .B1(
        n19486), .B2(n19568), .ZN(n19453) );
  OAI211_X1 U22446 ( .C1(n19571), .C2(n19459), .A(n19454), .B(n19453), .ZN(
        P2_U3110) );
  AOI22_X1 U22447 ( .A1(n19455), .A2(n19725), .B1(n19723), .B2(n19467), .ZN(
        n19458) );
  AOI22_X1 U22448 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19456), .B1(
        n19486), .B2(n19727), .ZN(n19457) );
  OAI211_X1 U22449 ( .C1(n19733), .C2(n19459), .A(n19458), .B(n19457), .ZN(
        P2_U3111) );
  INV_X1 U22450 ( .A(n19521), .ZN(n19509) );
  NOR2_X1 U22451 ( .A1(n19544), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19496) );
  INV_X1 U22452 ( .A(n19496), .ZN(n19499) );
  NOR2_X1 U22453 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19499), .ZN(
        n19485) );
  AOI22_X1 U22454 ( .A1(n19682), .A2(n19509), .B1(n19673), .B2(n19485), .ZN(
        n19471) );
  AOI21_X1 U22455 ( .B1(n19484), .B2(n19521), .A(n19868), .ZN(n19462) );
  NOR2_X1 U22456 ( .A1(n19462), .A2(n19636), .ZN(n19466) );
  OAI21_X1 U22457 ( .B1(n11999), .B2(n10692), .A(n19385), .ZN(n19463) );
  AOI21_X1 U22458 ( .B1(n19466), .B2(n19464), .A(n19463), .ZN(n19465) );
  OAI21_X1 U22459 ( .B1(n19485), .B2(n19465), .A(n19680), .ZN(n19488) );
  OAI21_X1 U22460 ( .B1(n19485), .B2(n19467), .A(n19466), .ZN(n19469) );
  OAI21_X1 U22461 ( .B1(n11999), .B2(n19485), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19468) );
  NAND2_X1 U22462 ( .A1(n19469), .A2(n19468), .ZN(n19487) );
  AOI22_X1 U22463 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19488), .B1(
        n19674), .B2(n19487), .ZN(n19470) );
  OAI211_X1 U22464 ( .C1(n19685), .C2(n19484), .A(n19471), .B(n19470), .ZN(
        P2_U3112) );
  AOI22_X1 U22465 ( .A1(n19646), .A2(n19486), .B1(n19686), .B2(n19485), .ZN(
        n19473) );
  AOI22_X1 U22466 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19488), .B1(
        n19687), .B2(n19487), .ZN(n19472) );
  OAI211_X1 U22467 ( .C1(n19649), .C2(n19521), .A(n19473), .B(n19472), .ZN(
        P2_U3113) );
  AOI22_X1 U22468 ( .A1(n19581), .A2(n19486), .B1(n19692), .B2(n19485), .ZN(
        n19475) );
  AOI22_X1 U22469 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19488), .B1(
        n19693), .B2(n19487), .ZN(n19474) );
  OAI211_X1 U22470 ( .C1(n19528), .C2(n19521), .A(n19475), .B(n19474), .ZN(
        P2_U3114) );
  AOI22_X1 U22471 ( .A1(n19700), .A2(n19509), .B1(n19698), .B2(n19485), .ZN(
        n19477) );
  AOI22_X1 U22472 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19488), .B1(
        n19699), .B2(n19487), .ZN(n19476) );
  OAI211_X1 U22473 ( .C1(n19703), .C2(n19484), .A(n19477), .B(n19476), .ZN(
        P2_U3115) );
  AOI22_X1 U22474 ( .A1(n19706), .A2(n19486), .B1(n19704), .B2(n19485), .ZN(
        n19479) );
  AOI22_X1 U22475 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19488), .B1(
        n19705), .B2(n19487), .ZN(n19478) );
  OAI211_X1 U22476 ( .C1(n19709), .C2(n19521), .A(n19479), .B(n19478), .ZN(
        P2_U3116) );
  AOI22_X1 U22477 ( .A1(n19711), .A2(n19486), .B1(n19238), .B2(n19485), .ZN(
        n19481) );
  AOI22_X1 U22478 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19488), .B1(
        n19710), .B2(n19487), .ZN(n19480) );
  OAI211_X1 U22479 ( .C1(n19714), .C2(n19521), .A(n19481), .B(n19480), .ZN(
        P2_U3117) );
  AOI22_X1 U22480 ( .A1(n19568), .A2(n19509), .B1(n19715), .B2(n19485), .ZN(
        n19483) );
  AOI22_X1 U22481 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19488), .B1(
        n19716), .B2(n19487), .ZN(n19482) );
  OAI211_X1 U22482 ( .C1(n19571), .C2(n19484), .A(n19483), .B(n19482), .ZN(
        P2_U3118) );
  AOI22_X1 U22483 ( .A1(n19665), .A2(n19486), .B1(n19723), .B2(n19485), .ZN(
        n19490) );
  AOI22_X1 U22484 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19488), .B1(
        n19725), .B2(n19487), .ZN(n19489) );
  OAI211_X1 U22485 ( .C1(n19670), .C2(n19521), .A(n19490), .B(n19489), .ZN(
        P2_U3119) );
  AOI22_X1 U22486 ( .A1(n19682), .A2(n19540), .B1(n19673), .B2(n19516), .ZN(
        n19502) );
  NOR2_X1 U22487 ( .A1(n19818), .A2(n19868), .ZN(n19676) );
  INV_X1 U22488 ( .A(n19676), .ZN(n19492) );
  OAI21_X1 U22489 ( .B1(n19492), .B2(n19491), .A(n19820), .ZN(n19500) );
  INV_X1 U22490 ( .A(n19516), .ZN(n19493) );
  OAI211_X1 U22491 ( .C1(n19494), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19493), 
        .B(n19636), .ZN(n19495) );
  OAI211_X1 U22492 ( .C1(n19500), .C2(n19496), .A(n19680), .B(n19495), .ZN(
        n19518) );
  OAI21_X1 U22493 ( .B1(n19497), .B2(n19516), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19498) );
  OAI21_X1 U22494 ( .B1(n19500), .B2(n19499), .A(n19498), .ZN(n19517) );
  AOI22_X1 U22495 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19518), .B1(
        n19674), .B2(n19517), .ZN(n19501) );
  OAI211_X1 U22496 ( .C1(n19685), .C2(n19521), .A(n19502), .B(n19501), .ZN(
        P2_U3120) );
  AOI22_X1 U22497 ( .A1(n19688), .A2(n19540), .B1(n19686), .B2(n19516), .ZN(
        n19504) );
  AOI22_X1 U22498 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19518), .B1(
        n19687), .B2(n19517), .ZN(n19503) );
  OAI211_X1 U22499 ( .C1(n19691), .C2(n19521), .A(n19504), .B(n19503), .ZN(
        P2_U3121) );
  AOI22_X1 U22500 ( .A1(n19694), .A2(n19540), .B1(n19692), .B2(n19516), .ZN(
        n19506) );
  AOI22_X1 U22501 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19518), .B1(
        n19693), .B2(n19517), .ZN(n19505) );
  OAI211_X1 U22502 ( .C1(n19697), .C2(n19521), .A(n19506), .B(n19505), .ZN(
        P2_U3122) );
  AOI22_X1 U22503 ( .A1(n19700), .A2(n19540), .B1(n19698), .B2(n19516), .ZN(
        n19508) );
  AOI22_X1 U22504 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19518), .B1(
        n19699), .B2(n19517), .ZN(n19507) );
  OAI211_X1 U22505 ( .C1(n19703), .C2(n19521), .A(n19508), .B(n19507), .ZN(
        P2_U3123) );
  AOI22_X1 U22506 ( .A1(n19706), .A2(n19509), .B1(n19704), .B2(n19516), .ZN(
        n19511) );
  AOI22_X1 U22507 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19518), .B1(
        n19705), .B2(n19517), .ZN(n19510) );
  OAI211_X1 U22508 ( .C1(n19709), .C2(n19537), .A(n19511), .B(n19510), .ZN(
        P2_U3124) );
  AOI22_X1 U22509 ( .A1(n19564), .A2(n19540), .B1(n19238), .B2(n19516), .ZN(
        n19513) );
  AOI22_X1 U22510 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19518), .B1(
        n19710), .B2(n19517), .ZN(n19512) );
  OAI211_X1 U22511 ( .C1(n19567), .C2(n19521), .A(n19513), .B(n19512), .ZN(
        P2_U3125) );
  AOI22_X1 U22512 ( .A1(n19568), .A2(n19540), .B1(n19715), .B2(n19516), .ZN(
        n19515) );
  AOI22_X1 U22513 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19518), .B1(
        n19716), .B2(n19517), .ZN(n19514) );
  OAI211_X1 U22514 ( .C1(n19571), .C2(n19521), .A(n19515), .B(n19514), .ZN(
        P2_U3126) );
  AOI22_X1 U22515 ( .A1(n19727), .A2(n19540), .B1(n19723), .B2(n19516), .ZN(
        n19520) );
  AOI22_X1 U22516 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19518), .B1(
        n19725), .B2(n19517), .ZN(n19519) );
  OAI211_X1 U22517 ( .C1(n19733), .C2(n19521), .A(n19520), .B(n19519), .ZN(
        P2_U3127) );
  AOI22_X1 U22518 ( .A1(n19539), .A2(n19687), .B1(n19686), .B2(n19538), .ZN(
        n19523) );
  AOI22_X1 U22519 ( .A1(n19540), .A2(n19646), .B1(n19560), .B2(n19688), .ZN(
        n19522) );
  OAI211_X1 U22520 ( .C1(n19525), .C2(n19524), .A(n19523), .B(n19522), .ZN(
        P2_U3129) );
  AOI22_X1 U22521 ( .A1(n19539), .A2(n19693), .B1(n19692), .B2(n19538), .ZN(
        n19527) );
  AOI22_X1 U22522 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19541), .B1(
        n19540), .B2(n19581), .ZN(n19526) );
  OAI211_X1 U22523 ( .C1(n19528), .C2(n19577), .A(n19527), .B(n19526), .ZN(
        P2_U3130) );
  AOI22_X1 U22524 ( .A1(n19539), .A2(n19699), .B1(n19698), .B2(n19538), .ZN(
        n19530) );
  AOI22_X1 U22525 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19541), .B1(
        n19560), .B2(n19700), .ZN(n19529) );
  OAI211_X1 U22526 ( .C1(n19703), .C2(n19537), .A(n19530), .B(n19529), .ZN(
        P2_U3131) );
  AOI22_X1 U22527 ( .A1(n19539), .A2(n19705), .B1(n19704), .B2(n19538), .ZN(
        n19532) );
  AOI22_X1 U22528 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19541), .B1(
        n19540), .B2(n19706), .ZN(n19531) );
  OAI211_X1 U22529 ( .C1(n19709), .C2(n19577), .A(n19532), .B(n19531), .ZN(
        P2_U3132) );
  AOI22_X1 U22530 ( .A1(n19539), .A2(n19710), .B1(n19238), .B2(n19538), .ZN(
        n19534) );
  AOI22_X1 U22531 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19541), .B1(
        n19540), .B2(n19711), .ZN(n19533) );
  OAI211_X1 U22532 ( .C1(n19714), .C2(n19577), .A(n19534), .B(n19533), .ZN(
        P2_U3133) );
  AOI22_X1 U22533 ( .A1(n19539), .A2(n19716), .B1(n19715), .B2(n19538), .ZN(
        n19536) );
  AOI22_X1 U22534 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19541), .B1(
        n19560), .B2(n19568), .ZN(n19535) );
  OAI211_X1 U22535 ( .C1(n19571), .C2(n19537), .A(n19536), .B(n19535), .ZN(
        P2_U3134) );
  AOI22_X1 U22536 ( .A1(n19539), .A2(n19725), .B1(n19723), .B2(n19538), .ZN(
        n19543) );
  AOI22_X1 U22537 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19541), .B1(
        n19540), .B2(n19665), .ZN(n19542) );
  OAI211_X1 U22538 ( .C1(n19670), .C2(n19577), .A(n19543), .B(n19542), .ZN(
        P2_U3135) );
  OR2_X1 U22539 ( .A1(n10670), .A2(n19544), .ZN(n19549) );
  OR2_X1 U22540 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19549), .ZN(n19546) );
  NOR2_X1 U22541 ( .A1(n19545), .A2(n19544), .ZN(n19572) );
  NOR3_X1 U22542 ( .A1(n12000), .A2(n19572), .A3(n10692), .ZN(n19548) );
  AOI21_X1 U22543 ( .B1(n10692), .B2(n19546), .A(n19548), .ZN(n19573) );
  AOI22_X1 U22544 ( .A1(n19573), .A2(n19674), .B1(n19673), .B2(n19572), .ZN(
        n19553) );
  NAND2_X1 U22545 ( .A1(n19676), .A2(n19547), .ZN(n19550) );
  AOI21_X1 U22546 ( .B1(n19550), .B2(n19549), .A(n19548), .ZN(n19551) );
  OAI211_X1 U22547 ( .C1(n19572), .C2(n19385), .A(n19551), .B(n19680), .ZN(
        n19574) );
  AOI22_X1 U22548 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19574), .B1(
        n19596), .B2(n19682), .ZN(n19552) );
  OAI211_X1 U22549 ( .C1(n19685), .C2(n19577), .A(n19553), .B(n19552), .ZN(
        P2_U3136) );
  AOI22_X1 U22550 ( .A1(n19573), .A2(n19687), .B1(n19686), .B2(n19572), .ZN(
        n19555) );
  AOI22_X1 U22551 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19574), .B1(
        n19596), .B2(n19688), .ZN(n19554) );
  OAI211_X1 U22552 ( .C1(n19691), .C2(n19577), .A(n19555), .B(n19554), .ZN(
        P2_U3137) );
  AOI22_X1 U22553 ( .A1(n19573), .A2(n19693), .B1(n19692), .B2(n19572), .ZN(
        n19557) );
  AOI22_X1 U22554 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19574), .B1(
        n19596), .B2(n19694), .ZN(n19556) );
  OAI211_X1 U22555 ( .C1(n19697), .C2(n19577), .A(n19557), .B(n19556), .ZN(
        P2_U3138) );
  AOI22_X1 U22556 ( .A1(n19573), .A2(n19699), .B1(n19698), .B2(n19572), .ZN(
        n19559) );
  AOI22_X1 U22557 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19574), .B1(
        n19596), .B2(n19700), .ZN(n19558) );
  OAI211_X1 U22558 ( .C1(n19703), .C2(n19577), .A(n19559), .B(n19558), .ZN(
        P2_U3139) );
  AOI22_X1 U22559 ( .A1(n19573), .A2(n19705), .B1(n19704), .B2(n19572), .ZN(
        n19562) );
  AOI22_X1 U22560 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19574), .B1(
        n19560), .B2(n19706), .ZN(n19561) );
  OAI211_X1 U22561 ( .C1(n19709), .C2(n19563), .A(n19562), .B(n19561), .ZN(
        P2_U3140) );
  AOI22_X1 U22562 ( .A1(n19573), .A2(n19710), .B1(n19238), .B2(n19572), .ZN(
        n19566) );
  AOI22_X1 U22563 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19574), .B1(
        n19596), .B2(n19564), .ZN(n19565) );
  OAI211_X1 U22564 ( .C1(n19567), .C2(n19577), .A(n19566), .B(n19565), .ZN(
        P2_U3141) );
  AOI22_X1 U22565 ( .A1(n19573), .A2(n19716), .B1(n19715), .B2(n19572), .ZN(
        n19570) );
  AOI22_X1 U22566 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19574), .B1(
        n19596), .B2(n19568), .ZN(n19569) );
  OAI211_X1 U22567 ( .C1(n19571), .C2(n19577), .A(n19570), .B(n19569), .ZN(
        P2_U3142) );
  AOI22_X1 U22568 ( .A1(n19573), .A2(n19725), .B1(n19723), .B2(n19572), .ZN(
        n19576) );
  AOI22_X1 U22569 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19574), .B1(
        n19596), .B2(n19727), .ZN(n19575) );
  OAI211_X1 U22570 ( .C1(n19733), .C2(n19577), .A(n19576), .B(n19575), .ZN(
        P2_U3143) );
  INV_X1 U22571 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n19580) );
  AOI22_X1 U22572 ( .A1(n19595), .A2(n19687), .B1(n19686), .B2(n19594), .ZN(
        n19579) );
  AOI22_X1 U22573 ( .A1(n19596), .A2(n19646), .B1(n19623), .B2(n19688), .ZN(
        n19578) );
  OAI211_X1 U22574 ( .C1(n19587), .C2(n19580), .A(n19579), .B(n19578), .ZN(
        P2_U3145) );
  INV_X1 U22575 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n19584) );
  AOI22_X1 U22576 ( .A1(n19595), .A2(n19693), .B1(n19692), .B2(n19594), .ZN(
        n19583) );
  AOI22_X1 U22577 ( .A1(n19596), .A2(n19581), .B1(n19623), .B2(n19694), .ZN(
        n19582) );
  OAI211_X1 U22578 ( .C1(n19587), .C2(n19584), .A(n19583), .B(n19582), .ZN(
        P2_U3146) );
  AOI22_X1 U22579 ( .A1(n19595), .A2(n19699), .B1(n19698), .B2(n19594), .ZN(
        n19586) );
  AOI22_X1 U22580 ( .A1(n19623), .A2(n19700), .B1(n19596), .B2(n19653), .ZN(
        n19585) );
  OAI211_X1 U22581 ( .C1(n19587), .C2(n10319), .A(n19586), .B(n19585), .ZN(
        P2_U3147) );
  AOI22_X1 U22582 ( .A1(n19595), .A2(n19705), .B1(n19704), .B2(n19594), .ZN(
        n19589) );
  AOI22_X1 U22583 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19597), .B1(
        n19596), .B2(n19706), .ZN(n19588) );
  OAI211_X1 U22584 ( .C1(n19709), .C2(n19630), .A(n19589), .B(n19588), .ZN(
        P2_U3148) );
  AOI22_X1 U22585 ( .A1(n19595), .A2(n19710), .B1(n19238), .B2(n19594), .ZN(
        n19591) );
  AOI22_X1 U22586 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19597), .B1(
        n19596), .B2(n19711), .ZN(n19590) );
  OAI211_X1 U22587 ( .C1(n19714), .C2(n19630), .A(n19591), .B(n19590), .ZN(
        P2_U3149) );
  AOI22_X1 U22588 ( .A1(n19595), .A2(n19716), .B1(n19715), .B2(n19594), .ZN(
        n19593) );
  AOI22_X1 U22589 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19597), .B1(
        n19596), .B2(n19717), .ZN(n19592) );
  OAI211_X1 U22590 ( .C1(n19722), .C2(n19630), .A(n19593), .B(n19592), .ZN(
        P2_U3150) );
  AOI22_X1 U22591 ( .A1(n19595), .A2(n19725), .B1(n19723), .B2(n19594), .ZN(
        n19599) );
  AOI22_X1 U22592 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19597), .B1(
        n19596), .B2(n19665), .ZN(n19598) );
  OAI211_X1 U22593 ( .C1(n19670), .C2(n19630), .A(n19599), .B(n19598), .ZN(
        P2_U3151) );
  OR2_X1 U22594 ( .A1(n19605), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19603) );
  NOR2_X1 U22595 ( .A1(n12376), .A2(n19605), .ZN(n19634) );
  INV_X1 U22596 ( .A(n19634), .ZN(n19600) );
  NAND3_X1 U22597 ( .A1(n19601), .A2(P2_STATE2_REG_2__SCAN_IN), .A3(n19600), 
        .ZN(n19607) );
  INV_X1 U22598 ( .A(n19607), .ZN(n19602) );
  AOI21_X1 U22599 ( .B1(n19603), .B2(n10692), .A(n19602), .ZN(n19626) );
  AOI22_X1 U22600 ( .A1(n19626), .A2(n19674), .B1(n19673), .B2(n19634), .ZN(
        n19612) );
  NAND2_X1 U22601 ( .A1(n19676), .A2(n19604), .ZN(n19606) );
  AOI21_X1 U22602 ( .B1(n19606), .B2(n19605), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n19608) );
  OAI211_X1 U22603 ( .C1(n19608), .C2(n19634), .A(n19680), .B(n19607), .ZN(
        n19627) );
  AOI22_X1 U22604 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19627), .B1(
        n19664), .B2(n19682), .ZN(n19611) );
  OAI211_X1 U22605 ( .C1(n19685), .C2(n19630), .A(n19612), .B(n19611), .ZN(
        P2_U3152) );
  INV_X1 U22606 ( .A(n19664), .ZN(n19652) );
  AOI22_X1 U22607 ( .A1(n19626), .A2(n19687), .B1(n19686), .B2(n19634), .ZN(
        n19614) );
  AOI22_X1 U22608 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19627), .B1(
        n19623), .B2(n19646), .ZN(n19613) );
  OAI211_X1 U22609 ( .C1(n19649), .C2(n19652), .A(n19614), .B(n19613), .ZN(
        P2_U3153) );
  AOI22_X1 U22610 ( .A1(n19626), .A2(n19693), .B1(n19692), .B2(n19634), .ZN(
        n19616) );
  AOI22_X1 U22611 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19627), .B1(
        n19664), .B2(n19694), .ZN(n19615) );
  OAI211_X1 U22612 ( .C1(n19697), .C2(n19630), .A(n19616), .B(n19615), .ZN(
        P2_U3154) );
  AOI22_X1 U22613 ( .A1(n19626), .A2(n19699), .B1(n19698), .B2(n19634), .ZN(
        n19618) );
  AOI22_X1 U22614 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19627), .B1(
        n19623), .B2(n19653), .ZN(n19617) );
  OAI211_X1 U22615 ( .C1(n19656), .C2(n19652), .A(n19618), .B(n19617), .ZN(
        P2_U3155) );
  AOI22_X1 U22616 ( .A1(n19626), .A2(n19705), .B1(n19704), .B2(n19634), .ZN(
        n19620) );
  AOI22_X1 U22617 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19627), .B1(
        n19623), .B2(n19706), .ZN(n19619) );
  OAI211_X1 U22618 ( .C1(n19709), .C2(n19652), .A(n19620), .B(n19619), .ZN(
        P2_U3156) );
  AOI22_X1 U22619 ( .A1(n19626), .A2(n19710), .B1(n19238), .B2(n19634), .ZN(
        n19622) );
  AOI22_X1 U22620 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19627), .B1(
        n19623), .B2(n19711), .ZN(n19621) );
  OAI211_X1 U22621 ( .C1(n19714), .C2(n19652), .A(n19622), .B(n19621), .ZN(
        P2_U3157) );
  AOI22_X1 U22622 ( .A1(n19626), .A2(n19716), .B1(n19715), .B2(n19634), .ZN(
        n19625) );
  AOI22_X1 U22623 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19627), .B1(
        n19623), .B2(n19717), .ZN(n19624) );
  OAI211_X1 U22624 ( .C1(n19722), .C2(n19652), .A(n19625), .B(n19624), .ZN(
        P2_U3158) );
  AOI22_X1 U22625 ( .A1(n19626), .A2(n19725), .B1(n19723), .B2(n19634), .ZN(
        n19629) );
  AOI22_X1 U22626 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19627), .B1(
        n19664), .B2(n19727), .ZN(n19628) );
  OAI211_X1 U22627 ( .C1(n19733), .C2(n19630), .A(n19629), .B(n19628), .ZN(
        P2_U3159) );
  AND3_X1 U22628 ( .A1(n12376), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        n19671), .ZN(n19663) );
  AOI22_X1 U22629 ( .A1(n19632), .A2(n19664), .B1(n19673), .B2(n19663), .ZN(
        n19644) );
  OAI21_X1 U22630 ( .B1(n19718), .B2(n19664), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19633) );
  NAND2_X1 U22631 ( .A1(n19633), .A2(n19820), .ZN(n19642) );
  NOR2_X1 U22632 ( .A1(n19663), .A2(n19634), .ZN(n19641) );
  INV_X1 U22633 ( .A(n19641), .ZN(n19639) );
  NAND2_X1 U22634 ( .A1(n12011), .A2(n19385), .ZN(n19637) );
  INV_X1 U22635 ( .A(n19663), .ZN(n19635) );
  NAND3_X1 U22636 ( .A1(n19637), .A2(n19636), .A3(n19635), .ZN(n19638) );
  OAI211_X1 U22637 ( .C1(n19642), .C2(n19639), .A(n19680), .B(n19638), .ZN(
        n19667) );
  OAI21_X1 U22638 ( .B1(n12011), .B2(n19663), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19640) );
  AOI22_X1 U22639 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19667), .B1(
        n19674), .B2(n19666), .ZN(n19643) );
  OAI211_X1 U22640 ( .C1(n19645), .C2(n19732), .A(n19644), .B(n19643), .ZN(
        P2_U3160) );
  AOI22_X1 U22641 ( .A1(n19646), .A2(n19664), .B1(n19686), .B2(n19663), .ZN(
        n19648) );
  AOI22_X1 U22642 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19667), .B1(
        n19687), .B2(n19666), .ZN(n19647) );
  OAI211_X1 U22643 ( .C1(n19649), .C2(n19732), .A(n19648), .B(n19647), .ZN(
        P2_U3161) );
  AOI22_X1 U22644 ( .A1(n19694), .A2(n19718), .B1(n19692), .B2(n19663), .ZN(
        n19651) );
  AOI22_X1 U22645 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19667), .B1(
        n19693), .B2(n19666), .ZN(n19650) );
  OAI211_X1 U22646 ( .C1(n19697), .C2(n19652), .A(n19651), .B(n19650), .ZN(
        P2_U3162) );
  AOI22_X1 U22647 ( .A1(n19653), .A2(n19664), .B1(n19698), .B2(n19663), .ZN(
        n19655) );
  AOI22_X1 U22648 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19667), .B1(
        n19699), .B2(n19666), .ZN(n19654) );
  OAI211_X1 U22649 ( .C1(n19656), .C2(n19732), .A(n19655), .B(n19654), .ZN(
        P2_U3163) );
  AOI22_X1 U22650 ( .A1(n19706), .A2(n19664), .B1(n19704), .B2(n19663), .ZN(
        n19658) );
  AOI22_X1 U22651 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19667), .B1(
        n19705), .B2(n19666), .ZN(n19657) );
  OAI211_X1 U22652 ( .C1(n19709), .C2(n19732), .A(n19658), .B(n19657), .ZN(
        P2_U3164) );
  AOI22_X1 U22653 ( .A1(n19711), .A2(n19664), .B1(n19238), .B2(n19663), .ZN(
        n19660) );
  AOI22_X1 U22654 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19667), .B1(
        n19710), .B2(n19666), .ZN(n19659) );
  OAI211_X1 U22655 ( .C1(n19714), .C2(n19732), .A(n19660), .B(n19659), .ZN(
        P2_U3165) );
  AOI22_X1 U22656 ( .A1(n19717), .A2(n19664), .B1(n19715), .B2(n19663), .ZN(
        n19662) );
  AOI22_X1 U22657 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19667), .B1(
        n19716), .B2(n19666), .ZN(n19661) );
  OAI211_X1 U22658 ( .C1(n19722), .C2(n19732), .A(n19662), .B(n19661), .ZN(
        P2_U3166) );
  AOI22_X1 U22659 ( .A1(n19665), .A2(n19664), .B1(n19723), .B2(n19663), .ZN(
        n19669) );
  AOI22_X1 U22660 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19667), .B1(
        n19725), .B2(n19666), .ZN(n19668) );
  OAI211_X1 U22661 ( .C1(n19670), .C2(n19732), .A(n19669), .B(n19668), .ZN(
        P2_U3167) );
  NAND2_X1 U22662 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19671), .ZN(
        n19678) );
  OR2_X1 U22663 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19678), .ZN(n19672) );
  NOR3_X1 U22664 ( .A1(n21051), .A2(n19724), .A3(n10692), .ZN(n19677) );
  AOI21_X1 U22665 ( .B1(n10692), .B2(n19672), .A(n19677), .ZN(n19726) );
  AOI22_X1 U22666 ( .A1(n19726), .A2(n19674), .B1(n19724), .B2(n19673), .ZN(
        n19684) );
  INV_X1 U22667 ( .A(n19815), .ZN(n19675) );
  NAND2_X1 U22668 ( .A1(n19676), .A2(n19675), .ZN(n19679) );
  AOI21_X1 U22669 ( .B1(n19679), .B2(n19678), .A(n19677), .ZN(n19681) );
  OAI211_X1 U22670 ( .C1(n19724), .C2(n19385), .A(n19681), .B(n19680), .ZN(
        n19729) );
  AOI22_X1 U22671 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19729), .B1(
        n19728), .B2(n19682), .ZN(n19683) );
  OAI211_X1 U22672 ( .C1(n19685), .C2(n19732), .A(n19684), .B(n19683), .ZN(
        P2_U3168) );
  AOI22_X1 U22673 ( .A1(n19726), .A2(n19687), .B1(n19724), .B2(n19686), .ZN(
        n19690) );
  AOI22_X1 U22674 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19729), .B1(
        n19728), .B2(n19688), .ZN(n19689) );
  OAI211_X1 U22675 ( .C1(n19691), .C2(n19732), .A(n19690), .B(n19689), .ZN(
        P2_U3169) );
  AOI22_X1 U22676 ( .A1(n19726), .A2(n19693), .B1(n19724), .B2(n19692), .ZN(
        n19696) );
  AOI22_X1 U22677 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19729), .B1(
        n19728), .B2(n19694), .ZN(n19695) );
  OAI211_X1 U22678 ( .C1(n19697), .C2(n19732), .A(n19696), .B(n19695), .ZN(
        P2_U3170) );
  AOI22_X1 U22679 ( .A1(n19726), .A2(n19699), .B1(n19724), .B2(n19698), .ZN(
        n19702) );
  AOI22_X1 U22680 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19729), .B1(
        n19728), .B2(n19700), .ZN(n19701) );
  OAI211_X1 U22681 ( .C1(n19703), .C2(n19732), .A(n19702), .B(n19701), .ZN(
        P2_U3171) );
  INV_X1 U22682 ( .A(n19728), .ZN(n19721) );
  AOI22_X1 U22683 ( .A1(n19726), .A2(n19705), .B1(n19724), .B2(n19704), .ZN(
        n19708) );
  AOI22_X1 U22684 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19729), .B1(
        n19718), .B2(n19706), .ZN(n19707) );
  OAI211_X1 U22685 ( .C1(n19709), .C2(n19721), .A(n19708), .B(n19707), .ZN(
        P2_U3172) );
  AOI22_X1 U22686 ( .A1(n19726), .A2(n19710), .B1(n19724), .B2(n19238), .ZN(
        n19713) );
  AOI22_X1 U22687 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19729), .B1(
        n19718), .B2(n19711), .ZN(n19712) );
  OAI211_X1 U22688 ( .C1(n19714), .C2(n19721), .A(n19713), .B(n19712), .ZN(
        P2_U3173) );
  AOI22_X1 U22689 ( .A1(n19726), .A2(n19716), .B1(n19724), .B2(n19715), .ZN(
        n19720) );
  AOI22_X1 U22690 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19729), .B1(
        n19718), .B2(n19717), .ZN(n19719) );
  OAI211_X1 U22691 ( .C1(n19722), .C2(n19721), .A(n19720), .B(n19719), .ZN(
        P2_U3174) );
  AOI22_X1 U22692 ( .A1(n19726), .A2(n19725), .B1(n19724), .B2(n19723), .ZN(
        n19731) );
  AOI22_X1 U22693 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19729), .B1(
        n19728), .B2(n19727), .ZN(n19730) );
  OAI211_X1 U22694 ( .C1(n19733), .C2(n19732), .A(n19731), .B(n19730), .ZN(
        P2_U3175) );
  AOI211_X1 U22695 ( .C1(n10692), .C2(n19865), .A(n19737), .B(n19734), .ZN(
        n19735) );
  INV_X1 U22696 ( .A(n19735), .ZN(n19740) );
  OAI211_X1 U22697 ( .C1(n19737), .C2(n19736), .A(n19865), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19739) );
  OAI211_X1 U22698 ( .C1(n19741), .C2(n19740), .A(n19739), .B(n19738), .ZN(
        P2_U3177) );
  AND2_X1 U22699 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19742), .ZN(
        P2_U3179) );
  AND2_X1 U22700 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19742), .ZN(
        P2_U3180) );
  AND2_X1 U22701 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19742), .ZN(
        P2_U3181) );
  AND2_X1 U22702 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19742), .ZN(
        P2_U3182) );
  AND2_X1 U22703 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19742), .ZN(
        P2_U3183) );
  AND2_X1 U22704 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19742), .ZN(
        P2_U3184) );
  AND2_X1 U22705 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19742), .ZN(
        P2_U3185) );
  AND2_X1 U22706 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19742), .ZN(
        P2_U3186) );
  AND2_X1 U22707 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19742), .ZN(
        P2_U3187) );
  AND2_X1 U22708 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19742), .ZN(
        P2_U3188) );
  NOR2_X1 U22709 ( .A1(n21026), .A2(n19808), .ZN(P2_U3189) );
  AND2_X1 U22710 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19742), .ZN(
        P2_U3190) );
  AND2_X1 U22711 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19742), .ZN(
        P2_U3191) );
  AND2_X1 U22712 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19742), .ZN(
        P2_U3192) );
  AND2_X1 U22713 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19742), .ZN(
        P2_U3193) );
  AND2_X1 U22714 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19742), .ZN(
        P2_U3194) );
  AND2_X1 U22715 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19742), .ZN(
        P2_U3195) );
  INV_X1 U22716 ( .A(P2_DATAWIDTH_REG_14__SCAN_IN), .ZN(n20880) );
  NOR2_X1 U22717 ( .A1(n20880), .A2(n19808), .ZN(P2_U3196) );
  AND2_X1 U22718 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19742), .ZN(
        P2_U3197) );
  AND2_X1 U22719 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19742), .ZN(
        P2_U3198) );
  AND2_X1 U22720 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19742), .ZN(
        P2_U3199) );
  AND2_X1 U22721 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19742), .ZN(
        P2_U3200) );
  AND2_X1 U22722 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19742), .ZN(P2_U3201) );
  AND2_X1 U22723 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19742), .ZN(P2_U3202) );
  AND2_X1 U22724 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19742), .ZN(P2_U3203) );
  AND2_X1 U22725 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19742), .ZN(P2_U3204) );
  NOR2_X1 U22726 ( .A1(n20925), .A2(n19808), .ZN(P2_U3205) );
  AND2_X1 U22727 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19742), .ZN(P2_U3206) );
  AND2_X1 U22728 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19742), .ZN(P2_U3207) );
  AND2_X1 U22729 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19742), .ZN(P2_U3208) );
  INV_X1 U22730 ( .A(NA), .ZN(n20650) );
  OAI21_X1 U22731 ( .B1(n20650), .B2(n19748), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19759) );
  INV_X1 U22732 ( .A(n19759), .ZN(n19746) );
  NOR2_X1 U22733 ( .A1(n19867), .A2(n19743), .ZN(n19753) );
  INV_X1 U22734 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19877) );
  NOR3_X1 U22735 ( .A1(n19753), .A2(n19877), .A3(n19747), .ZN(n19745) );
  OAI211_X1 U22736 ( .C1(HOLD), .C2(n19877), .A(n19880), .B(n19754), .ZN(
        n19744) );
  OAI21_X1 U22737 ( .B1(n19746), .B2(n19745), .A(n19744), .ZN(P2_U3209) );
  NOR2_X1 U22738 ( .A1(HOLD), .A2(n19747), .ZN(n19758) );
  AOI21_X1 U22739 ( .B1(n19760), .B2(n19748), .A(n19758), .ZN(n19751) );
  OAI22_X1 U22740 ( .A1(n19751), .A2(n19877), .B1(n19750), .B2(n19749), .ZN(
        n19752) );
  OR3_X1 U22741 ( .A1(n19871), .A2(n19753), .A3(n19752), .ZN(P2_U3210) );
  INV_X1 U22742 ( .A(n19753), .ZN(n19757) );
  OAI22_X1 U22743 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19754), .B1(NA), 
        .B2(n19757), .ZN(n19755) );
  OAI211_X1 U22744 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19755), .ZN(n19756) );
  OAI221_X1 U22745 ( .B1(n19759), .B2(n19758), .C1(n19759), .C2(n19757), .A(
        n19756), .ZN(P2_U3211) );
  INV_X2 U22746 ( .A(n19880), .ZN(n19879) );
  OAI222_X1 U22747 ( .A1(n19797), .A2(n14868), .B1(n19761), .B2(n19879), .C1(
        n10790), .C2(n19801), .ZN(P2_U3212) );
  OAI222_X1 U22748 ( .A1(n19797), .A2(n10790), .B1(n20803), .B2(n19879), .C1(
        n10803), .C2(n19801), .ZN(P2_U3213) );
  OAI222_X1 U22749 ( .A1(n19797), .A2(n10803), .B1(n19762), .B2(n19879), .C1(
        n10814), .C2(n19801), .ZN(P2_U3214) );
  OAI222_X1 U22750 ( .A1(n19801), .A2(n13974), .B1(n19763), .B2(n19879), .C1(
        n10814), .C2(n19797), .ZN(P2_U3215) );
  OAI222_X1 U22751 ( .A1(n19801), .A2(n19765), .B1(n19764), .B2(n19879), .C1(
        n13974), .C2(n19797), .ZN(P2_U3216) );
  OAI222_X1 U22752 ( .A1(n19801), .A2(n10824), .B1(n19766), .B2(n19879), .C1(
        n19765), .C2(n19797), .ZN(P2_U3217) );
  OAI222_X1 U22753 ( .A1(n19801), .A2(n10830), .B1(n19767), .B2(n19879), .C1(
        n10824), .C2(n19797), .ZN(P2_U3218) );
  OAI222_X1 U22754 ( .A1(n19801), .A2(n10836), .B1(n19768), .B2(n19879), .C1(
        n10830), .C2(n19797), .ZN(P2_U3219) );
  OAI222_X1 U22755 ( .A1(n19801), .A2(n10840), .B1(n20905), .B2(n19879), .C1(
        n10836), .C2(n19797), .ZN(P2_U3220) );
  OAI222_X1 U22756 ( .A1(n19801), .A2(n10843), .B1(n19769), .B2(n19879), .C1(
        n10840), .C2(n19797), .ZN(P2_U3221) );
  OAI222_X1 U22757 ( .A1(n19801), .A2(n10848), .B1(n19770), .B2(n19879), .C1(
        n10843), .C2(n19797), .ZN(P2_U3222) );
  OAI222_X1 U22758 ( .A1(n19801), .A2(n15187), .B1(n19771), .B2(n19879), .C1(
        n10848), .C2(n19797), .ZN(P2_U3223) );
  OAI222_X1 U22759 ( .A1(n19801), .A2(n10855), .B1(n19772), .B2(n19879), .C1(
        n15187), .C2(n19797), .ZN(P2_U3224) );
  OAI222_X1 U22760 ( .A1(n19801), .A2(n10863), .B1(n19773), .B2(n19879), .C1(
        n10855), .C2(n19797), .ZN(P2_U3225) );
  OAI222_X1 U22761 ( .A1(n19801), .A2(n19775), .B1(n19774), .B2(n19879), .C1(
        n10863), .C2(n19797), .ZN(P2_U3226) );
  OAI222_X1 U22762 ( .A1(n19801), .A2(n19777), .B1(n19776), .B2(n19879), .C1(
        n19775), .C2(n19797), .ZN(P2_U3227) );
  OAI222_X1 U22763 ( .A1(n19801), .A2(n10874), .B1(n19778), .B2(n19879), .C1(
        n19777), .C2(n19797), .ZN(P2_U3228) );
  OAI222_X1 U22764 ( .A1(n19801), .A2(n10877), .B1(n19779), .B2(n19879), .C1(
        n10874), .C2(n19797), .ZN(P2_U3229) );
  OAI222_X1 U22765 ( .A1(n19801), .A2(n10882), .B1(n19780), .B2(n19879), .C1(
        n10877), .C2(n19797), .ZN(P2_U3230) );
  OAI222_X1 U22766 ( .A1(n19801), .A2(n10886), .B1(n19781), .B2(n19879), .C1(
        n10882), .C2(n19797), .ZN(P2_U3231) );
  OAI222_X1 U22767 ( .A1(n19801), .A2(n19783), .B1(n19782), .B2(n19879), .C1(
        n10886), .C2(n19797), .ZN(P2_U3232) );
  OAI222_X1 U22768 ( .A1(n19801), .A2(n15102), .B1(n19784), .B2(n19879), .C1(
        n19783), .C2(n19797), .ZN(P2_U3233) );
  OAI222_X1 U22769 ( .A1(n19801), .A2(n19786), .B1(n19785), .B2(n19879), .C1(
        n15102), .C2(n19797), .ZN(P2_U3234) );
  OAI222_X1 U22770 ( .A1(n19801), .A2(n19788), .B1(n19787), .B2(n19879), .C1(
        n19786), .C2(n19797), .ZN(P2_U3235) );
  OAI222_X1 U22771 ( .A1(n19801), .A2(n10900), .B1(n19789), .B2(n19879), .C1(
        n19788), .C2(n19797), .ZN(P2_U3236) );
  OAI222_X1 U22772 ( .A1(n19801), .A2(n19792), .B1(n19790), .B2(n19879), .C1(
        n10900), .C2(n19797), .ZN(P2_U3237) );
  OAI222_X1 U22773 ( .A1(n19797), .A2(n19792), .B1(n19791), .B2(n19879), .C1(
        n19793), .C2(n19801), .ZN(P2_U3238) );
  OAI222_X1 U22774 ( .A1(n19801), .A2(n19795), .B1(n19794), .B2(n19879), .C1(
        n19793), .C2(n19797), .ZN(P2_U3239) );
  OAI222_X1 U22775 ( .A1(n19801), .A2(n19798), .B1(n19796), .B2(n19879), .C1(
        n19795), .C2(n19797), .ZN(P2_U3240) );
  INV_X1 U22776 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19800) );
  OAI222_X1 U22777 ( .A1(n19801), .A2(n19800), .B1(n19799), .B2(n19879), .C1(
        n19798), .C2(n19797), .ZN(P2_U3241) );
  OAI22_X1 U22778 ( .A1(n19880), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19879), .ZN(n19802) );
  INV_X1 U22779 ( .A(n19802), .ZN(P2_U3585) );
  MUX2_X1 U22780 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n19880), .Z(P2_U3586) );
  OAI22_X1 U22781 ( .A1(n19880), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19879), .ZN(n19803) );
  INV_X1 U22782 ( .A(n19803), .ZN(P2_U3587) );
  OAI22_X1 U22783 ( .A1(n19880), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19879), .ZN(n19804) );
  INV_X1 U22784 ( .A(n19804), .ZN(P2_U3588) );
  OAI21_X1 U22785 ( .B1(n19808), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19806), 
        .ZN(n19805) );
  INV_X1 U22786 ( .A(n19805), .ZN(P2_U3591) );
  OAI21_X1 U22787 ( .B1(n19808), .B2(n19807), .A(n19806), .ZN(P2_U3592) );
  OAI22_X1 U22788 ( .A1(n19818), .A2(n19810), .B1(n19816), .B2(n19809), .ZN(
        n19812) );
  OAI22_X1 U22789 ( .A1(n19813), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n19812), .B2(n19811), .ZN(n19814) );
  INV_X1 U22790 ( .A(n19814), .ZN(P2_U3596) );
  OAI21_X1 U22791 ( .B1(n19815), .B2(n19868), .A(n19820), .ZN(n19817) );
  NAND2_X1 U22792 ( .A1(n19817), .A2(n19816), .ZN(n19828) );
  INV_X1 U22793 ( .A(n19818), .ZN(n19822) );
  AOI222_X1 U22794 ( .A1(n19828), .A2(n19822), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19821), .C1(n19820), .C2(n19819), .ZN(n19823) );
  AOI22_X1 U22795 ( .A1(n19849), .A2(n19824), .B1(n19823), .B2(n19850), .ZN(
        P2_U3602) );
  INV_X1 U22796 ( .A(n19834), .ZN(n19826) );
  OAI21_X1 U22797 ( .B1(n19838), .B2(n19826), .A(n19825), .ZN(n19827) );
  AOI22_X1 U22798 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19829), .B1(n19828), 
        .B2(n19827), .ZN(n19830) );
  AOI22_X1 U22799 ( .A1(n19849), .A2(n12371), .B1(n19830), .B2(n19850), .ZN(
        P2_U3603) );
  INV_X1 U22800 ( .A(n19831), .ZN(n19832) );
  NAND2_X1 U22801 ( .A1(n19841), .A2(n19832), .ZN(n19837) );
  NAND2_X1 U22802 ( .A1(n19833), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19836) );
  NAND2_X1 U22803 ( .A1(n19838), .A2(n19834), .ZN(n19835) );
  OAI211_X1 U22804 ( .C1(n19838), .C2(n19837), .A(n19836), .B(n19835), .ZN(
        n19839) );
  INV_X1 U22805 ( .A(n19839), .ZN(n19840) );
  AOI22_X1 U22806 ( .A1(n19849), .A2(n10670), .B1(n19840), .B2(n19850), .ZN(
        P2_U3604) );
  INV_X1 U22807 ( .A(n19841), .ZN(n19845) );
  INV_X1 U22808 ( .A(n19842), .ZN(n19844) );
  OAI22_X1 U22809 ( .A1(n19846), .A2(n19845), .B1(n19844), .B2(n19843), .ZN(
        n19847) );
  AOI21_X1 U22810 ( .B1(n12376), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19847), 
        .ZN(n19848) );
  OAI22_X1 U22811 ( .A1(n12376), .A2(n19850), .B1(n19849), .B2(n19848), .ZN(
        P2_U3605) );
  INV_X1 U22812 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19851) );
  AOI22_X1 U22813 ( .A1(n19879), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19851), 
        .B2(n19880), .ZN(P2_U3608) );
  OAI22_X1 U22814 ( .A1(n19855), .A2(n19854), .B1(n19853), .B2(n19852), .ZN(
        n19856) );
  INV_X1 U22815 ( .A(n19856), .ZN(n19857) );
  NAND2_X1 U22816 ( .A1(n19858), .A2(n19857), .ZN(n19860) );
  MUX2_X1 U22817 ( .A(P2_MORE_REG_SCAN_IN), .B(n19860), .S(n19859), .Z(
        P2_U3609) );
  OAI21_X1 U22818 ( .B1(n19861), .B2(n10692), .A(n19385), .ZN(n19862) );
  OAI211_X1 U22819 ( .C1(n19865), .C2(n19864), .A(n19863), .B(n19862), .ZN(
        n19878) );
  AOI21_X1 U22820 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19867), .A(n19866), 
        .ZN(n19875) );
  NAND2_X1 U22821 ( .A1(n19869), .A2(n19868), .ZN(n19870) );
  NAND2_X1 U22822 ( .A1(n19871), .A2(n19870), .ZN(n19872) );
  AND3_X1 U22823 ( .A1(n19873), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n19872), 
        .ZN(n19874) );
  OAI21_X1 U22824 ( .B1(n19875), .B2(n19874), .A(n19878), .ZN(n19876) );
  OAI21_X1 U22825 ( .B1(n19878), .B2(n19877), .A(n19876), .ZN(P2_U3610) );
  OAI22_X1 U22826 ( .A1(n19880), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19879), .ZN(n19881) );
  INV_X1 U22827 ( .A(n19881), .ZN(P2_U3611) );
  INV_X1 U22828 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20655) );
  AOI21_X1 U22829 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n20658), .A(n20655), 
        .ZN(n19889) );
  INV_X1 U22830 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19882) );
  NAND2_X1 U22831 ( .A1(n20655), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20713) );
  AOI21_X1 U22832 ( .B1(n19889), .B2(n19882), .A(n20715), .ZN(P1_U2802) );
  NAND2_X1 U22833 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n19883), .ZN(n19887) );
  OAI21_X1 U22834 ( .B1(n19885), .B2(n19884), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19886) );
  OAI21_X1 U22835 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n19887), .A(n19886), 
        .ZN(P1_U2803) );
  NOR2_X1 U22836 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19890) );
  OAI21_X1 U22837 ( .B1(n19890), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20727), .ZN(
        n19888) );
  OAI21_X1 U22838 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20713), .A(n19888), 
        .ZN(P1_U2804) );
  NOR2_X1 U22839 ( .A1(n20715), .A2(n19889), .ZN(n20704) );
  OAI21_X1 U22840 ( .B1(BS16), .B2(n19890), .A(n20704), .ZN(n20702) );
  OAI21_X1 U22841 ( .B1(n20704), .B2(n20906), .A(n20702), .ZN(P1_U2805) );
  AOI21_X1 U22842 ( .B1(n19891), .B2(P1_FLUSH_REG_SCAN_IN), .A(n20064), .ZN(
        n19892) );
  INV_X1 U22843 ( .A(n19892), .ZN(P1_U2806) );
  NOR4_X1 U22844 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19896) );
  NOR4_X1 U22845 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_17__SCAN_IN), .A3(P1_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(n19895) );
  NOR4_X1 U22846 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19894) );
  NOR4_X1 U22847 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19893) );
  NAND4_X1 U22848 ( .A1(n19896), .A2(n19895), .A3(n19894), .A4(n19893), .ZN(
        n19902) );
  NOR4_X1 U22849 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_3__SCAN_IN), .A3(P1_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19900) );
  AOI211_X1 U22850 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_4__SCAN_IN), .B(
        P1_DATAWIDTH_REG_8__SCAN_IN), .ZN(n19899) );
  NOR4_X1 U22851 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_13__SCAN_IN), .A3(P1_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_15__SCAN_IN), .ZN(n19898) );
  NOR4_X1 U22852 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_9__SCAN_IN), .A3(P1_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_11__SCAN_IN), .ZN(n19897) );
  NAND4_X1 U22853 ( .A1(n19900), .A2(n19899), .A3(n19898), .A4(n19897), .ZN(
        n19901) );
  NOR2_X1 U22854 ( .A1(n19902), .A2(n19901), .ZN(n20709) );
  INV_X1 U22855 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19904) );
  NOR3_X1 U22856 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19905) );
  OAI21_X1 U22857 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19905), .A(n20709), .ZN(
        n19903) );
  OAI21_X1 U22858 ( .B1(n20709), .B2(n19904), .A(n19903), .ZN(P1_U2807) );
  INV_X1 U22859 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20703) );
  AOI21_X1 U22860 ( .B1(n20705), .B2(n20703), .A(n19905), .ZN(n19907) );
  INV_X1 U22861 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19906) );
  INV_X1 U22862 ( .A(n20709), .ZN(n20712) );
  AOI22_X1 U22863 ( .A1(n20709), .A2(n19907), .B1(n19906), .B2(n20712), .ZN(
        P1_U2808) );
  INV_X1 U22864 ( .A(n19908), .ZN(n19914) );
  NAND3_X1 U22865 ( .A1(n19982), .A2(n19915), .A3(n19909), .ZN(n19911) );
  AOI21_X1 U22866 ( .B1(n19991), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n19925), .ZN(n19910) );
  OAI211_X1 U22867 ( .C1(n19986), .C2(n19912), .A(n19911), .B(n19910), .ZN(
        n19913) );
  AOI21_X1 U22868 ( .B1(n19914), .B2(n19959), .A(n19913), .ZN(n19919) );
  INV_X1 U22869 ( .A(n19915), .ZN(n19916) );
  NAND2_X1 U22870 ( .A1(n19982), .A2(n19916), .ZN(n19930) );
  NAND2_X1 U22871 ( .A1(n19927), .A2(n19930), .ZN(n19922) );
  AOI22_X1 U22872 ( .A1(n19917), .A2(n19932), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n19922), .ZN(n19918) );
  OAI211_X1 U22873 ( .C1(n19920), .C2(n19965), .A(n19919), .B(n19918), .ZN(
        P1_U2833) );
  OAI22_X1 U22874 ( .A1(n20001), .A2(n19987), .B1(n20007), .B2(n19986), .ZN(
        n19921) );
  AOI21_X1 U22875 ( .B1(n19922), .B2(P1_REIP_REG_6__SCAN_IN), .A(n19921), .ZN(
        n19923) );
  INV_X1 U22876 ( .A(n19923), .ZN(n19924) );
  AOI211_X1 U22877 ( .C1(n19991), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n19925), .B(n19924), .ZN(n19934) );
  INV_X1 U22878 ( .A(n19937), .ZN(n19926) );
  AND2_X1 U22879 ( .A1(n19927), .A2(n19926), .ZN(n19928) );
  OR2_X1 U22880 ( .A1(n19929), .A2(n19928), .ZN(n19960) );
  NAND2_X1 U22881 ( .A1(n19960), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n19939) );
  NOR2_X1 U22882 ( .A1(n19939), .A2(n19930), .ZN(n19931) );
  AOI21_X1 U22883 ( .B1(n20005), .B2(n19932), .A(n19931), .ZN(n19933) );
  OAI211_X1 U22884 ( .C1(n19935), .C2(n19965), .A(n19934), .B(n19933), .ZN(
        P1_U2834) );
  OAI21_X1 U22885 ( .B1(n19969), .B2(n19937), .A(n19936), .ZN(n19938) );
  NAND2_X1 U22886 ( .A1(n19939), .A2(n19938), .ZN(n19946) );
  OAI22_X1 U22887 ( .A1(n19941), .A2(n19987), .B1(n19986), .B2(n19940), .ZN(
        n19942) );
  INV_X1 U22888 ( .A(n19942), .ZN(n19943) );
  NAND2_X1 U22889 ( .A1(n19953), .A2(n19943), .ZN(n19944) );
  AOI21_X1 U22890 ( .B1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n19991), .A(
        n19944), .ZN(n19945) );
  NAND2_X1 U22891 ( .A1(n19946), .A2(n19945), .ZN(n19947) );
  AOI21_X1 U22892 ( .B1(n19948), .B2(n19996), .A(n19947), .ZN(n19949) );
  OAI21_X1 U22893 ( .B1(n19950), .B2(n19965), .A(n19949), .ZN(P1_U2835) );
  NAND3_X1 U22894 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n19951) );
  NOR3_X1 U22895 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n19969), .A3(n19951), .ZN(
        n19958) );
  INV_X1 U22896 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19955) );
  AOI22_X1 U22897 ( .A1(n19952), .A2(n19983), .B1(n19971), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n19954) );
  OAI211_X1 U22898 ( .C1(n19956), .C2(n19955), .A(n19954), .B(n19953), .ZN(
        n19957) );
  AOI211_X1 U22899 ( .C1(n20069), .C2(n19959), .A(n19958), .B(n19957), .ZN(
        n19964) );
  INV_X1 U22900 ( .A(n19960), .ZN(n19961) );
  AOI22_X1 U22901 ( .A1(n19962), .A2(n19996), .B1(P1_REIP_REG_4__SCAN_IN), 
        .B2(n19961), .ZN(n19963) );
  OAI211_X1 U22902 ( .C1(n19966), .C2(n19965), .A(n19964), .B(n19963), .ZN(
        P1_U2836) );
  INV_X1 U22903 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n19981) );
  NAND2_X1 U22904 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_2__SCAN_IN), 
        .ZN(n19968) );
  AOI21_X1 U22905 ( .B1(n19982), .B2(n19968), .A(n19967), .ZN(n19999) );
  NAND2_X1 U22906 ( .A1(n20349), .A2(n19983), .ZN(n19973) );
  NOR3_X1 U22907 ( .A1(n19969), .A2(P1_REIP_REG_3__SCAN_IN), .A3(n19968), .ZN(
        n19970) );
  AOI21_X1 U22908 ( .B1(P1_EBX_REG_3__SCAN_IN), .B2(n19971), .A(n19970), .ZN(
        n19972) );
  OAI211_X1 U22909 ( .C1(n19974), .C2(n19987), .A(n19973), .B(n19972), .ZN(
        n19975) );
  AOI21_X1 U22910 ( .B1(n19991), .B2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n19975), .ZN(n19980) );
  INV_X1 U22911 ( .A(n19976), .ZN(n19977) );
  AOI22_X1 U22912 ( .A1(n19978), .A2(n19996), .B1(n19977), .B2(n19993), .ZN(
        n19979) );
  OAI211_X1 U22913 ( .C1(n19981), .C2(n19999), .A(n19980), .B(n19979), .ZN(
        P1_U2837) );
  AOI21_X1 U22914 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19982), .A(
        P1_REIP_REG_2__SCAN_IN), .ZN(n20000) );
  INV_X1 U22915 ( .A(n19983), .ZN(n19984) );
  NOR2_X1 U22916 ( .A1(n13425), .A2(n19984), .ZN(n19990) );
  OAI22_X1 U22917 ( .A1(n19988), .A2(n19987), .B1(n19986), .B2(n19985), .ZN(
        n19989) );
  AOI211_X1 U22918 ( .C1(n19991), .C2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n19990), .B(n19989), .ZN(n19998) );
  INV_X1 U22919 ( .A(n19992), .ZN(n19994) );
  AOI22_X1 U22920 ( .A1(n19996), .A2(n19995), .B1(n19994), .B2(n19993), .ZN(
        n19997) );
  OAI211_X1 U22921 ( .C1(n20000), .C2(n19999), .A(n19998), .B(n19997), .ZN(
        P1_U2838) );
  NOR2_X1 U22922 ( .A1(n20002), .A2(n20001), .ZN(n20003) );
  AOI21_X1 U22923 ( .B1(n20005), .B2(n20004), .A(n20003), .ZN(n20006) );
  OAI21_X1 U22924 ( .B1(n14350), .B2(n20007), .A(n20006), .ZN(P1_U2866) );
  INV_X1 U22925 ( .A(P1_UWORD_REG_1__SCAN_IN), .ZN(n20751) );
  INV_X1 U22926 ( .A(n20008), .ZN(n20010) );
  AOI22_X1 U22927 ( .A1(n20033), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n20010), 
        .B2(P1_EAX_REG_17__SCAN_IN), .ZN(n20009) );
  OAI21_X1 U22928 ( .B1(n20751), .B2(n20013), .A(n20009), .ZN(P1_U2919) );
  INV_X1 U22929 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n20951) );
  AOI22_X1 U22930 ( .A1(n20010), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20719), .ZN(n20011) );
  OAI21_X1 U22931 ( .B1(n20951), .B2(n20017), .A(n20011), .ZN(P1_U2920) );
  AOI22_X1 U22932 ( .A1(P1_EAX_REG_15__SCAN_IN), .A2(n20023), .B1(n20033), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20012) );
  OAI21_X1 U22933 ( .B1(n20014), .B2(n20013), .A(n20012), .ZN(P1_U2921) );
  AOI22_X1 U22934 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20015) );
  OAI21_X1 U22935 ( .B1(n14056), .B2(n20035), .A(n20015), .ZN(P1_U2922) );
  AOI22_X1 U22936 ( .A1(P1_EAX_REG_13__SCAN_IN), .A2(n20023), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20719), .ZN(n20016) );
  OAI21_X1 U22937 ( .B1(n20965), .B2(n20017), .A(n20016), .ZN(P1_U2923) );
  INV_X1 U22938 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20019) );
  AOI22_X1 U22939 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20018) );
  OAI21_X1 U22940 ( .B1(n20019), .B2(n20035), .A(n20018), .ZN(P1_U2924) );
  AOI22_X1 U22941 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20020) );
  OAI21_X1 U22942 ( .B1(n14047), .B2(n20035), .A(n20020), .ZN(P1_U2925) );
  AOI22_X1 U22943 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20021) );
  OAI21_X1 U22944 ( .B1(n13998), .B2(n20035), .A(n20021), .ZN(P1_U2926) );
  AOI22_X1 U22945 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20022) );
  OAI21_X1 U22946 ( .B1(n13937), .B2(n20035), .A(n20022), .ZN(P1_U2927) );
  AOI222_X1 U22947 ( .A1(n20719), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n20023), 
        .B2(P1_EAX_REG_8__SCAN_IN), .C1(P1_DATAO_REG_8__SCAN_IN), .C2(n20033), 
        .ZN(n20024) );
  INV_X1 U22948 ( .A(n20024), .ZN(P1_U2928) );
  AOI22_X1 U22949 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20025) );
  OAI21_X1 U22950 ( .B1(n13822), .B2(n20035), .A(n20025), .ZN(P1_U2929) );
  AOI22_X1 U22951 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20026) );
  OAI21_X1 U22952 ( .B1(n11399), .B2(n20035), .A(n20026), .ZN(P1_U2930) );
  AOI22_X1 U22953 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20027) );
  OAI21_X1 U22954 ( .B1(n13696), .B2(n20035), .A(n20027), .ZN(P1_U2931) );
  AOI22_X1 U22955 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20028) );
  OAI21_X1 U22956 ( .B1(n20029), .B2(n20035), .A(n20028), .ZN(P1_U2932) );
  AOI22_X1 U22957 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20030) );
  OAI21_X1 U22958 ( .B1(n11373), .B2(n20035), .A(n20030), .ZN(P1_U2933) );
  AOI22_X1 U22959 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20031) );
  OAI21_X1 U22960 ( .B1(n13580), .B2(n20035), .A(n20031), .ZN(P1_U2934) );
  AOI22_X1 U22961 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20032) );
  OAI21_X1 U22962 ( .B1(n11362), .B2(n20035), .A(n20032), .ZN(P1_U2935) );
  AOI22_X1 U22963 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20719), .B1(n20033), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20034) );
  OAI21_X1 U22964 ( .B1(n11353), .B2(n20035), .A(n20034), .ZN(P1_U2936) );
  AOI22_X1 U22965 ( .A1(n20056), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20055), .ZN(n20037) );
  NAND2_X1 U22966 ( .A1(n20043), .A2(n20036), .ZN(n20045) );
  NAND2_X1 U22967 ( .A1(n20037), .A2(n20045), .ZN(P1_U2946) );
  AOI22_X1 U22968 ( .A1(n20056), .A2(P1_EAX_REG_26__SCAN_IN), .B1(n20055), 
        .B2(P1_UWORD_REG_10__SCAN_IN), .ZN(n20039) );
  NAND2_X1 U22969 ( .A1(n20043), .A2(n20038), .ZN(n20047) );
  NAND2_X1 U22970 ( .A1(n20039), .A2(n20047), .ZN(P1_U2947) );
  AOI22_X1 U22971 ( .A1(n20056), .A2(P1_EAX_REG_27__SCAN_IN), .B1(n20055), 
        .B2(P1_UWORD_REG_11__SCAN_IN), .ZN(n20041) );
  NAND2_X1 U22972 ( .A1(n20043), .A2(n20040), .ZN(n20049) );
  NAND2_X1 U22973 ( .A1(n20041), .A2(n20049), .ZN(P1_U2948) );
  AOI22_X1 U22974 ( .A1(n20056), .A2(P1_EAX_REG_29__SCAN_IN), .B1(n20055), 
        .B2(P1_UWORD_REG_13__SCAN_IN), .ZN(n20044) );
  NAND2_X1 U22975 ( .A1(n20043), .A2(n20042), .ZN(n20053) );
  NAND2_X1 U22976 ( .A1(n20044), .A2(n20053), .ZN(P1_U2950) );
  AOI22_X1 U22977 ( .A1(n20056), .A2(P1_EAX_REG_9__SCAN_IN), .B1(n20055), .B2(
        P1_LWORD_REG_9__SCAN_IN), .ZN(n20046) );
  NAND2_X1 U22978 ( .A1(n20046), .A2(n20045), .ZN(P1_U2961) );
  AOI22_X1 U22979 ( .A1(n20056), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n20055), 
        .B2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20048) );
  NAND2_X1 U22980 ( .A1(n20048), .A2(n20047), .ZN(P1_U2962) );
  AOI22_X1 U22981 ( .A1(n20056), .A2(P1_EAX_REG_11__SCAN_IN), .B1(n20055), 
        .B2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20050) );
  NAND2_X1 U22982 ( .A1(n20050), .A2(n20049), .ZN(P1_U2963) );
  AOI22_X1 U22983 ( .A1(n20056), .A2(P1_EAX_REG_12__SCAN_IN), .B1(n20055), 
        .B2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20052) );
  NAND2_X1 U22984 ( .A1(n20052), .A2(n20051), .ZN(P1_U2964) );
  AOI22_X1 U22985 ( .A1(n20056), .A2(P1_EAX_REG_13__SCAN_IN), .B1(n20055), 
        .B2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20054) );
  NAND2_X1 U22986 ( .A1(n20054), .A2(n20053), .ZN(P1_U2965) );
  AOI22_X1 U22987 ( .A1(n20056), .A2(P1_EAX_REG_14__SCAN_IN), .B1(n20055), 
        .B2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20058) );
  NAND2_X1 U22988 ( .A1(n20058), .A2(n20057), .ZN(P1_U2966) );
  OR2_X1 U22989 ( .A1(n20060), .A2(n20059), .ZN(n20065) );
  OR2_X1 U22990 ( .A1(n20061), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n20062) );
  AND2_X1 U22991 ( .A1(n20063), .A2(n20062), .ZN(n20081) );
  AOI22_X1 U22992 ( .A1(n20065), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n20064), .B2(n20081), .ZN(n20067) );
  OR2_X1 U22993 ( .A1(n20066), .A2(n20711), .ZN(n20086) );
  OAI211_X1 U22994 ( .C1(n20068), .C2(n20106), .A(n20067), .B(n20086), .ZN(
        P1_U2999) );
  NAND2_X1 U22995 ( .A1(n20070), .A2(n20069), .ZN(n20071) );
  OAI211_X1 U22996 ( .C1(n20074), .C2(n20073), .A(n20072), .B(n20071), .ZN(
        n20075) );
  AOI21_X1 U22997 ( .B1(n20076), .B2(n20082), .A(n20075), .ZN(n20080) );
  OAI211_X1 U22998 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20078), .B(n20077), .ZN(n20079) );
  NAND2_X1 U22999 ( .A1(n20080), .A2(n20079), .ZN(P1_U3027) );
  NAND2_X1 U23000 ( .A1(n20082), .A2(n20081), .ZN(n20089) );
  INV_X1 U23001 ( .A(n20083), .ZN(n20084) );
  NAND2_X1 U23002 ( .A1(n20085), .A2(n20084), .ZN(n20087) );
  AND4_X1 U23003 ( .A1(n20089), .A2(n20088), .A3(n20087), .A4(n20086), .ZN(
        n20090) );
  OAI221_X1 U23004 ( .B1(n20093), .B2(n20092), .C1(n20093), .C2(n20091), .A(
        n20090), .ZN(P1_U3031) );
  AND2_X1 U23005 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n20094), .ZN(
        P1_U3032) );
  NAND2_X1 U23006 ( .A1(n20096), .A2(n20095), .ZN(n20217) );
  NAND2_X1 U23007 ( .A1(n20182), .A2(n13363), .ZN(n20488) );
  NAND2_X1 U23008 ( .A1(n20180), .A2(n20547), .ZN(n20099) );
  NAND2_X1 U23009 ( .A1(n13664), .A2(n20097), .ZN(n20585) );
  INV_X1 U23010 ( .A(n20585), .ZN(n20098) );
  NAND2_X1 U23011 ( .A1(n20547), .A2(n20906), .ZN(n20408) );
  OAI21_X1 U23012 ( .B1(n20099), .B2(n20634), .A(n20408), .ZN(n20114) );
  INV_X1 U23013 ( .A(n13425), .ZN(n20100) );
  OR2_X1 U23014 ( .A1(n20349), .A2(n20100), .ZN(n20185) );
  NOR2_X1 U23015 ( .A1(n20185), .A2(n20553), .ZN(n20111) );
  INV_X1 U23016 ( .A(n20411), .ZN(n20102) );
  INV_X1 U23017 ( .A(n20101), .ZN(n20350) );
  NOR2_X1 U23018 ( .A1(n20102), .A2(n20350), .ZN(n20243) );
  NOR2_X1 U23019 ( .A1(n20109), .A2(n20579), .ZN(n20413) );
  AOI22_X1 U23020 ( .A1(n20114), .A2(n20111), .B1(n20243), .B2(n20413), .ZN(
        n20156) );
  INV_X1 U23021 ( .A(n20584), .ZN(n20424) );
  NOR2_X2 U23022 ( .A1(n20149), .A2(n11249), .ZN(n20583) );
  NOR3_X1 U23023 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20160) );
  NAND2_X1 U23024 ( .A1(n20517), .A2(n20160), .ZN(n20112) );
  INV_X1 U23025 ( .A(n20112), .ZN(n20150) );
  NOR2_X2 U23026 ( .A1(n20106), .A2(n20105), .ZN(n20151) );
  AOI22_X1 U23027 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20151), .B1(DATAI_24_), 
        .B2(n20108), .ZN(n20593) );
  INV_X1 U23028 ( .A(n20593), .ZN(n20415) );
  AOI22_X1 U23029 ( .A1(n20583), .A2(n20150), .B1(n20634), .B2(n20415), .ZN(
        n20118) );
  INV_X1 U23030 ( .A(n20109), .ZN(n20110) );
  NOR2_X1 U23031 ( .A1(n20110), .A2(n20579), .ZN(n20299) );
  INV_X1 U23032 ( .A(n20111), .ZN(n20113) );
  AOI22_X1 U23033 ( .A1(n20114), .A2(n20113), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20112), .ZN(n20115) );
  OAI211_X1 U23034 ( .C1(n20243), .C2(n20640), .A(n20421), .B(n20115), .ZN(
        n20153) );
  AOI22_X1 U23035 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20151), .B1(DATAI_16_), 
        .B2(n20108), .ZN(n20116) );
  INV_X1 U23036 ( .A(n20116), .ZN(n20590) );
  AOI22_X1 U23037 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20153), .B1(
        n20152), .B2(n20590), .ZN(n20117) );
  OAI211_X1 U23038 ( .C1(n20156), .C2(n20424), .A(n20118), .B(n20117), .ZN(
        P1_U3033) );
  INV_X1 U23039 ( .A(n20595), .ZN(n20428) );
  NOR2_X2 U23040 ( .A1(n20149), .A2(n20120), .ZN(n20594) );
  INV_X1 U23041 ( .A(n20599), .ZN(n20425) );
  AOI22_X1 U23042 ( .A1(n20594), .A2(n20150), .B1(n20634), .B2(n20425), .ZN(
        n20123) );
  AOI22_X1 U23043 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20151), .B1(DATAI_17_), 
        .B2(n20108), .ZN(n20121) );
  INV_X1 U23044 ( .A(n20121), .ZN(n20596) );
  AOI22_X1 U23045 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20153), .B1(
        n20152), .B2(n20596), .ZN(n20122) );
  OAI211_X1 U23046 ( .C1(n20156), .C2(n20428), .A(n20123), .B(n20122), .ZN(
        P1_U3034) );
  INV_X1 U23047 ( .A(n20601), .ZN(n20432) );
  NOR2_X2 U23048 ( .A1(n20149), .A2(n20125), .ZN(n20600) );
  INV_X1 U23049 ( .A(n20605), .ZN(n20429) );
  AOI22_X1 U23050 ( .A1(n20600), .A2(n20150), .B1(n20634), .B2(n20429), .ZN(
        n20128) );
  AOI22_X1 U23051 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20151), .B1(DATAI_18_), 
        .B2(n20108), .ZN(n20126) );
  INV_X1 U23052 ( .A(n20126), .ZN(n20602) );
  AOI22_X1 U23053 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20153), .B1(
        n20152), .B2(n20602), .ZN(n20127) );
  OAI211_X1 U23054 ( .C1(n20156), .C2(n20432), .A(n20128), .B(n20127), .ZN(
        P1_U3035) );
  INV_X1 U23055 ( .A(n20607), .ZN(n20436) );
  NOR2_X2 U23056 ( .A1(n20149), .A2(n20130), .ZN(n20606) );
  INV_X1 U23057 ( .A(n20611), .ZN(n20433) );
  AOI22_X1 U23058 ( .A1(n20606), .A2(n20150), .B1(n20634), .B2(n20433), .ZN(
        n20133) );
  AOI22_X1 U23059 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20151), .B1(DATAI_19_), 
        .B2(n20108), .ZN(n20131) );
  INV_X1 U23060 ( .A(n20131), .ZN(n20608) );
  AOI22_X1 U23061 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20153), .B1(
        n20152), .B2(n20608), .ZN(n20132) );
  OAI211_X1 U23062 ( .C1(n20156), .C2(n20436), .A(n20133), .B(n20132), .ZN(
        P1_U3036) );
  INV_X1 U23063 ( .A(n20613), .ZN(n20440) );
  NOR2_X2 U23064 ( .A1(n20149), .A2(n11222), .ZN(n20612) );
  INV_X1 U23065 ( .A(n20617), .ZN(n20437) );
  AOI22_X1 U23066 ( .A1(n20612), .A2(n20150), .B1(n20634), .B2(n20437), .ZN(
        n20137) );
  AOI22_X1 U23067 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20151), .B1(DATAI_20_), 
        .B2(n20108), .ZN(n20135) );
  INV_X1 U23068 ( .A(n20135), .ZN(n20614) );
  AOI22_X1 U23069 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20153), .B1(
        n20152), .B2(n20614), .ZN(n20136) );
  OAI211_X1 U23070 ( .C1(n20156), .C2(n20440), .A(n20137), .B(n20136), .ZN(
        P1_U3037) );
  INV_X1 U23071 ( .A(n20619), .ZN(n20444) );
  NOR2_X2 U23072 ( .A1(n20149), .A2(n20139), .ZN(n20618) );
  INV_X1 U23073 ( .A(n20623), .ZN(n20441) );
  AOI22_X1 U23074 ( .A1(n20618), .A2(n20150), .B1(n20634), .B2(n20441), .ZN(
        n20142) );
  AOI22_X1 U23075 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20151), .B1(DATAI_21_), 
        .B2(n20108), .ZN(n20140) );
  INV_X1 U23076 ( .A(n20140), .ZN(n20620) );
  AOI22_X1 U23077 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20153), .B1(
        n20152), .B2(n20620), .ZN(n20141) );
  OAI211_X1 U23078 ( .C1(n20156), .C2(n20444), .A(n20142), .B(n20141), .ZN(
        P1_U3038) );
  INV_X1 U23079 ( .A(n20625), .ZN(n20448) );
  NOR2_X2 U23080 ( .A1(n20149), .A2(n11180), .ZN(n20624) );
  INV_X1 U23081 ( .A(n20629), .ZN(n20445) );
  AOI22_X1 U23082 ( .A1(n20624), .A2(n20150), .B1(n20634), .B2(n20445), .ZN(
        n20146) );
  AOI22_X1 U23083 ( .A1(DATAI_22_), .A2(n20108), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n20151), .ZN(n20144) );
  INV_X1 U23084 ( .A(n20144), .ZN(n20626) );
  AOI22_X1 U23085 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20153), .B1(
        n20152), .B2(n20626), .ZN(n20145) );
  OAI211_X1 U23086 ( .C1(n20156), .C2(n20448), .A(n20146), .B(n20145), .ZN(
        P1_U3039) );
  INV_X1 U23087 ( .A(n20632), .ZN(n20735) );
  NOR2_X2 U23088 ( .A1(n20149), .A2(n20148), .ZN(n20728) );
  AOI22_X1 U23089 ( .A1(DATAI_31_), .A2(n20108), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20151), .ZN(n20734) );
  INV_X1 U23090 ( .A(n20734), .ZN(n20542) );
  AOI22_X1 U23091 ( .A1(n20728), .A2(n20150), .B1(n20634), .B2(n20542), .ZN(
        n20155) );
  AOI22_X1 U23092 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20151), .B1(DATAI_23_), 
        .B2(n20108), .ZN(n20730) );
  INV_X1 U23093 ( .A(n20730), .ZN(n20633) );
  AOI22_X1 U23094 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20153), .B1(
        n20152), .B2(n20633), .ZN(n20154) );
  OAI211_X1 U23095 ( .C1(n20156), .C2(n20735), .A(n20155), .B(n20154), .ZN(
        P1_U3040) );
  INV_X1 U23096 ( .A(n20185), .ZN(n20213) );
  INV_X1 U23097 ( .A(n20377), .ZN(n20518) );
  INV_X1 U23098 ( .A(n20160), .ZN(n20157) );
  NOR2_X1 U23099 ( .A1(n20517), .A2(n20157), .ZN(n20175) );
  AOI21_X1 U23100 ( .B1(n20213), .B2(n20518), .A(n20175), .ZN(n20158) );
  OAI22_X1 U23101 ( .A1(n20158), .A2(n20581), .B1(n20157), .B2(n20579), .ZN(
        n20176) );
  AOI22_X1 U23102 ( .A1(n20584), .A2(n20176), .B1(n20583), .B2(n20175), .ZN(
        n20162) );
  OAI21_X1 U23103 ( .B1(n20217), .B2(n20906), .A(n20158), .ZN(n20159) );
  OAI221_X1 U23104 ( .B1(n20547), .B2(n20160), .C1(n20581), .C2(n20159), .A(
        n20587), .ZN(n20177) );
  OR2_X1 U23105 ( .A1(n20217), .A2(n20523), .ZN(n20183) );
  AOI22_X1 U23106 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20177), .B1(
        n20207), .B2(n20590), .ZN(n20161) );
  OAI211_X1 U23107 ( .C1(n20593), .C2(n20180), .A(n20162), .B(n20161), .ZN(
        P1_U3041) );
  AOI22_X1 U23108 ( .A1(n20595), .A2(n20176), .B1(n20594), .B2(n20175), .ZN(
        n20164) );
  AOI22_X1 U23109 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20177), .B1(
        n20207), .B2(n20596), .ZN(n20163) );
  OAI211_X1 U23110 ( .C1(n20599), .C2(n20180), .A(n20164), .B(n20163), .ZN(
        P1_U3042) );
  AOI22_X1 U23111 ( .A1(n20601), .A2(n20176), .B1(n20600), .B2(n20175), .ZN(
        n20166) );
  AOI22_X1 U23112 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20177), .B1(
        n20207), .B2(n20602), .ZN(n20165) );
  OAI211_X1 U23113 ( .C1(n20605), .C2(n20180), .A(n20166), .B(n20165), .ZN(
        P1_U3043) );
  AOI22_X1 U23114 ( .A1(n20607), .A2(n20176), .B1(n20606), .B2(n20175), .ZN(
        n20168) );
  AOI22_X1 U23115 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20177), .B1(
        n20207), .B2(n20608), .ZN(n20167) );
  OAI211_X1 U23116 ( .C1(n20611), .C2(n20180), .A(n20168), .B(n20167), .ZN(
        P1_U3044) );
  AOI22_X1 U23117 ( .A1(n20613), .A2(n20176), .B1(n20612), .B2(n20175), .ZN(
        n20170) );
  AOI22_X1 U23118 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20177), .B1(
        n20207), .B2(n20614), .ZN(n20169) );
  OAI211_X1 U23119 ( .C1(n20617), .C2(n20180), .A(n20170), .B(n20169), .ZN(
        P1_U3045) );
  AOI22_X1 U23120 ( .A1(n20619), .A2(n20176), .B1(n20618), .B2(n20175), .ZN(
        n20172) );
  AOI22_X1 U23121 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20177), .B1(
        n20207), .B2(n20620), .ZN(n20171) );
  OAI211_X1 U23122 ( .C1(n20623), .C2(n20180), .A(n20172), .B(n20171), .ZN(
        P1_U3046) );
  AOI22_X1 U23123 ( .A1(n20625), .A2(n20176), .B1(n20624), .B2(n20175), .ZN(
        n20174) );
  AOI22_X1 U23124 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20177), .B1(
        n20207), .B2(n20626), .ZN(n20173) );
  OAI211_X1 U23125 ( .C1(n20629), .C2(n20180), .A(n20174), .B(n20173), .ZN(
        P1_U3047) );
  AOI22_X1 U23126 ( .A1(n20632), .A2(n20176), .B1(n20728), .B2(n20175), .ZN(
        n20179) );
  AOI22_X1 U23127 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20177), .B1(
        n20207), .B2(n20633), .ZN(n20178) );
  OAI211_X1 U23128 ( .C1(n20734), .C2(n20180), .A(n20179), .B(n20178), .ZN(
        P1_U3048) );
  INV_X1 U23129 ( .A(n20406), .ZN(n20551) );
  OR2_X1 U23130 ( .A1(n20217), .A2(n20551), .ZN(n20191) );
  NAND3_X1 U23131 ( .A1(n20191), .A2(n20183), .A3(n20547), .ZN(n20184) );
  NAND2_X1 U23132 ( .A1(n20184), .A2(n20408), .ZN(n20189) );
  NOR2_X1 U23133 ( .A1(n20185), .A2(n13669), .ZN(n20186) );
  NOR2_X1 U23134 ( .A1(n20411), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20300) );
  AOI22_X1 U23135 ( .A1(n20189), .A2(n20186), .B1(n20413), .B2(n20300), .ZN(
        n20211) );
  NOR3_X1 U23136 ( .A1(n20414), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20218) );
  NAND2_X1 U23137 ( .A1(n20517), .A2(n20218), .ZN(n20187) );
  INV_X1 U23138 ( .A(n20187), .ZN(n20206) );
  AOI22_X1 U23139 ( .A1(n20207), .A2(n20415), .B1(n20583), .B2(n20206), .ZN(
        n20193) );
  INV_X1 U23140 ( .A(n20186), .ZN(n20188) );
  AOI22_X1 U23141 ( .A1(n20189), .A2(n20188), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20187), .ZN(n20190) );
  OAI21_X1 U23142 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20411), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20304) );
  NAND3_X1 U23143 ( .A1(n20421), .A2(n20190), .A3(n20304), .ZN(n20208) );
  AOI22_X1 U23144 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20208), .B1(
        n20237), .B2(n20590), .ZN(n20192) );
  OAI211_X1 U23145 ( .C1(n20211), .C2(n20424), .A(n20193), .B(n20192), .ZN(
        P1_U3049) );
  AOI22_X1 U23146 ( .A1(n20237), .A2(n20596), .B1(n20594), .B2(n20206), .ZN(
        n20195) );
  AOI22_X1 U23147 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20208), .B1(
        n20207), .B2(n20425), .ZN(n20194) );
  OAI211_X1 U23148 ( .C1(n20211), .C2(n20428), .A(n20195), .B(n20194), .ZN(
        P1_U3050) );
  AOI22_X1 U23149 ( .A1(n20237), .A2(n20602), .B1(n20600), .B2(n20206), .ZN(
        n20197) );
  AOI22_X1 U23150 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20208), .B1(
        n20207), .B2(n20429), .ZN(n20196) );
  OAI211_X1 U23151 ( .C1(n20211), .C2(n20432), .A(n20197), .B(n20196), .ZN(
        P1_U3051) );
  AOI22_X1 U23152 ( .A1(n20207), .A2(n20433), .B1(n20606), .B2(n20206), .ZN(
        n20199) );
  AOI22_X1 U23153 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20208), .B1(
        n20237), .B2(n20608), .ZN(n20198) );
  OAI211_X1 U23154 ( .C1(n20211), .C2(n20436), .A(n20199), .B(n20198), .ZN(
        P1_U3052) );
  AOI22_X1 U23155 ( .A1(n20207), .A2(n20437), .B1(n20612), .B2(n20206), .ZN(
        n20201) );
  AOI22_X1 U23156 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20208), .B1(
        n20237), .B2(n20614), .ZN(n20200) );
  OAI211_X1 U23157 ( .C1(n20211), .C2(n20440), .A(n20201), .B(n20200), .ZN(
        P1_U3053) );
  AOI22_X1 U23158 ( .A1(n20237), .A2(n20620), .B1(n20618), .B2(n20206), .ZN(
        n20203) );
  AOI22_X1 U23159 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20208), .B1(
        n20207), .B2(n20441), .ZN(n20202) );
  OAI211_X1 U23160 ( .C1(n20211), .C2(n20444), .A(n20203), .B(n20202), .ZN(
        P1_U3054) );
  AOI22_X1 U23161 ( .A1(n20237), .A2(n20626), .B1(n20624), .B2(n20206), .ZN(
        n20205) );
  AOI22_X1 U23162 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20208), .B1(
        n20207), .B2(n20445), .ZN(n20204) );
  OAI211_X1 U23163 ( .C1(n20211), .C2(n20448), .A(n20205), .B(n20204), .ZN(
        P1_U3055) );
  AOI22_X1 U23164 ( .A1(n20207), .A2(n20542), .B1(n20728), .B2(n20206), .ZN(
        n20210) );
  AOI22_X1 U23165 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20208), .B1(
        n20237), .B2(n20633), .ZN(n20209) );
  OAI211_X1 U23166 ( .C1(n20211), .C2(n20735), .A(n20210), .B(n20209), .ZN(
        P1_U3056) );
  AOI21_X1 U23167 ( .B1(n20213), .B2(n9837), .A(n10149), .ZN(n20220) );
  INV_X1 U23168 ( .A(n20220), .ZN(n20215) );
  INV_X1 U23169 ( .A(n20217), .ZN(n20214) );
  AOI21_X1 U23170 ( .B1(n20214), .B2(n20459), .A(n20581), .ZN(n20221) );
  AOI22_X1 U23171 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20218), .B1(n20215), 
        .B2(n20221), .ZN(n20242) );
  INV_X1 U23172 ( .A(n20463), .ZN(n20216) );
  AOI22_X1 U23173 ( .A1(n20238), .A2(n20590), .B1(n20583), .B2(n10149), .ZN(
        n20224) );
  OAI21_X1 U23174 ( .B1(n20547), .B2(n20218), .A(n20587), .ZN(n20219) );
  AOI21_X1 U23175 ( .B1(n20221), .B2(n20220), .A(n20219), .ZN(n20222) );
  AOI22_X1 U23176 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20239), .B1(
        n20237), .B2(n20415), .ZN(n20223) );
  OAI211_X1 U23177 ( .C1(n20242), .C2(n20424), .A(n20224), .B(n20223), .ZN(
        P1_U3057) );
  AOI22_X1 U23178 ( .A1(n20237), .A2(n20425), .B1(n20594), .B2(n10149), .ZN(
        n20226) );
  AOI22_X1 U23179 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20239), .B1(
        n20238), .B2(n20596), .ZN(n20225) );
  OAI211_X1 U23180 ( .C1(n20242), .C2(n20428), .A(n20226), .B(n20225), .ZN(
        P1_U3058) );
  AOI22_X1 U23181 ( .A1(n20238), .A2(n20602), .B1(n20600), .B2(n10149), .ZN(
        n20228) );
  AOI22_X1 U23182 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20239), .B1(
        n20237), .B2(n20429), .ZN(n20227) );
  OAI211_X1 U23183 ( .C1(n20242), .C2(n20432), .A(n20228), .B(n20227), .ZN(
        P1_U3059) );
  AOI22_X1 U23184 ( .A1(n20238), .A2(n20608), .B1(n20606), .B2(n10149), .ZN(
        n20230) );
  AOI22_X1 U23185 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20239), .B1(
        n20237), .B2(n20433), .ZN(n20229) );
  OAI211_X1 U23186 ( .C1(n20242), .C2(n20436), .A(n20230), .B(n20229), .ZN(
        P1_U3060) );
  AOI22_X1 U23187 ( .A1(n20238), .A2(n20614), .B1(n20612), .B2(n10149), .ZN(
        n20232) );
  AOI22_X1 U23188 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20239), .B1(
        n20237), .B2(n20437), .ZN(n20231) );
  OAI211_X1 U23189 ( .C1(n20242), .C2(n20440), .A(n20232), .B(n20231), .ZN(
        P1_U3061) );
  AOI22_X1 U23190 ( .A1(n20238), .A2(n20620), .B1(n20618), .B2(n10149), .ZN(
        n20234) );
  AOI22_X1 U23191 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20239), .B1(
        n20237), .B2(n20441), .ZN(n20233) );
  OAI211_X1 U23192 ( .C1(n20242), .C2(n20444), .A(n20234), .B(n20233), .ZN(
        P1_U3062) );
  AOI22_X1 U23193 ( .A1(n20238), .A2(n20626), .B1(n20624), .B2(n10149), .ZN(
        n20236) );
  AOI22_X1 U23194 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20239), .B1(
        n20237), .B2(n20445), .ZN(n20235) );
  OAI211_X1 U23195 ( .C1(n20242), .C2(n20448), .A(n20236), .B(n20235), .ZN(
        P1_U3063) );
  AOI22_X1 U23196 ( .A1(n20237), .A2(n20542), .B1(n20728), .B2(n10149), .ZN(
        n20241) );
  AOI22_X1 U23197 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20239), .B1(
        n20238), .B2(n20633), .ZN(n20240) );
  OAI211_X1 U23198 ( .C1(n20242), .C2(n20735), .A(n20241), .B(n20240), .ZN(
        P1_U3064) );
  INV_X1 U23199 ( .A(n20299), .ZN(n20550) );
  INV_X1 U23200 ( .A(n20243), .ZN(n20246) );
  NOR2_X1 U23201 ( .A1(n13425), .A2(n20244), .ZN(n20322) );
  NAND3_X1 U23202 ( .A1(n20322), .A2(n20547), .A3(n13669), .ZN(n20245) );
  OAI21_X1 U23203 ( .B1(n20550), .B2(n20246), .A(n20245), .ZN(n20266) );
  NOR3_X1 U23204 ( .A1(n20487), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20276) );
  INV_X1 U23205 ( .A(n20276), .ZN(n20272) );
  NOR2_X1 U23206 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20272), .ZN(
        n20265) );
  AOI22_X1 U23207 ( .A1(n20584), .A2(n20266), .B1(n20583), .B2(n20265), .ZN(
        n20252) );
  INV_X1 U23208 ( .A(n20488), .ZN(n20352) );
  AOI21_X1 U23209 ( .B1(n20271), .B2(n20297), .A(n20906), .ZN(n20247) );
  AOI21_X1 U23210 ( .B1(n20322), .B2(n13669), .A(n20247), .ZN(n20248) );
  NOR2_X1 U23211 ( .A1(n20248), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20250) );
  AOI22_X1 U23212 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20268), .B1(
        n20267), .B2(n20590), .ZN(n20251) );
  OAI211_X1 U23213 ( .C1(n20593), .C2(n20271), .A(n20252), .B(n20251), .ZN(
        P1_U3065) );
  AOI22_X1 U23214 ( .A1(n20595), .A2(n20266), .B1(n20594), .B2(n20265), .ZN(
        n20254) );
  AOI22_X1 U23215 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20268), .B1(
        n20267), .B2(n20596), .ZN(n20253) );
  OAI211_X1 U23216 ( .C1(n20599), .C2(n20271), .A(n20254), .B(n20253), .ZN(
        P1_U3066) );
  AOI22_X1 U23217 ( .A1(n20601), .A2(n20266), .B1(n20600), .B2(n20265), .ZN(
        n20256) );
  AOI22_X1 U23218 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20268), .B1(
        n20267), .B2(n20602), .ZN(n20255) );
  OAI211_X1 U23219 ( .C1(n20605), .C2(n20271), .A(n20256), .B(n20255), .ZN(
        P1_U3067) );
  AOI22_X1 U23220 ( .A1(n20607), .A2(n20266), .B1(n20606), .B2(n20265), .ZN(
        n20258) );
  AOI22_X1 U23221 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20268), .B1(
        n20267), .B2(n20608), .ZN(n20257) );
  OAI211_X1 U23222 ( .C1(n20611), .C2(n20271), .A(n20258), .B(n20257), .ZN(
        P1_U3068) );
  AOI22_X1 U23223 ( .A1(n20613), .A2(n20266), .B1(n20612), .B2(n20265), .ZN(
        n20260) );
  AOI22_X1 U23224 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20268), .B1(
        n20267), .B2(n20614), .ZN(n20259) );
  OAI211_X1 U23225 ( .C1(n20617), .C2(n20271), .A(n20260), .B(n20259), .ZN(
        P1_U3069) );
  AOI22_X1 U23226 ( .A1(n20619), .A2(n20266), .B1(n20618), .B2(n20265), .ZN(
        n20262) );
  AOI22_X1 U23227 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20268), .B1(
        n20267), .B2(n20620), .ZN(n20261) );
  OAI211_X1 U23228 ( .C1(n20623), .C2(n20271), .A(n20262), .B(n20261), .ZN(
        P1_U3070) );
  AOI22_X1 U23229 ( .A1(n20625), .A2(n20266), .B1(n20624), .B2(n20265), .ZN(
        n20264) );
  AOI22_X1 U23230 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20268), .B1(
        n20267), .B2(n20626), .ZN(n20263) );
  OAI211_X1 U23231 ( .C1(n20629), .C2(n20271), .A(n20264), .B(n20263), .ZN(
        P1_U3071) );
  AOI22_X1 U23232 ( .A1(n20632), .A2(n20266), .B1(n20728), .B2(n20265), .ZN(
        n20270) );
  AOI22_X1 U23233 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20268), .B1(
        n20267), .B2(n20633), .ZN(n20269) );
  OAI211_X1 U23234 ( .C1(n20734), .C2(n20271), .A(n20270), .B(n20269), .ZN(
        P1_U3072) );
  NOR2_X1 U23235 ( .A1(n20517), .A2(n20272), .ZN(n20292) );
  AOI21_X1 U23236 ( .B1(n20322), .B2(n20518), .A(n20292), .ZN(n20273) );
  OAI22_X1 U23237 ( .A1(n20273), .A2(n20581), .B1(n20272), .B2(n20579), .ZN(
        n20293) );
  AOI22_X1 U23238 ( .A1(n20584), .A2(n20293), .B1(n20583), .B2(n20292), .ZN(
        n20279) );
  INV_X1 U23239 ( .A(n20328), .ZN(n20274) );
  OAI21_X1 U23240 ( .B1(n20274), .B2(n20906), .A(n20273), .ZN(n20275) );
  OAI221_X1 U23241 ( .B1(n20547), .B2(n20276), .C1(n20581), .C2(n20275), .A(
        n20587), .ZN(n20294) );
  INV_X1 U23242 ( .A(n20523), .ZN(n20277) );
  AOI22_X1 U23243 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20294), .B1(
        n20319), .B2(n20590), .ZN(n20278) );
  OAI211_X1 U23244 ( .C1(n20593), .C2(n20297), .A(n20279), .B(n20278), .ZN(
        P1_U3073) );
  AOI22_X1 U23245 ( .A1(n20595), .A2(n20293), .B1(n20594), .B2(n20292), .ZN(
        n20281) );
  AOI22_X1 U23246 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20294), .B1(
        n20319), .B2(n20596), .ZN(n20280) );
  OAI211_X1 U23247 ( .C1(n20599), .C2(n20297), .A(n20281), .B(n20280), .ZN(
        P1_U3074) );
  AOI22_X1 U23248 ( .A1(n20601), .A2(n20293), .B1(n20600), .B2(n20292), .ZN(
        n20283) );
  AOI22_X1 U23249 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20294), .B1(
        n20319), .B2(n20602), .ZN(n20282) );
  OAI211_X1 U23250 ( .C1(n20605), .C2(n20297), .A(n20283), .B(n20282), .ZN(
        P1_U3075) );
  AOI22_X1 U23251 ( .A1(n20607), .A2(n20293), .B1(n20606), .B2(n20292), .ZN(
        n20285) );
  AOI22_X1 U23252 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20294), .B1(
        n20319), .B2(n20608), .ZN(n20284) );
  OAI211_X1 U23253 ( .C1(n20611), .C2(n20297), .A(n20285), .B(n20284), .ZN(
        P1_U3076) );
  AOI22_X1 U23254 ( .A1(n20613), .A2(n20293), .B1(n20612), .B2(n20292), .ZN(
        n20287) );
  AOI22_X1 U23255 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20294), .B1(
        n20319), .B2(n20614), .ZN(n20286) );
  OAI211_X1 U23256 ( .C1(n20617), .C2(n20297), .A(n20287), .B(n20286), .ZN(
        P1_U3077) );
  AOI22_X1 U23257 ( .A1(n20619), .A2(n20293), .B1(n20618), .B2(n20292), .ZN(
        n20289) );
  AOI22_X1 U23258 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20294), .B1(
        n20319), .B2(n20620), .ZN(n20288) );
  OAI211_X1 U23259 ( .C1(n20623), .C2(n20297), .A(n20289), .B(n20288), .ZN(
        P1_U3078) );
  AOI22_X1 U23260 ( .A1(n20625), .A2(n20293), .B1(n20624), .B2(n20292), .ZN(
        n20291) );
  AOI22_X1 U23261 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20294), .B1(
        n20319), .B2(n20626), .ZN(n20290) );
  OAI211_X1 U23262 ( .C1(n20629), .C2(n20297), .A(n20291), .B(n20290), .ZN(
        P1_U3079) );
  AOI22_X1 U23263 ( .A1(n20632), .A2(n20293), .B1(n20728), .B2(n20292), .ZN(
        n20296) );
  AOI22_X1 U23264 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20294), .B1(
        n20319), .B2(n20633), .ZN(n20295) );
  OAI211_X1 U23265 ( .C1(n20734), .C2(n20297), .A(n20296), .B(n20295), .ZN(
        P1_U3080) );
  INV_X1 U23266 ( .A(n20319), .ZN(n20733) );
  NAND3_X1 U23267 ( .A1(n20729), .A2(n20733), .A3(n20547), .ZN(n20298) );
  NAND2_X1 U23268 ( .A1(n20298), .A2(n20408), .ZN(n20303) );
  AND2_X1 U23269 ( .A1(n20322), .A2(n20553), .ZN(n20301) );
  NOR2_X1 U23270 ( .A1(n20323), .A2(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n20318) );
  AOI22_X1 U23271 ( .A1(n20583), .A2(n20318), .B1(n20319), .B2(n20415), .ZN(
        n20307) );
  INV_X1 U23272 ( .A(n20301), .ZN(n20302) );
  INV_X1 U23273 ( .A(n20318), .ZN(n20731) );
  AOI22_X1 U23274 ( .A1(n20303), .A2(n20302), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20731), .ZN(n20305) );
  NAND3_X1 U23275 ( .A1(n20556), .A2(n20305), .A3(n20304), .ZN(n20739) );
  AOI22_X1 U23276 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20739), .B1(
        n20345), .B2(n20590), .ZN(n20306) );
  OAI211_X1 U23277 ( .C1(n20736), .C2(n20424), .A(n20307), .B(n20306), .ZN(
        P1_U3081) );
  AOI22_X1 U23278 ( .A1(n20594), .A2(n20318), .B1(n20345), .B2(n20596), .ZN(
        n20309) );
  AOI22_X1 U23279 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20739), .B1(
        n20319), .B2(n20425), .ZN(n20308) );
  OAI211_X1 U23280 ( .C1(n20736), .C2(n20428), .A(n20309), .B(n20308), .ZN(
        P1_U3082) );
  AOI22_X1 U23281 ( .A1(n20600), .A2(n20318), .B1(n20345), .B2(n20602), .ZN(
        n20311) );
  AOI22_X1 U23282 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20739), .B1(
        n20319), .B2(n20429), .ZN(n20310) );
  OAI211_X1 U23283 ( .C1(n20736), .C2(n20432), .A(n20311), .B(n20310), .ZN(
        P1_U3083) );
  AOI22_X1 U23284 ( .A1(n20606), .A2(n20318), .B1(n20319), .B2(n20433), .ZN(
        n20313) );
  AOI22_X1 U23285 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20739), .B1(
        n20345), .B2(n20608), .ZN(n20312) );
  OAI211_X1 U23286 ( .C1(n20736), .C2(n20436), .A(n20313), .B(n20312), .ZN(
        P1_U3084) );
  AOI22_X1 U23287 ( .A1(n20612), .A2(n20318), .B1(n20345), .B2(n20614), .ZN(
        n20315) );
  AOI22_X1 U23288 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20739), .B1(
        n20319), .B2(n20437), .ZN(n20314) );
  OAI211_X1 U23289 ( .C1(n20736), .C2(n20440), .A(n20315), .B(n20314), .ZN(
        P1_U3085) );
  AOI22_X1 U23290 ( .A1(n20618), .A2(n20318), .B1(n20319), .B2(n20441), .ZN(
        n20317) );
  AOI22_X1 U23291 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20739), .B1(
        n20345), .B2(n20620), .ZN(n20316) );
  OAI211_X1 U23292 ( .C1(n20736), .C2(n20444), .A(n20317), .B(n20316), .ZN(
        P1_U3086) );
  AOI22_X1 U23293 ( .A1(n20624), .A2(n20318), .B1(n20345), .B2(n20626), .ZN(
        n20321) );
  AOI22_X1 U23294 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20739), .B1(
        n20319), .B2(n20445), .ZN(n20320) );
  OAI211_X1 U23295 ( .C1(n20736), .C2(n20448), .A(n20321), .B(n20320), .ZN(
        P1_U3087) );
  AOI21_X1 U23296 ( .B1(n20322), .B2(n9837), .A(n20343), .ZN(n20324) );
  OAI22_X1 U23297 ( .A1(n20324), .A2(n20581), .B1(n20323), .B2(n20579), .ZN(
        n20344) );
  AOI22_X1 U23298 ( .A1(n20584), .A2(n20344), .B1(n20583), .B2(n20343), .ZN(
        n20330) );
  INV_X1 U23299 ( .A(n20323), .ZN(n20327) );
  NAND2_X1 U23300 ( .A1(n20325), .A2(n20324), .ZN(n20326) );
  OAI221_X1 U23301 ( .B1(n20547), .B2(n20327), .C1(n20581), .C2(n20326), .A(
        n20587), .ZN(n20346) );
  AOI22_X1 U23302 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20346), .B1(
        n20353), .B2(n20590), .ZN(n20329) );
  OAI211_X1 U23303 ( .C1(n20593), .C2(n20729), .A(n20330), .B(n20329), .ZN(
        P1_U3089) );
  AOI22_X1 U23304 ( .A1(n20595), .A2(n20344), .B1(n20594), .B2(n20343), .ZN(
        n20332) );
  AOI22_X1 U23305 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20346), .B1(
        n20353), .B2(n20596), .ZN(n20331) );
  OAI211_X1 U23306 ( .C1(n20599), .C2(n20729), .A(n20332), .B(n20331), .ZN(
        P1_U3090) );
  AOI22_X1 U23307 ( .A1(n20601), .A2(n20344), .B1(n20600), .B2(n20343), .ZN(
        n20334) );
  AOI22_X1 U23308 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20346), .B1(
        n20353), .B2(n20602), .ZN(n20333) );
  OAI211_X1 U23309 ( .C1(n20605), .C2(n20729), .A(n20334), .B(n20333), .ZN(
        P1_U3091) );
  AOI22_X1 U23310 ( .A1(n20607), .A2(n20344), .B1(n20606), .B2(n20343), .ZN(
        n20336) );
  AOI22_X1 U23311 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20346), .B1(
        n20353), .B2(n20608), .ZN(n20335) );
  OAI211_X1 U23312 ( .C1(n20611), .C2(n20729), .A(n20336), .B(n20335), .ZN(
        P1_U3092) );
  AOI22_X1 U23313 ( .A1(n20613), .A2(n20344), .B1(n20612), .B2(n20343), .ZN(
        n20338) );
  AOI22_X1 U23314 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20346), .B1(
        n20353), .B2(n20614), .ZN(n20337) );
  OAI211_X1 U23315 ( .C1(n20617), .C2(n20729), .A(n20338), .B(n20337), .ZN(
        P1_U3093) );
  AOI22_X1 U23316 ( .A1(n20619), .A2(n20344), .B1(n20618), .B2(n20343), .ZN(
        n20340) );
  AOI22_X1 U23317 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20346), .B1(
        n20353), .B2(n20620), .ZN(n20339) );
  OAI211_X1 U23318 ( .C1(n20623), .C2(n20729), .A(n20340), .B(n20339), .ZN(
        P1_U3094) );
  AOI22_X1 U23319 ( .A1(n20625), .A2(n20344), .B1(n20624), .B2(n20343), .ZN(
        n20342) );
  AOI22_X1 U23320 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20346), .B1(
        n20353), .B2(n20626), .ZN(n20341) );
  OAI211_X1 U23321 ( .C1(n20629), .C2(n20729), .A(n20342), .B(n20341), .ZN(
        P1_U3095) );
  AOI22_X1 U23322 ( .A1(n20632), .A2(n20344), .B1(n20728), .B2(n20343), .ZN(
        n20348) );
  AOI22_X1 U23323 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20346), .B1(
        n20345), .B2(n20542), .ZN(n20347) );
  OAI211_X1 U23324 ( .C1(n20730), .C2(n20376), .A(n20348), .B(n20347), .ZN(
        P1_U3096) );
  NAND2_X1 U23325 ( .A1(n20349), .A2(n13425), .ZN(n20410) );
  INV_X1 U23326 ( .A(n20410), .ZN(n20456) );
  NOR3_X1 U23327 ( .A1(n20486), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20380) );
  INV_X1 U23328 ( .A(n20380), .ZN(n20382) );
  NOR2_X1 U23329 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20382), .ZN(
        n20371) );
  AOI21_X1 U23330 ( .B1(n20456), .B2(n13669), .A(n20371), .ZN(n20354) );
  INV_X1 U23331 ( .A(n20413), .ZN(n20351) );
  NAND2_X1 U23332 ( .A1(n20350), .A2(n20411), .ZN(n20494) );
  OAI22_X1 U23333 ( .A1(n20354), .A2(n20581), .B1(n20351), .B2(n20494), .ZN(
        n20372) );
  AOI22_X1 U23334 ( .A1(n20584), .A2(n20372), .B1(n20583), .B2(n20371), .ZN(
        n20358) );
  OAI21_X1 U23335 ( .B1(n20384), .B2(n20353), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20355) );
  NAND2_X1 U23336 ( .A1(n20355), .A2(n20354), .ZN(n20356) );
  AOI22_X1 U23337 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20373), .B1(
        n20384), .B2(n20590), .ZN(n20357) );
  OAI211_X1 U23338 ( .C1(n20593), .C2(n20376), .A(n20358), .B(n20357), .ZN(
        P1_U3097) );
  AOI22_X1 U23339 ( .A1(n20595), .A2(n20372), .B1(n20594), .B2(n20371), .ZN(
        n20360) );
  AOI22_X1 U23340 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20373), .B1(
        n20384), .B2(n20596), .ZN(n20359) );
  OAI211_X1 U23341 ( .C1(n20599), .C2(n20376), .A(n20360), .B(n20359), .ZN(
        P1_U3098) );
  AOI22_X1 U23342 ( .A1(n20601), .A2(n20372), .B1(n20600), .B2(n20371), .ZN(
        n20362) );
  AOI22_X1 U23343 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20373), .B1(
        n20384), .B2(n20602), .ZN(n20361) );
  OAI211_X1 U23344 ( .C1(n20605), .C2(n20376), .A(n20362), .B(n20361), .ZN(
        P1_U3099) );
  AOI22_X1 U23345 ( .A1(n20607), .A2(n20372), .B1(n20606), .B2(n20371), .ZN(
        n20364) );
  AOI22_X1 U23346 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20373), .B1(
        n20384), .B2(n20608), .ZN(n20363) );
  OAI211_X1 U23347 ( .C1(n20611), .C2(n20376), .A(n20364), .B(n20363), .ZN(
        P1_U3100) );
  AOI22_X1 U23348 ( .A1(n20613), .A2(n20372), .B1(n20612), .B2(n20371), .ZN(
        n20366) );
  AOI22_X1 U23349 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20373), .B1(
        n20384), .B2(n20614), .ZN(n20365) );
  OAI211_X1 U23350 ( .C1(n20617), .C2(n20376), .A(n20366), .B(n20365), .ZN(
        P1_U3101) );
  AOI22_X1 U23351 ( .A1(n20619), .A2(n20372), .B1(n20618), .B2(n20371), .ZN(
        n20368) );
  AOI22_X1 U23352 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20373), .B1(
        n20384), .B2(n20620), .ZN(n20367) );
  OAI211_X1 U23353 ( .C1(n20623), .C2(n20376), .A(n20368), .B(n20367), .ZN(
        P1_U3102) );
  AOI22_X1 U23354 ( .A1(n20625), .A2(n20372), .B1(n20624), .B2(n20371), .ZN(
        n20370) );
  AOI22_X1 U23355 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20373), .B1(
        n20384), .B2(n20626), .ZN(n20369) );
  OAI211_X1 U23356 ( .C1(n20629), .C2(n20376), .A(n20370), .B(n20369), .ZN(
        P1_U3103) );
  AOI22_X1 U23357 ( .A1(n20632), .A2(n20372), .B1(n20728), .B2(n20371), .ZN(
        n20375) );
  AOI22_X1 U23358 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20373), .B1(
        n20384), .B2(n20633), .ZN(n20374) );
  OAI211_X1 U23359 ( .C1(n20734), .C2(n20376), .A(n20375), .B(n20374), .ZN(
        P1_U3104) );
  OR2_X1 U23360 ( .A1(n20410), .A2(n20377), .ZN(n20379) );
  NOR2_X1 U23361 ( .A1(n20517), .A2(n20382), .ZN(n20400) );
  INV_X1 U23362 ( .A(n20400), .ZN(n20378) );
  AND2_X1 U23363 ( .A1(n20379), .A2(n20378), .ZN(n20383) );
  OAI21_X1 U23364 ( .B1(n20460), .B2(n20906), .A(n20383), .ZN(n20381) );
  OAI221_X1 U23365 ( .B1(n20381), .B2(n20581), .C1(n20380), .C2(n20547), .A(
        n20587), .ZN(n20402) );
  INV_X1 U23366 ( .A(n20402), .ZN(n20387) );
  INV_X1 U23367 ( .A(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n20885) );
  OAI22_X1 U23368 ( .A1(n20383), .A2(n20581), .B1(n20382), .B2(n20579), .ZN(
        n20401) );
  AOI22_X1 U23369 ( .A1(n20584), .A2(n20401), .B1(n20583), .B2(n20400), .ZN(
        n20386) );
  AOI22_X1 U23370 ( .A1(n20384), .A2(n20415), .B1(n20450), .B2(n20590), .ZN(
        n20385) );
  OAI211_X1 U23371 ( .C1(n20387), .C2(n20885), .A(n20386), .B(n20385), .ZN(
        P1_U3105) );
  AOI22_X1 U23372 ( .A1(n20595), .A2(n20401), .B1(n20594), .B2(n20400), .ZN(
        n20389) );
  AOI22_X1 U23373 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20402), .B1(
        n20450), .B2(n20596), .ZN(n20388) );
  OAI211_X1 U23374 ( .C1(n20599), .C2(n20405), .A(n20389), .B(n20388), .ZN(
        P1_U3106) );
  AOI22_X1 U23375 ( .A1(n20601), .A2(n20401), .B1(n20600), .B2(n20400), .ZN(
        n20391) );
  AOI22_X1 U23376 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20402), .B1(
        n20450), .B2(n20602), .ZN(n20390) );
  OAI211_X1 U23377 ( .C1(n20605), .C2(n20405), .A(n20391), .B(n20390), .ZN(
        P1_U3107) );
  AOI22_X1 U23378 ( .A1(n20607), .A2(n20401), .B1(n20606), .B2(n20400), .ZN(
        n20393) );
  AOI22_X1 U23379 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20402), .B1(
        n20450), .B2(n20608), .ZN(n20392) );
  OAI211_X1 U23380 ( .C1(n20611), .C2(n20405), .A(n20393), .B(n20392), .ZN(
        P1_U3108) );
  AOI22_X1 U23381 ( .A1(n20613), .A2(n20401), .B1(n20612), .B2(n20400), .ZN(
        n20395) );
  AOI22_X1 U23382 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20402), .B1(
        n20450), .B2(n20614), .ZN(n20394) );
  OAI211_X1 U23383 ( .C1(n20617), .C2(n20405), .A(n20395), .B(n20394), .ZN(
        P1_U3109) );
  AOI22_X1 U23384 ( .A1(n20619), .A2(n20401), .B1(n20618), .B2(n20400), .ZN(
        n20397) );
  AOI22_X1 U23385 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20402), .B1(
        n20450), .B2(n20620), .ZN(n20396) );
  OAI211_X1 U23386 ( .C1(n20623), .C2(n20405), .A(n20397), .B(n20396), .ZN(
        P1_U3110) );
  AOI22_X1 U23387 ( .A1(n20625), .A2(n20401), .B1(n20624), .B2(n20400), .ZN(
        n20399) );
  AOI22_X1 U23388 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20402), .B1(
        n20450), .B2(n20626), .ZN(n20398) );
  OAI211_X1 U23389 ( .C1(n20629), .C2(n20405), .A(n20399), .B(n20398), .ZN(
        P1_U3111) );
  AOI22_X1 U23390 ( .A1(n20632), .A2(n20401), .B1(n20728), .B2(n20400), .ZN(
        n20404) );
  AOI22_X1 U23391 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20402), .B1(
        n20450), .B2(n20633), .ZN(n20403) );
  OAI211_X1 U23392 ( .C1(n20734), .C2(n20405), .A(n20404), .B(n20403), .ZN(
        P1_U3112) );
  INV_X1 U23393 ( .A(n20450), .ZN(n20407) );
  NAND3_X1 U23394 ( .A1(n20407), .A2(n20547), .A3(n20480), .ZN(n20409) );
  NAND2_X1 U23395 ( .A1(n20409), .A2(n20408), .ZN(n20419) );
  NOR2_X1 U23396 ( .A1(n20410), .A2(n13669), .ZN(n20416) );
  OR2_X1 U23397 ( .A1(n20411), .A2(n20486), .ZN(n20549) );
  INV_X1 U23398 ( .A(n20549), .ZN(n20412) );
  NOR3_X1 U23399 ( .A1(n20486), .A2(n20414), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20462) );
  NAND2_X1 U23400 ( .A1(n20517), .A2(n20462), .ZN(n20417) );
  INV_X1 U23401 ( .A(n20417), .ZN(n20449) );
  AOI22_X1 U23402 ( .A1(n20450), .A2(n20415), .B1(n20583), .B2(n20449), .ZN(
        n20423) );
  INV_X1 U23403 ( .A(n20416), .ZN(n20418) );
  AOI22_X1 U23404 ( .A1(n20419), .A2(n20418), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20417), .ZN(n20420) );
  NAND2_X1 U23405 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20549), .ZN(n20555) );
  NAND3_X1 U23406 ( .A1(n20421), .A2(n20420), .A3(n20555), .ZN(n20451) );
  AOI22_X1 U23407 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20451), .B1(
        n20482), .B2(n20590), .ZN(n20422) );
  OAI211_X1 U23408 ( .C1(n20454), .C2(n20424), .A(n20423), .B(n20422), .ZN(
        P1_U3113) );
  AOI22_X1 U23409 ( .A1(n20482), .A2(n20596), .B1(n20594), .B2(n20449), .ZN(
        n20427) );
  AOI22_X1 U23410 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20451), .B1(
        n20450), .B2(n20425), .ZN(n20426) );
  OAI211_X1 U23411 ( .C1(n20454), .C2(n20428), .A(n20427), .B(n20426), .ZN(
        P1_U3114) );
  AOI22_X1 U23412 ( .A1(n20482), .A2(n20602), .B1(n20600), .B2(n20449), .ZN(
        n20431) );
  AOI22_X1 U23413 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20451), .B1(
        n20450), .B2(n20429), .ZN(n20430) );
  OAI211_X1 U23414 ( .C1(n20454), .C2(n20432), .A(n20431), .B(n20430), .ZN(
        P1_U3115) );
  AOI22_X1 U23415 ( .A1(n20450), .A2(n20433), .B1(n20606), .B2(n20449), .ZN(
        n20435) );
  AOI22_X1 U23416 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20451), .B1(
        n20482), .B2(n20608), .ZN(n20434) );
  OAI211_X1 U23417 ( .C1(n20454), .C2(n20436), .A(n20435), .B(n20434), .ZN(
        P1_U3116) );
  AOI22_X1 U23418 ( .A1(n20482), .A2(n20614), .B1(n20612), .B2(n20449), .ZN(
        n20439) );
  AOI22_X1 U23419 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20451), .B1(
        n20450), .B2(n20437), .ZN(n20438) );
  OAI211_X1 U23420 ( .C1(n20454), .C2(n20440), .A(n20439), .B(n20438), .ZN(
        P1_U3117) );
  AOI22_X1 U23421 ( .A1(n20450), .A2(n20441), .B1(n20618), .B2(n20449), .ZN(
        n20443) );
  AOI22_X1 U23422 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20451), .B1(
        n20482), .B2(n20620), .ZN(n20442) );
  OAI211_X1 U23423 ( .C1(n20454), .C2(n20444), .A(n20443), .B(n20442), .ZN(
        P1_U3118) );
  AOI22_X1 U23424 ( .A1(n20450), .A2(n20445), .B1(n20624), .B2(n20449), .ZN(
        n20447) );
  AOI22_X1 U23425 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20451), .B1(
        n20482), .B2(n20626), .ZN(n20446) );
  OAI211_X1 U23426 ( .C1(n20454), .C2(n20448), .A(n20447), .B(n20446), .ZN(
        P1_U3119) );
  AOI22_X1 U23427 ( .A1(n20450), .A2(n20542), .B1(n20728), .B2(n20449), .ZN(
        n20453) );
  AOI22_X1 U23428 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20451), .B1(
        n20482), .B2(n20633), .ZN(n20452) );
  OAI211_X1 U23429 ( .C1(n20454), .C2(n20735), .A(n20453), .B(n20452), .ZN(
        P1_U3120) );
  AOI21_X1 U23430 ( .B1(n20456), .B2(n9837), .A(n10143), .ZN(n20458) );
  INV_X1 U23431 ( .A(n20462), .ZN(n20457) );
  OAI22_X1 U23432 ( .A1(n20458), .A2(n20581), .B1(n20457), .B2(n20579), .ZN(
        n20481) );
  AOI22_X1 U23433 ( .A1(n20584), .A2(n20481), .B1(n20583), .B2(n10143), .ZN(
        n20466) );
  NAND2_X1 U23434 ( .A1(n20459), .A2(n20547), .ZN(n20586) );
  NOR2_X1 U23435 ( .A1(n20460), .A2(n20586), .ZN(n20461) );
  OAI21_X1 U23436 ( .B1(n20462), .B2(n20461), .A(n20587), .ZN(n20483) );
  AOI22_X1 U23437 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20483), .B1(
        n20477), .B2(n20590), .ZN(n20465) );
  OAI211_X1 U23438 ( .C1(n20593), .C2(n20480), .A(n20466), .B(n20465), .ZN(
        P1_U3121) );
  AOI22_X1 U23439 ( .A1(n20595), .A2(n20481), .B1(n20594), .B2(n10143), .ZN(
        n20468) );
  AOI22_X1 U23440 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20483), .B1(
        n20477), .B2(n20596), .ZN(n20467) );
  OAI211_X1 U23441 ( .C1(n20599), .C2(n20480), .A(n20468), .B(n20467), .ZN(
        P1_U3122) );
  AOI22_X1 U23442 ( .A1(n20601), .A2(n20481), .B1(n20600), .B2(n10143), .ZN(
        n20470) );
  AOI22_X1 U23443 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20483), .B1(
        n20477), .B2(n20602), .ZN(n20469) );
  OAI211_X1 U23444 ( .C1(n20605), .C2(n20480), .A(n20470), .B(n20469), .ZN(
        P1_U3123) );
  AOI22_X1 U23445 ( .A1(n20607), .A2(n20481), .B1(n20606), .B2(n10143), .ZN(
        n20472) );
  AOI22_X1 U23446 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20483), .B1(
        n20477), .B2(n20608), .ZN(n20471) );
  OAI211_X1 U23447 ( .C1(n20611), .C2(n20480), .A(n20472), .B(n20471), .ZN(
        P1_U3124) );
  AOI22_X1 U23448 ( .A1(n20613), .A2(n20481), .B1(n20612), .B2(n10143), .ZN(
        n20474) );
  AOI22_X1 U23449 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20483), .B1(
        n20477), .B2(n20614), .ZN(n20473) );
  OAI211_X1 U23450 ( .C1(n20617), .C2(n20480), .A(n20474), .B(n20473), .ZN(
        P1_U3125) );
  AOI22_X1 U23451 ( .A1(n20619), .A2(n20481), .B1(n20618), .B2(n10143), .ZN(
        n20476) );
  AOI22_X1 U23452 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20483), .B1(
        n20477), .B2(n20620), .ZN(n20475) );
  OAI211_X1 U23453 ( .C1(n20623), .C2(n20480), .A(n20476), .B(n20475), .ZN(
        P1_U3126) );
  AOI22_X1 U23454 ( .A1(n20625), .A2(n20481), .B1(n20624), .B2(n10143), .ZN(
        n20479) );
  AOI22_X1 U23455 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20483), .B1(
        n20477), .B2(n20626), .ZN(n20478) );
  OAI211_X1 U23456 ( .C1(n20629), .C2(n20480), .A(n20479), .B(n20478), .ZN(
        P1_U3127) );
  AOI22_X1 U23457 ( .A1(n20632), .A2(n20481), .B1(n20728), .B2(n10143), .ZN(
        n20485) );
  AOI22_X1 U23458 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20483), .B1(
        n20482), .B2(n20542), .ZN(n20484) );
  OAI211_X1 U23459 ( .C1(n20730), .C2(n20516), .A(n20485), .B(n20484), .ZN(
        P1_U3128) );
  NOR3_X1 U23460 ( .A1(n20487), .A2(n20486), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20522) );
  INV_X1 U23461 ( .A(n20522), .ZN(n20519) );
  NOR2_X1 U23462 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20519), .ZN(
        n20511) );
  AOI22_X1 U23463 ( .A1(n20583), .A2(n20511), .B1(n20543), .B2(n20590), .ZN(
        n20498) );
  NAND2_X1 U23464 ( .A1(n20516), .A2(n20539), .ZN(n20489) );
  AOI21_X1 U23465 ( .B1(n20489), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20581), 
        .ZN(n20493) );
  NAND2_X1 U23466 ( .A1(n10137), .A2(n13669), .ZN(n20495) );
  AOI22_X1 U23467 ( .A1(n20493), .A2(n20495), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20494), .ZN(n20491) );
  OAI211_X1 U23468 ( .C1(n20511), .C2(n20492), .A(n20556), .B(n20491), .ZN(
        n20513) );
  INV_X1 U23469 ( .A(n20493), .ZN(n20496) );
  OAI22_X1 U23470 ( .A1(n20496), .A2(n20495), .B1(n20550), .B2(n20494), .ZN(
        n20512) );
  AOI22_X1 U23471 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20513), .B1(
        n20584), .B2(n20512), .ZN(n20497) );
  OAI211_X1 U23472 ( .C1(n20593), .C2(n20516), .A(n20498), .B(n20497), .ZN(
        P1_U3129) );
  AOI22_X1 U23473 ( .A1(n20594), .A2(n20511), .B1(n20543), .B2(n20596), .ZN(
        n20500) );
  AOI22_X1 U23474 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20513), .B1(
        n20595), .B2(n20512), .ZN(n20499) );
  OAI211_X1 U23475 ( .C1(n20599), .C2(n20516), .A(n20500), .B(n20499), .ZN(
        P1_U3130) );
  AOI22_X1 U23476 ( .A1(n20600), .A2(n20511), .B1(n20543), .B2(n20602), .ZN(
        n20502) );
  AOI22_X1 U23477 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20513), .B1(
        n20601), .B2(n20512), .ZN(n20501) );
  OAI211_X1 U23478 ( .C1(n20605), .C2(n20516), .A(n20502), .B(n20501), .ZN(
        P1_U3131) );
  AOI22_X1 U23479 ( .A1(n20606), .A2(n20511), .B1(n20543), .B2(n20608), .ZN(
        n20504) );
  AOI22_X1 U23480 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20513), .B1(
        n20607), .B2(n20512), .ZN(n20503) );
  OAI211_X1 U23481 ( .C1(n20611), .C2(n20516), .A(n20504), .B(n20503), .ZN(
        P1_U3132) );
  AOI22_X1 U23482 ( .A1(n20612), .A2(n20511), .B1(n20543), .B2(n20614), .ZN(
        n20506) );
  AOI22_X1 U23483 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20513), .B1(
        n20613), .B2(n20512), .ZN(n20505) );
  OAI211_X1 U23484 ( .C1(n20617), .C2(n20516), .A(n20506), .B(n20505), .ZN(
        P1_U3133) );
  AOI22_X1 U23485 ( .A1(n20618), .A2(n20511), .B1(n20543), .B2(n20620), .ZN(
        n20508) );
  AOI22_X1 U23486 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20513), .B1(
        n20619), .B2(n20512), .ZN(n20507) );
  OAI211_X1 U23487 ( .C1(n20623), .C2(n20516), .A(n20508), .B(n20507), .ZN(
        P1_U3134) );
  AOI22_X1 U23488 ( .A1(n20624), .A2(n20511), .B1(n20543), .B2(n20626), .ZN(
        n20510) );
  AOI22_X1 U23489 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20513), .B1(
        n20625), .B2(n20512), .ZN(n20509) );
  OAI211_X1 U23490 ( .C1(n20629), .C2(n20516), .A(n20510), .B(n20509), .ZN(
        P1_U3135) );
  AOI22_X1 U23491 ( .A1(n20728), .A2(n20511), .B1(n20543), .B2(n20633), .ZN(
        n20515) );
  AOI22_X1 U23492 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20513), .B1(
        n20632), .B2(n20512), .ZN(n20514) );
  OAI211_X1 U23493 ( .C1(n20734), .C2(n20516), .A(n20515), .B(n20514), .ZN(
        P1_U3136) );
  NOR2_X1 U23494 ( .A1(n20517), .A2(n20519), .ZN(n20540) );
  AOI21_X1 U23495 ( .B1(n10137), .B2(n20518), .A(n20540), .ZN(n20520) );
  OAI22_X1 U23496 ( .A1(n20520), .A2(n20581), .B1(n20519), .B2(n20579), .ZN(
        n20541) );
  AOI22_X1 U23497 ( .A1(n20584), .A2(n20541), .B1(n20583), .B2(n20540), .ZN(
        n20525) );
  OAI21_X1 U23498 ( .B1(n20585), .B2(n20906), .A(n20520), .ZN(n20521) );
  OAI221_X1 U23499 ( .B1(n20547), .B2(n20522), .C1(n20581), .C2(n20521), .A(
        n20587), .ZN(n20544) );
  AOI22_X1 U23500 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20544), .B1(
        n20536), .B2(n20590), .ZN(n20524) );
  OAI211_X1 U23501 ( .C1(n20593), .C2(n20539), .A(n20525), .B(n20524), .ZN(
        P1_U3137) );
  AOI22_X1 U23502 ( .A1(n20595), .A2(n20541), .B1(n20594), .B2(n20540), .ZN(
        n20527) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20544), .B1(
        n20536), .B2(n20596), .ZN(n20526) );
  OAI211_X1 U23504 ( .C1(n20599), .C2(n20539), .A(n20527), .B(n20526), .ZN(
        P1_U3138) );
  AOI22_X1 U23505 ( .A1(n20601), .A2(n20541), .B1(n20600), .B2(n20540), .ZN(
        n20529) );
  AOI22_X1 U23506 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20544), .B1(
        n20536), .B2(n20602), .ZN(n20528) );
  OAI211_X1 U23507 ( .C1(n20605), .C2(n20539), .A(n20529), .B(n20528), .ZN(
        P1_U3139) );
  AOI22_X1 U23508 ( .A1(n20607), .A2(n20541), .B1(n20606), .B2(n20540), .ZN(
        n20531) );
  AOI22_X1 U23509 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20544), .B1(
        n20536), .B2(n20608), .ZN(n20530) );
  OAI211_X1 U23510 ( .C1(n20611), .C2(n20539), .A(n20531), .B(n20530), .ZN(
        P1_U3140) );
  AOI22_X1 U23511 ( .A1(n20613), .A2(n20541), .B1(n20612), .B2(n20540), .ZN(
        n20533) );
  AOI22_X1 U23512 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20544), .B1(
        n20536), .B2(n20614), .ZN(n20532) );
  OAI211_X1 U23513 ( .C1(n20617), .C2(n20539), .A(n20533), .B(n20532), .ZN(
        P1_U3141) );
  AOI22_X1 U23514 ( .A1(n20619), .A2(n20541), .B1(n20618), .B2(n20540), .ZN(
        n20535) );
  AOI22_X1 U23515 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20544), .B1(
        n20536), .B2(n20620), .ZN(n20534) );
  OAI211_X1 U23516 ( .C1(n20623), .C2(n20539), .A(n20535), .B(n20534), .ZN(
        P1_U3142) );
  AOI22_X1 U23517 ( .A1(n20625), .A2(n20541), .B1(n20624), .B2(n20540), .ZN(
        n20538) );
  AOI22_X1 U23518 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20544), .B1(
        n20536), .B2(n20626), .ZN(n20537) );
  OAI211_X1 U23519 ( .C1(n20629), .C2(n20539), .A(n20538), .B(n20537), .ZN(
        P1_U3143) );
  AOI22_X1 U23520 ( .A1(n20632), .A2(n20541), .B1(n20728), .B2(n20540), .ZN(
        n20546) );
  AOI22_X1 U23521 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20542), .ZN(n20545) );
  OAI211_X1 U23522 ( .C1(n20730), .C2(n20578), .A(n20546), .B(n20545), .ZN(
        P1_U3144) );
  NAND3_X1 U23523 ( .A1(n10137), .A2(n20553), .A3(n20547), .ZN(n20548) );
  OAI21_X1 U23524 ( .B1(n20550), .B2(n20549), .A(n20548), .ZN(n20573) );
  NOR2_X1 U23525 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20580), .ZN(
        n20572) );
  AOI22_X1 U23526 ( .A1(n20584), .A2(n20573), .B1(n20583), .B2(n20572), .ZN(
        n20559) );
  AOI21_X1 U23527 ( .B1(n20638), .B2(n20578), .A(n20906), .ZN(n20552) );
  AOI21_X1 U23528 ( .B1(n10137), .B2(n20553), .A(n20552), .ZN(n20554) );
  NOR2_X1 U23529 ( .A1(n20554), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20557) );
  OAI211_X1 U23530 ( .C1(n20572), .C2(n20557), .A(n20556), .B(n20555), .ZN(
        n20575) );
  AOI22_X1 U23531 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20575), .B1(
        n20574), .B2(n20590), .ZN(n20558) );
  OAI211_X1 U23532 ( .C1(n20593), .C2(n20578), .A(n20559), .B(n20558), .ZN(
        P1_U3145) );
  AOI22_X1 U23533 ( .A1(n20595), .A2(n20573), .B1(n20594), .B2(n20572), .ZN(
        n20561) );
  AOI22_X1 U23534 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20575), .B1(
        n20574), .B2(n20596), .ZN(n20560) );
  OAI211_X1 U23535 ( .C1(n20599), .C2(n20578), .A(n20561), .B(n20560), .ZN(
        P1_U3146) );
  AOI22_X1 U23536 ( .A1(n20601), .A2(n20573), .B1(n20600), .B2(n20572), .ZN(
        n20563) );
  AOI22_X1 U23537 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20575), .B1(
        n20574), .B2(n20602), .ZN(n20562) );
  OAI211_X1 U23538 ( .C1(n20605), .C2(n20578), .A(n20563), .B(n20562), .ZN(
        P1_U3147) );
  AOI22_X1 U23539 ( .A1(n20607), .A2(n20573), .B1(n20606), .B2(n20572), .ZN(
        n20565) );
  AOI22_X1 U23540 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20575), .B1(
        n20574), .B2(n20608), .ZN(n20564) );
  OAI211_X1 U23541 ( .C1(n20611), .C2(n20578), .A(n20565), .B(n20564), .ZN(
        P1_U3148) );
  AOI22_X1 U23542 ( .A1(n20613), .A2(n20573), .B1(n20612), .B2(n20572), .ZN(
        n20567) );
  AOI22_X1 U23543 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20575), .B1(
        n20574), .B2(n20614), .ZN(n20566) );
  OAI211_X1 U23544 ( .C1(n20617), .C2(n20578), .A(n20567), .B(n20566), .ZN(
        P1_U3149) );
  AOI22_X1 U23545 ( .A1(n20619), .A2(n20573), .B1(n20618), .B2(n20572), .ZN(
        n20569) );
  AOI22_X1 U23546 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20575), .B1(
        n20574), .B2(n20620), .ZN(n20568) );
  OAI211_X1 U23547 ( .C1(n20623), .C2(n20578), .A(n20569), .B(n20568), .ZN(
        P1_U3150) );
  AOI22_X1 U23548 ( .A1(n20625), .A2(n20573), .B1(n20624), .B2(n20572), .ZN(
        n20571) );
  AOI22_X1 U23549 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20575), .B1(
        n20574), .B2(n20626), .ZN(n20570) );
  OAI211_X1 U23550 ( .C1(n20629), .C2(n20578), .A(n20571), .B(n20570), .ZN(
        P1_U3151) );
  AOI22_X1 U23551 ( .A1(n20632), .A2(n20573), .B1(n20728), .B2(n20572), .ZN(
        n20577) );
  AOI22_X1 U23552 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20575), .B1(
        n20574), .B2(n20633), .ZN(n20576) );
  OAI211_X1 U23553 ( .C1(n20734), .C2(n20578), .A(n20577), .B(n20576), .ZN(
        P1_U3152) );
  AOI21_X1 U23554 ( .B1(n10137), .B2(n9837), .A(n20630), .ZN(n20582) );
  OAI22_X1 U23555 ( .A1(n20582), .A2(n20581), .B1(n20580), .B2(n20579), .ZN(
        n20631) );
  AOI22_X1 U23556 ( .A1(n20584), .A2(n20631), .B1(n20583), .B2(n20630), .ZN(
        n20592) );
  NOR2_X1 U23557 ( .A1(n20586), .A2(n20585), .ZN(n20588) );
  OAI21_X1 U23558 ( .B1(n20589), .B2(n20588), .A(n20587), .ZN(n20635) );
  AOI22_X1 U23559 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20635), .B1(
        n20634), .B2(n20590), .ZN(n20591) );
  OAI211_X1 U23560 ( .C1(n20593), .C2(n20638), .A(n20592), .B(n20591), .ZN(
        P1_U3153) );
  AOI22_X1 U23561 ( .A1(n20595), .A2(n20631), .B1(n20594), .B2(n20630), .ZN(
        n20598) );
  AOI22_X1 U23562 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20635), .B1(
        n20634), .B2(n20596), .ZN(n20597) );
  OAI211_X1 U23563 ( .C1(n20599), .C2(n20638), .A(n20598), .B(n20597), .ZN(
        P1_U3154) );
  AOI22_X1 U23564 ( .A1(n20601), .A2(n20631), .B1(n20600), .B2(n20630), .ZN(
        n20604) );
  AOI22_X1 U23565 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20635), .B1(
        n20634), .B2(n20602), .ZN(n20603) );
  OAI211_X1 U23566 ( .C1(n20605), .C2(n20638), .A(n20604), .B(n20603), .ZN(
        P1_U3155) );
  AOI22_X1 U23567 ( .A1(n20607), .A2(n20631), .B1(n20606), .B2(n20630), .ZN(
        n20610) );
  AOI22_X1 U23568 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20635), .B1(
        n20634), .B2(n20608), .ZN(n20609) );
  OAI211_X1 U23569 ( .C1(n20611), .C2(n20638), .A(n20610), .B(n20609), .ZN(
        P1_U3156) );
  AOI22_X1 U23570 ( .A1(n20613), .A2(n20631), .B1(n20612), .B2(n20630), .ZN(
        n20616) );
  AOI22_X1 U23571 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20635), .B1(
        n20634), .B2(n20614), .ZN(n20615) );
  OAI211_X1 U23572 ( .C1(n20617), .C2(n20638), .A(n20616), .B(n20615), .ZN(
        P1_U3157) );
  AOI22_X1 U23573 ( .A1(n20619), .A2(n20631), .B1(n20618), .B2(n20630), .ZN(
        n20622) );
  AOI22_X1 U23574 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20635), .B1(
        n20634), .B2(n20620), .ZN(n20621) );
  OAI211_X1 U23575 ( .C1(n20623), .C2(n20638), .A(n20622), .B(n20621), .ZN(
        P1_U3158) );
  AOI22_X1 U23576 ( .A1(n20625), .A2(n20631), .B1(n20624), .B2(n20630), .ZN(
        n20628) );
  AOI22_X1 U23577 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20635), .B1(
        n20634), .B2(n20626), .ZN(n20627) );
  OAI211_X1 U23578 ( .C1(n20629), .C2(n20638), .A(n20628), .B(n20627), .ZN(
        P1_U3159) );
  AOI22_X1 U23579 ( .A1(n20632), .A2(n20631), .B1(n20728), .B2(n20630), .ZN(
        n20637) );
  AOI22_X1 U23580 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20635), .B1(
        n20634), .B2(n20633), .ZN(n20636) );
  OAI211_X1 U23581 ( .C1(n20734), .C2(n20638), .A(n20637), .B(n20636), .ZN(
        P1_U3160) );
  NOR2_X1 U23582 ( .A1(n20639), .A2(n14146), .ZN(n20642) );
  AOI22_X1 U23583 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20642), .B1(n20641), 
        .B2(n20640), .ZN(P1_U3163) );
  AND2_X1 U23584 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20643), .ZN(
        P1_U3164) );
  AND2_X1 U23585 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20643), .ZN(
        P1_U3165) );
  AND2_X1 U23586 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20643), .ZN(
        P1_U3166) );
  AND2_X1 U23587 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20643), .ZN(
        P1_U3167) );
  AND2_X1 U23588 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20643), .ZN(
        P1_U3168) );
  AND2_X1 U23589 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20643), .ZN(
        P1_U3169) );
  AND2_X1 U23590 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20643), .ZN(
        P1_U3170) );
  AND2_X1 U23591 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20643), .ZN(
        P1_U3171) );
  AND2_X1 U23592 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20643), .ZN(
        P1_U3172) );
  AND2_X1 U23593 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20643), .ZN(
        P1_U3173) );
  AND2_X1 U23594 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20643), .ZN(
        P1_U3174) );
  AND2_X1 U23595 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20643), .ZN(
        P1_U3175) );
  AND2_X1 U23596 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20643), .ZN(
        P1_U3176) );
  AND2_X1 U23597 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20643), .ZN(
        P1_U3177) );
  AND2_X1 U23598 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20643), .ZN(
        P1_U3178) );
  AND2_X1 U23599 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20643), .ZN(
        P1_U3179) );
  AND2_X1 U23600 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20643), .ZN(
        P1_U3180) );
  AND2_X1 U23601 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20643), .ZN(
        P1_U3181) );
  AND2_X1 U23602 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20643), .ZN(
        P1_U3182) );
  AND2_X1 U23603 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20643), .ZN(
        P1_U3183) );
  AND2_X1 U23604 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20643), .ZN(
        P1_U3184) );
  AND2_X1 U23605 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20643), .ZN(
        P1_U3185) );
  AND2_X1 U23606 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20643), .ZN(P1_U3186) );
  INV_X1 U23607 ( .A(P1_DATAWIDTH_REG_8__SCAN_IN), .ZN(n20966) );
  NOR2_X1 U23608 ( .A1(n20704), .A2(n20966), .ZN(P1_U3187) );
  AND2_X1 U23609 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20643), .ZN(P1_U3188) );
  AND2_X1 U23610 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20643), .ZN(P1_U3189) );
  AND2_X1 U23611 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20643), .ZN(P1_U3190) );
  INV_X1 U23612 ( .A(P1_DATAWIDTH_REG_4__SCAN_IN), .ZN(n20742) );
  NOR2_X1 U23613 ( .A1(n20704), .A2(n20742), .ZN(P1_U3191) );
  AND2_X1 U23614 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20643), .ZN(P1_U3192) );
  AND2_X1 U23615 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20643), .ZN(P1_U3193) );
  AND2_X1 U23616 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20644), .ZN(n20657) );
  OAI21_X1 U23617 ( .B1(P1_STATE_REG_0__SCAN_IN), .B2(n20650), .A(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20645) );
  AOI211_X1 U23618 ( .C1(HOLD), .C2(P1_STATE_REG_1__SCAN_IN), .A(n20646), .B(
        n20645), .ZN(n20647) );
  OAI22_X1 U23619 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20657), .B1(n20715), 
        .B2(n20647), .ZN(P1_U3194) );
  INV_X1 U23620 ( .A(n20648), .ZN(n20651) );
  INV_X1 U23621 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20653) );
  NOR2_X1 U23622 ( .A1(n20655), .A2(n20653), .ZN(n20649) );
  OAI22_X1 U23623 ( .A1(n20651), .A2(n20650), .B1(P1_STATE_REG_2__SCAN_IN), 
        .B2(n20649), .ZN(n20656) );
  OAI211_X1 U23624 ( .C1(NA), .C2(n20718), .A(P1_STATE_REG_1__SCAN_IN), .B(
        n20658), .ZN(n20652) );
  OAI211_X1 U23625 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20653), .A(HOLD), .B(
        n20652), .ZN(n20654) );
  OAI22_X1 U23626 ( .A1(n20657), .A2(n20656), .B1(n20655), .B2(n20654), .ZN(
        P1_U3196) );
  OR2_X1 U23627 ( .A1(n20727), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20685) );
  NOR2_X1 U23628 ( .A1(n20658), .A2(n20727), .ZN(n20693) );
  INV_X1 U23629 ( .A(n20693), .ZN(n20682) );
  AOI222_X1 U23630 ( .A1(n9723), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20713), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n20695), .ZN(n20659) );
  INV_X1 U23631 ( .A(n20659), .ZN(P1_U3197) );
  AOI222_X1 U23632 ( .A1(n20695), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20727), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n9723), .ZN(n20660) );
  INV_X1 U23633 ( .A(n20660), .ZN(P1_U3198) );
  AOI222_X1 U23634 ( .A1(n20695), .A2(P1_REIP_REG_3__SCAN_IN), .B1(
        P1_ADDRESS_REG_2__SCAN_IN), .B2(n20713), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n9723), .ZN(n20661) );
  INV_X1 U23635 ( .A(n20661), .ZN(P1_U3199) );
  AOI222_X1 U23636 ( .A1(n20695), .A2(P1_REIP_REG_4__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20713), .C1(P1_REIP_REG_5__SCAN_IN), 
        .C2(n9723), .ZN(n20662) );
  INV_X1 U23637 ( .A(n20662), .ZN(P1_U3200) );
  AOI222_X1 U23638 ( .A1(n20695), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20713), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n9723), .ZN(n20663) );
  INV_X1 U23639 ( .A(n20663), .ZN(P1_U3201) );
  AOI222_X1 U23640 ( .A1(n20695), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20713), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n9723), .ZN(n20664) );
  INV_X1 U23641 ( .A(n20664), .ZN(P1_U3202) );
  AOI222_X1 U23642 ( .A1(n20695), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20713), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n9723), .ZN(n20665) );
  INV_X1 U23643 ( .A(n20665), .ZN(P1_U3203) );
  AOI22_X1 U23644 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n20727), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n9723), .ZN(n20666) );
  OAI21_X1 U23645 ( .B1(n20908), .B2(n20682), .A(n20666), .ZN(P1_U3204) );
  AOI22_X1 U23646 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(n20727), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20693), .ZN(n20667) );
  OAI21_X1 U23647 ( .B1(n20668), .B2(n20685), .A(n20667), .ZN(P1_U3205) );
  AOI222_X1 U23648 ( .A1(n9723), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20713), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20695), .ZN(n20669) );
  INV_X1 U23649 ( .A(n20669), .ZN(P1_U3206) );
  AOI222_X1 U23650 ( .A1(n9723), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20713), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n20695), .ZN(n20670) );
  INV_X1 U23651 ( .A(n20670), .ZN(P1_U3207) );
  AOI222_X1 U23652 ( .A1(n9723), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20713), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20695), .ZN(n20671) );
  INV_X1 U23653 ( .A(n20671), .ZN(P1_U3208) );
  AOI22_X1 U23654 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20727), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n9723), .ZN(n20672) );
  OAI21_X1 U23655 ( .B1(n20819), .B2(n20682), .A(n20672), .ZN(P1_U3209) );
  AOI22_X1 U23656 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20727), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20695), .ZN(n20673) );
  OAI21_X1 U23657 ( .B1(n14539), .B2(n20685), .A(n20673), .ZN(P1_U3210) );
  AOI22_X1 U23658 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(n20727), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n9723), .ZN(n20674) );
  OAI21_X1 U23659 ( .B1(n14539), .B2(n20682), .A(n20674), .ZN(P1_U3211) );
  AOI22_X1 U23660 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20727), .B1(
        P1_REIP_REG_16__SCAN_IN), .B2(n20693), .ZN(n20675) );
  OAI21_X1 U23661 ( .B1(n20676), .B2(n20685), .A(n20675), .ZN(P1_U3212) );
  AOI222_X1 U23662 ( .A1(n9723), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n20713), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20695), .ZN(n20677) );
  INV_X1 U23663 ( .A(n20677), .ZN(P1_U3213) );
  AOI222_X1 U23664 ( .A1(n20693), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20713), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n9723), .ZN(n20678) );
  INV_X1 U23665 ( .A(n20678), .ZN(P1_U3214) );
  AOI222_X1 U23666 ( .A1(n9723), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20713), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20695), .ZN(n20679) );
  INV_X1 U23667 ( .A(n20679), .ZN(P1_U3215) );
  AOI222_X1 U23668 ( .A1(n20693), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20713), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n9723), .ZN(n20680) );
  INV_X1 U23669 ( .A(n20680), .ZN(P1_U3216) );
  AOI22_X1 U23670 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(n20727), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(n9723), .ZN(n20681) );
  OAI21_X1 U23671 ( .B1(n20683), .B2(n20682), .A(n20681), .ZN(P1_U3217) );
  AOI22_X1 U23672 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20727), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(n20693), .ZN(n20684) );
  OAI21_X1 U23673 ( .B1(n20686), .B2(n20685), .A(n20684), .ZN(P1_U3218) );
  AOI222_X1 U23674 ( .A1(n20693), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20713), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n9723), .ZN(n20687) );
  INV_X1 U23675 ( .A(n20687), .ZN(P1_U3219) );
  AOI222_X1 U23676 ( .A1(n20693), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20713), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n9723), .ZN(n20688) );
  INV_X1 U23677 ( .A(n20688), .ZN(P1_U3220) );
  AOI222_X1 U23678 ( .A1(n20693), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20727), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n9723), .ZN(n20689) );
  INV_X1 U23679 ( .A(n20689), .ZN(P1_U3221) );
  AOI222_X1 U23680 ( .A1(n20695), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20713), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n9723), .ZN(n20690) );
  INV_X1 U23681 ( .A(n20690), .ZN(P1_U3222) );
  AOI222_X1 U23682 ( .A1(n20695), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20713), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n9723), .ZN(n20691) );
  INV_X1 U23683 ( .A(n20691), .ZN(P1_U3223) );
  AOI222_X1 U23684 ( .A1(n20695), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20713), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n9723), .ZN(n20692) );
  INV_X1 U23685 ( .A(n20692), .ZN(P1_U3224) );
  AOI222_X1 U23686 ( .A1(n20693), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20713), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n9723), .ZN(n20694) );
  INV_X1 U23687 ( .A(n20694), .ZN(P1_U3225) );
  AOI222_X1 U23688 ( .A1(n20695), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20713), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n9723), .ZN(n20696) );
  INV_X1 U23689 ( .A(n20696), .ZN(P1_U3226) );
  OAI22_X1 U23690 ( .A1(n20713), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20715), .ZN(n20697) );
  INV_X1 U23691 ( .A(n20697), .ZN(P1_U3458) );
  OAI22_X1 U23692 ( .A1(n20727), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20715), .ZN(n20698) );
  INV_X1 U23693 ( .A(n20698), .ZN(P1_U3459) );
  OAI22_X1 U23694 ( .A1(n20727), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20715), .ZN(n20699) );
  INV_X1 U23695 ( .A(n20699), .ZN(P1_U3460) );
  OAI22_X1 U23696 ( .A1(n20727), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20715), .ZN(n20700) );
  INV_X1 U23697 ( .A(n20700), .ZN(P1_U3461) );
  OAI21_X1 U23698 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20704), .A(n20702), 
        .ZN(n20701) );
  INV_X1 U23699 ( .A(n20701), .ZN(P1_U3464) );
  OAI21_X1 U23700 ( .B1(n20704), .B2(n20703), .A(n20702), .ZN(P1_U3465) );
  AOI21_X1 U23701 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20706) );
  AOI22_X1 U23702 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20706), .B2(n20705), .ZN(n20708) );
  INV_X1 U23703 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20707) );
  AOI22_X1 U23704 ( .A1(n20709), .A2(n20708), .B1(n20707), .B2(n20712), .ZN(
        P1_U3481) );
  INV_X1 U23705 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20898) );
  NOR2_X1 U23706 ( .A1(n20712), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n20710) );
  AOI22_X1 U23707 ( .A1(n20898), .A2(n20712), .B1(n20711), .B2(n20710), .ZN(
        P1_U3482) );
  AOI22_X1 U23708 ( .A1(n20715), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20714), 
        .B2(n20713), .ZN(P1_U3483) );
  AOI211_X1 U23709 ( .C1(n20719), .C2(n20718), .A(n20717), .B(n20716), .ZN(
        n20726) );
  OAI211_X1 U23710 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20721), .A(n20720), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20723) );
  AOI21_X1 U23711 ( .B1(n20723), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n20722), 
        .ZN(n20725) );
  NAND2_X1 U23712 ( .A1(n20726), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20724) );
  OAI21_X1 U23713 ( .B1(n20726), .B2(n20725), .A(n20724), .ZN(P1_U3485) );
  MUX2_X1 U23714 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n20727), .Z(P1_U3486) );
  INV_X1 U23715 ( .A(n20728), .ZN(n20732) );
  OAI22_X1 U23716 ( .A1(n20732), .A2(n20731), .B1(n20730), .B2(n20729), .ZN(
        n20738) );
  OAI22_X1 U23717 ( .A1(n20736), .A2(n20735), .B1(n20734), .B2(n20733), .ZN(
        n20737) );
  AOI211_X1 U23718 ( .C1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .C2(n20739), .A(
        n20738), .B(n20737), .ZN(n20986) );
  INV_X1 U23719 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n20741) );
  AOI22_X1 U23720 ( .A1(n20742), .A2(keyinput95), .B1(keyinput52), .B2(n20741), 
        .ZN(n20740) );
  OAI221_X1 U23721 ( .B1(n20742), .B2(keyinput95), .C1(n20741), .C2(keyinput52), .A(n20740), .ZN(n20746) );
  XOR2_X1 U23722 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B(keyinput78), .Z(
        n20745) );
  XNOR2_X1 U23723 ( .A(n20743), .B(keyinput49), .ZN(n20744) );
  OR3_X1 U23724 ( .A1(n20746), .A2(n20745), .A3(n20744), .ZN(n20755) );
  AOI22_X1 U23725 ( .A1(n20749), .A2(keyinput37), .B1(keyinput92), .B2(n20748), 
        .ZN(n20747) );
  OAI221_X1 U23726 ( .B1(n20749), .B2(keyinput37), .C1(n20748), .C2(keyinput92), .A(n20747), .ZN(n20754) );
  AOI22_X1 U23727 ( .A1(n20752), .A2(keyinput80), .B1(keyinput19), .B2(n20751), 
        .ZN(n20750) );
  OAI221_X1 U23728 ( .B1(n20752), .B2(keyinput80), .C1(n20751), .C2(keyinput19), .A(n20750), .ZN(n20753) );
  NOR3_X1 U23729 ( .A1(n20755), .A2(n20754), .A3(n20753), .ZN(n20801) );
  AOI22_X1 U23730 ( .A1(n11353), .A2(keyinput16), .B1(keyinput36), .B2(n20757), 
        .ZN(n20756) );
  OAI221_X1 U23731 ( .B1(n11353), .B2(keyinput16), .C1(n20757), .C2(keyinput36), .A(n20756), .ZN(n20768) );
  AOI22_X1 U23732 ( .A1(n20760), .A2(keyinput108), .B1(keyinput28), .B2(n20759), .ZN(n20758) );
  OAI221_X1 U23733 ( .B1(n20760), .B2(keyinput108), .C1(n20759), .C2(
        keyinput28), .A(n20758), .ZN(n20767) );
  INV_X1 U23734 ( .A(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n20762) );
  AOI22_X1 U23735 ( .A1(n21022), .A2(keyinput64), .B1(n20762), .B2(keyinput11), 
        .ZN(n20761) );
  OAI221_X1 U23736 ( .B1(n21022), .B2(keyinput64), .C1(n20762), .C2(keyinput11), .A(n20761), .ZN(n20766) );
  XNOR2_X1 U23737 ( .A(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B(keyinput17), .ZN(
        n20764) );
  XNOR2_X1 U23738 ( .A(keyinput87), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), 
        .ZN(n20763) );
  NAND2_X1 U23739 ( .A1(n20764), .A2(n20763), .ZN(n20765) );
  NOR4_X1 U23740 ( .A1(n20768), .A2(n20767), .A3(n20766), .A4(n20765), .ZN(
        n20800) );
  INV_X1 U23741 ( .A(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n20771) );
  AOI22_X1 U23742 ( .A1(n20771), .A2(keyinput44), .B1(keyinput123), .B2(n20770), .ZN(n20769) );
  OAI221_X1 U23743 ( .B1(n20771), .B2(keyinput44), .C1(n20770), .C2(
        keyinput123), .A(n20769), .ZN(n20781) );
  AOI22_X1 U23744 ( .A1(n21021), .A2(keyinput105), .B1(keyinput10), .B2(n20773), .ZN(n20772) );
  OAI221_X1 U23745 ( .B1(n21021), .B2(keyinput105), .C1(n20773), .C2(
        keyinput10), .A(n20772), .ZN(n20780) );
  AOI22_X1 U23746 ( .A1(n21026), .A2(keyinput110), .B1(n20775), .B2(keyinput45), .ZN(n20774) );
  OAI221_X1 U23747 ( .B1(n21026), .B2(keyinput110), .C1(n20775), .C2(
        keyinput45), .A(n20774), .ZN(n20779) );
  INV_X1 U23748 ( .A(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n20777) );
  INV_X1 U23749 ( .A(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n20993) );
  AOI22_X1 U23750 ( .A1(n20777), .A2(keyinput85), .B1(n20993), .B2(keyinput75), 
        .ZN(n20776) );
  OAI221_X1 U23751 ( .B1(n20777), .B2(keyinput85), .C1(n20993), .C2(keyinput75), .A(n20776), .ZN(n20778) );
  NOR4_X1 U23752 ( .A1(n20781), .A2(n20780), .A3(n20779), .A4(n20778), .ZN(
        n20799) );
  AOI22_X1 U23753 ( .A1(n20784), .A2(keyinput101), .B1(keyinput102), .B2(
        n20783), .ZN(n20782) );
  OAI221_X1 U23754 ( .B1(n20784), .B2(keyinput101), .C1(n20783), .C2(
        keyinput102), .A(n20782), .ZN(n20797) );
  AOI22_X1 U23755 ( .A1(n20787), .A2(keyinput2), .B1(n20786), .B2(keyinput53), 
        .ZN(n20785) );
  OAI221_X1 U23756 ( .B1(n20787), .B2(keyinput2), .C1(n20786), .C2(keyinput53), 
        .A(n20785), .ZN(n20796) );
  AOI22_X1 U23757 ( .A1(n20790), .A2(keyinput58), .B1(n20789), .B2(keyinput50), 
        .ZN(n20788) );
  OAI221_X1 U23758 ( .B1(n20790), .B2(keyinput58), .C1(n20789), .C2(keyinput50), .A(n20788), .ZN(n20795) );
  INV_X1 U23759 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n20793) );
  AOI22_X1 U23760 ( .A1(n20793), .A2(keyinput1), .B1(n20792), .B2(keyinput7), 
        .ZN(n20791) );
  OAI221_X1 U23761 ( .B1(n20793), .B2(keyinput1), .C1(n20792), .C2(keyinput7), 
        .A(n20791), .ZN(n20794) );
  NOR4_X1 U23762 ( .A1(n20797), .A2(n20796), .A3(n20795), .A4(n20794), .ZN(
        n20798) );
  NAND4_X1 U23763 ( .A1(n20801), .A2(n20800), .A3(n20799), .A4(n20798), .ZN(
        n20984) );
  AOI22_X1 U23764 ( .A1(n20804), .A2(keyinput54), .B1(n20803), .B2(keyinput20), 
        .ZN(n20802) );
  OAI221_X1 U23765 ( .B1(n20804), .B2(keyinput54), .C1(n20803), .C2(keyinput20), .A(n20802), .ZN(n20817) );
  INV_X1 U23766 ( .A(DATAI_6_), .ZN(n20807) );
  AOI22_X1 U23767 ( .A1(n20807), .A2(keyinput109), .B1(keyinput104), .B2(
        n20806), .ZN(n20805) );
  OAI221_X1 U23768 ( .B1(n20807), .B2(keyinput109), .C1(n20806), .C2(
        keyinput104), .A(n20805), .ZN(n20816) );
  INV_X1 U23769 ( .A(DATAI_30_), .ZN(n20809) );
  AOI22_X1 U23770 ( .A1(n20810), .A2(keyinput51), .B1(keyinput48), .B2(n20809), 
        .ZN(n20808) );
  OAI221_X1 U23771 ( .B1(n20810), .B2(keyinput51), .C1(n20809), .C2(keyinput48), .A(n20808), .ZN(n20815) );
  AOI22_X1 U23772 ( .A1(n20813), .A2(keyinput79), .B1(keyinput35), .B2(n20812), 
        .ZN(n20811) );
  OAI221_X1 U23773 ( .B1(n20813), .B2(keyinput79), .C1(n20812), .C2(keyinput35), .A(n20811), .ZN(n20814) );
  NOR4_X1 U23774 ( .A1(n20817), .A2(n20816), .A3(n20815), .A4(n20814), .ZN(
        n20862) );
  AOI22_X1 U23775 ( .A1(n20820), .A2(keyinput124), .B1(keyinput22), .B2(n20819), .ZN(n20818) );
  OAI221_X1 U23776 ( .B1(n20820), .B2(keyinput124), .C1(n20819), .C2(
        keyinput22), .A(n20818), .ZN(n20832) );
  AOI22_X1 U23777 ( .A1(n20823), .A2(keyinput120), .B1(n20822), .B2(keyinput77), .ZN(n20821) );
  OAI221_X1 U23778 ( .B1(n20823), .B2(keyinput120), .C1(n20822), .C2(
        keyinput77), .A(n20821), .ZN(n20831) );
  AOI22_X1 U23779 ( .A1(n20826), .A2(keyinput82), .B1(n20825), .B2(keyinput67), 
        .ZN(n20824) );
  OAI221_X1 U23780 ( .B1(n20826), .B2(keyinput82), .C1(n20825), .C2(keyinput67), .A(n20824), .ZN(n20830) );
  INV_X1 U23781 ( .A(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n20990) );
  AOI22_X1 U23782 ( .A1(n20828), .A2(keyinput71), .B1(n20990), .B2(keyinput107), .ZN(n20827) );
  OAI221_X1 U23783 ( .B1(n20828), .B2(keyinput71), .C1(n20990), .C2(
        keyinput107), .A(n20827), .ZN(n20829) );
  NOR4_X1 U23784 ( .A1(n20832), .A2(n20831), .A3(n20830), .A4(n20829), .ZN(
        n20861) );
  AOI22_X1 U23785 ( .A1(n20835), .A2(keyinput72), .B1(n20834), .B2(keyinput113), .ZN(n20833) );
  OAI221_X1 U23786 ( .B1(n20835), .B2(keyinput72), .C1(n20834), .C2(
        keyinput113), .A(n20833), .ZN(n20846) );
  INV_X1 U23787 ( .A(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n20838) );
  AOI22_X1 U23788 ( .A1(n20838), .A2(keyinput43), .B1(keyinput114), .B2(n20837), .ZN(n20836) );
  OAI221_X1 U23789 ( .B1(n20838), .B2(keyinput43), .C1(n20837), .C2(
        keyinput114), .A(n20836), .ZN(n20845) );
  AOI22_X1 U23790 ( .A1(n20840), .A2(keyinput12), .B1(n21011), .B2(keyinput23), 
        .ZN(n20839) );
  OAI221_X1 U23791 ( .B1(n20840), .B2(keyinput12), .C1(n21011), .C2(keyinput23), .A(n20839), .ZN(n20844) );
  INV_X1 U23792 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n21024) );
  INV_X1 U23793 ( .A(DATAI_28_), .ZN(n20842) );
  AOI22_X1 U23794 ( .A1(n21024), .A2(keyinput86), .B1(n20842), .B2(keyinput31), 
        .ZN(n20841) );
  OAI221_X1 U23795 ( .B1(n21024), .B2(keyinput86), .C1(n20842), .C2(keyinput31), .A(n20841), .ZN(n20843) );
  NOR4_X1 U23796 ( .A1(n20846), .A2(n20845), .A3(n20844), .A4(n20843), .ZN(
        n20860) );
  AOI22_X1 U23797 ( .A1(n20848), .A2(keyinput6), .B1(n12092), .B2(keyinput57), 
        .ZN(n20847) );
  OAI221_X1 U23798 ( .B1(n20848), .B2(keyinput6), .C1(n12092), .C2(keyinput57), 
        .A(n20847), .ZN(n20858) );
  AOI22_X1 U23799 ( .A1(n20851), .A2(keyinput30), .B1(keyinput56), .B2(n20850), 
        .ZN(n20849) );
  OAI221_X1 U23800 ( .B1(n20851), .B2(keyinput30), .C1(n20850), .C2(keyinput56), .A(n20849), .ZN(n20857) );
  AOI22_X1 U23801 ( .A1(n20853), .A2(keyinput70), .B1(keyinput65), .B2(n14366), 
        .ZN(n20852) );
  OAI221_X1 U23802 ( .B1(n20853), .B2(keyinput70), .C1(n14366), .C2(keyinput65), .A(n20852), .ZN(n20856) );
  AOI22_X1 U23803 ( .A1(n21023), .A2(keyinput88), .B1(n12527), .B2(keyinput42), 
        .ZN(n20854) );
  OAI221_X1 U23804 ( .B1(n21023), .B2(keyinput88), .C1(n12527), .C2(keyinput42), .A(n20854), .ZN(n20855) );
  NOR4_X1 U23805 ( .A1(n20858), .A2(n20857), .A3(n20856), .A4(n20855), .ZN(
        n20859) );
  NAND4_X1 U23806 ( .A1(n20862), .A2(n20861), .A3(n20860), .A4(n20859), .ZN(
        n20983) );
  AOI22_X1 U23807 ( .A1(n20865), .A2(keyinput96), .B1(n20864), .B2(keyinput15), 
        .ZN(n20863) );
  OAI221_X1 U23808 ( .B1(n20865), .B2(keyinput96), .C1(n20864), .C2(keyinput15), .A(n20863), .ZN(n20877) );
  INV_X1 U23809 ( .A(DATAI_26_), .ZN(n20867) );
  AOI22_X1 U23810 ( .A1(n20868), .A2(keyinput24), .B1(keyinput116), .B2(n20867), .ZN(n20866) );
  OAI221_X1 U23811 ( .B1(n20868), .B2(keyinput24), .C1(n20867), .C2(
        keyinput116), .A(n20866), .ZN(n20876) );
  AOI22_X1 U23812 ( .A1(n14165), .A2(keyinput84), .B1(n20870), .B2(keyinput103), .ZN(n20869) );
  OAI221_X1 U23813 ( .B1(n14165), .B2(keyinput84), .C1(n20870), .C2(
        keyinput103), .A(n20869), .ZN(n20875) );
  XOR2_X1 U23814 ( .A(n20871), .B(keyinput27), .Z(n20873) );
  XNOR2_X1 U23815 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(keyinput76), 
        .ZN(n20872) );
  NAND2_X1 U23816 ( .A1(n20873), .A2(n20872), .ZN(n20874) );
  NOR4_X1 U23817 ( .A1(n20877), .A2(n20876), .A3(n20875), .A4(n20874), .ZN(
        n20920) );
  INV_X1 U23818 ( .A(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n20994) );
  AOI22_X1 U23819 ( .A1(n20994), .A2(keyinput5), .B1(keyinput126), .B2(n21020), 
        .ZN(n20878) );
  OAI221_X1 U23820 ( .B1(n20994), .B2(keyinput5), .C1(n21020), .C2(keyinput126), .A(n20878), .ZN(n20891) );
  AOI22_X1 U23821 ( .A1(n20881), .A2(keyinput73), .B1(keyinput69), .B2(n20880), 
        .ZN(n20879) );
  OAI221_X1 U23822 ( .B1(n20881), .B2(keyinput73), .C1(n20880), .C2(keyinput69), .A(n20879), .ZN(n20890) );
  AOI22_X1 U23823 ( .A1(n20884), .A2(keyinput125), .B1(n20883), .B2(keyinput41), .ZN(n20882) );
  OAI221_X1 U23824 ( .B1(n20884), .B2(keyinput125), .C1(n20883), .C2(
        keyinput41), .A(n20882), .ZN(n20889) );
  XOR2_X1 U23825 ( .A(n20885), .B(keyinput34), .Z(n20887) );
  XNOR2_X1 U23826 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B(keyinput8), .ZN(
        n20886) );
  NAND2_X1 U23827 ( .A1(n20887), .A2(n20886), .ZN(n20888) );
  NOR4_X1 U23828 ( .A1(n20891), .A2(n20890), .A3(n20889), .A4(n20888), .ZN(
        n20919) );
  INV_X1 U23829 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n20893) );
  AOI22_X1 U23830 ( .A1(n20894), .A2(keyinput18), .B1(n20893), .B2(keyinput29), 
        .ZN(n20892) );
  OAI221_X1 U23831 ( .B1(n20894), .B2(keyinput18), .C1(n20893), .C2(keyinput29), .A(n20892), .ZN(n20903) );
  AOI22_X1 U23832 ( .A1(n21025), .A2(keyinput46), .B1(n21028), .B2(keyinput122), .ZN(n20895) );
  OAI221_X1 U23833 ( .B1(n21025), .B2(keyinput46), .C1(n21028), .C2(
        keyinput122), .A(n20895), .ZN(n20902) );
  AOI22_X1 U23834 ( .A1(n9999), .A2(keyinput39), .B1(n21010), .B2(keyinput121), 
        .ZN(n20896) );
  OAI221_X1 U23835 ( .B1(n9999), .B2(keyinput39), .C1(n21010), .C2(keyinput121), .A(n20896), .ZN(n20901) );
  INV_X1 U23836 ( .A(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n20899) );
  AOI22_X1 U23837 ( .A1(n20899), .A2(keyinput59), .B1(keyinput9), .B2(n20898), 
        .ZN(n20897) );
  OAI221_X1 U23838 ( .B1(n20899), .B2(keyinput59), .C1(n20898), .C2(keyinput9), 
        .A(n20897), .ZN(n20900) );
  NOR4_X1 U23839 ( .A1(n20903), .A2(n20902), .A3(n20901), .A4(n20900), .ZN(
        n20918) );
  AOI22_X1 U23840 ( .A1(n20906), .A2(keyinput3), .B1(n20905), .B2(keyinput66), 
        .ZN(n20904) );
  OAI221_X1 U23841 ( .B1(n20906), .B2(keyinput3), .C1(n20905), .C2(keyinput66), 
        .A(n20904), .ZN(n20916) );
  INV_X1 U23842 ( .A(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n20987) );
  AOI22_X1 U23843 ( .A1(n20908), .A2(keyinput74), .B1(n20987), .B2(keyinput112), .ZN(n20907) );
  OAI221_X1 U23844 ( .B1(n20908), .B2(keyinput74), .C1(n20987), .C2(
        keyinput112), .A(n20907), .ZN(n20915) );
  AOI22_X1 U23845 ( .A1(n20992), .A2(keyinput111), .B1(n20910), .B2(keyinput63), .ZN(n20909) );
  OAI221_X1 U23846 ( .B1(n20992), .B2(keyinput111), .C1(n20910), .C2(
        keyinput63), .A(n20909), .ZN(n20914) );
  INV_X1 U23847 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n20912) );
  AOI22_X1 U23848 ( .A1(n20912), .A2(keyinput117), .B1(n10713), .B2(keyinput62), .ZN(n20911) );
  OAI221_X1 U23849 ( .B1(n20912), .B2(keyinput117), .C1(n10713), .C2(
        keyinput62), .A(n20911), .ZN(n20913) );
  NOR4_X1 U23850 ( .A1(n20916), .A2(n20915), .A3(n20914), .A4(n20913), .ZN(
        n20917) );
  NAND4_X1 U23851 ( .A1(n20920), .A2(n20919), .A3(n20918), .A4(n20917), .ZN(
        n20982) );
  AOI22_X1 U23852 ( .A1(n20922), .A2(keyinput115), .B1(n13580), .B2(keyinput60), .ZN(n20921) );
  OAI221_X1 U23853 ( .B1(n20922), .B2(keyinput115), .C1(n13580), .C2(
        keyinput60), .A(n20921), .ZN(n20934) );
  AOI22_X1 U23854 ( .A1(n20925), .A2(keyinput100), .B1(n20924), .B2(keyinput4), 
        .ZN(n20923) );
  OAI221_X1 U23855 ( .B1(n20925), .B2(keyinput100), .C1(n20924), .C2(keyinput4), .A(n20923), .ZN(n20933) );
  AOI22_X1 U23856 ( .A1(n21009), .A2(keyinput106), .B1(n20927), .B2(keyinput97), .ZN(n20926) );
  OAI221_X1 U23857 ( .B1(n21009), .B2(keyinput106), .C1(n20927), .C2(
        keyinput97), .A(n20926), .ZN(n20932) );
  INV_X1 U23858 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n20929) );
  AOI22_X1 U23859 ( .A1(n20930), .A2(keyinput13), .B1(n20929), .B2(keyinput99), 
        .ZN(n20928) );
  OAI221_X1 U23860 ( .B1(n20930), .B2(keyinput13), .C1(n20929), .C2(keyinput99), .A(n20928), .ZN(n20931) );
  NOR4_X1 U23861 ( .A1(n20934), .A2(n20933), .A3(n20932), .A4(n20931), .ZN(
        n20980) );
  INV_X1 U23862 ( .A(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n20936) );
  AOI22_X1 U23863 ( .A1(n11941), .A2(keyinput68), .B1(keyinput55), .B2(n20936), 
        .ZN(n20935) );
  OAI221_X1 U23864 ( .B1(n11941), .B2(keyinput68), .C1(n20936), .C2(keyinput55), .A(n20935), .ZN(n20948) );
  AOI22_X1 U23865 ( .A1(n20939), .A2(keyinput21), .B1(n20938), .B2(keyinput83), 
        .ZN(n20937) );
  OAI221_X1 U23866 ( .B1(n20939), .B2(keyinput21), .C1(n20938), .C2(keyinput83), .A(n20937), .ZN(n20947) );
  AOI22_X1 U23867 ( .A1(n20942), .A2(keyinput33), .B1(n20941), .B2(keyinput40), 
        .ZN(n20940) );
  OAI221_X1 U23868 ( .B1(n20942), .B2(keyinput33), .C1(n20941), .C2(keyinput40), .A(n20940), .ZN(n20946) );
  INV_X1 U23869 ( .A(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n20944) );
  AOI22_X1 U23870 ( .A1(n20944), .A2(keyinput47), .B1(keyinput93), .B2(n21008), 
        .ZN(n20943) );
  OAI221_X1 U23871 ( .B1(n20944), .B2(keyinput47), .C1(n21008), .C2(keyinput93), .A(n20943), .ZN(n20945) );
  NOR4_X1 U23872 ( .A1(n20948), .A2(n20947), .A3(n20946), .A4(n20945), .ZN(
        n20979) );
  AOI22_X1 U23873 ( .A1(n20951), .A2(keyinput118), .B1(keyinput32), .B2(n20950), .ZN(n20949) );
  OAI221_X1 U23874 ( .B1(n20951), .B2(keyinput118), .C1(n20950), .C2(
        keyinput32), .A(n20949), .ZN(n20963) );
  INV_X1 U23875 ( .A(DATAI_4_), .ZN(n20953) );
  AOI22_X1 U23876 ( .A1(n20954), .A2(keyinput127), .B1(n20953), .B2(keyinput98), .ZN(n20952) );
  OAI221_X1 U23877 ( .B1(n20954), .B2(keyinput127), .C1(n20953), .C2(
        keyinput98), .A(n20952), .ZN(n20962) );
  AOI22_X1 U23878 ( .A1(n20957), .A2(keyinput38), .B1(keyinput14), .B2(n20956), 
        .ZN(n20955) );
  OAI221_X1 U23879 ( .B1(n20957), .B2(keyinput38), .C1(n20956), .C2(keyinput14), .A(n20955), .ZN(n20961) );
  AOI22_X1 U23880 ( .A1(n20959), .A2(keyinput90), .B1(keyinput89), .B2(n20991), 
        .ZN(n20958) );
  OAI221_X1 U23881 ( .B1(n20959), .B2(keyinput90), .C1(n20991), .C2(keyinput89), .A(n20958), .ZN(n20960) );
  NOR4_X1 U23882 ( .A1(n20963), .A2(n20962), .A3(n20961), .A4(n20960), .ZN(
        n20978) );
  AOI22_X1 U23883 ( .A1(n20966), .A2(keyinput91), .B1(n20965), .B2(keyinput25), 
        .ZN(n20964) );
  OAI221_X1 U23884 ( .B1(n20966), .B2(keyinput91), .C1(n20965), .C2(keyinput25), .A(n20964), .ZN(n20976) );
  AOI22_X1 U23885 ( .A1(n21027), .A2(keyinput81), .B1(n10499), .B2(keyinput119), .ZN(n20967) );
  OAI221_X1 U23886 ( .B1(n21027), .B2(keyinput81), .C1(n10499), .C2(
        keyinput119), .A(n20967), .ZN(n20975) );
  AOI22_X1 U23887 ( .A1(n20969), .A2(keyinput94), .B1(keyinput0), .B2(n11852), 
        .ZN(n20968) );
  OAI221_X1 U23888 ( .B1(n20969), .B2(keyinput94), .C1(n11852), .C2(keyinput0), 
        .A(n20968), .ZN(n20974) );
  AOI22_X1 U23889 ( .A1(n20972), .A2(keyinput26), .B1(n20971), .B2(keyinput61), 
        .ZN(n20970) );
  OAI221_X1 U23890 ( .B1(n20972), .B2(keyinput26), .C1(n20971), .C2(keyinput61), .A(n20970), .ZN(n20973) );
  NOR4_X1 U23891 ( .A1(n20976), .A2(n20975), .A3(n20974), .A4(n20973), .ZN(
        n20977) );
  NAND4_X1 U23892 ( .A1(n20980), .A2(n20979), .A3(n20978), .A4(n20977), .ZN(
        n20981) );
  NOR4_X1 U23893 ( .A1(n20984), .A2(n20983), .A3(n20982), .A4(n20981), .ZN(
        n20985) );
  XNOR2_X1 U23894 ( .A(n20986), .B(n20985), .ZN(n21050) );
  NAND4_X1 U23895 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20989), .A3(
        n20988), .A4(n20987), .ZN(n21003) );
  NOR4_X1 U23896 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_5__2__SCAN_IN), .A3(n20991), .A4(n20990), .ZN(n21001)
         );
  NOR4_X1 U23897 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_10__1__SCAN_IN), .A3(n20993), .A4(n20992), .ZN(n21000) );
  NAND4_X1 U23898 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_14__7__SCAN_IN), .A3(P3_EBX_REG_26__SCAN_IN), .A4(
        P3_REIP_REG_5__SCAN_IN), .ZN(n20998) );
  NAND4_X1 U23899 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A3(
        P3_INSTQUEUE_REG_9__7__SCAN_IN), .A4(n20994), .ZN(n20997) );
  NAND4_X1 U23900 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_15__3__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A4(BUF2_REG_1__SCAN_IN), .ZN(
        n20996) );
  NAND4_X1 U23901 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_STATE_REG_0__SCAN_IN), .A3(BUF2_REG_2__SCAN_IN), .A4(
        P3_EBX_REG_15__SCAN_IN), .ZN(n20995) );
  NOR4_X1 U23902 ( .A1(n20998), .A2(n20997), .A3(n20996), .A4(n20995), .ZN(
        n20999) );
  NAND3_X1 U23903 ( .A1(n21001), .A2(n21000), .A3(n20999), .ZN(n21002) );
  NOR4_X1 U23904 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(
        P1_INSTQUEUE_REG_7__7__SCAN_IN), .A3(n21003), .A4(n21002), .ZN(n21048)
         );
  NAND4_X1 U23905 ( .A1(P1_EAX_REG_2__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_UWORD_REG_1__SCAN_IN), .A4(
        P2_LWORD_REG_10__SCAN_IN), .ZN(n21007) );
  NAND4_X1 U23906 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_8__SCAN_IN), .A3(P3_ADDRESS_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_4__SCAN_IN), .ZN(n21006) );
  NAND4_X1 U23907 ( .A1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A3(P2_UWORD_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_5__SCAN_IN), .ZN(n21005) );
  NAND4_X1 U23908 ( .A1(P2_EAX_REG_25__SCAN_IN), .A2(P1_EBX_REG_19__SCAN_IN), 
        .A3(P2_LWORD_REG_4__SCAN_IN), .A4(P2_LWORD_REG_9__SCAN_IN), .ZN(n21004) );
  NOR4_X1 U23909 ( .A1(n21007), .A2(n21006), .A3(n21005), .A4(n21004), .ZN(
        n21047) );
  NAND4_X1 U23910 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_REIP_REG_13__SCAN_IN), .A3(DATAI_30_), .A4(P3_EAX_REG_0__SCAN_IN), 
        .ZN(n21015) );
  NAND4_X1 U23911 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_8__5__SCAN_IN), .A3(BUF2_REG_27__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n21014) );
  NAND4_X1 U23912 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(
        P1_DATAO_REG_16__SCAN_IN), .A3(n21009), .A4(n21008), .ZN(n21013) );
  NAND4_X1 U23913 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(DATAI_26_), .A3(
        n21011), .A4(n21010), .ZN(n21012) );
  NOR4_X1 U23914 ( .A1(n21015), .A2(n21014), .A3(n21013), .A4(n21012), .ZN(
        n21046) );
  NOR4_X1 U23915 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_EAX_REG_4__SCAN_IN), .A3(P1_EBX_REG_29__SCAN_IN), .A4(
        BUF1_REG_0__SCAN_IN), .ZN(n21019) );
  NOR4_X1 U23916 ( .A1(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A3(P1_EAX_REG_0__SCAN_IN), .A4(
        DATAI_4_), .ZN(n21018) );
  NOR4_X1 U23917 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(P3_REIP_REG_8__SCAN_IN), .A4(
        P3_UWORD_REG_5__SCAN_IN), .ZN(n21017) );
  NOR4_X1 U23918 ( .A1(P2_EBX_REG_12__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_8__5__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), 
        .A4(P3_DATAWIDTH_REG_12__SCAN_IN), .ZN(n21016) );
  NAND4_X1 U23919 ( .A1(n21019), .A2(n21018), .A3(n21017), .A4(n21016), .ZN(
        n21044) );
  NOR4_X1 U23920 ( .A1(n21023), .A2(n21022), .A3(n21021), .A4(n21020), .ZN(
        n21032) );
  NOR4_X1 U23921 ( .A1(n21027), .A2(n21026), .A3(n21025), .A4(n21024), .ZN(
        n21031) );
  NOR4_X1 U23922 ( .A1(DATAI_6_), .A2(P3_DATAO_REG_2__SCAN_IN), .A3(
        P3_DATAO_REG_7__SCAN_IN), .A4(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(
        n21030) );
  NOR4_X1 U23923 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(P3_ADDRESS_REG_8__SCAN_IN), .A3(P3_DATAO_REG_0__SCAN_IN), .A4(n21028), .ZN(n21029) );
  NAND4_X1 U23924 ( .A1(n21032), .A2(n21031), .A3(n21030), .A4(n21029), .ZN(
        n21043) );
  NOR4_X1 U23925 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(
        P2_EBX_REG_19__SCAN_IN), .A3(P2_EBX_REG_23__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n21036) );
  NOR4_X1 U23926 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_13__3__SCAN_IN), .A3(P2_INSTQUEUE_REG_3__2__SCAN_IN), 
        .A4(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n21035) );
  NOR4_X1 U23927 ( .A1(BUF1_REG_30__SCAN_IN), .A2(P1_EAX_REG_30__SCAN_IN), 
        .A3(P1_REIP_REG_11__SCAN_IN), .A4(DATAI_28_), .ZN(n21034) );
  NOR4_X1 U23928 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_21__SCAN_IN), .A3(P1_EAX_REG_28__SCAN_IN), .A4(
        P1_REIP_REG_8__SCAN_IN), .ZN(n21033) );
  NAND4_X1 U23929 ( .A1(n21036), .A2(n21035), .A3(n21034), .A4(n21033), .ZN(
        n21042) );
  NOR4_X1 U23930 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .A3(P3_EBX_REG_17__SCAN_IN), .A4(
        P3_EBX_REG_1__SCAN_IN), .ZN(n21040) );
  NOR4_X1 U23931 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(
        P3_INSTQUEUE_REG_6__0__SCAN_IN), .A3(P3_INSTQUEUE_REG_11__6__SCAN_IN), 
        .A4(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n21039) );
  NOR4_X1 U23932 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_2__0__SCAN_IN), .A3(P2_INSTQUEUE_REG_12__5__SCAN_IN), 
        .A4(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n21038) );
  NOR4_X1 U23933 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_EBX_REG_19__SCAN_IN), .A3(P2_DATAO_REG_25__SCAN_IN), .A4(
        P2_DATAO_REG_29__SCAN_IN), .ZN(n21037) );
  NAND4_X1 U23934 ( .A1(n21040), .A2(n21039), .A3(n21038), .A4(n21037), .ZN(
        n21041) );
  NOR4_X1 U23935 ( .A1(n21044), .A2(n21043), .A3(n21042), .A4(n21041), .ZN(
        n21045) );
  NAND4_X1 U23936 ( .A1(n21048), .A2(n21047), .A3(n21046), .A4(n21045), .ZN(
        n21049) );
  XNOR2_X1 U23937 ( .A(n21050), .B(n21049), .ZN(P1_U3088) );
  AND2_X2 U11580 ( .A1(n13460), .A2(n10926), .ZN(n11261) );
  AND2_X1 U11578 ( .A1(n10927), .A2(n13468), .ZN(n11090) );
  AND2_X1 U11626 ( .A1(n10028), .A2(n10027), .ZN(n11182) );
  NOR2_X1 U11627 ( .A1(n14478), .A2(n20956), .ZN(n14490) );
  INV_X2 U11290 ( .A(n14160), .ZN(n14545) );
  CLKBUF_X1 U11162 ( .A(n11297), .Z(n11642) );
  CLKBUF_X2 U11198 ( .A(n10630), .Z(n12707) );
  CLKBUF_X1 U11229 ( .A(n10908), .Z(n9751) );
  CLKBUF_X1 U11239 ( .A(n10735), .Z(n19223) );
  CLKBUF_X1 U11245 ( .A(n15032), .Z(n15053) );
  AND2_X2 U11258 ( .A1(n15108), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9739) );
  CLKBUF_X1 U11685 ( .A(n15137), .Z(n15138) );
  CLKBUF_X1 U12394 ( .A(n16423), .Z(n16424) );
  AND2_X1 U14312 ( .A1(n11911), .A2(n11921), .ZN(n21051) );
  CLKBUF_X1 U14345 ( .A(n11261), .Z(n11262) );
endmodule

