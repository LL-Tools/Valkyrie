

module b14_C_gen_AntiSAT_k_256_5 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, 
        keyinput_f67, keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, 
        keyinput_f72, keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, 
        keyinput_f77, keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, 
        keyinput_f82, keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, 
        keyinput_f87, keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, 
        keyinput_f92, keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, 
        keyinput_f97, keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101, 
        keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105, 
        keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109, 
        keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113, 
        keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117, 
        keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121, 
        keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125, 
        keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67, 
        keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72, 
        keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77, 
        keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82, 
        keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87, 
        keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92, 
        keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97, 
        keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101, 
        keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105, 
        keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109, 
        keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113, 
        keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117, 
        keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121, 
        keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125, 
        keyinput_g126, keyinput_g127, U3352, U3351, U3350, U3349, U3348, U3347, 
        U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, 
        U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, 
        U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, 
        U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, 
        U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, 
        U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, 
        U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, 
        U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, 
        U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, 
        U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, 
        U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, 
        U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, 
        U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, 
        U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, 
        U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, 
        U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, 
        U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, 
        U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, 
        U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, 
        U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, 
        U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, 
        U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, 
        U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, 
        U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_f64, keyinput_f65, keyinput_f66, keyinput_f67,
         keyinput_f68, keyinput_f69, keyinput_f70, keyinput_f71, keyinput_f72,
         keyinput_f73, keyinput_f74, keyinput_f75, keyinput_f76, keyinput_f77,
         keyinput_f78, keyinput_f79, keyinput_f80, keyinput_f81, keyinput_f82,
         keyinput_f83, keyinput_f84, keyinput_f85, keyinput_f86, keyinput_f87,
         keyinput_f88, keyinput_f89, keyinput_f90, keyinput_f91, keyinput_f92,
         keyinput_f93, keyinput_f94, keyinput_f95, keyinput_f96, keyinput_f97,
         keyinput_f98, keyinput_f99, keyinput_f100, keyinput_f101,
         keyinput_f102, keyinput_f103, keyinput_f104, keyinput_f105,
         keyinput_f106, keyinput_f107, keyinput_f108, keyinput_f109,
         keyinput_f110, keyinput_f111, keyinput_f112, keyinput_f113,
         keyinput_f114, keyinput_f115, keyinput_f116, keyinput_f117,
         keyinput_f118, keyinput_f119, keyinput_f120, keyinput_f121,
         keyinput_f122, keyinput_f123, keyinput_f124, keyinput_f125,
         keyinput_f126, keyinput_f127, keyinput_g0, keyinput_g1, keyinput_g2,
         keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7,
         keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12,
         keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17,
         keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22,
         keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27,
         keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32,
         keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37,
         keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42,
         keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47,
         keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52,
         keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57,
         keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62,
         keyinput_g63, keyinput_g64, keyinput_g65, keyinput_g66, keyinput_g67,
         keyinput_g68, keyinput_g69, keyinput_g70, keyinput_g71, keyinput_g72,
         keyinput_g73, keyinput_g74, keyinput_g75, keyinput_g76, keyinput_g77,
         keyinput_g78, keyinput_g79, keyinput_g80, keyinput_g81, keyinput_g82,
         keyinput_g83, keyinput_g84, keyinput_g85, keyinput_g86, keyinput_g87,
         keyinput_g88, keyinput_g89, keyinput_g90, keyinput_g91, keyinput_g92,
         keyinput_g93, keyinput_g94, keyinput_g95, keyinput_g96, keyinput_g97,
         keyinput_g98, keyinput_g99, keyinput_g100, keyinput_g101,
         keyinput_g102, keyinput_g103, keyinput_g104, keyinput_g105,
         keyinput_g106, keyinput_g107, keyinput_g108, keyinput_g109,
         keyinput_g110, keyinput_g111, keyinput_g112, keyinput_g113,
         keyinput_g114, keyinput_g115, keyinput_g116, keyinput_g117,
         keyinput_g118, keyinput_g119, keyinput_g120, keyinput_g121,
         keyinput_g122, keyinput_g123, keyinput_g124, keyinput_g125,
         keyinput_g126, keyinput_g127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2235, n2236, n2237, n2238, n2239, n2240, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
         n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505,
         n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
         n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
         n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
         n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
         n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555,
         n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
         n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
         n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
         n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
         n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
         n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
         n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
         n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
         n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
         n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
         n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
         n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
         n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
         n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
         n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
         n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
         n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785,
         n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
         n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805,
         n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
         n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825,
         n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835,
         n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845,
         n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
         n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140;

  AOI211_X1 U2476 ( .C1(n2289), .C2(n4592), .A(n4086), .B(n3331), .ZN(n3350)
         );
  INV_X1 U2477 ( .A(n3766), .ZN(n3152) );
  BUF_X2 U2478 ( .A(n2939), .Z(n3763) );
  CLKBUF_X2 U2479 ( .A(n2479), .Z(n3915) );
  NOR2_X2 U2480 ( .A1(n4738), .A2(n2252), .ZN(n2958) );
  CLKBUF_X1 U2481 ( .A(n2753), .Z(n2242) );
  INV_X2 U2482 ( .A(n4713), .ZN(n4209) );
  AND4_X1 U2483 ( .A1(n2743), .A2(n5042), .A3(n5040), .A4(n2741), .ZN(n2258)
         );
  INV_X1 U2485 ( .A(n3374), .ZN(n3421) );
  INV_X1 U2486 ( .A(n2252), .ZN(n3069) );
  CLKBUF_X3 U2487 ( .A(n2493), .Z(n2240) );
  INV_X1 U2488 ( .A(n2939), .ZN(n3143) );
  AND3_X4 U2489 ( .A1(n2375), .A2(n2290), .A3(n2432), .ZN(n2535) );
  NAND2_X1 U2490 ( .A1(n4558), .A2(n3232), .ZN(n2487) );
  NAND2_X2 U2491 ( .A1(n3081), .A2(n3080), .ZN(n3842) );
  OAI211_X2 U2492 ( .C1(n3900), .C2(n4578), .A(n4580), .B(n3901), .ZN(n3081)
         );
  XNOR2_X2 U2493 ( .A(n3193), .B(n3955), .ZN(n4136) );
  AOI21_X2 U2494 ( .B1(n3192), .B2(n3953), .A(n3191), .ZN(n3193) );
  NAND2_X2 U2495 ( .A1(n3791), .A2(IR_REG_31__SCAN_IN), .ZN(n2284) );
  BUF_X4 U2496 ( .A(n3069), .Z(n2244) );
  INV_X1 U2497 ( .A(n3763), .ZN(n2235) );
  INV_X2 U2498 ( .A(n3763), .ZN(n2236) );
  OAI21_X1 U2499 ( .B1(n4301), .B2(n4283), .A(n2279), .ZN(n2278) );
  NAND2_X1 U2500 ( .A1(n4325), .A2(n2280), .ZN(n4301) );
  NAND2_X1 U2501 ( .A1(n3682), .A2(n2271), .ZN(n3740) );
  NAND2_X1 U2502 ( .A1(n4002), .A2(n4004), .ZN(n3433) );
  NAND2_X2 U2503 ( .A1(n2476), .A2(n2935), .ZN(n3995) );
  CLKBUF_X1 U2504 ( .A(n2477), .Z(n3912) );
  OAI21_X2 U2505 ( .B1(n2668), .B2(IR_REG_18__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2746) );
  INV_X2 U2506 ( .A(IR_REG_19__SCAN_IN), .ZN(n2741) );
  OR2_X1 U2507 ( .A1(n3822), .A2(n3823), .ZN(n2418) );
  CLKBUF_X1 U2508 ( .A(n3796), .Z(n3872) );
  NAND2_X1 U2509 ( .A1(n2286), .A2(n2703), .ZN(n4183) );
  NAND2_X1 U2510 ( .A1(n4245), .A2(n2269), .ZN(n4221) );
  NAND2_X1 U2511 ( .A1(n4246), .A2(n4252), .ZN(n4245) );
  OR2_X1 U2512 ( .A1(n4491), .A2(n4495), .ZN(n4384) );
  NOR2_X2 U2513 ( .A1(n4174), .A2(n3892), .ZN(n4175) );
  NAND2_X1 U2514 ( .A1(n3611), .A2(n3968), .ZN(n3613) );
  OR2_X2 U2515 ( .A1(n3493), .A2(n3966), .ZN(n3492) );
  AND2_X1 U2516 ( .A1(n4140), .A2(n3784), .ZN(n3191) );
  NAND2_X1 U2517 ( .A1(n2528), .A2(n2527), .ZN(n3465) );
  NAND2_X1 U2518 ( .A1(n2282), .A2(n3433), .ZN(n3436) );
  OR2_X2 U2519 ( .A1(n3740), .A2(n4468), .ZN(n4366) );
  NAND2_X1 U2520 ( .A1(n3379), .A2(n2495), .ZN(n3370) );
  NAND2_X1 U2521 ( .A1(n3380), .A2(n3957), .ZN(n3379) );
  NAND2_X1 U2522 ( .A1(n2765), .A2(n3355), .ZN(n3354) );
  NAND3_X2 U2523 ( .A1(n2511), .A2(n2510), .A3(n2509), .ZN(n4084) );
  NAND4_X1 U2524 ( .A1(n2534), .A2(n2533), .A3(n2532), .A4(n2531), .ZN(n4082)
         );
  INV_X1 U2525 ( .A(n2934), .ZN(n2476) );
  NAND4_X2 U2526 ( .A1(n2499), .A2(n2498), .A3(n2497), .A4(n2496), .ZN(n4085)
         );
  NAND4_X2 U2527 ( .A1(n2471), .A2(n2470), .A3(n2469), .A4(n2468), .ZN(n2934)
         );
  CLKBUF_X3 U2528 ( .A(n3912), .Z(n2735) );
  INV_X2 U2529 ( .A(n2461), .ZN(n2758) );
  CLKBUF_X3 U2530 ( .A(n2478), .Z(n2715) );
  NAND2_X1 U2531 ( .A1(n2809), .A2(n4559), .ZN(n3215) );
  NAND2_X1 U2532 ( .A1(n2319), .A2(IR_REG_31__SCAN_IN), .ZN(n2460) );
  XNOR2_X1 U2533 ( .A(n2751), .B(IR_REG_22__SCAN_IN), .ZN(n4561) );
  NAND2_X1 U2534 ( .A1(n2293), .A2(IR_REG_31__SCAN_IN), .ZN(n2866) );
  NOR2_X1 U2535 ( .A1(n2427), .A2(n2287), .ZN(n2425) );
  NOR2_X1 U2536 ( .A1(n2449), .A2(IR_REG_12__SCAN_IN), .ZN(n2295) );
  AND2_X1 U2537 ( .A1(n2491), .A2(n2377), .ZN(n2375) );
  INV_X1 U2538 ( .A(IR_REG_16__SCAN_IN), .ZN(n5042) );
  INV_X1 U2539 ( .A(IR_REG_24__SCAN_IN), .ZN(n2803) );
  INV_X1 U2540 ( .A(IR_REG_6__SCAN_IN), .ZN(n2545) );
  NOR2_X1 U2541 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2447)
         );
  NOR2_X1 U2542 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2446)
         );
  NOR2_X1 U2543 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2448)
         );
  INV_X2 U2544 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U2545 ( .A(IR_REG_2__SCAN_IN), .ZN(n2491) );
  INV_X1 U2546 ( .A(IR_REG_4__SCAN_IN), .ZN(n2515) );
  NAND2_X1 U2547 ( .A1(n3636), .A2(n2619), .ZN(n2237) );
  NAND2_X1 U2548 ( .A1(n3636), .A2(n2619), .ZN(n3731) );
  OR2_X4 U2549 ( .A1(n3181), .A2(n2921), .ZN(n2939) );
  OAI21_X2 U2550 ( .B1(n4149), .B2(n2731), .A(n2730), .ZN(n3192) );
  NOR2_X1 U2551 ( .A1(n4558), .A2(n3232), .ZN(n2478) );
  NAND2_X1 U2552 ( .A1(n4558), .A2(n2285), .ZN(n2479) );
  OAI21_X1 U2553 ( .B1(n2395), .B2(n2393), .A(n2391), .ZN(n3851) );
  XNOR2_X1 U2554 ( .A(n2746), .B(IR_REG_19__SCAN_IN), .ZN(n4563) );
  NOR2_X2 U2555 ( .A1(n4327), .A2(n3806), .ZN(n2294) );
  NAND2_X1 U2556 ( .A1(n2278), .A2(n3981), .ZN(n4263) );
  NAND2_X2 U2557 ( .A1(n2397), .A2(n2396), .ZN(n3625) );
  NOR2_X1 U2558 ( .A1(n4558), .A2(n3232), .ZN(n2238) );
  AOI21_X4 U2559 ( .B1(n3832), .B2(n2259), .A(n2373), .ZN(n3514) );
  AND2_X2 U2560 ( .A1(n3852), .A2(n3135), .ZN(n3822) );
  NAND2_X1 U2561 ( .A1(n2742), .A2(IR_REG_31__SCAN_IN), .ZN(n2744) );
  INV_X1 U2562 ( .A(n2487), .ZN(n2239) );
  NOR2_X2 U2563 ( .A1(n3582), .A2(n3555), .ZN(n2254) );
  NOR2_X2 U2564 ( .A1(n3078), .A2(n3077), .ZN(n3900) );
  AOI21_X2 U2565 ( .B1(n3064), .B2(n2276), .A(n3063), .ZN(n3078) );
  XNOR2_X1 U2566 ( .A(n2744), .B(n2743), .ZN(n2753) );
  INV_X4 U2567 ( .A(IR_REG_0__SCAN_IN), .ZN(n2289) );
  INV_X2 U2568 ( .A(n3367), .ZN(n3307) );
  NAND2_X2 U2569 ( .A1(n3613), .A2(n2592), .ZN(n3636) );
  NAND2_X2 U2570 ( .A1(n2753), .A2(n2757), .ZN(n2921) );
  MUX2_X2 U2571 ( .A(n3211), .B(n3210), .S(n4759), .Z(n3213) );
  MUX2_X2 U2572 ( .A(n3204), .B(n3210), .S(n4770), .Z(n3209) );
  NOR2_X4 U2573 ( .A1(n2567), .A2(n2450), .ZN(n2749) );
  NAND2_X2 U2574 ( .A1(n2535), .A2(n2440), .ZN(n2567) );
  OAI21_X2 U2575 ( .B1(n3625), .B2(n3626), .A(n3627), .ZN(n3704) );
  OR2_X1 U2576 ( .A1(n2949), .A2(n3301), .ZN(n3996) );
  NAND3_X2 U2577 ( .A1(n2433), .A2(n2490), .A3(n2288), .ZN(n2949) );
  NAND2_X2 U2578 ( .A1(n3995), .A2(n3993), .ZN(n2765) );
  BUF_X1 U2579 ( .A(n4386), .Z(n2243) );
  NAND2_X2 U2580 ( .A1(n3834), .A2(n3833), .ZN(n3832) );
  AOI21_X2 U2581 ( .B1(n4344), .B2(n2661), .A(n2660), .ZN(n4324) );
  AOI21_X2 U2582 ( .B1(n4263), .B2(n2686), .A(n2277), .ZN(n4246) );
  AOI21_X2 U2583 ( .B1(n4221), .B2(n2696), .A(n2695), .ZN(n4199) );
  AOI21_X2 U2584 ( .B1(n3492), .B2(n2571), .A(n2430), .ZN(n3690) );
  NAND2_X1 U2585 ( .A1(n4363), .A2(n4373), .ZN(n4362) );
  AOI21_X2 U2586 ( .B1(n3654), .B2(n2635), .A(n2270), .ZN(n4363) );
  XNOR2_X2 U2587 ( .A(n2460), .B(IR_REG_29__SCAN_IN), .ZN(n3232) );
  AND2_X1 U2588 ( .A1(n2439), .A2(n2545), .ZN(n2440) );
  NOR2_X1 U2589 ( .A1(IR_REG_8__SCAN_IN), .A2(IR_REG_7__SCAN_IN), .ZN(n2439)
         );
  NAND2_X1 U2590 ( .A1(n2262), .A2(n2793), .ZN(n2333) );
  AND2_X2 U2591 ( .A1(n5057), .A2(n2289), .ZN(n2290) );
  INV_X1 U2592 ( .A(n3770), .ZN(n2410) );
  OAI22_X1 U2593 ( .A1(n3307), .A2(n2939), .B1(n3215), .B2(n2289), .ZN(n2922)
         );
  INV_X1 U2594 ( .A(n3215), .ZN(n3181) );
  INV_X1 U2595 ( .A(n2345), .ZN(n2340) );
  AOI21_X1 U2596 ( .B1(REG1_REG_5__SCAN_IN), .B2(n3218), .A(n3234), .ZN(n2881)
         );
  AOI21_X1 U2597 ( .B1(n3252), .B2(n3248), .A(n3247), .ZN(n2884) );
  OR2_X1 U2598 ( .A1(n4660), .A2(n2857), .ZN(n2859) );
  OR2_X1 U2599 ( .A1(n4189), .A2(n3951), .ZN(n4167) );
  AND2_X1 U2600 ( .A1(n3980), .A2(n4284), .ZN(n2279) );
  NAND2_X1 U2601 ( .A1(n2318), .A2(n2749), .ZN(n2319) );
  AND2_X1 U2602 ( .A1(n2425), .A2(n2265), .ZN(n2318) );
  NOR2_X1 U2603 ( .A1(n2867), .A2(n2868), .ZN(n4113) );
  NOR2_X1 U2604 ( .A1(n4028), .A2(n2317), .ZN(n2316) );
  INV_X1 U2605 ( .A(n4022), .ZN(n2314) );
  INV_X1 U2606 ( .A(IR_REG_13__SCAN_IN), .ZN(n2442) );
  AND2_X1 U2607 ( .A1(n3924), .A2(n2309), .ZN(n2308) );
  NAND2_X1 U2608 ( .A1(n4225), .A2(n2310), .ZN(n2309) );
  INV_X1 U2609 ( .A(n4034), .ZN(n2310) );
  NAND2_X1 U2610 ( .A1(n2308), .A2(n2311), .ZN(n2307) );
  INV_X1 U2611 ( .A(n4225), .ZN(n2311) );
  OR2_X1 U2612 ( .A1(n2622), .A2(n2621), .ZN(n3728) );
  NAND2_X1 U2613 ( .A1(n2768), .A2(n4004), .ZN(n2324) );
  NOR2_X1 U2614 ( .A1(n4005), .A2(n2325), .ZN(n2321) );
  AOI21_X1 U2615 ( .B1(n2333), .B2(n2331), .A(n3935), .ZN(n2330) );
  NOR2_X1 U2616 ( .A1(n2334), .A2(n3933), .ZN(n2331) );
  NOR2_X1 U2617 ( .A1(n2808), .A2(n2826), .ZN(n2821) );
  INV_X1 U2618 ( .A(n2806), .ZN(n2808) );
  NAND2_X1 U2619 ( .A1(n2451), .A2(n2426), .ZN(n2287) );
  INV_X1 U2620 ( .A(IR_REG_26__SCAN_IN), .ZN(n2426) );
  NAND2_X1 U2621 ( .A1(n2428), .A2(n2453), .ZN(n2427) );
  INV_X1 U2622 ( .A(IR_REG_25__SCAN_IN), .ZN(n2453) );
  INV_X1 U2623 ( .A(n2452), .ZN(n2428) );
  INV_X1 U2624 ( .A(IR_REG_23__SCAN_IN), .ZN(n2810) );
  AOI21_X1 U2625 ( .B1(n2421), .B2(n2268), .A(n2420), .ZN(n2419) );
  INV_X1 U2626 ( .A(n3889), .ZN(n2420) );
  NOR2_X1 U2627 ( .A1(n2424), .A2(n2422), .ZN(n2421) );
  INV_X1 U2628 ( .A(n3824), .ZN(n2422) );
  NOR2_X1 U2629 ( .A1(n2724), .A2(n3174), .ZN(n2732) );
  AOI21_X1 U2630 ( .B1(n2413), .B2(n2423), .A(n2246), .ZN(n2412) );
  XOR2_X1 U2631 ( .A(n3769), .B(n3768), .Z(n3770) );
  INV_X1 U2632 ( .A(n3029), .ZN(n2400) );
  INV_X1 U2633 ( .A(n2402), .ZN(n2401) );
  OAI21_X1 U2634 ( .B1(n3023), .B2(n2403), .A(n3590), .ZN(n2402) );
  INV_X1 U2635 ( .A(n2399), .ZN(n2398) );
  OAI21_X1 U2636 ( .B1(n3023), .B2(n2400), .A(n3589), .ZN(n2399) );
  INV_X1 U2637 ( .A(n3124), .ZN(n2393) );
  AOI21_X1 U2638 ( .B1(n2392), .B2(n3124), .A(n2261), .ZN(n2391) );
  XNOR2_X1 U2639 ( .A(n3046), .B(n3152), .ZN(n3705) );
  XNOR2_X1 U2640 ( .A(n2947), .B(n3152), .ZN(n2953) );
  NOR2_X1 U2641 ( .A1(n2611), .A2(n4861), .ZN(n2625) );
  NOR2_X1 U2642 ( .A1(n3222), .A2(n2825), .ZN(n2809) );
  NOR2_X1 U2643 ( .A1(n2835), .A2(n2363), .ZN(n4092) );
  NAND2_X1 U2644 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n2363) );
  INV_X1 U2645 ( .A(n2290), .ZN(n2473) );
  NAND2_X1 U2646 ( .A1(n2346), .A2(n4566), .ZN(n2345) );
  NOR2_X1 U2647 ( .A1(n3237), .A2(n2342), .ZN(n2842) );
  NOR2_X1 U2648 ( .A1(n2344), .A2(n2343), .ZN(n2342) );
  XNOR2_X1 U2649 ( .A(n2881), .B(n2372), .ZN(n3263) );
  NOR2_X1 U2650 ( .A1(n3263), .A2(n3262), .ZN(n3261) );
  OAI22_X1 U2651 ( .A1(n3268), .A2(n2887), .B1(n2886), .B2(n2885), .ZN(n4598)
         );
  NAND2_X1 U2652 ( .A1(n4598), .A2(n4599), .ZN(n4597) );
  XNOR2_X1 U2653 ( .A(n2848), .B(n2847), .ZN(n4610) );
  XNOR2_X1 U2654 ( .A(n2891), .B(n2851), .ZN(n4631) );
  NAND2_X1 U2655 ( .A1(n4631), .A2(REG1_REG_12__SCAN_IN), .ZN(n4630) );
  OR2_X1 U2656 ( .A1(n4653), .A2(n3743), .ZN(n2358) );
  NAND2_X1 U2657 ( .A1(n4669), .A2(n2860), .ZN(n4678) );
  OR2_X1 U2658 ( .A1(n4673), .A2(REG1_REG_16__SCAN_IN), .ZN(n2370) );
  NAND2_X1 U2659 ( .A1(n4678), .A2(n4680), .ZN(n4679) );
  AND2_X1 U2660 ( .A1(n2792), .A2(n2793), .ZN(n4150) );
  NOR2_X1 U2661 ( .A1(n4439), .A2(n4429), .ZN(n2277) );
  NAND2_X1 U2662 ( .A1(n2281), .A2(n4328), .ZN(n2280) );
  INV_X1 U2663 ( .A(n4455), .ZN(n2281) );
  OR2_X1 U2664 ( .A1(n4467), .A2(n3741), .ZN(n3917) );
  NOR2_X1 U2665 ( .A1(n2560), .A2(n2559), .ZN(n2572) );
  OR2_X1 U2666 ( .A1(n2263), .A2(n2435), .ZN(n2430) );
  INV_X1 U2667 ( .A(n2302), .ZN(n2301) );
  OAI21_X1 U2668 ( .B1(n4012), .B2(n2303), .A(n4011), .ZN(n2302) );
  INV_X1 U2669 ( .A(n3437), .ZN(n2327) );
  INV_X1 U2670 ( .A(n4375), .ZN(n4312) );
  AND2_X1 U2671 ( .A1(n4570), .A2(n2863), .ZN(n4478) );
  OR2_X1 U2672 ( .A1(n4570), .A2(n3162), .ZN(n4481) );
  NAND2_X1 U2673 ( .A1(n3359), .A2(n3307), .ZN(n3390) );
  OR2_X1 U2674 ( .A1(n3309), .A2(n4561), .ZN(n4733) );
  AND2_X1 U2675 ( .A1(n3215), .A2(n4716), .ZN(n3279) );
  NAND2_X1 U2676 ( .A1(n2810), .A2(n2803), .ZN(n2452) );
  AND2_X1 U2677 ( .A1(n2447), .A2(n2448), .ZN(n2298) );
  INV_X1 U2678 ( .A(n2500), .ZN(n2376) );
  OR2_X1 U2679 ( .A1(n3182), .A2(n3175), .ZN(n3875) );
  AOI21_X1 U2680 ( .B1(n2380), .B2(n2382), .A(n2274), .ZN(n2378) );
  OR2_X1 U2681 ( .A1(n3182), .A2(n3173), .ZN(n4571) );
  AOI21_X1 U2682 ( .B1(n4479), .B2(n3764), .A(n3068), .ZN(n4578) );
  NAND2_X1 U2683 ( .A1(n2721), .A2(n2720), .ZN(n4393) );
  OR2_X1 U2684 ( .A1(n2487), .A2(n3317), .ZN(n2481) );
  XNOR2_X1 U2685 ( .A(n2492), .B(n2491), .ZN(n3333) );
  NAND2_X1 U2686 ( .A1(n2473), .A2(IR_REG_31__SCAN_IN), .ZN(n2492) );
  OR2_X1 U2687 ( .A1(n4673), .A2(n2369), .ZN(n2367) );
  OR2_X1 U2688 ( .A1(n4685), .A2(REG1_REG_16__SCAN_IN), .ZN(n2369) );
  OR2_X1 U2689 ( .A1(n2251), .A2(n4685), .ZN(n2368) );
  OR2_X1 U2690 ( .A1(n4113), .A2(n4112), .ZN(n4115) );
  INV_X1 U2691 ( .A(n4640), .ZN(n4677) );
  INV_X1 U2692 ( .A(n2328), .ZN(n3196) );
  AOI21_X1 U2693 ( .B1(n4167), .B2(n2334), .A(n2329), .ZN(n2328) );
  INV_X1 U2694 ( .A(n4563), .ZN(n4123) );
  OR2_X1 U2695 ( .A1(n3786), .A2(n4556), .ZN(n2830) );
  AND2_X1 U2696 ( .A1(n3873), .A2(n2249), .ZN(n2394) );
  NAND2_X1 U2697 ( .A1(n2297), .A2(n2296), .ZN(n2449) );
  INV_X1 U2698 ( .A(IR_REG_9__SCAN_IN), .ZN(n2297) );
  INV_X1 U2699 ( .A(n2394), .ZN(n2392) );
  AND2_X1 U2700 ( .A1(n3797), .A2(n3798), .ZN(n3124) );
  INV_X1 U2701 ( .A(n3565), .ZN(n3023) );
  NOR2_X1 U2702 ( .A1(n3881), .A2(n2389), .ZN(n2388) );
  NAND2_X1 U2703 ( .A1(n3339), .A2(n2362), .ZN(n2839) );
  OR2_X1 U2704 ( .A1(n3333), .A2(n2837), .ZN(n2362) );
  OR2_X1 U2705 ( .A1(n4342), .A2(n4222), .ZN(n4303) );
  INV_X1 U2706 ( .A(n2316), .ZN(n2315) );
  AND2_X1 U2707 ( .A1(n4033), .A2(n2313), .ZN(n2312) );
  NAND2_X1 U2708 ( .A1(n2316), .A2(n2314), .ZN(n2313) );
  OR2_X1 U2709 ( .A1(n3733), .A2(n3728), .ZN(n3730) );
  AND2_X1 U2710 ( .A1(n3727), .A2(n3949), .ZN(n2619) );
  OR2_X1 U2711 ( .A1(n4206), .A2(n4190), .ZN(n4174) );
  OR2_X1 U2712 ( .A1(n2617), .A2(IR_REG_14__SCAN_IN), .ZN(n2632) );
  CLKBUF_X1 U2713 ( .A(n2616), .Z(n2617) );
  AND2_X1 U2714 ( .A1(n2386), .A2(n2384), .ZN(n2383) );
  INV_X1 U2715 ( .A(n3883), .ZN(n2384) );
  INV_X1 U2716 ( .A(n2419), .ZN(n2415) );
  XNOR2_X1 U2717 ( .A(n2967), .B(n3152), .ZN(n2971) );
  NAND2_X1 U2718 ( .A1(n2966), .A2(n2965), .ZN(n2967) );
  INV_X1 U2719 ( .A(n3099), .ZN(n2390) );
  AOI21_X1 U2720 ( .B1(n2383), .B2(n2381), .A(n3805), .ZN(n2380) );
  INV_X1 U2721 ( .A(n2388), .ZN(n2381) );
  INV_X1 U2722 ( .A(n2383), .ZN(n2382) );
  AND2_X1 U2723 ( .A1(n3112), .A2(n3111), .ZN(n3864) );
  AND2_X1 U2724 ( .A1(n3040), .A2(n3041), .ZN(n3626) );
  NAND2_X1 U2725 ( .A1(n3024), .A2(n3023), .ZN(n3563) );
  NAND2_X1 U2726 ( .A1(n2387), .A2(n3844), .ZN(n2386) );
  INV_X1 U2727 ( .A(n3881), .ZN(n2387) );
  NAND2_X1 U2728 ( .A1(n3842), .A2(n2388), .ZN(n2385) );
  NAND2_X1 U2729 ( .A1(n2519), .A2(REG3_REG_5__SCAN_IN), .ZN(n2529) );
  NOR2_X1 U2730 ( .A1(n2529), .A2(n3259), .ZN(n2538) );
  OR4_X1 U2731 ( .A1(n3932), .A2(n3935), .A3(n3934), .A4(n3936), .ZN(n3943) );
  OAI21_X1 U2732 ( .B1(n3333), .B2(REG2_REG_2__SCAN_IN), .A(n2836), .ZN(n3337)
         );
  NAND2_X1 U2733 ( .A1(n2365), .A2(n2876), .ZN(n2877) );
  NOR2_X1 U2734 ( .A1(n3245), .A2(n2351), .ZN(n2349) );
  NOR2_X1 U2735 ( .A1(n3245), .A2(n2372), .ZN(n2348) );
  AND2_X1 U2736 ( .A1(n2353), .A2(n2352), .ZN(n2844) );
  NAND2_X1 U2737 ( .A1(n2883), .A2(REG2_REG_7__SCAN_IN), .ZN(n2352) );
  XNOR2_X1 U2738 ( .A(n2844), .B(n2886), .ZN(n3269) );
  NAND2_X1 U2739 ( .A1(n4597), .A2(n2888), .ZN(n2889) );
  NAND2_X1 U2740 ( .A1(n4600), .A2(n2846), .ZN(n2848) );
  NAND2_X1 U2741 ( .A1(n4610), .A2(REG2_REG_10__SCAN_IN), .ZN(n4609) );
  NAND2_X1 U2742 ( .A1(n4621), .A2(n2850), .ZN(n2852) );
  NAND2_X1 U2743 ( .A1(n4646), .A2(n2893), .ZN(n2895) );
  AND3_X1 U2744 ( .A1(n2368), .A2(n2275), .A3(n2367), .ZN(n2903) );
  AND2_X1 U2745 ( .A1(n2793), .A2(n4053), .ZN(n2334) );
  INV_X1 U2746 ( .A(n2333), .ZN(n2329) );
  INV_X1 U2747 ( .A(n4393), .ZN(n4157) );
  OR2_X1 U2748 ( .A1(n2725), .A2(n2732), .ZN(n4156) );
  AND2_X1 U2749 ( .A1(n2724), .A2(n2714), .ZN(n4178) );
  AND2_X1 U2750 ( .A1(n2307), .A2(n2786), .ZN(n2306) );
  NAND2_X1 U2751 ( .A1(n2691), .A2(REG3_REG_23__SCAN_IN), .ZN(n2697) );
  NOR2_X1 U2752 ( .A1(n2677), .A2(n2676), .ZN(n2687) );
  OR2_X1 U2753 ( .A1(n4303), .A2(n4223), .ZN(n4280) );
  NAND2_X1 U2754 ( .A1(n2662), .A2(REG3_REG_19__SCAN_IN), .ZN(n2669) );
  NOR2_X1 U2755 ( .A1(n2646), .A2(n2645), .ZN(n2647) );
  NAND2_X1 U2756 ( .A1(n2780), .A2(n4034), .ZN(n4342) );
  NAND2_X1 U2757 ( .A1(n4362), .A2(n2644), .ZN(n4344) );
  NAND2_X1 U2758 ( .A1(n4469), .A2(n4377), .ZN(n2644) );
  NAND2_X1 U2759 ( .A1(n2625), .A2(REG3_REG_15__SCAN_IN), .ZN(n2636) );
  NAND2_X1 U2760 ( .A1(n3734), .A2(n3733), .ZN(n3735) );
  OR2_X1 U2761 ( .A1(n2593), .A2(n3630), .ZN(n2603) );
  OR2_X1 U2762 ( .A1(n2603), .A2(n2602), .ZN(n2611) );
  NAND2_X1 U2763 ( .A1(n3610), .A2(n4026), .ZN(n3645) );
  NAND2_X1 U2764 ( .A1(n2771), .A2(n4022), .ZN(n3610) );
  NAND2_X1 U2765 ( .A1(n2538), .A2(REG3_REG_7__SCAN_IN), .ZN(n2548) );
  NAND2_X1 U2766 ( .A1(n2769), .A2(n4012), .ZN(n3573) );
  AND2_X1 U2767 ( .A1(n4006), .A2(n4012), .ZN(n3966) );
  INV_X1 U2768 ( .A(n2992), .ZN(n3516) );
  NAND2_X1 U2769 ( .A1(n2322), .A2(n2320), .ZN(n3463) );
  INV_X1 U2770 ( .A(n2323), .ZN(n2322) );
  OAI21_X1 U2771 ( .B1(n2324), .B2(n4005), .A(n4020), .ZN(n2323) );
  AND2_X1 U2772 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2519) );
  OAI21_X1 U2773 ( .B1(n2765), .B2(n3356), .A(n3995), .ZN(n3382) );
  NAND2_X1 U2774 ( .A1(n2493), .A2(DATAI_0_), .ZN(n2291) );
  NOR3_X1 U2775 ( .A1(n3206), .A2(n4389), .A3(n3205), .ZN(n4386) );
  OAI21_X1 U2776 ( .B1(n4167), .B2(n2332), .A(n2330), .ZN(n2337) );
  NAND2_X1 U2777 ( .A1(n2333), .A2(n3194), .ZN(n2332) );
  NAND2_X1 U2778 ( .A1(n4152), .A2(n3771), .ZN(n3206) );
  AND2_X2 U2779 ( .A1(n4175), .A2(n4154), .ZN(n4152) );
  AND2_X1 U2780 ( .A1(n2740), .A2(n2739), .ZN(n4396) );
  OR2_X1 U2781 ( .A1(n3780), .A2(n2758), .ZN(n2740) );
  INV_X1 U2782 ( .A(n3827), .ZN(n4190) );
  NAND2_X1 U2783 ( .A1(n4238), .A2(n4207), .ZN(n4206) );
  AND2_X1 U2784 ( .A1(n2245), .A2(n4236), .ZN(n4238) );
  AND2_X1 U2785 ( .A1(n4265), .A2(n4256), .ZN(n2245) );
  NOR2_X1 U2786 ( .A1(n4287), .A2(n4429), .ZN(n4265) );
  NAND2_X1 U2787 ( .A1(n2294), .A2(n4292), .ZN(n4287) );
  NAND2_X1 U2788 ( .A1(n4348), .A2(n4328), .ZN(n4327) );
  AND2_X1 U2789 ( .A1(n4367), .A2(n4357), .ZN(n4348) );
  NOR2_X2 U2790 ( .A1(n4366), .A2(n4377), .ZN(n4367) );
  INV_X1 U2791 ( .A(n3708), .ZN(n3681) );
  AND2_X1 U2792 ( .A1(n3682), .A2(n3681), .ZN(n3742) );
  OR2_X1 U2793 ( .A1(n3688), .A2(n3592), .ZN(n3637) );
  MUX2_X1 U2794 ( .A(n4629), .B(DATAI_12_), .S(n2240), .Z(n3715) );
  INV_X1 U2795 ( .A(n3692), .ZN(n3689) );
  NAND2_X1 U2796 ( .A1(n2254), .A2(n3689), .ZN(n3688) );
  OR2_X1 U2797 ( .A1(n3306), .A2(n2242), .ZN(n4309) );
  INV_X1 U2798 ( .A(n4309), .ZN(n4477) );
  OAI21_X1 U2799 ( .B1(n3227), .B2(D_REG_0__SCAN_IN), .A(n3229), .ZN(n3311) );
  INV_X1 U2800 ( .A(n2821), .ZN(n3227) );
  INV_X1 U2801 ( .A(IR_REG_7__SCAN_IN), .ZN(n2554) );
  INV_X1 U2802 ( .A(IR_REG_5__SCAN_IN), .ZN(n2377) );
  NAND2_X1 U2803 ( .A1(n2361), .A2(n2360), .ZN(n2474) );
  NAND2_X1 U2804 ( .A1(n5057), .A2(IR_REG_31__SCAN_IN), .ZN(n2360) );
  NAND2_X1 U2805 ( .A1(n2472), .A2(IR_REG_1__SCAN_IN), .ZN(n2361) );
  NOR2_X1 U2806 ( .A1(n3453), .A2(n3452), .ZN(n2373) );
  NAND2_X1 U2807 ( .A1(n3453), .A2(n3452), .ZN(n2374) );
  NAND2_X1 U2808 ( .A1(n2416), .A2(n2419), .ZN(n3762) );
  AND2_X1 U2809 ( .A1(n2412), .A2(n2410), .ZN(n2409) );
  OAI21_X1 U2810 ( .B1(n2412), .B2(n3770), .A(n2407), .ZN(n2406) );
  NAND2_X1 U2811 ( .A1(n2412), .A2(n2408), .ZN(n2407) );
  NAND2_X1 U2812 ( .A1(n2414), .A2(n2410), .ZN(n2408) );
  NAND2_X1 U2813 ( .A1(n2413), .A2(n3770), .ZN(n2411) );
  AOI22_X1 U2814 ( .A1(n2401), .A2(n2403), .B1(n2398), .B2(n2400), .ZN(n2396)
         );
  INV_X1 U2815 ( .A(n4571), .ZN(n3905) );
  INV_X1 U2816 ( .A(n3852), .ZN(n3853) );
  INV_X1 U2817 ( .A(n3875), .ZN(n4577) );
  NAND2_X1 U2818 ( .A1(n3563), .A2(n3029), .ZN(n3588) );
  CLKBUF_X1 U2819 ( .A(n3297), .Z(n3298) );
  NAND2_X1 U2820 ( .A1(n3832), .A2(n2983), .ZN(n3455) );
  NAND2_X1 U2821 ( .A1(n2418), .A2(n3824), .ZN(n3891) );
  INV_X1 U2822 ( .A(n3861), .ZN(n4581) );
  NAND2_X1 U2823 ( .A1(n2708), .A2(n2707), .ZN(n4211) );
  INV_X1 U2824 ( .A(n4193), .ZN(n4233) );
  AND2_X1 U2825 ( .A1(n2683), .A2(n2682), .ZN(n2684) );
  NAND4_X1 U2826 ( .A1(n2667), .A2(n2666), .A3(n2665), .A4(n2664), .ZN(n4332)
         );
  NAND4_X1 U2827 ( .A1(n2466), .A2(n2465), .A3(n2464), .A4(n2463), .ZN(n4455)
         );
  NAND4_X1 U2828 ( .A1(n2653), .A2(n2652), .A3(n2651), .A4(n2650), .ZN(n4576)
         );
  NAND4_X1 U2829 ( .A1(n2631), .A2(n2630), .A3(n2629), .A4(n2628), .ZN(n4479)
         );
  NAND4_X1 U2830 ( .A1(n2615), .A2(n2614), .A3(n2613), .A4(n2612), .ZN(n4467)
         );
  NAND4_X1 U2831 ( .A1(n2608), .A2(n2607), .A3(n2606), .A4(n2605), .ZN(n4075)
         );
  NAND4_X1 U2832 ( .A1(n2589), .A2(n2588), .A3(n2587), .A4(n2586), .ZN(n4077)
         );
  NAND4_X1 U2833 ( .A1(n2578), .A2(n2577), .A3(n2576), .A4(n2575), .ZN(n4078)
         );
  NAND4_X1 U2834 ( .A1(n2566), .A2(n2565), .A3(n2564), .A4(n2563), .ZN(n4079)
         );
  NAND4_X1 U2835 ( .A1(n2553), .A2(n2552), .A3(n2551), .A4(n2550), .ZN(n4080)
         );
  OR2_X1 U2836 ( .A1(n2479), .A2(n2837), .ZN(n2433) );
  OAI21_X1 U2837 ( .B1(n4092), .B2(n3336), .A(n3337), .ZN(n3339) );
  NAND2_X1 U2838 ( .A1(n4684), .A2(n2364), .ZN(n3341) );
  AND2_X1 U2839 ( .A1(n3345), .A2(n2880), .ZN(n3236) );
  OAI21_X1 U2840 ( .B1(n3344), .B2(n2247), .A(n2338), .ZN(n3237) );
  NAND2_X1 U2841 ( .A1(n2340), .A2(n2339), .ZN(n2338) );
  INV_X1 U2842 ( .A(n3238), .ZN(n2339) );
  INV_X1 U2843 ( .A(n2341), .ZN(n3239) );
  OAI21_X1 U2844 ( .B1(n3344), .B2(n2841), .A(n2345), .ZN(n2341) );
  NOR2_X1 U2845 ( .A1(n3261), .A2(n2371), .ZN(n3252) );
  AND2_X1 U2846 ( .A1(n2882), .A2(n4565), .ZN(n2371) );
  AND2_X1 U2847 ( .A1(n2350), .A2(n2354), .ZN(n3246) );
  NAND2_X1 U2848 ( .A1(n3258), .A2(REG2_REG_6__SCAN_IN), .ZN(n2350) );
  NAND2_X1 U2849 ( .A1(n4601), .A2(n4602), .ZN(n4600) );
  XNOR2_X1 U2850 ( .A(n2889), .B(n2847), .ZN(n4615) );
  NAND2_X1 U2851 ( .A1(n4615), .A2(REG1_REG_10__SCAN_IN), .ZN(n4614) );
  NAND2_X1 U2852 ( .A1(n4622), .A2(n4623), .ZN(n4621) );
  XNOR2_X1 U2853 ( .A(n2852), .B(n2851), .ZN(n4633) );
  NAND2_X1 U2854 ( .A1(n4633), .A2(REG2_REG_12__SCAN_IN), .ZN(n4632) );
  AND2_X1 U2855 ( .A1(n4593), .A2(n4066), .ZN(n4640) );
  NAND2_X1 U2856 ( .A1(n4630), .A2(n2892), .ZN(n4647) );
  NAND2_X1 U2857 ( .A1(n4647), .A2(n4648), .ZN(n4646) );
  XNOR2_X1 U2858 ( .A(n2895), .B(n4723), .ZN(n4657) );
  INV_X1 U2859 ( .A(n2358), .ZN(n4652) );
  NAND2_X1 U2860 ( .A1(n2359), .A2(REG2_REG_14__SCAN_IN), .ZN(n2356) );
  NAND2_X1 U2861 ( .A1(n2855), .A2(n2359), .ZN(n2355) );
  INV_X1 U2862 ( .A(n4661), .ZN(n2359) );
  INV_X1 U2863 ( .A(n2855), .ZN(n2357) );
  XNOR2_X1 U2864 ( .A(n2859), .B(n4720), .ZN(n4670) );
  NAND2_X1 U2865 ( .A1(n4679), .A2(n2347), .ZN(n2867) );
  NAND2_X1 U2866 ( .A1(n4718), .A2(n2649), .ZN(n2347) );
  NAND2_X1 U2867 ( .A1(n4167), .A2(n4053), .ZN(n2335) );
  NAND2_X1 U2868 ( .A1(n4209), .A2(n3365), .ZN(n4317) );
  NAND2_X1 U2869 ( .A1(n2300), .A2(n2301), .ZN(n3541) );
  INV_X1 U2870 ( .A(n3497), .ZN(n3472) );
  INV_X1 U2871 ( .A(n4382), .ZN(n4347) );
  NAND2_X1 U2872 ( .A1(n2326), .A2(n4004), .ZN(n3401) );
  NAND2_X1 U2873 ( .A1(n2327), .A2(n4002), .ZN(n2326) );
  OR2_X1 U2874 ( .A1(n3168), .A2(n4733), .ZN(n4369) );
  INV_X2 U2875 ( .A(n4767), .ZN(n4770) );
  XNOR2_X1 U2876 ( .A(n2243), .B(n4128), .ZN(n4495) );
  INV_X2 U2877 ( .A(n4757), .ZN(n4759) );
  INV_X1 U2878 ( .A(n4714), .ZN(n4715) );
  INV_X1 U2879 ( .A(n2293), .ZN(n2457) );
  XNOR2_X1 U2880 ( .A(n2807), .B(IR_REG_26__SCAN_IN), .ZN(n4559) );
  NOR2_X1 U2881 ( .A1(n2801), .A2(n2452), .ZN(n2798) );
  AND2_X1 U2882 ( .A1(n2862), .A2(STATE_REG_SCAN_IN), .ZN(n4716) );
  INV_X1 U2883 ( .A(IR_REG_21__SCAN_IN), .ZN(n2747) );
  INV_X1 U2884 ( .A(n4111), .ZN(n4717) );
  INV_X1 U2885 ( .A(n2898), .ZN(n4720) );
  INV_X1 U2886 ( .A(n2872), .ZN(n4727) );
  NAND2_X1 U2887 ( .A1(n2368), .A2(n2367), .ZN(n4686) );
  XNOR2_X1 U2888 ( .A(n4115), .B(n4114), .ZN(n4127) );
  OR2_X1 U2889 ( .A1(n4143), .A2(n4491), .ZN(n3208) );
  AND2_X1 U2890 ( .A1(n2918), .A2(n2429), .ZN(n2919) );
  AND2_X1 U2891 ( .A1(n2830), .A2(n2431), .ZN(n2831) );
  NAND2_X1 U2892 ( .A1(n2916), .A2(n4759), .ZN(n2832) );
  AOI21_X1 U2893 ( .B1(n3842), .B2(n3843), .A(n3844), .ZN(n3880) );
  NAND2_X1 U2894 ( .A1(n2376), .A2(n2432), .ZN(n2524) );
  INV_X1 U2895 ( .A(IR_REG_31__SCAN_IN), .ZN(n2797) );
  NOR2_X1 U2896 ( .A1(n3760), .A2(n3759), .ZN(n2246) );
  OR2_X1 U2897 ( .A1(n3238), .A2(n2841), .ZN(n2247) );
  OR2_X1 U2898 ( .A1(n2398), .A2(n2401), .ZN(n2248) );
  NAND2_X1 U2899 ( .A1(n2685), .A2(n2684), .ZN(n4439) );
  OR2_X1 U2900 ( .A1(n3814), .A2(n3813), .ZN(n2249) );
  AND2_X1 U2901 ( .A1(n2301), .A2(n2304), .ZN(n2250) );
  OR2_X1 U2902 ( .A1(n2898), .A2(n2899), .ZN(n2251) );
  NAND2_X1 U2903 ( .A1(n2379), .A2(n2378), .ZN(n3812) );
  NAND2_X1 U2904 ( .A1(n2921), .A2(n3215), .ZN(n2252) );
  OR2_X1 U2905 ( .A1(n2801), .A2(n2427), .ZN(n2253) );
  OAI21_X1 U2906 ( .B1(n2493), .B2(n2289), .A(n2291), .ZN(n3367) );
  OR2_X1 U2907 ( .A1(n3761), .A2(n2415), .ZN(n2414) );
  NAND2_X1 U2908 ( .A1(n3003), .A2(n3002), .ZN(n2255) );
  OR2_X1 U2909 ( .A1(n3206), .A2(n3205), .ZN(n2256) );
  AND2_X1 U2910 ( .A1(n2385), .A2(n2383), .ZN(n2257) );
  INV_X1 U2911 ( .A(n3232), .ZN(n2285) );
  NAND2_X1 U2912 ( .A1(n3796), .A2(n3124), .ZN(n3795) );
  AND2_X1 U2913 ( .A1(n2983), .A2(n2374), .ZN(n2259) );
  AND2_X1 U2914 ( .A1(n2385), .A2(n2386), .ZN(n2260) );
  INV_X1 U2915 ( .A(IR_REG_28__SCAN_IN), .ZN(n2755) );
  INV_X1 U2916 ( .A(n3935), .ZN(n3195) );
  OR2_X1 U2917 ( .A1(n3133), .A2(n3129), .ZN(n2261) );
  INV_X1 U2918 ( .A(n2414), .ZN(n2413) );
  NAND2_X1 U2919 ( .A1(n4150), .A2(n3974), .ZN(n2262) );
  INV_X1 U2920 ( .A(IR_REG_22__SCAN_IN), .ZN(n2451) );
  NOR2_X1 U2921 ( .A1(n4079), .A2(n3555), .ZN(n2263) );
  AND2_X1 U2922 ( .A1(n2335), .A2(n3974), .ZN(n2264) );
  AND2_X1 U2923 ( .A1(n2456), .A2(n2755), .ZN(n2265) );
  AND2_X1 U2924 ( .A1(n2370), .A2(n2251), .ZN(n2266) );
  AND2_X1 U2925 ( .A1(n2395), .A2(n2249), .ZN(n2267) );
  INV_X1 U2926 ( .A(n4565), .ZN(n2372) );
  INV_X1 U2927 ( .A(n3955), .ZN(n2336) );
  INV_X1 U2928 ( .A(n3823), .ZN(n2424) );
  INV_X1 U2929 ( .A(n4004), .ZN(n2325) );
  OR2_X1 U2930 ( .A1(n3149), .A2(n3148), .ZN(n2268) );
  OR2_X1 U2931 ( .A1(n4273), .A2(n4256), .ZN(n2269) );
  INV_X1 U2932 ( .A(n2294), .ZN(n4314) );
  NOR2_X1 U2933 ( .A1(n4479), .A2(n4468), .ZN(n2270) );
  AND2_X1 U2934 ( .A1(n3681), .A2(n3741), .ZN(n2271) );
  AND2_X1 U2935 ( .A1(n2358), .A2(n2357), .ZN(n2272) );
  INV_X1 U2936 ( .A(n2423), .ZN(n2417) );
  NAND2_X1 U2937 ( .A1(n2268), .A2(n3824), .ZN(n2423) );
  NAND2_X1 U2938 ( .A1(n2237), .A2(n3730), .ZN(n2273) );
  AND2_X1 U2939 ( .A1(n2390), .A2(n3098), .ZN(n2274) );
  INV_X1 U2940 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2343) );
  INV_X1 U2941 ( .A(n4013), .ZN(n2303) );
  INV_X1 U2942 ( .A(n2757), .ZN(n3990) );
  INV_X1 U2943 ( .A(n2487), .ZN(n2461) );
  INV_X1 U2944 ( .A(n4026), .ZN(n2317) );
  INV_X1 U2945 ( .A(n3843), .ZN(n2389) );
  INV_X1 U2946 ( .A(n4292), .ZN(n4438) );
  INV_X1 U2947 ( .A(n4018), .ZN(n2304) );
  INV_X1 U2948 ( .A(REG2_REG_6__SCAN_IN), .ZN(n2351) );
  OR2_X1 U2949 ( .A1(REG1_REG_17__SCAN_IN), .A2(n2901), .ZN(n2275) );
  NAND2_X1 U2950 ( .A1(n2457), .A2(n2456), .ZN(n2754) );
  NOR2_X1 U2951 ( .A1(n3486), .A2(n3516), .ZN(n2828) );
  NAND2_X1 U2952 ( .A1(n3059), .A2(n3060), .ZN(n2276) );
  INV_X1 U2953 ( .A(IR_REG_10__SCAN_IN), .ZN(n2296) );
  INV_X1 U2954 ( .A(IR_REG_20__SCAN_IN), .ZN(n2743) );
  INV_X1 U2955 ( .A(IR_REG_3__SCAN_IN), .ZN(n2512) );
  INV_X1 U2956 ( .A(n3434), .ZN(n2282) );
  NAND2_X1 U2957 ( .A1(n2283), .A2(n2502), .ZN(n3434) );
  NAND2_X1 U2958 ( .A1(n3370), .A2(n2501), .ZN(n2283) );
  NOR2_X1 U2959 ( .A1(n2285), .A2(n4558), .ZN(n2477) );
  XNOR2_X2 U2960 ( .A(n2284), .B(IR_REG_30__SCAN_IN), .ZN(n4558) );
  OAI21_X2 U2961 ( .B1(n4165), .B2(n2723), .A(n2722), .ZN(n4149) );
  OAI21_X2 U2962 ( .B1(n4183), .B2(n2710), .A(n2709), .ZN(n4165) );
  NAND2_X1 U2963 ( .A1(n4199), .A2(n2702), .ZN(n2286) );
  OAI22_X2 U2964 ( .A1(n3465), .A2(n2537), .B1(n3497), .B2(n4082), .ZN(n3493)
         );
  NAND2_X1 U2965 ( .A1(n3143), .A2(n2949), .ZN(n2946) );
  AND2_X1 U2966 ( .A1(n2489), .A2(n2488), .ZN(n2288) );
  NAND2_X1 U2967 ( .A1(n2290), .A2(n2491), .ZN(n2500) );
  NOR2_X2 U2968 ( .A1(n3389), .A2(n3390), .ZN(n3392) );
  INV_X1 U2969 ( .A(n2828), .ZN(n3580) );
  NAND2_X1 U2970 ( .A1(n2828), .A2(n2292), .ZN(n3582) );
  INV_X1 U2971 ( .A(n3579), .ZN(n2292) );
  NAND2_X1 U2972 ( .A1(n2425), .A2(n2749), .ZN(n2293) );
  NAND2_X1 U2973 ( .A1(n2866), .A2(n2755), .ZN(n2454) );
  AND2_X2 U2974 ( .A1(n2515), .A2(n2512), .ZN(n2432) );
  NAND4_X1 U2975 ( .A1(n2298), .A2(n2295), .A3(n2258), .A4(n2446), .ZN(n2450)
         );
  INV_X1 U2976 ( .A(n2769), .ZN(n2299) );
  NAND2_X1 U2977 ( .A1(n2299), .A2(n4013), .ZN(n2300) );
  NAND2_X1 U2978 ( .A1(n2300), .A2(n2250), .ZN(n2770) );
  NAND2_X1 U2979 ( .A1(n2305), .A2(n2306), .ZN(n2790) );
  NAND2_X1 U2980 ( .A1(n2780), .A2(n2308), .ZN(n2305) );
  OAI21_X1 U2981 ( .B1(n2771), .B2(n2315), .A(n2312), .ZN(n3734) );
  INV_X1 U2982 ( .A(n2319), .ZN(n2459) );
  NAND2_X1 U2983 ( .A1(n3437), .A2(n2321), .ZN(n2320) );
  XNOR2_X1 U2984 ( .A(n2337), .B(n2336), .ZN(n3201) );
  INV_X1 U2985 ( .A(n3218), .ZN(n2344) );
  INV_X1 U2986 ( .A(n2840), .ZN(n2346) );
  NAND2_X1 U2987 ( .A1(n2843), .A2(n4565), .ZN(n2354) );
  AOI22_X1 U2988 ( .A1(n3258), .A2(n2349), .B1(n2843), .B2(n2348), .ZN(n2353)
         );
  INV_X1 U2989 ( .A(n2353), .ZN(n3244) );
  XNOR2_X1 U2990 ( .A(n2854), .B(n4723), .ZN(n4653) );
  OAI21_X1 U2991 ( .B1(n4653), .B2(n2356), .A(n2355), .ZN(n4660) );
  INV_X2 U2992 ( .A(IR_REG_1__SCAN_IN), .ZN(n5057) );
  AND2_X1 U2993 ( .A1(n2366), .A2(n2365), .ZN(n2364) );
  NAND2_X1 U2994 ( .A1(n3334), .A2(n3335), .ZN(n2365) );
  OR2_X1 U2995 ( .A1(n3334), .A2(n3335), .ZN(n2366) );
  INV_X1 U2996 ( .A(n2370), .ZN(n4674) );
  NAND2_X1 U2997 ( .A1(n3842), .A2(n2380), .ZN(n2379) );
  NAND2_X1 U2998 ( .A1(n3114), .A2(n3113), .ZN(n2395) );
  NAND2_X1 U2999 ( .A1(n2395), .A2(n2394), .ZN(n3796) );
  NAND2_X1 U3000 ( .A1(n3024), .A2(n2248), .ZN(n2397) );
  NAND2_X1 U3001 ( .A1(n3029), .A2(n2404), .ZN(n2403) );
  INV_X1 U3002 ( .A(n3589), .ZN(n2404) );
  NAND2_X1 U3003 ( .A1(n3822), .A2(n2409), .ZN(n2405) );
  OAI211_X1 U3004 ( .C1(n3822), .C2(n2411), .A(n2405), .B(n2406), .ZN(n3777)
         );
  NAND2_X1 U3005 ( .A1(n3822), .A2(n2417), .ZN(n2416) );
  NAND2_X1 U3006 ( .A1(n2749), .A2(n2451), .ZN(n2801) );
  MUX2_X2 U3007 ( .A(n2455), .B(n2454), .S(n2456), .Z(n2493) );
  NAND2_X1 U3008 ( .A1(n2444), .A2(n2437), .ZN(n2668) );
  INV_X1 U3009 ( .A(n2609), .ZN(n2443) );
  NAND2_X1 U3010 ( .A1(n2478), .A2(REG0_REG_0__SCAN_IN), .ZN(n2482) );
  NAND2_X1 U3011 ( .A1(n2238), .A2(REG0_REG_1__SCAN_IN), .ZN(n2469) );
  OR2_X1 U3012 ( .A1(n4770), .A2(n2917), .ZN(n2429) );
  INV_X1 U3013 ( .A(n4586), .ZN(n3185) );
  AND2_X2 U3014 ( .A1(n3315), .A2(n4369), .ZN(n4713) );
  INV_X1 U3015 ( .A(n4629), .ZN(n2851) );
  OR2_X1 U3016 ( .A1(n4759), .A2(n2829), .ZN(n2431) );
  OR2_X1 U3017 ( .A1(n3215), .A2(n2928), .ZN(n2434) );
  INV_X1 U3018 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2559) );
  NOR2_X1 U3019 ( .A1(n2570), .A2(n3538), .ZN(n2435) );
  OR2_X1 U3020 ( .A1(n4075), .A2(n3708), .ZN(n2436) );
  AND3_X1 U3021 ( .A1(n2448), .A2(n5042), .A3(n5040), .ZN(n2437) );
  AND2_X1 U3022 ( .A1(n2611), .A2(n4861), .ZN(n2438) );
  INV_X1 U3023 ( .A(n3751), .ZN(n3063) );
  INV_X1 U3024 ( .A(n3706), .ZN(n3048) );
  AND2_X1 U3025 ( .A1(n3947), .A2(n4200), .ZN(n4045) );
  AND2_X1 U3026 ( .A1(n3975), .A2(n4166), .ZN(n4053) );
  INV_X1 U3027 ( .A(IR_REG_27__SCAN_IN), .ZN(n2456) );
  INV_X1 U3028 ( .A(n3132), .ZN(n3129) );
  INV_X1 U3029 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4861) );
  INV_X1 U3030 ( .A(n4608), .ZN(n2847) );
  AND2_X1 U3031 ( .A1(n4576), .A2(n4454), .ZN(n2660) );
  INV_X1 U3032 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3259) );
  OR2_X1 U3033 ( .A1(n2866), .A2(n2755), .ZN(n2455) );
  INV_X1 U3034 ( .A(n2616), .ZN(n2444) );
  CLKBUF_X3 U3035 ( .A(n2958), .Z(n3764) );
  OR2_X1 U3036 ( .A1(n2713), .A2(n2711), .ZN(n2724) );
  OR2_X1 U3037 ( .A1(n2669), .A2(n4873), .ZN(n2677) );
  INV_X1 U3038 ( .A(n4102), .ZN(n2838) );
  AND2_X1 U3039 ( .A1(n4396), .A2(n3784), .ZN(n3935) );
  AND2_X1 U3040 ( .A1(n4279), .A2(n2784), .ZN(n4225) );
  AND2_X1 U3041 ( .A1(n2647), .A2(REG3_REG_18__SCAN_IN), .ZN(n2662) );
  AND2_X1 U3042 ( .A1(n2623), .A2(n3730), .ZN(n2624) );
  AND2_X1 U3043 ( .A1(n3917), .A2(n3918), .ZN(n3733) );
  NAND2_X1 U3044 ( .A1(n2583), .A2(REG3_REG_11__SCAN_IN), .ZN(n2593) );
  INV_X1 U3045 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4859) );
  AND2_X1 U3046 ( .A1(n2757), .A2(n4561), .ZN(n2863) );
  INV_X1 U3047 ( .A(n4271), .ZN(n4429) );
  INV_X1 U3048 ( .A(n3618), .ZN(n3592) );
  INV_X1 U3049 ( .A(n3301), .ZN(n3389) );
  INV_X1 U3050 ( .A(n3761), .ZN(n3155) );
  AND2_X1 U3051 ( .A1(n2572), .A2(REG3_REG_10__SCAN_IN), .ZN(n2583) );
  XNOR2_X1 U3052 ( .A(n2938), .B(n3766), .ZN(n2943) );
  OR2_X1 U3053 ( .A1(n2697), .A2(n5033), .ZN(n2713) );
  AND2_X1 U3054 ( .A1(n3094), .A2(n3093), .ZN(n3883) );
  OR2_X1 U3055 ( .A1(n4210), .A2(n2758), .ZN(n2701) );
  NAND2_X1 U3056 ( .A1(n2879), .A2(n4566), .ZN(n2880) );
  NAND2_X1 U3057 ( .A1(n3346), .A2(REG1_REG_4__SCAN_IN), .ZN(n3345) );
  INV_X1 U3058 ( .A(REG3_REG_12__SCAN_IN), .ZN(n3630) );
  NAND2_X1 U3059 ( .A1(n2853), .A2(n4632), .ZN(n4642) );
  AND2_X1 U3060 ( .A1(n4111), .A2(REG2_REG_18__SCAN_IN), .ZN(n4112) );
  INV_X1 U3061 ( .A(n4481), .ZN(n4411) );
  INV_X1 U3062 ( .A(n4430), .ZN(n4273) );
  AND2_X1 U3063 ( .A1(n3956), .A2(n4226), .ZN(n4264) );
  OR2_X1 U3064 ( .A1(n2548), .A2(n4859), .ZN(n2560) );
  INV_X1 U3065 ( .A(n3433), .ZN(n3967) );
  INV_X1 U3066 ( .A(n4177), .ZN(n3892) );
  INV_X1 U3067 ( .A(n4573), .ZN(n4377) );
  INV_X1 U3068 ( .A(n4478), .ZN(n4415) );
  OR2_X1 U3069 ( .A1(n2546), .A2(n2797), .ZN(n2555) );
  NAND2_X1 U3070 ( .A1(n3186), .A2(n3185), .ZN(n3187) );
  INV_X1 U3071 ( .A(n3795), .ZN(n3800) );
  OR2_X1 U3072 ( .A1(n2636), .A2(n4931), .ZN(n2646) );
  AND2_X1 U3073 ( .A1(n2687), .A2(REG3_REG_22__SCAN_IN), .ZN(n2691) );
  AND3_X1 U3074 ( .A1(n2701), .A2(n2700), .A3(n2699), .ZN(n4193) );
  AND2_X1 U3075 ( .A1(n2508), .A2(n2507), .ZN(n2509) );
  AND2_X1 U3076 ( .A1(n2906), .A2(n2865), .ZN(n4593) );
  AND2_X1 U3077 ( .A1(n4593), .A2(n2902), .ZN(n4684) );
  INV_X1 U3078 ( .A(n4362), .ZN(n4365) );
  NAND2_X1 U3079 ( .A1(n4063), .A2(n2794), .ZN(n4375) );
  INV_X1 U3080 ( .A(n4317), .ZN(n4707) );
  OR2_X1 U3081 ( .A1(n3786), .A2(n4491), .ZN(n2918) );
  INV_X1 U3082 ( .A(n4491), .ZN(n4408) );
  INV_X1 U3083 ( .A(n4559), .ZN(n2826) );
  AND2_X1 U3084 ( .A1(n2634), .A2(n2642), .ZN(n2870) );
  AND2_X1 U3085 ( .A1(n2906), .A2(n2905), .ZN(n4683) );
  AND2_X1 U3086 ( .A1(n3184), .A2(n3183), .ZN(n4586) );
  INV_X1 U3087 ( .A(n4396), .ZN(n4140) );
  OAI211_X1 U3088 ( .C1(n4239), .C2(n2758), .A(n2694), .B(n2693), .ZN(n4412)
         );
  NAND4_X1 U3089 ( .A1(n2641), .A2(n2640), .A3(n2639), .A4(n2638), .ZN(n4469)
         );
  NAND2_X1 U3090 ( .A1(n2912), .A2(n2911), .ZN(n2913) );
  NAND2_X1 U3091 ( .A1(n4209), .A2(n3399), .ZN(n4382) );
  NAND2_X1 U3092 ( .A1(n4770), .A2(n4738), .ZN(n4491) );
  OR2_X1 U3093 ( .A1(n2915), .A2(n3311), .ZN(n4767) );
  OR2_X1 U3094 ( .A1(n4143), .A2(n4556), .ZN(n3212) );
  NAND2_X1 U3095 ( .A1(n4759), .A2(n4738), .ZN(n4556) );
  OR2_X1 U3096 ( .A1(n2915), .A2(n2827), .ZN(n4757) );
  INV_X1 U3097 ( .A(n2894), .ZN(n4723) );
  NAND2_X1 U3098 ( .A1(n2832), .A2(n2831), .ZN(U3514) );
  NOR2_X1 U3099 ( .A1(n2567), .A2(n2449), .ZN(n2590) );
  NOR2_X1 U3100 ( .A1(IR_REG_12__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2441)
         );
  NAND2_X1 U3101 ( .A1(n2590), .A2(n2441), .ZN(n2609) );
  NAND2_X1 U3102 ( .A1(n2443), .A2(n2442), .ZN(n2616) );
  INV_X2 U3103 ( .A(IR_REG_15__SCAN_IN), .ZN(n5040) );
  NAND2_X1 U3104 ( .A1(n2668), .A2(IR_REG_31__SCAN_IN), .ZN(n2445) );
  XNOR2_X1 U3105 ( .A(n2445), .B(IR_REG_18__SCAN_IN), .ZN(n4111) );
  INV_X1 U3106 ( .A(DATAI_18_), .ZN(n4796) );
  MUX2_X1 U3107 ( .A(n4717), .B(n4796), .S(n2240), .Z(n4328) );
  INV_X1 U3108 ( .A(n4328), .ZN(n4331) );
  INV_X1 U3109 ( .A(IR_REG_29__SCAN_IN), .ZN(n2458) );
  NAND2_X1 U3110 ( .A1(n2459), .A2(n2458), .ZN(n3791) );
  NAND2_X1 U3111 ( .A1(n2715), .A2(REG0_REG_18__SCAN_IN), .ZN(n2466) );
  NAND2_X1 U3112 ( .A1(n2735), .A2(REG1_REG_18__SCAN_IN), .ZN(n2465) );
  INV_X1 U3113 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2602) );
  INV_X1 U3114 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4931) );
  INV_X1 U3115 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2645) );
  NOR2_X1 U3116 ( .A1(n2647), .A2(REG3_REG_18__SCAN_IN), .ZN(n2462) );
  OR2_X1 U3117 ( .A1(n2662), .A2(n2462), .ZN(n4337) );
  OR2_X1 U3118 ( .A1(n2758), .A2(n4337), .ZN(n2464) );
  INV_X1 U3119 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4338) );
  OR2_X1 U3120 ( .A1(n3915), .A2(n4338), .ZN(n2463) );
  NAND2_X1 U3121 ( .A1(n2477), .A2(REG1_REG_1__SCAN_IN), .ZN(n2471) );
  INV_X1 U3122 ( .A(n2479), .ZN(n2467) );
  NAND2_X1 U3123 ( .A1(n2467), .A2(REG2_REG_1__SCAN_IN), .ZN(n2470) );
  NAND2_X1 U3124 ( .A1(n2239), .A2(REG3_REG_1__SCAN_IN), .ZN(n2468) );
  NAND2_X1 U3125 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2472)
         );
  NAND2_X1 U3126 ( .A1(n2474), .A2(n2473), .ZN(n4091) );
  INV_X1 U3127 ( .A(DATAI_1_), .ZN(n2475) );
  MUX2_X1 U3128 ( .A(n4091), .B(n2475), .S(n2493), .Z(n3359) );
  NAND2_X1 U3129 ( .A1(n2934), .A2(n3359), .ZN(n3993) );
  NAND2_X1 U3130 ( .A1(n3912), .A2(REG1_REG_0__SCAN_IN), .ZN(n2483) );
  INV_X1 U3131 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3317) );
  INV_X1 U3132 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3327) );
  OR2_X1 U3133 ( .A1(n2479), .A2(n3327), .ZN(n2480) );
  NAND4_X2 U3134 ( .A1(n2483), .A2(n2482), .A3(n2481), .A4(n2480), .ZN(n2925)
         );
  AND2_X1 U3135 ( .A1(n2925), .A2(n3367), .ZN(n3355) );
  CLKBUF_X1 U3136 ( .A(n2934), .Z(n2484) );
  NAND2_X1 U3137 ( .A1(n2484), .A2(n2935), .ZN(n2485) );
  AND2_X2 U3138 ( .A1(n3354), .A2(n2485), .ZN(n3380) );
  NAND2_X1 U3139 ( .A1(n3912), .A2(REG1_REG_2__SCAN_IN), .ZN(n2490) );
  NAND2_X1 U3140 ( .A1(n2478), .A2(REG0_REG_2__SCAN_IN), .ZN(n2489) );
  INV_X1 U3141 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2486) );
  OR2_X1 U3142 ( .A1(n2487), .A2(n2486), .ZN(n2488) );
  INV_X1 U3143 ( .A(DATAI_2_), .ZN(n2494) );
  MUX2_X1 U3144 ( .A(n3333), .B(n2494), .S(n2493), .Z(n3301) );
  NAND2_X1 U3145 ( .A1(n2949), .A2(n3301), .ZN(n3999) );
  NAND2_X1 U3146 ( .A1(n3996), .A2(n3999), .ZN(n3957) );
  OR2_X1 U3147 ( .A1(n2949), .A2(n3389), .ZN(n2495) );
  NAND2_X1 U31480 ( .A1(n2735), .A2(REG1_REG_3__SCAN_IN), .ZN(n2499) );
  NAND2_X1 U31490 ( .A1(n2715), .A2(REG0_REG_3__SCAN_IN), .ZN(n2498) );
  OR2_X1 U3150 ( .A1(n2758), .A2(REG3_REG_3__SCAN_IN), .ZN(n2497) );
  INV_X1 U3151 ( .A(REG2_REG_3__SCAN_IN), .ZN(n4104) );
  OR2_X1 U3152 ( .A1(n3915), .A2(n4104), .ZN(n2496) );
  NAND2_X1 U3153 ( .A1(n2500), .A2(IR_REG_31__SCAN_IN), .ZN(n2513) );
  XNOR2_X1 U3154 ( .A(n2513), .B(IR_REG_3__SCAN_IN), .ZN(n4102) );
  MUX2_X1 U3155 ( .A(n4102), .B(DATAI_3_), .S(n2493), .Z(n3374) );
  NAND2_X1 U3156 ( .A1(n4085), .A2(n3374), .ZN(n2501) );
  OR2_X1 U3157 ( .A1(n4085), .A2(n3374), .ZN(n2502) );
  NAND2_X1 U3158 ( .A1(n2735), .A2(REG1_REG_4__SCAN_IN), .ZN(n2511) );
  INV_X1 U3159 ( .A(REG2_REG_4__SCAN_IN), .ZN(n2841) );
  OR2_X1 U3160 ( .A1(n3915), .A2(n2841), .ZN(n2510) );
  INV_X1 U3161 ( .A(n2519), .ZN(n2506) );
  INV_X1 U3162 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2504) );
  INV_X1 U3163 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2503) );
  NAND2_X1 U3164 ( .A1(n2504), .A2(n2503), .ZN(n2505) );
  NAND2_X1 U3165 ( .A1(n2506), .A2(n2505), .ZN(n3447) );
  OR2_X1 U3166 ( .A1(n2758), .A2(n3447), .ZN(n2508) );
  NAND2_X1 U3167 ( .A1(n2715), .A2(REG0_REG_4__SCAN_IN), .ZN(n2507) );
  NAND2_X1 U3168 ( .A1(n2513), .A2(n2512), .ZN(n2514) );
  NAND2_X1 U3169 ( .A1(n2514), .A2(IR_REG_31__SCAN_IN), .ZN(n2516) );
  XNOR2_X1 U3170 ( .A(n2516), .B(n2515), .ZN(n3349) );
  INV_X1 U3171 ( .A(DATAI_4_), .ZN(n2517) );
  MUX2_X1 U3172 ( .A(n3349), .B(n2517), .S(n2240), .Z(n3445) );
  OR2_X1 U3173 ( .A1(n4084), .A2(n3445), .ZN(n4002) );
  NAND2_X1 U3174 ( .A1(n4084), .A2(n3445), .ZN(n4004) );
  INV_X1 U3175 ( .A(n3445), .ZN(n3438) );
  NAND2_X1 U3176 ( .A1(n4084), .A2(n3438), .ZN(n2518) );
  NAND2_X1 U3177 ( .A1(n3436), .A2(n2518), .ZN(n3400) );
  NAND2_X1 U3178 ( .A1(n2715), .A2(REG0_REG_5__SCAN_IN), .ZN(n2523) );
  NAND2_X1 U3179 ( .A1(n2735), .A2(REG1_REG_5__SCAN_IN), .ZN(n2522) );
  OAI21_X1 U3180 ( .B1(n2519), .B2(REG3_REG_5__SCAN_IN), .A(n2529), .ZN(n3837)
         );
  OR2_X1 U3181 ( .A1(n2758), .A2(n3837), .ZN(n2521) );
  OR2_X1 U3182 ( .A1(n3915), .A2(n2343), .ZN(n2520) );
  NAND4_X1 U3183 ( .A1(n2523), .A2(n2522), .A3(n2521), .A4(n2520), .ZN(n4083)
         );
  NAND2_X1 U3184 ( .A1(n2524), .A2(IR_REG_31__SCAN_IN), .ZN(n2525) );
  XNOR2_X1 U3185 ( .A(n2525), .B(IR_REG_5__SCAN_IN), .ZN(n3218) );
  MUX2_X1 U3186 ( .A(n3218), .B(DATAI_5_), .S(n2240), .Z(n3836) );
  OR2_X1 U3187 ( .A1(n4083), .A2(n3836), .ZN(n2526) );
  NAND2_X1 U3188 ( .A1(n3400), .A2(n2526), .ZN(n2528) );
  NAND2_X1 U3189 ( .A1(n4083), .A2(n3836), .ZN(n2527) );
  NAND2_X1 U3190 ( .A1(n2715), .A2(REG0_REG_6__SCAN_IN), .ZN(n2534) );
  NAND2_X1 U3191 ( .A1(n2735), .A2(REG1_REG_6__SCAN_IN), .ZN(n2533) );
  AND2_X1 U3192 ( .A1(n2529), .A2(n3259), .ZN(n2530) );
  OR2_X1 U3193 ( .A1(n2530), .A2(n2538), .ZN(n3471) );
  OR2_X1 U3194 ( .A1(n2758), .A2(n3471), .ZN(n2532) );
  OR2_X1 U3195 ( .A1(n3915), .A2(n2351), .ZN(n2531) );
  OR2_X1 U3196 ( .A1(n2535), .A2(n2797), .ZN(n2536) );
  XNOR2_X1 U3197 ( .A(n2536), .B(IR_REG_6__SCAN_IN), .ZN(n4565) );
  MUX2_X1 U3198 ( .A(n4565), .B(DATAI_6_), .S(n2240), .Z(n3497) );
  AND2_X1 U3199 ( .A1(n4082), .A2(n3497), .ZN(n2537) );
  NAND2_X1 U3200 ( .A1(n2715), .A2(REG0_REG_7__SCAN_IN), .ZN(n2544) );
  NAND2_X1 U3201 ( .A1(n2735), .A2(REG1_REG_7__SCAN_IN), .ZN(n2543) );
  OR2_X1 U3202 ( .A1(n2538), .A2(REG3_REG_7__SCAN_IN), .ZN(n2539) );
  NAND2_X1 U3203 ( .A1(n2548), .A2(n2539), .ZN(n3519) );
  OR2_X1 U3204 ( .A1(n2758), .A2(n3519), .ZN(n2542) );
  INV_X1 U3205 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2540) );
  OR2_X1 U3206 ( .A1(n3915), .A2(n2540), .ZN(n2541) );
  NAND4_X1 U3207 ( .A1(n2544), .A2(n2543), .A3(n2542), .A4(n2541), .ZN(n4081)
         );
  AND2_X1 U3208 ( .A1(n2535), .A2(n2545), .ZN(n2546) );
  XNOR2_X1 U3209 ( .A(n2555), .B(n2554), .ZN(n3254) );
  INV_X1 U32100 ( .A(DATAI_7_), .ZN(n2547) );
  MUX2_X1 U32110 ( .A(n3254), .B(n2547), .S(n2240), .Z(n2992) );
  OR2_X1 U32120 ( .A1(n4081), .A2(n2992), .ZN(n4006) );
  NAND2_X1 U32130 ( .A1(n4081), .A2(n2992), .ZN(n4012) );
  NAND2_X1 U32140 ( .A1(n4081), .A2(n3516), .ZN(n3571) );
  NAND2_X1 U32150 ( .A1(n2735), .A2(REG1_REG_8__SCAN_IN), .ZN(n2553) );
  NAND2_X1 U32160 ( .A1(n2715), .A2(REG0_REG_8__SCAN_IN), .ZN(n2552) );
  NAND2_X1 U32170 ( .A1(n2548), .A2(n4859), .ZN(n2549) );
  AND2_X1 U32180 ( .A1(n2560), .A2(n2549), .ZN(n4698) );
  INV_X1 U32190 ( .A(n4698), .ZN(n3533) );
  OR2_X1 U32200 ( .A1(n2758), .A2(n3533), .ZN(n2551) );
  INV_X1 U32210 ( .A(REG2_REG_8__SCAN_IN), .ZN(n2845) );
  OR2_X1 U32220 ( .A1(n3915), .A2(n2845), .ZN(n2550) );
  NAND2_X1 U32230 ( .A1(n2555), .A2(n2554), .ZN(n2556) );
  NAND2_X1 U32240 ( .A1(n2556), .A2(IR_REG_31__SCAN_IN), .ZN(n2557) );
  XNOR2_X1 U32250 ( .A(n2557), .B(IR_REG_8__SCAN_IN), .ZN(n4564) );
  MUX2_X1 U32260 ( .A(n4564), .B(DATAI_8_), .S(n2240), .Z(n3579) );
  NAND2_X1 U32270 ( .A1(n4080), .A2(n3579), .ZN(n2558) );
  AND2_X1 U32280 ( .A1(n3571), .A2(n2558), .ZN(n3537) );
  NAND2_X1 U32290 ( .A1(n2735), .A2(REG1_REG_9__SCAN_IN), .ZN(n2566) );
  NAND2_X1 U32300 ( .A1(n2715), .A2(REG0_REG_9__SCAN_IN), .ZN(n2565) );
  AND2_X1 U32310 ( .A1(n2560), .A2(n2559), .ZN(n2561) );
  OR2_X1 U32320 ( .A1(n2561), .A2(n2572), .ZN(n3558) );
  OR2_X1 U32330 ( .A1(n2758), .A2(n3558), .ZN(n2564) );
  INV_X1 U32340 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2562) );
  OR2_X1 U32350 ( .A1(n3915), .A2(n2562), .ZN(n2563) );
  NAND2_X1 U32360 ( .A1(n2567), .A2(IR_REG_31__SCAN_IN), .ZN(n2568) );
  XNOR2_X1 U32370 ( .A(n2568), .B(IR_REG_9__SCAN_IN), .ZN(n2874) );
  MUX2_X1 U32380 ( .A(n2874), .B(DATAI_9_), .S(n2240), .Z(n3555) );
  AND2_X1 U32390 ( .A1(n4079), .A2(n3555), .ZN(n2570) );
  INV_X1 U32400 ( .A(n2570), .ZN(n2569) );
  AND2_X1 U32410 ( .A1(n3537), .A2(n2569), .ZN(n2571) );
  OR2_X1 U32420 ( .A1(n4080), .A2(n3579), .ZN(n3538) );
  NAND2_X1 U32430 ( .A1(n2735), .A2(REG1_REG_10__SCAN_IN), .ZN(n2578) );
  NAND2_X1 U32440 ( .A1(n2715), .A2(REG0_REG_10__SCAN_IN), .ZN(n2577) );
  NOR2_X1 U32450 ( .A1(n2572), .A2(REG3_REG_10__SCAN_IN), .ZN(n2573) );
  OR2_X1 U32460 ( .A1(n2583), .A2(n2573), .ZN(n4690) );
  OR2_X1 U32470 ( .A1(n2758), .A2(n4690), .ZN(n2576) );
  INV_X1 U32480 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2574) );
  OR2_X1 U32490 ( .A1(n3915), .A2(n2574), .ZN(n2575) );
  OR2_X1 U32500 ( .A1(n2567), .A2(IR_REG_9__SCAN_IN), .ZN(n2579) );
  NAND2_X1 U32510 ( .A1(n2579), .A2(IR_REG_31__SCAN_IN), .ZN(n2580) );
  XNOR2_X1 U32520 ( .A(n2580), .B(IR_REG_10__SCAN_IN), .ZN(n4608) );
  MUX2_X1 U32530 ( .A(n4608), .B(DATAI_10_), .S(n2240), .Z(n3692) );
  OR2_X1 U32540 ( .A1(n4078), .A2(n3692), .ZN(n2582) );
  AND2_X1 U32550 ( .A1(n4078), .A2(n3692), .ZN(n2581) );
  AOI21_X1 U32560 ( .B1(n3690), .B2(n2582), .A(n2581), .ZN(n3611) );
  NAND2_X1 U32570 ( .A1(n2715), .A2(REG0_REG_11__SCAN_IN), .ZN(n2589) );
  NAND2_X1 U32580 ( .A1(n2735), .A2(REG1_REG_11__SCAN_IN), .ZN(n2588) );
  OR2_X1 U32590 ( .A1(n2583), .A2(REG3_REG_11__SCAN_IN), .ZN(n2584) );
  NAND2_X1 U32600 ( .A1(n2593), .A2(n2584), .ZN(n3620) );
  OR2_X1 U32610 ( .A1(n2758), .A2(n3620), .ZN(n2587) );
  INV_X1 U32620 ( .A(REG2_REG_11__SCAN_IN), .ZN(n2585) );
  OR2_X1 U32630 ( .A1(n3915), .A2(n2585), .ZN(n2586) );
  OR2_X1 U32640 ( .A1(n2590), .A2(n2797), .ZN(n2599) );
  XNOR2_X1 U32650 ( .A(n2599), .B(IR_REG_11__SCAN_IN), .ZN(n2872) );
  INV_X1 U32660 ( .A(DATAI_11_), .ZN(n2591) );
  MUX2_X1 U32670 ( .A(n4727), .B(n2591), .S(n2240), .Z(n3618) );
  OR2_X1 U32680 ( .A1(n4077), .A2(n3618), .ZN(n3644) );
  NAND2_X1 U32690 ( .A1(n4077), .A2(n3618), .ZN(n4026) );
  NAND2_X1 U32700 ( .A1(n3644), .A2(n4026), .ZN(n3968) );
  OR2_X1 U32710 ( .A1(n4077), .A2(n3592), .ZN(n2592) );
  NAND2_X1 U32720 ( .A1(n2715), .A2(REG0_REG_12__SCAN_IN), .ZN(n2598) );
  NAND2_X1 U32730 ( .A1(n2735), .A2(REG1_REG_12__SCAN_IN), .ZN(n2597) );
  NAND2_X1 U32740 ( .A1(n2593), .A2(n3630), .ZN(n2594) );
  NAND2_X1 U32750 ( .A1(n2603), .A2(n2594), .ZN(n3639) );
  OR2_X1 U32760 ( .A1(n2758), .A2(n3639), .ZN(n2596) );
  INV_X1 U32770 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3640) );
  OR2_X1 U32780 ( .A1(n3915), .A2(n3640), .ZN(n2595) );
  NAND4_X1 U32790 ( .A1(n2598), .A2(n2597), .A3(n2596), .A4(n2595), .ZN(n4076)
         );
  INV_X1 U32800 ( .A(IR_REG_11__SCAN_IN), .ZN(n4847) );
  NAND2_X1 U32810 ( .A1(n2599), .A2(n4847), .ZN(n2600) );
  NAND2_X1 U32820 ( .A1(n2600), .A2(IR_REG_31__SCAN_IN), .ZN(n2601) );
  XNOR2_X1 U32830 ( .A(n2601), .B(IR_REG_12__SCAN_IN), .ZN(n4629) );
  NAND2_X1 U32840 ( .A1(n4076), .A2(n3715), .ZN(n3664) );
  NAND2_X1 U32850 ( .A1(n2735), .A2(REG1_REG_13__SCAN_IN), .ZN(n2608) );
  NAND2_X1 U32860 ( .A1(n2715), .A2(REG0_REG_13__SCAN_IN), .ZN(n2607) );
  NAND2_X1 U32870 ( .A1(n2603), .A2(n2602), .ZN(n2604) );
  NAND2_X1 U32880 ( .A1(n2611), .A2(n2604), .ZN(n3711) );
  OR2_X1 U32890 ( .A1(n2758), .A2(n3711), .ZN(n2606) );
  INV_X1 U32900 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3683) );
  OR2_X1 U32910 ( .A1(n3915), .A2(n3683), .ZN(n2605) );
  NAND2_X1 U32920 ( .A1(n2609), .A2(IR_REG_31__SCAN_IN), .ZN(n2610) );
  XNOR2_X1 U32930 ( .A(n2610), .B(IR_REG_13__SCAN_IN), .ZN(n4724) );
  MUX2_X1 U32940 ( .A(n4724), .B(DATAI_13_), .S(n2240), .Z(n3708) );
  NAND2_X1 U32950 ( .A1(n4075), .A2(n3708), .ZN(n2620) );
  AND2_X1 U32960 ( .A1(n3664), .A2(n2620), .ZN(n3727) );
  NAND2_X1 U32970 ( .A1(n2715), .A2(REG0_REG_14__SCAN_IN), .ZN(n2615) );
  NAND2_X1 U32980 ( .A1(n2735), .A2(REG1_REG_14__SCAN_IN), .ZN(n2614) );
  OR2_X1 U32990 ( .A1(n2438), .A2(n2625), .ZN(n3755) );
  OR2_X1 U33000 ( .A1(n2758), .A2(n3755), .ZN(n2613) );
  INV_X1 U33010 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3743) );
  OR2_X1 U33020 ( .A1(n3915), .A2(n3743), .ZN(n2612) );
  NAND2_X1 U33030 ( .A1(n2617), .A2(IR_REG_31__SCAN_IN), .ZN(n2618) );
  XNOR2_X1 U33040 ( .A(n2618), .B(IR_REG_14__SCAN_IN), .ZN(n2894) );
  INV_X1 U33050 ( .A(DATAI_14_), .ZN(n4722) );
  MUX2_X1 U33060 ( .A(n4723), .B(n4722), .S(n2240), .Z(n3741) );
  NAND2_X1 U33070 ( .A1(n4467), .A2(n3741), .ZN(n3918) );
  INV_X1 U33080 ( .A(n3733), .ZN(n3949) );
  INV_X1 U33090 ( .A(n3741), .ZN(n4476) );
  OR2_X1 U33100 ( .A1(n4467), .A2(n4476), .ZN(n2623) );
  INV_X1 U33110 ( .A(n2620), .ZN(n2622) );
  OR2_X1 U33120 ( .A1(n4076), .A2(n3715), .ZN(n3665) );
  AND2_X1 U33130 ( .A1(n3665), .A2(n2436), .ZN(n2621) );
  NAND2_X1 U33140 ( .A1(n3731), .A2(n2624), .ZN(n3654) );
  NAND2_X1 U33150 ( .A1(n2715), .A2(REG0_REG_15__SCAN_IN), .ZN(n2631) );
  NAND2_X1 U33160 ( .A1(n2735), .A2(REG1_REG_15__SCAN_IN), .ZN(n2630) );
  OR2_X1 U33170 ( .A1(n2625), .A2(REG3_REG_15__SCAN_IN), .ZN(n2626) );
  NAND2_X1 U33180 ( .A1(n2636), .A2(n2626), .ZN(n3908) );
  OR2_X1 U33190 ( .A1(n2758), .A2(n3908), .ZN(n2629) );
  INV_X1 U33200 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2627) );
  OR2_X1 U33210 ( .A1(n3915), .A2(n2627), .ZN(n2628) );
  NAND2_X1 U33220 ( .A1(n2632), .A2(IR_REG_31__SCAN_IN), .ZN(n2656) );
  INV_X1 U33230 ( .A(n2656), .ZN(n2633) );
  NAND2_X1 U33240 ( .A1(n2633), .A2(IR_REG_15__SCAN_IN), .ZN(n2634) );
  NAND2_X1 U33250 ( .A1(n2656), .A2(n5040), .ZN(n2642) );
  MUX2_X1 U33260 ( .A(n2870), .B(DATAI_15_), .S(n2240), .Z(n4468) );
  NAND2_X1 U33270 ( .A1(n4479), .A2(n4468), .ZN(n2635) );
  NAND2_X1 U33280 ( .A1(n2735), .A2(REG1_REG_16__SCAN_IN), .ZN(n2641) );
  NAND2_X1 U33290 ( .A1(n2715), .A2(REG0_REG_16__SCAN_IN), .ZN(n2640) );
  NAND2_X1 U33300 ( .A1(n2636), .A2(n4931), .ZN(n2637) );
  NAND2_X1 U33310 ( .A1(n2646), .A2(n2637), .ZN(n4585) );
  OR2_X1 U33320 ( .A1(n2758), .A2(n4585), .ZN(n2639) );
  INV_X1 U33330 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4370) );
  OR2_X1 U33340 ( .A1(n3915), .A2(n4370), .ZN(n2638) );
  NAND2_X1 U33350 ( .A1(n2642), .A2(IR_REG_31__SCAN_IN), .ZN(n2643) );
  XNOR2_X1 U33360 ( .A(n2643), .B(IR_REG_16__SCAN_IN), .ZN(n2898) );
  INV_X1 U33370 ( .A(DATAI_16_), .ZN(n4719) );
  MUX2_X1 U33380 ( .A(n4720), .B(n4719), .S(n2240), .Z(n4573) );
  OR2_X1 U33390 ( .A1(n4469), .A2(n4573), .ZN(n4038) );
  NAND2_X1 U33400 ( .A1(n4469), .A2(n4573), .ZN(n4034) );
  NAND2_X1 U33410 ( .A1(n4038), .A2(n4034), .ZN(n4373) );
  NAND2_X1 U33420 ( .A1(n2735), .A2(REG1_REG_17__SCAN_IN), .ZN(n2653) );
  NAND2_X1 U33430 ( .A1(n2715), .A2(REG0_REG_17__SCAN_IN), .ZN(n2652) );
  AND2_X1 U33440 ( .A1(n2646), .A2(n2645), .ZN(n2648) );
  OR2_X1 U33450 ( .A1(n2648), .A2(n2647), .ZN(n4352) );
  OR2_X1 U33460 ( .A1(n2758), .A2(n4352), .ZN(n2651) );
  INV_X1 U33470 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2649) );
  OR2_X1 U33480 ( .A1(n3915), .A2(n2649), .ZN(n2650) );
  INV_X1 U33490 ( .A(n4576), .ZN(n4334) );
  OR2_X1 U33500 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2654)
         );
  NAND2_X1 U33510 ( .A1(IR_REG_31__SCAN_IN), .A2(n2654), .ZN(n2655) );
  NAND2_X1 U33520 ( .A1(n2656), .A2(n2655), .ZN(n2658) );
  INV_X1 U3353 ( .A(IR_REG_17__SCAN_IN), .ZN(n2657) );
  XNOR2_X1 U33540 ( .A(n2658), .B(n2657), .ZN(n2901) );
  INV_X1 U3355 ( .A(n2901), .ZN(n4718) );
  INV_X1 U3356 ( .A(DATAI_17_), .ZN(n2659) );
  MUX2_X1 U3357 ( .A(n4718), .B(n2659), .S(n2240), .Z(n4357) );
  NAND2_X1 U3358 ( .A1(n4334), .A2(n4357), .ZN(n2661) );
  INV_X1 U3359 ( .A(n4357), .ZN(n4454) );
  OR2_X1 U3360 ( .A1(n4455), .A2(n4328), .ZN(n4304) );
  NAND2_X1 U3361 ( .A1(n4455), .A2(n4328), .ZN(n4305) );
  NAND2_X1 U3362 ( .A1(n4304), .A2(n4305), .ZN(n4330) );
  NAND2_X1 U3363 ( .A1(n4324), .A2(n4330), .ZN(n4325) );
  NAND2_X1 U3364 ( .A1(n2735), .A2(REG1_REG_19__SCAN_IN), .ZN(n2667) );
  NAND2_X1 U3365 ( .A1(n2715), .A2(REG0_REG_19__SCAN_IN), .ZN(n2666) );
  OR2_X1 U3366 ( .A1(n2662), .A2(REG3_REG_19__SCAN_IN), .ZN(n2663) );
  NAND2_X1 U3367 ( .A1(n2669), .A2(n2663), .ZN(n4318) );
  OR2_X1 U3368 ( .A1(n2758), .A2(n4318), .ZN(n2665) );
  INV_X1 U3369 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4319) );
  OR2_X1 U3370 ( .A1(n3915), .A2(n4319), .ZN(n2664) );
  MUX2_X1 U3371 ( .A(n4563), .B(DATAI_19_), .S(n2240), .Z(n3806) );
  NOR2_X1 U3372 ( .A1(n4332), .A2(n3806), .ZN(n4283) );
  NAND2_X1 U3373 ( .A1(n4332), .A2(n3806), .ZN(n4284) );
  NAND2_X1 U3374 ( .A1(n2715), .A2(REG0_REG_20__SCAN_IN), .ZN(n2675) );
  NAND2_X1 U3375 ( .A1(n2735), .A2(REG1_REG_20__SCAN_IN), .ZN(n2674) );
  INV_X1 U3376 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4873) );
  NAND2_X1 U3377 ( .A1(n2669), .A2(n4873), .ZN(n2670) );
  NAND2_X1 U3378 ( .A1(n2677), .A2(n2670), .ZN(n4288) );
  OR2_X1 U3379 ( .A1(n2758), .A2(n4288), .ZN(n2673) );
  INV_X1 U3380 ( .A(REG2_REG_20__SCAN_IN), .ZN(n2671) );
  OR2_X1 U3381 ( .A1(n3915), .A2(n2671), .ZN(n2672) );
  NAND4_X1 U3382 ( .A1(n2675), .A2(n2674), .A3(n2673), .A4(n2672), .ZN(n4272)
         );
  NAND2_X1 U3383 ( .A1(n2240), .A2(DATAI_20_), .ZN(n4292) );
  NAND2_X1 U3384 ( .A1(n4272), .A2(n4438), .ZN(n3980) );
  OR2_X1 U3385 ( .A1(n4272), .A2(n4438), .ZN(n3981) );
  INV_X1 U3386 ( .A(REG3_REG_21__SCAN_IN), .ZN(n2676) );
  AND2_X1 U3387 ( .A1(n2677), .A2(n2676), .ZN(n2678) );
  OR2_X1 U3388 ( .A1(n2678), .A2(n2687), .ZN(n4268) );
  INV_X1 U3389 ( .A(REG2_REG_21__SCAN_IN), .ZN(n2679) );
  OR2_X1 U3390 ( .A1(n3915), .A2(n2679), .ZN(n2680) );
  OAI21_X1 U3391 ( .B1(n4268), .B2(n2758), .A(n2680), .ZN(n2681) );
  INV_X1 U3392 ( .A(n2681), .ZN(n2685) );
  NAND2_X1 U3393 ( .A1(n2715), .A2(REG0_REG_21__SCAN_IN), .ZN(n2683) );
  NAND2_X1 U3394 ( .A1(n2735), .A2(REG1_REG_21__SCAN_IN), .ZN(n2682) );
  NAND2_X1 U3395 ( .A1(n2240), .A2(DATAI_21_), .ZN(n4271) );
  NAND2_X1 U3396 ( .A1(n4439), .A2(n4429), .ZN(n2686) );
  INV_X1 U3397 ( .A(n4439), .ZN(n4294) );
  NOR2_X1 U3398 ( .A1(n2687), .A2(REG3_REG_22__SCAN_IN), .ZN(n2688) );
  OR2_X1 U3399 ( .A1(n2691), .A2(n2688), .ZN(n4248) );
  AOI22_X1 U3400 ( .A1(n2735), .A2(REG1_REG_22__SCAN_IN), .B1(n2715), .B2(
        REG0_REG_22__SCAN_IN), .ZN(n2690) );
  INV_X1 U3401 ( .A(REG2_REG_22__SCAN_IN), .ZN(n4249) );
  OR2_X1 U3402 ( .A1(n3915), .A2(n4249), .ZN(n2689) );
  OAI211_X1 U3403 ( .C1(n4248), .C2(n2758), .A(n2690), .B(n2689), .ZN(n4430)
         );
  NAND2_X1 U3404 ( .A1(n2240), .A2(DATAI_22_), .ZN(n4256) );
  OR2_X1 U3405 ( .A1(n4430), .A2(n4256), .ZN(n4228) );
  NAND2_X1 U3406 ( .A1(n4430), .A2(n4256), .ZN(n2787) );
  NAND2_X1 U3407 ( .A1(n4228), .A2(n2787), .ZN(n4252) );
  OR2_X1 U3408 ( .A1(n2691), .A2(REG3_REG_23__SCAN_IN), .ZN(n2692) );
  NAND2_X1 U3409 ( .A1(n2697), .A2(n2692), .ZN(n4239) );
  AOI22_X1 U3410 ( .A1(n2735), .A2(REG1_REG_23__SCAN_IN), .B1(n2715), .B2(
        REG0_REG_23__SCAN_IN), .ZN(n2694) );
  INV_X1 U3411 ( .A(REG2_REG_23__SCAN_IN), .ZN(n4240) );
  OR2_X1 U3412 ( .A1(n3915), .A2(n4240), .ZN(n2693) );
  INV_X1 U3413 ( .A(n4412), .ZN(n4212) );
  NAND2_X1 U3414 ( .A1(n2240), .A2(DATAI_23_), .ZN(n4236) );
  NAND2_X1 U3415 ( .A1(n4212), .A2(n4236), .ZN(n2696) );
  NOR2_X1 U3416 ( .A1(n4212), .A2(n4236), .ZN(n2695) );
  INV_X1 U3417 ( .A(REG3_REG_24__SCAN_IN), .ZN(n5033) );
  NAND2_X1 U3418 ( .A1(n2697), .A2(n5033), .ZN(n2698) );
  NAND2_X1 U3419 ( .A1(n2713), .A2(n2698), .ZN(n4210) );
  AOI22_X1 U3420 ( .A1(n2735), .A2(REG1_REG_24__SCAN_IN), .B1(n2715), .B2(
        REG0_REG_24__SCAN_IN), .ZN(n2700) );
  INV_X1 U3421 ( .A(REG2_REG_24__SCAN_IN), .ZN(n4208) );
  OR2_X1 U3422 ( .A1(n3915), .A2(n4208), .ZN(n2699) );
  NAND2_X1 U3423 ( .A1(n2240), .A2(DATAI_24_), .ZN(n4207) );
  INV_X1 U3424 ( .A(n4207), .ZN(n4410) );
  NAND2_X1 U3425 ( .A1(n4233), .A2(n4410), .ZN(n2702) );
  NAND2_X1 U3426 ( .A1(n4193), .A2(n4207), .ZN(n2703) );
  XNOR2_X1 U3427 ( .A(n2713), .B(REG3_REG_25__SCAN_IN), .ZN(n4185) );
  NAND2_X1 U3428 ( .A1(n4185), .A2(n2461), .ZN(n2708) );
  INV_X1 U3429 ( .A(REG2_REG_25__SCAN_IN), .ZN(n4186) );
  NAND2_X1 U3430 ( .A1(n2735), .A2(REG1_REG_25__SCAN_IN), .ZN(n2705) );
  NAND2_X1 U3431 ( .A1(n2715), .A2(REG0_REG_25__SCAN_IN), .ZN(n2704) );
  OAI211_X1 U3432 ( .C1(n4186), .C2(n3915), .A(n2705), .B(n2704), .ZN(n2706)
         );
  INV_X1 U3433 ( .A(n2706), .ZN(n2707) );
  NAND2_X1 U3434 ( .A1(n2240), .A2(DATAI_25_), .ZN(n3827) );
  NOR2_X1 U3435 ( .A1(n4211), .A2(n4190), .ZN(n2710) );
  NAND2_X1 U3436 ( .A1(n4211), .A2(n4190), .ZN(n2709) );
  NAND2_X1 U3437 ( .A1(REG3_REG_25__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2711) );
  INV_X1 U3438 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3826) );
  INV_X1 U3439 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2712) );
  OAI21_X1 U3440 ( .B1(n2713), .B2(n3826), .A(n2712), .ZN(n2714) );
  NAND2_X1 U3441 ( .A1(n4178), .A2(n2461), .ZN(n2721) );
  INV_X1 U3442 ( .A(REG2_REG_26__SCAN_IN), .ZN(n2718) );
  NAND2_X1 U3443 ( .A1(n2715), .A2(REG0_REG_26__SCAN_IN), .ZN(n2717) );
  NAND2_X1 U3444 ( .A1(n2735), .A2(REG1_REG_26__SCAN_IN), .ZN(n2716) );
  OAI211_X1 U3445 ( .C1(n2718), .C2(n3915), .A(n2717), .B(n2716), .ZN(n2719)
         );
  INV_X1 U3446 ( .A(n2719), .ZN(n2720) );
  NAND2_X1 U3447 ( .A1(n2240), .A2(DATAI_26_), .ZN(n4177) );
  NOR2_X1 U3448 ( .A1(n4157), .A2(n4177), .ZN(n2723) );
  NAND2_X1 U3449 ( .A1(n4157), .A2(n4177), .ZN(n2722) );
  INV_X1 U3450 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3174) );
  AND2_X1 U3451 ( .A1(n2724), .A2(n3174), .ZN(n2725) );
  INV_X1 U3452 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4155) );
  NAND2_X1 U3453 ( .A1(n2735), .A2(REG1_REG_27__SCAN_IN), .ZN(n2727) );
  NAND2_X1 U3454 ( .A1(n2715), .A2(REG0_REG_27__SCAN_IN), .ZN(n2726) );
  OAI211_X1 U3455 ( .C1(n4155), .C2(n3915), .A(n2727), .B(n2726), .ZN(n2728)
         );
  INV_X1 U3456 ( .A(n2728), .ZN(n2729) );
  OAI21_X1 U3457 ( .B1(n4156), .B2(n2758), .A(n2729), .ZN(n4074) );
  NAND2_X1 U34580 ( .A1(n2240), .A2(DATAI_27_), .ZN(n4154) );
  INV_X1 U34590 ( .A(n4154), .ZN(n4392) );
  NOR2_X1 U3460 ( .A1(n4074), .A2(n4392), .ZN(n2731) );
  NAND2_X1 U3461 ( .A1(n4074), .A2(n4392), .ZN(n2730) );
  NAND2_X1 U3462 ( .A1(n2732), .A2(REG3_REG_28__SCAN_IN), .ZN(n4142) );
  INV_X1 U3463 ( .A(n2732), .ZN(n2733) );
  INV_X1 U3464 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3772) );
  NAND2_X1 U3465 ( .A1(n2733), .A2(n3772), .ZN(n2734) );
  NAND2_X1 U3466 ( .A1(n4142), .A2(n2734), .ZN(n3780) );
  INV_X1 U34670 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3779) );
  NAND2_X1 U3468 ( .A1(n2715), .A2(REG0_REG_28__SCAN_IN), .ZN(n2737) );
  NAND2_X1 U34690 ( .A1(n2735), .A2(REG1_REG_28__SCAN_IN), .ZN(n2736) );
  OAI211_X1 U3470 ( .C1(n3779), .C2(n3915), .A(n2737), .B(n2736), .ZN(n2738)
         );
  INV_X1 U34710 ( .A(n2738), .ZN(n2739) );
  NAND2_X1 U3472 ( .A1(n2240), .A2(DATAI_28_), .ZN(n3771) );
  INV_X1 U34730 ( .A(n3771), .ZN(n3784) );
  NAND2_X1 U3474 ( .A1(n4140), .A2(n3771), .ZN(n3194) );
  NAND2_X1 U34750 ( .A1(n3195), .A2(n3194), .ZN(n3953) );
  XNOR2_X1 U3476 ( .A(n3192), .B(n3953), .ZN(n3790) );
  NAND2_X1 U34770 ( .A1(n2746), .A2(n2741), .ZN(n2742) );
  OAI21_X1 U3478 ( .B1(IR_REG_19__SCAN_IN), .B2(IR_REG_20__SCAN_IN), .A(
        IR_REG_31__SCAN_IN), .ZN(n2745) );
  NAND2_X1 U34790 ( .A1(n2746), .A2(n2745), .ZN(n2748) );
  XNOR2_X2 U3480 ( .A(n2748), .B(n2747), .ZN(n2757) );
  INV_X1 U34810 ( .A(n2749), .ZN(n2750) );
  NAND2_X1 U3482 ( .A1(n2750), .A2(IR_REG_31__SCAN_IN), .ZN(n2751) );
  XNOR2_X1 U34830 ( .A(n2921), .B(n4561), .ZN(n2752) );
  NAND2_X1 U3484 ( .A1(n2752), .A2(n4123), .ZN(n3738) );
  NAND2_X1 U34850 ( .A1(n2242), .A2(n4563), .ZN(n3309) );
  NAND2_X1 U3486 ( .A1(n3738), .A2(n4733), .ZN(n4745) );
  INV_X1 U34870 ( .A(n4745), .ZN(n4452) );
  NAND2_X1 U3488 ( .A1(n2754), .A2(IR_REG_31__SCAN_IN), .ZN(n2756) );
  XNOR2_X1 U34890 ( .A(n2756), .B(n2755), .ZN(n4570) );
  INV_X1 U3490 ( .A(n2863), .ZN(n3162) );
  OR2_X1 U34910 ( .A1(n4142), .A2(n2758), .ZN(n2763) );
  INV_X1 U3492 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4137) );
  NAND2_X1 U34930 ( .A1(n2715), .A2(REG0_REG_29__SCAN_IN), .ZN(n2760) );
  NAND2_X1 U3494 ( .A1(n2735), .A2(REG1_REG_29__SCAN_IN), .ZN(n2759) );
  OAI211_X1 U34950 ( .C1(n4137), .C2(n3915), .A(n2760), .B(n2759), .ZN(n2761)
         );
  INV_X1 U3496 ( .A(n2761), .ZN(n2762) );
  NAND2_X1 U34970 ( .A1(n2763), .A2(n2762), .ZN(n4073) );
  INV_X1 U3498 ( .A(n4073), .ZN(n3781) );
  INV_X1 U34990 ( .A(n4561), .ZN(n2930) );
  NAND2_X1 U3500 ( .A1(n3990), .A2(n2930), .ZN(n3306) );
  OAI22_X1 U35010 ( .A1(n3781), .A2(n4415), .B1(n3771), .B2(n4309), .ZN(n2764)
         );
  AOI21_X1 U3502 ( .B1(n4411), .B2(n4074), .A(n2764), .ZN(n2796) );
  OR2_X1 U35030 ( .A1(n2925), .A2(n3307), .ZN(n3356) );
  INV_X1 U3504 ( .A(n3957), .ZN(n3381) );
  NAND2_X1 U35050 ( .A1(n3382), .A2(n3381), .ZN(n2766) );
  NAND2_X1 U35060 ( .A1(n2766), .A2(n3996), .ZN(n3372) );
  OR2_X1 U35070 ( .A1(n4085), .A2(n3421), .ZN(n4001) );
  NAND2_X1 U35080 ( .A1(n4085), .A2(n3421), .ZN(n3998) );
  AND2_X1 U35090 ( .A1(n4001), .A2(n3998), .ZN(n3371) );
  NAND2_X1 U35100 ( .A1(n3372), .A2(n3371), .ZN(n2767) );
  NAND2_X1 U35110 ( .A1(n2767), .A2(n4001), .ZN(n3437) );
  INV_X1 U35120 ( .A(n4002), .ZN(n2768) );
  INV_X1 U35130 ( .A(n3836), .ZN(n3478) );
  AND2_X1 U35140 ( .A1(n4083), .A2(n3478), .ZN(n4005) );
  OR2_X1 U35150 ( .A1(n4083), .A2(n3478), .ZN(n4020) );
  NAND2_X1 U35160 ( .A1(n4082), .A2(n3472), .ZN(n3462) );
  NOR2_X1 U35170 ( .A1(n4082), .A2(n3472), .ZN(n4007) );
  AOI21_X1 U35180 ( .B1(n3463), .B2(n3462), .A(n4007), .ZN(n3487) );
  NAND2_X1 U35190 ( .A1(n3487), .A2(n4006), .ZN(n2769) );
  OR2_X1 U35200 ( .A1(n4080), .A2(n2292), .ZN(n4013) );
  NAND2_X1 U35210 ( .A1(n4080), .A2(n2292), .ZN(n4011) );
  INV_X1 U35220 ( .A(n3555), .ZN(n3598) );
  AND2_X1 U35230 ( .A1(n4079), .A2(n3598), .ZN(n4018) );
  OR2_X1 U35240 ( .A1(n4079), .A2(n3598), .ZN(n4014) );
  NAND2_X1 U35250 ( .A1(n2770), .A2(n4014), .ZN(n3691) );
  NAND2_X1 U35260 ( .A1(n4078), .A2(n3689), .ZN(n4027) );
  NAND2_X1 U35270 ( .A1(n3691), .A2(n4027), .ZN(n2771) );
  OR2_X1 U35280 ( .A1(n4078), .A2(n3689), .ZN(n4022) );
  INV_X1 U35290 ( .A(n3715), .ZN(n2772) );
  NAND2_X1 U35300 ( .A1(n4076), .A2(n2772), .ZN(n3671) );
  NAND2_X1 U35310 ( .A1(n4075), .A2(n3681), .ZN(n3667) );
  NAND2_X1 U35320 ( .A1(n3671), .A2(n3667), .ZN(n4028) );
  INV_X1 U35330 ( .A(n4028), .ZN(n2775) );
  OR2_X1 U35340 ( .A1(n4076), .A2(n2772), .ZN(n3670) );
  NAND2_X1 U35350 ( .A1(n3644), .A2(n3670), .ZN(n2774) );
  OR2_X1 U35360 ( .A1(n4075), .A2(n3681), .ZN(n3668) );
  INV_X1 U35370 ( .A(n3668), .ZN(n2773) );
  AOI21_X1 U35380 ( .B1(n2775), .B2(n2774), .A(n2773), .ZN(n4033) );
  INV_X1 U35390 ( .A(n4468), .ZN(n3659) );
  OR2_X1 U35400 ( .A1(n4479), .A2(n3659), .ZN(n3920) );
  NAND2_X1 U35410 ( .A1(n4479), .A2(n3659), .ZN(n3919) );
  NAND2_X1 U35420 ( .A1(n3920), .A2(n3919), .ZN(n3948) );
  INV_X1 U35430 ( .A(n3917), .ZN(n2776) );
  NOR2_X1 U35440 ( .A1(n3948), .A2(n2776), .ZN(n2777) );
  NAND2_X1 U35450 ( .A1(n3735), .A2(n2777), .ZN(n2778) );
  NAND2_X1 U35460 ( .A1(n2778), .A2(n3919), .ZN(n4374) );
  INV_X1 U35470 ( .A(n4373), .ZN(n2779) );
  NAND2_X1 U35480 ( .A1(n4374), .A2(n2779), .ZN(n2780) );
  INV_X1 U35490 ( .A(n3806), .ZN(n4315) );
  NAND2_X1 U35500 ( .A1(n4332), .A2(n4315), .ZN(n2781) );
  AND2_X1 U35510 ( .A1(n4305), .A2(n2781), .ZN(n2785) );
  OR2_X1 U35520 ( .A1(n4576), .A2(n4357), .ZN(n4302) );
  NAND2_X1 U35530 ( .A1(n4304), .A2(n4302), .ZN(n2783) );
  NOR2_X1 U35540 ( .A1(n4332), .A2(n4315), .ZN(n2782) );
  AOI21_X1 U35550 ( .B1(n2785), .B2(n2783), .A(n2782), .ZN(n4279) );
  OR2_X1 U35560 ( .A1(n4272), .A2(n4292), .ZN(n2784) );
  INV_X1 U35570 ( .A(n2785), .ZN(n4223) );
  AND2_X1 U35580 ( .A1(n4576), .A2(n4357), .ZN(n4222) );
  OR2_X1 U35590 ( .A1(n4223), .A2(n4222), .ZN(n4037) );
  AND2_X1 U35600 ( .A1(n4272), .A2(n4292), .ZN(n4224) );
  AOI21_X1 U35610 ( .B1(n4225), .B2(n4037), .A(n4224), .ZN(n3924) );
  OR2_X1 U35620 ( .A1(n4439), .A2(n4271), .ZN(n4226) );
  NAND2_X1 U35630 ( .A1(n4228), .A2(n4226), .ZN(n4043) );
  INV_X1 U35640 ( .A(n4043), .ZN(n2786) );
  NAND2_X1 U35650 ( .A1(n4412), .A2(n4236), .ZN(n2788) );
  NAND2_X1 U35660 ( .A1(n2788), .A2(n2787), .ZN(n4046) );
  AND2_X1 U35670 ( .A1(n4439), .A2(n4271), .ZN(n4041) );
  AND2_X1 U35680 ( .A1(n4228), .A2(n4041), .ZN(n2789) );
  NOR2_X1 U35690 ( .A1(n4046), .A2(n2789), .ZN(n3927) );
  NAND2_X1 U35700 ( .A1(n2790), .A2(n3927), .ZN(n4201) );
  NAND2_X1 U35710 ( .A1(n4193), .A2(n4410), .ZN(n3947) );
  OR2_X1 U35720 ( .A1(n4412), .A2(n4236), .ZN(n4200) );
  NAND2_X1 U35730 ( .A1(n4201), .A2(n4045), .ZN(n2791) );
  NAND2_X1 U35740 ( .A1(n4233), .A2(n4207), .ZN(n3946) );
  NAND2_X1 U35750 ( .A1(n2791), .A2(n3946), .ZN(n4189) );
  AND2_X1 U35760 ( .A1(n4211), .A2(n3827), .ZN(n3951) );
  NAND2_X1 U35770 ( .A1(n4157), .A2(n3892), .ZN(n3975) );
  OR2_X1 U35780 ( .A1(n4211), .A2(n3827), .ZN(n4166) );
  NAND2_X1 U35790 ( .A1(n4393), .A2(n4177), .ZN(n3974) );
  AND2_X1 U35800 ( .A1(n4074), .A2(n4154), .ZN(n4051) );
  INV_X1 U35810 ( .A(n4051), .ZN(n2792) );
  OR2_X1 U3582 ( .A1(n4074), .A2(n4154), .ZN(n2793) );
  INV_X1 U3583 ( .A(n2793), .ZN(n3934) );
  XNOR2_X1 U3584 ( .A(n3196), .B(n3953), .ZN(n2795) );
  INV_X1 U3585 ( .A(n2242), .ZN(n4562) );
  NAND2_X1 U3586 ( .A1(n4562), .A2(n2757), .ZN(n4063) );
  NAND2_X1 U3587 ( .A1(n4563), .A2(n4561), .ZN(n2794) );
  NAND2_X1 U3588 ( .A1(n2795), .A2(n4375), .ZN(n3778) );
  OAI211_X1 U3589 ( .C1(n3790), .C2(n4452), .A(n2796), .B(n3778), .ZN(n2916)
         );
  OR2_X1 U3590 ( .A1(n2798), .A2(n2797), .ZN(n2799) );
  MUX2_X1 U3591 ( .A(IR_REG_31__SCAN_IN), .B(n2799), .S(IR_REG_25__SCAN_IN), 
        .Z(n2800) );
  NAND2_X1 U3592 ( .A1(n2800), .A2(n2253), .ZN(n3222) );
  NAND2_X1 U3593 ( .A1(n3222), .A2(B_REG_SCAN_IN), .ZN(n2805) );
  NAND2_X1 U3594 ( .A1(n2801), .A2(IR_REG_31__SCAN_IN), .ZN(n2811) );
  NAND2_X1 U3595 ( .A1(n2811), .A2(n2810), .ZN(n2802) );
  NAND2_X1 U3596 ( .A1(n2802), .A2(IR_REG_31__SCAN_IN), .ZN(n2804) );
  XNOR2_X1 U3597 ( .A(n2804), .B(n2803), .ZN(n2825) );
  INV_X1 U3598 ( .A(n2825), .ZN(n4560) );
  MUX2_X1 U3599 ( .A(n2805), .B(B_REG_SCAN_IN), .S(n4560), .Z(n2806) );
  NAND2_X1 U3600 ( .A1(n2253), .A2(IR_REG_31__SCAN_IN), .ZN(n2807) );
  NOR2_X1 U3601 ( .A1(n3227), .A2(D_REG_1__SCAN_IN), .ZN(n3158) );
  AND2_X1 U3602 ( .A1(n2826), .A2(n3222), .ZN(n3228) );
  XNOR2_X1 U3603 ( .A(n2811), .B(n2810), .ZN(n2862) );
  NAND2_X1 U3604 ( .A1(n2242), .A2(n4123), .ZN(n3160) );
  NAND2_X1 U3605 ( .A1(n3160), .A2(n2863), .ZN(n3312) );
  OAI211_X1 U3606 ( .C1(n4733), .C2(n2757), .A(n3279), .B(n3312), .ZN(n2812)
         );
  INV_X1 U3607 ( .A(n2812), .ZN(n2824) );
  NOR4_X1 U3608 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n2816) );
  NOR4_X1 U3609 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_2__SCAN_IN), .A3(
        D_REG_29__SCAN_IN), .A4(D_REG_6__SCAN_IN), .ZN(n2815) );
  NOR4_X1 U3610 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2814) );
  NOR4_X1 U3611 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_20__SCAN_IN), .A3(
        D_REG_13__SCAN_IN), .A4(D_REG_16__SCAN_IN), .ZN(n2813) );
  NAND4_X1 U3612 ( .A1(n2816), .A2(n2815), .A3(n2814), .A4(n2813), .ZN(n2823)
         );
  NOR2_X1 U3613 ( .A1(D_REG_30__SCAN_IN), .A2(D_REG_25__SCAN_IN), .ZN(n2820)
         );
  NOR4_X1 U3614 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_23__SCAN_IN), .ZN(n2819) );
  NOR4_X1 U3615 ( .A1(D_REG_3__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_28__SCAN_IN), .ZN(n2818) );
  NOR4_X1 U3616 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_11__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2817) );
  NAND4_X1 U3617 ( .A1(n2820), .A2(n2819), .A3(n2818), .A4(n2817), .ZN(n2822)
         );
  OAI21_X1 U3618 ( .B1(n2823), .B2(n2822), .A(n2821), .ZN(n3157) );
  OAI211_X1 U3619 ( .C1(n3158), .C2(n3228), .A(n2824), .B(n3157), .ZN(n2915)
         );
  NAND2_X1 U3620 ( .A1(n2826), .A2(n2825), .ZN(n3229) );
  INV_X1 U3621 ( .A(n3311), .ZN(n2827) );
  AND2_X2 U3622 ( .A1(n3392), .A2(n3421), .ZN(n3446) );
  NAND2_X1 U3623 ( .A1(n3446), .A2(n3445), .ZN(n3444) );
  NOR2_X2 U3624 ( .A1(n3444), .A2(n3836), .ZN(n3466) );
  NAND2_X1 U3625 ( .A1(n3466), .A2(n3472), .ZN(n3486) );
  NOR2_X4 U3626 ( .A1(n3637), .A2(n3715), .ZN(n3682) );
  OAI21_X1 U3627 ( .B1(n4152), .B2(n3771), .A(n3206), .ZN(n3786) );
  INV_X1 U3628 ( .A(n3306), .ZN(n3161) );
  INV_X1 U3630 ( .A(REG0_REG_28__SCAN_IN), .ZN(n2829) );
  AOI22_X1 U3631 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4717), .B1(n4111), .B2(
        n4338), .ZN(n2868) );
  NOR2_X1 U3632 ( .A1(REG2_REG_17__SCAN_IN), .A2(n2901), .ZN(n2833) );
  AOI21_X1 U3633 ( .B1(REG2_REG_17__SCAN_IN), .B2(n2901), .A(n2833), .ZN(n4680) );
  INV_X1 U3634 ( .A(n4724), .ZN(n4651) );
  NOR2_X1 U3635 ( .A1(n3683), .A2(n4651), .ZN(n4639) );
  NAND2_X1 U3636 ( .A1(REG2_REG_11__SCAN_IN), .A2(n2872), .ZN(n2850) );
  AOI22_X1 U3637 ( .A1(REG2_REG_11__SCAN_IN), .A2(n2872), .B1(n4727), .B2(
        n2585), .ZN(n4623) );
  NAND2_X1 U3638 ( .A1(n2874), .A2(REG2_REG_9__SCAN_IN), .ZN(n2846) );
  INV_X1 U3639 ( .A(n2874), .ZN(n4729) );
  AOI22_X1 U3640 ( .A1(n2874), .A2(REG2_REG_9__SCAN_IN), .B1(n2562), .B2(n4729), .ZN(n4602) );
  INV_X1 U3641 ( .A(n3254), .ZN(n2883) );
  INV_X1 U3642 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2837) );
  INV_X1 U3643 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2834) );
  MUX2_X1 U3644 ( .A(REG2_REG_1__SCAN_IN), .B(n2834), .S(n4091), .Z(n2835) );
  NOR2_X1 U3645 ( .A1(n4091), .A2(n2834), .ZN(n3336) );
  NAND2_X1 U3646 ( .A1(n3333), .A2(REG2_REG_2__SCAN_IN), .ZN(n2836) );
  XNOR2_X1 U3647 ( .A(n2839), .B(n2838), .ZN(n4105) );
  AOI22_X1 U3648 ( .A1(n4105), .A2(REG2_REG_3__SCAN_IN), .B1(n4102), .B2(n2839), .ZN(n2840) );
  XNOR2_X1 U3649 ( .A(n2840), .B(n3349), .ZN(n3344) );
  MUX2_X1 U3650 ( .A(n2343), .B(REG2_REG_5__SCAN_IN), .S(n3218), .Z(n3238) );
  XNOR2_X1 U3651 ( .A(n2842), .B(n4565), .ZN(n3258) );
  INV_X1 U3652 ( .A(n2842), .ZN(n2843) );
  MUX2_X1 U3653 ( .A(REG2_REG_7__SCAN_IN), .B(n2540), .S(n3254), .Z(n3245) );
  INV_X1 U3654 ( .A(n4564), .ZN(n2886) );
  OAI22_X1 U3655 ( .A1(n3269), .A2(n2845), .B1(n2844), .B2(n2886), .ZN(n4601)
         );
  NAND2_X1 U3656 ( .A1(n4608), .A2(n2848), .ZN(n2849) );
  NAND2_X1 U3657 ( .A1(n2849), .A2(n4609), .ZN(n4622) );
  NAND2_X1 U3658 ( .A1(n4629), .A2(n2852), .ZN(n2853) );
  OAI22_X1 U3659 ( .A1(n4639), .A2(n4642), .B1(REG2_REG_13__SCAN_IN), .B2(
        n4724), .ZN(n2854) );
  NOR2_X1 U3660 ( .A1(n4723), .A2(n2854), .ZN(n2855) );
  NAND2_X1 U3661 ( .A1(REG2_REG_15__SCAN_IN), .A2(n2870), .ZN(n2856) );
  OAI21_X1 U3662 ( .B1(REG2_REG_15__SCAN_IN), .B2(n2870), .A(n2856), .ZN(n4661) );
  AND2_X1 U3663 ( .A1(n2870), .A2(REG2_REG_15__SCAN_IN), .ZN(n2857) );
  INV_X1 U3664 ( .A(n2859), .ZN(n2858) );
  NAND2_X1 U3665 ( .A1(n2858), .A2(n4720), .ZN(n2860) );
  NAND2_X1 U3666 ( .A1(n4670), .A2(n4370), .ZN(n4669) );
  OR2_X1 U3667 ( .A1(n2862), .A2(U3149), .ZN(n4070) );
  INV_X1 U3668 ( .A(n4070), .ZN(n2861) );
  OR2_X1 U3669 ( .A1(n3279), .A2(n2861), .ZN(n2906) );
  NAND2_X1 U3670 ( .A1(n2863), .A2(n2862), .ZN(n2864) );
  NAND2_X1 U3671 ( .A1(n2240), .A2(n2864), .ZN(n2905) );
  INV_X1 U3672 ( .A(n2905), .ZN(n2865) );
  XNOR2_X1 U3673 ( .A(n2866), .B(IR_REG_27__SCAN_IN), .ZN(n4591) );
  INV_X1 U3674 ( .A(n4591), .ZN(n2902) );
  NOR2_X1 U3675 ( .A1(n4570), .A2(n2902), .ZN(n4066) );
  AOI211_X1 U3676 ( .C1(n2868), .C2(n2867), .A(n4113), .B(n4677), .ZN(n2914)
         );
  INV_X1 U3677 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4117) );
  AOI22_X1 U3678 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4111), .B1(n4717), .B2(
        n4117), .ZN(n2904) );
  NAND2_X1 U3679 ( .A1(REG1_REG_15__SCAN_IN), .A2(n2870), .ZN(n2897) );
  INV_X1 U3680 ( .A(n2870), .ZN(n4721) );
  INV_X1 U3681 ( .A(REG1_REG_15__SCAN_IN), .ZN(n2869) );
  AOI22_X1 U3682 ( .A1(REG1_REG_15__SCAN_IN), .A2(n2870), .B1(n4721), .B2(
        n2869), .ZN(n4666) );
  NAND2_X1 U3683 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4724), .ZN(n2893) );
  INV_X1 U3684 ( .A(REG1_REG_13__SCAN_IN), .ZN(n2871) );
  AOI22_X1 U3685 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4724), .B1(n4651), .B2(
        n2871), .ZN(n4648) );
  INV_X1 U3686 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4768) );
  AOI22_X1 U3687 ( .A1(REG1_REG_11__SCAN_IN), .A2(n2872), .B1(n4727), .B2(
        n4768), .ZN(n4620) );
  NAND2_X1 U3688 ( .A1(n2874), .A2(REG1_REG_9__SCAN_IN), .ZN(n2888) );
  INV_X1 U3689 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2873) );
  AOI22_X1 U3690 ( .A1(n2874), .A2(REG1_REG_9__SCAN_IN), .B1(n2873), .B2(n4729), .ZN(n4599) );
  XNOR2_X1 U3691 ( .A(n4091), .B(REG1_REG_1__SCAN_IN), .ZN(n4089) );
  AND2_X1 U3692 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n4088)
         );
  NAND2_X1 U3693 ( .A1(n4089), .A2(n4088), .ZN(n4087) );
  INV_X1 U3694 ( .A(n4091), .ZN(n4568) );
  NAND2_X1 U3695 ( .A1(n4568), .A2(REG1_REG_1__SCAN_IN), .ZN(n2875) );
  NAND2_X1 U3696 ( .A1(n4087), .A2(n2875), .ZN(n3334) );
  XNOR2_X1 U3697 ( .A(n3333), .B(REG1_REG_2__SCAN_IN), .ZN(n3335) );
  INV_X1 U3698 ( .A(n3333), .ZN(n4567) );
  NAND2_X1 U3699 ( .A1(n4567), .A2(REG1_REG_2__SCAN_IN), .ZN(n2876) );
  XNOR2_X1 U3700 ( .A(n2877), .B(n2838), .ZN(n4101) );
  NAND2_X1 U3701 ( .A1(n4101), .A2(REG1_REG_3__SCAN_IN), .ZN(n4100) );
  NAND2_X1 U3702 ( .A1(n2877), .A2(n4102), .ZN(n2878) );
  NAND2_X1 U3703 ( .A1(n4100), .A2(n2878), .ZN(n2879) );
  XNOR2_X1 U3704 ( .A(n2879), .B(n3349), .ZN(n3346) );
  INV_X1 U3705 ( .A(n3349), .ZN(n4566) );
  XNOR2_X1 U3706 ( .A(n3218), .B(REG1_REG_5__SCAN_IN), .ZN(n3235) );
  NOR2_X1 U3707 ( .A1(n3236), .A2(n3235), .ZN(n3234) );
  INV_X1 U3708 ( .A(n2881), .ZN(n2882) );
  INV_X1 U3709 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3262) );
  NAND2_X1 U3710 ( .A1(n2883), .A2(REG1_REG_7__SCAN_IN), .ZN(n3248) );
  NOR2_X1 U3711 ( .A1(n2883), .A2(REG1_REG_7__SCAN_IN), .ZN(n3247) );
  XNOR2_X1 U3712 ( .A(n2884), .B(n4564), .ZN(n3268) );
  INV_X1 U3713 ( .A(REG1_REG_8__SCAN_IN), .ZN(n2887) );
  INV_X1 U3714 ( .A(n2884), .ZN(n2885) );
  NAND2_X1 U3715 ( .A1(n4608), .A2(n2889), .ZN(n2890) );
  NAND2_X1 U3716 ( .A1(n2890), .A2(n4614), .ZN(n4619) );
  NAND2_X1 U3717 ( .A1(n4620), .A2(n4619), .ZN(n4618) );
  OAI21_X1 U3718 ( .B1(n4727), .B2(n4768), .A(n4618), .ZN(n2891) );
  NAND2_X1 U3719 ( .A1(n4629), .A2(n2891), .ZN(n2892) );
  NAND2_X1 U3720 ( .A1(n2894), .A2(n2895), .ZN(n2896) );
  NAND2_X1 U3721 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4657), .ZN(n4656) );
  NAND2_X1 U3722 ( .A1(n2896), .A2(n4656), .ZN(n4665) );
  NAND2_X1 U3723 ( .A1(n4666), .A2(n4665), .ZN(n4664) );
  NAND2_X1 U3724 ( .A1(n2897), .A2(n4664), .ZN(n2899) );
  XNOR2_X1 U3725 ( .A(n2899), .B(n2898), .ZN(n4673) );
  INV_X1 U3726 ( .A(REG1_REG_17__SCAN_IN), .ZN(n2900) );
  AOI22_X1 U3727 ( .A1(n4718), .A2(REG1_REG_17__SCAN_IN), .B1(n2900), .B2(
        n2901), .ZN(n4685) );
  NAND2_X1 U3728 ( .A1(n2903), .A2(n2904), .ZN(n4116) );
  OAI211_X1 U3729 ( .C1(n2904), .C2(n2903), .A(n4684), .B(n4116), .ZN(n2912)
         );
  NAND2_X1 U3730 ( .A1(n4593), .A2(n4570), .ZN(n4689) );
  INV_X1 U3731 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2907) );
  NOR2_X1 U3732 ( .A1(STATE_REG_SCAN_IN), .A2(n2907), .ZN(n2908) );
  AOI21_X1 U3733 ( .B1(n4683), .B2(ADDR_REG_18__SCAN_IN), .A(n2908), .ZN(n2909) );
  OAI21_X1 U3734 ( .B1(n4689), .B2(n4717), .A(n2909), .ZN(n2910) );
  INV_X1 U3735 ( .A(n2910), .ZN(n2911) );
  OR2_X1 U3736 ( .A1(n2914), .A2(n2913), .ZN(U3258) );
  NAND2_X1 U3737 ( .A1(n2916), .A2(n4770), .ZN(n2920) );
  INV_X1 U3738 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2917) );
  NAND2_X1 U3739 ( .A1(n2920), .A2(n2919), .ZN(U3546) );
  NAND2_X1 U3740 ( .A1(n2925), .A2(n2958), .ZN(n2924) );
  INV_X1 U3741 ( .A(n2922), .ZN(n2923) );
  NAND2_X1 U3742 ( .A1(n2924), .A2(n2923), .ZN(n3291) );
  NAND2_X1 U3743 ( .A1(n2925), .A2(n3143), .ZN(n2927) );
  NAND2_X1 U3744 ( .A1(n3367), .A2(n3069), .ZN(n2926) );
  NAND2_X1 U3745 ( .A1(n2927), .A2(n2926), .ZN(n2932) );
  INV_X1 U3746 ( .A(n2932), .ZN(n2929) );
  INV_X1 U3747 ( .A(REG1_REG_0__SCAN_IN), .ZN(n2928) );
  NAND2_X1 U3748 ( .A1(n2929), .A2(n2434), .ZN(n3292) );
  NAND2_X1 U3749 ( .A1(n3291), .A2(n3292), .ZN(n3290) );
  NOR2_X1 U3750 ( .A1(n4563), .A2(n2930), .ZN(n3170) );
  INV_X1 U3751 ( .A(n3170), .ZN(n2931) );
  NAND2_X4 U3752 ( .A1(n2921), .A2(n2931), .ZN(n3766) );
  OR2_X1 U3753 ( .A1(n2932), .A2(n3766), .ZN(n2933) );
  NAND2_X1 U3754 ( .A1(n3290), .A2(n2933), .ZN(n3282) );
  NAND2_X1 U3755 ( .A1(n2934), .A2(n3143), .ZN(n2937) );
  INV_X1 U3756 ( .A(n3359), .ZN(n2935) );
  NAND2_X1 U3757 ( .A1(n2935), .A2(n3069), .ZN(n2936) );
  NAND2_X1 U3758 ( .A1(n2937), .A2(n2936), .ZN(n2938) );
  NOR2_X1 U3759 ( .A1(n3359), .A2(n2939), .ZN(n2940) );
  AOI21_X1 U3760 ( .B1(n2934), .B2(n2958), .A(n2940), .ZN(n2941) );
  XNOR2_X1 U3761 ( .A(n2943), .B(n2941), .ZN(n3283) );
  NAND2_X1 U3762 ( .A1(n3282), .A2(n3283), .ZN(n3281) );
  INV_X1 U3763 ( .A(n2941), .ZN(n2942) );
  NAND2_X1 U3764 ( .A1(n2943), .A2(n2942), .ZN(n2944) );
  NAND2_X1 U3765 ( .A1(n3281), .A2(n2944), .ZN(n3296) );
  INV_X1 U3766 ( .A(n3296), .ZN(n2951) );
  NAND2_X1 U3767 ( .A1(n3389), .A2(n2244), .ZN(n2945) );
  NAND2_X1 U3768 ( .A1(n2946), .A2(n2945), .ZN(n2947) );
  NOR2_X1 U3769 ( .A1(n3301), .A2(n3763), .ZN(n2948) );
  AOI21_X1 U3770 ( .B1(n2949), .B2(n2958), .A(n2948), .ZN(n2952) );
  XNOR2_X1 U3771 ( .A(n2953), .B(n2952), .ZN(n3295) );
  INV_X1 U3772 ( .A(n3295), .ZN(n2950) );
  NAND2_X1 U3773 ( .A1(n2951), .A2(n2950), .ZN(n3297) );
  NAND2_X1 U3774 ( .A1(n2953), .A2(n2952), .ZN(n2954) );
  NAND2_X1 U3775 ( .A1(n3297), .A2(n2954), .ZN(n3321) );
  NAND2_X1 U3776 ( .A1(n4085), .A2(n2235), .ZN(n2956) );
  NAND2_X1 U3777 ( .A1(n3374), .A2(n2244), .ZN(n2955) );
  NAND2_X1 U3778 ( .A1(n2956), .A2(n2955), .ZN(n2957) );
  XNOR2_X1 U3779 ( .A(n2957), .B(n3766), .ZN(n2960) );
  NOR2_X1 U3780 ( .A1(n3421), .A2(n3763), .ZN(n2959) );
  AOI21_X1 U3781 ( .B1(n4085), .B2(n3764), .A(n2959), .ZN(n2961) );
  XNOR2_X1 U3782 ( .A(n2960), .B(n2961), .ZN(n3322) );
  NAND2_X1 U3783 ( .A1(n3321), .A2(n3322), .ZN(n2964) );
  INV_X1 U3784 ( .A(n2960), .ZN(n2962) );
  NAND2_X1 U3785 ( .A1(n2962), .A2(n2961), .ZN(n2963) );
  NAND2_X1 U3786 ( .A1(n2964), .A2(n2963), .ZN(n3410) );
  INV_X1 U3787 ( .A(n3410), .ZN(n2970) );
  NAND2_X1 U3788 ( .A1(n4084), .A2(n2235), .ZN(n2966) );
  NAND2_X1 U3789 ( .A1(n3438), .A2(n2244), .ZN(n2965) );
  NOR2_X1 U3790 ( .A1(n3445), .A2(n3763), .ZN(n2968) );
  AOI21_X1 U3791 ( .B1(n4084), .B2(n3764), .A(n2968), .ZN(n2972) );
  XNOR2_X1 U3792 ( .A(n2971), .B(n2972), .ZN(n3413) );
  INV_X1 U3793 ( .A(n3413), .ZN(n2969) );
  NAND2_X1 U3794 ( .A1(n2970), .A2(n2969), .ZN(n3411) );
  INV_X1 U3795 ( .A(n2971), .ZN(n2974) );
  INV_X1 U3796 ( .A(n2972), .ZN(n2973) );
  NAND2_X1 U3797 ( .A1(n2974), .A2(n2973), .ZN(n2975) );
  NAND2_X1 U3798 ( .A1(n3411), .A2(n2975), .ZN(n3834) );
  NAND2_X1 U3799 ( .A1(n4083), .A2(n2236), .ZN(n2977) );
  NAND2_X1 U3800 ( .A1(n3836), .A2(n2244), .ZN(n2976) );
  NAND2_X1 U3801 ( .A1(n2977), .A2(n2976), .ZN(n2978) );
  XNOR2_X1 U3802 ( .A(n2978), .B(n3766), .ZN(n2982) );
  NOR2_X1 U3803 ( .A1(n3478), .A2(n3763), .ZN(n2979) );
  AOI21_X1 U3804 ( .B1(n4083), .B2(n3764), .A(n2979), .ZN(n2980) );
  XNOR2_X1 U3805 ( .A(n2982), .B(n2980), .ZN(n3833) );
  INV_X1 U3806 ( .A(n2980), .ZN(n2981) );
  NAND2_X1 U3807 ( .A1(n2982), .A2(n2981), .ZN(n2983) );
  NAND2_X1 U3808 ( .A1(n4082), .A2(n3764), .ZN(n2985) );
  NAND2_X1 U3809 ( .A1(n3497), .A2(n2236), .ZN(n2984) );
  NAND2_X1 U3810 ( .A1(n2985), .A2(n2984), .ZN(n3452) );
  NAND2_X1 U3811 ( .A1(n4082), .A2(n2236), .ZN(n2987) );
  NAND2_X1 U3812 ( .A1(n3497), .A2(n2244), .ZN(n2986) );
  NAND2_X1 U3813 ( .A1(n2987), .A2(n2986), .ZN(n2988) );
  XNOR2_X1 U3814 ( .A(n2988), .B(n3766), .ZN(n3453) );
  NAND2_X1 U3815 ( .A1(n4081), .A2(n2236), .ZN(n2990) );
  NAND2_X1 U3816 ( .A1(n3516), .A2(n2244), .ZN(n2989) );
  NAND2_X1 U3817 ( .A1(n2990), .A2(n2989), .ZN(n2991) );
  XNOR2_X1 U3818 ( .A(n2991), .B(n3766), .ZN(n3006) );
  NOR2_X1 U3819 ( .A1(n2992), .A2(n3763), .ZN(n2993) );
  AOI21_X1 U3820 ( .B1(n4081), .B2(n3764), .A(n2993), .ZN(n3004) );
  XNOR2_X1 U3821 ( .A(n3006), .B(n3004), .ZN(n3523) );
  NAND2_X1 U3822 ( .A1(n4080), .A2(n2236), .ZN(n2995) );
  NAND2_X1 U3823 ( .A1(n3579), .A2(n2244), .ZN(n2994) );
  NAND2_X1 U3824 ( .A1(n2995), .A2(n2994), .ZN(n2996) );
  XNOR2_X1 U3825 ( .A(n2996), .B(n3766), .ZN(n3003) );
  INV_X1 U3826 ( .A(n3003), .ZN(n3000) );
  NAND2_X1 U3827 ( .A1(n4080), .A2(n3764), .ZN(n2998) );
  NAND2_X1 U3828 ( .A1(n3579), .A2(n2236), .ZN(n2997) );
  NAND2_X1 U3829 ( .A1(n2998), .A2(n2997), .ZN(n3002) );
  INV_X1 U3830 ( .A(n3002), .ZN(n2999) );
  NAND2_X1 U3831 ( .A1(n3000), .A2(n2999), .ZN(n3526) );
  AND2_X1 U3832 ( .A1(n3523), .A2(n3526), .ZN(n3001) );
  NAND2_X1 U3833 ( .A1(n3514), .A2(n3001), .ZN(n3552) );
  INV_X1 U3834 ( .A(n3526), .ZN(n3008) );
  INV_X1 U3835 ( .A(n3004), .ZN(n3005) );
  NAND2_X1 U3836 ( .A1(n3006), .A2(n3005), .ZN(n3524) );
  AND2_X1 U3837 ( .A1(n2255), .A2(n3524), .ZN(n3007) );
  OR2_X1 U3838 ( .A1(n3008), .A2(n3007), .ZN(n3551) );
  NAND2_X1 U3839 ( .A1(n4079), .A2(n2236), .ZN(n3010) );
  NAND2_X1 U3840 ( .A1(n3555), .A2(n2244), .ZN(n3009) );
  NAND2_X1 U3841 ( .A1(n3010), .A2(n3009), .ZN(n3011) );
  XNOR2_X1 U3842 ( .A(n3011), .B(n3766), .ZN(n3014) );
  NOR2_X1 U3843 ( .A1(n3598), .A2(n3763), .ZN(n3012) );
  AOI21_X1 U3844 ( .B1(n4079), .B2(n3764), .A(n3012), .ZN(n3015) );
  XNOR2_X1 U3845 ( .A(n3014), .B(n3015), .ZN(n3553) );
  AND2_X1 U3846 ( .A1(n3551), .A2(n3553), .ZN(n3013) );
  NAND2_X1 U3847 ( .A1(n3552), .A2(n3013), .ZN(n3018) );
  INV_X1 U3848 ( .A(n3014), .ZN(n3016) );
  NAND2_X1 U3849 ( .A1(n3016), .A2(n3015), .ZN(n3017) );
  NAND2_X1 U3850 ( .A1(n3018), .A2(n3017), .ZN(n3562) );
  INV_X1 U3851 ( .A(n3562), .ZN(n3024) );
  NAND2_X1 U3852 ( .A1(n4078), .A2(n2236), .ZN(n3020) );
  NAND2_X1 U3853 ( .A1(n3692), .A2(n2244), .ZN(n3019) );
  NAND2_X1 U3854 ( .A1(n3020), .A2(n3019), .ZN(n3021) );
  XNOR2_X1 U3855 ( .A(n3021), .B(n3152), .ZN(n3025) );
  NOR2_X1 U3856 ( .A1(n3689), .A2(n3763), .ZN(n3022) );
  AOI21_X1 U3857 ( .B1(n4078), .B2(n3764), .A(n3022), .ZN(n3026) );
  XNOR2_X1 U3858 ( .A(n3025), .B(n3026), .ZN(n3565) );
  INV_X1 U3859 ( .A(n3025), .ZN(n3028) );
  INV_X1 U3860 ( .A(n3026), .ZN(n3027) );
  NAND2_X1 U3861 ( .A1(n3028), .A2(n3027), .ZN(n3029) );
  NAND2_X1 U3862 ( .A1(n4077), .A2(n3764), .ZN(n3031) );
  NAND2_X1 U3863 ( .A1(n3592), .A2(n2236), .ZN(n3030) );
  NAND2_X1 U3864 ( .A1(n3031), .A2(n3030), .ZN(n3589) );
  NAND2_X1 U3865 ( .A1(n4077), .A2(n2236), .ZN(n3033) );
  NAND2_X1 U3866 ( .A1(n3592), .A2(n2244), .ZN(n3032) );
  NAND2_X1 U3867 ( .A1(n3033), .A2(n3032), .ZN(n3034) );
  XNOR2_X1 U3868 ( .A(n3034), .B(n3766), .ZN(n3590) );
  NAND2_X1 U3869 ( .A1(n4076), .A2(n2236), .ZN(n3036) );
  NAND2_X1 U3870 ( .A1(n3715), .A2(n2244), .ZN(n3035) );
  NAND2_X1 U3871 ( .A1(n3036), .A2(n3035), .ZN(n3037) );
  XNOR2_X1 U3872 ( .A(n3037), .B(n3766), .ZN(n3040) );
  NAND2_X1 U3873 ( .A1(n4076), .A2(n3764), .ZN(n3039) );
  NAND2_X1 U3874 ( .A1(n3715), .A2(n2236), .ZN(n3038) );
  NAND2_X1 U3875 ( .A1(n3039), .A2(n3038), .ZN(n3041) );
  INV_X1 U3876 ( .A(n3040), .ZN(n3043) );
  INV_X1 U3877 ( .A(n3041), .ZN(n3042) );
  NAND2_X1 U3878 ( .A1(n3043), .A2(n3042), .ZN(n3627) );
  NAND2_X1 U3879 ( .A1(n4075), .A2(n2236), .ZN(n3045) );
  NAND2_X1 U3880 ( .A1(n3708), .A2(n2244), .ZN(n3044) );
  NAND2_X1 U3881 ( .A1(n3045), .A2(n3044), .ZN(n3046) );
  NAND2_X1 U3882 ( .A1(n3704), .A2(n3705), .ZN(n3049) );
  NOR2_X1 U3883 ( .A1(n3681), .A2(n3763), .ZN(n3047) );
  AOI21_X1 U3884 ( .B1(n4075), .B2(n3764), .A(n3047), .ZN(n3706) );
  NAND2_X1 U3885 ( .A1(n3049), .A2(n3048), .ZN(n3053) );
  INV_X1 U3886 ( .A(n3704), .ZN(n3051) );
  INV_X1 U3887 ( .A(n3705), .ZN(n3050) );
  NAND2_X1 U3888 ( .A1(n3051), .A2(n3050), .ZN(n3052) );
  NAND2_X1 U3889 ( .A1(n3053), .A2(n3052), .ZN(n3750) );
  INV_X1 U3890 ( .A(n3750), .ZN(n3064) );
  NAND2_X1 U3891 ( .A1(n4467), .A2(n2236), .ZN(n3055) );
  NAND2_X1 U3892 ( .A1(n4476), .A2(n2244), .ZN(n3054) );
  NAND2_X1 U3893 ( .A1(n3055), .A2(n3054), .ZN(n3056) );
  XNOR2_X1 U3894 ( .A(n3056), .B(n3766), .ZN(n3059) );
  NAND2_X1 U3895 ( .A1(n4467), .A2(n3764), .ZN(n3058) );
  NAND2_X1 U3896 ( .A1(n4476), .A2(n2236), .ZN(n3057) );
  NAND2_X1 U3897 ( .A1(n3058), .A2(n3057), .ZN(n3060) );
  INV_X1 U3898 ( .A(n3059), .ZN(n3062) );
  INV_X1 U3899 ( .A(n3060), .ZN(n3061) );
  NAND2_X1 U3900 ( .A1(n3062), .A2(n3061), .ZN(n3751) );
  NAND2_X1 U3901 ( .A1(n4479), .A2(n2236), .ZN(n3066) );
  NAND2_X1 U3902 ( .A1(n4468), .A2(n2244), .ZN(n3065) );
  NAND2_X1 U3903 ( .A1(n3066), .A2(n3065), .ZN(n3067) );
  XNOR2_X1 U3904 ( .A(n3067), .B(n3766), .ZN(n3077) );
  NOR2_X1 U3905 ( .A1(n3659), .A2(n3763), .ZN(n3068) );
  NAND2_X1 U3906 ( .A1(n4469), .A2(n2236), .ZN(n3071) );
  NAND2_X1 U3907 ( .A1(n4377), .A2(n2244), .ZN(n3070) );
  NAND2_X1 U3908 ( .A1(n3071), .A2(n3070), .ZN(n3072) );
  XNOR2_X1 U3909 ( .A(n3072), .B(n3766), .ZN(n3076) );
  NAND2_X1 U3910 ( .A1(n4469), .A2(n3764), .ZN(n3074) );
  NAND2_X1 U3911 ( .A1(n4377), .A2(n2236), .ZN(n3073) );
  NAND2_X1 U3912 ( .A1(n3074), .A2(n3073), .ZN(n3075) );
  NOR2_X1 U3913 ( .A1(n3076), .A2(n3075), .ZN(n3079) );
  AOI21_X1 U3914 ( .B1(n3076), .B2(n3075), .A(n3079), .ZN(n4580) );
  NAND2_X1 U3915 ( .A1(n3078), .A2(n3077), .ZN(n3901) );
  INV_X1 U3916 ( .A(n3079), .ZN(n3080) );
  NAND2_X1 U3917 ( .A1(n4576), .A2(n2236), .ZN(n3083) );
  NAND2_X1 U3918 ( .A1(n4454), .A2(n2244), .ZN(n3082) );
  NAND2_X1 U3919 ( .A1(n3083), .A2(n3082), .ZN(n3084) );
  XNOR2_X1 U3920 ( .A(n3084), .B(n3766), .ZN(n3088) );
  NAND2_X1 U3921 ( .A1(n4576), .A2(n3764), .ZN(n3086) );
  NAND2_X1 U3922 ( .A1(n4454), .A2(n2236), .ZN(n3085) );
  NAND2_X1 U3923 ( .A1(n3086), .A2(n3085), .ZN(n3087) );
  NAND2_X1 U3924 ( .A1(n3088), .A2(n3087), .ZN(n3843) );
  NOR2_X1 U3925 ( .A1(n3088), .A2(n3087), .ZN(n3844) );
  NAND2_X1 U3926 ( .A1(n4455), .A2(n2236), .ZN(n3090) );
  NAND2_X1 U3927 ( .A1(n4331), .A2(n2244), .ZN(n3089) );
  NAND2_X1 U3928 ( .A1(n3090), .A2(n3089), .ZN(n3091) );
  XNOR2_X1 U3929 ( .A(n3091), .B(n3152), .ZN(n3094) );
  NOR2_X1 U3930 ( .A1(n4328), .A2(n3763), .ZN(n3092) );
  AOI21_X1 U3931 ( .B1(n4455), .B2(n3764), .A(n3092), .ZN(n3093) );
  NOR2_X1 U3932 ( .A1(n3094), .A2(n3093), .ZN(n3881) );
  AOI22_X1 U3933 ( .A1(n4332), .A2(n3764), .B1(n2236), .B2(n3806), .ZN(n3098)
         );
  NAND2_X1 U3934 ( .A1(n4332), .A2(n2236), .ZN(n3096) );
  NAND2_X1 U3935 ( .A1(n3806), .A2(n2244), .ZN(n3095) );
  NAND2_X1 U3936 ( .A1(n3096), .A2(n3095), .ZN(n3097) );
  XNOR2_X1 U3937 ( .A(n3097), .B(n3766), .ZN(n3099) );
  XOR2_X1 U3938 ( .A(n3098), .B(n3099), .Z(n3805) );
  NAND2_X1 U3939 ( .A1(n4272), .A2(n2236), .ZN(n3101) );
  NAND2_X1 U3940 ( .A1(n4438), .A2(n2244), .ZN(n3100) );
  NAND2_X1 U3941 ( .A1(n3101), .A2(n3100), .ZN(n3102) );
  XNOR2_X1 U3942 ( .A(n3102), .B(n3766), .ZN(n3109) );
  NAND2_X1 U3943 ( .A1(n4272), .A2(n3764), .ZN(n3104) );
  NAND2_X1 U3944 ( .A1(n2236), .A2(n4438), .ZN(n3103) );
  NAND2_X1 U3945 ( .A1(n3104), .A2(n3103), .ZN(n3110) );
  NAND2_X1 U3946 ( .A1(n3109), .A2(n3110), .ZN(n3863) );
  NAND2_X1 U3947 ( .A1(n3812), .A2(n3863), .ZN(n3114) );
  NOR2_X1 U3948 ( .A1(n3763), .A2(n4271), .ZN(n3105) );
  AOI21_X1 U3949 ( .B1(n4439), .B2(n3764), .A(n3105), .ZN(n3813) );
  NAND2_X1 U3950 ( .A1(n4439), .A2(n2236), .ZN(n3107) );
  NAND2_X1 U3951 ( .A1(n4429), .A2(n2244), .ZN(n3106) );
  NAND2_X1 U3952 ( .A1(n3107), .A2(n3106), .ZN(n3108) );
  XNOR2_X1 U3953 ( .A(n3108), .B(n3152), .ZN(n3814) );
  INV_X1 U3954 ( .A(n3109), .ZN(n3112) );
  INV_X1 U3955 ( .A(n3110), .ZN(n3111) );
  AOI21_X1 U3956 ( .B1(n3813), .B2(n3814), .A(n3864), .ZN(n3113) );
  OAI22_X1 U3957 ( .A1(n4273), .A2(n3765), .B1(n3763), .B2(n4256), .ZN(n3121)
         );
  OAI22_X1 U3958 ( .A1(n4273), .A2(n3763), .B1(n2252), .B2(n4256), .ZN(n3115)
         );
  XNOR2_X1 U3959 ( .A(n3115), .B(n3766), .ZN(n3120) );
  XOR2_X1 U3960 ( .A(n3121), .B(n3120), .Z(n3873) );
  NAND2_X1 U3961 ( .A1(n4412), .A2(n2236), .ZN(n3117) );
  INV_X1 U3962 ( .A(n4236), .ZN(n3945) );
  NAND2_X1 U3963 ( .A1(n3945), .A2(n2244), .ZN(n3116) );
  NAND2_X1 U3964 ( .A1(n3117), .A2(n3116), .ZN(n3118) );
  XNOR2_X1 U3965 ( .A(n3118), .B(n3766), .ZN(n3125) );
  NOR2_X1 U3966 ( .A1(n3763), .A2(n4236), .ZN(n3119) );
  AOI21_X1 U3967 ( .B1(n4412), .B2(n3764), .A(n3119), .ZN(n3126) );
  XNOR2_X1 U3968 ( .A(n3125), .B(n3126), .ZN(n3797) );
  INV_X1 U3969 ( .A(n3120), .ZN(n3123) );
  INV_X1 U3970 ( .A(n3121), .ZN(n3122) );
  NAND2_X1 U3971 ( .A1(n3123), .A2(n3122), .ZN(n3798) );
  INV_X1 U3972 ( .A(n3125), .ZN(n3127) );
  OR2_X1 U3973 ( .A1(n3127), .A2(n3126), .ZN(n3131) );
  NAND2_X1 U3974 ( .A1(n3795), .A2(n3131), .ZN(n3130) );
  NOR2_X1 U3975 ( .A1(n3763), .A2(n4207), .ZN(n3128) );
  AOI21_X1 U3976 ( .B1(n4233), .B2(n3764), .A(n3128), .ZN(n3132) );
  NAND2_X1 U3977 ( .A1(n3130), .A2(n3129), .ZN(n3852) );
  INV_X1 U3978 ( .A(n3131), .ZN(n3133) );
  OAI22_X1 U3979 ( .A1(n4193), .A2(n2939), .B1(n2252), .B2(n4207), .ZN(n3134)
         );
  XNOR2_X1 U3980 ( .A(n3134), .B(n3766), .ZN(n3855) );
  NAND2_X1 U3981 ( .A1(n3851), .A2(n3855), .ZN(n3135) );
  NAND2_X1 U3982 ( .A1(n4211), .A2(n2236), .ZN(n3137) );
  NAND2_X1 U3983 ( .A1(n4190), .A2(n2244), .ZN(n3136) );
  NAND2_X1 U3984 ( .A1(n3137), .A2(n3136), .ZN(n3138) );
  XNOR2_X1 U3985 ( .A(n3138), .B(n3766), .ZN(n3142) );
  NAND2_X1 U3986 ( .A1(n4211), .A2(n3764), .ZN(n3140) );
  NAND2_X1 U3987 ( .A1(n2236), .A2(n4190), .ZN(n3139) );
  NAND2_X1 U3988 ( .A1(n3140), .A2(n3139), .ZN(n3141) );
  NOR2_X1 U3989 ( .A1(n3142), .A2(n3141), .ZN(n3823) );
  NAND2_X1 U3990 ( .A1(n3142), .A2(n3141), .ZN(n3824) );
  NAND2_X1 U3991 ( .A1(n4393), .A2(n2236), .ZN(n3145) );
  NAND2_X1 U3992 ( .A1(n3892), .A2(n2244), .ZN(n3144) );
  NAND2_X1 U3993 ( .A1(n3145), .A2(n3144), .ZN(n3146) );
  XNOR2_X1 U3994 ( .A(n3146), .B(n3152), .ZN(n3149) );
  NOR2_X1 U3995 ( .A1(n3763), .A2(n4177), .ZN(n3147) );
  AOI21_X1 U3996 ( .B1(n4393), .B2(n3764), .A(n3147), .ZN(n3148) );
  NAND2_X1 U3997 ( .A1(n3149), .A2(n3148), .ZN(n3889) );
  NAND2_X1 U3998 ( .A1(n4074), .A2(n2236), .ZN(n3151) );
  NAND2_X1 U3999 ( .A1(n4392), .A2(n2244), .ZN(n3150) );
  NAND2_X1 U4000 ( .A1(n3151), .A2(n3150), .ZN(n3153) );
  XNOR2_X1 U4001 ( .A(n3153), .B(n3152), .ZN(n3760) );
  NOR2_X1 U4002 ( .A1(n2939), .A2(n4154), .ZN(n3154) );
  AOI21_X1 U4003 ( .B1(n4074), .B2(n3764), .A(n3154), .ZN(n3759) );
  XNOR2_X1 U4004 ( .A(n3760), .B(n3759), .ZN(n3761) );
  XNOR2_X1 U4005 ( .A(n3762), .B(n3155), .ZN(n3166) );
  INV_X1 U4006 ( .A(n3228), .ZN(n3156) );
  AND2_X1 U4007 ( .A1(n3157), .A2(n3156), .ZN(n3313) );
  NOR2_X1 U4008 ( .A1(n3311), .A2(n3158), .ZN(n3159) );
  NAND2_X1 U4009 ( .A1(n3313), .A2(n3159), .ZN(n3182) );
  INV_X1 U4010 ( .A(n3182), .ZN(n3165) );
  INV_X1 U4011 ( .A(n3279), .ZN(n3310) );
  NAND2_X1 U4012 ( .A1(n3161), .A2(n3160), .ZN(n3163) );
  NAND2_X1 U4013 ( .A1(n3163), .A2(n3162), .ZN(n3178) );
  NOR2_X1 U4014 ( .A1(n3310), .A2(n3178), .ZN(n3164) );
  NAND2_X1 U4015 ( .A1(n3165), .A2(n3164), .ZN(n3861) );
  NAND2_X1 U4016 ( .A1(n3166), .A2(n4581), .ZN(n3190) );
  NAND2_X1 U4017 ( .A1(n4477), .A2(n3279), .ZN(n3167) );
  OR2_X1 U4018 ( .A1(n3182), .A2(n3167), .ZN(n3169) );
  NAND2_X1 U4019 ( .A1(n3279), .A2(n3990), .ZN(n3168) );
  NAND2_X1 U4020 ( .A1(n3169), .A2(n4369), .ZN(n3904) );
  NAND2_X1 U4021 ( .A1(n3170), .A2(n4716), .ZN(n3171) );
  NOR2_X1 U4022 ( .A1(n3763), .A2(n3171), .ZN(n4067) );
  INV_X1 U4023 ( .A(n4570), .ZN(n3172) );
  NAND2_X1 U4024 ( .A1(n4067), .A2(n3172), .ZN(n3173) );
  OAI22_X1 U4025 ( .A1(n4157), .A2(n4571), .B1(STATE_REG_SCAN_IN), .B2(n3174), 
        .ZN(n3177) );
  NAND2_X1 U4026 ( .A1(n4067), .A2(n4570), .ZN(n3175) );
  NOR2_X1 U4027 ( .A1(n4396), .A2(n3875), .ZN(n3176) );
  AOI211_X1 U4028 ( .C1(n4392), .C2(n3904), .A(n3177), .B(n3176), .ZN(n3188)
         );
  INV_X1 U4029 ( .A(n4156), .ZN(n3186) );
  NAND2_X1 U4030 ( .A1(n3178), .A2(n4309), .ZN(n3179) );
  NAND2_X1 U4031 ( .A1(n3182), .A2(n3179), .ZN(n3180) );
  NAND2_X1 U4032 ( .A1(n3180), .A2(n3312), .ZN(n3277) );
  OAI21_X1 U4033 ( .B1(n3277), .B2(n3181), .A(STATE_REG_SCAN_IN), .ZN(n3184)
         );
  NAND2_X1 U4034 ( .A1(n3182), .A2(n4067), .ZN(n3278) );
  AND2_X1 U4035 ( .A1(n3278), .A2(n4070), .ZN(n3183) );
  AND2_X1 U4036 ( .A1(n3188), .A2(n3187), .ZN(n3189) );
  NAND2_X1 U4037 ( .A1(n3190), .A2(n3189), .ZN(U3211) );
  INV_X1 U4038 ( .A(REG1_REG_29__SCAN_IN), .ZN(n3204) );
  NAND2_X1 U4039 ( .A1(n2493), .A2(DATAI_29_), .ZN(n4138) );
  XNOR2_X1 U4040 ( .A(n4073), .B(n4138), .ZN(n3955) );
  INV_X1 U4041 ( .A(n3194), .ZN(n3933) );
  NAND2_X1 U4042 ( .A1(n4591), .A2(B_REG_SCAN_IN), .ZN(n3197) );
  AND2_X1 U40430 ( .A1(n4478), .A2(n3197), .ZN(n4129) );
  INV_X1 U4044 ( .A(REG2_REG_30__SCAN_IN), .ZN(n3200) );
  NAND2_X1 U4045 ( .A1(n2735), .A2(REG1_REG_30__SCAN_IN), .ZN(n3199) );
  NAND2_X1 U4046 ( .A1(n2715), .A2(REG0_REG_30__SCAN_IN), .ZN(n3198) );
  OAI211_X1 U4047 ( .C1(n3915), .C2(n3200), .A(n3199), .B(n3198), .ZN(n4072)
         );
  AOI22_X1 U4048 ( .A1(n3201), .A2(n4375), .B1(n4129), .B2(n4072), .ZN(n4141)
         );
  NAND2_X1 U4049 ( .A1(n4140), .A2(n4411), .ZN(n3202) );
  OAI211_X1 U4050 ( .C1(n4138), .C2(n4309), .A(n4141), .B(n3202), .ZN(n3203)
         );
  AOI21_X1 U4051 ( .B1(n4136), .B2(n4745), .A(n3203), .ZN(n3210) );
  INV_X1 U4052 ( .A(n3206), .ZN(n3207) );
  INV_X1 U4053 ( .A(n4138), .ZN(n3205) );
  OAI21_X2 U4054 ( .B1(n3207), .B2(n4138), .A(n2256), .ZN(n4143) );
  NAND2_X1 U4055 ( .A1(n3209), .A2(n3208), .ZN(U3547) );
  INV_X1 U4056 ( .A(REG0_REG_29__SCAN_IN), .ZN(n3211) );
  NAND2_X1 U4057 ( .A1(n3213), .A2(n3212), .ZN(U3515) );
  INV_X1 U4058 ( .A(n4716), .ZN(n3214) );
  OR2_X2 U4059 ( .A1(n3215), .A2(n3214), .ZN(n4086) );
  INV_X1 U4060 ( .A(n4086), .ZN(U4043) );
  INV_X1 U4061 ( .A(DATAI_3_), .ZN(n3216) );
  MUX2_X1 U4062 ( .A(n3216), .B(n2838), .S(STATE_REG_SCAN_IN), .Z(n3217) );
  INV_X1 U4063 ( .A(n3217), .ZN(U3349) );
  INV_X1 U4064 ( .A(DATAI_5_), .ZN(n3219) );
  MUX2_X1 U4065 ( .A(n2344), .B(n3219), .S(U3149), .Z(n3220) );
  INV_X1 U4066 ( .A(n3220), .ZN(U3347) );
  MUX2_X1 U4067 ( .A(n3254), .B(n2547), .S(U3149), .Z(n3221) );
  INV_X1 U4068 ( .A(n3221), .ZN(U3345) );
  INV_X1 U4069 ( .A(DATAI_25_), .ZN(n4864) );
  INV_X1 U4070 ( .A(n3222), .ZN(n3223) );
  NAND2_X1 U4071 ( .A1(n3223), .A2(STATE_REG_SCAN_IN), .ZN(n3224) );
  OAI21_X1 U4072 ( .B1(STATE_REG_SCAN_IN), .B2(n4864), .A(n3224), .ZN(U3327)
         );
  INV_X1 U4073 ( .A(DATAI_27_), .ZN(n5099) );
  NAND2_X1 U4074 ( .A1(n4591), .A2(STATE_REG_SCAN_IN), .ZN(n3225) );
  OAI21_X1 U4075 ( .B1(STATE_REG_SCAN_IN), .B2(n5099), .A(n3225), .ZN(U3325)
         );
  INV_X1 U4076 ( .A(DATAI_21_), .ZN(n5032) );
  NAND2_X1 U4077 ( .A1(n2757), .A2(STATE_REG_SCAN_IN), .ZN(n3226) );
  OAI21_X1 U4078 ( .B1(STATE_REG_SCAN_IN), .B2(n5032), .A(n3226), .ZN(U3331)
         );
  NAND2_X1 U4079 ( .A1(n3227), .A2(n3279), .ZN(n4714) );
  INV_X1 U4080 ( .A(D_REG_1__SCAN_IN), .ZN(n5118) );
  AOI22_X1 U4081 ( .A1(n4714), .A2(n5118), .B1(n3228), .B2(n4716), .ZN(U3459)
         );
  INV_X1 U4082 ( .A(D_REG_0__SCAN_IN), .ZN(n3231) );
  INV_X1 U4083 ( .A(n3229), .ZN(n3230) );
  AOI22_X1 U4084 ( .A1(n4714), .A2(n3231), .B1(n3230), .B2(n4716), .ZN(U3458)
         );
  INV_X1 U4085 ( .A(DATAI_29_), .ZN(n4903) );
  NAND2_X1 U4086 ( .A1(n3232), .A2(STATE_REG_SCAN_IN), .ZN(n3233) );
  OAI21_X1 U4087 ( .B1(STATE_REG_SCAN_IN), .B2(n4903), .A(n3233), .ZN(U3323)
         );
  NOR2_X1 U4088 ( .A1(n4683), .A2(U4043), .ZN(U3148) );
  INV_X1 U4089 ( .A(n4684), .ZN(n3275) );
  AOI211_X1 U4090 ( .C1(n3236), .C2(n3235), .A(n3234), .B(n3275), .ZN(n3243)
         );
  AOI211_X1 U4091 ( .C1(n3239), .C2(n3238), .A(n3237), .B(n4677), .ZN(n3242)
         );
  INV_X1 U4092 ( .A(REG3_REG_5__SCAN_IN), .ZN(n4886) );
  NOR2_X1 U4093 ( .A1(STATE_REG_SCAN_IN), .A2(n4886), .ZN(n3835) );
  AOI21_X1 U4094 ( .B1(n4683), .B2(ADDR_REG_5__SCAN_IN), .A(n3835), .ZN(n3240)
         );
  OAI21_X1 U4095 ( .B1(n4689), .B2(n2344), .A(n3240), .ZN(n3241) );
  OR3_X1 U4096 ( .A1(n3243), .A2(n3242), .A3(n3241), .ZN(U3245) );
  AOI211_X1 U4097 ( .C1(n3246), .C2(n3245), .A(n4677), .B(n3244), .ZN(n3257)
         );
  INV_X1 U4098 ( .A(n3247), .ZN(n3249) );
  NAND2_X1 U4099 ( .A1(n3249), .A2(n3248), .ZN(n3251) );
  OAI21_X1 U4100 ( .B1(n3252), .B2(n3251), .A(n4684), .ZN(n3250) );
  AOI21_X1 U4101 ( .B1(n3252), .B2(n3251), .A(n3250), .ZN(n3256) );
  INV_X1 U4102 ( .A(REG3_REG_7__SCAN_IN), .ZN(n5039) );
  NOR2_X1 U4103 ( .A1(STATE_REG_SCAN_IN), .A2(n5039), .ZN(n3515) );
  AOI21_X1 U4104 ( .B1(n4683), .B2(ADDR_REG_7__SCAN_IN), .A(n3515), .ZN(n3253)
         );
  OAI21_X1 U4105 ( .B1(n4689), .B2(n3254), .A(n3253), .ZN(n3255) );
  OR3_X1 U4106 ( .A1(n3257), .A2(n3256), .A3(n3255), .ZN(U3247) );
  XNOR2_X1 U4107 ( .A(n3258), .B(REG2_REG_6__SCAN_IN), .ZN(n3267) );
  INV_X1 U4108 ( .A(n4689), .ZN(n4103) );
  NOR2_X1 U4109 ( .A1(STATE_REG_SCAN_IN), .A2(n3259), .ZN(n3456) );
  AOI21_X1 U4110 ( .B1(n4683), .B2(ADDR_REG_6__SCAN_IN), .A(n3456), .ZN(n3260)
         );
  INV_X1 U4111 ( .A(n3260), .ZN(n3265) );
  AOI211_X1 U4112 ( .C1(n3263), .C2(n3262), .A(n3275), .B(n3261), .ZN(n3264)
         );
  AOI211_X1 U4113 ( .C1(n4103), .C2(n4565), .A(n3265), .B(n3264), .ZN(n3266)
         );
  OAI21_X1 U4114 ( .B1(n3267), .B2(n4677), .A(n3266), .ZN(U3246) );
  XOR2_X1 U4115 ( .A(REG1_REG_8__SCAN_IN), .B(n3268), .Z(n3276) );
  XNOR2_X1 U4116 ( .A(REG2_REG_8__SCAN_IN), .B(n3269), .ZN(n3270) );
  NAND2_X1 U4117 ( .A1(n4640), .A2(n3270), .ZN(n3271) );
  NAND2_X1 U4118 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3529) );
  NAND2_X1 U4119 ( .A1(n3271), .A2(n3529), .ZN(n3272) );
  AOI21_X1 U4120 ( .B1(n4683), .B2(ADDR_REG_8__SCAN_IN), .A(n3272), .ZN(n3274)
         );
  NAND2_X1 U4121 ( .A1(n4103), .A2(n4564), .ZN(n3273) );
  OAI211_X1 U4122 ( .C1(n3276), .C2(n3275), .A(n3274), .B(n3273), .ZN(U3248)
         );
  INV_X1 U4123 ( .A(n3277), .ZN(n3280) );
  NAND3_X1 U4124 ( .A1(n3280), .A2(n3279), .A3(n3278), .ZN(n3303) );
  INV_X1 U4125 ( .A(n3303), .ZN(n3289) );
  INV_X1 U4126 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3288) );
  OAI211_X1 U4127 ( .C1(n3283), .C2(n3282), .A(n3281), .B(n4581), .ZN(n3287)
         );
  INV_X1 U4128 ( .A(n2925), .ZN(n3284) );
  INV_X1 U4129 ( .A(n2949), .ZN(n3427) );
  OAI22_X1 U4130 ( .A1(n3284), .A2(n4571), .B1(n3427), .B2(n3875), .ZN(n3285)
         );
  AOI21_X1 U4131 ( .B1(n2935), .B2(n3904), .A(n3285), .ZN(n3286) );
  OAI211_X1 U4132 ( .C1(n3289), .C2(n3288), .A(n3287), .B(n3286), .ZN(U3219)
         );
  OAI21_X1 U4133 ( .B1(n3292), .B2(n3291), .A(n3290), .ZN(n3329) );
  INV_X1 U4134 ( .A(n3904), .ZN(n4574) );
  OAI22_X1 U4135 ( .A1(n4574), .A2(n3307), .B1(n2476), .B2(n3875), .ZN(n3293)
         );
  AOI21_X1 U4136 ( .B1(REG3_REG_0__SCAN_IN), .B2(n3303), .A(n3293), .ZN(n3294)
         );
  OAI21_X1 U4137 ( .B1(n3329), .B2(n3861), .A(n3294), .ZN(U3229) );
  INV_X1 U4138 ( .A(n3298), .ZN(n3299) );
  AOI21_X1 U4139 ( .B1(n3295), .B2(n3296), .A(n3299), .ZN(n3305) );
  AOI22_X1 U4140 ( .A1(n4577), .A2(n4085), .B1(n3905), .B2(n2484), .ZN(n3300)
         );
  OAI21_X1 U4141 ( .B1(n4574), .B2(n3301), .A(n3300), .ZN(n3302) );
  AOI21_X1 U4142 ( .B1(REG3_REG_2__SCAN_IN), .B2(n3303), .A(n3302), .ZN(n3304)
         );
  OAI21_X1 U4143 ( .B1(n3305), .B2(n3861), .A(n3304), .ZN(U3234) );
  NOR2_X1 U4144 ( .A1(n3307), .A2(n3306), .ZN(n4731) );
  INV_X1 U4145 ( .A(n3738), .ZN(n3697) );
  NAND2_X1 U4146 ( .A1(n2925), .A2(n3307), .ZN(n3992) );
  NAND2_X1 U4147 ( .A1(n3356), .A2(n3992), .ZN(n4732) );
  OAI21_X1 U4148 ( .B1(n3697), .B2(n4375), .A(n4732), .ZN(n3308) );
  OAI21_X1 U4149 ( .B1(n2476), .B2(n4415), .A(n3308), .ZN(n4730) );
  AOI21_X1 U4150 ( .B1(n4731), .B2(n3309), .A(n4730), .ZN(n3320) );
  OAI21_X1 U4151 ( .B1(n5118), .B2(n3310), .A(n4714), .ZN(n3314) );
  NAND4_X1 U4152 ( .A1(n3314), .A2(n3313), .A3(n3312), .A4(n3311), .ZN(n3315)
         );
  OR2_X1 U4153 ( .A1(n2921), .A2(n4123), .ZN(n3398) );
  INV_X1 U4154 ( .A(n3398), .ZN(n3316) );
  NAND2_X1 U4155 ( .A1(n4209), .A2(n3316), .ZN(n3451) );
  INV_X1 U4156 ( .A(n3451), .ZN(n4708) );
  OAI22_X1 U4157 ( .A1(n4209), .A2(n3327), .B1(n3317), .B2(n4369), .ZN(n3318)
         );
  AOI21_X1 U4158 ( .B1(n4708), .B2(n4732), .A(n3318), .ZN(n3319) );
  OAI21_X1 U4159 ( .B1(n3320), .B2(n4713), .A(n3319), .ZN(U3290) );
  XOR2_X1 U4160 ( .A(n3321), .B(n3322), .Z(n3326) );
  INV_X1 U4161 ( .A(n4084), .ZN(n3422) );
  OAI22_X1 U4162 ( .A1(n3427), .A2(n4571), .B1(n3422), .B2(n3875), .ZN(n3324)
         );
  MUX2_X1 U4163 ( .A(n3185), .B(U3149), .S(REG3_REG_3__SCAN_IN), .Z(n3323) );
  AOI211_X1 U4164 ( .C1(n3374), .C2(n3904), .A(n3324), .B(n3323), .ZN(n3325)
         );
  OAI21_X1 U4165 ( .B1(n3326), .B2(n3861), .A(n3325), .ZN(U3215) );
  AND2_X1 U4166 ( .A1(n4591), .A2(n3327), .ZN(n3328) );
  OR2_X1 U4167 ( .A1(n4570), .A2(n3328), .ZN(n4592) );
  NAND2_X1 U4168 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n4090) );
  NOR2_X1 U4169 ( .A1(n3329), .A2(n4591), .ZN(n3330) );
  AOI211_X1 U4170 ( .C1(n4591), .C2(n4090), .A(n4570), .B(n3330), .ZN(n3331)
         );
  AOI22_X1 U4171 ( .A1(n4683), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3332) );
  OAI21_X1 U4172 ( .B1(n4689), .B2(n3333), .A(n3332), .ZN(n3343) );
  OR3_X1 U4173 ( .A1(n4092), .A2(n3337), .A3(n3336), .ZN(n3338) );
  NAND3_X1 U4174 ( .A1(n4640), .A2(n3339), .A3(n3338), .ZN(n3340) );
  NAND2_X1 U4175 ( .A1(n3341), .A2(n3340), .ZN(n3342) );
  OR3_X1 U4176 ( .A1(n3350), .A2(n3343), .A3(n3342), .ZN(U3242) );
  XNOR2_X1 U4177 ( .A(n3344), .B(REG2_REG_4__SCAN_IN), .ZN(n3352) );
  OAI211_X1 U4178 ( .C1(REG1_REG_4__SCAN_IN), .C2(n3346), .A(n4684), .B(n3345), 
        .ZN(n3348) );
  AND2_X1 U4179 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3414) );
  AOI21_X1 U4180 ( .B1(n4683), .B2(ADDR_REG_4__SCAN_IN), .A(n3414), .ZN(n3347)
         );
  OAI211_X1 U4181 ( .C1(n4689), .C2(n3349), .A(n3348), .B(n3347), .ZN(n3351)
         );
  AOI211_X1 U4182 ( .C1(n4640), .C2(n3352), .A(n3351), .B(n3350), .ZN(n3353)
         );
  INV_X1 U4183 ( .A(n3353), .ZN(U3244) );
  OAI21_X1 U4184 ( .B1(n2765), .B2(n3355), .A(n3354), .ZN(n4734) );
  INV_X1 U4185 ( .A(n3356), .ZN(n3994) );
  XNOR2_X1 U4186 ( .A(n2765), .B(n3994), .ZN(n3363) );
  OR2_X1 U4187 ( .A1(n4734), .A2(n3738), .ZN(n3362) );
  NAND2_X1 U4188 ( .A1(n2925), .A2(n4411), .ZN(n3358) );
  NAND2_X1 U4189 ( .A1(n2949), .A2(n4478), .ZN(n3357) );
  OAI211_X1 U4190 ( .C1(n4309), .C2(n3359), .A(n3358), .B(n3357), .ZN(n3360)
         );
  INV_X1 U4191 ( .A(n3360), .ZN(n3361) );
  OAI211_X1 U4192 ( .C1(n4312), .C2(n3363), .A(n3362), .B(n3361), .ZN(n4735)
         );
  MUX2_X1 U4193 ( .A(n4735), .B(REG2_REG_1__SCAN_IN), .S(n4713), .Z(n3364) );
  INV_X1 U4194 ( .A(n3364), .ZN(n3369) );
  AND2_X1 U4195 ( .A1(n4738), .A2(n4123), .ZN(n3365) );
  INV_X1 U4196 ( .A(n3390), .ZN(n3366) );
  AOI21_X1 U4197 ( .B1(n3367), .B2(n2935), .A(n3366), .ZN(n4737) );
  INV_X1 U4198 ( .A(n4369), .ZN(n4705) );
  AOI22_X1 U4199 ( .A1(n4707), .A2(n4737), .B1(REG3_REG_1__SCAN_IN), .B2(n4705), .ZN(n3368) );
  OAI211_X1 U4200 ( .C1(n4734), .C2(n3451), .A(n3369), .B(n3368), .ZN(U3289)
         );
  INV_X1 U4201 ( .A(n3371), .ZN(n3958) );
  XNOR2_X1 U4202 ( .A(n3370), .B(n3958), .ZN(n3419) );
  XNOR2_X1 U4203 ( .A(n3372), .B(n3371), .ZN(n3373) );
  NAND2_X1 U4204 ( .A1(n3373), .A2(n4375), .ZN(n3420) );
  AOI22_X1 U4205 ( .A1(n4084), .A2(n4478), .B1(n4477), .B2(n3374), .ZN(n3375)
         );
  OAI211_X1 U4206 ( .C1(n3427), .C2(n4481), .A(n3420), .B(n3375), .ZN(n3376)
         );
  AOI21_X1 U4207 ( .B1(n4745), .B2(n3419), .A(n3376), .ZN(n3397) );
  NOR2_X1 U4208 ( .A1(n3392), .A2(n3421), .ZN(n3377) );
  NOR2_X1 U4209 ( .A1(n3377), .A2(n3446), .ZN(n3423) );
  INV_X1 U4210 ( .A(n4556), .ZN(n4509) );
  AOI22_X1 U4211 ( .A1(n3423), .A2(n4509), .B1(REG0_REG_3__SCAN_IN), .B2(n4757), .ZN(n3378) );
  OAI21_X1 U4212 ( .B1(n3397), .B2(n4757), .A(n3378), .ZN(U3473) );
  INV_X1 U4213 ( .A(n4733), .ZN(n4756) );
  OAI21_X1 U4214 ( .B1(n3380), .B2(n3957), .A(n3379), .ZN(n4709) );
  XNOR2_X1 U4215 ( .A(n3382), .B(n3381), .ZN(n3387) );
  INV_X1 U4216 ( .A(n4085), .ZN(n3385) );
  NAND2_X1 U4217 ( .A1(n4709), .A2(n3697), .ZN(n3384) );
  AOI22_X1 U4218 ( .A1(n2484), .A2(n4411), .B1(n3389), .B2(n4477), .ZN(n3383)
         );
  OAI211_X1 U4219 ( .C1(n3385), .C2(n4415), .A(n3384), .B(n3383), .ZN(n3386)
         );
  AOI21_X1 U4220 ( .B1(n3387), .B2(n4375), .A(n3386), .ZN(n4712) );
  INV_X1 U4221 ( .A(n4712), .ZN(n3388) );
  AOI21_X1 U4222 ( .B1(n4756), .B2(n4709), .A(n3388), .ZN(n3395) );
  AND2_X1 U4223 ( .A1(n3390), .A2(n3389), .ZN(n3391) );
  NOR2_X1 U4224 ( .A1(n3392), .A2(n3391), .ZN(n4706) );
  AOI22_X1 U4225 ( .A1(n4408), .A2(n4706), .B1(n4767), .B2(REG1_REG_2__SCAN_IN), .ZN(n3393) );
  OAI21_X1 U4226 ( .B1(n3395), .B2(n4767), .A(n3393), .ZN(U3520) );
  AOI22_X1 U4227 ( .A1(n4509), .A2(n4706), .B1(n4757), .B2(REG0_REG_2__SCAN_IN), .ZN(n3394) );
  OAI21_X1 U4228 ( .B1(n3395), .B2(n4757), .A(n3394), .ZN(U3471) );
  AOI22_X1 U4229 ( .A1(n3423), .A2(n4408), .B1(REG1_REG_3__SCAN_IN), .B2(n4767), .ZN(n3396) );
  OAI21_X1 U4230 ( .B1(n3397), .B2(n4767), .A(n3396), .ZN(U3521) );
  NAND2_X1 U4231 ( .A1(n3738), .A2(n3398), .ZN(n3399) );
  XNOR2_X1 U4232 ( .A(n4083), .B(n3478), .ZN(n3986) );
  XNOR2_X1 U4233 ( .A(n3400), .B(n3986), .ZN(n3483) );
  XOR2_X1 U4234 ( .A(n3986), .B(n3401), .Z(n3402) );
  NOR2_X1 U4235 ( .A1(n3402), .A2(n4312), .ZN(n3480) );
  AND2_X1 U4236 ( .A1(n3444), .A2(n3836), .ZN(n3403) );
  NOR2_X1 U4237 ( .A1(n3466), .A2(n3403), .ZN(n3510) );
  NAND2_X1 U4238 ( .A1(n3510), .A2(n4707), .ZN(n3407) );
  NAND2_X1 U4239 ( .A1(n4209), .A2(n4477), .ZN(n4356) );
  INV_X1 U4240 ( .A(n4356), .ZN(n4215) );
  OAI22_X1 U4241 ( .A1(n4209), .A2(n2343), .B1(n3837), .B2(n4369), .ZN(n3404)
         );
  AOI21_X1 U4242 ( .B1(n3836), .B2(n4215), .A(n3404), .ZN(n3406) );
  NAND2_X1 U4243 ( .A1(n4209), .A2(n4478), .ZN(n4293) );
  INV_X1 U4244 ( .A(n4293), .ZN(n4351) );
  AND2_X1 U4245 ( .A1(n4209), .A2(n4411), .ZN(n4350) );
  AOI22_X1 U4246 ( .A1(n4351), .A2(n4082), .B1(n4350), .B2(n4084), .ZN(n3405)
         );
  NAND3_X1 U4247 ( .A1(n3407), .A2(n3406), .A3(n3405), .ZN(n3408) );
  AOI21_X1 U4248 ( .B1(n3480), .B2(n4209), .A(n3408), .ZN(n3409) );
  OAI21_X1 U4249 ( .B1(n4382), .B2(n3483), .A(n3409), .ZN(U3285) );
  INV_X1 U4250 ( .A(n3411), .ZN(n3412) );
  AOI211_X1 U4251 ( .C1(n3413), .C2(n3410), .A(n3861), .B(n3412), .ZN(n3418)
         );
  AOI21_X1 U4252 ( .B1(n4577), .B2(n4083), .A(n3414), .ZN(n3416) );
  AOI22_X1 U4253 ( .A1(n3905), .A2(n4085), .B1(n3904), .B2(n3438), .ZN(n3415)
         );
  OAI211_X1 U4254 ( .C1(n4586), .C2(n3447), .A(n3416), .B(n3415), .ZN(n3417)
         );
  OR2_X1 U4255 ( .A1(n3418), .A2(n3417), .ZN(U3227) );
  INV_X1 U4256 ( .A(n3419), .ZN(n3432) );
  INV_X1 U4257 ( .A(n3420), .ZN(n3430) );
  OAI22_X1 U4258 ( .A1(n3422), .A2(n4293), .B1(n4356), .B2(n3421), .ZN(n3429)
         );
  INV_X1 U4259 ( .A(n4350), .ZN(n4291) );
  NAND2_X1 U4260 ( .A1(n3423), .A2(n4707), .ZN(n3426) );
  OAI22_X1 U4261 ( .A1(n4209), .A2(n4104), .B1(REG3_REG_3__SCAN_IN), .B2(n4369), .ZN(n3424) );
  INV_X1 U4262 ( .A(n3424), .ZN(n3425) );
  OAI211_X1 U4263 ( .C1(n3427), .C2(n4291), .A(n3426), .B(n3425), .ZN(n3428)
         );
  AOI211_X1 U4264 ( .C1(n3430), .C2(n4209), .A(n3429), .B(n3428), .ZN(n3431)
         );
  OAI21_X1 U4265 ( .B1(n3432), .B2(n4382), .A(n3431), .ZN(U3287) );
  NAND2_X1 U4266 ( .A1(n3434), .A2(n3967), .ZN(n3435) );
  NAND2_X1 U4267 ( .A1(n3436), .A2(n3435), .ZN(n4739) );
  XNOR2_X1 U4268 ( .A(n3437), .B(n3967), .ZN(n3442) );
  AOI22_X1 U4269 ( .A1(n4085), .A2(n4411), .B1(n3438), .B2(n4477), .ZN(n3440)
         );
  NAND2_X1 U4270 ( .A1(n4083), .A2(n4478), .ZN(n3439) );
  OAI211_X1 U4271 ( .C1(n4739), .C2(n3738), .A(n3440), .B(n3439), .ZN(n3441)
         );
  AOI21_X1 U4272 ( .B1(n3442), .B2(n4375), .A(n3441), .ZN(n3443) );
  INV_X1 U4273 ( .A(n3443), .ZN(n4741) );
  OAI211_X1 U4274 ( .C1(n3446), .C2(n3445), .A(n4738), .B(n3444), .ZN(n4740)
         );
  OAI22_X1 U4275 ( .A1(n4740), .A2(n4563), .B1(n4369), .B2(n3447), .ZN(n3448)
         );
  OAI21_X1 U4276 ( .B1(n4741), .B2(n3448), .A(n4209), .ZN(n3450) );
  NAND2_X1 U4277 ( .A1(n4713), .A2(REG2_REG_4__SCAN_IN), .ZN(n3449) );
  OAI211_X1 U4278 ( .C1(n4739), .C2(n3451), .A(n3450), .B(n3449), .ZN(U3286)
         );
  XNOR2_X1 U4279 ( .A(n3453), .B(n3452), .ZN(n3454) );
  XNOR2_X1 U4280 ( .A(n3455), .B(n3454), .ZN(n3460) );
  AOI21_X1 U4281 ( .B1(n4577), .B2(n4081), .A(n3456), .ZN(n3458) );
  AOI22_X1 U4282 ( .A1(n3905), .A2(n4083), .B1(n3904), .B2(n3497), .ZN(n3457)
         );
  OAI211_X1 U4283 ( .C1(n4586), .C2(n3471), .A(n3458), .B(n3457), .ZN(n3459)
         );
  AOI21_X1 U4284 ( .B1(n3460), .B2(n4581), .A(n3459), .ZN(n3461) );
  INV_X1 U4285 ( .A(n3461), .ZN(U3236) );
  INV_X1 U4286 ( .A(n3462), .ZN(n4017) );
  OR2_X1 U4287 ( .A1(n4007), .A2(n4017), .ZN(n3964) );
  XOR2_X1 U4288 ( .A(n3964), .B(n3463), .Z(n3464) );
  NAND2_X1 U4289 ( .A1(n3464), .A2(n4375), .ZN(n3499) );
  XOR2_X1 U4290 ( .A(n3964), .B(n3465), .Z(n3502) );
  NAND2_X1 U4291 ( .A1(n3502), .A2(n4347), .ZN(n3477) );
  INV_X1 U4292 ( .A(n3466), .ZN(n3468) );
  INV_X1 U4293 ( .A(n3486), .ZN(n3467) );
  AOI21_X1 U4294 ( .B1(n3497), .B2(n3468), .A(n3467), .ZN(n3506) );
  NAND2_X1 U4295 ( .A1(n4350), .A2(n4083), .ZN(n3470) );
  NAND2_X1 U4296 ( .A1(n4713), .A2(REG2_REG_6__SCAN_IN), .ZN(n3469) );
  OAI211_X1 U4297 ( .C1(n4369), .C2(n3471), .A(n3470), .B(n3469), .ZN(n3475)
         );
  INV_X1 U4298 ( .A(n4081), .ZN(n3473) );
  OAI22_X1 U4299 ( .A1(n3473), .A2(n4293), .B1(n4356), .B2(n3472), .ZN(n3474)
         );
  AOI211_X1 U4300 ( .C1(n3506), .C2(n4707), .A(n3475), .B(n3474), .ZN(n3476)
         );
  OAI211_X1 U4301 ( .C1(n4713), .C2(n3499), .A(n3477), .B(n3476), .ZN(U3284)
         );
  INV_X1 U4302 ( .A(n4082), .ZN(n3479) );
  OAI22_X1 U4303 ( .A1(n3479), .A2(n4415), .B1(n4309), .B2(n3478), .ZN(n3481)
         );
  AOI211_X1 U4304 ( .C1(n4411), .C2(n4084), .A(n3481), .B(n3480), .ZN(n3482)
         );
  OAI21_X1 U4305 ( .B1(n4452), .B2(n3483), .A(n3482), .ZN(n3509) );
  INV_X1 U4306 ( .A(n3509), .ZN(n3485) );
  AOI22_X1 U4307 ( .A1(n3510), .A2(n4509), .B1(REG0_REG_5__SCAN_IN), .B2(n4757), .ZN(n3484) );
  OAI21_X1 U4308 ( .B1(n3485), .B2(n4757), .A(n3484), .ZN(U3477) );
  INV_X1 U4309 ( .A(n4738), .ZN(n4751) );
  AOI211_X1 U4310 ( .C1(n3516), .C2(n3486), .A(n4751), .B(n2828), .ZN(n4747)
         );
  XNOR2_X1 U4311 ( .A(n3487), .B(n3966), .ZN(n3490) );
  AOI22_X1 U4312 ( .A1(n4080), .A2(n4478), .B1(n4477), .B2(n3516), .ZN(n3489)
         );
  NAND2_X1 U4313 ( .A1(n4082), .A2(n4411), .ZN(n3488) );
  OAI211_X1 U4314 ( .C1(n3490), .C2(n4312), .A(n3489), .B(n3488), .ZN(n4749)
         );
  AOI21_X1 U4315 ( .B1(n4747), .B2(n4123), .A(n4749), .ZN(n3496) );
  OAI22_X1 U4316 ( .A1(n4209), .A2(n2540), .B1(n3519), .B2(n4369), .ZN(n3491)
         );
  INV_X1 U4317 ( .A(n3491), .ZN(n3495) );
  NAND2_X1 U4318 ( .A1(n3493), .A2(n3966), .ZN(n4746) );
  NAND3_X1 U4319 ( .A1(n3492), .A2(n4746), .A3(n4347), .ZN(n3494) );
  OAI211_X1 U4320 ( .C1(n3496), .C2(n4713), .A(n3495), .B(n3494), .ZN(U3283)
         );
  INV_X1 U4321 ( .A(n4083), .ZN(n3500) );
  AOI22_X1 U4322 ( .A1(n4081), .A2(n4478), .B1(n3497), .B2(n4477), .ZN(n3498)
         );
  OAI211_X1 U4323 ( .C1(n3500), .C2(n4481), .A(n3499), .B(n3498), .ZN(n3501)
         );
  AOI21_X1 U4324 ( .B1(n3502), .B2(n4745), .A(n3501), .ZN(n3508) );
  INV_X1 U4325 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3503) );
  NOR2_X1 U4326 ( .A1(n4759), .A2(n3503), .ZN(n3504) );
  AOI21_X1 U4327 ( .B1(n3506), .B2(n4509), .A(n3504), .ZN(n3505) );
  OAI21_X1 U4328 ( .B1(n3508), .B2(n4757), .A(n3505), .ZN(U3479) );
  AOI22_X1 U4329 ( .A1(n3506), .A2(n4408), .B1(n4767), .B2(REG1_REG_6__SCAN_IN), .ZN(n3507) );
  OAI21_X1 U4330 ( .B1(n3508), .B2(n4767), .A(n3507), .ZN(U3524) );
  INV_X1 U4331 ( .A(REG1_REG_5__SCAN_IN), .ZN(n3513) );
  NAND2_X1 U4332 ( .A1(n3509), .A2(n4770), .ZN(n3512) );
  NAND2_X1 U4333 ( .A1(n3510), .A2(n4408), .ZN(n3511) );
  OAI211_X1 U4334 ( .C1(n4770), .C2(n3513), .A(n3512), .B(n3511), .ZN(U3523)
         );
  XOR2_X1 U4335 ( .A(n3514), .B(n3523), .Z(n3521) );
  AOI21_X1 U4336 ( .B1(n4577), .B2(n4080), .A(n3515), .ZN(n3518) );
  AOI22_X1 U4337 ( .A1(n3905), .A2(n4082), .B1(n3904), .B2(n3516), .ZN(n3517)
         );
  OAI211_X1 U4338 ( .C1(n4586), .C2(n3519), .A(n3518), .B(n3517), .ZN(n3520)
         );
  AOI21_X1 U4339 ( .B1(n3521), .B2(n4581), .A(n3520), .ZN(n3522) );
  INV_X1 U4340 ( .A(n3522), .ZN(U3210) );
  NAND2_X1 U4341 ( .A1(n3514), .A2(n3523), .ZN(n3525) );
  NAND2_X1 U4342 ( .A1(n3525), .A2(n3524), .ZN(n3528) );
  NAND2_X1 U4343 ( .A1(n2255), .A2(n3526), .ZN(n3527) );
  XNOR2_X1 U4344 ( .A(n3528), .B(n3527), .ZN(n3535) );
  INV_X1 U4345 ( .A(n3529), .ZN(n3530) );
  AOI21_X1 U4346 ( .B1(n4577), .B2(n4079), .A(n3530), .ZN(n3532) );
  AOI22_X1 U4347 ( .A1(n3905), .A2(n4081), .B1(n3904), .B2(n3579), .ZN(n3531)
         );
  OAI211_X1 U4348 ( .C1(n4586), .C2(n3533), .A(n3532), .B(n3531), .ZN(n3534)
         );
  AOI21_X1 U4349 ( .B1(n3535), .B2(n4581), .A(n3534), .ZN(n3536) );
  INV_X1 U4350 ( .A(n3536), .ZN(U3218) );
  NAND2_X1 U4351 ( .A1(n3492), .A2(n3537), .ZN(n3539) );
  AND2_X1 U4352 ( .A1(n3539), .A2(n3538), .ZN(n3540) );
  NAND2_X1 U4353 ( .A1(n2304), .A2(n4014), .ZN(n3965) );
  XNOR2_X1 U4354 ( .A(n3540), .B(n3965), .ZN(n3603) );
  XOR2_X1 U4355 ( .A(n3965), .B(n3541), .Z(n3542) );
  NOR2_X1 U4356 ( .A1(n3542), .A2(n4312), .ZN(n3600) );
  NAND2_X1 U4357 ( .A1(n3600), .A2(n4209), .ZN(n3550) );
  AND2_X1 U4358 ( .A1(n3582), .A2(n3555), .ZN(n3543) );
  NOR2_X1 U4359 ( .A1(n2254), .A2(n3543), .ZN(n3607) );
  OAI22_X1 U4360 ( .A1(n3558), .A2(n4369), .B1(n2562), .B2(n4209), .ZN(n3547)
         );
  INV_X1 U4361 ( .A(n4078), .ZN(n3599) );
  NAND2_X1 U4362 ( .A1(n4350), .A2(n4080), .ZN(n3545) );
  OR2_X1 U4363 ( .A1(n4356), .A2(n3598), .ZN(n3544) );
  OAI211_X1 U4364 ( .C1(n3599), .C2(n4293), .A(n3545), .B(n3544), .ZN(n3546)
         );
  OR2_X1 U4365 ( .A1(n3547), .A2(n3546), .ZN(n3548) );
  AOI21_X1 U4366 ( .B1(n3607), .B2(n4707), .A(n3548), .ZN(n3549) );
  OAI211_X1 U4367 ( .C1(n3603), .C2(n4382), .A(n3550), .B(n3549), .ZN(U3281)
         );
  AND2_X1 U4368 ( .A1(n3552), .A2(n3551), .ZN(n3554) );
  XNOR2_X1 U4369 ( .A(n3554), .B(n3553), .ZN(n3560) );
  NOR2_X1 U4370 ( .A1(STATE_REG_SCAN_IN), .A2(n2559), .ZN(n4606) );
  AOI21_X1 U4371 ( .B1(n4577), .B2(n4078), .A(n4606), .ZN(n3557) );
  AOI22_X1 U4372 ( .A1(n3905), .A2(n4080), .B1(n3904), .B2(n3555), .ZN(n3556)
         );
  OAI211_X1 U4373 ( .C1(n4586), .C2(n3558), .A(n3557), .B(n3556), .ZN(n3559)
         );
  AOI21_X1 U4374 ( .B1(n3560), .B2(n4581), .A(n3559), .ZN(n3561) );
  INV_X1 U4375 ( .A(n3561), .ZN(U3228) );
  INV_X1 U4376 ( .A(n3563), .ZN(n3564) );
  AOI211_X1 U4377 ( .C1(n3565), .C2(n3562), .A(n3861), .B(n3564), .ZN(n3570)
         );
  NAND2_X1 U4378 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4611) );
  INV_X1 U4379 ( .A(n4611), .ZN(n3566) );
  AOI21_X1 U4380 ( .B1(n3905), .B2(n4079), .A(n3566), .ZN(n3568) );
  AOI22_X1 U4381 ( .A1(n4577), .A2(n4077), .B1(n3904), .B2(n3692), .ZN(n3567)
         );
  OAI211_X1 U4382 ( .C1(n4586), .C2(n4690), .A(n3568), .B(n3567), .ZN(n3569)
         );
  OR2_X1 U4383 ( .A1(n3570), .A2(n3569), .ZN(U3214) );
  NAND2_X1 U4384 ( .A1(n4013), .A2(n4011), .ZN(n3961) );
  NAND2_X1 U4385 ( .A1(n3492), .A2(n3571), .ZN(n3572) );
  XOR2_X1 U4386 ( .A(n3961), .B(n3572), .Z(n4701) );
  INV_X1 U4387 ( .A(n4701), .ZN(n3578) );
  XOR2_X1 U4388 ( .A(n3961), .B(n3573), .Z(n3576) );
  AOI22_X1 U4389 ( .A1(n4081), .A2(n4411), .B1(n3579), .B2(n4477), .ZN(n3575)
         );
  NAND2_X1 U4390 ( .A1(n4079), .A2(n4478), .ZN(n3574) );
  OAI211_X1 U4391 ( .C1(n3576), .C2(n4312), .A(n3575), .B(n3574), .ZN(n3577)
         );
  AOI21_X1 U4392 ( .B1(n4701), .B2(n3697), .A(n3577), .ZN(n4704) );
  OAI21_X1 U4393 ( .B1(n4733), .B2(n3578), .A(n4704), .ZN(n3586) );
  NAND2_X1 U4394 ( .A1(n3580), .A2(n3579), .ZN(n3581) );
  NAND2_X1 U4395 ( .A1(n3582), .A2(n3581), .ZN(n4699) );
  INV_X1 U4396 ( .A(REG0_REG_8__SCAN_IN), .ZN(n4900) );
  OAI22_X1 U4397 ( .A1(n4699), .A2(n4556), .B1(n4759), .B2(n4900), .ZN(n3583)
         );
  AOI21_X1 U4398 ( .B1(n3586), .B2(n4759), .A(n3583), .ZN(n3584) );
  INV_X1 U4399 ( .A(n3584), .ZN(U3483) );
  OAI22_X1 U4400 ( .A1(n4699), .A2(n4491), .B1(n4770), .B2(n2887), .ZN(n3585)
         );
  AOI21_X1 U4401 ( .B1(n3586), .B2(n4770), .A(n3585), .ZN(n3587) );
  INV_X1 U4402 ( .A(n3587), .ZN(U3526) );
  XNOR2_X1 U4403 ( .A(n3590), .B(n3589), .ZN(n3591) );
  XNOR2_X1 U4404 ( .A(n3588), .B(n3591), .ZN(n3596) );
  AND2_X1 U4405 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4627) );
  AOI21_X1 U4406 ( .B1(n3905), .B2(n4078), .A(n4627), .ZN(n3594) );
  AOI22_X1 U4407 ( .A1(n4577), .A2(n4076), .B1(n3904), .B2(n3592), .ZN(n3593)
         );
  OAI211_X1 U4408 ( .C1(n4586), .C2(n3620), .A(n3594), .B(n3593), .ZN(n3595)
         );
  AOI21_X1 U4409 ( .B1(n3596), .B2(n4581), .A(n3595), .ZN(n3597) );
  INV_X1 U4410 ( .A(n3597), .ZN(U3233) );
  OAI22_X1 U4411 ( .A1(n3599), .A2(n4415), .B1(n4309), .B2(n3598), .ZN(n3601)
         );
  AOI211_X1 U4412 ( .C1(n4411), .C2(n4080), .A(n3601), .B(n3600), .ZN(n3602)
         );
  OAI21_X1 U4413 ( .B1(n4452), .B2(n3603), .A(n3602), .ZN(n3606) );
  INV_X1 U4414 ( .A(n3606), .ZN(n3605) );
  AOI22_X1 U4415 ( .A1(n3607), .A2(n4509), .B1(REG0_REG_9__SCAN_IN), .B2(n4757), .ZN(n3604) );
  OAI21_X1 U4416 ( .B1(n3605), .B2(n4757), .A(n3604), .ZN(U3485) );
  NAND2_X1 U4417 ( .A1(n3606), .A2(n4770), .ZN(n3609) );
  NAND2_X1 U4418 ( .A1(n3607), .A2(n4408), .ZN(n3608) );
  OAI211_X1 U4419 ( .C1(n4770), .C2(n2873), .A(n3609), .B(n3608), .ZN(U3527)
         );
  XNOR2_X1 U4420 ( .A(n3610), .B(n3968), .ZN(n3617) );
  OR2_X1 U4421 ( .A1(n3611), .A2(n3968), .ZN(n3612) );
  NAND2_X1 U4422 ( .A1(n3613), .A2(n3612), .ZN(n4755) );
  NAND2_X1 U4423 ( .A1(n4755), .A2(n3697), .ZN(n3616) );
  INV_X1 U4424 ( .A(n4076), .ZN(n3679) );
  OAI22_X1 U4425 ( .A1(n3679), .A2(n4415), .B1(n4309), .B2(n3618), .ZN(n3614)
         );
  AOI21_X1 U4426 ( .B1(n4411), .B2(n4078), .A(n3614), .ZN(n3615) );
  OAI211_X1 U4427 ( .C1(n4312), .C2(n3617), .A(n3616), .B(n3615), .ZN(n4753)
         );
  INV_X1 U4428 ( .A(n4753), .ZN(n3624) );
  INV_X1 U4429 ( .A(n3688), .ZN(n3619) );
  OAI21_X1 U4430 ( .B1(n3619), .B2(n3618), .A(n3637), .ZN(n4752) );
  NOR2_X1 U4431 ( .A1(n4752), .A2(n4317), .ZN(n3622) );
  OAI22_X1 U4432 ( .A1(n4209), .A2(n2585), .B1(n3620), .B2(n4369), .ZN(n3621)
         );
  AOI211_X1 U4433 ( .C1(n4755), .C2(n4708), .A(n3622), .B(n3621), .ZN(n3623)
         );
  OAI21_X1 U4434 ( .B1(n3624), .B2(n4713), .A(n3623), .ZN(U3279) );
  INV_X1 U4435 ( .A(n3626), .ZN(n3628) );
  NAND2_X1 U4436 ( .A1(n3628), .A2(n3627), .ZN(n3629) );
  XNOR2_X1 U4437 ( .A(n3625), .B(n3629), .ZN(n3634) );
  NOR2_X1 U4438 ( .A1(STATE_REG_SCAN_IN), .A2(n3630), .ZN(n4637) );
  AOI21_X1 U4439 ( .B1(n3905), .B2(n4077), .A(n4637), .ZN(n3632) );
  AOI22_X1 U4440 ( .A1(n4577), .A2(n4075), .B1(n3904), .B2(n3715), .ZN(n3631)
         );
  OAI211_X1 U4441 ( .C1(n4586), .C2(n3639), .A(n3632), .B(n3631), .ZN(n3633)
         );
  AOI21_X1 U4442 ( .B1(n3634), .B2(n4581), .A(n3633), .ZN(n3635) );
  INV_X1 U4443 ( .A(n3635), .ZN(U3221) );
  NAND2_X1 U4444 ( .A1(n3670), .A2(n3671), .ZN(n3963) );
  XNOR2_X1 U4445 ( .A(n3636), .B(n3963), .ZN(n3720) );
  AND2_X1 U4446 ( .A1(n3637), .A2(n3715), .ZN(n3638) );
  OR2_X1 U4447 ( .A1(n3638), .A2(n3682), .ZN(n3726) );
  OAI22_X1 U4448 ( .A1(n4209), .A2(n3640), .B1(n3639), .B2(n4369), .ZN(n3641)
         );
  AOI21_X1 U4449 ( .B1(n3715), .B2(n4215), .A(n3641), .ZN(n3643) );
  AOI22_X1 U4450 ( .A1(n4351), .A2(n4075), .B1(n4350), .B2(n4077), .ZN(n3642)
         );
  OAI211_X1 U4451 ( .C1(n3726), .C2(n4317), .A(n3643), .B(n3642), .ZN(n3649)
         );
  NAND2_X1 U4452 ( .A1(n3645), .A2(n3644), .ZN(n3673) );
  INV_X1 U4453 ( .A(n3963), .ZN(n3646) );
  XNOR2_X1 U4454 ( .A(n3673), .B(n3646), .ZN(n3647) );
  NAND2_X1 U4455 ( .A1(n3647), .A2(n4375), .ZN(n3718) );
  NOR2_X1 U4456 ( .A1(n3718), .A2(n4713), .ZN(n3648) );
  AOI211_X1 U4457 ( .C1(n4347), .C2(n3720), .A(n3649), .B(n3648), .ZN(n3650)
         );
  INV_X1 U4458 ( .A(n3650), .ZN(U3278) );
  NAND2_X1 U4459 ( .A1(n3735), .A2(n3917), .ZN(n3652) );
  INV_X1 U4460 ( .A(n3948), .ZN(n3651) );
  XNOR2_X1 U4461 ( .A(n3652), .B(n3651), .ZN(n3653) );
  NAND2_X1 U4462 ( .A1(n3653), .A2(n4375), .ZN(n4471) );
  XNOR2_X1 U4463 ( .A(n3654), .B(n3948), .ZN(n4474) );
  NAND2_X1 U4464 ( .A1(n4474), .A2(n4347), .ZN(n3663) );
  INV_X1 U4465 ( .A(n3740), .ZN(n3655) );
  OAI21_X1 U4466 ( .B1(n3655), .B2(n3659), .A(n4366), .ZN(n4548) );
  INV_X1 U4467 ( .A(n4548), .ZN(n3661) );
  AOI22_X1 U4468 ( .A1(n4351), .A2(n4469), .B1(n4350), .B2(n4467), .ZN(n3658)
         );
  INV_X1 U4469 ( .A(n3908), .ZN(n3656) );
  AOI22_X1 U4470 ( .A1(n4713), .A2(REG2_REG_15__SCAN_IN), .B1(n3656), .B2(
        n4705), .ZN(n3657) );
  OAI211_X1 U4471 ( .C1(n3659), .C2(n4356), .A(n3658), .B(n3657), .ZN(n3660)
         );
  AOI21_X1 U4472 ( .B1(n3661), .B2(n4707), .A(n3660), .ZN(n3662) );
  OAI211_X1 U4473 ( .C1(n4713), .C2(n4471), .A(n3663), .B(n3662), .ZN(U3275)
         );
  NAND2_X1 U4474 ( .A1(n3636), .A2(n3664), .ZN(n3666) );
  NAND2_X1 U4475 ( .A1(n3666), .A2(n3665), .ZN(n3669) );
  AND2_X1 U4476 ( .A1(n3668), .A2(n3667), .ZN(n3984) );
  INV_X1 U4477 ( .A(n3984), .ZN(n3674) );
  XNOR2_X1 U4478 ( .A(n3669), .B(n3674), .ZN(n4489) );
  INV_X1 U4479 ( .A(n4489), .ZN(n3687) );
  INV_X1 U4480 ( .A(n3670), .ZN(n3672) );
  OAI21_X1 U4481 ( .B1(n3673), .B2(n3672), .A(n3671), .ZN(n3675) );
  XNOR2_X1 U4482 ( .A(n3675), .B(n3674), .ZN(n3676) );
  NAND2_X1 U4483 ( .A1(n3676), .A2(n4375), .ZN(n3678) );
  AOI22_X1 U4484 ( .A1(n4467), .A2(n4478), .B1(n4477), .B2(n3708), .ZN(n3677)
         );
  OAI211_X1 U4485 ( .C1(n3679), .C2(n4481), .A(n3678), .B(n3677), .ZN(n4488)
         );
  INV_X1 U4486 ( .A(n3742), .ZN(n3680) );
  OAI21_X1 U4487 ( .B1(n3682), .B2(n3681), .A(n3680), .ZN(n4557) );
  NOR2_X1 U4488 ( .A1(n4557), .A2(n4317), .ZN(n3685) );
  OAI22_X1 U4489 ( .A1(n4209), .A2(n3683), .B1(n3711), .B2(n4369), .ZN(n3684)
         );
  AOI211_X1 U4490 ( .C1(n4488), .C2(n4209), .A(n3685), .B(n3684), .ZN(n3686)
         );
  OAI21_X1 U4491 ( .B1(n3687), .B2(n4382), .A(n3686), .ZN(U3277) );
  OAI21_X1 U4492 ( .B1(n2254), .B2(n3689), .A(n3688), .ZN(n4692) );
  INV_X1 U4493 ( .A(REG0_REG_10__SCAN_IN), .ZN(n3699) );
  NAND2_X1 U4494 ( .A1(n4022), .A2(n4027), .ZN(n3962) );
  XOR2_X1 U4495 ( .A(n3690), .B(n3962), .Z(n4694) );
  XNOR2_X1 U4496 ( .A(n3691), .B(n3962), .ZN(n3695) );
  AOI22_X1 U4497 ( .A1(n4079), .A2(n4411), .B1(n3692), .B2(n4477), .ZN(n3694)
         );
  NAND2_X1 U4498 ( .A1(n4077), .A2(n4478), .ZN(n3693) );
  OAI211_X1 U4499 ( .C1(n3695), .C2(n4312), .A(n3694), .B(n3693), .ZN(n3696)
         );
  AOI21_X1 U4500 ( .B1(n4694), .B2(n3697), .A(n3696), .ZN(n4697) );
  INV_X1 U4501 ( .A(n4697), .ZN(n3698) );
  AOI21_X1 U4502 ( .B1(n4756), .B2(n4694), .A(n3698), .ZN(n3701) );
  MUX2_X1 U4503 ( .A(n3699), .B(n3701), .S(n4759), .Z(n3700) );
  OAI21_X1 U4504 ( .B1(n4692), .B2(n4556), .A(n3700), .ZN(U3487) );
  INV_X1 U4505 ( .A(REG1_REG_10__SCAN_IN), .ZN(n3702) );
  MUX2_X1 U4506 ( .A(n3702), .B(n3701), .S(n4770), .Z(n3703) );
  OAI21_X1 U4507 ( .B1(n4692), .B2(n4491), .A(n3703), .ZN(U3528) );
  XOR2_X1 U4508 ( .A(n3706), .B(n3705), .Z(n3707) );
  XNOR2_X1 U4509 ( .A(n3704), .B(n3707), .ZN(n3713) );
  NOR2_X1 U4510 ( .A1(STATE_REG_SCAN_IN), .A2(n2602), .ZN(n4645) );
  AOI21_X1 U4511 ( .B1(n3905), .B2(n4076), .A(n4645), .ZN(n3710) );
  AOI22_X1 U4512 ( .A1(n4577), .A2(n4467), .B1(n3904), .B2(n3708), .ZN(n3709)
         );
  OAI211_X1 U4513 ( .C1(n4586), .C2(n3711), .A(n3710), .B(n3709), .ZN(n3712)
         );
  AOI21_X1 U4514 ( .B1(n3713), .B2(n4581), .A(n3712), .ZN(n3714) );
  INV_X1 U4515 ( .A(n3714), .ZN(U3231) );
  INV_X1 U4516 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3721) );
  AOI22_X1 U4517 ( .A1(n4075), .A2(n4478), .B1(n4477), .B2(n3715), .ZN(n3717)
         );
  NAND2_X1 U4518 ( .A1(n4077), .A2(n4411), .ZN(n3716) );
  NAND3_X1 U4519 ( .A1(n3718), .A2(n3717), .A3(n3716), .ZN(n3719) );
  AOI21_X1 U4520 ( .B1(n3720), .B2(n4745), .A(n3719), .ZN(n3723) );
  MUX2_X1 U4521 ( .A(n3721), .B(n3723), .S(n4759), .Z(n3722) );
  OAI21_X1 U4522 ( .B1(n3726), .B2(n4556), .A(n3722), .ZN(U3491) );
  INV_X1 U4523 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3724) );
  MUX2_X1 U4524 ( .A(n3724), .B(n3723), .S(n4770), .Z(n3725) );
  OAI21_X1 U4525 ( .B1(n4491), .B2(n3726), .A(n3725), .ZN(U3530) );
  NAND2_X1 U4526 ( .A1(n3636), .A2(n3727), .ZN(n3729) );
  AND2_X1 U4527 ( .A1(n3729), .A2(n3728), .ZN(n3732) );
  AOI21_X1 U4528 ( .B1(n3733), .B2(n3732), .A(n2273), .ZN(n3739) );
  INV_X1 U4529 ( .A(n3734), .ZN(n3921) );
  INV_X1 U4530 ( .A(n3735), .ZN(n3736) );
  AOI21_X1 U4531 ( .B1(n3921), .B2(n3949), .A(n3736), .ZN(n3737) );
  OAI22_X1 U4532 ( .A1(n3739), .A2(n3738), .B1(n4312), .B2(n3737), .ZN(n4483)
         );
  INV_X1 U4533 ( .A(n4483), .ZN(n3749) );
  INV_X1 U4534 ( .A(n3739), .ZN(n4485) );
  OAI21_X1 U4535 ( .B1(n3742), .B2(n3741), .A(n3740), .ZN(n4552) );
  OAI22_X1 U4536 ( .A1(n4209), .A2(n3743), .B1(n3755), .B2(n4369), .ZN(n3745)
         );
  INV_X1 U4537 ( .A(n4075), .ZN(n4482) );
  INV_X1 U4538 ( .A(n4479), .ZN(n4572) );
  OAI22_X1 U4539 ( .A1(n4291), .A2(n4482), .B1(n4572), .B2(n4293), .ZN(n3744)
         );
  AOI211_X1 U4540 ( .C1(n4476), .C2(n4215), .A(n3745), .B(n3744), .ZN(n3746)
         );
  OAI21_X1 U4541 ( .B1(n4552), .B2(n4317), .A(n3746), .ZN(n3747) );
  AOI21_X1 U4542 ( .B1(n4485), .B2(n4708), .A(n3747), .ZN(n3748) );
  OAI21_X1 U4543 ( .B1(n3749), .B2(n4713), .A(n3748), .ZN(U3276) );
  NAND2_X1 U4544 ( .A1(n2276), .A2(n3751), .ZN(n3752) );
  XNOR2_X1 U4545 ( .A(n3750), .B(n3752), .ZN(n3757) );
  AND2_X1 U4546 ( .A1(REG3_REG_14__SCAN_IN), .A2(U3149), .ZN(n4655) );
  AOI21_X1 U4547 ( .B1(n4577), .B2(n4479), .A(n4655), .ZN(n3754) );
  AOI22_X1 U4548 ( .A1(n3905), .A2(n4075), .B1(n3904), .B2(n4476), .ZN(n3753)
         );
  OAI211_X1 U4549 ( .C1(n4586), .C2(n3755), .A(n3754), .B(n3753), .ZN(n3756)
         );
  AOI21_X1 U4550 ( .B1(n3757), .B2(n4581), .A(n3756), .ZN(n3758) );
  INV_X1 U4551 ( .A(n3758), .ZN(U3212) );
  OAI22_X1 U4552 ( .A1(n4396), .A2(n2939), .B1(n2252), .B2(n3771), .ZN(n3769)
         );
  INV_X1 U4553 ( .A(n3764), .ZN(n3765) );
  OAI22_X1 U4554 ( .A1(n4396), .A2(n3765), .B1(n2939), .B2(n3771), .ZN(n3767)
         );
  XNOR2_X1 U4555 ( .A(n3767), .B(n3766), .ZN(n3768) );
  INV_X1 U4556 ( .A(n3780), .ZN(n3775) );
  OAI22_X1 U4557 ( .A1(n3781), .A2(n3875), .B1(n4574), .B2(n3771), .ZN(n3774)
         );
  INV_X1 U4558 ( .A(n4074), .ZN(n4170) );
  OAI22_X1 U4559 ( .A1(n4170), .A2(n4571), .B1(STATE_REG_SCAN_IN), .B2(n3772), 
        .ZN(n3773) );
  AOI211_X1 U4560 ( .C1(n3775), .C2(n3185), .A(n3774), .B(n3773), .ZN(n3776)
         );
  OAI21_X1 U4561 ( .B1(n3777), .B2(n3861), .A(n3776), .ZN(U3217) );
  INV_X1 U4562 ( .A(n3778), .ZN(n3788) );
  OAI22_X1 U4563 ( .A1(n3780), .A2(n4369), .B1(n3779), .B2(n4209), .ZN(n3783)
         );
  OAI22_X1 U4564 ( .A1(n4170), .A2(n4291), .B1(n3781), .B2(n4293), .ZN(n3782)
         );
  AOI211_X1 U4565 ( .C1(n3784), .C2(n4215), .A(n3783), .B(n3782), .ZN(n3785)
         );
  OAI21_X1 U4566 ( .B1(n3786), .B2(n4317), .A(n3785), .ZN(n3787) );
  AOI21_X1 U4567 ( .B1(n3788), .B2(n4209), .A(n3787), .ZN(n3789) );
  OAI21_X1 U4568 ( .B1(n3790), .B2(n4382), .A(n3789), .ZN(U3262) );
  INV_X1 U4569 ( .A(IR_REG_30__SCAN_IN), .ZN(n3792) );
  NAND3_X1 U4570 ( .A1(n3792), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3794) );
  INV_X1 U4571 ( .A(DATAI_31_), .ZN(n3793) );
  OAI22_X1 U4572 ( .A1(n3791), .A2(n3794), .B1(STATE_REG_SCAN_IN), .B2(n3793), 
        .ZN(U3321) );
  AOI21_X1 U4573 ( .B1(n3872), .B2(n3798), .A(n3797), .ZN(n3799) );
  NOR3_X1 U4574 ( .A1(n3800), .A2(n3799), .A3(n3861), .ZN(n3804) );
  AOI22_X1 U4575 ( .A1(n4233), .A2(n4577), .B1(n3945), .B2(n3904), .ZN(n3802)
         );
  AOI22_X1 U4576 ( .A1(n4430), .A2(n3905), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n3801) );
  OAI211_X1 U4577 ( .C1(n4586), .C2(n4239), .A(n3802), .B(n3801), .ZN(n3803)
         );
  OR2_X1 U4578 ( .A1(n3804), .A2(n3803), .ZN(U3213) );
  XNOR2_X1 U4579 ( .A(n2257), .B(n3805), .ZN(n3810) );
  AND2_X1 U4580 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4121) );
  AOI21_X1 U4581 ( .B1(n3905), .B2(n4455), .A(n4121), .ZN(n3808) );
  AOI22_X1 U4582 ( .A1(n4577), .A2(n4272), .B1(n3904), .B2(n3806), .ZN(n3807)
         );
  OAI211_X1 U4583 ( .C1(n4586), .C2(n4318), .A(n3808), .B(n3807), .ZN(n3809)
         );
  AOI21_X1 U4584 ( .B1(n3810), .B2(n4581), .A(n3809), .ZN(n3811) );
  INV_X1 U4585 ( .A(n3811), .ZN(U3216) );
  OAI21_X1 U4586 ( .B1(n3812), .B2(n3864), .A(n3863), .ZN(n3816) );
  XNOR2_X1 U4587 ( .A(n3814), .B(n3813), .ZN(n3815) );
  XNOR2_X1 U4588 ( .A(n3816), .B(n3815), .ZN(n3820) );
  AOI22_X1 U4589 ( .A1(n3905), .A2(n4272), .B1(REG3_REG_21__SCAN_IN), .B2(
        U3149), .ZN(n3818) );
  AOI22_X1 U4590 ( .A1(n4430), .A2(n4577), .B1(n3904), .B2(n4429), .ZN(n3817)
         );
  OAI211_X1 U4591 ( .C1(n4586), .C2(n4268), .A(n3818), .B(n3817), .ZN(n3819)
         );
  AOI21_X1 U4592 ( .B1(n3820), .B2(n4581), .A(n3819), .ZN(n3821) );
  INV_X1 U4593 ( .A(n3821), .ZN(U3220) );
  NAND2_X1 U4594 ( .A1(n2424), .A2(n3824), .ZN(n3825) );
  XNOR2_X1 U4595 ( .A(n3822), .B(n3825), .ZN(n3831) );
  OAI22_X1 U4596 ( .A1(n4193), .A2(n4571), .B1(STATE_REG_SCAN_IN), .B2(n3826), 
        .ZN(n3829) );
  OAI22_X1 U4597 ( .A1(n4157), .A2(n3875), .B1(n4574), .B2(n3827), .ZN(n3828)
         );
  AOI211_X1 U4598 ( .C1(n4185), .C2(n3185), .A(n3829), .B(n3828), .ZN(n3830)
         );
  OAI21_X1 U4599 ( .B1(n3831), .B2(n3861), .A(n3830), .ZN(U3222) );
  OAI211_X1 U4600 ( .C1(n3834), .C2(n3833), .A(n3832), .B(n4581), .ZN(n3841)
         );
  AOI21_X1 U4601 ( .B1(n3905), .B2(n4084), .A(n3835), .ZN(n3840) );
  AOI22_X1 U4602 ( .A1(n4577), .A2(n4082), .B1(n3904), .B2(n3836), .ZN(n3839)
         );
  OR2_X1 U4603 ( .A1(n4586), .A2(n3837), .ZN(n3838) );
  NAND4_X1 U4604 ( .A1(n3841), .A2(n3840), .A3(n3839), .A4(n3838), .ZN(U3224)
         );
  NOR2_X1 U4605 ( .A1(n3844), .A2(n2389), .ZN(n3845) );
  XNOR2_X1 U4606 ( .A(n3842), .B(n3845), .ZN(n3849) );
  NOR2_X1 U4607 ( .A1(STATE_REG_SCAN_IN), .A2(n2645), .ZN(n4682) );
  AOI21_X1 U4608 ( .B1(n3905), .B2(n4469), .A(n4682), .ZN(n3847) );
  AOI22_X1 U4609 ( .A1(n4577), .A2(n4455), .B1(n3904), .B2(n4454), .ZN(n3846)
         );
  OAI211_X1 U4610 ( .C1(n4586), .C2(n4352), .A(n3847), .B(n3846), .ZN(n3848)
         );
  AOI21_X1 U4611 ( .B1(n3849), .B2(n4581), .A(n3848), .ZN(n3850) );
  INV_X1 U4612 ( .A(n3850), .ZN(U3225) );
  INV_X1 U4613 ( .A(n3851), .ZN(n3854) );
  NOR2_X1 U4614 ( .A1(n3854), .A2(n3853), .ZN(n3856) );
  XNOR2_X1 U4615 ( .A(n3856), .B(n3855), .ZN(n3862) );
  AOI22_X1 U4616 ( .A1(n4412), .A2(n3905), .B1(REG3_REG_24__SCAN_IN), .B2(
        U3149), .ZN(n3857) );
  OAI21_X1 U4617 ( .B1(n4574), .B2(n4207), .A(n3857), .ZN(n3859) );
  NOR2_X1 U4618 ( .A1(n4586), .A2(n4210), .ZN(n3858) );
  AOI211_X1 U4619 ( .C1(n4577), .C2(n4211), .A(n3859), .B(n3858), .ZN(n3860)
         );
  OAI21_X1 U4620 ( .B1(n3862), .B2(n3861), .A(n3860), .ZN(U3226) );
  INV_X1 U4621 ( .A(n3863), .ZN(n3865) );
  NOR2_X1 U4622 ( .A1(n3865), .A2(n3864), .ZN(n3866) );
  XNOR2_X1 U4623 ( .A(n3812), .B(n3866), .ZN(n3870) );
  AOI22_X1 U4624 ( .A1(n3905), .A2(n4332), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n3868) );
  AOI22_X1 U4625 ( .A1(n4577), .A2(n4439), .B1(n3904), .B2(n4438), .ZN(n3867)
         );
  OAI211_X1 U4626 ( .C1(n4586), .C2(n4288), .A(n3868), .B(n3867), .ZN(n3869)
         );
  AOI21_X1 U4627 ( .B1(n3870), .B2(n4581), .A(n3869), .ZN(n3871) );
  INV_X1 U4628 ( .A(n3871), .ZN(U3230) );
  OAI21_X1 U4629 ( .B1(n3873), .B2(n2267), .A(n3872), .ZN(n3874) );
  NAND2_X1 U4630 ( .A1(n3874), .A2(n4581), .ZN(n3879) );
  NOR2_X1 U4631 ( .A1(n4294), .A2(n4571), .ZN(n3877) );
  OAI22_X1 U4632 ( .A1(n4212), .A2(n3875), .B1(n4574), .B2(n4256), .ZN(n3876)
         );
  AOI211_X1 U4633 ( .C1(REG3_REG_22__SCAN_IN), .C2(U3149), .A(n3877), .B(n3876), .ZN(n3878) );
  OAI211_X1 U4634 ( .C1(n4586), .C2(n4248), .A(n3879), .B(n3878), .ZN(U3232)
         );
  OAI21_X1 U4635 ( .B1(n3881), .B2(n3883), .A(n3880), .ZN(n3882) );
  OAI21_X1 U4636 ( .B1(n2260), .B2(n3883), .A(n3882), .ZN(n3887) );
  AOI22_X1 U4637 ( .A1(n3905), .A2(n4576), .B1(REG3_REG_18__SCAN_IN), .B2(
        U3149), .ZN(n3885) );
  AOI22_X1 U4638 ( .A1(n4577), .A2(n4332), .B1(n3904), .B2(n4331), .ZN(n3884)
         );
  OAI211_X1 U4639 ( .C1(n4586), .C2(n4337), .A(n3885), .B(n3884), .ZN(n3886)
         );
  AOI21_X1 U4640 ( .B1(n3887), .B2(n4581), .A(n3886), .ZN(n3888) );
  INV_X1 U4641 ( .A(n3888), .ZN(U3235) );
  NAND2_X1 U4642 ( .A1(n2268), .A2(n3889), .ZN(n3890) );
  XNOR2_X1 U4643 ( .A(n3891), .B(n3890), .ZN(n3898) );
  AOI22_X1 U4644 ( .A1(n4074), .A2(n4577), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3896) );
  NAND2_X1 U4645 ( .A1(n3185), .A2(n4178), .ZN(n3895) );
  NAND2_X1 U4646 ( .A1(n4211), .A2(n3905), .ZN(n3894) );
  NAND2_X1 U4647 ( .A1(n3904), .A2(n3892), .ZN(n3893) );
  NAND4_X1 U4648 ( .A1(n3896), .A2(n3895), .A3(n3894), .A4(n3893), .ZN(n3897)
         );
  AOI21_X1 U4649 ( .B1(n3898), .B2(n4581), .A(n3897), .ZN(n3899) );
  INV_X1 U4650 ( .A(n3899), .ZN(U3237) );
  INV_X1 U4651 ( .A(n3901), .ZN(n3902) );
  NOR2_X1 U4652 ( .A1(n3900), .A2(n3902), .ZN(n3903) );
  XNOR2_X1 U4653 ( .A(n3903), .B(n4578), .ZN(n3910) );
  AND2_X1 U4654 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4663) );
  AOI21_X1 U4655 ( .B1(n4577), .B2(n4469), .A(n4663), .ZN(n3907) );
  AOI22_X1 U4656 ( .A1(n3905), .A2(n4467), .B1(n3904), .B2(n4468), .ZN(n3906)
         );
  OAI211_X1 U4657 ( .C1(n4586), .C2(n3908), .A(n3907), .B(n3906), .ZN(n3909)
         );
  AOI21_X1 U4658 ( .B1(n3910), .B2(n4581), .A(n3909), .ZN(n3911) );
  INV_X1 U4659 ( .A(n3911), .ZN(U3238) );
  NAND2_X1 U4660 ( .A1(n2240), .A2(DATAI_31_), .ZN(n4128) );
  INV_X1 U4661 ( .A(n4128), .ZN(n4131) );
  NAND2_X1 U4662 ( .A1(n2240), .A2(DATAI_30_), .ZN(n3940) );
  AND2_X1 U4663 ( .A1(n4072), .A2(n3940), .ZN(n3977) );
  INV_X1 U4664 ( .A(REG2_REG_31__SCAN_IN), .ZN(n4133) );
  NAND2_X1 U4665 ( .A1(n2735), .A2(REG1_REG_31__SCAN_IN), .ZN(n3914) );
  NAND2_X1 U4666 ( .A1(n2715), .A2(REG0_REG_31__SCAN_IN), .ZN(n3913) );
  OAI211_X1 U4667 ( .C1(n3915), .C2(n4133), .A(n3914), .B(n3913), .ZN(n4130)
         );
  NOR2_X1 U4668 ( .A1(n4130), .A2(n4128), .ZN(n3976) );
  INV_X1 U4669 ( .A(n3946), .ZN(n3916) );
  NOR2_X1 U4670 ( .A1(n3951), .A2(n3916), .ZN(n4049) );
  INV_X1 U4671 ( .A(n4049), .ZN(n3930) );
  AND2_X1 U4672 ( .A1(n3917), .A2(n3920), .ZN(n4032) );
  NAND2_X1 U4673 ( .A1(n3919), .A2(n3918), .ZN(n4016) );
  AND2_X1 U4674 ( .A1(n4016), .A2(n3920), .ZN(n4031) );
  AOI21_X1 U4675 ( .B1(n3921), .B2(n4032), .A(n4031), .ZN(n3923) );
  INV_X1 U4676 ( .A(n4038), .ZN(n3922) );
  OAI21_X1 U4677 ( .B1(n3923), .B2(n3922), .A(n4034), .ZN(n3926) );
  INV_X1 U4678 ( .A(n3924), .ZN(n3925) );
  AOI21_X1 U4679 ( .B1(n3926), .B2(n4225), .A(n3925), .ZN(n3928) );
  OAI21_X1 U4680 ( .B1(n3928), .B2(n4043), .A(n3927), .ZN(n3929) );
  OAI221_X1 U4681 ( .B1(n3930), .B2(n4045), .C1(n3930), .C2(n3929), .A(n4053), 
        .ZN(n3932) );
  NAND2_X1 U4682 ( .A1(n4130), .A2(n4128), .ZN(n4057) );
  OR2_X1 U4683 ( .A1(n4072), .A2(n3940), .ZN(n3931) );
  AND2_X1 U4684 ( .A1(n4057), .A2(n3931), .ZN(n3983) );
  OAI21_X1 U4685 ( .B1(n4073), .B2(n4138), .A(n3983), .ZN(n3936) );
  INV_X1 U4686 ( .A(n4150), .ZN(n3939) );
  AOI21_X1 U4687 ( .B1(n4073), .B2(n4138), .A(n3933), .ZN(n3937) );
  NAND2_X1 U4688 ( .A1(n3937), .A2(n3974), .ZN(n4050) );
  OR2_X1 U4689 ( .A1(n3935), .A2(n3934), .ZN(n3938) );
  AOI21_X1 U4690 ( .B1(n3938), .B2(n3937), .A(n3936), .ZN(n4054) );
  OAI21_X1 U4691 ( .B1(n3939), .B2(n4050), .A(n4054), .ZN(n3942) );
  INV_X1 U4692 ( .A(n4130), .ZN(n3941) );
  INV_X1 U4693 ( .A(n3940), .ZN(n4389) );
  AOI22_X1 U4694 ( .A1(n3943), .A2(n3942), .B1(n3941), .B2(n4389), .ZN(n3944)
         );
  AOI211_X1 U4695 ( .C1(n4131), .C2(n3977), .A(n3976), .B(n3944), .ZN(n4064)
         );
  XNOR2_X1 U4696 ( .A(n4412), .B(n3945), .ZN(n4229) );
  XNOR2_X1 U4697 ( .A(n4332), .B(n4315), .ZN(n4300) );
  INV_X1 U4698 ( .A(n4300), .ZN(n4307) );
  NAND2_X1 U4699 ( .A1(n3947), .A2(n3946), .ZN(n4202) );
  NOR4_X1 U4700 ( .A1(n4202), .A2(n3949), .A3(n3948), .A4(n4732), .ZN(n3950)
         );
  NAND4_X1 U4701 ( .A1(n4150), .A2(n4229), .A3(n4307), .A4(n3950), .ZN(n3954)
         );
  INV_X1 U4702 ( .A(n3951), .ZN(n3952) );
  NAND2_X1 U4703 ( .A1(n3952), .A2(n4166), .ZN(n4188) );
  NOR3_X1 U4704 ( .A1(n3954), .A2(n3953), .A3(n4188), .ZN(n3989) );
  INV_X1 U4705 ( .A(n4041), .ZN(n3956) );
  INV_X1 U4706 ( .A(n4264), .ZN(n3959) );
  NOR4_X1 U4707 ( .A1(n3959), .A2(n3958), .A3(n3957), .A4(n2765), .ZN(n3973)
         );
  INV_X1 U4708 ( .A(n4222), .ZN(n3960) );
  NAND2_X1 U4709 ( .A1(n3960), .A2(n4302), .ZN(n4345) );
  NOR4_X1 U4710 ( .A1(n4345), .A2(n3963), .A3(n3962), .A4(n3961), .ZN(n3972)
         );
  NOR4_X1 U4711 ( .A1(n4252), .A2(n3965), .A3(n3964), .A4(n4373), .ZN(n3971)
         );
  INV_X1 U4712 ( .A(n3966), .ZN(n3969) );
  NOR4_X1 U4713 ( .A1(n3969), .A2(n3433), .A3(n4330), .A4(n3968), .ZN(n3970)
         );
  NAND4_X1 U4714 ( .A1(n3973), .A2(n3972), .A3(n3971), .A4(n3970), .ZN(n3987)
         );
  NAND2_X1 U4715 ( .A1(n3975), .A2(n3974), .ZN(n4168) );
  INV_X1 U4716 ( .A(n3976), .ZN(n3979) );
  INV_X1 U4717 ( .A(n3977), .ZN(n3978) );
  NAND2_X1 U4718 ( .A1(n3979), .A2(n3978), .ZN(n4058) );
  INV_X1 U4719 ( .A(n4058), .ZN(n3982) );
  NAND2_X1 U4720 ( .A1(n3981), .A2(n3980), .ZN(n4285) );
  NAND4_X1 U4721 ( .A1(n3984), .A2(n3983), .A3(n3982), .A4(n4285), .ZN(n3985)
         );
  NOR4_X1 U4722 ( .A1(n3987), .A2(n4168), .A3(n3986), .A4(n3985), .ZN(n3988)
         );
  NAND3_X1 U4723 ( .A1(n3989), .A2(n2336), .A3(n3988), .ZN(n3991) );
  NAND2_X1 U4724 ( .A1(n3991), .A2(n3990), .ZN(n4061) );
  OAI211_X1 U4725 ( .C1(n3994), .C2(n2757), .A(n3993), .B(n3992), .ZN(n3997)
         );
  NAND3_X1 U4726 ( .A1(n3997), .A2(n3996), .A3(n3995), .ZN(n4000) );
  NAND3_X1 U4727 ( .A1(n4000), .A2(n3999), .A3(n3998), .ZN(n4003) );
  NAND3_X1 U4728 ( .A1(n4003), .A2(n4002), .A3(n4001), .ZN(n4010) );
  NOR3_X1 U4729 ( .A1(n4017), .A2(n2325), .A3(n4005), .ZN(n4009) );
  INV_X1 U4730 ( .A(n4006), .ZN(n4008) );
  AOI211_X1 U4731 ( .C1(n4010), .C2(n4009), .A(n4008), .B(n4007), .ZN(n4015)
         );
  NAND2_X1 U4732 ( .A1(n4012), .A2(n4011), .ZN(n4019) );
  OAI211_X1 U4733 ( .C1(n4015), .C2(n4019), .A(n4014), .B(n4013), .ZN(n4025)
         );
  NOR2_X1 U4734 ( .A1(n4016), .A2(n4018), .ZN(n4024) );
  OR4_X1 U4735 ( .A1(n4020), .A2(n4019), .A3(n4018), .A4(n4017), .ZN(n4021) );
  AOI21_X1 U4736 ( .B1(n4022), .B2(n4021), .A(n4031), .ZN(n4023) );
  AOI21_X1 U4737 ( .B1(n4025), .B2(n4024), .A(n4023), .ZN(n4030) );
  INV_X1 U4738 ( .A(n4027), .ZN(n4029) );
  NOR4_X1 U4739 ( .A1(n4030), .A2(n2317), .A3(n4029), .A4(n4028), .ZN(n4036)
         );
  AOI21_X1 U4740 ( .B1(n4033), .B2(n4032), .A(n4031), .ZN(n4035) );
  OAI21_X1 U4741 ( .B1(n4036), .B2(n4035), .A(n4034), .ZN(n4039) );
  AOI21_X1 U4742 ( .B1(n4039), .B2(n4038), .A(n4037), .ZN(n4040) );
  INV_X1 U4743 ( .A(n4040), .ZN(n4042) );
  AOI211_X1 U4744 ( .C1(n4042), .C2(n4225), .A(n4041), .B(n4224), .ZN(n4044)
         );
  NOR2_X1 U4745 ( .A1(n4044), .A2(n4043), .ZN(n4047) );
  OAI21_X1 U4746 ( .B1(n4047), .B2(n4046), .A(n4045), .ZN(n4048) );
  NAND2_X1 U4747 ( .A1(n4049), .A2(n4048), .ZN(n4052) );
  AOI211_X1 U4748 ( .C1(n4053), .C2(n4052), .A(n4051), .B(n4050), .ZN(n4056)
         );
  INV_X1 U4749 ( .A(n4054), .ZN(n4055) );
  NOR2_X1 U4750 ( .A1(n4056), .A2(n4055), .ZN(n4059) );
  OAI21_X1 U4751 ( .B1(n4059), .B2(n4058), .A(n4057), .ZN(n4060) );
  MUX2_X1 U4752 ( .A(n4061), .B(n4060), .S(n2242), .Z(n4062) );
  OAI21_X1 U4753 ( .B1(n4064), .B2(n4063), .A(n4062), .ZN(n4065) );
  XNOR2_X1 U4754 ( .A(n4065), .B(n4123), .ZN(n4071) );
  NAND2_X1 U4755 ( .A1(n4067), .A2(n4066), .ZN(n4068) );
  OAI211_X1 U4756 ( .C1(n4561), .C2(n4070), .A(n4068), .B(B_REG_SCAN_IN), .ZN(
        n4069) );
  OAI21_X1 U4757 ( .B1(n4071), .B2(n4070), .A(n4069), .ZN(U3239) );
  MUX2_X1 U4758 ( .A(DATAO_REG_31__SCAN_IN), .B(n4130), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4759 ( .A(DATAO_REG_30__SCAN_IN), .B(n4072), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4760 ( .A(n4073), .B(DATAO_REG_29__SCAN_IN), .S(n4086), .Z(U3579)
         );
  MUX2_X1 U4761 ( .A(n4140), .B(DATAO_REG_28__SCAN_IN), .S(n4086), .Z(U3578)
         );
  MUX2_X1 U4762 ( .A(n4074), .B(DATAO_REG_27__SCAN_IN), .S(n4086), .Z(U3577)
         );
  MUX2_X1 U4763 ( .A(n4393), .B(DATAO_REG_26__SCAN_IN), .S(n4086), .Z(U3576)
         );
  MUX2_X1 U4764 ( .A(n4211), .B(DATAO_REG_25__SCAN_IN), .S(n4086), .Z(U3575)
         );
  MUX2_X1 U4765 ( .A(n4233), .B(DATAO_REG_24__SCAN_IN), .S(n4086), .Z(U3574)
         );
  MUX2_X1 U4766 ( .A(DATAO_REG_23__SCAN_IN), .B(n4412), .S(U4043), .Z(U3573)
         );
  MUX2_X1 U4767 ( .A(DATAO_REG_22__SCAN_IN), .B(n4430), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4768 ( .A(DATAO_REG_21__SCAN_IN), .B(n4439), .S(U4043), .Z(U3571)
         );
  MUX2_X1 U4769 ( .A(n4272), .B(DATAO_REG_20__SCAN_IN), .S(n4086), .Z(U3570)
         );
  MUX2_X1 U4770 ( .A(n4332), .B(DATAO_REG_19__SCAN_IN), .S(n4086), .Z(U3569)
         );
  MUX2_X1 U4771 ( .A(n4455), .B(DATAO_REG_18__SCAN_IN), .S(n4086), .Z(U3568)
         );
  MUX2_X1 U4772 ( .A(n4576), .B(DATAO_REG_17__SCAN_IN), .S(n4086), .Z(U3567)
         );
  MUX2_X1 U4773 ( .A(n4469), .B(DATAO_REG_16__SCAN_IN), .S(n4086), .Z(U3566)
         );
  MUX2_X1 U4774 ( .A(n4479), .B(DATAO_REG_15__SCAN_IN), .S(n4086), .Z(U3565)
         );
  MUX2_X1 U4775 ( .A(n4467), .B(DATAO_REG_14__SCAN_IN), .S(n4086), .Z(U3564)
         );
  MUX2_X1 U4776 ( .A(n4075), .B(DATAO_REG_13__SCAN_IN), .S(n4086), .Z(U3563)
         );
  MUX2_X1 U4777 ( .A(n4076), .B(DATAO_REG_12__SCAN_IN), .S(n4086), .Z(U3562)
         );
  MUX2_X1 U4778 ( .A(n4077), .B(DATAO_REG_11__SCAN_IN), .S(n4086), .Z(U3561)
         );
  MUX2_X1 U4779 ( .A(n4078), .B(DATAO_REG_10__SCAN_IN), .S(n4086), .Z(U3560)
         );
  MUX2_X1 U4780 ( .A(n4079), .B(DATAO_REG_9__SCAN_IN), .S(n4086), .Z(U3559) );
  MUX2_X1 U4781 ( .A(n4080), .B(DATAO_REG_8__SCAN_IN), .S(n4086), .Z(U3558) );
  MUX2_X1 U4782 ( .A(n4081), .B(DATAO_REG_7__SCAN_IN), .S(n4086), .Z(U3557) );
  MUX2_X1 U4783 ( .A(n4082), .B(DATAO_REG_6__SCAN_IN), .S(n4086), .Z(U3556) );
  MUX2_X1 U4784 ( .A(n4083), .B(DATAO_REG_5__SCAN_IN), .S(n4086), .Z(U3555) );
  MUX2_X1 U4785 ( .A(n4084), .B(DATAO_REG_4__SCAN_IN), .S(n4086), .Z(U3554) );
  MUX2_X1 U4786 ( .A(n4085), .B(DATAO_REG_3__SCAN_IN), .S(n4086), .Z(U3553) );
  MUX2_X1 U4787 ( .A(n2949), .B(DATAO_REG_2__SCAN_IN), .S(n4086), .Z(U3552) );
  MUX2_X1 U4788 ( .A(n2484), .B(DATAO_REG_1__SCAN_IN), .S(n4086), .Z(U3551) );
  MUX2_X1 U4789 ( .A(n2925), .B(DATAO_REG_0__SCAN_IN), .S(n4086), .Z(U3550) );
  OAI211_X1 U4790 ( .C1(n4089), .C2(n4088), .A(n4684), .B(n4087), .ZN(n4099)
         );
  INV_X1 U4791 ( .A(n4090), .ZN(n4095) );
  MUX2_X1 U4792 ( .A(n2834), .B(REG2_REG_1__SCAN_IN), .S(n4091), .Z(n4094) );
  INV_X1 U4793 ( .A(n4092), .ZN(n4093) );
  OAI211_X1 U4794 ( .C1(n4095), .C2(n4094), .A(n4640), .B(n4093), .ZN(n4098)
         );
  NAND2_X1 U4795 ( .A1(n4103), .A2(n4568), .ZN(n4097) );
  AOI22_X1 U4796 ( .A1(n4683), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n4096) );
  NAND4_X1 U4797 ( .A1(n4099), .A2(n4098), .A3(n4097), .A4(n4096), .ZN(U3241)
         );
  OAI211_X1 U4798 ( .C1(REG1_REG_3__SCAN_IN), .C2(n4101), .A(n4684), .B(n4100), 
        .ZN(n4110) );
  NAND2_X1 U4799 ( .A1(n4103), .A2(n4102), .ZN(n4109) );
  AOI22_X1 U4800 ( .A1(n4683), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n4108) );
  XNOR2_X1 U4801 ( .A(n4105), .B(n4104), .ZN(n4106) );
  NAND2_X1 U4802 ( .A1(n4640), .A2(n4106), .ZN(n4107) );
  NAND4_X1 U4803 ( .A1(n4110), .A2(n4109), .A3(n4108), .A4(n4107), .ZN(U3243)
         );
  MUX2_X1 U4804 ( .A(REG2_REG_19__SCAN_IN), .B(n4319), .S(n4563), .Z(n4114) );
  OAI21_X1 U4805 ( .B1(n4717), .B2(n4117), .A(n4116), .ZN(n4120) );
  INV_X1 U4806 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4118) );
  MUX2_X1 U4807 ( .A(n4118), .B(REG1_REG_19__SCAN_IN), .S(n4563), .Z(n4119) );
  XNOR2_X1 U4808 ( .A(n4120), .B(n4119), .ZN(n4125) );
  AOI21_X1 U4809 ( .B1(n4683), .B2(ADDR_REG_19__SCAN_IN), .A(n4121), .ZN(n4122) );
  OAI21_X1 U4810 ( .B1(n4689), .B2(n4123), .A(n4122), .ZN(n4124) );
  AOI21_X1 U4811 ( .B1(n4125), .B2(n4684), .A(n4124), .ZN(n4126) );
  OAI21_X1 U4812 ( .B1(n4127), .B2(n4677), .A(n4126), .ZN(U3259) );
  NAND2_X1 U4813 ( .A1(n4130), .A2(n4129), .ZN(n4387) );
  NAND2_X1 U4814 ( .A1(n4131), .A2(n4477), .ZN(n4132) );
  NAND2_X1 U4815 ( .A1(n4387), .A2(n4132), .ZN(n4492) );
  NOR2_X1 U4816 ( .A1(n4209), .A2(n4133), .ZN(n4134) );
  AOI21_X1 U4817 ( .B1(n4209), .B2(n4492), .A(n4134), .ZN(n4135) );
  OAI21_X1 U4818 ( .B1(n4495), .B2(n4317), .A(n4135), .ZN(U3260) );
  INV_X1 U4819 ( .A(n4136), .ZN(n4148) );
  OAI22_X1 U4820 ( .A1(n4356), .A2(n4138), .B1(n4137), .B2(n4209), .ZN(n4139)
         );
  AOI21_X1 U4821 ( .B1(n4140), .B2(n4350), .A(n4139), .ZN(n4147) );
  INV_X1 U4822 ( .A(n4141), .ZN(n4145) );
  OAI22_X1 U4823 ( .A1(n4143), .A2(n4317), .B1(n4142), .B2(n4369), .ZN(n4144)
         );
  OAI21_X1 U4824 ( .B1(n4145), .B2(n4144), .A(n4209), .ZN(n4146) );
  OAI211_X1 U4825 ( .C1(n4148), .C2(n4382), .A(n4147), .B(n4146), .ZN(U3354)
         );
  XOR2_X1 U4826 ( .A(n4150), .B(n4149), .Z(n4398) );
  INV_X1 U4827 ( .A(n4398), .ZN(n4164) );
  XNOR2_X1 U4828 ( .A(n2264), .B(n4150), .ZN(n4151) );
  NAND2_X1 U4829 ( .A1(n4151), .A2(n4375), .ZN(n4395) );
  INV_X1 U4830 ( .A(n4395), .ZN(n4162) );
  INV_X1 U4831 ( .A(n4152), .ZN(n4153) );
  OAI21_X1 U4832 ( .B1(n4175), .B2(n4154), .A(n4153), .ZN(n4502) );
  OAI22_X1 U4833 ( .A1(n4156), .A2(n4369), .B1(n4155), .B2(n4209), .ZN(n4159)
         );
  OAI22_X1 U4834 ( .A1(n4396), .A2(n4293), .B1(n4157), .B2(n4291), .ZN(n4158)
         );
  AOI211_X1 U4835 ( .C1(n4392), .C2(n4215), .A(n4159), .B(n4158), .ZN(n4160)
         );
  OAI21_X1 U4836 ( .B1(n4502), .B2(n4317), .A(n4160), .ZN(n4161) );
  AOI21_X1 U4837 ( .B1(n4162), .B2(n4209), .A(n4161), .ZN(n4163) );
  OAI21_X1 U4838 ( .B1(n4164), .B2(n4382), .A(n4163), .ZN(U3263) );
  XOR2_X1 U4839 ( .A(n4168), .B(n4165), .Z(n4402) );
  INV_X1 U4840 ( .A(n4402), .ZN(n4182) );
  NAND2_X1 U4841 ( .A1(n4167), .A2(n4166), .ZN(n4169) );
  XNOR2_X1 U4842 ( .A(n4169), .B(n4168), .ZN(n4173) );
  OAI22_X1 U4843 ( .A1(n4170), .A2(n4415), .B1(n4309), .B2(n4177), .ZN(n4171)
         );
  AOI21_X1 U4844 ( .B1(n4411), .B2(n4211), .A(n4171), .ZN(n4172) );
  OAI21_X1 U4845 ( .B1(n4173), .B2(n4312), .A(n4172), .ZN(n4401) );
  INV_X1 U4846 ( .A(n4174), .ZN(n4184) );
  INV_X1 U4847 ( .A(n4175), .ZN(n4176) );
  OAI21_X1 U4848 ( .B1(n4184), .B2(n4177), .A(n4176), .ZN(n4506) );
  AOI22_X1 U4849 ( .A1(n4178), .A2(n4705), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4713), .ZN(n4179) );
  OAI21_X1 U4850 ( .B1(n4506), .B2(n4317), .A(n4179), .ZN(n4180) );
  AOI21_X1 U4851 ( .B1(n4401), .B2(n4209), .A(n4180), .ZN(n4181) );
  OAI21_X1 U4852 ( .B1(n4182), .B2(n4382), .A(n4181), .ZN(U3264) );
  XOR2_X1 U4853 ( .A(n4188), .B(n4183), .Z(n4406) );
  AOI21_X1 U4854 ( .B1(n4190), .B2(n4206), .A(n4184), .ZN(n4510) );
  INV_X1 U4855 ( .A(n4185), .ZN(n4187) );
  OAI22_X1 U4856 ( .A1(n4187), .A2(n4369), .B1(n4186), .B2(n4209), .ZN(n4197)
         );
  XNOR2_X1 U4857 ( .A(n4189), .B(n4188), .ZN(n4195) );
  NAND2_X1 U4858 ( .A1(n4393), .A2(n4478), .ZN(n4192) );
  NAND2_X1 U4859 ( .A1(n4190), .A2(n4477), .ZN(n4191) );
  OAI211_X1 U4860 ( .C1(n4193), .C2(n4481), .A(n4192), .B(n4191), .ZN(n4194)
         );
  AOI21_X1 U4861 ( .B1(n4195), .B2(n4375), .A(n4194), .ZN(n4405) );
  NOR2_X1 U4862 ( .A1(n4405), .A2(n4713), .ZN(n4196) );
  AOI211_X1 U4863 ( .C1(n4510), .C2(n4707), .A(n4197), .B(n4196), .ZN(n4198)
         );
  OAI21_X1 U4864 ( .B1(n4406), .B2(n4382), .A(n4198), .ZN(U3265) );
  XNOR2_X1 U4865 ( .A(n4199), .B(n4202), .ZN(n4418) );
  INV_X1 U4866 ( .A(n4418), .ZN(n4220) );
  NAND2_X1 U4867 ( .A1(n4201), .A2(n4200), .ZN(n4204) );
  INV_X1 U4868 ( .A(n4202), .ZN(n4203) );
  XNOR2_X1 U4869 ( .A(n4204), .B(n4203), .ZN(n4205) );
  NAND2_X1 U4870 ( .A1(n4205), .A2(n4375), .ZN(n4414) );
  INV_X1 U4871 ( .A(n4414), .ZN(n4218) );
  OAI21_X1 U4872 ( .B1(n4238), .B2(n4207), .A(n4206), .ZN(n4515) );
  OAI22_X1 U4873 ( .A1(n4210), .A2(n4369), .B1(n4209), .B2(n4208), .ZN(n4214)
         );
  INV_X1 U4874 ( .A(n4211), .ZN(n4416) );
  OAI22_X1 U4875 ( .A1(n4416), .A2(n4293), .B1(n4212), .B2(n4291), .ZN(n4213)
         );
  AOI211_X1 U4876 ( .C1(n4410), .C2(n4215), .A(n4214), .B(n4213), .ZN(n4216)
         );
  OAI21_X1 U4877 ( .B1(n4515), .B2(n4317), .A(n4216), .ZN(n4217) );
  AOI21_X1 U4878 ( .B1(n4218), .B2(n4209), .A(n4217), .ZN(n4219) );
  OAI21_X1 U4879 ( .B1(n4220), .B2(n4382), .A(n4219), .ZN(U3266) );
  XNOR2_X1 U4880 ( .A(n4221), .B(n4229), .ZN(n4422) );
  INV_X1 U4881 ( .A(n4422), .ZN(n4244) );
  AOI21_X1 U4882 ( .B1(n4280), .B2(n4225), .A(n4224), .ZN(n4261) );
  INV_X1 U4883 ( .A(n4226), .ZN(n4227) );
  AOI21_X1 U4884 ( .B1(n4261), .B2(n4264), .A(n4227), .ZN(n4253) );
  OAI21_X1 U4885 ( .B1(n4253), .B2(n4252), .A(n4228), .ZN(n4231) );
  INV_X1 U4886 ( .A(n4229), .ZN(n4230) );
  XNOR2_X1 U4887 ( .A(n4231), .B(n4230), .ZN(n4235) );
  OAI22_X1 U4888 ( .A1(n4273), .A2(n4481), .B1(n4309), .B2(n4236), .ZN(n4232)
         );
  AOI21_X1 U4889 ( .B1(n4233), .B2(n4478), .A(n4232), .ZN(n4234) );
  OAI21_X1 U4890 ( .B1(n4235), .B2(n4312), .A(n4234), .ZN(n4421) );
  NOR2_X1 U4891 ( .A1(n2245), .A2(n4236), .ZN(n4237) );
  OR2_X1 U4892 ( .A1(n4238), .A2(n4237), .ZN(n4519) );
  NOR2_X1 U4893 ( .A1(n4519), .A2(n4317), .ZN(n4242) );
  OAI22_X1 U4894 ( .A1(n4209), .A2(n4240), .B1(n4239), .B2(n4369), .ZN(n4241)
         );
  AOI211_X1 U4895 ( .C1(n4421), .C2(n4209), .A(n4242), .B(n4241), .ZN(n4243)
         );
  OAI21_X1 U4896 ( .B1(n4244), .B2(n4382), .A(n4243), .ZN(U3267) );
  OAI21_X1 U4897 ( .B1(n4246), .B2(n4252), .A(n4245), .ZN(n4426) );
  NOR2_X1 U4898 ( .A1(n4265), .A2(n4256), .ZN(n4247) );
  OR2_X1 U4899 ( .A1(n2245), .A2(n4247), .ZN(n4523) );
  INV_X1 U4900 ( .A(n4523), .ZN(n4251) );
  OAI22_X1 U4901 ( .A1(n4209), .A2(n4249), .B1(n4248), .B2(n4369), .ZN(n4250)
         );
  AOI21_X1 U4902 ( .B1(n4251), .B2(n4707), .A(n4250), .ZN(n4260) );
  XNOR2_X1 U4903 ( .A(n4253), .B(n4252), .ZN(n4258) );
  NAND2_X1 U4904 ( .A1(n4412), .A2(n4478), .ZN(n4255) );
  NAND2_X1 U4905 ( .A1(n4439), .A2(n4411), .ZN(n4254) );
  OAI211_X1 U4906 ( .C1(n4309), .C2(n4256), .A(n4255), .B(n4254), .ZN(n4257)
         );
  AOI21_X1 U4907 ( .B1(n4258), .B2(n4375), .A(n4257), .ZN(n4425) );
  OR2_X1 U4908 ( .A1(n4425), .A2(n4713), .ZN(n4259) );
  OAI211_X1 U4909 ( .C1(n4426), .C2(n4382), .A(n4260), .B(n4259), .ZN(U3268)
         );
  XNOR2_X1 U4910 ( .A(n4261), .B(n4264), .ZN(n4262) );
  NAND2_X1 U4911 ( .A1(n4262), .A2(n4375), .ZN(n4432) );
  XOR2_X1 U4912 ( .A(n4264), .B(n4263), .Z(n4435) );
  NAND2_X1 U4913 ( .A1(n4435), .A2(n4347), .ZN(n4278) );
  INV_X1 U4914 ( .A(n4287), .ZN(n4267) );
  INV_X1 U4915 ( .A(n4265), .ZN(n4266) );
  OAI21_X1 U4916 ( .B1(n4267), .B2(n4271), .A(n4266), .ZN(n4527) );
  INV_X1 U4917 ( .A(n4527), .ZN(n4276) );
  INV_X1 U4918 ( .A(n4268), .ZN(n4269) );
  AOI22_X1 U4919 ( .A1(n4713), .A2(REG2_REG_21__SCAN_IN), .B1(n4269), .B2(
        n4705), .ZN(n4270) );
  OAI21_X1 U4920 ( .B1(n4271), .B2(n4356), .A(n4270), .ZN(n4275) );
  INV_X1 U4921 ( .A(n4272), .ZN(n4433) );
  OAI22_X1 U4922 ( .A1(n4291), .A2(n4433), .B1(n4273), .B2(n4293), .ZN(n4274)
         );
  AOI211_X1 U4923 ( .C1(n4276), .C2(n4707), .A(n4275), .B(n4274), .ZN(n4277)
         );
  OAI211_X1 U4924 ( .C1(n4713), .C2(n4432), .A(n4278), .B(n4277), .ZN(U3269)
         );
  NAND2_X1 U4925 ( .A1(n4280), .A2(n4279), .ZN(n4281) );
  XNOR2_X1 U4926 ( .A(n4281), .B(n4285), .ZN(n4282) );
  NAND2_X1 U4927 ( .A1(n4282), .A2(n4375), .ZN(n4441) );
  AOI21_X1 U4928 ( .B1(n4301), .B2(n4284), .A(n4283), .ZN(n4286) );
  XNOR2_X1 U4929 ( .A(n4286), .B(n4285), .ZN(n4444) );
  NAND2_X1 U4930 ( .A1(n4444), .A2(n4347), .ZN(n4299) );
  OAI21_X1 U4931 ( .B1(n2294), .B2(n4292), .A(n4287), .ZN(n4531) );
  INV_X1 U4932 ( .A(n4531), .ZN(n4297) );
  INV_X1 U4933 ( .A(n4332), .ZN(n4442) );
  INV_X1 U4934 ( .A(n4288), .ZN(n4289) );
  AOI22_X1 U4935 ( .A1(n4713), .A2(REG2_REG_20__SCAN_IN), .B1(n4289), .B2(
        n4705), .ZN(n4290) );
  OAI21_X1 U4936 ( .B1(n4291), .B2(n4442), .A(n4290), .ZN(n4296) );
  OAI22_X1 U4937 ( .A1(n4294), .A2(n4293), .B1(n4356), .B2(n4292), .ZN(n4295)
         );
  AOI211_X1 U4938 ( .C1(n4297), .C2(n4707), .A(n4296), .B(n4295), .ZN(n4298)
         );
  OAI211_X1 U4939 ( .C1(n4713), .C2(n4441), .A(n4299), .B(n4298), .ZN(U3270)
         );
  XNOR2_X1 U4940 ( .A(n4301), .B(n4300), .ZN(n4448) );
  INV_X1 U4941 ( .A(n4448), .ZN(n4323) );
  NAND2_X1 U4942 ( .A1(n4303), .A2(n4302), .ZN(n4329) );
  INV_X1 U4943 ( .A(n4304), .ZN(n4306) );
  OAI21_X1 U4944 ( .B1(n4329), .B2(n4306), .A(n4305), .ZN(n4308) );
  XNOR2_X1 U4945 ( .A(n4308), .B(n4307), .ZN(n4313) );
  OAI22_X1 U4946 ( .A1(n4433), .A2(n4415), .B1(n4315), .B2(n4309), .ZN(n4310)
         );
  AOI21_X1 U4947 ( .B1(n4411), .B2(n4455), .A(n4310), .ZN(n4311) );
  OAI21_X1 U4948 ( .B1(n4313), .B2(n4312), .A(n4311), .ZN(n4447) );
  INV_X1 U4949 ( .A(n4327), .ZN(n4316) );
  OAI21_X1 U4950 ( .B1(n4316), .B2(n4315), .A(n4314), .ZN(n4535) );
  NOR2_X1 U4951 ( .A1(n4535), .A2(n4317), .ZN(n4321) );
  OAI22_X1 U4952 ( .A1(n4209), .A2(n4319), .B1(n4318), .B2(n4369), .ZN(n4320)
         );
  AOI211_X1 U4953 ( .C1(n4447), .C2(n4209), .A(n4321), .B(n4320), .ZN(n4322)
         );
  OAI21_X1 U4954 ( .B1(n4323), .B2(n4382), .A(n4322), .ZN(U3271) );
  OAI21_X1 U4955 ( .B1(n4324), .B2(n4330), .A(n4325), .ZN(n4326) );
  INV_X1 U4956 ( .A(n4326), .ZN(n4453) );
  OAI211_X1 U4957 ( .C1(n4348), .C2(n4328), .A(n4738), .B(n4327), .ZN(n4450)
         );
  XOR2_X1 U4958 ( .A(n4330), .B(n4329), .Z(n4336) );
  AOI22_X1 U4959 ( .A1(n4332), .A2(n4478), .B1(n4331), .B2(n4477), .ZN(n4333)
         );
  OAI21_X1 U4960 ( .B1(n4334), .B2(n4481), .A(n4333), .ZN(n4335) );
  AOI21_X1 U4961 ( .B1(n4336), .B2(n4375), .A(n4335), .ZN(n4451) );
  OAI21_X1 U4962 ( .B1(n4563), .B2(n4450), .A(n4451), .ZN(n4340) );
  OAI22_X1 U4963 ( .A1(n4209), .A2(n4338), .B1(n4337), .B2(n4369), .ZN(n4339)
         );
  AOI21_X1 U4964 ( .B1(n4340), .B2(n4209), .A(n4339), .ZN(n4341) );
  OAI21_X1 U4965 ( .B1(n4453), .B2(n4382), .A(n4341), .ZN(U3272) );
  XNOR2_X1 U4966 ( .A(n4342), .B(n4345), .ZN(n4343) );
  NAND2_X1 U4967 ( .A1(n4343), .A2(n4375), .ZN(n4457) );
  INV_X1 U4968 ( .A(n4344), .ZN(n4346) );
  XNOR2_X1 U4969 ( .A(n4346), .B(n4345), .ZN(n4460) );
  NAND2_X1 U4970 ( .A1(n4460), .A2(n4347), .ZN(n4361) );
  INV_X1 U4971 ( .A(n4348), .ZN(n4349) );
  OAI21_X1 U4972 ( .B1(n4367), .B2(n4357), .A(n4349), .ZN(n4540) );
  INV_X1 U4973 ( .A(n4540), .ZN(n4359) );
  AOI22_X1 U4974 ( .A1(n4351), .A2(n4455), .B1(n4350), .B2(n4469), .ZN(n4355)
         );
  INV_X1 U4975 ( .A(n4352), .ZN(n4353) );
  AOI22_X1 U4976 ( .A1(n4713), .A2(REG2_REG_17__SCAN_IN), .B1(n4353), .B2(
        n4705), .ZN(n4354) );
  OAI211_X1 U4977 ( .C1(n4357), .C2(n4356), .A(n4355), .B(n4354), .ZN(n4358)
         );
  AOI21_X1 U4978 ( .B1(n4359), .B2(n4707), .A(n4358), .ZN(n4360) );
  OAI211_X1 U4979 ( .C1(n4713), .C2(n4457), .A(n4361), .B(n4360), .ZN(U3273)
         );
  NOR2_X1 U4980 ( .A1(n4363), .A2(n4373), .ZN(n4364) );
  OR2_X1 U4981 ( .A1(n4365), .A2(n4364), .ZN(n4462) );
  AND2_X1 U4982 ( .A1(n4366), .A2(n4377), .ZN(n4368) );
  OR2_X1 U4983 ( .A1(n4368), .A2(n4367), .ZN(n4544) );
  INV_X1 U4984 ( .A(n4544), .ZN(n4372) );
  OAI22_X1 U4985 ( .A1(n4209), .A2(n4370), .B1(n4585), .B2(n4369), .ZN(n4371)
         );
  AOI21_X1 U4986 ( .B1(n4372), .B2(n4707), .A(n4371), .ZN(n4381) );
  XNOR2_X1 U4987 ( .A(n4374), .B(n4373), .ZN(n4376) );
  NAND2_X1 U4988 ( .A1(n4376), .A2(n4375), .ZN(n4379) );
  AOI22_X1 U4989 ( .A1(n4576), .A2(n4478), .B1(n4477), .B2(n4377), .ZN(n4378)
         );
  OAI211_X1 U4990 ( .C1(n4572), .C2(n4481), .A(n4379), .B(n4378), .ZN(n4463)
         );
  NAND2_X1 U4991 ( .A1(n4463), .A2(n4209), .ZN(n4380) );
  OAI211_X1 U4992 ( .C1(n4462), .C2(n4382), .A(n4381), .B(n4380), .ZN(U3274)
         );
  INV_X1 U4993 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4385) );
  NAND2_X1 U4994 ( .A1(n4492), .A2(n4770), .ZN(n4383) );
  OAI211_X1 U4995 ( .C1(n4770), .C2(n4385), .A(n4384), .B(n4383), .ZN(U3549)
         );
  AOI21_X1 U4996 ( .B1(n4389), .B2(n2256), .A(n2243), .ZN(n4587) );
  INV_X1 U4997 ( .A(n4587), .ZN(n4498) );
  INV_X1 U4998 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4390) );
  INV_X1 U4999 ( .A(n4387), .ZN(n4388) );
  AOI21_X1 U5000 ( .B1(n4389), .B2(n4477), .A(n4388), .ZN(n4589) );
  MUX2_X1 U5001 ( .A(n4390), .B(n4589), .S(n4770), .Z(n4391) );
  OAI21_X1 U5002 ( .B1(n4498), .B2(n4491), .A(n4391), .ZN(U3548) );
  INV_X1 U5003 ( .A(REG1_REG_27__SCAN_IN), .ZN(n4399) );
  AOI22_X1 U5004 ( .A1(n4393), .A2(n4411), .B1(n4392), .B2(n4477), .ZN(n4394)
         );
  OAI211_X1 U5005 ( .C1(n4396), .C2(n4415), .A(n4395), .B(n4394), .ZN(n4397)
         );
  AOI21_X1 U5006 ( .B1(n4398), .B2(n4745), .A(n4397), .ZN(n4499) );
  MUX2_X1 U5007 ( .A(n4399), .B(n4499), .S(n4770), .Z(n4400) );
  OAI21_X1 U5008 ( .B1(n4491), .B2(n4502), .A(n4400), .ZN(U3545) );
  INV_X1 U5009 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4403) );
  AOI21_X1 U5010 ( .B1(n4402), .B2(n4745), .A(n4401), .ZN(n4503) );
  MUX2_X1 U5011 ( .A(n4403), .B(n4503), .S(n4770), .Z(n4404) );
  OAI21_X1 U5012 ( .B1(n4491), .B2(n4506), .A(n4404), .ZN(U3544) );
  OAI21_X1 U5013 ( .B1(n4406), .B2(n4452), .A(n4405), .ZN(n4507) );
  MUX2_X1 U5014 ( .A(REG1_REG_25__SCAN_IN), .B(n4507), .S(n4770), .Z(n4407) );
  AOI21_X1 U5015 ( .B1(n4408), .B2(n4510), .A(n4407), .ZN(n4409) );
  INV_X1 U5016 ( .A(n4409), .ZN(U3543) );
  INV_X1 U5017 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4419) );
  AOI22_X1 U5018 ( .A1(n4412), .A2(n4411), .B1(n4477), .B2(n4410), .ZN(n4413)
         );
  OAI211_X1 U5019 ( .C1(n4416), .C2(n4415), .A(n4414), .B(n4413), .ZN(n4417)
         );
  AOI21_X1 U5020 ( .B1(n4418), .B2(n4745), .A(n4417), .ZN(n4512) );
  MUX2_X1 U5021 ( .A(n4419), .B(n4512), .S(n4770), .Z(n4420) );
  OAI21_X1 U5022 ( .B1(n4491), .B2(n4515), .A(n4420), .ZN(U3542) );
  INV_X1 U5023 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4423) );
  AOI21_X1 U5024 ( .B1(n4422), .B2(n4745), .A(n4421), .ZN(n4516) );
  MUX2_X1 U5025 ( .A(n4423), .B(n4516), .S(n4770), .Z(n4424) );
  OAI21_X1 U5026 ( .B1(n4491), .B2(n4519), .A(n4424), .ZN(U3541) );
  OAI21_X1 U5027 ( .B1(n4426), .B2(n4452), .A(n4425), .ZN(n4520) );
  MUX2_X1 U5028 ( .A(REG1_REG_22__SCAN_IN), .B(n4520), .S(n4770), .Z(n4427) );
  INV_X1 U5029 ( .A(n4427), .ZN(n4428) );
  OAI21_X1 U5030 ( .B1(n4491), .B2(n4523), .A(n4428), .ZN(U3540) );
  INV_X1 U5031 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4436) );
  AOI22_X1 U5032 ( .A1(n4430), .A2(n4478), .B1(n4477), .B2(n4429), .ZN(n4431)
         );
  OAI211_X1 U5033 ( .C1(n4433), .C2(n4481), .A(n4432), .B(n4431), .ZN(n4434)
         );
  AOI21_X1 U5034 ( .B1(n4435), .B2(n4745), .A(n4434), .ZN(n4524) );
  MUX2_X1 U5035 ( .A(n4436), .B(n4524), .S(n4770), .Z(n4437) );
  OAI21_X1 U5036 ( .B1(n4491), .B2(n4527), .A(n4437), .ZN(U3539) );
  INV_X1 U5037 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4445) );
  AOI22_X1 U5038 ( .A1(n4439), .A2(n4478), .B1(n4438), .B2(n4477), .ZN(n4440)
         );
  OAI211_X1 U5039 ( .C1(n4442), .C2(n4481), .A(n4441), .B(n4440), .ZN(n4443)
         );
  AOI21_X1 U5040 ( .B1(n4444), .B2(n4745), .A(n4443), .ZN(n4528) );
  MUX2_X1 U5041 ( .A(n4445), .B(n4528), .S(n4770), .Z(n4446) );
  OAI21_X1 U5042 ( .B1(n4491), .B2(n4531), .A(n4446), .ZN(U3538) );
  AOI21_X1 U5043 ( .B1(n4448), .B2(n4745), .A(n4447), .ZN(n4532) );
  MUX2_X1 U5044 ( .A(n4118), .B(n4532), .S(n4770), .Z(n4449) );
  OAI21_X1 U5045 ( .B1(n4491), .B2(n4535), .A(n4449), .ZN(U3537) );
  OAI211_X1 U5046 ( .C1(n4453), .C2(n4452), .A(n4451), .B(n4450), .ZN(n4536)
         );
  MUX2_X1 U5047 ( .A(REG1_REG_18__SCAN_IN), .B(n4536), .S(n4770), .Z(U3536) );
  INV_X1 U5048 ( .A(n4469), .ZN(n4458) );
  AOI22_X1 U5049 ( .A1(n4455), .A2(n4478), .B1(n4477), .B2(n4454), .ZN(n4456)
         );
  OAI211_X1 U5050 ( .C1(n4458), .C2(n4481), .A(n4457), .B(n4456), .ZN(n4459)
         );
  AOI21_X1 U5051 ( .B1(n4460), .B2(n4745), .A(n4459), .ZN(n4537) );
  MUX2_X1 U5052 ( .A(n2900), .B(n4537), .S(n4770), .Z(n4461) );
  OAI21_X1 U5053 ( .B1(n4491), .B2(n4540), .A(n4461), .ZN(U3535) );
  INV_X1 U5054 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4465) );
  INV_X1 U5055 ( .A(n4462), .ZN(n4464) );
  AOI21_X1 U5056 ( .B1(n4464), .B2(n4745), .A(n4463), .ZN(n4541) );
  MUX2_X1 U5057 ( .A(n4465), .B(n4541), .S(n4770), .Z(n4466) );
  OAI21_X1 U5058 ( .B1(n4491), .B2(n4544), .A(n4466), .ZN(U3534) );
  INV_X1 U5059 ( .A(n4467), .ZN(n4472) );
  AOI22_X1 U5060 ( .A1(n4469), .A2(n4478), .B1(n4477), .B2(n4468), .ZN(n4470)
         );
  OAI211_X1 U5061 ( .C1(n4472), .C2(n4481), .A(n4471), .B(n4470), .ZN(n4473)
         );
  AOI21_X1 U5062 ( .B1(n4474), .B2(n4745), .A(n4473), .ZN(n4545) );
  MUX2_X1 U5063 ( .A(n2869), .B(n4545), .S(n4770), .Z(n4475) );
  OAI21_X1 U5064 ( .B1(n4491), .B2(n4548), .A(n4475), .ZN(U3533) );
  INV_X1 U5065 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4486) );
  AOI22_X1 U5066 ( .A1(n4479), .A2(n4478), .B1(n4477), .B2(n4476), .ZN(n4480)
         );
  OAI21_X1 U5067 ( .B1(n4482), .B2(n4481), .A(n4480), .ZN(n4484) );
  AOI211_X1 U5068 ( .C1(n4756), .C2(n4485), .A(n4484), .B(n4483), .ZN(n4549)
         );
  MUX2_X1 U5069 ( .A(n4486), .B(n4549), .S(n4770), .Z(n4487) );
  OAI21_X1 U5070 ( .B1(n4491), .B2(n4552), .A(n4487), .ZN(U3532) );
  AOI21_X1 U5071 ( .B1(n4489), .B2(n4745), .A(n4488), .ZN(n4553) );
  MUX2_X1 U5072 ( .A(n2871), .B(n4553), .S(n4770), .Z(n4490) );
  OAI21_X1 U5073 ( .B1(n4491), .B2(n4557), .A(n4490), .ZN(U3531) );
  NAND2_X1 U5074 ( .A1(n4492), .A2(n4759), .ZN(n4494) );
  NAND2_X1 U5075 ( .A1(n4757), .A2(REG0_REG_31__SCAN_IN), .ZN(n4493) );
  OAI211_X1 U5076 ( .C1(n4495), .C2(n4556), .A(n4494), .B(n4493), .ZN(U3517)
         );
  INV_X1 U5077 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4496) );
  MUX2_X1 U5078 ( .A(n4496), .B(n4589), .S(n4759), .Z(n4497) );
  OAI21_X1 U5079 ( .B1(n4498), .B2(n4556), .A(n4497), .ZN(U3516) );
  INV_X1 U5080 ( .A(REG0_REG_27__SCAN_IN), .ZN(n4500) );
  MUX2_X1 U5081 ( .A(n4500), .B(n4499), .S(n4759), .Z(n4501) );
  OAI21_X1 U5082 ( .B1(n4502), .B2(n4556), .A(n4501), .ZN(U3513) );
  INV_X1 U5083 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4504) );
  MUX2_X1 U5084 ( .A(n4504), .B(n4503), .S(n4759), .Z(n4505) );
  OAI21_X1 U5085 ( .B1(n4506), .B2(n4556), .A(n4505), .ZN(U3512) );
  MUX2_X1 U5086 ( .A(REG0_REG_25__SCAN_IN), .B(n4507), .S(n4759), .Z(n4508) );
  AOI21_X1 U5087 ( .B1(n4510), .B2(n4509), .A(n4508), .ZN(n4511) );
  INV_X1 U5088 ( .A(n4511), .ZN(U3511) );
  INV_X1 U5089 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4513) );
  MUX2_X1 U5090 ( .A(n4513), .B(n4512), .S(n4759), .Z(n4514) );
  OAI21_X1 U5091 ( .B1(n4515), .B2(n4556), .A(n4514), .ZN(U3510) );
  INV_X1 U5092 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4517) );
  MUX2_X1 U5093 ( .A(n4517), .B(n4516), .S(n4759), .Z(n4518) );
  OAI21_X1 U5094 ( .B1(n4519), .B2(n4556), .A(n4518), .ZN(U3509) );
  MUX2_X1 U5095 ( .A(REG0_REG_22__SCAN_IN), .B(n4520), .S(n4759), .Z(n4521) );
  INV_X1 U5096 ( .A(n4521), .ZN(n4522) );
  OAI21_X1 U5097 ( .B1(n4523), .B2(n4556), .A(n4522), .ZN(U3508) );
  INV_X1 U5098 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4525) );
  MUX2_X1 U5099 ( .A(n4525), .B(n4524), .S(n4759), .Z(n4526) );
  OAI21_X1 U5100 ( .B1(n4527), .B2(n4556), .A(n4526), .ZN(U3507) );
  INV_X1 U5101 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4529) );
  MUX2_X1 U5102 ( .A(n4529), .B(n4528), .S(n4759), .Z(n4530) );
  OAI21_X1 U5103 ( .B1(n4531), .B2(n4556), .A(n4530), .ZN(U3506) );
  INV_X1 U5104 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4533) );
  MUX2_X1 U5105 ( .A(n4533), .B(n4532), .S(n4759), .Z(n4534) );
  OAI21_X1 U5106 ( .B1(n4535), .B2(n4556), .A(n4534), .ZN(U3505) );
  MUX2_X1 U5107 ( .A(REG0_REG_18__SCAN_IN), .B(n4536), .S(n4759), .Z(U3503) );
  INV_X1 U5108 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4538) );
  MUX2_X1 U5109 ( .A(n4538), .B(n4537), .S(n4759), .Z(n4539) );
  OAI21_X1 U5110 ( .B1(n4540), .B2(n4556), .A(n4539), .ZN(U3501) );
  INV_X1 U5111 ( .A(REG0_REG_16__SCAN_IN), .ZN(n4542) );
  MUX2_X1 U5112 ( .A(n4542), .B(n4541), .S(n4759), .Z(n4543) );
  OAI21_X1 U5113 ( .B1(n4544), .B2(n4556), .A(n4543), .ZN(U3499) );
  INV_X1 U5114 ( .A(REG0_REG_15__SCAN_IN), .ZN(n4546) );
  MUX2_X1 U5115 ( .A(n4546), .B(n4545), .S(n4759), .Z(n4547) );
  OAI21_X1 U5116 ( .B1(n4548), .B2(n4556), .A(n4547), .ZN(U3497) );
  INV_X1 U5117 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4550) );
  MUX2_X1 U5118 ( .A(n4550), .B(n4549), .S(n4759), .Z(n4551) );
  OAI21_X1 U5119 ( .B1(n4552), .B2(n4556), .A(n4551), .ZN(U3495) );
  INV_X1 U5120 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4554) );
  MUX2_X1 U5121 ( .A(n4554), .B(n4553), .S(n4759), .Z(n4555) );
  OAI21_X1 U5122 ( .B1(n4557), .B2(n4556), .A(n4555), .ZN(U3493) );
  MUX2_X1 U5123 ( .A(DATAI_30_), .B(n4558), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U5124 ( .A(DATAI_26_), .B(n4559), .S(STATE_REG_SCAN_IN), .Z(U3326)
         );
  MUX2_X1 U5125 ( .A(DATAI_24_), .B(n4560), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U5126 ( .A(DATAI_22_), .B(n4561), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U5127 ( .A(DATAI_20_), .B(n4562), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5128 ( .A(DATAI_19_), .B(n4563), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U5129 ( .A(n4564), .B(DATAI_8_), .S(U3149), .Z(U3344) );
  MUX2_X1 U5130 ( .A(n4565), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5131 ( .A(DATAI_4_), .B(n4566), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5132 ( .A(n4567), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5133 ( .A(n4568), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  INV_X1 U5134 ( .A(DATAI_28_), .ZN(n4569) );
  AOI22_X1 U5135 ( .A1(STATE_REG_SCAN_IN), .A2(n4570), .B1(n4569), .B2(U3149), 
        .ZN(U3324) );
  NOR2_X1 U5136 ( .A1(STATE_REG_SCAN_IN), .A2(n4931), .ZN(n4672) );
  OAI22_X1 U5137 ( .A1(n4574), .A2(n4573), .B1(n4572), .B2(n4571), .ZN(n4575)
         );
  AOI211_X1 U5138 ( .C1(n4577), .C2(n4576), .A(n4672), .B(n4575), .ZN(n4584)
         );
  AOI21_X1 U5139 ( .B1(n4578), .B2(n3901), .A(n3900), .ZN(n4579) );
  XOR2_X1 U5140 ( .A(n4580), .B(n4579), .Z(n4582) );
  NAND2_X1 U5141 ( .A1(n4582), .A2(n4581), .ZN(n4583) );
  OAI211_X1 U5142 ( .C1(n4586), .C2(n4585), .A(n4584), .B(n4583), .ZN(U3223)
         );
  AOI22_X1 U5143 ( .A1(n4587), .A2(n4707), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4713), .ZN(n4588) );
  OAI21_X1 U5144 ( .B1(n4713), .B2(n4589), .A(n4588), .ZN(U3261) );
  INV_X1 U5145 ( .A(n4592), .ZN(n4590) );
  OAI211_X1 U5146 ( .C1(REG1_REG_0__SCAN_IN), .C2(n4591), .A(n4593), .B(n4590), 
        .ZN(n4596) );
  AOI22_X1 U5147 ( .A1(n4593), .A2(n4592), .B1(n4684), .B2(n2928), .ZN(n4595)
         );
  AOI22_X1 U5148 ( .A1(ADDR_REG_0__SCAN_IN), .A2(n4683), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n4594) );
  OAI221_X1 U5149 ( .B1(IR_REG_0__SCAN_IN), .B2(n4596), .C1(n2289), .C2(n4595), 
        .A(n4594), .ZN(U3240) );
  OAI211_X1 U5150 ( .C1(n4599), .C2(n4598), .A(n4684), .B(n4597), .ZN(n4604)
         );
  OAI211_X1 U5151 ( .C1(n4602), .C2(n4601), .A(n4640), .B(n4600), .ZN(n4603)
         );
  OAI211_X1 U5152 ( .C1(n4689), .C2(n4729), .A(n4604), .B(n4603), .ZN(n4605)
         );
  AOI211_X1 U5153 ( .C1(n4683), .C2(ADDR_REG_9__SCAN_IN), .A(n4606), .B(n4605), 
        .ZN(n4607) );
  INV_X1 U5154 ( .A(n4607), .ZN(U3249) );
  OAI211_X1 U5155 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4610), .A(n4640), .B(n4609), .ZN(n4612) );
  NAND2_X1 U5156 ( .A1(n4612), .A2(n4611), .ZN(n4613) );
  AOI21_X1 U5157 ( .B1(n4683), .B2(ADDR_REG_10__SCAN_IN), .A(n4613), .ZN(n4617) );
  OAI211_X1 U5158 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4615), .A(n4684), .B(n4614), .ZN(n4616) );
  OAI211_X1 U5159 ( .C1(n4689), .C2(n2847), .A(n4617), .B(n4616), .ZN(U3250)
         );
  OAI211_X1 U5160 ( .C1(n4620), .C2(n4619), .A(n4684), .B(n4618), .ZN(n4625)
         );
  OAI211_X1 U5161 ( .C1(n4623), .C2(n4622), .A(n4640), .B(n4621), .ZN(n4624)
         );
  OAI211_X1 U5162 ( .C1(n4689), .C2(n4727), .A(n4625), .B(n4624), .ZN(n4626)
         );
  AOI211_X1 U5163 ( .C1(n4683), .C2(ADDR_REG_11__SCAN_IN), .A(n4627), .B(n4626), .ZN(n4628) );
  INV_X1 U5164 ( .A(n4628), .ZN(U3251) );
  OAI211_X1 U5165 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4631), .A(n4684), .B(n4630), .ZN(n4635) );
  OAI211_X1 U5166 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4633), .A(n4640), .B(n4632), .ZN(n4634) );
  OAI211_X1 U5167 ( .C1(n4689), .C2(n2851), .A(n4635), .B(n4634), .ZN(n4636)
         );
  AOI211_X1 U5168 ( .C1(n4683), .C2(ADDR_REG_12__SCAN_IN), .A(n4637), .B(n4636), .ZN(n4638) );
  INV_X1 U5169 ( .A(n4638), .ZN(U3252) );
  AOI21_X1 U5170 ( .B1(n3683), .B2(n4651), .A(n4639), .ZN(n4643) );
  OAI21_X1 U5171 ( .B1(n4643), .B2(n4642), .A(n4640), .ZN(n4641) );
  AOI21_X1 U5172 ( .B1(n4643), .B2(n4642), .A(n4641), .ZN(n4644) );
  AOI211_X1 U5173 ( .C1(n4683), .C2(ADDR_REG_13__SCAN_IN), .A(n4645), .B(n4644), .ZN(n4650) );
  OAI211_X1 U5174 ( .C1(n4648), .C2(n4647), .A(n4684), .B(n4646), .ZN(n4649)
         );
  OAI211_X1 U5175 ( .C1(n4689), .C2(n4651), .A(n4650), .B(n4649), .ZN(U3253)
         );
  AOI211_X1 U5176 ( .C1(n3743), .C2(n4653), .A(n4652), .B(n4677), .ZN(n4654)
         );
  AOI211_X1 U5177 ( .C1(n4683), .C2(ADDR_REG_14__SCAN_IN), .A(n4655), .B(n4654), .ZN(n4659) );
  OAI211_X1 U5178 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4657), .A(n4684), .B(n4656), .ZN(n4658) );
  OAI211_X1 U5179 ( .C1(n4689), .C2(n4723), .A(n4659), .B(n4658), .ZN(U3254)
         );
  AOI211_X1 U5180 ( .C1(n2272), .C2(n4661), .A(n4660), .B(n4677), .ZN(n4662)
         );
  AOI211_X1 U5181 ( .C1(n4683), .C2(ADDR_REG_15__SCAN_IN), .A(n4663), .B(n4662), .ZN(n4668) );
  OAI211_X1 U5182 ( .C1(n4666), .C2(n4665), .A(n4684), .B(n4664), .ZN(n4667)
         );
  OAI211_X1 U5183 ( .C1(n4689), .C2(n4721), .A(n4668), .B(n4667), .ZN(U3255)
         );
  AOI221_X1 U5184 ( .B1(n4670), .B2(n4669), .C1(n4370), .C2(n4669), .A(n4677), 
        .ZN(n4671) );
  AOI211_X1 U5185 ( .C1(n4683), .C2(ADDR_REG_16__SCAN_IN), .A(n4672), .B(n4671), .ZN(n4676) );
  OAI221_X1 U5186 ( .B1(n4674), .B2(REG1_REG_16__SCAN_IN), .C1(n4674), .C2(
        n4673), .A(n4684), .ZN(n4675) );
  OAI211_X1 U5187 ( .C1(n4689), .C2(n4720), .A(n4676), .B(n4675), .ZN(U3256)
         );
  AOI221_X1 U5188 ( .B1(n4680), .B2(n4679), .C1(n4678), .C2(n4679), .A(n4677), 
        .ZN(n4681) );
  AOI211_X1 U5189 ( .C1(n4683), .C2(ADDR_REG_17__SCAN_IN), .A(n4682), .B(n4681), .ZN(n4688) );
  OAI221_X1 U5190 ( .B1(n4686), .B2(n2266), .C1(n4686), .C2(n4685), .A(n4684), 
        .ZN(n4687) );
  OAI211_X1 U5191 ( .C1(n4718), .C2(n4689), .A(n4688), .B(n4687), .ZN(U3257)
         );
  INV_X1 U5192 ( .A(n4690), .ZN(n4691) );
  AOI22_X1 U5193 ( .A1(n4691), .A2(n4705), .B1(REG2_REG_10__SCAN_IN), .B2(
        n4713), .ZN(n4696) );
  INV_X1 U5194 ( .A(n4692), .ZN(n4693) );
  AOI22_X1 U5195 ( .A1(n4694), .A2(n4708), .B1(n4707), .B2(n4693), .ZN(n4695)
         );
  OAI211_X1 U5196 ( .C1(n4713), .C2(n4697), .A(n4696), .B(n4695), .ZN(U3280)
         );
  AOI22_X1 U5197 ( .A1(n4698), .A2(n4705), .B1(REG2_REG_8__SCAN_IN), .B2(n4713), .ZN(n4703) );
  INV_X1 U5198 ( .A(n4699), .ZN(n4700) );
  AOI22_X1 U5199 ( .A1(n4701), .A2(n4708), .B1(n4707), .B2(n4700), .ZN(n4702)
         );
  OAI211_X1 U5200 ( .C1(n4713), .C2(n4704), .A(n4703), .B(n4702), .ZN(U3282)
         );
  AOI22_X1 U5201 ( .A1(REG2_REG_2__SCAN_IN), .A2(n4713), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4705), .ZN(n4711) );
  AOI22_X1 U5202 ( .A1(n4709), .A2(n4708), .B1(n4707), .B2(n4706), .ZN(n4710)
         );
  OAI211_X1 U5203 ( .C1(n4713), .C2(n4712), .A(n4711), .B(n4710), .ZN(U3288)
         );
  INV_X1 U5204 ( .A(D_REG_31__SCAN_IN), .ZN(n4914) );
  NOR2_X1 U5205 ( .A1(n4715), .A2(n4914), .ZN(U3291) );
  AND2_X1 U5206 ( .A1(n4714), .A2(D_REG_30__SCAN_IN), .ZN(U3292) );
  INV_X1 U5207 ( .A(D_REG_29__SCAN_IN), .ZN(n4920) );
  NOR2_X1 U5208 ( .A1(n4715), .A2(n4920), .ZN(U3293) );
  INV_X1 U5209 ( .A(D_REG_28__SCAN_IN), .ZN(n4910) );
  NOR2_X1 U5210 ( .A1(n4715), .A2(n4910), .ZN(U3294) );
  INV_X1 U5211 ( .A(D_REG_27__SCAN_IN), .ZN(n5087) );
  NOR2_X1 U5212 ( .A1(n4715), .A2(n5087), .ZN(U3295) );
  INV_X1 U5213 ( .A(D_REG_26__SCAN_IN), .ZN(n5055) );
  NOR2_X1 U5214 ( .A1(n4715), .A2(n5055), .ZN(U3296) );
  AND2_X1 U5215 ( .A1(n4714), .A2(D_REG_25__SCAN_IN), .ZN(U3297) );
  INV_X1 U5216 ( .A(D_REG_24__SCAN_IN), .ZN(n4799) );
  NOR2_X1 U5217 ( .A1(n4715), .A2(n4799), .ZN(U3298) );
  AND2_X1 U5218 ( .A1(n4714), .A2(D_REG_23__SCAN_IN), .ZN(U3299) );
  INV_X1 U5219 ( .A(D_REG_22__SCAN_IN), .ZN(n5056) );
  NOR2_X1 U5220 ( .A1(n4715), .A2(n5056), .ZN(U3300) );
  INV_X1 U5221 ( .A(D_REG_21__SCAN_IN), .ZN(n4877) );
  NOR2_X1 U5222 ( .A1(n4715), .A2(n4877), .ZN(U3301) );
  INV_X1 U5223 ( .A(D_REG_20__SCAN_IN), .ZN(n5071) );
  NOR2_X1 U5224 ( .A1(n4715), .A2(n5071), .ZN(U3302) );
  INV_X1 U5225 ( .A(D_REG_19__SCAN_IN), .ZN(n5077) );
  NOR2_X1 U5226 ( .A1(n4715), .A2(n5077), .ZN(U3303) );
  INV_X1 U5227 ( .A(D_REG_18__SCAN_IN), .ZN(n5078) );
  NOR2_X1 U5228 ( .A1(n4715), .A2(n5078), .ZN(U3304) );
  AND2_X1 U5229 ( .A1(n4714), .A2(D_REG_17__SCAN_IN), .ZN(U3305) );
  INV_X1 U5230 ( .A(D_REG_16__SCAN_IN), .ZN(n5074) );
  NOR2_X1 U5231 ( .A1(n4715), .A2(n5074), .ZN(U3306) );
  INV_X1 U5232 ( .A(D_REG_15__SCAN_IN), .ZN(n5081) );
  NOR2_X1 U5233 ( .A1(n4715), .A2(n5081), .ZN(U3307) );
  AND2_X1 U5234 ( .A1(n4714), .A2(D_REG_14__SCAN_IN), .ZN(U3308) );
  INV_X1 U5235 ( .A(D_REG_13__SCAN_IN), .ZN(n5075) );
  NOR2_X1 U5236 ( .A1(n4715), .A2(n5075), .ZN(U3309) );
  INV_X1 U5237 ( .A(D_REG_12__SCAN_IN), .ZN(n4846) );
  NOR2_X1 U5238 ( .A1(n4715), .A2(n4846), .ZN(U3310) );
  AND2_X1 U5239 ( .A1(n4714), .A2(D_REG_11__SCAN_IN), .ZN(U3311) );
  INV_X1 U5240 ( .A(D_REG_10__SCAN_IN), .ZN(n5072) );
  NOR2_X1 U5241 ( .A1(n4715), .A2(n5072), .ZN(U3312) );
  INV_X1 U5242 ( .A(D_REG_9__SCAN_IN), .ZN(n4933) );
  NOR2_X1 U5243 ( .A1(n4715), .A2(n4933), .ZN(U3313) );
  INV_X1 U5244 ( .A(D_REG_8__SCAN_IN), .ZN(n5052) );
  NOR2_X1 U5245 ( .A1(n4715), .A2(n5052), .ZN(U3314) );
  INV_X1 U5246 ( .A(D_REG_7__SCAN_IN), .ZN(n5088) );
  NOR2_X1 U5247 ( .A1(n4715), .A2(n5088), .ZN(U3315) );
  INV_X1 U5248 ( .A(D_REG_6__SCAN_IN), .ZN(n5061) );
  NOR2_X1 U5249 ( .A1(n4715), .A2(n5061), .ZN(U3316) );
  INV_X1 U5250 ( .A(D_REG_5__SCAN_IN), .ZN(n5080) );
  NOR2_X1 U5251 ( .A1(n4715), .A2(n5080), .ZN(U3317) );
  INV_X1 U5252 ( .A(D_REG_4__SCAN_IN), .ZN(n5053) );
  NOR2_X1 U5253 ( .A1(n4715), .A2(n5053), .ZN(U3318) );
  INV_X1 U5254 ( .A(D_REG_3__SCAN_IN), .ZN(n4884) );
  NOR2_X1 U5255 ( .A1(n4715), .A2(n4884), .ZN(U3319) );
  INV_X1 U5256 ( .A(D_REG_2__SCAN_IN), .ZN(n4922) );
  NOR2_X1 U5257 ( .A1(n4715), .A2(n4922), .ZN(U3320) );
  INV_X1 U5258 ( .A(DATAI_23_), .ZN(n5117) );
  AOI21_X1 U5259 ( .B1(U3149), .B2(n5117), .A(n4716), .ZN(U3329) );
  AOI22_X1 U5260 ( .A1(STATE_REG_SCAN_IN), .A2(n4717), .B1(n4796), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5261 ( .A1(STATE_REG_SCAN_IN), .A2(n4718), .B1(n2659), .B2(U3149), 
        .ZN(U3335) );
  AOI22_X1 U5262 ( .A1(STATE_REG_SCAN_IN), .A2(n4720), .B1(n4719), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5263 ( .A(DATAI_15_), .ZN(n4999) );
  AOI22_X1 U5264 ( .A1(STATE_REG_SCAN_IN), .A2(n4721), .B1(n4999), .B2(U3149), 
        .ZN(U3337) );
  AOI22_X1 U5265 ( .A1(STATE_REG_SCAN_IN), .A2(n4723), .B1(n4722), .B2(U3149), 
        .ZN(U3338) );
  OAI22_X1 U5266 ( .A1(U3149), .A2(n4724), .B1(DATAI_13_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4725) );
  INV_X1 U5267 ( .A(n4725), .ZN(U3339) );
  INV_X1 U5268 ( .A(DATAI_12_), .ZN(n4726) );
  AOI22_X1 U5269 ( .A1(STATE_REG_SCAN_IN), .A2(n2851), .B1(n4726), .B2(U3149), 
        .ZN(U3340) );
  AOI22_X1 U5270 ( .A1(STATE_REG_SCAN_IN), .A2(n4727), .B1(n2591), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5271 ( .A(DATAI_10_), .ZN(n5102) );
  AOI22_X1 U5272 ( .A1(STATE_REG_SCAN_IN), .A2(n2847), .B1(n5102), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5273 ( .A(DATAI_9_), .ZN(n4728) );
  AOI22_X1 U5274 ( .A1(STATE_REG_SCAN_IN), .A2(n4729), .B1(n4728), .B2(U3149), 
        .ZN(U3343) );
  AOI211_X1 U5275 ( .C1(n4756), .C2(n4732), .A(n4731), .B(n4730), .ZN(n4760)
         );
  INV_X1 U5276 ( .A(REG0_REG_0__SCAN_IN), .ZN(n4870) );
  AOI22_X1 U5277 ( .A1(n4759), .A2(n4760), .B1(n4870), .B2(n4757), .ZN(U3467)
         );
  NOR2_X1 U5278 ( .A1(n4734), .A2(n4733), .ZN(n4736) );
  AOI211_X1 U5279 ( .C1(n4738), .C2(n4737), .A(n4736), .B(n4735), .ZN(n4762)
         );
  INV_X1 U5280 ( .A(REG0_REG_1__SCAN_IN), .ZN(n5043) );
  AOI22_X1 U5281 ( .A1(n4759), .A2(n4762), .B1(n5043), .B2(n4757), .ZN(U3469)
         );
  INV_X1 U5282 ( .A(n4739), .ZN(n4743) );
  INV_X1 U5283 ( .A(n4740), .ZN(n4742) );
  AOI211_X1 U5284 ( .C1(n4743), .C2(n4756), .A(n4742), .B(n4741), .ZN(n4764)
         );
  INV_X1 U5285 ( .A(REG0_REG_4__SCAN_IN), .ZN(n4744) );
  AOI22_X1 U5286 ( .A1(n4759), .A2(n4764), .B1(n4744), .B2(n4757), .ZN(U3475)
         );
  AND3_X1 U5287 ( .A1(n3492), .A2(n4746), .A3(n4745), .ZN(n4748) );
  NOR3_X1 U5288 ( .A1(n4749), .A2(n4748), .A3(n4747), .ZN(n4766) );
  INV_X1 U5289 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4750) );
  AOI22_X1 U5290 ( .A1(n4759), .A2(n4766), .B1(n4750), .B2(n4757), .ZN(U3481)
         );
  NOR2_X1 U5291 ( .A1(n4752), .A2(n4751), .ZN(n4754) );
  AOI211_X1 U5292 ( .C1(n4756), .C2(n4755), .A(n4754), .B(n4753), .ZN(n4769)
         );
  INV_X1 U5293 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4758) );
  AOI22_X1 U5294 ( .A1(n4759), .A2(n4769), .B1(n4758), .B2(n4757), .ZN(U3489)
         );
  AOI22_X1 U5295 ( .A1(n4770), .A2(n4760), .B1(n2928), .B2(n4767), .ZN(U3518)
         );
  INV_X1 U5296 ( .A(REG1_REG_1__SCAN_IN), .ZN(n4761) );
  AOI22_X1 U5297 ( .A1(n4770), .A2(n4762), .B1(n4761), .B2(n4767), .ZN(U3519)
         );
  INV_X1 U5298 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4763) );
  AOI22_X1 U5299 ( .A1(n4770), .A2(n4764), .B1(n4763), .B2(n4767), .ZN(U3522)
         );
  INV_X1 U5300 ( .A(REG1_REG_7__SCAN_IN), .ZN(n4765) );
  AOI22_X1 U5301 ( .A1(n4770), .A2(n4766), .B1(n4765), .B2(n4767), .ZN(U3525)
         );
  AOI22_X1 U5302 ( .A1(n4770), .A2(n4769), .B1(n4768), .B2(n4767), .ZN(U3529)
         );
  OAI22_X1 U5303 ( .A1(DATAI_28_), .A2(keyinput_g3), .B1(keyinput_g0), .B2(
        DATAI_31_), .ZN(n4771) );
  AOI221_X1 U5304 ( .B1(DATAI_28_), .B2(keyinput_g3), .C1(DATAI_31_), .C2(
        keyinput_g0), .A(n4771), .ZN(n4778) );
  OAI22_X1 U5305 ( .A1(IR_REG_23__SCAN_IN), .A2(keyinput_g78), .B1(
        keyinput_g14), .B2(DATAI_17_), .ZN(n4772) );
  AOI221_X1 U5306 ( .B1(IR_REG_23__SCAN_IN), .B2(keyinput_g78), .C1(DATAI_17_), 
        .C2(keyinput_g14), .A(n4772), .ZN(n4777) );
  OAI22_X1 U5307 ( .A1(D_REG_6__SCAN_IN), .A2(keyinput_g93), .B1(DATAI_27_), 
        .B2(keyinput_g4), .ZN(n4773) );
  AOI221_X1 U5308 ( .B1(D_REG_6__SCAN_IN), .B2(keyinput_g93), .C1(keyinput_g4), 
        .C2(DATAI_27_), .A(n4773), .ZN(n4776) );
  OAI22_X1 U5309 ( .A1(IR_REG_22__SCAN_IN), .A2(keyinput_g77), .B1(
        keyinput_g23), .B2(DATAI_8_), .ZN(n4774) );
  AOI221_X1 U5310 ( .B1(IR_REG_22__SCAN_IN), .B2(keyinput_g77), .C1(DATAI_8_), 
        .C2(keyinput_g23), .A(n4774), .ZN(n4775) );
  NAND4_X1 U5311 ( .A1(n4778), .A2(n4777), .A3(n4776), .A4(n4775), .ZN(n4809)
         );
  OAI22_X1 U5312 ( .A1(REG3_REG_12__SCAN_IN), .A2(keyinput_g44), .B1(
        keyinput_g123), .B2(REG0_REG_4__SCAN_IN), .ZN(n4779) );
  AOI221_X1 U5313 ( .B1(REG3_REG_12__SCAN_IN), .B2(keyinput_g44), .C1(
        REG0_REG_4__SCAN_IN), .C2(keyinput_g123), .A(n4779), .ZN(n4786) );
  OAI22_X1 U5314 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput_g52), .B1(DATAI_26_), 
        .B2(keyinput_g5), .ZN(n4780) );
  AOI221_X1 U5315 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput_g52), .C1(
        keyinput_g5), .C2(DATAI_26_), .A(n4780), .ZN(n4785) );
  OAI22_X1 U5316 ( .A1(IR_REG_6__SCAN_IN), .A2(keyinput_g61), .B1(keyinput_g43), .B2(REG3_REG_21__SCAN_IN), .ZN(n4781) );
  AOI221_X1 U5317 ( .B1(IR_REG_6__SCAN_IN), .B2(keyinput_g61), .C1(
        REG3_REG_21__SCAN_IN), .C2(keyinput_g43), .A(n4781), .ZN(n4784) );
  OAI22_X1 U5318 ( .A1(IR_REG_27__SCAN_IN), .A2(keyinput_g82), .B1(DATAI_9_), 
        .B2(keyinput_g22), .ZN(n4782) );
  AOI221_X1 U5319 ( .B1(IR_REG_27__SCAN_IN), .B2(keyinput_g82), .C1(
        keyinput_g22), .C2(DATAI_9_), .A(n4782), .ZN(n4783) );
  NAND4_X1 U5320 ( .A1(n4786), .A2(n4785), .A3(n4784), .A4(n4783), .ZN(n4808)
         );
  OAI22_X1 U5321 ( .A1(IR_REG_26__SCAN_IN), .A2(keyinput_g81), .B1(
        IR_REG_21__SCAN_IN), .B2(keyinput_g76), .ZN(n4787) );
  AOI221_X1 U5322 ( .B1(IR_REG_26__SCAN_IN), .B2(keyinput_g81), .C1(
        keyinput_g76), .C2(IR_REG_21__SCAN_IN), .A(n4787), .ZN(n4794) );
  OAI22_X1 U5323 ( .A1(IR_REG_13__SCAN_IN), .A2(keyinput_g68), .B1(
        keyinput_g15), .B2(DATAI_16_), .ZN(n4788) );
  AOI221_X1 U5324 ( .B1(IR_REG_13__SCAN_IN), .B2(keyinput_g68), .C1(DATAI_16_), 
        .C2(keyinput_g15), .A(n4788), .ZN(n4793) );
  OAI22_X1 U5325 ( .A1(D_REG_26__SCAN_IN), .A2(keyinput_g113), .B1(
        keyinput_g31), .B2(DATAI_0_), .ZN(n4789) );
  AOI221_X1 U5326 ( .B1(D_REG_26__SCAN_IN), .B2(keyinput_g113), .C1(DATAI_0_), 
        .C2(keyinput_g31), .A(n4789), .ZN(n4792) );
  OAI22_X1 U5327 ( .A1(IR_REG_17__SCAN_IN), .A2(keyinput_g72), .B1(
        keyinput_g98), .B2(D_REG_11__SCAN_IN), .ZN(n4790) );
  AOI221_X1 U5328 ( .B1(IR_REG_17__SCAN_IN), .B2(keyinput_g72), .C1(
        D_REG_11__SCAN_IN), .C2(keyinput_g98), .A(n4790), .ZN(n4791) );
  NAND4_X1 U5329 ( .A1(n4794), .A2(n4793), .A3(n4792), .A4(n4791), .ZN(n4807)
         );
  AOI22_X1 U5330 ( .A1(n4796), .A2(keyinput_g13), .B1(n5032), .B2(keyinput_g10), .ZN(n4795) );
  OAI221_X1 U5331 ( .B1(n4796), .B2(keyinput_g13), .C1(n5032), .C2(
        keyinput_g10), .A(n4795), .ZN(n4805) );
  AOI22_X1 U5332 ( .A1(n2289), .A2(keyinput_g55), .B1(keyinput_g114), .B2(
        n5087), .ZN(n4797) );
  OAI221_X1 U5333 ( .B1(n2289), .B2(keyinput_g55), .C1(n5087), .C2(
        keyinput_g114), .A(n4797), .ZN(n4804) );
  AOI22_X1 U5334 ( .A1(IR_REG_16__SCAN_IN), .A2(keyinput_g71), .B1(n4799), 
        .B2(keyinput_g111), .ZN(n4798) );
  OAI221_X1 U5335 ( .B1(IR_REG_16__SCAN_IN), .B2(keyinput_g71), .C1(n4799), 
        .C2(keyinput_g111), .A(n4798), .ZN(n4803) );
  XNOR2_X1 U5336 ( .A(IR_REG_28__SCAN_IN), .B(keyinput_g83), .ZN(n4801) );
  XNOR2_X1 U5337 ( .A(REG3_REG_24__SCAN_IN), .B(keyinput_g49), .ZN(n4800) );
  NAND2_X1 U5338 ( .A1(n4801), .A2(n4800), .ZN(n4802) );
  OR4_X1 U5339 ( .A1(n4805), .A2(n4804), .A3(n4803), .A4(n4802), .ZN(n4806) );
  NOR4_X1 U5340 ( .A1(n4809), .A2(n4808), .A3(n4807), .A4(n4806), .ZN(n5138)
         );
  OAI22_X1 U5341 ( .A1(D_REG_17__SCAN_IN), .A2(keyinput_g104), .B1(
        D_REG_14__SCAN_IN), .B2(keyinput_g101), .ZN(n4810) );
  AOI221_X1 U5342 ( .B1(D_REG_17__SCAN_IN), .B2(keyinput_g104), .C1(
        keyinput_g101), .C2(D_REG_14__SCAN_IN), .A(n4810), .ZN(n4817) );
  OAI22_X1 U5343 ( .A1(DATAI_14_), .A2(keyinput_g17), .B1(DATAI_13_), .B2(
        keyinput_g18), .ZN(n4811) );
  AOI221_X1 U5344 ( .B1(DATAI_14_), .B2(keyinput_g17), .C1(keyinput_g18), .C2(
        DATAI_13_), .A(n4811), .ZN(n4816) );
  OAI22_X1 U5345 ( .A1(DATAI_12_), .A2(keyinput_g19), .B1(DATAI_11_), .B2(
        keyinput_g20), .ZN(n4812) );
  AOI221_X1 U5346 ( .B1(DATAI_12_), .B2(keyinput_g19), .C1(keyinput_g20), .C2(
        DATAI_11_), .A(n4812), .ZN(n4815) );
  OAI22_X1 U5347 ( .A1(DATAI_7_), .A2(keyinput_g24), .B1(DATAI_5_), .B2(
        keyinput_g26), .ZN(n4813) );
  AOI221_X1 U5348 ( .B1(DATAI_7_), .B2(keyinput_g24), .C1(keyinput_g26), .C2(
        DATAI_5_), .A(n4813), .ZN(n4814) );
  NAND4_X1 U5349 ( .A1(n4817), .A2(n4816), .A3(n4815), .A4(n4814), .ZN(n4948)
         );
  OAI22_X1 U5350 ( .A1(DATAI_3_), .A2(keyinput_g28), .B1(keyinput_g29), .B2(
        DATAI_2_), .ZN(n4818) );
  AOI221_X1 U5351 ( .B1(DATAI_3_), .B2(keyinput_g28), .C1(DATAI_2_), .C2(
        keyinput_g29), .A(n4818), .ZN(n4843) );
  OAI22_X1 U5352 ( .A1(D_REG_25__SCAN_IN), .A2(keyinput_g112), .B1(
        D_REG_23__SCAN_IN), .B2(keyinput_g110), .ZN(n4819) );
  AOI221_X1 U5353 ( .B1(D_REG_25__SCAN_IN), .B2(keyinput_g112), .C1(
        keyinput_g110), .C2(D_REG_23__SCAN_IN), .A(n4819), .ZN(n4822) );
  OAI22_X1 U5354 ( .A1(D_REG_30__SCAN_IN), .A2(keyinput_g117), .B1(
        keyinput_g42), .B2(REG3_REG_1__SCAN_IN), .ZN(n4820) );
  AOI221_X1 U5355 ( .B1(D_REG_30__SCAN_IN), .B2(keyinput_g117), .C1(
        REG3_REG_1__SCAN_IN), .C2(keyinput_g42), .A(n4820), .ZN(n4821) );
  OAI211_X1 U5356 ( .C1(n5078), .C2(keyinput_g105), .A(n4822), .B(n4821), .ZN(
        n4823) );
  AOI21_X1 U5357 ( .B1(n5078), .B2(keyinput_g105), .A(n4823), .ZN(n4842) );
  AOI22_X1 U5358 ( .A1(REG0_REG_3__SCAN_IN), .A2(keyinput_g122), .B1(
        REG0_REG_5__SCAN_IN), .B2(keyinput_g124), .ZN(n4824) );
  OAI221_X1 U5359 ( .B1(REG0_REG_3__SCAN_IN), .B2(keyinput_g122), .C1(
        REG0_REG_5__SCAN_IN), .C2(keyinput_g124), .A(n4824), .ZN(n4831) );
  AOI22_X1 U5360 ( .A1(REG0_REG_6__SCAN_IN), .A2(keyinput_g125), .B1(
        REG0_REG_7__SCAN_IN), .B2(keyinput_g126), .ZN(n4825) );
  OAI221_X1 U5361 ( .B1(REG0_REG_6__SCAN_IN), .B2(keyinput_g125), .C1(
        REG0_REG_7__SCAN_IN), .C2(keyinput_g126), .A(n4825), .ZN(n4830) );
  AOI22_X1 U5362 ( .A1(REG3_REG_4__SCAN_IN), .A2(keyinput_g50), .B1(
        IR_REG_4__SCAN_IN), .B2(keyinput_g59), .ZN(n4826) );
  OAI221_X1 U5363 ( .B1(REG3_REG_4__SCAN_IN), .B2(keyinput_g50), .C1(
        IR_REG_4__SCAN_IN), .C2(keyinput_g59), .A(n4826), .ZN(n4829) );
  AOI22_X1 U5364 ( .A1(D_REG_10__SCAN_IN), .A2(keyinput_g97), .B1(
        IR_REG_2__SCAN_IN), .B2(keyinput_g57), .ZN(n4827) );
  OAI221_X1 U5365 ( .B1(D_REG_10__SCAN_IN), .B2(keyinput_g97), .C1(
        IR_REG_2__SCAN_IN), .C2(keyinput_g57), .A(n4827), .ZN(n4828) );
  NOR4_X1 U5366 ( .A1(n4831), .A2(n4830), .A3(n4829), .A4(n4828), .ZN(n4841)
         );
  AOI22_X1 U5367 ( .A1(REG3_REG_19__SCAN_IN), .A2(keyinput_g39), .B1(
        D_REG_0__SCAN_IN), .B2(keyinput_g87), .ZN(n4832) );
  OAI221_X1 U5368 ( .B1(REG3_REG_19__SCAN_IN), .B2(keyinput_g39), .C1(
        D_REG_0__SCAN_IN), .C2(keyinput_g87), .A(n4832), .ZN(n4839) );
  AOI22_X1 U5369 ( .A1(REG3_REG_23__SCAN_IN), .A2(keyinput_g36), .B1(
        IR_REG_29__SCAN_IN), .B2(keyinput_g84), .ZN(n4833) );
  OAI221_X1 U5370 ( .B1(REG3_REG_23__SCAN_IN), .B2(keyinput_g36), .C1(
        IR_REG_29__SCAN_IN), .C2(keyinput_g84), .A(n4833), .ZN(n4838) );
  AOI22_X1 U5371 ( .A1(DATAI_15_), .A2(keyinput_g16), .B1(IR_REG_9__SCAN_IN), 
        .B2(keyinput_g64), .ZN(n4834) );
  OAI221_X1 U5372 ( .B1(DATAI_15_), .B2(keyinput_g16), .C1(IR_REG_9__SCAN_IN), 
        .C2(keyinput_g64), .A(n4834), .ZN(n4837) );
  AOI22_X1 U5373 ( .A1(IR_REG_8__SCAN_IN), .A2(keyinput_g63), .B1(
        IR_REG_24__SCAN_IN), .B2(keyinput_g79), .ZN(n4835) );
  OAI221_X1 U5374 ( .B1(IR_REG_8__SCAN_IN), .B2(keyinput_g63), .C1(
        IR_REG_24__SCAN_IN), .C2(keyinput_g79), .A(n4835), .ZN(n4836) );
  NOR4_X1 U5375 ( .A1(n4839), .A2(n4838), .A3(n4837), .A4(n4836), .ZN(n4840)
         );
  NAND4_X1 U5376 ( .A1(n4843), .A2(n4842), .A3(n4841), .A4(n4840), .ZN(n4947)
         );
  INV_X1 U5377 ( .A(DATAI_6_), .ZN(n4845) );
  AOI22_X1 U5378 ( .A1(n5117), .A2(keyinput_g8), .B1(keyinput_g25), .B2(n4845), 
        .ZN(n4844) );
  OAI221_X1 U5379 ( .B1(n5117), .B2(keyinput_g8), .C1(n4845), .C2(keyinput_g25), .A(n4844), .ZN(n4850) );
  XNOR2_X1 U5380 ( .A(n4846), .B(keyinput_g99), .ZN(n4849) );
  XNOR2_X1 U5381 ( .A(n4847), .B(keyinput_g66), .ZN(n4848) );
  OR3_X1 U5382 ( .A1(n4850), .A2(n4849), .A3(n4848), .ZN(n4855) );
  AOI22_X1 U5383 ( .A1(n2741), .A2(keyinput_g74), .B1(keyinput_g94), .B2(n5088), .ZN(n4851) );
  OAI221_X1 U5384 ( .B1(n2741), .B2(keyinput_g74), .C1(n5088), .C2(
        keyinput_g94), .A(n4851), .ZN(n4854) );
  AOI22_X1 U5385 ( .A1(n2645), .A2(keyinput_g48), .B1(n5080), .B2(keyinput_g92), .ZN(n4852) );
  OAI221_X1 U5386 ( .B1(n2645), .B2(keyinput_g48), .C1(n5080), .C2(
        keyinput_g92), .A(n4852), .ZN(n4853) );
  NOR3_X1 U5387 ( .A1(n4855), .A2(n4854), .A3(n4853), .ZN(n4897) );
  INV_X1 U5388 ( .A(DATAI_22_), .ZN(n4857) );
  AOI22_X1 U5389 ( .A1(n4857), .A2(keyinput_g9), .B1(n2512), .B2(keyinput_g58), 
        .ZN(n4856) );
  OAI221_X1 U5390 ( .B1(n4857), .B2(keyinput_g9), .C1(n2512), .C2(keyinput_g58), .A(n4856), .ZN(n4868) );
  AOI22_X1 U5391 ( .A1(n4859), .A2(keyinput_g41), .B1(n5081), .B2(
        keyinput_g102), .ZN(n4858) );
  OAI221_X1 U5392 ( .B1(n4859), .B2(keyinput_g41), .C1(n5081), .C2(
        keyinput_g102), .A(n4858), .ZN(n4867) );
  INV_X1 U5393 ( .A(DATAI_19_), .ZN(n4862) );
  AOI22_X1 U5394 ( .A1(n4862), .A2(keyinput_g12), .B1(n4861), .B2(keyinput_g35), .ZN(n4860) );
  OAI221_X1 U5395 ( .B1(n4862), .B2(keyinput_g12), .C1(n4861), .C2(
        keyinput_g35), .A(n4860), .ZN(n4866) );
  AOI22_X1 U5396 ( .A1(n3792), .A2(keyinput_g85), .B1(keyinput_g6), .B2(n4864), 
        .ZN(n4863) );
  OAI221_X1 U5397 ( .B1(n3792), .B2(keyinput_g85), .C1(n4864), .C2(keyinput_g6), .A(n4863), .ZN(n4865) );
  NOR4_X1 U5398 ( .A1(n4868), .A2(n4867), .A3(n4866), .A4(n4865), .ZN(n4896)
         );
  INV_X1 U5399 ( .A(DATAI_24_), .ZN(n4871) );
  AOI22_X1 U5400 ( .A1(n4871), .A2(keyinput_g7), .B1(n4870), .B2(keyinput_g119), .ZN(n4869) );
  OAI221_X1 U5401 ( .B1(n4871), .B2(keyinput_g7), .C1(n4870), .C2(
        keyinput_g119), .A(n4869), .ZN(n4881) );
  AOI22_X1 U5402 ( .A1(n2296), .A2(keyinput_g65), .B1(keyinput_g53), .B2(n4873), .ZN(n4872) );
  OAI221_X1 U5403 ( .B1(n2296), .B2(keyinput_g65), .C1(n4873), .C2(
        keyinput_g53), .A(n4872), .ZN(n4880) );
  INV_X1 U5404 ( .A(REG0_REG_2__SCAN_IN), .ZN(n4875) );
  AOI22_X1 U5405 ( .A1(n5071), .A2(keyinput_g107), .B1(keyinput_g121), .B2(
        n4875), .ZN(n4874) );
  OAI221_X1 U5406 ( .B1(n5071), .B2(keyinput_g107), .C1(n4875), .C2(
        keyinput_g121), .A(n4874), .ZN(n4879) );
  AOI22_X1 U5407 ( .A1(n5118), .A2(keyinput_g88), .B1(keyinput_g108), .B2(
        n4877), .ZN(n4876) );
  OAI221_X1 U5408 ( .B1(n5118), .B2(keyinput_g88), .C1(n4877), .C2(
        keyinput_g108), .A(n4876), .ZN(n4878) );
  NOR4_X1 U5409 ( .A1(n4881), .A2(n4880), .A3(n4879), .A4(n4878), .ZN(n4895)
         );
  INV_X1 U5410 ( .A(DATAI_30_), .ZN(n4883) );
  AOI22_X1 U5411 ( .A1(n4884), .A2(keyinput_g90), .B1(keyinput_g1), .B2(n4883), 
        .ZN(n4882) );
  OAI221_X1 U5412 ( .B1(n4884), .B2(keyinput_g90), .C1(n4883), .C2(keyinput_g1), .A(n4882), .ZN(n4893) );
  AOI22_X1 U5413 ( .A1(n5040), .A2(keyinput_g70), .B1(keyinput_g47), .B2(n4886), .ZN(n4885) );
  OAI221_X1 U5414 ( .B1(n5040), .B2(keyinput_g70), .C1(n4886), .C2(
        keyinput_g47), .A(n4885), .ZN(n4892) );
  XNOR2_X1 U5415 ( .A(IR_REG_18__SCAN_IN), .B(keyinput_g73), .ZN(n4889) );
  XNOR2_X1 U5416 ( .A(REG3_REG_27__SCAN_IN), .B(keyinput_g34), .ZN(n4888) );
  XNOR2_X1 U5417 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_g60), .ZN(n4887) );
  NAND3_X1 U5418 ( .A1(n4889), .A2(n4888), .A3(n4887), .ZN(n4891) );
  XNOR2_X1 U5419 ( .A(n5052), .B(keyinput_g95), .ZN(n4890) );
  NOR4_X1 U5420 ( .A1(n4893), .A2(n4892), .A3(n4891), .A4(n4890), .ZN(n4894)
         );
  NAND4_X1 U5421 ( .A1(n4897), .A2(n4896), .A3(n4895), .A4(n4894), .ZN(n4946)
         );
  AOI22_X1 U5422 ( .A1(n5053), .A2(keyinput_g91), .B1(keyinput_g54), .B2(n2602), .ZN(n4898) );
  OAI221_X1 U5423 ( .B1(n5053), .B2(keyinput_g91), .C1(n2602), .C2(
        keyinput_g54), .A(n4898), .ZN(n4907) );
  AOI22_X1 U5424 ( .A1(n2743), .A2(keyinput_g75), .B1(keyinput_g127), .B2(
        n4900), .ZN(n4899) );
  OAI221_X1 U5425 ( .B1(n2743), .B2(keyinput_g75), .C1(n4900), .C2(
        keyinput_g127), .A(n4899), .ZN(n4906) );
  AOI22_X1 U5426 ( .A1(n2475), .A2(keyinput_g30), .B1(n5039), .B2(keyinput_g33), .ZN(n4901) );
  OAI221_X1 U5427 ( .B1(n2475), .B2(keyinput_g30), .C1(n5039), .C2(
        keyinput_g33), .A(n4901), .ZN(n4905) );
  AOI22_X1 U5428 ( .A1(n5056), .A2(keyinput_g109), .B1(keyinput_g2), .B2(n4903), .ZN(n4902) );
  OAI221_X1 U5429 ( .B1(n5056), .B2(keyinput_g109), .C1(n4903), .C2(
        keyinput_g2), .A(n4902), .ZN(n4904) );
  NOR4_X1 U5430 ( .A1(n4907), .A2(n4906), .A3(n4905), .A4(n4904), .ZN(n4944)
         );
  AOI22_X1 U5431 ( .A1(n5043), .A2(keyinput_g120), .B1(n2559), .B2(
        keyinput_g51), .ZN(n4908) );
  OAI221_X1 U5432 ( .B1(n5043), .B2(keyinput_g120), .C1(n2559), .C2(
        keyinput_g51), .A(n4908), .ZN(n4918) );
  INV_X1 U5433 ( .A(DATAI_20_), .ZN(n5101) );
  AOI22_X1 U5434 ( .A1(n5101), .A2(keyinput_g11), .B1(n4910), .B2(
        keyinput_g115), .ZN(n4909) );
  OAI221_X1 U5435 ( .B1(n5101), .B2(keyinput_g11), .C1(n4910), .C2(
        keyinput_g115), .A(n4909), .ZN(n4917) );
  XNOR2_X1 U5436 ( .A(IR_REG_14__SCAN_IN), .B(keyinput_g69), .ZN(n4913) );
  XNOR2_X1 U5437 ( .A(DATAI_4_), .B(keyinput_g27), .ZN(n4912) );
  XNOR2_X1 U5438 ( .A(DATAI_10_), .B(keyinput_g21), .ZN(n4911) );
  NAND3_X1 U5439 ( .A1(n4913), .A2(n4912), .A3(n4911), .ZN(n4916) );
  XNOR2_X1 U5440 ( .A(n4914), .B(keyinput_g118), .ZN(n4915) );
  NOR4_X1 U5441 ( .A1(n4918), .A2(n4917), .A3(n4916), .A4(n4915), .ZN(n4943)
         );
  AOI22_X1 U5442 ( .A1(n4920), .A2(keyinput_g116), .B1(keyinput_g103), .B2(
        n5074), .ZN(n4919) );
  OAI221_X1 U5443 ( .B1(n4920), .B2(keyinput_g116), .C1(n5074), .C2(
        keyinput_g103), .A(n4919), .ZN(n4929) );
  AOI22_X1 U5444 ( .A1(n5057), .A2(keyinput_g56), .B1(keyinput_g89), .B2(n4922), .ZN(n4921) );
  OAI221_X1 U5445 ( .B1(n5057), .B2(keyinput_g56), .C1(n4922), .C2(
        keyinput_g89), .A(n4921), .ZN(n4928) );
  XNOR2_X1 U5446 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput_g37), .ZN(n4926) );
  XNOR2_X1 U5447 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_g86), .ZN(n4925) );
  XNOR2_X1 U5448 ( .A(IR_REG_25__SCAN_IN), .B(keyinput_g80), .ZN(n4924) );
  XNOR2_X1 U5449 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_g38), .ZN(n4923) );
  NAND4_X1 U5450 ( .A1(n4926), .A2(n4925), .A3(n4924), .A4(n4923), .ZN(n4927)
         );
  NOR3_X1 U5451 ( .A1(n4929), .A2(n4928), .A3(n4927), .ZN(n4942) );
  AOI22_X1 U5452 ( .A1(n4931), .A2(keyinput_g46), .B1(n5077), .B2(
        keyinput_g106), .ZN(n4930) );
  OAI221_X1 U5453 ( .B1(n4931), .B2(keyinput_g46), .C1(n5077), .C2(
        keyinput_g106), .A(n4930), .ZN(n4940) );
  AOI22_X1 U5454 ( .A1(n5075), .A2(keyinput_g100), .B1(n4933), .B2(
        keyinput_g96), .ZN(n4932) );
  OAI221_X1 U5455 ( .B1(n5075), .B2(keyinput_g100), .C1(n4933), .C2(
        keyinput_g96), .A(n4932), .ZN(n4939) );
  XOR2_X1 U5456 ( .A(n3772), .B(keyinput_g40), .Z(n4937) );
  XNOR2_X1 U5457 ( .A(IR_REG_7__SCAN_IN), .B(keyinput_g62), .ZN(n4936) );
  XNOR2_X1 U5458 ( .A(REG3_REG_25__SCAN_IN), .B(keyinput_g45), .ZN(n4935) );
  XNOR2_X1 U5459 ( .A(IR_REG_12__SCAN_IN), .B(keyinput_g67), .ZN(n4934) );
  NAND4_X1 U5460 ( .A1(n4937), .A2(n4936), .A3(n4935), .A4(n4934), .ZN(n4938)
         );
  NOR3_X1 U5461 ( .A1(n4940), .A2(n4939), .A3(n4938), .ZN(n4941) );
  NAND4_X1 U5462 ( .A1(n4944), .A2(n4943), .A3(n4942), .A4(n4941), .ZN(n4945)
         );
  NOR4_X1 U5463 ( .A1(n4948), .A2(n4947), .A3(n4946), .A4(n4945), .ZN(n5137)
         );
  OAI22_X1 U5464 ( .A1(DATAI_12_), .A2(keyinput_f19), .B1(DATAI_11_), .B2(
        keyinput_f20), .ZN(n4949) );
  AOI221_X1 U5465 ( .B1(DATAI_12_), .B2(keyinput_f19), .C1(keyinput_f20), .C2(
        DATAI_11_), .A(n4949), .ZN(n4956) );
  OAI22_X1 U5466 ( .A1(DATAI_9_), .A2(keyinput_f22), .B1(DATAI_8_), .B2(
        keyinput_f23), .ZN(n4950) );
  AOI221_X1 U5467 ( .B1(DATAI_9_), .B2(keyinput_f22), .C1(keyinput_f23), .C2(
        DATAI_8_), .A(n4950), .ZN(n4955) );
  OAI22_X1 U5468 ( .A1(DATAI_7_), .A2(keyinput_f24), .B1(DATAI_5_), .B2(
        keyinput_f26), .ZN(n4951) );
  AOI221_X1 U5469 ( .B1(DATAI_7_), .B2(keyinput_f24), .C1(keyinput_f26), .C2(
        DATAI_5_), .A(n4951), .ZN(n4954) );
  OAI22_X1 U5470 ( .A1(REG0_REG_3__SCAN_IN), .A2(keyinput_f122), .B1(
        REG0_REG_4__SCAN_IN), .B2(keyinput_f123), .ZN(n4952) );
  AOI221_X1 U5471 ( .B1(REG0_REG_3__SCAN_IN), .B2(keyinput_f122), .C1(
        keyinput_f123), .C2(REG0_REG_4__SCAN_IN), .A(n4952), .ZN(n4953) );
  NAND4_X1 U5472 ( .A1(n4956), .A2(n4955), .A3(n4954), .A4(n4953), .ZN(n4984)
         );
  OAI22_X1 U5473 ( .A1(REG0_REG_6__SCAN_IN), .A2(keyinput_f125), .B1(
        keyinput_f124), .B2(REG0_REG_5__SCAN_IN), .ZN(n4957) );
  AOI221_X1 U5474 ( .B1(REG0_REG_6__SCAN_IN), .B2(keyinput_f125), .C1(
        REG0_REG_5__SCAN_IN), .C2(keyinput_f124), .A(n4957), .ZN(n4964) );
  OAI22_X1 U5475 ( .A1(IR_REG_11__SCAN_IN), .A2(keyinput_f66), .B1(
        keyinput_f126), .B2(REG0_REG_7__SCAN_IN), .ZN(n4958) );
  AOI221_X1 U5476 ( .B1(IR_REG_11__SCAN_IN), .B2(keyinput_f66), .C1(
        REG0_REG_7__SCAN_IN), .C2(keyinput_f126), .A(n4958), .ZN(n4963) );
  OAI22_X1 U5477 ( .A1(IR_REG_13__SCAN_IN), .A2(keyinput_f68), .B1(
        IR_REG_6__SCAN_IN), .B2(keyinput_f61), .ZN(n4959) );
  AOI221_X1 U5478 ( .B1(IR_REG_13__SCAN_IN), .B2(keyinput_f68), .C1(
        keyinput_f61), .C2(IR_REG_6__SCAN_IN), .A(n4959), .ZN(n4962) );
  OAI22_X1 U5479 ( .A1(IR_REG_4__SCAN_IN), .A2(keyinput_f59), .B1(keyinput_f47), .B2(REG3_REG_5__SCAN_IN), .ZN(n4960) );
  AOI221_X1 U5480 ( .B1(IR_REG_4__SCAN_IN), .B2(keyinput_f59), .C1(
        REG3_REG_5__SCAN_IN), .C2(keyinput_f47), .A(n4960), .ZN(n4961) );
  NAND4_X1 U5481 ( .A1(n4964), .A2(n4963), .A3(n4962), .A4(n4961), .ZN(n4983)
         );
  OAI22_X1 U5482 ( .A1(IR_REG_3__SCAN_IN), .A2(keyinput_f58), .B1(DATAI_0_), 
        .B2(keyinput_f31), .ZN(n4965) );
  AOI221_X1 U5483 ( .B1(IR_REG_3__SCAN_IN), .B2(keyinput_f58), .C1(
        keyinput_f31), .C2(DATAI_0_), .A(n4965), .ZN(n4972) );
  OAI22_X1 U5484 ( .A1(IR_REG_2__SCAN_IN), .A2(keyinput_f57), .B1(
        keyinput_f119), .B2(REG0_REG_0__SCAN_IN), .ZN(n4966) );
  AOI221_X1 U5485 ( .B1(IR_REG_2__SCAN_IN), .B2(keyinput_f57), .C1(
        REG0_REG_0__SCAN_IN), .C2(keyinput_f119), .A(n4966), .ZN(n4971) );
  OAI22_X1 U5486 ( .A1(REG3_REG_9__SCAN_IN), .A2(keyinput_f51), .B1(
        keyinput_f127), .B2(REG0_REG_8__SCAN_IN), .ZN(n4967) );
  AOI221_X1 U5487 ( .B1(REG3_REG_9__SCAN_IN), .B2(keyinput_f51), .C1(
        REG0_REG_8__SCAN_IN), .C2(keyinput_f127), .A(n4967), .ZN(n4970) );
  OAI22_X1 U5488 ( .A1(D_REG_9__SCAN_IN), .A2(keyinput_f96), .B1(
        D_REG_3__SCAN_IN), .B2(keyinput_f90), .ZN(n4968) );
  AOI221_X1 U5489 ( .B1(D_REG_9__SCAN_IN), .B2(keyinput_f96), .C1(keyinput_f90), .C2(D_REG_3__SCAN_IN), .A(n4968), .ZN(n4969) );
  NAND4_X1 U5490 ( .A1(n4972), .A2(n4971), .A3(n4970), .A4(n4969), .ZN(n4982)
         );
  OAI22_X1 U5491 ( .A1(D_REG_21__SCAN_IN), .A2(keyinput_f108), .B1(
        D_REG_12__SCAN_IN), .B2(keyinput_f99), .ZN(n4973) );
  AOI221_X1 U5492 ( .B1(D_REG_21__SCAN_IN), .B2(keyinput_f108), .C1(
        keyinput_f99), .C2(D_REG_12__SCAN_IN), .A(n4973), .ZN(n4980) );
  OAI22_X1 U5493 ( .A1(D_REG_28__SCAN_IN), .A2(keyinput_f115), .B1(
        D_REG_31__SCAN_IN), .B2(keyinput_f118), .ZN(n4974) );
  AOI221_X1 U5494 ( .B1(D_REG_28__SCAN_IN), .B2(keyinput_f115), .C1(
        keyinput_f118), .C2(D_REG_31__SCAN_IN), .A(n4974), .ZN(n4979) );
  OAI22_X1 U5495 ( .A1(D_REG_2__SCAN_IN), .A2(keyinput_f89), .B1(
        D_REG_29__SCAN_IN), .B2(keyinput_f116), .ZN(n4975) );
  AOI221_X1 U5496 ( .B1(D_REG_2__SCAN_IN), .B2(keyinput_f89), .C1(
        keyinput_f116), .C2(D_REG_29__SCAN_IN), .A(n4975), .ZN(n4978) );
  OAI22_X1 U5497 ( .A1(D_REG_0__SCAN_IN), .A2(keyinput_f87), .B1(
        IR_REG_29__SCAN_IN), .B2(keyinput_f84), .ZN(n4976) );
  AOI221_X1 U5498 ( .B1(D_REG_0__SCAN_IN), .B2(keyinput_f87), .C1(keyinput_f84), .C2(IR_REG_29__SCAN_IN), .A(n4976), .ZN(n4977) );
  NAND4_X1 U5499 ( .A1(n4980), .A2(n4979), .A3(n4978), .A4(n4977), .ZN(n4981)
         );
  NOR4_X1 U5500 ( .A1(n4984), .A2(n4983), .A3(n4982), .A4(n4981), .ZN(n5131)
         );
  OAI22_X1 U5501 ( .A1(REG3_REG_21__SCAN_IN), .A2(keyinput_f43), .B1(
        REG3_REG_20__SCAN_IN), .B2(keyinput_f53), .ZN(n4985) );
  AOI221_X1 U5502 ( .B1(REG3_REG_21__SCAN_IN), .B2(keyinput_f43), .C1(
        keyinput_f53), .C2(REG3_REG_20__SCAN_IN), .A(n4985), .ZN(n4992) );
  OAI22_X1 U5503 ( .A1(DATAI_31_), .A2(keyinput_f0), .B1(DATAI_30_), .B2(
        keyinput_f1), .ZN(n4986) );
  AOI221_X1 U5504 ( .B1(DATAI_31_), .B2(keyinput_f0), .C1(keyinput_f1), .C2(
        DATAI_30_), .A(n4986), .ZN(n4991) );
  OAI22_X1 U5505 ( .A1(DATAI_29_), .A2(keyinput_f2), .B1(keyinput_f3), .B2(
        DATAI_28_), .ZN(n4987) );
  AOI221_X1 U5506 ( .B1(DATAI_29_), .B2(keyinput_f2), .C1(DATAI_28_), .C2(
        keyinput_f3), .A(n4987), .ZN(n4990) );
  OAI22_X1 U5507 ( .A1(REG3_REG_3__SCAN_IN), .A2(keyinput_f38), .B1(
        keyinput_f5), .B2(DATAI_26_), .ZN(n4988) );
  AOI221_X1 U5508 ( .B1(REG3_REG_3__SCAN_IN), .B2(keyinput_f38), .C1(DATAI_26_), .C2(keyinput_f5), .A(n4988), .ZN(n4989) );
  NAND4_X1 U5509 ( .A1(n4992), .A2(n4991), .A3(n4990), .A4(n4989), .ZN(n5129)
         );
  OAI22_X1 U5510 ( .A1(DATAI_3_), .A2(keyinput_f28), .B1(keyinput_f29), .B2(
        DATAI_2_), .ZN(n4993) );
  AOI221_X1 U5511 ( .B1(DATAI_3_), .B2(keyinput_f28), .C1(DATAI_2_), .C2(
        keyinput_f29), .A(n4993), .ZN(n5019) );
  OAI22_X1 U5512 ( .A1(REG3_REG_28__SCAN_IN), .A2(keyinput_f40), .B1(
        keyinput_f34), .B2(REG3_REG_27__SCAN_IN), .ZN(n4994) );
  AOI221_X1 U5513 ( .B1(REG3_REG_28__SCAN_IN), .B2(keyinput_f40), .C1(
        REG3_REG_27__SCAN_IN), .C2(keyinput_f34), .A(n4994), .ZN(n4997) );
  OAI22_X1 U5514 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput_f52), .B1(
        keyinput_f27), .B2(DATAI_4_), .ZN(n4995) );
  AOI221_X1 U5515 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput_f52), .C1(DATAI_4_), 
        .C2(keyinput_f27), .A(n4995), .ZN(n4996) );
  OAI211_X1 U5516 ( .C1(n4999), .C2(keyinput_f16), .A(n4997), .B(n4996), .ZN(
        n4998) );
  AOI21_X1 U5517 ( .B1(n4999), .B2(keyinput_f16), .A(n4998), .ZN(n5018) );
  AOI22_X1 U5518 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput_f42), .B1(
        REG3_REG_14__SCAN_IN), .B2(keyinput_f35), .ZN(n5000) );
  OAI221_X1 U5519 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput_f42), .C1(
        REG3_REG_14__SCAN_IN), .C2(keyinput_f35), .A(n5000), .ZN(n5007) );
  AOI22_X1 U5520 ( .A1(D_REG_25__SCAN_IN), .A2(keyinput_f112), .B1(
        D_REG_30__SCAN_IN), .B2(keyinput_f117), .ZN(n5001) );
  OAI221_X1 U5521 ( .B1(D_REG_25__SCAN_IN), .B2(keyinput_f112), .C1(
        D_REG_30__SCAN_IN), .C2(keyinput_f117), .A(n5001), .ZN(n5006) );
  AOI22_X1 U5522 ( .A1(D_REG_23__SCAN_IN), .A2(keyinput_f110), .B1(
        D_REG_24__SCAN_IN), .B2(keyinput_f111), .ZN(n5002) );
  OAI221_X1 U5523 ( .B1(D_REG_23__SCAN_IN), .B2(keyinput_f110), .C1(
        D_REG_24__SCAN_IN), .C2(keyinput_f111), .A(n5002), .ZN(n5005) );
  AOI22_X1 U5524 ( .A1(D_REG_14__SCAN_IN), .A2(keyinput_f101), .B1(
        D_REG_17__SCAN_IN), .B2(keyinput_f104), .ZN(n5003) );
  OAI221_X1 U5525 ( .B1(D_REG_14__SCAN_IN), .B2(keyinput_f101), .C1(
        D_REG_17__SCAN_IN), .C2(keyinput_f104), .A(n5003), .ZN(n5004) );
  NOR4_X1 U5526 ( .A1(n5007), .A2(n5006), .A3(n5005), .A4(n5004), .ZN(n5017)
         );
  AOI22_X1 U5527 ( .A1(IR_REG_30__SCAN_IN), .A2(keyinput_f85), .B1(
        D_REG_11__SCAN_IN), .B2(keyinput_f98), .ZN(n5008) );
  OAI221_X1 U5528 ( .B1(IR_REG_30__SCAN_IN), .B2(keyinput_f85), .C1(
        D_REG_11__SCAN_IN), .C2(keyinput_f98), .A(n5008), .ZN(n5015) );
  AOI22_X1 U5529 ( .A1(IR_REG_17__SCAN_IN), .A2(keyinput_f72), .B1(
        IR_REG_31__SCAN_IN), .B2(keyinput_f86), .ZN(n5009) );
  OAI221_X1 U5530 ( .B1(IR_REG_17__SCAN_IN), .B2(keyinput_f72), .C1(
        IR_REG_31__SCAN_IN), .C2(keyinput_f86), .A(n5009), .ZN(n5014) );
  AOI22_X1 U5531 ( .A1(DATAI_16_), .A2(keyinput_f15), .B1(IR_REG_14__SCAN_IN), 
        .B2(keyinput_f69), .ZN(n5010) );
  OAI221_X1 U5532 ( .B1(DATAI_16_), .B2(keyinput_f15), .C1(IR_REG_14__SCAN_IN), 
        .C2(keyinput_f69), .A(n5010), .ZN(n5013) );
  AOI22_X1 U5533 ( .A1(DATAI_13_), .A2(keyinput_f18), .B1(DATAI_14_), .B2(
        keyinput_f17), .ZN(n5011) );
  OAI221_X1 U5534 ( .B1(DATAI_13_), .B2(keyinput_f18), .C1(DATAI_14_), .C2(
        keyinput_f17), .A(n5011), .ZN(n5012) );
  NOR4_X1 U5535 ( .A1(n5015), .A2(n5014), .A3(n5013), .A4(n5012), .ZN(n5016)
         );
  NAND4_X1 U5536 ( .A1(n5019), .A2(n5018), .A3(n5017), .A4(n5016), .ZN(n5128)
         );
  AOI22_X1 U5537 ( .A1(DATAI_1_), .A2(keyinput_f30), .B1(IR_REG_26__SCAN_IN), 
        .B2(keyinput_f81), .ZN(n5020) );
  OAI221_X1 U5538 ( .B1(DATAI_1_), .B2(keyinput_f30), .C1(IR_REG_26__SCAN_IN), 
        .C2(keyinput_f81), .A(n5020), .ZN(n5027) );
  AOI22_X1 U5539 ( .A1(REG0_REG_2__SCAN_IN), .A2(keyinput_f121), .B1(
        IR_REG_21__SCAN_IN), .B2(keyinput_f76), .ZN(n5021) );
  OAI221_X1 U5540 ( .B1(REG0_REG_2__SCAN_IN), .B2(keyinput_f121), .C1(
        IR_REG_21__SCAN_IN), .C2(keyinput_f76), .A(n5021), .ZN(n5026) );
  AOI22_X1 U5541 ( .A1(DATAI_25_), .A2(keyinput_f6), .B1(IR_REG_10__SCAN_IN), 
        .B2(keyinput_f65), .ZN(n5022) );
  OAI221_X1 U5542 ( .B1(DATAI_25_), .B2(keyinput_f6), .C1(IR_REG_10__SCAN_IN), 
        .C2(keyinput_f65), .A(n5022), .ZN(n5025) );
  AOI22_X1 U5543 ( .A1(DATAI_24_), .A2(keyinput_f7), .B1(DATAI_19_), .B2(
        keyinput_f12), .ZN(n5023) );
  OAI221_X1 U5544 ( .B1(DATAI_24_), .B2(keyinput_f7), .C1(DATAI_19_), .C2(
        keyinput_f12), .A(n5023), .ZN(n5024) );
  NOR4_X1 U5545 ( .A1(n5027), .A2(n5026), .A3(n5025), .A4(n5024), .ZN(n5069)
         );
  AOI22_X1 U5546 ( .A1(DATAI_18_), .A2(keyinput_f13), .B1(IR_REG_28__SCAN_IN), 
        .B2(keyinput_f83), .ZN(n5028) );
  OAI221_X1 U5547 ( .B1(DATAI_18_), .B2(keyinput_f13), .C1(IR_REG_28__SCAN_IN), 
        .C2(keyinput_f83), .A(n5028), .ZN(n5037) );
  AOI22_X1 U5548 ( .A1(DATAI_22_), .A2(keyinput_f9), .B1(REG3_REG_8__SCAN_IN), 
        .B2(keyinput_f41), .ZN(n5029) );
  OAI221_X1 U5549 ( .B1(DATAI_22_), .B2(keyinput_f9), .C1(REG3_REG_8__SCAN_IN), 
        .C2(keyinput_f41), .A(n5029), .ZN(n5036) );
  AOI22_X1 U5550 ( .A1(REG3_REG_10__SCAN_IN), .A2(keyinput_f37), .B1(
        IR_REG_25__SCAN_IN), .B2(keyinput_f80), .ZN(n5030) );
  OAI221_X1 U5551 ( .B1(REG3_REG_10__SCAN_IN), .B2(keyinput_f37), .C1(
        IR_REG_25__SCAN_IN), .C2(keyinput_f80), .A(n5030), .ZN(n5035) );
  AOI22_X1 U5552 ( .A1(n5033), .A2(keyinput_f49), .B1(keyinput_f10), .B2(n5032), .ZN(n5031) );
  OAI221_X1 U5553 ( .B1(n5033), .B2(keyinput_f49), .C1(n5032), .C2(
        keyinput_f10), .A(n5031), .ZN(n5034) );
  NOR4_X1 U5554 ( .A1(n5037), .A2(n5036), .A3(n5035), .A4(n5034), .ZN(n5068)
         );
  AOI22_X1 U5555 ( .A1(n2602), .A2(keyinput_f54), .B1(keyinput_f33), .B2(n5039), .ZN(n5038) );
  OAI221_X1 U5556 ( .B1(n2602), .B2(keyinput_f54), .C1(n5039), .C2(
        keyinput_f33), .A(n5038), .ZN(n5050) );
  AOI22_X1 U5557 ( .A1(n5042), .A2(keyinput_f71), .B1(keyinput_f70), .B2(n5040), .ZN(n5041) );
  OAI221_X1 U5558 ( .B1(n5042), .B2(keyinput_f71), .C1(n5040), .C2(
        keyinput_f70), .A(n5041), .ZN(n5049) );
  XOR2_X1 U5559 ( .A(n2289), .B(keyinput_f55), .Z(n5047) );
  XOR2_X1 U5560 ( .A(n5043), .B(keyinput_f120), .Z(n5046) );
  XNOR2_X1 U5561 ( .A(IR_REG_27__SCAN_IN), .B(keyinput_f82), .ZN(n5045) );
  XNOR2_X1 U5562 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_f50), .ZN(n5044) );
  NAND4_X1 U5563 ( .A1(n5047), .A2(n5046), .A3(n5045), .A4(n5044), .ZN(n5048)
         );
  NOR3_X1 U5564 ( .A1(n5050), .A2(n5049), .A3(n5048), .ZN(n5067) );
  AOI22_X1 U5565 ( .A1(n5053), .A2(keyinput_f91), .B1(keyinput_f95), .B2(n5052), .ZN(n5051) );
  OAI221_X1 U5566 ( .B1(n5053), .B2(keyinput_f91), .C1(n5052), .C2(
        keyinput_f95), .A(n5051), .ZN(n5065) );
  AOI22_X1 U5567 ( .A1(n5056), .A2(keyinput_f109), .B1(keyinput_f113), .B2(
        n5055), .ZN(n5054) );
  OAI221_X1 U5568 ( .B1(n5056), .B2(keyinput_f109), .C1(n5055), .C2(
        keyinput_f113), .A(n5054), .ZN(n5064) );
  XOR2_X1 U5569 ( .A(n5057), .B(keyinput_f56), .Z(n5060) );
  XNOR2_X1 U5570 ( .A(IR_REG_7__SCAN_IN), .B(keyinput_f62), .ZN(n5059) );
  XNOR2_X1 U5571 ( .A(IR_REG_18__SCAN_IN), .B(keyinput_f73), .ZN(n5058) );
  NAND3_X1 U5572 ( .A1(n5060), .A2(n5059), .A3(n5058), .ZN(n5063) );
  XNOR2_X1 U5573 ( .A(n5061), .B(keyinput_f93), .ZN(n5062) );
  NOR4_X1 U5574 ( .A1(n5065), .A2(n5064), .A3(n5063), .A4(n5062), .ZN(n5066)
         );
  NAND4_X1 U5575 ( .A1(n5069), .A2(n5068), .A3(n5067), .A4(n5066), .ZN(n5127)
         );
  AOI22_X1 U5576 ( .A1(n5072), .A2(keyinput_f97), .B1(keyinput_f107), .B2(
        n5071), .ZN(n5070) );
  OAI221_X1 U5577 ( .B1(n5072), .B2(keyinput_f97), .C1(n5071), .C2(
        keyinput_f107), .A(n5070), .ZN(n5085) );
  AOI22_X1 U5578 ( .A1(n5075), .A2(keyinput_f100), .B1(keyinput_f103), .B2(
        n5074), .ZN(n5073) );
  OAI221_X1 U5579 ( .B1(n5075), .B2(keyinput_f100), .C1(n5074), .C2(
        keyinput_f103), .A(n5073), .ZN(n5084) );
  AOI22_X1 U5580 ( .A1(n5078), .A2(keyinput_f105), .B1(keyinput_f106), .B2(
        n5077), .ZN(n5076) );
  OAI221_X1 U5581 ( .B1(n5078), .B2(keyinput_f105), .C1(n5077), .C2(
        keyinput_f106), .A(n5076), .ZN(n5083) );
  AOI22_X1 U5582 ( .A1(n5081), .A2(keyinput_f102), .B1(keyinput_f92), .B2(
        n5080), .ZN(n5079) );
  OAI221_X1 U5583 ( .B1(n5081), .B2(keyinput_f102), .C1(n5080), .C2(
        keyinput_f92), .A(n5079), .ZN(n5082) );
  NOR4_X1 U5584 ( .A1(n5085), .A2(n5084), .A3(n5083), .A4(n5082), .ZN(n5125)
         );
  AOI22_X1 U5585 ( .A1(n5088), .A2(keyinput_f94), .B1(keyinput_f114), .B2(
        n5087), .ZN(n5086) );
  OAI221_X1 U5586 ( .B1(n5088), .B2(keyinput_f94), .C1(n5087), .C2(
        keyinput_f114), .A(n5086), .ZN(n5097) );
  INV_X1 U5587 ( .A(REG3_REG_19__SCAN_IN), .ZN(n5090) );
  AOI22_X1 U5588 ( .A1(n2645), .A2(keyinput_f48), .B1(n5090), .B2(keyinput_f39), .ZN(n5089) );
  OAI221_X1 U5589 ( .B1(n2645), .B2(keyinput_f48), .C1(n5090), .C2(
        keyinput_f39), .A(n5089), .ZN(n5096) );
  XNOR2_X1 U5590 ( .A(REG3_REG_25__SCAN_IN), .B(keyinput_f45), .ZN(n5094) );
  XNOR2_X1 U5591 ( .A(IR_REG_12__SCAN_IN), .B(keyinput_f67), .ZN(n5093) );
  XNOR2_X1 U5592 ( .A(IR_REG_9__SCAN_IN), .B(keyinput_f64), .ZN(n5092) );
  XNOR2_X1 U5593 ( .A(REG3_REG_23__SCAN_IN), .B(keyinput_f36), .ZN(n5091) );
  NAND4_X1 U5594 ( .A1(n5094), .A2(n5093), .A3(n5092), .A4(n5091), .ZN(n5095)
         );
  NOR3_X1 U5595 ( .A1(n5097), .A2(n5096), .A3(n5095), .ZN(n5124) );
  AOI22_X1 U5596 ( .A1(n5099), .A2(keyinput_f4), .B1(keyinput_f14), .B2(n2659), 
        .ZN(n5098) );
  OAI221_X1 U5597 ( .B1(n5099), .B2(keyinput_f4), .C1(n2659), .C2(keyinput_f14), .A(n5098), .ZN(n5109) );
  AOI22_X1 U5598 ( .A1(n5102), .A2(keyinput_f21), .B1(n5101), .B2(keyinput_f11), .ZN(n5100) );
  OAI221_X1 U5599 ( .B1(n5102), .B2(keyinput_f21), .C1(n5101), .C2(
        keyinput_f11), .A(n5100), .ZN(n5108) );
  XNOR2_X1 U5600 ( .A(REG3_REG_16__SCAN_IN), .B(keyinput_f46), .ZN(n5106) );
  XNOR2_X1 U5601 ( .A(IR_REG_23__SCAN_IN), .B(keyinput_f78), .ZN(n5105) );
  XNOR2_X1 U5602 ( .A(IR_REG_22__SCAN_IN), .B(keyinput_f77), .ZN(n5104) );
  XNOR2_X1 U5603 ( .A(REG3_REG_12__SCAN_IN), .B(keyinput_f44), .ZN(n5103) );
  NAND4_X1 U5604 ( .A1(n5106), .A2(n5105), .A3(n5104), .A4(n5103), .ZN(n5107)
         );
  NOR3_X1 U5605 ( .A1(n5109), .A2(n5108), .A3(n5107), .ZN(n5123) );
  XOR2_X1 U5606 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_f63), .Z(n5111) );
  XOR2_X1 U5607 ( .A(DATAI_6_), .B(keyinput_f25), .Z(n5110) );
  NOR2_X1 U5608 ( .A1(n5111), .A2(n5110), .ZN(n5115) );
  XNOR2_X1 U5609 ( .A(keyinput_f75), .B(IR_REG_20__SCAN_IN), .ZN(n5114) );
  XNOR2_X1 U5610 ( .A(IR_REG_24__SCAN_IN), .B(keyinput_f79), .ZN(n5113) );
  XNOR2_X1 U5611 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_f60), .ZN(n5112) );
  NAND4_X1 U5612 ( .A1(n5115), .A2(n5114), .A3(n5113), .A4(n5112), .ZN(n5121)
         );
  AOI22_X1 U5613 ( .A1(n2741), .A2(keyinput_f74), .B1(keyinput_f8), .B2(n5117), 
        .ZN(n5116) );
  OAI221_X1 U5614 ( .B1(n2741), .B2(keyinput_f74), .C1(n5117), .C2(keyinput_f8), .A(n5116), .ZN(n5120) );
  XNOR2_X1 U5615 ( .A(n5118), .B(keyinput_f88), .ZN(n5119) );
  NOR3_X1 U5616 ( .A1(n5121), .A2(n5120), .A3(n5119), .ZN(n5122) );
  NAND4_X1 U5617 ( .A1(n5125), .A2(n5124), .A3(n5123), .A4(n5122), .ZN(n5126)
         );
  NOR4_X1 U5618 ( .A1(n5129), .A2(n5128), .A3(n5127), .A4(n5126), .ZN(n5130)
         );
  NAND2_X1 U5619 ( .A1(n5131), .A2(n5130), .ZN(n5133) );
  AOI21_X1 U5620 ( .B1(keyinput_f32), .B2(n5133), .A(keyinput_g32), .ZN(n5135)
         );
  INV_X1 U5621 ( .A(keyinput_f32), .ZN(n5132) );
  AOI21_X1 U5622 ( .B1(n5133), .B2(n5132), .A(U3149), .ZN(n5134) );
  AOI22_X1 U5623 ( .A1(U3149), .A2(n5135), .B1(keyinput_g32), .B2(n5134), .ZN(
        n5136) );
  AOI21_X1 U5624 ( .B1(n5138), .B2(n5137), .A(n5136), .ZN(n5140) );
  AOI22_X1 U5625 ( .A1(STATE_REG_SCAN_IN), .A2(IR_REG_0__SCAN_IN), .B1(
        DATAI_0_), .B2(U3149), .ZN(n5139) );
  XNOR2_X1 U5626 ( .A(n5140), .B(n5139), .ZN(U3352) );
  AND2_X1 U2484 ( .A1(n3161), .A2(n2242), .ZN(n4738) );
endmodule

