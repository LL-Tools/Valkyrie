

module b17_C_SARLock_k_64_1 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, U355, U356, U357, U358, 
        U359, U360, U361, U362, U363, U364, U366, U367, U368, U369, U370, U371, 
        U372, U373, U374, U375, U347, U348, U349, U350, U351, U352, U353, U354, 
        U365, U376, U247, U246, U245, U244, U243, U242, U241, U240, U239, U238, 
        U237, U236, U235, U234, U233, U232, U231, U230, U229, U228, U227, U226, 
        U225, U224, U223, U222, U221, U220, U219, U218, U217, U216, U251, U252, 
        U253, U254, U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, 
        U265, U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276, 
        U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274, 
        P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, 
        P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, 
        P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, 
        P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, 
        P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, 
        P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, 
        P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, 
        P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, 
        P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, 
        P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, 
        P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, 
        P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, 
        P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, 
        P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, 
        P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, 
        P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, 
        P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, 
        P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, 
        P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, 
        P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, 
        P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, 
        P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, 
        P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, 
        P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, 
        P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, 
        P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, 
        P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, 
        P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, 
        P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, 
        P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, 
        P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, 
        P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, 
        P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, 
        P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, 
        P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, 
        P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, 
        P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, 
        P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, 
        P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, 
        P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, 
        P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, 
        P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, 
        P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, 
        P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, 
        P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, 
        P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, 
        P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, 
        P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, 
        P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, 
        P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, 
        P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, 
        P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, 
        P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, 
        P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, 
        P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, 
        P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, 
        P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, 
        P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, 
        P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, 
        P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, 
        P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, 
        P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, 
        P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, 
        P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, 
        P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, 
        P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, 
        P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, 
        P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, 
        P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, 
        P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, 
        P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, 
        P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, 
        P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, 
        P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, 
        P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, 
        P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, 
        P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, 
        P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, 
        P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, 
        P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, 
        P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, 
        P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, 
        P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, 
        P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, 
        P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, 
        P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, 
        P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, 
        P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, 
        P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, 
        P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, 
        P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, 
        P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, 
        P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, 
        P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, 
        P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, 
        P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, 
        P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, 
        P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, 
        P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, 
        P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, 
        P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, 
        P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, 
        P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, 
        P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, 
        P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, 
        P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, 
        P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, 
        P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, 
        P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, 
        P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, 
        P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, 
        P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, 
        P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, 
        P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, 
        P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, 
        P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, 
        P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, 
        P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, 
        P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, 
        P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, 
        P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, 
        P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, 
        P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, 
        P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, 
        P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, 
        P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, 
        P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, 
        P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, 
        P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, 
        P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, 
        P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, 
        P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, 
        P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, 
        P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, 
        P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, 
        P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, 
        P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, 
        P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, 
        P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, 
        P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, 
        P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, 
        P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, 
        P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, 
        P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, 
        P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, 
        P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, 
        P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, 
        P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, 
        P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, 
        P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, 
        P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, 
        P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, 
        P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, 
        P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, 
        P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, 
        P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, 
        P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, 
        P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, 
        P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, 
        P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, 
        P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, 
        P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, 
        P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, 
        P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, 
        P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, 
        P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, 
        P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, 
        P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, 
        P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, 
        P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, 
        P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, 
        P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, 
        P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, 
        P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, 
        P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, 
        P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, 
        P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, 
        P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, 
        P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, 
        P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, 
        P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, 
        P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, 
        P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, 
        P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, 
        P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, 
        P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, 
        P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, 
        P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, 
        P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, 
        P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, 
        P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, 
        P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, 
        P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9591, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
         n9602, n9603, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13960, n13961, n13962, n13963, n13964,
         n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972,
         n13973, n13974, n13975, n13976, n13977, n13978, n13979, n13980,
         n13981, n13982, n13983, n13984, n13985, n13986, n13987, n13988,
         n13989, n13990, n13991, n13992, n13993, n13994, n13995, n13996,
         n13997, n13998, n13999, n14000, n14001, n14002, n14003, n14004,
         n14005, n14006, n14007, n14008, n14009, n14010, n14011, n14012,
         n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14020,
         n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028,
         n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
         n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044,
         n14045, n14046, n14047, n14048, n14049, n14050, n14051, n14052,
         n14053, n14054, n14055, n14056, n14057, n14058, n14059, n14060,
         n14061, n14062, n14063, n14064, n14065, n14066, n14067, n14068,
         n14069, n14070, n14071, n14072, n14073, n14074, n14075, n14076,
         n14077, n14078, n14079, n14080, n14081, n14082, n14083, n14084,
         n14085, n14086, n14087, n14088, n14089, n14090, n14091, n14092,
         n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100,
         n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
         n14109, n14110, n14111, n14112, n14113, n14114, n14115, n14116,
         n14117, n14118, n14119, n14120, n14121, n14122, n14123, n14124,
         n14125, n14126, n14127, n14128, n14129, n14130, n14131, n14132,
         n14133, n14134, n14135, n14136, n14137, n14138, n14139, n14140,
         n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148,
         n14149, n14150, n14151, n14152, n14153, n14154, n14155, n14156,
         n14157, n14158, n14159, n14160, n14161, n14162, n14163, n14164,
         n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
         n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180,
         n14181, n14182, n14183, n14184, n14185, n14186, n14187, n14188,
         n14189, n14190, n14191, n14192, n14193, n14194, n14195, n14196,
         n14197, n14198, n14199, n14200, n14201, n14202, n14203, n14204,
         n14205, n14206, n14207, n14208, n14209, n14210, n14211, n14212,
         n14213, n14214, n14215, n14216, n14217, n14218, n14219, n14220,
         n14221, n14222, n14223, n14224, n14225, n14226, n14227, n14228,
         n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
         n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244,
         n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252,
         n14253, n14254, n14255, n14256, n14257, n14258, n14259, n14260,
         n14261, n14262, n14263, n14264, n14265, n14266, n14267, n14268,
         n14269, n14270, n14271, n14272, n14273, n14274, n14275, n14276,
         n14277, n14278, n14279, n14280, n14281, n14282, n14283, n14284,
         n14285, n14286, n14287, n14288, n14289, n14290, n14291, n14292,
         n14293, n14294, n14295, n14296, n14297, n14298, n14299, n14300,
         n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
         n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316,
         n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324,
         n14325, n14326, n14327, n14328, n14329, n14330, n14331, n14332,
         n14333, n14334, n14335, n14336, n14337, n14338, n14339, n14340,
         n14341, n14342, n14343, n14344, n14345, n14346, n14347, n14348,
         n14349, n14350, n14351, n14352, n14353, n14354, n14355, n14356,
         n14357, n14358, n14359, n14360, n14361, n14362, n14363, n14364,
         n14365, n14366, n14367, n14368, n14369, n14370, n14371, n14372,
         n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
         n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388,
         n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396,
         n14397, n14398, n14399, n14400, n14401, n14402, n14403, n14404,
         n14405, n14406, n14407, n14408, n14409, n14410, n14411, n14412,
         n14413, n14414, n14415, n14416, n14417, n14418, n14419, n14420,
         n14421, n14422, n14423, n14424, n14425, n14426, n14427, n14428,
         n14429, n14430, n14431, n14432, n14433, n14434, n14435, n14436,
         n14437, n14438, n14439, n14440, n14441, n14442, n14443, n14444,
         n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
         n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460,
         n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468,
         n14469, n14470, n14471, n14472, n14473, n14474, n14475, n14476,
         n14477, n14478, n14479, n14480, n14481, n14482, n14483, n14484,
         n14485, n14486, n14487, n14488, n14489, n14490, n14491, n14492,
         n14493, n14494, n14495, n14496, n14497, n14498, n14499, n14500,
         n14501, n14502, n14503, n14504, n14505, n14506, n14507, n14508,
         n14509, n14510, n14511, n14512, n14513, n14514, n14515, n14516,
         n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
         n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532,
         n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540,
         n14541, n14542, n14543, n14544, n14545, n14546, n14547, n14548,
         n14549, n14550, n14551, n14552, n14553, n14554, n14555, n14556,
         n14557, n14558, n14559, n14560, n14561, n14562, n14563, n14564,
         n14565, n14566, n14567, n14568, n14569, n14570, n14571, n14572,
         n14573, n14574, n14575, n14576, n14577, n14578, n14579, n14580,
         n14581, n14582, n14583, n14584, n14585, n14586, n14587, n14588,
         n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
         n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604,
         n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612,
         n14613, n14614, n14615, n14616, n14617, n14618, n14619, n14620,
         n14621, n14622, n14623, n14624, n14625, n14626, n14627, n14628,
         n14629, n14630, n14631, n14632, n14633, n14634, n14635, n14636,
         n14637, n14638, n14639, n14640, n14641, n14642, n14643, n14644,
         n14645, n14646, n14647, n14648, n14649, n14650, n14651, n14652,
         n14653, n14654, n14655, n14656, n14657, n14658, n14659, n14660,
         n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
         n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676,
         n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684,
         n14685, n14686, n14687, n14688, n14689, n14690, n14691, n14692,
         n14693, n14694, n14695, n14696, n14697, n14698, n14699, n14700,
         n14701, n14702, n14703, n14704, n14705, n14706, n14707, n14708,
         n14709, n14710, n14711, n14712, n14713, n14714, n14715, n14716,
         n14717, n14718, n14719, n14720, n14721, n14722, n14723, n14724,
         n14725, n14726, n14727, n14728, n14729, n14730, n14731, n14732,
         n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
         n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748,
         n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756,
         n14757, n14758, n14759, n14760, n14761, n14762, n14763, n14764,
         n14765, n14766, n14767, n14768, n14769, n14770, n14771, n14772,
         n14773, n14774, n14775, n14776, n14777, n14778, n14779, n14780,
         n14781, n14782, n14783, n14784, n14785, n14786, n14787, n14788,
         n14789, n14790, n14791, n14792, n14793, n14794, n14795, n14796,
         n14797, n14798, n14799, n14800, n14801, n14802, n14803, n14804,
         n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
         n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820,
         n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828,
         n14829, n14830, n14831, n14832, n14833, n14834, n14835, n14836,
         n14837, n14838, n14839, n14840, n14841, n14842, n14843, n14844,
         n14845, n14846, n14847, n14848, n14849, n14850, n14851, n14852,
         n14853, n14854, n14855, n14856, n14857, n14858, n14859, n14860,
         n14861, n14862, n14863, n14864, n14865, n14866, n14867, n14868,
         n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
         n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884,
         n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892,
         n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900,
         n14901, n14902, n14903, n14904, n14905, n14906, n14907, n14908,
         n14909, n14910, n14911, n14912, n14913, n14914, n14915, n14916,
         n14917, n14918, n14919, n14920, n14921, n14922, n14923, n14924,
         n14925, n14926, n14927, n14928, n14929, n14930, n14931, n14932,
         n14933, n14934, n14935, n14936, n14937, n14938, n14939, n14940,
         n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
         n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956,
         n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964,
         n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972,
         n14973, n14974, n14975, n14976, n14977, n14978, n14979, n14980,
         n14981, n14982, n14983, n14984, n14985, n14986, n14987, n14988,
         n14989, n14990, n14991, n14992, n14993, n14994, n14995, n14996,
         n14997, n14998, n14999, n15000, n15001, n15002, n15003, n15004,
         n15005, n15006, n15007, n15008, n15009, n15010, n15011, n15012,
         n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
         n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028,
         n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036,
         n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044,
         n15045, n15046, n15047, n15048, n15049, n15050, n15051, n15052,
         n15053, n15054, n15055, n15056, n15057, n15058, n15059, n15060,
         n15061, n15062, n15063, n15064, n15065, n15066, n15067, n15068,
         n15069, n15070, n15071, n15072, n15073, n15074, n15075, n15076,
         n15077, n15078, n15079, n15080, n15081, n15082, n15083, n15084,
         n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
         n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100,
         n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108,
         n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116,
         n15117, n15118, n15119, n15120, n15121, n15122, n15123, n15124,
         n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132,
         n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140,
         n15141, n15142, n15143, n15144, n15145, n15146, n15147, n15148,
         n15149, n15150, n15151, n15152, n15153, n15154, n15155, n15156,
         n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
         n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172,
         n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180,
         n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188,
         n15189, n15190, n15191, n15192, n15193, n15194, n15195, n15196,
         n15197, n15198, n15199, n15200, n15201, n15202, n15203, n15204,
         n15205, n15206, n15207, n15208, n15209, n15210, n15211, n15212,
         n15213, n15214, n15215, n15216, n15217, n15218, n15219, n15220,
         n15221, n15222, n15223, n15224, n15225, n15226, n15227, n15228,
         n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
         n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244,
         n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252,
         n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260,
         n15261, n15262, n15263, n15264, n15265, n15266, n15267, n15268,
         n15269, n15270, n15271, n15272, n15273, n15274, n15275, n15276,
         n15277, n15278, n15279, n15280, n15281, n15282, n15283, n15284,
         n15285, n15286, n15287, n15288, n15289, n15290, n15291, n15292,
         n15293, n15294, n15295, n15296, n15297, n15298, n15299, n15300,
         n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
         n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316,
         n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324,
         n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332,
         n15333, n15334, n15335, n15336, n15337, n15338, n15339, n15340,
         n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
         n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356,
         n15357, n15358, n15359, n15360, n15361, n15362, n15363, n15364,
         n15365, n15366, n15367, n15368, n15369, n15370, n15371, n15372,
         n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
         n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388,
         n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396,
         n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404,
         n15405, n15406, n15407, n15408, n15409, n15410, n15411, n15412,
         n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
         n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428,
         n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15436,
         n15437, n15438, n15439, n15440, n15441, n15442, n15443, n15444,
         n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
         n15453, n15454, n15455, n15456, n15457, n15458, n15459, n15460,
         n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468,
         n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476,
         n15477, n15478, n15479, n15480, n15481, n15482, n15483, n15484,
         n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
         n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500,
         n15501, n15502, n15503, n15504, n15505, n15506, n15507, n15508,
         n15509, n15510, n15511, n15512, n15513, n15514, n15515, n15516,
         n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524,
         n15525, n15526, n15527, n15528, n15529, n15530, n15531, n15532,
         n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540,
         n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548,
         n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
         n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
         n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572,
         n15573, n15574, n15575, n15576, n15577, n15578, n15579, n15580,
         n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588,
         n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596,
         n15597, n15598, n15599, n15600, n15601, n15602, n15603, n15604,
         n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612,
         n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620,
         n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
         n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
         n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644,
         n15645, n15646, n15647, n15648, n15649, n15650, n15651, n15652,
         n15653, n15654, n15655, n15656, n15657, n15658, n15659, n15660,
         n15661, n15662, n15663, n15664, n15665, n15666, n15667, n15668,
         n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676,
         n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684,
         n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692,
         n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
         n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
         n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716,
         n15717, n15718, n15719, n15720, n15721, n15722, n15723, n15724,
         n15725, n15726, n15727, n15728, n15729, n15730, n15731, n15732,
         n15733, n15734, n15735, n15736, n15737, n15738, n15739, n15740,
         n15741, n15742, n15743, n15744, n15745, n15746, n15747, n15748,
         n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
         n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764,
         n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
         n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780,
         n15781, n15782, n15783, n15784, n15785, n15786, n15787, n15788,
         n15789, n15790, n15791, n15792, n15793, n15794, n15795, n15796,
         n15797, n15798, n15799, n15800, n15801, n15802, n15803, n15804,
         n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812,
         n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820,
         n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828,
         n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836,
         n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
         n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852,
         n15853, n15854, n15855, n15856, n15857, n15858, n15859, n15860,
         n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868,
         n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876,
         n15877, n15878, n15879, n15880, n15881, n15882, n15883, n15884,
         n15885, n15886, n15887, n15888, n15889, n15890, n15891, n15892,
         n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900,
         n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908,
         n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
         n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924,
         n15925, n15926, n15927, n15928, n15929, n15930, n15931, n15932,
         n15933, n15934, n15935, n15936, n15937, n15938, n15939, n15940,
         n15941, n15942, n15943, n15944, n15945, n15946, n15947, n15948,
         n15949, n15950, n15951, n15952, n15953, n15954, n15955, n15956,
         n15957, n15958, n15959, n15960, n15961, n15962, n15963, n15964,
         n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972,
         n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980,
         n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
         n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996,
         n15997, n15998, n15999, n16000, n16001, n16002, n16003, n16004,
         n16005, n16006, n16007, n16008, n16009, n16010, n16011, n16012,
         n16013, n16014, n16015, n16016, n16017, n16018, n16019, n16020,
         n16021, n16022, n16023, n16024, n16025, n16026, n16027, n16028,
         n16029, n16030, n16031, n16032, n16033, n16034, n16035, n16036,
         n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044,
         n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052,
         n16053, n16054, n16055, n16056, n16057, n16058, n16059, n16060,
         n16061, n16062, n16063, n16064, n16065, n16066, n16067, n16068,
         n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076,
         n16077, n16078, n16079, n16080, n16081, n16082, n16083, n16084,
         n16085, n16086, n16087, n16088, n16089, n16090, n16091, n16092,
         n16093, n16094, n16095, n16096, n16097, n16098, n16099, n16100,
         n16101, n16102, n16103, n16104, n16105, n16106, n16107, n16108,
         n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
         n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124,
         n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132,
         n16133, n16134, n16135, n16136, n16137, n16138, n16139, n16140,
         n16141, n16142, n16143, n16144, n16145, n16146, n16147, n16148,
         n16149, n16150, n16151, n16152, n16153, n16154, n16155, n16156,
         n16157, n16158, n16159, n16160, n16161, n16162, n16163, n16164,
         n16165, n16166, n16167, n16168, n16169, n16170, n16171, n16172,
         n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180,
         n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188,
         n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196,
         n16197, n16198, n16199, n16200, n16201, n16202, n16203, n16204,
         n16205, n16206, n16207, n16208, n16209, n16210, n16211, n16212,
         n16213, n16214, n16215, n16216, n16217, n16218, n16219, n16220,
         n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228,
         n16229, n16230, n16231, n16232, n16233, n16234, n16235, n16236,
         n16237, n16238, n16239, n16240, n16241, n16242, n16243, n16244,
         n16245, n16246, n16247, n16248, n16249, n16250, n16251, n16252,
         n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260,
         n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
         n16269, n16270, n16271, n16272, n16273, n16274, n16275, n16276,
         n16277, n16278, n16279, n16280, n16281, n16282, n16283, n16284,
         n16285, n16286, n16287, n16288, n16289, n16290, n16291, n16292,
         n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300,
         n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16308,
         n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316,
         n16317, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
         n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332,
         n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340,
         n16341, n16342, n16343, n16344, n16345, n16346, n16347, n16348,
         n16349, n16350, n16351, n16352, n16353, n16354, n16355, n16356,
         n16357, n16358, n16359, n16360, n16361, n16362, n16363, n16364,
         n16365, n16366, n16367, n16368, n16369, n16370, n16371, n16372,
         n16373, n16374, n16375, n16376, n16377, n16378, n16379, n16380,
         n16381, n16382, n16383, n16384, n16385, n16386, n16387, n16388,
         n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396,
         n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404,
         n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412,
         n16413, n16414, n16415, n16416, n16417, n16418, n16419, n16420,
         n16421, n16422, n16423, n16424, n16425, n16426, n16427, n16428,
         n16429, n16430, n16431, n16432, n16433, n16434, n16435, n16436,
         n16437, n16438, n16439, n16440, n16441, n16442, n16443, n16444,
         n16445, n16446, n16447, n16448, n16449, n16450, n16451, n16452,
         n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
         n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468,
         n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476,
         n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484,
         n16485, n16486, n16487, n16488, n16489, n16490, n16491, n16492,
         n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
         n16501, n16502, n16503, n16504, n16505, n16506, n16507, n16508,
         n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516,
         n16517, n16518, n16519, n16520, n16521, n16522, n16523, n16524,
         n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
         n16533, n16534, n16535, n16536, n16537, n16538, n16539, n16540,
         n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548,
         n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556,
         n16557, n16558, n16559, n16560, n16561, n16562, n16563, n16564,
         n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572,
         n16573, n16574, n16575, n16576, n16577, n16578, n16579, n16580,
         n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
         n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596,
         n16597, n16598, n16599, n16600, n16601, n16602, n16603, n16604,
         n16605, n16606, n16607, n16608, n16609, n16610, n16611, n16612,
         n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620,
         n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628,
         n16629, n16630, n16631, n16632, n16633, n16634, n16635, n16636,
         n16637, n16638, n16639, n16640, n16641, n16642, n16643, n16644,
         n16645, n16646, n16647, n16648, n16649, n16650, n16651, n16652,
         n16653, n16654, n16655, n16656, n16657, n16658, n16659, n16660,
         n16661, n16662, n16663, n16664, n16665, n16666, n16667, n16668,
         n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
         n16677, n16678, n16679, n16680, n16681, n16682, n16683, n16684,
         n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692,
         n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700,
         n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
         n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716,
         n16717, n16718, n16719, n16720, n16721, n16722, n16723, n16724,
         n16725, n16726, n16727, n16728, n16729, n16730, n16731, n16732,
         n16733, n16734, n16735, n16736, n16737, n16738, n16739, n16740,
         n16741, n16742, n16743, n16744, n16745, n16746, n16747, n16748,
         n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756,
         n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
         n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772,
         n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780,
         n16781, n16782, n16783, n16784, n16785, n16786, n16787, n16788,
         n16789, n16790, n16791, n16792, n16793, n16794, n16795, n16796,
         n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804,
         n16805, n16806, n16807, n16808, n16809, n16810, n16811, n16812,
         n16813, n16814, n16815, n16816, n16817, n16818, n16819, n16820,
         n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
         n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836,
         n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844,
         n16845, n16846, n16847, n16848, n16849, n16850, n16851, n16852,
         n16853, n16854, n16855, n16856, n16857, n16858, n16859, n16860,
         n16861, n16862, n16863, n16864, n16865, n16866, n16867, n16868,
         n16869, n16870, n16871, n16872, n16873, n16874, n16875, n16876,
         n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
         n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892,
         n16893, n16894, n16895, n16896, n16897, n16898, n16899, n16900,
         n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908,
         n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916,
         n16917, n16918, n16919, n16920, n16921, n16922, n16923, n16924,
         n16925, n16926, n16927, n16928, n16929, n16930, n16931, n16932,
         n16933, n16934, n16935, n16936, n16937, n16938, n16939, n16940,
         n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948,
         n16949, n16950, n16951, n16952, n16953, n16954, n16955, n16956,
         n16957, n16958, n16959, n16960, n16961, n16962, n16963, n16964,
         n16965, n16966, n16967, n16968, n16969, n16970, n16971, n16972,
         n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980,
         n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988,
         n16989, n16990, n16991, n16992, n16993, n16994, n16995, n16996,
         n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004,
         n17005, n17006, n17007, n17008, n17009, n17010, n17011, n17012,
         n17013, n17014, n17015, n17016, n17017, n17018, n17019, n17020,
         n17021, n17022, n17023, n17024, n17025, n17026, n17027, n17028,
         n17029, n17030, n17031, n17032, n17033, n17034, n17035, n17036,
         n17037, n17038, n17039, n17040, n17041, n17042, n17043, n17044,
         n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052,
         n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060,
         n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
         n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076,
         n17077, n17078, n17079, n17080, n17081, n17082, n17083, n17084,
         n17085, n17086, n17087, n17088, n17089, n17090, n17091, n17092,
         n17093, n17094, n17095, n17096, n17097, n17098, n17099, n17100,
         n17101, n17102, n17103, n17104, n17105, n17106, n17107, n17108,
         n17109, n17110, n17111, n17112, n17113, n17114, n17115, n17116,
         n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124,
         n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132,
         n17133, n17134, n17135, n17136, n17137, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
         n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
         n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
         n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
         n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
         n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
         n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
         n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
         n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
         n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
         n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
         n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
         n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
         n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
         n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
         n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349,
         n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
         n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
         n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
         n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
         n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
         n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
         n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
         n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
         n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
         n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
         n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
         n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
         n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
         n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
         n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
         n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
         n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
         n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
         n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
         n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
         n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
         n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
         n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
         n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845,
         n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
         n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
         n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
         n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
         n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
         n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
         n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
         n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
         n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
         n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
         n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
         n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
         n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
         n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
         n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
         n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
         n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
         n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
         n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
         n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
         n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
         n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
         n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
         n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
         n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
         n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
         n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
         n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
         n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
         n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
         n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
         n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
         n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
         n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
         n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
         n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
         n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
         n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
         n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
         n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
         n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
         n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
         n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
         n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
         n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
         n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
         n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
         n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
         n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
         n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
         n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
         n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
         n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
         n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
         n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
         n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
         n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
         n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
         n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
         n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
         n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
         n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
         n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
         n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
         n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
         n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
         n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
         n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
         n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
         n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
         n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
         n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
         n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
         n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
         n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
         n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
         n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
         n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
         n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
         n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
         n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
         n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
         n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
         n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
         n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
         n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
         n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
         n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
         n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
         n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
         n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
         n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
         n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
         n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
         n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
         n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
         n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
         n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
         n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
         n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
         n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
         n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
         n18982, n18983, n18984, n18985, n18986, n18987, n18989, n18990,
         n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
         n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006,
         n19007, n19008, n19009, n19010, n19011, n19012, n19013, n19014,
         n19015, n19016, n19017, n19018, n19019, n19020, n19021, n19022,
         n19023, n19024, n19025, n19026, n19027, n19028, n19029, n19030,
         n19031, n19032, n19033, n19034, n19035, n19036, n19037, n19038,
         n19039, n19040, n19041, n19042, n19043, n19044, n19045, n19046,
         n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
         n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062,
         n19063, n19064, n19065, n19066, n19067, n19068, n19069, n19070,
         n19071, n19072, n19073, n19074, n19075, n19076, n19077, n19078,
         n19079, n19080, n19081, n19082, n19083, n19084, n19085, n19086,
         n19087, n19088, n19089, n19090, n19091, n19092, n19093, n19094,
         n19095, n19096, n19097, n19098, n19099, n19100, n19101, n19102,
         n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110,
         n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118,
         n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126,
         n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134,
         n19135, n19136, n19137, n19138, n19139, n19140, n19141, n19142,
         n19143, n19144, n19145, n19146, n19147, n19148, n19149, n19150,
         n19151, n19152, n19153, n19154, n19155, n19156, n19157, n19158,
         n19159, n19160, n19161, n19162, n19163, n19164, n19165, n19166,
         n19167, n19168, n19169, n19170, n19171, n19172, n19173, n19174,
         n19175, n19176, n19177, n19178, n19179, n19180, n19181, n19182,
         n19183, n19184, n19185, n19186, n19187, n19188, n19189, n19190,
         n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198,
         n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206,
         n19207, n19208, n19209, n19210, n19211, n19212, n19213, n19214,
         n19215, n19216, n19217, n19218, n19219, n19220, n19221, n19222,
         n19223, n19224, n19225, n19226, n19227, n19228, n19229, n19230,
         n19231, n19232, n19233, n19234, n19235, n19236, n19237, n19238,
         n19239, n19240, n19241, n19242, n19243, n19244, n19245, n19246,
         n19247, n19248, n19249, n19250, n19251, n19252, n19253, n19254,
         n19255, n19256, n19257, n19258, n19259, n19260, n19261, n19262,
         n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270,
         n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278,
         n19279, n19280, n19281, n19282, n19283, n19284, n19285, n19286,
         n19287, n19288, n19289, n19290, n19291, n19292, n19293, n19294,
         n19295, n19296, n19297, n19298, n19299, n19300, n19301, n19302,
         n19303, n19304, n19305, n19306, n19307, n19308, n19309, n19310,
         n19311, n19312, n19313, n19314, n19315, n19316, n19317, n19318,
         n19319, n19320, n19321, n19322, n19323, n19324, n19325, n19326,
         n19327, n19328, n19329, n19330, n19331, n19332, n19333, n19334,
         n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342,
         n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350,
         n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358,
         n19359, n19360, n19361, n19362, n19363, n19364, n19365, n19366,
         n19367, n19368, n19369, n19370, n19371, n19372, n19373, n19374,
         n19375, n19376, n19377, n19378, n19379, n19380, n19381, n19382,
         n19383, n19384, n19385, n19386, n19387, n19388, n19389, n19390,
         n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398,
         n19399, n19400, n19401, n19402, n19403, n19404, n19405, n19406,
         n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414,
         n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422,
         n19423, n19424, n19425, n19426, n19427, n19428, n19429, n19430,
         n19431, n19432, n19433, n19434, n19435, n19436, n19437, n19438,
         n19439, n19440, n19441, n19442, n19443, n19444, n19445, n19446,
         n19447, n19448, n19449, n19450, n19451, n19452, n19453, n19454,
         n19455, n19456, n19457, n19458, n19459, n19460, n19461, n19462,
         n19463, n19464, n19465, n19466, n19467, n19468, n19469, n19470,
         n19471, n19472, n19473, n19474, n19475, n19476, n19477, n19478,
         n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486,
         n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494,
         n19495, n19496, n19497, n19498, n19499, n19500, n19501, n19502,
         n19503, n19504, n19505, n19506, n19507, n19508, n19509, n19510,
         n19511, n19512, n19513, n19514, n19515, n19516, n19517, n19518,
         n19519, n19520, n19521, n19522, n19523, n19524, n19525, n19526,
         n19527, n19528, n19529, n19530, n19531, n19532, n19533, n19534,
         n19535, n19536, n19537, n19538, n19539, n19540, n19541, n19542,
         n19543, n19544, n19545, n19546, n19547, n19548, n19549, n19550,
         n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558,
         n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566,
         n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574,
         n19575, n19576, n19577, n19578, n19579, n19580, n19581, n19582,
         n19583, n19584, n19585, n19586, n19587, n19588, n19589, n19590,
         n19591, n19592, n19593, n19594, n19595, n19596, n19597, n19598,
         n19599, n19600, n19601, n19602, n19603, n19604, n19605, n19606,
         n19607, n19608, n19609, n19610, n19611, n19612, n19613, n19614,
         n19615, n19616, n19617, n19618, n19619, n19620, n19621, n19622,
         n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630,
         n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638,
         n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
         n19647, n19648, n19649, n19650, n19651, n19652, n19653, n19654,
         n19655, n19656, n19657, n19658, n19659, n19660, n19661, n19662,
         n19663, n19664, n19665, n19666, n19667, n19668, n19669, n19670,
         n19671, n19672, n19673, n19674, n19675, n19676, n19677, n19678,
         n19679, n19680, n19681, n19682, n19683, n19684, n19685, n19686,
         n19687, n19688, n19689, n19690, n19691, n19692, n19693, n19694,
         n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702,
         n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710,
         n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718,
         n19719, n19720, n19721, n19722, n19723, n19724, n19725, n19726,
         n19727, n19728, n19729, n19730, n19731, n19732, n19733, n19734,
         n19735, n19736, n19737, n19738, n19739, n19740, n19741, n19742,
         n19743, n19744, n19745, n19746, n19747, n19748, n19749, n19750,
         n19751, n19752, n19753, n19754, n19755, n19756, n19757, n19758,
         n19759, n19760, n19761, n19762, n19763, n19764, n19765, n19766,
         n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774,
         n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
         n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790,
         n19791, n19792, n19793, n19794, n19795, n19796, n19797, n19798,
         n19799, n19800, n19801, n19802, n19803, n19804, n19805, n19806,
         n19807, n19808, n19809, n19810, n19811, n19812, n19813, n19814,
         n19815, n19816, n19817, n19818, n19819, n19820, n19821, n19822,
         n19823, n19824, n19825, n19826, n19827, n19828, n19829, n19830,
         n19831, n19832, n19833, n19834, n19835, n19836, n19837, n19838,
         n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846,
         n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
         n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862,
         n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870,
         n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878,
         n19879, n19880, n19881, n19882, n19883, n19884, n19885, n19886,
         n19887, n19888, n19889, n19890, n19891, n19892, n19893, n19894,
         n19895, n19896, n19897, n19898, n19899, n19900, n19901, n19902,
         n19903, n19904, n19905, n19906, n19907, n19908, n19909, n19910,
         n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918,
         n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926,
         n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934,
         n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942,
         n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950,
         n19951, n19952, n19953, n19954, n19955, n19956, n19957, n19958,
         n19959, n19960, n19961, n19962, n19963, n19964, n19965, n19966,
         n19967, n19968, n19969, n19970, n19971, n19972, n19973, n19974,
         n19975, n19976, n19977, n19978, n19979, n19980, n19981, n19982,
         n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990,
         n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
         n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006,
         n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014,
         n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022,
         n20023, n20024, n20025, n20026, n20027, n20028, n20029, n20030,
         n20031, n20032, n20033, n20034, n20035, n20036, n20037, n20038,
         n20039, n20040, n20041, n20042, n20043, n20044, n20045, n20046,
         n20047, n20048, n20049, n20050, n20051, n20052, n20053, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086,
         n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094,
         n20095, n20096, n20097, n20098, n20099, n20100, n20101, n20102,
         n20103, n20104, n20105, n20106, n20107, n20108, n20109, n20110,
         n20111, n20112, n20113, n20114, n20115, n20116, n20117, n20118,
         n20119, n20120, n20121, n20122, n20123, n20124, n20125, n20126,
         n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134,
         n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142,
         n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150,
         n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158,
         n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166,
         n20167, n20168, n20169, n20170, n20171, n20172, n20173, n20174,
         n20175, n20176, n20177, n20178, n20179, n20180, n20181, n20182,
         n20183, n20184, n20185, n20186, n20187, n20188, n20189, n20190,
         n20191, n20192, n20193, n20194, n20195, n20196, n20197, n20198,
         n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206,
         n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
         n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222,
         n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230,
         n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238,
         n20239, n20240, n20241, n20242, n20243, n20244, n20245, n20246,
         n20247, n20248, n20249, n20250, n20251, n20252, n20253, n20254,
         n20255, n20256, n20257, n20258, n20259, n20260, n20261, n20262,
         n20263, n20264, n20265, n20266, n20267, n20268, n20269, n20270,
         n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278,
         n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
         n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294,
         n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302,
         n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310,
         n20311, n20312, n20313, n20314, n20315, n20316, n20317, n20318,
         n20319, n20320, n20321, n20322, n20323, n20324, n20325, n20326,
         n20327, n20328, n20329, n20330, n20331, n20332, n20333, n20334,
         n20335, n20336, n20337, n20338, n20339, n20340, n20341, n20342,
         n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350,
         n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
         n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366,
         n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374,
         n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382,
         n20383, n20384, n20385, n20386, n20387, n20388, n20389, n20390,
         n20391, n20392, n20393, n20394, n20395, n20396, n20397, n20398,
         n20399, n20400, n20401, n20402, n20403, n20404, n20405, n20406,
         n20407, n20408, n20409, n20410, n20411, n20412, n20413, n20414,
         n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422,
         n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
         n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438,
         n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446,
         n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454,
         n20455, n20456, n20457, n20458, n20459, n20460, n20461, n20462,
         n20463, n20464, n20465, n20466, n20467, n20468, n20469, n20470,
         n20471, n20472, n20473, n20474, n20475, n20476, n20477, n20478,
         n20479, n20480, n20481, n20482, n20483, n20484, n20485, n20486,
         n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494,
         n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
         n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20510,
         n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518,
         n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526,
         n20527, n20528, n20529, n20530, n20531, n20532, n20533, n20534,
         n20535, n20536, n20537, n20538, n20539, n20540, n20541, n20542,
         n20543, n20544, n20545, n20546, n20547, n20548, n20549, n20550,
         n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
         n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566,
         n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574,
         n20575, n20576, n20577, n20578, n20579, n20580, n20581, n20582,
         n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590,
         n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598,
         n20599, n20600, n20601, n20602, n20603, n20604, n20605, n20606,
         n20607, n20608, n20609, n20610, n20611, n20612, n20613, n20614,
         n20615, n20616, n20617, n20618, n20619, n20620, n20621, n20622,
         n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
         n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638,
         n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646,
         n20647, n20648, n20649, n20650, n20651, n20652, n20653, n20654,
         n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662,
         n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670,
         n20671, n20672, n20673, n20674, n20675, n20676, n20677, n20678,
         n20679, n20680, n20681, n20682, n20683, n20684, n20685, n20686,
         n20687, n20688, n20689, n20690, n20691, n20692, n20693, n20694,
         n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
         n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710,
         n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718,
         n20719, n20720, n20721, n20722, n20723, n20724, n20725, n20726,
         n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734,
         n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742,
         n20743, n20744, n20745, n20746, n20747, n20748, n20749, n20750,
         n20751, n20752, n20753, n20754, n20755, n20756, n20757, n20758,
         n20759, n20760, n20761, n20762, n20763, n20764, n20765, n20766,
         n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774,
         n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782,
         n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790,
         n20791, n20792, n20793, n20794, n20795, n20796, n20797, n20798,
         n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806,
         n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814,
         n20815, n20816, n20817, n20818, n20819, n20820, n20821, n20822,
         n20823, n20824, n20825, n20826, n20827, n20828, n20829, n20830,
         n20831, n20832, n20833, n20834, n20835, n20836, n20837, n20838,
         n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846,
         n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854,
         n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862,
         n20863, n20864, n20865, n20866, n20867, n20868, n20869, n20870,
         n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878,
         n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886,
         n20887, n20888, n20889, n20890, n20891, n20892, n20893, n20894,
         n20895, n20896, n20897, n20898, n20899, n20900, n20901, n20902,
         n20903, n20904, n20905, n20906, n20907, n20908, n20909, n20910,
         n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918,
         n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926,
         n20927, n20928, n20929;

  NOR2_X1 U11037 ( .A1(n9773), .A2(n9772), .ZN(n9771) );
  INV_X1 U11038 ( .A(n17822), .ZN(n17794) );
  CLKBUF_X1 U11039 ( .A(n15068), .Z(n9593) );
  CLKBUF_X1 U11040 ( .A(n14291), .Z(n13781) );
  AND2_X1 U11041 ( .A1(n10011), .A2(n10286), .ZN(n19309) );
  NAND3_X1 U11042 ( .A1(n11305), .A2(n11304), .A3(n11303), .ZN(n17292) );
  AND2_X1 U11043 ( .A1(n12498), .A2(n10286), .ZN(n10284) );
  BUF_X1 U11044 ( .A(n12519), .Z(n19178) );
  INV_X2 U11045 ( .A(n12437), .ZN(n18182) );
  NAND2_X1 U11046 ( .A1(n10251), .A2(n10255), .ZN(n13963) );
  INV_X4 U11047 ( .A(n17159), .ZN(n12941) );
  OR2_X1 U11048 ( .A1(n10246), .A2(n10245), .ZN(n10258) );
  INV_X1 U11049 ( .A(n11441), .ZN(n17161) );
  BUF_X1 U11050 ( .A(n10340), .Z(n12666) );
  AND2_X1 U11051 ( .A1(n10300), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12631) );
  AND2_X1 U11052 ( .A1(n12678), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12545) );
  CLKBUF_X1 U11053 ( .A(n10339), .Z(n12650) );
  CLKBUF_X2 U11054 ( .A(n11462), .Z(n17144) );
  CLKBUF_X2 U11055 ( .A(n11410), .Z(n9597) );
  CLKBUF_X1 U11056 ( .A(n11306), .Z(n9623) );
  CLKBUF_X2 U11057 ( .A(n11398), .Z(n17156) );
  CLKBUF_X2 U11058 ( .A(n11410), .Z(n9596) );
  BUF_X1 U11059 ( .A(n16916), .Z(n17154) );
  CLKBUF_X3 U11060 ( .A(n17107), .Z(n9603) );
  INV_X4 U11061 ( .A(n9591), .ZN(n9602) );
  CLKBUF_X2 U11062 ( .A(n12293), .Z(n9631) );
  CLKBUF_X1 U11064 ( .A(n10293), .Z(n12817) );
  INV_X2 U11065 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16304) );
  INV_X2 U11066 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n16301) );
  AND2_X1 U11067 ( .A1(n11487), .A2(n13347), .ZN(n11808) );
  AND2_X1 U11068 ( .A1(n9793), .A2(n11484), .ZN(n12293) );
  AND2_X1 U11069 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13377) );
  OAI211_X1 U11070 ( .C1(n10165), .C2(n10164), .A(n10163), .B(n10664), .ZN(
        n10856) );
  NAND2_X1 U11071 ( .A1(n11626), .A2(n11620), .ZN(n13400) );
  AND3_X1 U11072 ( .A1(n11569), .A2(n14596), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12385) );
  AND2_X1 U11073 ( .A1(n12678), .A2(n16304), .ZN(n12660) );
  AND4_X1 U11074 ( .A1(n10290), .A2(n10289), .A3(n10288), .A4(n10287), .ZN(
        n10291) );
  AND2_X1 U11075 ( .A1(n11486), .A2(n13377), .ZN(n11691) );
  OR2_X1 U11076 ( .A1(n10521), .A2(n12848), .ZN(n10609) );
  NAND2_X1 U11077 ( .A1(n10471), .A2(n10465), .ZN(n10505) );
  INV_X1 U11078 ( .A(n10733), .ZN(n11182) );
  INV_X2 U11079 ( .A(n10891), .ZN(n11160) );
  INV_X2 U11080 ( .A(n19823), .ZN(n10664) );
  AND3_X1 U11081 ( .A1(n13670), .A2(n10282), .A3(n19178), .ZN(n10371) );
  AND2_X1 U11082 ( .A1(n10284), .A2(n10283), .ZN(n14102) );
  CLKBUF_X3 U11084 ( .A(n11349), .Z(n9607) );
  NOR2_X1 U11085 ( .A1(n15855), .A2(n14732), .ZN(n9613) );
  INV_X2 U11086 ( .A(n14596), .ZN(n20105) );
  NOR2_X1 U11087 ( .A1(n10505), .A2(n9876), .ZN(n10529) );
  NOR2_X1 U11088 ( .A1(n15454), .A2(n9970), .ZN(n15228) );
  INV_X1 U11089 ( .A(n10371), .ZN(n19277) );
  AND2_X1 U11090 ( .A1(n10284), .A2(n10282), .ZN(n14040) );
  AOI21_X1 U11091 ( .B1(n15728), .B2(n15727), .A(n16406), .ZN(n15729) );
  NOR2_X2 U11092 ( .A1(n17322), .A2(n12960), .ZN(n17730) );
  CLKBUF_X2 U11093 ( .A(n13574), .Z(n14522) );
  NOR2_X1 U11094 ( .A1(n15855), .A2(n14717), .ZN(n14726) );
  INV_X1 U11095 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11478) );
  NOR2_X1 U11096 ( .A1(n15454), .A2(n15443), .ZN(n15250) );
  NAND2_X1 U11097 ( .A1(n10602), .A2(n9771), .ZN(n15241) );
  NOR2_X1 U11098 ( .A1(n14047), .A2(n19312), .ZN(n19421) );
  XNOR2_X1 U11099 ( .A(n12422), .B(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n16805) );
  INV_X1 U11100 ( .A(n17292), .ZN(n18193) );
  INV_X1 U11101 ( .A(n17666), .ZN(n17675) );
  INV_X1 U11102 ( .A(n19927), .ZN(n19940) );
  INV_X2 U11103 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18793) );
  OR2_X1 U11104 ( .A1(n11291), .A2(n11289), .ZN(n9591) );
  NOR3_X2 U11105 ( .A1(n17284), .A2(n17250), .A3(n17210), .ZN(n17246) );
  INV_X1 U11106 ( .A(n19829), .ZN(n11085) );
  XNOR2_X2 U11107 ( .A(n13627), .B(n13634), .ZN(n13626) );
  XNOR2_X1 U11109 ( .A(n11764), .B(n11763), .ZN(n15068) );
  NAND2_X1 U11110 ( .A1(n10208), .A2(n10196), .ZN(n9594) );
  INV_X2 U11111 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13968) );
  OAI22_X2 U11113 ( .A1(n10748), .A2(n13604), .B1(n13937), .B2(n13826), .ZN(
        n10200) );
  NOR2_X1 U11115 ( .A1(n11294), .A2(n11293), .ZN(n11410) );
  AND2_X1 U11116 ( .A1(n9972), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9598) );
  INV_X1 U11117 ( .A(n9598), .ZN(n9599) );
  AND2_X2 U11118 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13676) );
  NOR2_X1 U11119 ( .A1(n11293), .A2(n11289), .ZN(n11398) );
  INV_X4 U11120 ( .A(n10128), .ZN(n12699) );
  INV_X2 U11121 ( .A(n10127), .ZN(n9601) );
  INV_X2 U11122 ( .A(n18629), .ZN(n18616) );
  OAI21_X4 U11123 ( .B1(n18609), .B2(n18619), .A(n18608), .ZN(n18629) );
  NAND2_X1 U11124 ( .A1(n9748), .A2(n10591), .ZN(n15267) );
  AND2_X1 U11125 ( .A1(n9921), .A2(n17829), .ZN(n16407) );
  NAND2_X1 U11126 ( .A1(n9956), .A2(n14499), .ZN(n14503) );
  AND2_X1 U11127 ( .A1(n11834), .A2(n11833), .ZN(n13638) );
  NAND2_X1 U11128 ( .A1(n10077), .A2(n12530), .ZN(n13652) );
  AND2_X1 U11129 ( .A1(n9841), .A2(n9691), .ZN(n10077) );
  INV_X1 U11130 ( .A(n11807), .ZN(n11821) );
  AND2_X1 U11131 ( .A1(n9614), .A2(n9615), .ZN(n13564) );
  INV_X4 U11132 ( .A(n17721), .ZN(n17731) );
  AOI21_X1 U11133 ( .B1(n10271), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A(
        n10270), .ZN(n10272) );
  NAND2_X2 U11134 ( .A1(n19175), .A2(n15537), .ZN(n15671) );
  NOR2_X1 U11135 ( .A1(n17321), .A2(n17396), .ZN(n17316) );
  OR3_X1 U11136 ( .A1(n10285), .A2(n10286), .A3(n15666), .ZN(n14185) );
  NOR2_X2 U11137 ( .A1(n9732), .A2(n18052), .ZN(n18594) );
  NOR2_X2 U11138 ( .A1(n13110), .A2(n19829), .ZN(n11114) );
  INV_X2 U11139 ( .A(n18089), .ZN(n18110) );
  NAND2_X1 U11141 ( .A1(n18631), .A2(n18616), .ZN(n18089) );
  AOI21_X1 U11142 ( .B1(n15810), .B2(n15809), .A(n18811), .ZN(n17207) );
  OAI211_X1 U11143 ( .C1(n18622), .C2(n15698), .A(n18596), .B(n18815), .ZN(
        n15810) );
  NOR2_X1 U11144 ( .A1(n17758), .A2(n9924), .ZN(n17752) );
  NOR2_X2 U11145 ( .A1(n12982), .A2(n18619), .ZN(n18622) );
  NAND2_X1 U11147 ( .A1(n12983), .A2(n12982), .ZN(n18605) );
  AND2_X1 U11148 ( .A1(n10469), .A2(n10468), .ZN(n10471) );
  NOR4_X2 U11149 ( .A1(n12437), .A2(n12991), .A3(n18160), .A4(n12436), .ZN(
        n17415) );
  NAND2_X2 U11151 ( .A1(n11558), .A2(n10079), .ZN(n11634) );
  AND3_X1 U11152 ( .A1(n11616), .A2(n13417), .A3(n13395), .ZN(n11617) );
  INV_X2 U11154 ( .A(n11569), .ZN(n11626) );
  NOR2_X1 U11155 ( .A1(n9809), .A2(n9808), .ZN(n9807) );
  AND4_X1 U11156 ( .A1(n11597), .A2(n11596), .A3(n11595), .A4(n11594), .ZN(
        n11614) );
  AND4_X1 U11157 ( .A1(n11580), .A2(n11579), .A3(n11578), .A4(n11577), .ZN(
        n11591) );
  AND4_X1 U11158 ( .A1(n10152), .A2(n10151), .A3(n10150), .A4(n10149), .ZN(
        n10153) );
  BUF_X2 U11159 ( .A(n11744), .Z(n12254) );
  CLKBUF_X3 U11160 ( .A(n11327), .Z(n9606) );
  CLKBUF_X2 U11161 ( .A(n11513), .Z(n12233) );
  CLKBUF_X3 U11162 ( .A(n11403), .Z(n9605) );
  CLKBUF_X2 U11163 ( .A(n11602), .Z(n12161) );
  BUF_X1 U11164 ( .A(n11295), .Z(n9622) );
  CLKBUF_X2 U11165 ( .A(n11462), .Z(n17052) );
  NAND2_X1 U11166 ( .A1(n9730), .A2(n9729), .ZN(n16958) );
  INV_X4 U11167 ( .A(n9652), .ZN(n17160) );
  BUF_X2 U11168 ( .A(n11658), .Z(n12300) );
  CLKBUF_X2 U11169 ( .A(n11593), .Z(n12228) );
  NOR2_X1 U11170 ( .A1(n11294), .A2(n11296), .ZN(n11295) );
  CLKBUF_X2 U11171 ( .A(n11808), .Z(n12207) );
  AND2_X2 U11172 ( .A1(n9793), .A2(n11485), .ZN(n12278) );
  AND2_X2 U11173 ( .A1(n11484), .A2(n13377), .ZN(n11737) );
  CLKBUF_X2 U11175 ( .A(n12249), .Z(n12295) );
  INV_X2 U11176 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10080) );
  NOR2_X4 U11177 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13964) );
  NAND2_X1 U11178 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18618) );
  AOI21_X1 U11179 ( .B1(n14830), .B2(n10059), .A(n14419), .ZN(n14420) );
  AOI21_X1 U11180 ( .B1(n15004), .B2(n20093), .A(n9819), .ZN(n14883) );
  XNOR2_X1 U11181 ( .A(n14880), .B(n15009), .ZN(n15004) );
  NAND2_X1 U11182 ( .A1(n15242), .A2(n15241), .ZN(n15435) );
  OR2_X1 U11183 ( .A1(n12485), .A2(n19174), .ZN(n12486) );
  AND2_X1 U11184 ( .A1(n15587), .A2(n15366), .ZN(n15594) );
  OAI21_X1 U11185 ( .B1(n15347), .B2(n11107), .A(n15332), .ZN(n15320) );
  AND2_X1 U11186 ( .A1(n14920), .A2(n14919), .ZN(n14933) );
  NAND2_X1 U11187 ( .A1(n9720), .A2(n9719), .ZN(n15235) );
  INV_X1 U11188 ( .A(n15454), .ZN(n9720) );
  INV_X1 U11189 ( .A(n9613), .ZN(n14731) );
  INV_X1 U11190 ( .A(n15331), .ZN(n15347) );
  NAND2_X1 U11191 ( .A1(n15961), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14412) );
  NAND2_X1 U11192 ( .A1(n9739), .A2(n10059), .ZN(n15962) );
  AND2_X1 U11193 ( .A1(n9920), .A2(n9918), .ZN(n16399) );
  NAND2_X1 U11194 ( .A1(n14889), .A2(n9740), .ZN(n9739) );
  NAND2_X1 U11195 ( .A1(n9747), .A2(n10597), .ZN(n15258) );
  OR2_X1 U11196 ( .A1(n15134), .A2(n15133), .ZN(n15131) );
  INV_X1 U11197 ( .A(n9815), .ZN(n14906) );
  OAI21_X1 U11198 ( .B1(n15267), .B2(n10017), .A(n10015), .ZN(n10601) );
  AND3_X2 U11199 ( .A1(n9968), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n9641), .ZN(n11131) );
  OR2_X1 U11200 ( .A1(n12738), .A2(n12737), .ZN(n10058) );
  AND2_X1 U11201 ( .A1(n15391), .A2(n10736), .ZN(n10737) );
  NAND2_X1 U11202 ( .A1(n16407), .A2(n17466), .ZN(n15728) );
  NAND2_X1 U11203 ( .A1(n15145), .A2(n9699), .ZN(n12736) );
  NOR2_X1 U11204 ( .A1(n9969), .A2(n9713), .ZN(n9967) );
  OR2_X1 U11205 ( .A1(n17492), .A2(n9922), .ZN(n9921) );
  NAND2_X1 U11206 ( .A1(n14503), .A2(n10722), .ZN(n10723) );
  NAND2_X1 U11207 ( .A1(n9657), .A2(n9636), .ZN(n9813) );
  OAI211_X1 U11208 ( .C1(n10467), .C2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n9757), .B(n9756), .ZN(n14171) );
  AOI21_X1 U11210 ( .B1(n16014), .B2(n10032), .A(n10031), .ZN(n10033) );
  XNOR2_X1 U11211 ( .A(n10735), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16253) );
  AND2_X1 U11212 ( .A1(n10623), .A2(n10615), .ZN(n15239) );
  OR2_X1 U11213 ( .A1(n9638), .A2(n12718), .ZN(n10057) );
  AND2_X1 U11214 ( .A1(n10071), .A2(n14144), .ZN(n10047) );
  NAND2_X1 U11215 ( .A1(n9760), .A2(n10504), .ZN(n14170) );
  AND3_X2 U11216 ( .A1(n13639), .A2(n13725), .A3(n13791), .ZN(n9618) );
  AND2_X1 U11217 ( .A1(n15975), .A2(n15973), .ZN(n14922) );
  NOR2_X1 U11218 ( .A1(n9746), .A2(n14918), .ZN(n10048) );
  INV_X2 U11220 ( .A(n13814), .ZN(n12536) );
  INV_X1 U11221 ( .A(n13876), .ZN(n11880) );
  NAND2_X1 U11222 ( .A1(n14407), .A2(n15985), .ZN(n14918) );
  OR2_X1 U11223 ( .A1(n14912), .A2(n10049), .ZN(n9746) );
  NAND2_X1 U11224 ( .A1(n13698), .A2(n10710), .ZN(n19144) );
  OAI21_X1 U11225 ( .B1(n13717), .B2(n13716), .A(n13715), .ZN(n13838) );
  NAND2_X1 U11226 ( .A1(n13700), .A2(n13699), .ZN(n13698) );
  XNOR2_X1 U11227 ( .A(n11875), .B(n10053), .ZN(n14135) );
  NAND2_X1 U11228 ( .A1(n13562), .A2(n11779), .ZN(n13572) );
  NAND2_X1 U11229 ( .A1(n11821), .A2(n11822), .ZN(n11846) );
  NAND2_X1 U11230 ( .A1(n11821), .A2(n9647), .ZN(n14149) );
  OR2_X1 U11231 ( .A1(n10405), .A2(n10404), .ZN(n10422) );
  NOR2_X1 U11232 ( .A1(n13932), .A2(n13933), .ZN(n14031) );
  NAND2_X1 U11233 ( .A1(n9937), .A2(n11797), .ZN(n11807) );
  INV_X1 U11234 ( .A(n17815), .ZN(n17827) );
  NAND2_X1 U11235 ( .A1(n17688), .A2(n17693), .ZN(n17676) );
  NAND2_X1 U11236 ( .A1(n17322), .A2(n17797), .ZN(n17734) );
  OR2_X1 U11237 ( .A1(n10573), .A2(n10553), .ZN(n18863) );
  AND3_X1 U11238 ( .A1(n10281), .A2(n10280), .A3(n9662), .ZN(n10290) );
  NAND2_X1 U11239 ( .A1(n10574), .A2(n10609), .ZN(n10573) );
  INV_X1 U11240 ( .A(n10363), .ZN(n19491) );
  NAND2_X1 U11241 ( .A1(n13521), .A2(n12524), .ZN(n13511) );
  AND2_X1 U11242 ( .A1(n10267), .A2(n10278), .ZN(n19433) );
  AND2_X1 U11243 ( .A1(n15794), .A2(n15019), .ZN(n15057) );
  AND2_X1 U11244 ( .A1(n10011), .A2(n19178), .ZN(n19197) );
  AND2_X1 U11245 ( .A1(n10267), .A2(n10283), .ZN(n19460) );
  NAND2_X1 U11246 ( .A1(n14578), .A2(n13289), .ZN(n15055) );
  OAI21_X1 U11247 ( .B1(n9738), .B2(n9860), .A(n9859), .ZN(n13080) );
  CLKBUF_X1 U11248 ( .A(n13421), .Z(n20491) );
  AND2_X1 U11249 ( .A1(n13529), .A2(n12512), .ZN(n13517) );
  OR3_X1 U11250 ( .A1(n10285), .A2(n15666), .A3(n19178), .ZN(n19380) );
  NOR2_X2 U11251 ( .A1(n19829), .A2(n14068), .ZN(n14064) );
  NAND2_X1 U11252 ( .A1(n13264), .A2(n13263), .ZN(n13289) );
  NAND2_X1 U11253 ( .A1(n11685), .A2(n11684), .ZN(n11713) );
  XOR2_X1 U11254 ( .A(n12961), .B(n12962), .Z(n17740) );
  OR2_X1 U11255 ( .A1(n11730), .A2(n11731), .ZN(n11728) );
  NAND2_X1 U11256 ( .A1(n11703), .A2(n11702), .ZN(n11704) );
  XNOR2_X1 U11257 ( .A(n10235), .B(n10234), .ZN(n10248) );
  NAND2_X1 U11258 ( .A1(n17772), .A2(n12955), .ZN(n17759) );
  NOR2_X1 U11259 ( .A1(n10230), .A2(n10229), .ZN(n10235) );
  NAND3_X1 U11260 ( .A1(n10189), .A2(n9754), .A3(n10202), .ZN(n10225) );
  AOI21_X1 U11261 ( .B1(n11153), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10242), .ZN(n10743) );
  AND2_X1 U11262 ( .A1(n10201), .A2(n10188), .ZN(n9754) );
  INV_X1 U11263 ( .A(n17415), .ZN(n15697) );
  NAND2_X1 U11264 ( .A1(n9656), .A2(n9849), .ZN(n12488) );
  OAI21_X1 U11265 ( .B1(n10213), .B2(n10178), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n10182) );
  NAND2_X1 U11266 ( .A1(n10843), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10208) );
  OAI21_X1 U11267 ( .B1(n10748), .B2(n10217), .A(n10076), .ZN(n10218) );
  CLKBUF_X1 U11268 ( .A(n10748), .Z(n10826) );
  AND2_X1 U11269 ( .A1(n15707), .A2(n12431), .ZN(n12436) );
  AND3_X1 U11270 ( .A1(n10177), .A2(n11252), .A3(n10176), .ZN(n10178) );
  INV_X1 U11271 ( .A(n12990), .ZN(n18169) );
  NOR2_X1 U11272 ( .A1(n17336), .A2(n12939), .ZN(n12937) );
  NAND2_X1 U11273 ( .A1(n11622), .A2(n11621), .ZN(n13349) );
  AND2_X1 U11274 ( .A1(n11628), .A2(n11627), .ZN(n11644) );
  INV_X1 U11275 ( .A(n18187), .ZN(n17211) );
  AND2_X1 U11276 ( .A1(n9723), .A2(n9774), .ZN(n10662) );
  AND2_X1 U11277 ( .A1(n14588), .A2(n14522), .ZN(n13175) );
  NAND2_X1 U11278 ( .A1(n11626), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n14146) );
  NAND3_X1 U11279 ( .A1(n12950), .A2(n12949), .A3(n12948), .ZN(n15811) );
  INV_X2 U11280 ( .A(n11633), .ZN(n11558) );
  AND2_X1 U11281 ( .A1(n11632), .A2(n11631), .ZN(n12345) );
  INV_X1 U11282 ( .A(n17341), .ZN(n13015) );
  AOI21_X1 U11283 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19775), .A(
        n10461), .ZN(n10640) );
  NAND2_X1 U11284 ( .A1(n13907), .A2(n13246), .ZN(n13574) );
  AND2_X1 U11285 ( .A1(n13295), .A2(n10161), .ZN(n12847) );
  NAND2_X1 U11286 ( .A1(n10060), .A2(n9925), .ZN(n17346) );
  AND2_X2 U11287 ( .A1(n14596), .A2(n13907), .ZN(n14467) );
  INV_X1 U11288 ( .A(n14046), .ZN(n12860) );
  NAND2_X1 U11289 ( .A1(n9810), .A2(n9807), .ZN(n13359) );
  NAND2_X2 U11290 ( .A1(n10107), .A2(n10106), .ZN(n14046) );
  INV_X1 U11291 ( .A(n11620), .ZN(n11630) );
  INV_X1 U11292 ( .A(n10448), .ZN(n10161) );
  AND2_X1 U11293 ( .A1(n19823), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19830) );
  AND4_X1 U11294 ( .A1(n12905), .A2(n12904), .A3(n12902), .A4(n9670), .ZN(
        n9925) );
  NAND4_X2 U11295 ( .A1(n11544), .A2(n11543), .A3(n11542), .A4(n11541), .ZN(
        n11569) );
  NAND2_X1 U11296 ( .A1(n9869), .A2(n9867), .ZN(n10448) );
  NAND2_X1 U11297 ( .A1(n10112), .A2(n16304), .ZN(n10118) );
  AND4_X1 U11298 ( .A1(n11584), .A2(n11583), .A3(n11582), .A4(n11581), .ZN(
        n11590) );
  AND4_X1 U11299 ( .A1(n11536), .A2(n11535), .A3(n11534), .A4(n11533), .ZN(
        n11542) );
  NOR2_X2 U11300 ( .A1(n20099), .A2(n20102), .ZN(n20100) );
  AND4_X1 U11301 ( .A1(n11532), .A2(n11531), .A3(n11530), .A4(n11529), .ZN(
        n11543) );
  NAND2_X1 U11302 ( .A1(n10153), .A2(n16304), .ZN(n10160) );
  NOR2_X1 U11303 ( .A1(n9812), .A2(n9811), .ZN(n9810) );
  AND4_X1 U11304 ( .A1(n11500), .A2(n11499), .A3(n11498), .A4(n11497), .ZN(
        n11511) );
  AND4_X1 U11305 ( .A1(n11540), .A2(n11539), .A3(n11538), .A4(n11537), .ZN(
        n11541) );
  AND4_X1 U11306 ( .A1(n11496), .A2(n11495), .A3(n11494), .A4(n11493), .ZN(
        n11512) );
  INV_X1 U11307 ( .A(n11295), .ZN(n16985) );
  AND4_X1 U11308 ( .A1(n11528), .A2(n11527), .A3(n11526), .A4(n11525), .ZN(
        n11544) );
  AND4_X1 U11309 ( .A1(n11606), .A2(n11605), .A3(n11604), .A4(n11603), .ZN(
        n11612) );
  AND4_X1 U11310 ( .A1(n11601), .A2(n11600), .A3(n11599), .A4(n11598), .ZN(
        n11613) );
  AND4_X1 U11311 ( .A1(n11588), .A2(n11587), .A3(n11586), .A4(n11585), .ZN(
        n11589) );
  AND4_X1 U11312 ( .A1(n11576), .A2(n11575), .A3(n11574), .A4(n11573), .ZN(
        n11592) );
  AND4_X1 U11313 ( .A1(n11610), .A2(n11609), .A3(n11608), .A4(n11607), .ZN(
        n11611) );
  AND4_X1 U11314 ( .A1(n10111), .A2(n10110), .A3(n10109), .A4(n10108), .ZN(
        n10112) );
  INV_X1 U11315 ( .A(n11480), .ZN(n9811) );
  NAND4_X1 U11316 ( .A1(n10116), .A2(n10115), .A3(n10114), .A4(n10113), .ZN(
        n10117) );
  AND4_X1 U11317 ( .A1(n11508), .A2(n11507), .A3(n11506), .A4(n11505), .ZN(
        n11509) );
  AND4_X1 U11318 ( .A1(n11504), .A2(n11503), .A3(n11502), .A4(n11501), .ZN(
        n11510) );
  NAND2_X2 U11319 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19837), .ZN(n19751) );
  NAND2_X2 U11320 ( .A1(n19837), .A2(n19700), .ZN(n19750) );
  AND2_X1 U11321 ( .A1(n10083), .A2(n16304), .ZN(n9870) );
  AND2_X1 U11322 ( .A1(n10088), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9868) );
  INV_X2 U11323 ( .A(n16507), .ZN(U215) );
  INV_X2 U11324 ( .A(n9612), .ZN(n12551) );
  NAND2_X2 U11325 ( .A1(n18822), .A2(n18690), .ZN(n18738) );
  AND2_X1 U11326 ( .A1(n9961), .A2(n9960), .ZN(n10115) );
  AND3_X1 U11327 ( .A1(n9779), .A2(n9778), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n9974) );
  AND2_X1 U11328 ( .A1(n10121), .A2(n16304), .ZN(n9976) );
  AND2_X1 U11329 ( .A1(n10154), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10158) );
  AOI22_X1 U11330 ( .A1(n12293), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9627), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11520) );
  AND2_X2 U11331 ( .A1(n12831), .A2(n16304), .ZN(n12665) );
  CLKBUF_X3 U11332 ( .A(n11492), .Z(n12202) );
  AND2_X2 U11333 ( .A1(n12832), .A2(n16304), .ZN(n10320) );
  BUF_X2 U11334 ( .A(n10293), .Z(n12686) );
  INV_X2 U11335 ( .A(n16511), .ZN(n16513) );
  BUF_X4 U11336 ( .A(n10300), .Z(n12831) );
  AND2_X2 U11337 ( .A1(n12832), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12552) );
  OR2_X1 U11338 ( .A1(n11292), .A2(n18618), .ZN(n12876) );
  NAND3_X1 U11339 ( .A1(n18793), .A2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n18612), .ZN(n17159) );
  OR2_X1 U11340 ( .A1(n11289), .A2(n11292), .ZN(n9652) );
  NAND2_X1 U11341 ( .A1(n18793), .A2(n18786), .ZN(n16880) );
  AND2_X1 U11342 ( .A1(n11235), .A2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11234) );
  INV_X2 U11343 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11718) );
  AND2_X1 U11344 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11485) );
  INV_X1 U11346 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19802) );
  AND2_X2 U11347 ( .A1(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n9972) );
  NAND2_X1 U11348 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11291) );
  XNOR2_X1 U11349 ( .A(n11780), .B(n20259), .ZN(n20735) );
  INV_X1 U11350 ( .A(n17513), .ZN(n9609) );
  AOI211_X2 U11351 ( .C1(n15832), .C2(n19927), .A(n15831), .B(n15830), .ZN(
        n15833) );
  INV_X1 U11352 ( .A(n13733), .ZN(n9610) );
  NOR2_X1 U11353 ( .A1(n13652), .A2(n12532), .ZN(n13729) );
  AND2_X1 U11354 ( .A1(n12225), .A2(n9611), .ZN(n14623) );
  INV_X1 U11355 ( .A(n14637), .ZN(n9611) );
  NAND2_X1 U11356 ( .A1(n12829), .A2(n16304), .ZN(n9612) );
  NAND2_X1 U11357 ( .A1(n15068), .A2(n9617), .ZN(n9614) );
  OR2_X2 U11358 ( .A1(n9616), .A2(n11768), .ZN(n9615) );
  INV_X1 U11359 ( .A(n13392), .ZN(n9616) );
  AND2_X1 U11360 ( .A1(n12003), .A2(n13392), .ZN(n9617) );
  NAND2_X2 U11361 ( .A1(n13572), .A2(n13571), .ZN(n13570) );
  OAI21_X2 U11362 ( .B1(n15125), .B2(n12795), .A(n15120), .ZN(n14571) );
  NOR2_X2 U11363 ( .A1(n15127), .A2(n15126), .ZN(n15125) );
  INV_X1 U11364 ( .A(n9618), .ZN(n13790) );
  OAI22_X2 U11365 ( .A1(n18016), .A2(n17827), .B1(n17734), .B2(n18014), .ZN(
        n17717) );
  NAND2_X2 U11366 ( .A1(n18110), .A2(n18108), .ZN(n18052) );
  NOR2_X4 U11367 ( .A1(n13570), .A2(n13638), .ZN(n13639) );
  AND2_X2 U11368 ( .A1(n10225), .A2(n10205), .ZN(n10253) );
  OR2_X4 U11369 ( .A1(n15259), .A2(n15461), .ZN(n15454) );
  NAND2_X2 U11370 ( .A1(n11131), .A2(n10740), .ZN(n15259) );
  OR2_X1 U11371 ( .A1(n15217), .A2(n15216), .ZN(n15414) );
  AND2_X1 U11372 ( .A1(n12699), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10934) );
  AND2_X1 U11373 ( .A1(n14536), .A2(n14907), .ZN(n9619) );
  AND2_X1 U11374 ( .A1(n14906), .A2(n14907), .ZN(n14890) );
  INV_X1 U11375 ( .A(n20372), .ZN(n9620) );
  NAND2_X1 U11376 ( .A1(n11798), .A2(n11756), .ZN(n20371) );
  XNOR2_X1 U11377 ( .A(n11713), .B(n11711), .ZN(n11761) );
  NAND2_X2 U11378 ( .A1(n13840), .A2(n13839), .ZN(n14127) );
  INV_X4 U11379 ( .A(n10885), .ZN(n10173) );
  NAND2_X2 U11380 ( .A1(n9975), .A2(n9973), .ZN(n10885) );
  INV_X2 U11381 ( .A(n14840), .ZN(n14859) );
  AND2_X2 U11382 ( .A1(n14860), .A2(n14869), .ZN(n14840) );
  XNOR2_X2 U11383 ( .A(n10731), .B(n10729), .ZN(n14265) );
  NAND3_X2 U11384 ( .A1(n10725), .A2(n9963), .A3(n9962), .ZN(n10731) );
  NOR2_X2 U11385 ( .A1(n14571), .A2(n14570), .ZN(n14569) );
  NAND2_X2 U11386 ( .A1(n11716), .A2(n11636), .ZN(n11722) );
  NAND2_X2 U11387 ( .A1(n9938), .A2(n11620), .ZN(n11633) );
  INV_X4 U11388 ( .A(n11547), .ZN(n9938) );
  NAND2_X1 U11389 ( .A1(n11807), .A2(n11799), .ZN(n20730) );
  NOR2_X1 U11390 ( .A1(n16880), .A2(n11293), .ZN(n11306) );
  AND2_X1 U11391 ( .A1(n11487), .A2(n13377), .ZN(n9624) );
  AOI21_X2 U11392 ( .B1(n14481), .B2(n14608), .A(n14480), .ZN(n14835) );
  AND2_X1 U11393 ( .A1(n9815), .A2(n9715), .ZN(n14889) );
  NAND2_X2 U11394 ( .A1(n14397), .A2(n14396), .ZN(n14426) );
  XNOR2_X2 U11395 ( .A(n13711), .B(n13720), .ZN(n13710) );
  NAND2_X2 U11396 ( .A1(n13629), .A2(n13628), .ZN(n13711) );
  NAND2_X2 U11397 ( .A1(n20149), .A2(n11735), .ZN(n13348) );
  INV_X1 U11398 ( .A(n10059), .ZN(n9625) );
  INV_X4 U11399 ( .A(n10059), .ZN(n9626) );
  INV_X2 U11400 ( .A(n10059), .ZN(n15987) );
  AND2_X4 U11401 ( .A1(n13347), .A2(n11485), .ZN(n11492) );
  AND2_X1 U11402 ( .A1(n11483), .A2(n11487), .ZN(n9627) );
  AND2_X1 U11403 ( .A1(n11483), .A2(n11487), .ZN(n9628) );
  AND2_X1 U11404 ( .A1(n9793), .A2(n11485), .ZN(n9629) );
  AND2_X1 U11405 ( .A1(n9793), .A2(n11485), .ZN(n9630) );
  NAND2_X1 U11406 ( .A1(n12502), .A2(n12501), .ZN(n12527) );
  AND4_X1 U11407 ( .A1(n14046), .A2(n14059), .A3(n10184), .A4(n14014), .ZN(
        n9774) );
  OR2_X1 U11408 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20098), .ZN(
        n12330) );
  NAND2_X1 U11409 ( .A1(n13964), .A2(n16301), .ZN(n10127) );
  NAND2_X1 U11410 ( .A1(n9722), .A2(n10475), .ZN(n10726) );
  INV_X1 U11411 ( .A(n10477), .ZN(n9722) );
  NAND2_X1 U11412 ( .A1(n15837), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13906) );
  INV_X1 U11413 ( .A(n12043), .ZN(n12311) );
  NOR2_X1 U11414 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13895) );
  INV_X1 U11415 ( .A(n12319), .ZN(n12043) );
  AND2_X1 U11416 ( .A1(n14475), .A2(n14467), .ZN(n14466) );
  NAND2_X1 U11417 ( .A1(n14522), .A2(n14467), .ZN(n14472) );
  INV_X1 U11418 ( .A(n20756), .ZN(n10040) );
  NAND2_X2 U11419 ( .A1(n14146), .A2(n11784), .ZN(n12357) );
  INV_X1 U11420 ( .A(n11798), .ZN(n9937) );
  INV_X1 U11421 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9717) );
  INV_X1 U11422 ( .A(n15552), .ZN(n10004) );
  INV_X1 U11423 ( .A(n15635), .ZN(n10020) );
  NAND2_X1 U11424 ( .A1(n10728), .A2(n10423), .ZN(n10734) );
  INV_X1 U11425 ( .A(n10726), .ZN(n10728) );
  OAI21_X1 U11426 ( .B1(n15393), .B2(n16253), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n9969) );
  INV_X1 U11427 ( .A(n11164), .ZN(n11078) );
  NOR2_X1 U11428 ( .A1(n10901), .A2(n10900), .ZN(n10908) );
  NAND2_X1 U11429 ( .A1(n16328), .A2(n10173), .ZN(n13216) );
  OAI21_X1 U11430 ( .B1(n11372), .B2(n11371), .A(n12441), .ZN(n12997) );
  INV_X1 U11431 ( .A(n14589), .ZN(n14579) );
  INV_X1 U11432 ( .A(n19845), .ZN(n14598) );
  INV_X1 U11433 ( .A(n13574), .ZN(n14475) );
  XNOR2_X1 U11434 ( .A(n9626), .B(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14907) );
  OR2_X1 U11435 ( .A1(n11206), .A2(n15231), .ZN(n11207) );
  NAND2_X1 U11436 ( .A1(n10877), .A2(n19794), .ZN(n11164) );
  NAND2_X1 U11437 ( .A1(n15241), .A2(n9770), .ZN(n9769) );
  INV_X1 U11438 ( .A(n12458), .ZN(n9770) );
  XNOR2_X1 U11439 ( .A(n9769), .B(n9768), .ZN(n15227) );
  INV_X1 U11440 ( .A(n12459), .ZN(n9768) );
  NAND2_X1 U11441 ( .A1(n15510), .A2(n10740), .ZN(n15442) );
  NAND2_X1 U11442 ( .A1(n15280), .A2(n10577), .ZN(n9748) );
  NAND2_X1 U11443 ( .A1(n14273), .A2(n9683), .ZN(n15627) );
  NAND2_X1 U11444 ( .A1(n9777), .A2(n9774), .ZN(n19810) );
  NAND2_X2 U11445 ( .A1(n10118), .A2(n10117), .ZN(n13295) );
  INV_X1 U11446 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19528) );
  OR2_X1 U11447 ( .A1(n11375), .A2(n9830), .ZN(n9829) );
  NOR3_X1 U11448 ( .A1(n12425), .A2(n17292), .A3(n12434), .ZN(n11375) );
  AND2_X1 U11449 ( .A1(n15699), .A2(n18598), .ZN(n9830) );
  OAI21_X1 U11450 ( .B1(n16026), .B2(n14881), .A(n15001), .ZN(n9821) );
  AND2_X2 U11451 ( .A1(n11718), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9793) );
  NAND2_X1 U11452 ( .A1(n10371), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10010) );
  NOR2_X1 U11453 ( .A1(n10457), .A2(n10456), .ZN(n10461) );
  AOI21_X1 U11454 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n18641), .A(
        n11362), .ZN(n11363) );
  NOR2_X1 U11455 ( .A1(n11366), .A2(n11365), .ZN(n11362) );
  NAND2_X1 U11456 ( .A1(n11821), .A2(n9946), .ZN(n11871) );
  INV_X1 U11457 ( .A(n9801), .ZN(n9795) );
  NAND2_X1 U11458 ( .A1(n12327), .A2(n12326), .ZN(n12331) );
  OR3_X1 U11459 ( .A1(n12372), .A2(n12371), .A3(n12370), .ZN(n12373) );
  INV_X1 U11460 ( .A(n13550), .ZN(n15737) );
  INV_X1 U11461 ( .A(n10226), .ZN(n10230) );
  NAND2_X1 U11462 ( .A1(n10233), .A2(n10232), .ZN(n10234) );
  NAND2_X1 U11463 ( .A1(n10853), .A2(n10126), .ZN(n10215) );
  NOR2_X1 U11464 ( .A1(n10364), .A2(n9753), .ZN(n9752) );
  OR2_X1 U11465 ( .A1(n10347), .A2(n10346), .ZN(n10462) );
  NAND2_X1 U11466 ( .A1(n12678), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n9778) );
  NAND2_X1 U11467 ( .A1(n12677), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n9779) );
  NAND2_X1 U11468 ( .A1(n10267), .A2(n10282), .ZN(n10363) );
  NAND2_X1 U11469 ( .A1(n10284), .A2(n10278), .ZN(n10362) );
  NAND2_X1 U11470 ( .A1(n9781), .A2(n9780), .ZN(n10652) );
  NAND2_X1 U11471 ( .A1(n11252), .A2(n10658), .ZN(n9780) );
  OR2_X1 U11472 ( .A1(n10649), .A2(n9782), .ZN(n9781) );
  NOR2_X1 U11473 ( .A1(n17329), .A2(n12936), .ZN(n12957) );
  INV_X1 U11474 ( .A(n17326), .ZN(n12956) );
  NOR2_X1 U11475 ( .A1(n12331), .A2(n12330), .ZN(n12383) );
  AND2_X1 U11476 ( .A1(n14622), .A2(n14609), .ZN(n9950) );
  NOR2_X1 U11477 ( .A1(n14753), .A2(n9954), .ZN(n9953) );
  INV_X1 U11478 ( .A(n14357), .ZN(n9954) );
  NAND2_X1 U11479 ( .A1(n12011), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12314) );
  INV_X1 U11480 ( .A(n14092), .ZN(n9945) );
  INV_X1 U11481 ( .A(n13977), .ZN(n11895) );
  INV_X1 U11482 ( .A(n13895), .ZN(n12317) );
  CLKBUF_X1 U11483 ( .A(n13895), .Z(n12290) );
  NOR2_X1 U11484 ( .A1(n9893), .A2(n14745), .ZN(n9892) );
  NOR2_X1 U11485 ( .A1(n9896), .A2(n14304), .ZN(n9895) );
  INV_X1 U11486 ( .A(n14683), .ZN(n9896) );
  INV_X1 U11487 ( .A(n11872), .ZN(n9745) );
  NOR2_X1 U11488 ( .A1(n13985), .A2(n9890), .ZN(n9889) );
  INV_X1 U11489 ( .A(n14123), .ZN(n9890) );
  INV_X1 U11490 ( .A(n14466), .ZN(n14474) );
  AND3_X1 U11491 ( .A1(n11700), .A2(n11699), .A3(n11698), .ZN(n11711) );
  OR2_X1 U11492 ( .A1(n14146), .A2(n11683), .ZN(n11684) );
  NAND2_X1 U11493 ( .A1(n10046), .A2(n11679), .ZN(n11771) );
  NAND2_X1 U11494 ( .A1(n20105), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11784) );
  INV_X1 U11495 ( .A(n13469), .ZN(n13468) );
  AND2_X1 U11496 ( .A1(n9658), .A2(n9872), .ZN(n9871) );
  INV_X1 U11497 ( .A(n10509), .ZN(n10506) );
  AND2_X1 U11498 ( .A1(n12659), .A2(n9644), .ZN(n9847) );
  AND2_X1 U11499 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12503) );
  NAND2_X1 U11500 ( .A1(n10244), .A2(n10243), .ZN(n10742) );
  INV_X1 U11501 ( .A(n15135), .ZN(n9992) );
  NAND2_X1 U11502 ( .A1(n9995), .A2(n9994), .ZN(n9993) );
  INV_X1 U11503 ( .A(n12464), .ZN(n9995) );
  INV_X1 U11504 ( .A(n13071), .ZN(n9994) );
  INV_X1 U11505 ( .A(n13072), .ZN(n10008) );
  INV_X1 U11506 ( .A(n13087), .ZN(n9997) );
  AND2_X1 U11507 ( .A1(n13084), .A2(n15166), .ZN(n9986) );
  AND2_X1 U11508 ( .A1(n9979), .A2(n14030), .ZN(n9978) );
  INV_X1 U11509 ( .A(n14089), .ZN(n9979) );
  AND2_X1 U11510 ( .A1(n9982), .A2(n13747), .ZN(n9981) );
  INV_X1 U11511 ( .A(n10050), .ZN(n10030) );
  NAND2_X1 U11512 ( .A1(n14171), .A2(n14170), .ZN(n9755) );
  OR2_X1 U11513 ( .A1(n10360), .A2(n10359), .ZN(n10702) );
  NAND2_X2 U11514 ( .A1(n10184), .A2(n10212), .ZN(n10848) );
  OR2_X1 U11515 ( .A1(n12753), .A2(n12520), .ZN(n12521) );
  NOR2_X1 U11516 ( .A1(n10285), .A2(n13963), .ZN(n10011) );
  INV_X1 U11517 ( .A(n19380), .ZN(n10271) );
  AND4_X1 U11518 ( .A1(n10092), .A2(n10091), .A3(n10090), .A4(n10089), .ZN(
        n10097) );
  NOR2_X1 U11519 ( .A1(n11296), .A2(n16880), .ZN(n17107) );
  NOR2_X1 U11520 ( .A1(n11296), .A2(n11289), .ZN(n11403) );
  NAND2_X1 U11521 ( .A1(n12989), .A2(n16520), .ZN(n15700) );
  NAND2_X1 U11522 ( .A1(n9923), .A2(n9707), .ZN(n9922) );
  INV_X1 U11523 ( .A(n17512), .ZN(n9923) );
  INV_X1 U11524 ( .A(n9934), .ZN(n9932) );
  NAND2_X1 U11525 ( .A1(n12957), .A2(n12956), .ZN(n12960) );
  NAND2_X1 U11526 ( .A1(n12937), .A2(n13025), .ZN(n12936) );
  OR2_X1 U11527 ( .A1(n12992), .A2(n18609), .ZN(n12434) );
  NAND2_X1 U11528 ( .A1(n18169), .A2(n18173), .ZN(n18609) );
  OR3_X1 U11529 ( .A1(n20758), .A2(n13898), .A3(n13897), .ZN(n15837) );
  OR2_X1 U11530 ( .A1(n16141), .A2(n13896), .ZN(n13897) );
  AND2_X1 U11531 ( .A1(n20752), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12318) );
  AND2_X1 U11532 ( .A1(n13895), .A2(n14882), .ZN(n12197) );
  OR2_X1 U11533 ( .A1(n12180), .A2(n15858), .ZN(n12181) );
  NOR2_X1 U11534 ( .A1(n12027), .A2(n12026), .ZN(n12028) );
  NOR2_X1 U11535 ( .A1(n14840), .A2(n14415), .ZN(n14418) );
  NAND2_X1 U11536 ( .A1(n9743), .A2(n9741), .ZN(n14830) );
  NAND2_X1 U11537 ( .A1(n14417), .A2(n9744), .ZN(n9743) );
  NAND2_X1 U11538 ( .A1(n14859), .A2(n9742), .ZN(n9741) );
  INV_X1 U11539 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n9744) );
  NOR2_X1 U11540 ( .A1(n14635), .A2(n14619), .ZN(n14620) );
  OR2_X1 U11541 ( .A1(n15797), .A2(n14733), .ZN(n14735) );
  AND2_X1 U11542 ( .A1(n14371), .A2(n14370), .ZN(n14756) );
  AND2_X1 U11543 ( .A1(n14331), .A2(n14330), .ZN(n14332) );
  OR2_X1 U11544 ( .A1(n14317), .A2(n14316), .ZN(n15908) );
  INV_X1 U11545 ( .A(n13799), .ZN(n13796) );
  INV_X1 U11546 ( .A(n13798), .ZN(n13797) );
  OR2_X1 U11547 ( .A1(n11773), .A2(n10042), .ZN(n10036) );
  NOR2_X1 U11548 ( .A1(n10045), .A2(n10040), .ZN(n10038) );
  OR2_X1 U11549 ( .A1(n12377), .A2(n12350), .ZN(n12392) );
  AND2_X1 U11550 ( .A1(n9593), .A2(n20103), .ZN(n20456) );
  NOR2_X1 U11551 ( .A1(n20730), .A2(n20372), .ZN(n20457) );
  OR2_X1 U11552 ( .A1(n9593), .A2(n20103), .ZN(n20487) );
  NAND2_X1 U11553 ( .A1(n20756), .A2(n20104), .ZN(n20265) );
  NAND2_X1 U11554 ( .A1(n10616), .A2(n10617), .ZN(n10629) );
  INV_X1 U11555 ( .A(n11181), .ZN(n10616) );
  NOR2_X1 U11558 ( .A1(n16324), .A2(n16361), .ZN(n13102) );
  NOR2_X1 U11559 ( .A1(n12528), .A2(n9843), .ZN(n9842) );
  INV_X1 U11560 ( .A(n12525), .ZN(n9843) );
  AND2_X1 U11561 ( .A1(n12527), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12528) );
  INV_X1 U11562 ( .A(n11059), .ZN(n11161) );
  NOR2_X1 U11563 ( .A1(n11255), .A2(n11081), .ZN(n11166) );
  NAND2_X1 U11564 ( .A1(n10002), .A2(n9708), .ZN(n18999) );
  INV_X1 U11565 ( .A(n10909), .ZN(n9998) );
  AND2_X1 U11566 ( .A1(n9862), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9861) );
  INV_X1 U11567 ( .A(n10253), .ZN(n10256) );
  NOR2_X1 U11568 ( .A1(n10624), .A2(n10013), .ZN(n10626) );
  OR2_X1 U11569 ( .A1(n15442), .A2(n11095), .ZN(n12480) );
  OR2_X1 U11570 ( .A1(n13067), .A2(n10733), .ZN(n12459) );
  INV_X1 U11571 ( .A(n10012), .ZN(n9772) );
  INV_X1 U11572 ( .A(n10603), .ZN(n9773) );
  NAND2_X1 U11573 ( .A1(n10602), .A2(n10603), .ZN(n15249) );
  NAND2_X1 U11574 ( .A1(n15295), .A2(n9863), .ZN(n10587) );
  AND2_X1 U11575 ( .A1(n11102), .A2(n9864), .ZN(n9863) );
  NOR2_X1 U11576 ( .A1(n9865), .A2(n11107), .ZN(n9864) );
  NOR2_X1 U11577 ( .A1(n15522), .A2(n11094), .ZN(n15510) );
  AND2_X1 U11578 ( .A1(n11058), .A2(n11057), .ZN(n15552) );
  NOR2_X1 U11579 ( .A1(n15601), .A2(n15582), .ZN(n14200) );
  AND2_X1 U11580 ( .A1(n14200), .A2(n9678), .ZN(n15555) );
  NAND2_X1 U11581 ( .A1(n10870), .A2(n14269), .ZN(n15534) );
  NAND2_X1 U11582 ( .A1(n15615), .A2(n15602), .ZN(n15601) );
  INV_X1 U11583 ( .A(n14266), .ZN(n10023) );
  INV_X1 U11584 ( .A(n10026), .ZN(n10025) );
  OAI21_X1 U11585 ( .B1(n10050), .B2(n10027), .A(n10528), .ZN(n10026) );
  NAND2_X1 U11586 ( .A1(n10028), .A2(n16254), .ZN(n10027) );
  INV_X1 U11587 ( .A(n15641), .ZN(n10005) );
  AND2_X1 U11588 ( .A1(n10955), .A2(n13803), .ZN(n10006) );
  AND2_X1 U11589 ( .A1(n15344), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15624) );
  OR2_X1 U11590 ( .A1(n10734), .A2(n10733), .ZN(n10735) );
  INV_X1 U11591 ( .A(n10736), .ZN(n15393) );
  NAND2_X1 U11592 ( .A1(n10932), .A2(n10063), .ZN(n14273) );
  NAND2_X1 U11593 ( .A1(n10721), .A2(n10720), .ZN(n10725) );
  NAND2_X2 U11594 ( .A1(n10173), .A2(n19823), .ZN(n19809) );
  NAND2_X1 U11595 ( .A1(n10701), .A2(n19673), .ZN(n11088) );
  NAND2_X1 U11596 ( .A1(n12506), .A2(n12505), .ZN(n13299) );
  XNOR2_X1 U11597 ( .A(n12523), .B(n12521), .ZN(n13516) );
  NAND2_X1 U11598 ( .A1(n19076), .A2(n19796), .ZN(n19312) );
  OR2_X1 U11599 ( .A1(n19782), .A2(n14180), .ZN(n19487) );
  NOR2_X2 U11600 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19764) );
  NAND2_X1 U11601 ( .A1(n19782), .A2(n14180), .ZN(n19562) );
  NAND2_X1 U11602 ( .A1(n10168), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10107) );
  OR2_X1 U11603 ( .A1(n19076), .A2(n19796), .ZN(n19488) );
  NAND2_X1 U11604 ( .A1(n11117), .A2(n11116), .ZN(n19533) );
  NOR2_X1 U11605 ( .A1(n14040), .A2(n14039), .ZN(n14045) );
  NAND2_X1 U11606 ( .A1(n9790), .A2(n10654), .ZN(n16328) );
  INV_X1 U11607 ( .A(n10655), .ZN(n9790) );
  NAND2_X1 U11608 ( .A1(n12997), .A2(n12998), .ZN(n18596) );
  NOR2_X1 U11609 ( .A1(n16549), .A2(n16547), .ZN(n16548) );
  NAND2_X1 U11610 ( .A1(n16668), .A2(n9904), .ZN(n16647) );
  NAND2_X1 U11611 ( .A1(n16805), .A2(n9905), .ZN(n9904) );
  INV_X1 U11612 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n9905) );
  NAND2_X1 U11613 ( .A1(n9829), .A2(n9681), .ZN(n11397) );
  NOR2_X1 U11614 ( .A1(n11293), .A2(n18618), .ZN(n11327) );
  INV_X1 U11615 ( .A(n18160), .ZN(n18814) );
  AND2_X1 U11616 ( .A1(n13003), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12421) );
  NOR2_X1 U11617 ( .A1(n17467), .A2(n17468), .ZN(n13000) );
  NOR2_X1 U11618 ( .A1(n17586), .A2(n9902), .ZN(n9901) );
  NOR2_X1 U11619 ( .A1(n17618), .A2(n17619), .ZN(n17605) );
  NAND2_X1 U11620 ( .A1(n9913), .A2(n9907), .ZN(n17618) );
  AND2_X1 U11621 ( .A1(n16721), .A2(n9908), .ZN(n9907) );
  NOR2_X1 U11622 ( .A1(n9910), .A2(n9909), .ZN(n9908) );
  NAND2_X1 U11623 ( .A1(n9912), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n9909) );
  OAI22_X1 U11624 ( .A1(n15777), .A2(n16393), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n17656), .ZN(n9919) );
  NOR2_X1 U11625 ( .A1(n9928), .A2(n9634), .ZN(n12964) );
  INV_X1 U11626 ( .A(n9929), .ZN(n9927) );
  NOR2_X1 U11627 ( .A1(n9634), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n9929) );
  NOR2_X1 U11628 ( .A1(n17730), .A2(n18063), .ZN(n17729) );
  AOI21_X1 U11629 ( .B1(n11374), .B2(n11373), .A(n12997), .ZN(n18598) );
  NAND2_X1 U11630 ( .A1(n19840), .A2(n19841), .ZN(n20758) );
  NAND2_X1 U11631 ( .A1(n16021), .A2(n14882), .ZN(n9822) );
  OR2_X1 U11632 ( .A1(n20093), .A2(n13404), .ZN(n16026) );
  INV_X1 U11633 ( .A(n16022), .ZN(n20102) );
  INV_X1 U11634 ( .A(n16068), .ZN(n16142) );
  OR2_X1 U11635 ( .A1(n20729), .A2(n20343), .ZN(n20370) );
  AND2_X1 U11636 ( .A1(n15760), .A2(n15759), .ZN(n15775) );
  NAND2_X1 U11637 ( .A1(n9835), .A2(n9834), .ZN(n16168) );
  NAND2_X1 U11638 ( .A1(n9838), .A2(n11249), .ZN(n9834) );
  OR2_X1 U11639 ( .A1(n16183), .A2(n11247), .ZN(n9835) );
  NOR2_X1 U11642 ( .A1(n16194), .A2(n11247), .ZN(n13066) );
  NOR2_X1 U11643 ( .A1(n13080), .A2(n11247), .ZN(n13052) );
  OR2_X1 U11644 ( .A1(n11258), .A2(n11257), .ZN(n18984) );
  INV_X1 U11645 ( .A(n19796), .ZN(n19030) );
  XNOR2_X1 U11646 ( .A(n11159), .B(n11158), .ZN(n14392) );
  AND2_X1 U11647 ( .A1(n15074), .A2(n9990), .ZN(n11159) );
  XNOR2_X1 U11648 ( .A(n9718), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n12494) );
  NAND2_X1 U11649 ( .A1(n15216), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9718) );
  AND2_X1 U11650 ( .A1(n16193), .A2(n16290), .ZN(n9881) );
  INV_X1 U11651 ( .A(n19179), .ZN(n16290) );
  INV_X1 U11652 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18661) );
  NOR2_X2 U11653 ( .A1(n18763), .A2(n16862), .ZN(n16876) );
  INV_X1 U11654 ( .A(n16848), .ZN(n16887) );
  NOR3_X1 U11655 ( .A1(n16898), .A2(n16897), .A3(n16942), .ZN(n16935) );
  NOR2_X1 U11656 ( .A1(n17009), .A2(n17011), .ZN(n16996) );
  AND2_X1 U11657 ( .A1(n17292), .A2(n17206), .ZN(n17203) );
  NAND2_X1 U11658 ( .A1(n17218), .A2(n17340), .ZN(n9735) );
  OR2_X1 U11659 ( .A1(n17349), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n9734) );
  INV_X1 U11660 ( .A(n17218), .ZN(n17214) );
  NAND2_X1 U11661 ( .A1(n17223), .A2(P3_EAX_REG_29__SCAN_IN), .ZN(n17218) );
  INV_X1 U11662 ( .A(n17256), .ZN(n17283) );
  NAND2_X1 U11663 ( .A1(n18630), .A2(n17207), .ZN(n17342) );
  NAND2_X1 U11664 ( .A1(n17207), .A2(P3_EAX_REG_1__SCAN_IN), .ZN(n17350) );
  NAND2_X1 U11665 ( .A1(n12345), .A2(n10056), .ZN(n13254) );
  NAND2_X1 U11666 ( .A1(n10455), .A2(n10454), .ZN(n10457) );
  OR2_X1 U11667 ( .A1(n10453), .A2(n10452), .ZN(n10455) );
  OAI21_X1 U11668 ( .B1(n12780), .B2(n9784), .A(n9783), .ZN(n9782) );
  NAND2_X1 U11669 ( .A1(n9785), .A2(n10659), .ZN(n9784) );
  AOI21_X1 U11670 ( .B1(n11252), .B2(n10644), .A(n10658), .ZN(n9783) );
  INV_X1 U11671 ( .A(n19830), .ZN(n9785) );
  INV_X1 U11672 ( .A(n12355), .ZN(n12337) );
  NOR2_X1 U11673 ( .A1(n11845), .A2(n9947), .ZN(n9946) );
  OR2_X1 U11674 ( .A1(n11844), .A2(n11843), .ZN(n13844) );
  OR2_X1 U11675 ( .A1(n11697), .A2(n11696), .ZN(n13470) );
  INV_X1 U11676 ( .A(n14151), .ZN(n11683) );
  NAND2_X1 U11677 ( .A1(n20105), .A2(n13426), .ZN(n11640) );
  NOR2_X1 U11678 ( .A1(n13400), .A2(n14596), .ZN(n13279) );
  INV_X1 U11679 ( .A(n11481), .ZN(n9812) );
  AND3_X1 U11680 ( .A1(n16339), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A3(
        n10640), .ZN(n10651) );
  INV_X1 U11681 ( .A(n10237), .ZN(n9766) );
  AND2_X1 U11682 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11124) );
  NOR2_X1 U11683 ( .A1(n10629), .A2(n10628), .ZN(n10633) );
  INV_X1 U11684 ( .A(n10597), .ZN(n10017) );
  NAND2_X1 U11685 ( .A1(n10198), .A2(n19829), .ZN(n10194) );
  AND2_X1 U11686 ( .A1(n13025), .A2(n13024), .ZN(n13009) );
  AOI21_X1 U11687 ( .B1(n18178), .B2(n12437), .A(n12993), .ZN(n12426) );
  AOI21_X1 U11688 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18636), .A(
        n11360), .ZN(n11366) );
  NAND2_X1 U11689 ( .A1(n9731), .A2(n18169), .ZN(n12993) );
  NAND2_X1 U11690 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18768), .ZN(
        n11296) );
  INV_X1 U11691 ( .A(n12314), .ZN(n12287) );
  NOR2_X1 U11692 ( .A1(n9952), .A2(n14747), .ZN(n9951) );
  INV_X1 U11693 ( .A(n9953), .ZN(n9952) );
  INV_X1 U11694 ( .A(n14149), .ZN(n11875) );
  NOR2_X1 U11695 ( .A1(n11801), .A2(n11800), .ZN(n11825) );
  INV_X1 U11696 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11800) );
  NOR2_X1 U11697 ( .A1(n14415), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9742) );
  INV_X1 U11698 ( .A(n14713), .ZN(n9900) );
  OR2_X1 U11699 ( .A1(n14721), .A2(n14728), .ZN(n9899) );
  INV_X1 U11700 ( .A(n14398), .ZN(n9818) );
  NOR2_X1 U11701 ( .A1(n15987), .A2(n14400), .ZN(n10049) );
  INV_X1 U11702 ( .A(n14399), .ZN(n9817) );
  NAND2_X1 U11703 ( .A1(n14953), .A2(n14399), .ZN(n14940) );
  NAND2_X1 U11704 ( .A1(n13399), .A2(n13398), .ZN(n9804) );
  NAND2_X1 U11705 ( .A1(n13411), .A2(n13410), .ZN(n13413) );
  INV_X1 U11706 ( .A(n11770), .ZN(n10045) );
  AOI21_X1 U11707 ( .B1(n13175), .B2(n11646), .A(n11645), .ZN(n11649) );
  NAND2_X1 U11708 ( .A1(n11724), .A2(n11723), .ZN(n11730) );
  AND2_X1 U11709 ( .A1(n12329), .A2(n12330), .ZN(n12351) );
  OR2_X1 U11710 ( .A1(n12331), .A2(n12328), .ZN(n12329) );
  AOI21_X1 U11711 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n20756), .A(
        n12388), .ZN(n12389) );
  NAND2_X1 U11712 ( .A1(n12385), .A2(n14145), .ZN(n12377) );
  INV_X1 U11713 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20424) );
  OAI21_X1 U11714 ( .B1(n13556), .B2(n16159), .A(n15767), .ZN(n20104) );
  INV_X1 U11715 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20488) );
  AND2_X1 U11716 ( .A1(n10676), .A2(n10675), .ZN(n10868) );
  NAND2_X1 U11717 ( .A1(n19809), .A2(n10659), .ZN(n10447) );
  NAND2_X1 U11718 ( .A1(n10559), .A2(n10609), .ZN(n10556) );
  NOR2_X1 U11719 ( .A1(n10564), .A2(n9874), .ZN(n9873) );
  INV_X1 U11720 ( .A(n10536), .ZN(n9874) );
  NAND2_X1 U11721 ( .A1(n10530), .A2(n13749), .ZN(n10538) );
  AND2_X1 U11722 ( .A1(n10529), .A2(n13739), .ZN(n10530) );
  NAND2_X1 U11723 ( .A1(n10450), .A2(n10449), .ZN(n10487) );
  NAND2_X1 U11724 ( .A1(n12848), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10449) );
  NAND2_X1 U11725 ( .A1(n10680), .A2(n10886), .ZN(n10450) );
  INV_X1 U11726 ( .A(n12753), .ZN(n12776) );
  NAND2_X1 U11727 ( .A1(n12497), .A2(n13295), .ZN(n12753) );
  NOR2_X1 U11728 ( .A1(n12780), .A2(n19822), .ZN(n12497) );
  OR2_X1 U11729 ( .A1(n10388), .A2(n10387), .ZN(n10922) );
  NOR2_X1 U11730 ( .A1(n11207), .A2(n11203), .ZN(n11204) );
  AND2_X1 U11731 ( .A1(n9682), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9862) );
  NOR2_X1 U11732 ( .A1(n9635), .A2(n9853), .ZN(n9852) );
  NOR2_X1 U11733 ( .A1(n16245), .A2(n9855), .ZN(n9854) );
  AND2_X1 U11734 ( .A1(n11123), .A2(n11234), .ZN(n11231) );
  NAND2_X1 U11735 ( .A1(n15417), .A2(n10014), .ZN(n10013) );
  INV_X1 U11736 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n10014) );
  INV_X1 U11737 ( .A(n15190), .ZN(n10009) );
  NAND2_X1 U11738 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n9971) );
  NAND2_X1 U11739 ( .A1(n14255), .A2(n9700), .ZN(n13089) );
  AND2_X1 U11740 ( .A1(n11061), .A2(n11060), .ZN(n11136) );
  INV_X1 U11741 ( .A(n10510), .ZN(n10028) );
  AND2_X1 U11742 ( .A1(n10434), .A2(n10433), .ZN(n10440) );
  AND4_X1 U11743 ( .A1(n10427), .A2(n10426), .A3(n10425), .A4(n10424), .ZN(
        n10442) );
  AND4_X1 U11744 ( .A1(n10438), .A2(n10437), .A3(n10436), .A4(n10435), .ZN(
        n10439) );
  OR2_X1 U11745 ( .A1(n10734), .A2(n10732), .ZN(n10736) );
  INV_X1 U11746 ( .A(n13648), .ZN(n9987) );
  NOR2_X1 U11747 ( .A1(n10909), .A2(n9999), .ZN(n10001) );
  NAND2_X1 U11748 ( .A1(n10000), .A2(n13768), .ZN(n9999) );
  INV_X1 U11749 ( .A(n19000), .ZN(n10000) );
  AND2_X1 U11750 ( .A1(n10762), .A2(n9989), .ZN(n9988) );
  INV_X1 U11751 ( .A(n13587), .ZN(n9989) );
  NAND2_X1 U11752 ( .A1(n9964), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9963) );
  INV_X1 U11753 ( .A(n10724), .ZN(n9964) );
  OR2_X1 U11754 ( .A1(n10926), .A2(n10925), .ZN(n10928) );
  OR2_X1 U11755 ( .A1(n10419), .A2(n10418), .ZN(n10929) );
  INV_X1 U11756 ( .A(n13505), .ZN(n10762) );
  AND2_X1 U11757 ( .A1(n10333), .A2(n10361), .ZN(n9721) );
  INV_X1 U11758 ( .A(n9958), .ZN(n9957) );
  XNOR2_X1 U11759 ( .A(n10477), .B(n10712), .ZN(n10718) );
  INV_X1 U11760 ( .A(n10475), .ZN(n10712) );
  OR2_X1 U11761 ( .A1(n13340), .A2(n10708), .ZN(n10709) );
  NAND2_X1 U11762 ( .A1(n10334), .A2(n10333), .ZN(n10711) );
  NOR2_X2 U11763 ( .A1(n10487), .A2(n10495), .ZN(n10486) );
  AND3_X1 U11764 ( .A1(n10460), .A2(n10459), .A3(n10458), .ZN(n10484) );
  OR2_X1 U11765 ( .A1(n10319), .A2(n10318), .ZN(n10884) );
  NAND2_X1 U11766 ( .A1(n12678), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n9961) );
  AOI21_X1 U11767 ( .B1(n12677), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A(
        n16304), .ZN(n9960) );
  OR2_X1 U11768 ( .A1(n10893), .A2(n10892), .ZN(n10899) );
  NAND2_X1 U11769 ( .A1(n12860), .A2(n19794), .ZN(n11059) );
  INV_X1 U11770 ( .A(n12518), .ZN(n12510) );
  OAI21_X1 U11771 ( .B1(n13295), .B2(n19822), .A(n19794), .ZN(n12516) );
  AND2_X1 U11772 ( .A1(n10259), .A2(n10258), .ZN(n10282) );
  NAND2_X1 U11773 ( .A1(n10143), .A2(n16304), .ZN(n10174) );
  NAND2_X1 U11774 ( .A1(n10148), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10175) );
  NAND2_X1 U11775 ( .A1(n10284), .A2(n10276), .ZN(n19564) );
  NAND2_X1 U11776 ( .A1(n9792), .A2(n9791), .ZN(n10655) );
  NAND2_X1 U11777 ( .A1(n16339), .A2(n19822), .ZN(n9791) );
  NAND2_X1 U11778 ( .A1(n10653), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n9792) );
  NAND2_X1 U11779 ( .A1(n18160), .A2(n9732), .ZN(n9731) );
  NAND2_X1 U11780 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18793), .ZN(
        n11294) );
  NAND2_X1 U11781 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11361), .ZN(
        n11292) );
  INV_X1 U11782 ( .A(n11291), .ZN(n9729) );
  INV_X1 U11783 ( .A(n16880), .ZN(n9730) );
  NOR2_X1 U11784 ( .A1(n11294), .A2(n11292), .ZN(n11349) );
  NAND2_X1 U11785 ( .A1(n18768), .A2(n11361), .ZN(n11293) );
  NAND2_X1 U11786 ( .A1(n10062), .A2(n9935), .ZN(n9934) );
  NOR2_X1 U11787 ( .A1(n17729), .A2(n18055), .ZN(n16366) );
  NAND2_X1 U11788 ( .A1(n17750), .A2(n12959), .ZN(n12961) );
  INV_X1 U11789 ( .A(n15837), .ZN(n15918) );
  NAND2_X1 U11790 ( .A1(n13915), .A2(n15761), .ZN(n15911) );
  AND2_X1 U11791 ( .A1(n13982), .A2(n13981), .ZN(n13984) );
  AND2_X1 U11792 ( .A1(n14815), .A2(n13415), .ZN(n13418) );
  NAND2_X1 U11793 ( .A1(n9665), .A2(n12003), .ZN(n11852) );
  AND2_X1 U11794 ( .A1(n11630), .A2(n11631), .ZN(n13417) );
  AND2_X1 U11795 ( .A1(n12292), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13899) );
  AND2_X1 U11796 ( .A1(n9950), .A2(n9949), .ZN(n9948) );
  INV_X1 U11797 ( .A(n14481), .ZN(n9949) );
  NOR2_X1 U11798 ( .A1(n12265), .A2(n14864), .ZN(n12266) );
  NOR2_X1 U11799 ( .A1(n12140), .A2(n15823), .ZN(n12115) );
  NAND2_X1 U11800 ( .A1(n12115), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12218) );
  NOR2_X1 U11801 ( .A1(n12176), .A2(n15845), .ZN(n12141) );
  NAND2_X1 U11802 ( .A1(n12141), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12140) );
  AND2_X1 U11803 ( .A1(n14891), .A2(n15025), .ZN(n9740) );
  AND2_X1 U11804 ( .A1(n12080), .A2(n12079), .ZN(n14738) );
  NOR2_X1 U11805 ( .A1(n12060), .A2(n14927), .ZN(n12062) );
  AND2_X1 U11806 ( .A1(n14358), .A2(n9951), .ZN(n14748) );
  NAND2_X1 U11807 ( .A1(n14358), .A2(n9953), .ZN(n14754) );
  AND2_X1 U11808 ( .A1(n12030), .A2(n12029), .ZN(n14357) );
  NAND2_X1 U11809 ( .A1(n14358), .A2(n14357), .ZN(n14752) );
  NAND2_X1 U11810 ( .A1(n11994), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12027) );
  INV_X1 U11811 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12026) );
  NOR2_X1 U11812 ( .A1(n11978), .A2(n14687), .ZN(n11994) );
  NAND2_X1 U11813 ( .A1(n14678), .A2(n11977), .ZN(n14680) );
  AND2_X1 U11814 ( .A1(n11928), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11929) );
  NOR2_X1 U11815 ( .A1(n14315), .A2(n14314), .ZN(n14676) );
  NOR2_X1 U11816 ( .A1(n11912), .A2(n11911), .ZN(n11928) );
  AOI21_X1 U11817 ( .B1(n19871), .B2(n13895), .A(n11910), .ZN(n14092) );
  CLKBUF_X1 U11818 ( .A(n14094), .Z(n14095) );
  AND3_X1 U11819 ( .A1(n11894), .A2(n11893), .A3(n11892), .ZN(n13977) );
  NAND2_X1 U11820 ( .A1(n11876), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11896) );
  NAND2_X1 U11821 ( .A1(n11880), .A2(n9618), .ZN(n13875) );
  AND2_X1 U11822 ( .A1(n11863), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n11876) );
  NAND2_X1 U11823 ( .A1(n13639), .A2(n13725), .ZN(n9940) );
  AND2_X1 U11824 ( .A1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n11825), .ZN(
        n11848) );
  NAND2_X1 U11825 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n11801) );
  AOI21_X1 U11826 ( .B1(n11760), .B2(n11975), .A(n9944), .ZN(n9943) );
  INV_X1 U11827 ( .A(n11779), .ZN(n9944) );
  NAND2_X1 U11828 ( .A1(n14672), .A2(n14647), .ZN(n14649) );
  OR2_X1 U11829 ( .A1(n14649), .A2(n14633), .ZN(n14635) );
  NOR2_X1 U11830 ( .A1(n14735), .A2(n9897), .ZN(n14672) );
  OR3_X1 U11831 ( .A1(n9899), .A2(n9900), .A3(n9898), .ZN(n9897) );
  INV_X1 U11832 ( .A(n14670), .ZN(n9898) );
  NOR3_X1 U11833 ( .A1(n14735), .A2(n9899), .A3(n9900), .ZN(n14715) );
  NOR2_X1 U11834 ( .A1(n14735), .A2(n9899), .ZN(n14722) );
  AND2_X1 U11835 ( .A1(n14452), .A2(n14451), .ZN(n14733) );
  INV_X1 U11836 ( .A(n15800), .ZN(n9891) );
  NAND2_X1 U11837 ( .A1(n14756), .A2(n9646), .ZN(n15799) );
  NAND2_X1 U11838 ( .A1(n14756), .A2(n14757), .ZN(n14760) );
  AND2_X1 U11839 ( .A1(n15910), .A2(n9690), .ZN(n14371) );
  INV_X1 U11840 ( .A(n14332), .ZN(n9894) );
  NAND2_X1 U11841 ( .A1(n15910), .A2(n9895), .ZN(n14333) );
  NOR2_X1 U11842 ( .A1(n15908), .A2(n15907), .ZN(n15910) );
  NAND2_X1 U11843 ( .A1(n15910), .A2(n14683), .ZN(n14682) );
  AND2_X1 U11844 ( .A1(n14295), .A2(n14294), .ZN(n14316) );
  INV_X1 U11845 ( .A(n14167), .ZN(n9887) );
  NAND2_X1 U11846 ( .A1(n9888), .A2(n9889), .ZN(n14166) );
  NOR2_X1 U11847 ( .A1(n13986), .A2(n13985), .ZN(n14124) );
  NOR2_X1 U11848 ( .A1(n13582), .A2(n9884), .ZN(n9883) );
  INV_X1 U11849 ( .A(n13786), .ZN(n9884) );
  NOR2_X1 U11850 ( .A1(n9885), .A2(n13582), .ZN(n13787) );
  NAND2_X1 U11851 ( .A1(n13488), .A2(n13580), .ZN(n13645) );
  INV_X1 U11852 ( .A(n13582), .ZN(n13488) );
  AND2_X1 U11853 ( .A1(n15057), .A2(n15055), .ZN(n16131) );
  NAND2_X1 U11854 ( .A1(n10044), .A2(n11770), .ZN(n10043) );
  NAND2_X1 U11855 ( .A1(n10041), .A2(n10040), .ZN(n10039) );
  INV_X1 U11856 ( .A(n11679), .ZN(n10044) );
  NAND2_X1 U11857 ( .A1(n11639), .A2(n11638), .ZN(n9936) );
  NAND2_X1 U11858 ( .A1(n11722), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11639) );
  OR2_X1 U11859 ( .A1(n11713), .A2(n11712), .ZN(n11714) );
  XNOR2_X1 U11860 ( .A(n11753), .B(n11752), .ZN(n11755) );
  OAI22_X1 U11861 ( .A1(n13421), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n13468), 
        .B2(n14146), .ZN(n11753) );
  NAND2_X1 U11862 ( .A1(n20735), .A2(n20756), .ZN(n11796) );
  AND3_X1 U11863 ( .A1(n13370), .A2(n13369), .A3(n13368), .ZN(n13550) );
  INV_X1 U11864 ( .A(n20456), .ZN(n20343) );
  AOI21_X1 U11865 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20519), .A(n20265), 
        .ZN(n20606) );
  OR2_X1 U11866 ( .A1(n20603), .A2(n20343), .ZN(n20107) );
  INV_X1 U11867 ( .A(n14561), .ZN(n15767) );
  OR2_X1 U11868 ( .A1(n16183), .A2(n11247), .ZN(n9837) );
  NOR2_X1 U11869 ( .A1(n13065), .A2(n11247), .ZN(n16184) );
  NAND2_X1 U11870 ( .A1(n10573), .A2(n10572), .ZN(n10593) );
  NOR2_X2 U11871 ( .A1(n10548), .A2(n10543), .ZN(n10550) );
  NAND2_X1 U11872 ( .A1(n10556), .A2(n10554), .ZN(n10546) );
  NAND2_X1 U11873 ( .A1(n10537), .A2(n9658), .ZN(n10557) );
  NOR2_X1 U11874 ( .A1(n18911), .A2(n11243), .ZN(n14203) );
  NAND2_X1 U11875 ( .A1(n14203), .A2(n14202), .ZN(n18896) );
  NAND2_X1 U11876 ( .A1(n18947), .A2(n18950), .ZN(n18928) );
  NAND2_X1 U11877 ( .A1(n13801), .A2(n15395), .ZN(n18954) );
  NOR2_X1 U11878 ( .A1(n18961), .A2(n18963), .ZN(n13801) );
  NAND2_X1 U11879 ( .A1(n10506), .A2(n9875), .ZN(n9876) );
  NOR2_X1 U11880 ( .A1(n10507), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n9875) );
  NAND2_X1 U11881 ( .A1(n9880), .A2(n9878), .ZN(n10514) );
  AND2_X1 U11882 ( .A1(n10506), .A2(n9879), .ZN(n9878) );
  NAND2_X1 U11883 ( .A1(n18987), .A2(n18990), .ZN(n13752) );
  NOR2_X1 U11884 ( .A1(n19007), .A2(n19140), .ZN(n18987) );
  NAND2_X1 U11885 ( .A1(n13765), .A2(n13766), .ZN(n19007) );
  NOR2_X1 U11886 ( .A1(n13831), .A2(n13687), .ZN(n13765) );
  AND2_X1 U11887 ( .A1(n9703), .A2(n9984), .ZN(n9983) );
  INV_X1 U11888 ( .A(n15151), .ZN(n9984) );
  NOR2_X1 U11889 ( .A1(n13929), .A2(n13928), .ZN(n12535) );
  OR2_X1 U11890 ( .A1(n10966), .A2(n10965), .ZN(n13655) );
  NOR2_X1 U11891 ( .A1(n9840), .A2(n12529), .ZN(n9839) );
  INV_X1 U11892 ( .A(n15119), .ZN(n12795) );
  AND2_X1 U11893 ( .A1(n15458), .A2(n9711), .ZN(n12476) );
  INV_X1 U11894 ( .A(n12474), .ZN(n10007) );
  OR2_X1 U11895 ( .A1(n9847), .A2(n12718), .ZN(n9845) );
  AND2_X1 U11896 ( .A1(n9847), .A2(n12718), .ZN(n9846) );
  AND2_X1 U11897 ( .A1(n19069), .A2(n12861), .ZN(n13301) );
  AND2_X1 U11898 ( .A1(n13217), .A2(n19828), .ZN(n19109) );
  OAI21_X1 U11899 ( .B1(n12858), .B2(n12857), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13190) );
  INV_X1 U11900 ( .A(n13190), .ZN(n13863) );
  OAI21_X1 U11901 ( .B1(n11207), .B2(n9850), .A(n11202), .ZN(n9849) );
  NAND2_X1 U11902 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n11201), .ZN(
        n9850) );
  AND2_X1 U11903 ( .A1(n11190), .A2(n9862), .ZN(n11212) );
  AND2_X1 U11904 ( .A1(n11119), .A2(n15166), .ZN(n15168) );
  OR2_X1 U11905 ( .A1(n18900), .A2(n10560), .ZN(n15330) );
  NAND2_X1 U11906 ( .A1(n15346), .A2(n10064), .ZN(n15331) );
  AND2_X1 U11907 ( .A1(n14031), .A2(n9693), .ZN(n14244) );
  INV_X1 U11908 ( .A(n14234), .ZN(n9977) );
  NOR2_X1 U11909 ( .A1(n11228), .A2(n9635), .ZN(n11245) );
  NAND2_X1 U11910 ( .A1(n9851), .A2(n9854), .ZN(n11244) );
  NAND2_X1 U11911 ( .A1(n13746), .A2(n9684), .ZN(n13932) );
  INV_X1 U11912 ( .A(n13889), .ZN(n9980) );
  NOR2_X1 U11913 ( .A1(n13658), .A2(n13734), .ZN(n13746) );
  INV_X1 U11914 ( .A(n11231), .ZN(n11239) );
  AOI21_X1 U11915 ( .B1(n10747), .B2(n10746), .A(n10745), .ZN(n13599) );
  AND2_X1 U11916 ( .A1(n13599), .A2(n13598), .ZN(n13607) );
  INV_X1 U11917 ( .A(n10248), .ZN(n10249) );
  NOR2_X1 U11918 ( .A1(n9991), .A2(n9709), .ZN(n9990) );
  OR2_X1 U11919 ( .A1(n9993), .A2(n9992), .ZN(n9991) );
  INV_X1 U11920 ( .A(n10828), .ZN(n11157) );
  NOR2_X1 U11921 ( .A1(n15137), .A2(n9993), .ZN(n12466) );
  NAND2_X1 U11922 ( .A1(n15458), .A2(n9701), .ZN(n15192) );
  NAND2_X1 U11923 ( .A1(n15458), .A2(n9702), .ZN(n13074) );
  OR2_X1 U11924 ( .A1(n9971), .A2(n15417), .ZN(n9970) );
  OR2_X1 U11925 ( .A1(n15137), .A2(n13071), .ZN(n13069) );
  AND2_X1 U11926 ( .A1(n14255), .A2(n9710), .ZN(n15456) );
  INV_X1 U11927 ( .A(n13059), .ZN(n9996) );
  AND2_X1 U11928 ( .A1(n15456), .A2(n15455), .ZN(n15458) );
  NAND2_X1 U11929 ( .A1(n15267), .A2(n15268), .ZN(n9747) );
  NAND2_X1 U11930 ( .A1(n11119), .A2(n9703), .ZN(n15152) );
  AND2_X1 U11931 ( .A1(n15313), .A2(n15266), .ZN(n15277) );
  NOR2_X1 U11932 ( .A1(n11137), .A2(n11136), .ZN(n14255) );
  NAND2_X1 U11933 ( .A1(n9866), .A2(n10582), .ZN(n15295) );
  INV_X1 U11934 ( .A(n18863), .ZN(n9866) );
  NAND2_X1 U11935 ( .A1(n15542), .A2(n9714), .ZN(n15522) );
  AND2_X1 U11936 ( .A1(n14200), .A2(n9694), .ZN(n15100) );
  INV_X1 U11937 ( .A(n15101), .ZN(n10003) );
  NAND2_X1 U11938 ( .A1(n14200), .A2(n9645), .ZN(n15102) );
  NOR2_X1 U11939 ( .A1(n15570), .A2(n15573), .ZN(n15542) );
  NOR2_X1 U11940 ( .A1(n15627), .A2(n15616), .ZN(n15615) );
  NAND2_X1 U11941 ( .A1(n13746), .A2(n9981), .ZN(n13888) );
  NAND2_X1 U11942 ( .A1(n13746), .A2(n13747), .ZN(n13817) );
  AOI21_X1 U11943 ( .B1(n10029), .B2(n9632), .A(n9706), .ZN(n10019) );
  NAND2_X1 U11944 ( .A1(n9755), .A2(n9639), .ZN(n10018) );
  NAND2_X1 U11945 ( .A1(n10024), .A2(n16254), .ZN(n15377) );
  NAND2_X1 U11946 ( .A1(n14266), .A2(n10510), .ZN(n10024) );
  NAND2_X1 U11947 ( .A1(n16283), .A2(n11092), .ZN(n15657) );
  INV_X1 U11948 ( .A(n9969), .ZN(n9966) );
  AND2_X1 U11949 ( .A1(n10763), .A2(n9680), .ZN(n13657) );
  INV_X1 U11950 ( .A(n15671), .ZN(n14269) );
  AND2_X1 U11951 ( .A1(n10951), .A2(n10950), .ZN(n16277) );
  AND2_X1 U11952 ( .A1(n14273), .A2(n10955), .ZN(n16275) );
  NAND2_X1 U11953 ( .A1(n10763), .A2(n9988), .ZN(n13649) );
  NAND2_X1 U11954 ( .A1(n19162), .A2(n11091), .ZN(n14174) );
  NAND2_X1 U11955 ( .A1(n10763), .A2(n10762), .ZN(n13588) );
  INV_X1 U11956 ( .A(n19182), .ZN(n10870) );
  AND2_X1 U11957 ( .A1(n13229), .A2(n13228), .ZN(n13231) );
  OR2_X1 U11958 ( .A1(n11088), .A2(n10862), .ZN(n15537) );
  OR2_X1 U11959 ( .A1(n11088), .A2(n16325), .ZN(n19175) );
  INV_X1 U11960 ( .A(n19564), .ZN(n19570) );
  NOR2_X2 U11961 ( .A1(n13863), .A2(n13862), .ZN(n14072) );
  NOR2_X2 U11962 ( .A1(n13861), .A2(n13862), .ZN(n14073) );
  NAND2_X1 U11963 ( .A1(n9655), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9776) );
  NAND2_X1 U11964 ( .A1(n10097), .A2(n16304), .ZN(n9775) );
  INV_X1 U11965 ( .A(n14073), .ZN(n14058) );
  INV_X1 U11966 ( .A(n14072), .ZN(n14057) );
  OR2_X1 U11967 ( .A1(n19076), .A2(n19030), .ZN(n19523) );
  OR2_X1 U11968 ( .A1(n10661), .A2(n10684), .ZN(n16324) );
  NAND2_X1 U11969 ( .A1(n19822), .A2(n13937), .ZN(n19818) );
  CLKBUF_X1 U11970 ( .A(n10662), .Z(n16352) );
  INV_X1 U11971 ( .A(n9731), .ZN(n12989) );
  NOR2_X1 U11972 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16723), .ZN(n16715) );
  AND2_X1 U11973 ( .A1(n9913), .A2(n9911), .ZN(n16712) );
  AND2_X1 U11974 ( .A1(n16721), .A2(n9906), .ZN(n9911) );
  NOR2_X1 U11975 ( .A1(n17662), .A2(n9910), .ZN(n9906) );
  NOR2_X1 U11976 ( .A1(n18595), .A2(n17355), .ZN(n18806) );
  NOR2_X1 U11977 ( .A1(n16896), .A2(n16895), .ZN(n9824) );
  NAND2_X1 U11978 ( .A1(n16996), .A2(P3_EBX_REG_20__SCAN_IN), .ZN(n16981) );
  NOR2_X1 U11979 ( .A1(n17171), .A2(n16780), .ZN(n17122) );
  AOI21_X1 U11980 ( .B1(n15700), .B2(n18654), .A(n18812), .ZN(n17356) );
  INV_X1 U11981 ( .A(n17412), .ZN(n17357) );
  INV_X1 U11982 ( .A(n17355), .ZN(n17414) );
  INV_X1 U11983 ( .A(n13003), .ZN(n12412) );
  AND2_X1 U11984 ( .A1(n13000), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13003) );
  NOR2_X1 U11985 ( .A1(n17504), .A2(n17505), .ZN(n17494) );
  NOR2_X1 U11986 ( .A1(n17507), .A2(n12415), .ZN(n17464) );
  NAND2_X1 U11987 ( .A1(n17605), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n17585) );
  AOI21_X1 U11988 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17548), .A(
        n18539), .ZN(n17661) );
  AND2_X1 U11989 ( .A1(n16721), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n9914) );
  NOR2_X1 U11990 ( .A1(n17746), .A2(n9910), .ZN(n17722) );
  AND2_X1 U11991 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17782) );
  INV_X1 U11992 ( .A(n9921), .ZN(n12975) );
  NOR2_X1 U11993 ( .A1(n17493), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17492) );
  NAND2_X1 U11994 ( .A1(n17573), .A2(n12971), .ZN(n17518) );
  AOI21_X1 U11995 ( .B1(n17615), .B2(n17524), .A(n12969), .ZN(n12970) );
  INV_X1 U11996 ( .A(n17831), .ZN(n17936) );
  AND2_X1 U11997 ( .A1(n16366), .A2(n17965), .ZN(n17647) );
  NAND2_X1 U11998 ( .A1(n17739), .A2(n9926), .ZN(n17698) );
  NOR3_X1 U11999 ( .A1(n9927), .A2(n17730), .A3(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n9926) );
  NOR2_X1 U12000 ( .A1(n13039), .A2(n17727), .ZN(n18016) );
  INV_X1 U12001 ( .A(n16366), .ZN(n18014) );
  NAND3_X1 U12002 ( .A1(n12874), .A2(n12873), .A3(n12872), .ZN(n16409) );
  NOR2_X1 U12003 ( .A1(n17728), .A2(n18055), .ZN(n17727) );
  AOI21_X1 U12004 ( .B1(n17759), .B2(n17760), .A(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n9924) );
  NAND2_X1 U12005 ( .A1(n17752), .A2(n17751), .ZN(n17750) );
  NOR2_X1 U12006 ( .A1(n17759), .A2(n17760), .ZN(n17758) );
  AND2_X1 U12007 ( .A1(n9832), .A2(n9831), .ZN(n15699) );
  NOR2_X1 U12008 ( .A1(n15707), .A2(n18610), .ZN(n9831) );
  NOR2_X1 U12009 ( .A1(n15711), .A2(n15695), .ZN(n16410) );
  XNOR2_X1 U12010 ( .A(n12952), .B(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n17806) );
  XNOR2_X1 U12011 ( .A(n17346), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n17813) );
  AOI21_X1 U12012 ( .B1(n18164), .B2(n12439), .A(n12985), .ZN(n12983) );
  INV_X1 U12013 ( .A(n15811), .ZN(n17821) );
  NAND2_X1 U12014 ( .A1(n14386), .A2(n18158), .ZN(n18262) );
  AOI22_X1 U12015 ( .A1(n18598), .A2(n18594), .B1(n16410), .B2(n18599), .ZN(
        n18603) );
  CLKBUF_X1 U12016 ( .A(n13190), .Z(n13861) );
  INV_X2 U12017 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20752) );
  INV_X1 U12018 ( .A(n19926), .ZN(n19941) );
  INV_X1 U12019 ( .A(n19938), .ZN(n19895) );
  AND2_X1 U12020 ( .A1(n15837), .A2(n13910), .ZN(n19927) );
  INV_X1 U12021 ( .A(n15911), .ZN(n19881) );
  AND2_X1 U12022 ( .A1(n13915), .A2(n13913), .ZN(n19938) );
  INV_X1 U12023 ( .A(n14761), .ZN(n15941) );
  AND2_X2 U12024 ( .A1(n13315), .A2(n14598), .ZN(n15945) );
  INV_X1 U12025 ( .A(n11631), .ZN(n20141) );
  INV_X1 U12026 ( .A(n14828), .ZN(n15949) );
  AND2_X1 U12027 ( .A1(n13418), .A2(n20101), .ZN(n15948) );
  INV_X1 U12028 ( .A(n14815), .ZN(n15946) );
  OR2_X1 U12029 ( .A1(n15947), .A2(n13418), .ZN(n14826) );
  NAND2_X2 U12030 ( .A1(n12394), .A2(n12393), .ZN(n14815) );
  INV_X1 U12031 ( .A(n15949), .ZN(n14814) );
  INV_X1 U12032 ( .A(n14826), .ZN(n14379) );
  CLKBUF_X1 U12033 ( .A(n19968), .Z(n20761) );
  CLKBUF_X1 U12034 ( .A(n19967), .Z(n19962) );
  OAI21_X1 U12035 ( .B1(n14607), .B2(n14609), .A(n14608), .ZN(n14846) );
  INV_X1 U12036 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15845) );
  INV_X1 U12037 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n14900) );
  INV_X1 U12038 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n14927) );
  AND2_X1 U12039 ( .A1(n13391), .A2(n20602), .ZN(n16022) );
  INV_X1 U12040 ( .A(n16026), .ZN(n20091) );
  XNOR2_X1 U12041 ( .A(n14527), .B(n14526), .ZN(n14703) );
  NOR2_X1 U12042 ( .A1(n14418), .A2(n14417), .ZN(n14831) );
  AND2_X1 U12043 ( .A1(n16034), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14993) );
  NAND2_X1 U12044 ( .A1(n16010), .A2(n14144), .ZN(n14394) );
  INV_X1 U12045 ( .A(n16103), .ZN(n16141) );
  NAND2_X1 U12046 ( .A1(n10034), .A2(n14129), .ZN(n16016) );
  NAND2_X1 U12047 ( .A1(n14127), .A2(n14126), .ZN(n10034) );
  NAND2_X1 U12048 ( .A1(n13289), .A2(n13286), .ZN(n16068) );
  INV_X1 U12049 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20519) );
  INV_X1 U12050 ( .A(n11762), .ZN(n11763) );
  INV_X1 U12052 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20738) );
  OR2_X1 U12053 ( .A1(n9620), .A2(n11797), .ZN(n20729) );
  INV_X1 U12054 ( .A(n20602), .ZN(n20728) );
  INV_X1 U12055 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14562) );
  INV_X1 U12056 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16154) );
  NOR2_X1 U12057 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n16151) );
  OAI22_X1 U12058 ( .A1(n20117), .A2(n20116), .B1(n20432), .B2(n20260), .ZN(
        n20145) );
  INV_X1 U12059 ( .A(n20336), .ZN(n20338) );
  NOR2_X1 U12060 ( .A1(n20519), .A2(n20345), .ZN(n20365) );
  OAI211_X1 U12061 ( .C1(n20394), .C2(n20493), .A(n20430), .B(n20378), .ZN(
        n20396) );
  AND2_X1 U12062 ( .A1(n20457), .A2(n20546), .ZN(n20483) );
  OAI211_X1 U12063 ( .C1(n20587), .C2(n20557), .A(n20556), .B(n20555), .ZN(
        n20590) );
  NOR2_X1 U12064 ( .A1(n20519), .A2(n20604), .ZN(n20648) );
  INV_X1 U12065 ( .A(n20107), .ZN(n20653) );
  NAND2_X1 U12066 ( .A1(n13902), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20660) );
  INV_X1 U12067 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20493) );
  AOI221_X1 U12068 ( .B1(n20756), .B2(n13902), .C1(n15766), .C2(n13902), .A(
        n16158), .ZN(n16162) );
  NAND2_X1 U12069 ( .A1(n16165), .A2(n9736), .ZN(n11286) );
  AND2_X1 U12070 ( .A1(n9838), .A2(n9737), .ZN(n9736) );
  AND2_X1 U12071 ( .A1(n16166), .A2(n18993), .ZN(n9737) );
  INV_X1 U12072 ( .A(n9837), .ZN(n11248) );
  NOR2_X1 U12073 ( .A1(n11247), .A2(n16206), .ZN(n15085) );
  NAND2_X1 U12074 ( .A1(n15287), .A2(n11219), .ZN(n9860) );
  INV_X1 U12075 ( .A(n18876), .ZN(n9738) );
  NOR2_X1 U12076 ( .A1(n18876), .A2(n11247), .ZN(n18865) );
  NOR2_X1 U12077 ( .A1(n18865), .A2(n18866), .ZN(n18864) );
  OAI21_X1 U12078 ( .B1(n18896), .B2(n18898), .A(n11225), .ZN(n18890) );
  NOR2_X1 U12079 ( .A1(n18954), .A2(n18956), .ZN(n18947) );
  INV_X1 U12080 ( .A(n18978), .ZN(n19017) );
  INV_X1 U12081 ( .A(n19028), .ZN(n18997) );
  INV_X1 U12082 ( .A(n18984), .ZN(n19022) );
  NOR2_X1 U12083 ( .A1(n13524), .A2(n10909), .ZN(n13769) );
  OR2_X1 U12084 ( .A1(n11258), .A2(n11266), .ZN(n19004) );
  INV_X1 U12085 ( .A(n19004), .ZN(n19020) );
  OR2_X1 U12086 ( .A1(n10993), .A2(n10992), .ZN(n13813) );
  INV_X1 U12087 ( .A(n15124), .ZN(n15150) );
  XNOR2_X1 U12088 ( .A(n13510), .B(n13511), .ZN(n19076) );
  INV_X1 U12089 ( .A(n19787), .ZN(n14180) );
  NAND2_X2 U12090 ( .A1(n13499), .A2(n19673), .ZN(n15169) );
  NAND2_X1 U12091 ( .A1(n19069), .A2(n12849), .ZN(n15206) );
  AND2_X1 U12092 ( .A1(n13301), .A2(n13863), .ZN(n19039) );
  NAND2_X1 U12093 ( .A1(n12846), .A2(n12845), .ZN(n19069) );
  NAND2_X1 U12094 ( .A1(n12843), .A2(n19673), .ZN(n12846) );
  NAND2_X1 U12095 ( .A1(n12526), .A2(n12525), .ZN(n13596) );
  AND2_X1 U12096 ( .A1(n19046), .A2(n19103), .ZN(n19082) );
  OR2_X1 U12097 ( .A1(n19037), .A2(n13301), .ZN(n19071) );
  NAND2_X1 U12098 ( .A1(n19069), .A2(n12847), .ZN(n19103) );
  AND2_X1 U12099 ( .A1(n13112), .A2(n19829), .ZN(n13211) );
  INV_X1 U12100 ( .A(n13211), .ZN(n13225) );
  XNOR2_X1 U12101 ( .A(n11250), .B(n11151), .ZN(n16172) );
  INV_X1 U12102 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16245) );
  INV_X1 U12103 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n16274) );
  INV_X1 U12104 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13690) );
  NAND2_X1 U12105 ( .A1(n13110), .A2(n11121), .ZN(n19154) );
  INV_X1 U12106 ( .A(n19141), .ZN(n15396) );
  INV_X1 U12107 ( .A(n11114), .ZN(n19147) );
  NOR2_X1 U12108 ( .A1(n9787), .A2(n9786), .ZN(n11173) );
  NOR3_X1 U12109 ( .A1(n12480), .A2(n11168), .A3(n9788), .ZN(n9787) );
  OAI21_X1 U12110 ( .B1(n15172), .B2(n19185), .A(n11169), .ZN(n9786) );
  NAND2_X1 U12111 ( .A1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n9789), .ZN(
        n9788) );
  INV_X1 U12112 ( .A(n11098), .ZN(n11099) );
  INV_X1 U12113 ( .A(n9769), .ZN(n12460) );
  NAND2_X1 U12114 ( .A1(n14200), .A2(n14199), .ZN(n15553) );
  NAND2_X1 U12115 ( .A1(n10021), .A2(n10025), .ZN(n15637) );
  NAND2_X1 U12116 ( .A1(n10023), .A2(n10022), .ZN(n10021) );
  AND2_X1 U12117 ( .A1(n14273), .A2(n9679), .ZN(n15629) );
  NOR2_X1 U12118 ( .A1(n10526), .A2(n15657), .ZN(n15647) );
  NAND2_X1 U12119 ( .A1(n14273), .A2(n10006), .ZN(n15642) );
  NOR2_X1 U12120 ( .A1(n14174), .A2(n14173), .ZN(n16283) );
  NAND2_X1 U12121 ( .A1(n9965), .A2(n10724), .ZN(n14169) );
  NAND2_X1 U12122 ( .A1(n10725), .A2(n10723), .ZN(n9965) );
  NOR2_X1 U12123 ( .A1(n16298), .A2(n16299), .ZN(n19162) );
  INV_X1 U12124 ( .A(n19185), .ZN(n16296) );
  OR2_X1 U12125 ( .A1(n11088), .A2(n10844), .ZN(n19179) );
  OR2_X1 U12126 ( .A1(n11088), .A2(n11087), .ZN(n19185) );
  OR2_X1 U12127 ( .A1(n13299), .A2(n13298), .ZN(n19796) );
  INV_X1 U12128 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19793) );
  NAND2_X1 U12129 ( .A1(n13529), .A2(n13528), .ZN(n19787) );
  OR2_X1 U12130 ( .A1(n13527), .A2(n13526), .ZN(n13528) );
  AND2_X1 U12131 ( .A1(n13521), .A2(n13520), .ZN(n19782) );
  AND2_X1 U12132 ( .A1(n13166), .A2(n13165), .ZN(n13975) );
  OR3_X1 U12133 ( .A1(n19196), .A2(n19565), .A3(n19195), .ZN(n19219) );
  NOR2_X1 U12134 ( .A1(n19193), .A2(n19312), .ZN(n19241) );
  OR3_X1 U12135 ( .A1(n19386), .A2(n19565), .A3(n19385), .ZN(n19404) );
  AND2_X1 U12136 ( .A1(n19274), .A2(n14037), .ZN(n19444) );
  INV_X1 U12137 ( .A(n19444), .ZN(n19458) );
  INV_X1 U12138 ( .A(n19580), .ZN(n19606) );
  INV_X1 U12139 ( .A(n19552), .ZN(n19595) );
  OAI21_X1 U12140 ( .B1(n14104), .B2(n14108), .A(n14103), .ZN(n19631) );
  INV_X1 U12141 ( .A(n19216), .ZN(n19627) );
  INV_X1 U12142 ( .A(n19283), .ZN(n19574) );
  INV_X1 U12143 ( .A(n19540), .ZN(n19639) );
  INV_X1 U12144 ( .A(n19543), .ZN(n19646) );
  INV_X1 U12145 ( .A(n19586), .ZN(n19645) );
  INV_X1 U12146 ( .A(n19289), .ZN(n19644) );
  INV_X1 U12147 ( .A(n19546), .ZN(n19652) );
  INV_X1 U12148 ( .A(n19589), .ZN(n19651) );
  INV_X1 U12149 ( .A(n19207), .ZN(n19649) );
  INV_X1 U12150 ( .A(n19295), .ZN(n19656) );
  INV_X1 U12151 ( .A(n19298), .ZN(n19594) );
  INV_X1 U12152 ( .A(n19516), .ZN(n19666) );
  INV_X1 U12153 ( .A(n19603), .ZN(n19668) );
  INV_X1 U12154 ( .A(n14189), .ZN(n19663) );
  NOR2_X2 U12155 ( .A1(n19488), .A2(n14047), .ZN(n19669) );
  NOR2_X1 U12156 ( .A1(n14045), .A2(n14044), .ZN(n19665) );
  INV_X1 U12157 ( .A(n19673), .ZN(n16361) );
  AND2_X1 U12158 ( .A1(n16328), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16356) );
  INV_X2 U12159 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19794) );
  NAND2_X1 U12160 ( .A1(n16805), .A2(n9664), .ZN(n16668) );
  INV_X1 U12161 ( .A(n16668), .ZN(n16655) );
  NOR2_X1 U12162 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16680), .ZN(n16664) );
  NOR2_X1 U12163 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16820), .ZN(n16806) );
  NOR2_X2 U12164 ( .A1(n18653), .A2(n12452), .ZN(n16843) );
  INV_X1 U12165 ( .A(n16843), .ZN(n16879) );
  NAND4_X1 U12166 ( .A1(n18141), .A2(n18827), .A3(n18667), .A4(n18658), .ZN(
        n16891) );
  NAND2_X1 U12167 ( .A1(n16954), .A2(n9823), .ZN(n16942) );
  AND2_X1 U12168 ( .A1(n9650), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n9823) );
  NOR2_X1 U12169 ( .A1(n16894), .A2(n16970), .ZN(n16954) );
  NAND2_X1 U12170 ( .A1(n17039), .A2(n10054), .ZN(n17009) );
  NOR2_X1 U12171 ( .A1(n17063), .A2(n16703), .ZN(n17039) );
  NAND2_X1 U12172 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17067), .ZN(n17063) );
  NOR2_X1 U12173 ( .A1(n16724), .A2(n17104), .ZN(n17067) );
  NAND2_X1 U12174 ( .A1(n17117), .A2(P3_EBX_REG_12__SCAN_IN), .ZN(n17104) );
  NAND2_X1 U12175 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17122), .ZN(n17118) );
  NOR2_X1 U12176 ( .A1(n17118), .A2(n17119), .ZN(n17117) );
  NAND2_X1 U12177 ( .A1(n17187), .A2(n9825), .ZN(n17171) );
  NOR2_X1 U12178 ( .A1(n9827), .A2(n9828), .ZN(n9825) );
  NAND2_X1 U12179 ( .A1(n17187), .A2(P3_EBX_REG_5__SCAN_IN), .ZN(n17178) );
  NOR2_X1 U12180 ( .A1(n11397), .A2(n11396), .ZN(n17184) );
  AND2_X1 U12181 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n17184), .ZN(n17187) );
  INV_X1 U12182 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17190) );
  INV_X2 U12183 ( .A(n17203), .ZN(n17197) );
  INV_X1 U12184 ( .A(n11397), .ZN(n17206) );
  NOR2_X1 U12185 ( .A1(n17362), .A2(n17227), .ZN(n17223) );
  NAND2_X1 U12186 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17231), .ZN(n17227) );
  NAND2_X1 U12187 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(P3_EAX_REG_25__SCAN_IN), 
        .ZN(n9727) );
  NOR3_X1 U12188 ( .A1(n17245), .A2(n17292), .A3(n9728), .ZN(n17236) );
  NOR2_X1 U12189 ( .A1(n17379), .A2(n17277), .ZN(n17271) );
  INV_X1 U12190 ( .A(n17287), .ZN(n17276) );
  NAND2_X1 U12191 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17288), .ZN(n17284) );
  NAND4_X1 U12192 ( .A1(n17316), .A2(P3_EAX_REG_14__SCAN_IN), .A3(
        P3_EAX_REG_13__SCAN_IN), .A4(n17209), .ZN(n17294) );
  NAND2_X1 U12193 ( .A1(n9726), .A2(n9724), .ZN(n17321) );
  NOR2_X1 U12194 ( .A1(n17208), .A2(n9725), .ZN(n9724) );
  INV_X1 U12195 ( .A(n17350), .ZN(n9726) );
  NOR2_X1 U12196 ( .A1(n12935), .A2(n12934), .ZN(n17326) );
  INV_X1 U12197 ( .A(n13010), .ZN(n17329) );
  NOR2_X1 U12198 ( .A1(n12925), .A2(n12924), .ZN(n17333) );
  INV_X1 U12199 ( .A(n13013), .ZN(n17336) );
  NOR2_X1 U12200 ( .A1(n12915), .A2(n12914), .ZN(n17341) );
  INV_X1 U12201 ( .A(n17348), .ZN(n17345) );
  INV_X1 U12202 ( .A(n9829), .ZN(n15808) );
  NOR2_X1 U12203 ( .A1(n18630), .A2(n17340), .ZN(n17348) );
  INV_X1 U12204 ( .A(n17342), .ZN(n17347) );
  CLKBUF_X1 U12206 ( .A(n17459), .Z(n17453) );
  INV_X1 U12207 ( .A(n17462), .ZN(n17454) );
  OAI211_X1 U12208 ( .C1(n18815), .C2(n18164), .A(n17415), .B(n17414), .ZN(
        n17459) );
  NOR2_X1 U12209 ( .A1(n17453), .A2(n18164), .ZN(n17460) );
  INV_X1 U12210 ( .A(n13000), .ZN(n16378) );
  AND2_X1 U12211 ( .A1(n17605), .A2(n9695), .ZN(n17534) );
  INV_X1 U12212 ( .A(n17734), .ZN(n17690) );
  NAND2_X1 U12213 ( .A1(n17749), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n17746) );
  NOR2_X1 U12214 ( .A1(n17766), .A2(n17765), .ZN(n17749) );
  INV_X2 U12215 ( .A(n18264), .ZN(n18539) );
  NAND2_X1 U12216 ( .A1(n17782), .A2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n17766) );
  INV_X1 U12217 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17765) );
  INV_X1 U12218 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17793) );
  INV_X1 U12219 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17811) );
  NAND2_X1 U12220 ( .A1(n12978), .A2(n12981), .ZN(n9920) );
  NAND2_X1 U12221 ( .A1(n9919), .A2(n9663), .ZN(n9918) );
  NOR2_X1 U12222 ( .A1(n18016), .A2(n17831), .ZN(n17971) );
  INV_X1 U12223 ( .A(n18062), .ZN(n17987) );
  NOR3_X1 U12224 ( .A1(n9928), .A2(n17730), .A3(n9927), .ZN(n17710) );
  NAND2_X1 U12225 ( .A1(n17739), .A2(n9929), .ZN(n13007) );
  AOI21_X2 U12226 ( .B1(n15716), .B2(n15715), .A(n18811), .ZN(n18125) );
  NAND2_X1 U12227 ( .A1(n18826), .A2(n15699), .ZN(n18108) );
  NOR2_X1 U12228 ( .A1(n18135), .A2(n18125), .ZN(n18121) );
  INV_X1 U12229 ( .A(n18121), .ZN(n18126) );
  NOR2_X1 U12230 ( .A1(n17995), .A2(n18142), .ZN(n18138) );
  NOR2_X1 U12231 ( .A1(n18600), .A2(n18142), .ZN(n18140) );
  INV_X1 U12232 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18641) );
  INV_X1 U12233 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20792) );
  INV_X1 U12234 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18768) );
  AOI211_X1 U12235 ( .C1(n18652), .C2(n18628), .A(n18159), .B(n15703), .ZN(
        n18794) );
  INV_X1 U12236 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18604) );
  INV_X1 U12237 ( .A(n18794), .ZN(n18791) );
  INV_X1 U12238 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18763) );
  NAND2_X1 U12239 ( .A1(n18688), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18823) );
  AND2_X1 U12240 ( .A1(n12404), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n20099)
         );
  NAND2_X1 U12242 ( .A1(n9822), .A2(n9820), .ZN(n9819) );
  INV_X1 U12243 ( .A(n9821), .ZN(n9820) );
  AND2_X1 U12244 ( .A1(n16175), .A2(n16176), .ZN(n9833) );
  OR4_X1 U12245 ( .A1(n13079), .A2(n13078), .A3(n13077), .A4(n13076), .ZN(
        P2_U2828) );
  NAND2_X1 U12246 ( .A1(n12494), .A2(n16261), .ZN(n12495) );
  OAI21_X1 U12247 ( .B1(n15435), .B2(n19157), .A(n9668), .ZN(P2_U3020) );
  OR3_X1 U12248 ( .A1(n16539), .A2(n16538), .A3(n16689), .ZN(n10073) );
  AOI211_X1 U12249 ( .C1(n16543), .C2(n16865), .A(n16542), .B(n16541), .ZN(
        n16546) );
  OAI21_X1 U12250 ( .B1(n11474), .B2(P3_EBX_REG_28__SCAN_IN), .A(n11473), .ZN(
        n11475) );
  AOI21_X1 U12251 ( .B1(n9733), .B2(P3_EAX_REG_31__SCAN_IN), .A(n9685), .ZN(
        n17212) );
  NAND2_X1 U12252 ( .A1(n9735), .A2(n9734), .ZN(n9733) );
  NAND2_X1 U12253 ( .A1(n9917), .A2(n9915), .ZN(P3_U2831) );
  AOI21_X1 U12254 ( .B1(n16400), .B2(n17987), .A(n9916), .ZN(n9915) );
  NAND2_X1 U12255 ( .A1(n16399), .A2(n18058), .ZN(n9917) );
  OAI21_X1 U12256 ( .B1(n16402), .B2(n18090), .A(n16401), .ZN(n9916) );
  AND2_X1 U12257 ( .A1(n10025), .A2(n10020), .ZN(n9632) );
  AND2_X1 U12258 ( .A1(n12536), .A2(n9644), .ZN(n9633) );
  INV_X1 U12259 ( .A(n11306), .ZN(n11441) );
  NAND2_X1 U12260 ( .A1(n13964), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10128) );
  AND2_X1 U12261 ( .A1(n12962), .A2(n12961), .ZN(n9634) );
  NAND2_X1 U12262 ( .A1(n9968), .A2(n9967), .ZN(n15335) );
  INV_X1 U12263 ( .A(n10173), .ZN(n19829) );
  INV_X2 U12264 ( .A(n11085), .ZN(n12780) );
  NOR2_X1 U12265 ( .A1(n11296), .A2(n18618), .ZN(n16916) );
  INV_X1 U12266 ( .A(n13249), .ZN(n20103) );
  NAND2_X1 U12267 ( .A1(n9854), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n9635) );
  AND2_X1 U12268 ( .A1(n10048), .A2(n9626), .ZN(n9636) );
  OR2_X1 U12269 ( .A1(n15549), .A2(n10583), .ZN(n9637) );
  NAND2_X1 U12270 ( .A1(n12536), .A2(n9847), .ZN(n9638) );
  AND2_X1 U12271 ( .A1(n9759), .A2(n9632), .ZN(n9639) );
  INV_X1 U12272 ( .A(n10507), .ZN(n9879) );
  INV_X1 U12273 ( .A(n10029), .ZN(n10022) );
  NAND2_X1 U12274 ( .A1(n10030), .A2(n16254), .ZN(n10029) );
  AND2_X1 U12275 ( .A1(n10039), .A2(n10043), .ZN(n9640) );
  AND2_X1 U12276 ( .A1(n9967), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9641) );
  AND2_X1 U12277 ( .A1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n11124), .ZN(
        n9642) );
  AND2_X1 U12278 ( .A1(n9680), .A2(n13656), .ZN(n9643) );
  NAND2_X1 U12279 ( .A1(n9841), .A2(n13593), .ZN(n13500) );
  INV_X1 U12280 ( .A(n13524), .ZN(n10002) );
  NAND2_X1 U12281 ( .A1(n12536), .A2(n12535), .ZN(n13930) );
  AND2_X1 U12282 ( .A1(n12535), .A2(n9848), .ZN(n9644) );
  AND2_X1 U12283 ( .A1(n9678), .A2(n14226), .ZN(n9645) );
  AND2_X1 U12284 ( .A1(n9892), .A2(n14740), .ZN(n9646) );
  INV_X1 U12285 ( .A(n11822), .ZN(n9947) );
  AND2_X1 U12286 ( .A1(n9946), .A2(n9745), .ZN(n9647) );
  AND2_X1 U12287 ( .A1(n9901), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9648) );
  AND2_X1 U12288 ( .A1(n9889), .A2(n9887), .ZN(n9649) );
  INV_X1 U12289 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n9910) );
  NAND2_X1 U12290 ( .A1(n9913), .A2(n9914), .ZN(n16736) );
  AND2_X1 U12291 ( .A1(n9824), .A2(P3_EBX_REG_25__SCAN_IN), .ZN(n9650) );
  OR2_X1 U12292 ( .A1(n11291), .A2(n18618), .ZN(n9651) );
  INV_X1 U12293 ( .A(n9732), .ZN(n18164) );
  OR2_X1 U12294 ( .A1(n11395), .A2(n11394), .ZN(n9732) );
  AND2_X1 U12295 ( .A1(n9968), .A2(n9966), .ZN(n15344) );
  OR2_X1 U12296 ( .A1(n14242), .A2(n14308), .ZN(n9653) );
  NAND2_X1 U12297 ( .A1(n15392), .A2(n10737), .ZN(n9968) );
  AND2_X1 U12298 ( .A1(n10537), .A2(n9873), .ZN(n10562) );
  NAND2_X1 U12299 ( .A1(n11119), .A2(n9986), .ZN(n13056) );
  OR3_X1 U12301 ( .A1(n17245), .A2(n17292), .A3(n9727), .ZN(n9654) );
  NOR2_X1 U12302 ( .A1(n14709), .A2(n12181), .ZN(n14662) );
  AND4_X1 U12303 ( .A1(n10096), .A2(n10095), .A3(n10094), .A4(n10093), .ZN(
        n9655) );
  OR2_X1 U12305 ( .A1(n14406), .A2(n14405), .ZN(n9657) );
  OR2_X2 U12306 ( .A1(n11557), .A2(n11556), .ZN(n11631) );
  AND2_X1 U12307 ( .A1(n9873), .A2(n10542), .ZN(n9658) );
  AND2_X1 U12308 ( .A1(n15075), .A2(n15076), .ZN(n15074) );
  NAND2_X1 U12309 ( .A1(n10422), .A2(n10421), .ZN(n10727) );
  INV_X1 U12310 ( .A(n10727), .ZN(n10423) );
  AND4_X1 U12311 ( .A1(n11650), .A2(n11649), .A3(n13280), .A4(n11648), .ZN(
        n9659) );
  NOR2_X1 U12312 ( .A1(n13716), .A2(n15018), .ZN(n9660) );
  NOR2_X1 U12313 ( .A1(n15436), .A2(n9881), .ZN(n9661) );
  OR2_X1 U12314 ( .A1(n10362), .A2(n10279), .ZN(n9662) );
  OR2_X1 U12315 ( .A1(n15776), .A2(n15782), .ZN(n9663) );
  NOR2_X1 U12316 ( .A1(n10651), .A2(n10650), .ZN(n10682) );
  NAND2_X1 U12317 ( .A1(n16653), .A2(n16693), .ZN(n9664) );
  AND2_X1 U12318 ( .A1(n11847), .A2(n11871), .ZN(n9665) );
  AND2_X1 U12319 ( .A1(n19019), .A2(n10256), .ZN(n10276) );
  AND3_X1 U12320 ( .A1(n11644), .A2(n13273), .A3(n11640), .ZN(n9666) );
  NAND3_X1 U12321 ( .A1(n11571), .A2(n11572), .A3(n11570), .ZN(n9667) );
  AND2_X1 U12322 ( .A1(n9882), .A2(n9661), .ZN(n9668) );
  AND2_X1 U12323 ( .A1(n9968), .A2(n9641), .ZN(n15322) );
  AND2_X1 U12324 ( .A1(n9755), .A2(n9759), .ZN(n14266) );
  NAND2_X1 U12325 ( .A1(n10537), .A2(n10536), .ZN(n10541) );
  AND2_X1 U12326 ( .A1(n10334), .A2(n9721), .ZN(n10475) );
  NAND2_X1 U12327 ( .A1(n10448), .A2(n13295), .ZN(n10668) );
  INV_X1 U12328 ( .A(n10668), .ZN(n9723) );
  AND2_X1 U12329 ( .A1(n10457), .A2(n10456), .ZN(n9669) );
  INV_X1 U12330 ( .A(n12519), .ZN(n10286) );
  OR2_X1 U12331 ( .A1(n16985), .A2(n12903), .ZN(n9670) );
  INV_X1 U12332 ( .A(n10042), .ZN(n10041) );
  NAND2_X1 U12333 ( .A1(n11679), .A2(n10045), .ZN(n10042) );
  AND2_X1 U12334 ( .A1(n9640), .A2(n9660), .ZN(n9671) );
  NAND2_X1 U12335 ( .A1(n12459), .A2(n15417), .ZN(n9672) );
  OR2_X1 U12336 ( .A1(n14134), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16014) );
  AND2_X2 U12337 ( .A1(n10258), .A2(n10252), .ZN(n19019) );
  NAND2_X1 U12338 ( .A1(n10173), .A2(n19794), .ZN(n10891) );
  INV_X1 U12339 ( .A(n11039), .ZN(n10888) );
  INV_X1 U12341 ( .A(n11617), .ZN(n13259) );
  NAND2_X1 U12342 ( .A1(n17605), .A2(n9648), .ZN(n12410) );
  AND3_X1 U12343 ( .A1(n11123), .A2(n9642), .A3(n11234), .ZN(n11230) );
  AND2_X1 U12344 ( .A1(n16954), .A2(n9650), .ZN(n9673) );
  AND2_X1 U12345 ( .A1(n16954), .A2(n9824), .ZN(n9674) );
  AND2_X1 U12346 ( .A1(n16954), .A2(P3_EBX_REG_23__SCAN_IN), .ZN(n9675) );
  NOR2_X1 U12348 ( .A1(n11228), .A2(n16245), .ZN(n11226) );
  NAND2_X1 U12350 ( .A1(n15458), .A2(n15079), .ZN(n15078) );
  OR2_X1 U12351 ( .A1(n17676), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9676) );
  AND2_X1 U12352 ( .A1(n17605), .A2(n9901), .ZN(n9677) );
  NOR2_X1 U12353 ( .A1(n9653), .A2(n11118), .ZN(n11119) );
  AND2_X1 U12354 ( .A1(n11119), .A2(n9983), .ZN(n15075) );
  NAND2_X1 U12355 ( .A1(n14031), .A2(n14030), .ZN(n14032) );
  NAND2_X1 U12356 ( .A1(n17292), .A2(n12433), .ZN(n12991) );
  INV_X1 U12357 ( .A(n12991), .ZN(n9832) );
  AND2_X1 U12358 ( .A1(n10004), .A2(n14199), .ZN(n9678) );
  AND2_X1 U12359 ( .A1(n10006), .A2(n10005), .ZN(n9679) );
  AND2_X1 U12360 ( .A1(n9988), .A2(n9987), .ZN(n9680) );
  NOR3_X1 U12361 ( .A1(n18160), .A2(n18164), .A3(n18811), .ZN(n9681) );
  INV_X1 U12362 ( .A(n17730), .ZN(n17656) );
  NAND2_X1 U12364 ( .A1(n14255), .A2(n14254), .ZN(n13086) );
  AND2_X1 U12365 ( .A1(n11189), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9682) );
  INV_X1 U12366 ( .A(n11797), .ZN(n20258) );
  NAND2_X1 U12367 ( .A1(n11796), .A2(n11795), .ZN(n11797) );
  AND2_X1 U12368 ( .A1(n9679), .A2(n15628), .ZN(n9683) );
  AND2_X1 U12369 ( .A1(n9981), .A2(n9980), .ZN(n9684) );
  AND2_X1 U12370 ( .A1(n17283), .A2(BUF2_REG_31__SCAN_IN), .ZN(n9685) );
  INV_X1 U12371 ( .A(n13581), .ZN(n13580) );
  NAND2_X1 U12372 ( .A1(n14031), .A2(n9978), .ZN(n14088) );
  OR2_X1 U12373 ( .A1(n14735), .A2(n14728), .ZN(n9686) );
  INV_X1 U12374 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n15382) );
  OR2_X1 U12375 ( .A1(n13639), .A2(n13725), .ZN(n9687) );
  NOR2_X1 U12376 ( .A1(n9626), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9688) );
  AND2_X1 U12377 ( .A1(n13760), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9689) );
  AND2_X1 U12378 ( .A1(n9895), .A2(n9894), .ZN(n9690) );
  AND2_X1 U12379 ( .A1(n9839), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n9691)
         );
  AND2_X1 U12380 ( .A1(n9951), .A2(n14738), .ZN(n9692) );
  AND2_X1 U12381 ( .A1(n9978), .A2(n9977), .ZN(n9693) );
  AND2_X1 U12382 ( .A1(n9645), .A2(n10003), .ZN(n9694) );
  AND2_X1 U12383 ( .A1(n9648), .A2(n17545), .ZN(n9695) );
  AND2_X1 U12384 ( .A1(n11895), .A2(n9945), .ZN(n9696) );
  AND2_X1 U12385 ( .A1(n9646), .A2(n9891), .ZN(n9697) );
  INV_X1 U12386 ( .A(n9886), .ZN(n9885) );
  NOR2_X1 U12387 ( .A1(n13581), .A2(n13644), .ZN(n9886) );
  NOR2_X1 U12388 ( .A1(n11212), .A2(n11211), .ZN(n9698) );
  INV_X1 U12389 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n9903) );
  INV_X1 U12390 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n9902) );
  AND2_X1 U12391 ( .A1(n9841), .A2(n9839), .ZN(n13502) );
  INV_X1 U12392 ( .A(n14753), .ZN(n9955) );
  NAND2_X1 U12393 ( .A1(n11617), .A2(n14596), .ZN(n13095) );
  NOR2_X1 U12394 ( .A1(n11221), .A2(n15309), .ZN(n11125) );
  AND2_X1 U12395 ( .A1(n11190), .A2(n11189), .ZN(n11213) );
  NAND2_X1 U12396 ( .A1(n13797), .A2(n13796), .ZN(n13986) );
  INV_X1 U12397 ( .A(n13986), .ZN(n9888) );
  OR2_X1 U12398 ( .A1(n12718), .A2(n12717), .ZN(n9699) );
  INV_X2 U12399 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n20756) );
  INV_X1 U12400 ( .A(n14029), .ZN(n9848) );
  AND2_X1 U12401 ( .A1(n9997), .A2(n14254), .ZN(n9700) );
  AND2_X1 U12402 ( .A1(n10009), .A2(n15079), .ZN(n9701) );
  AND2_X1 U12403 ( .A1(n9701), .A2(n10008), .ZN(n9702) );
  AND2_X1 U12404 ( .A1(n11190), .A2(n9682), .ZN(n11210) );
  INV_X1 U12405 ( .A(n17739), .ZN(n9928) );
  INV_X1 U12406 ( .A(n13057), .ZN(n9985) );
  INV_X1 U12407 ( .A(n12778), .ZN(n9856) );
  AND2_X1 U12408 ( .A1(n9986), .A2(n9985), .ZN(n9703) );
  AND2_X1 U12409 ( .A1(n14756), .A2(n9892), .ZN(n9704) );
  NAND2_X1 U12410 ( .A1(n13466), .A2(n13397), .ZN(n9800) );
  AND2_X1 U12411 ( .A1(n17207), .A2(n17292), .ZN(n17317) );
  INV_X2 U12412 ( .A(n17317), .ZN(n17340) );
  AND2_X2 U12413 ( .A1(n12686), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12626) );
  AND2_X1 U12414 ( .A1(n10002), .A2(n10001), .ZN(n9705) );
  AND2_X1 U12415 ( .A1(n10535), .A2(n10534), .ZN(n9706) );
  NAND2_X1 U12416 ( .A1(n17730), .A2(n17834), .ZN(n9707) );
  INV_X1 U12417 ( .A(n9827), .ZN(n9826) );
  AND2_X1 U12418 ( .A1(n9998), .A2(n13768), .ZN(n9708) );
  INV_X1 U12419 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n9789) );
  NAND2_X1 U12420 ( .A1(n11152), .A2(n11251), .ZN(n9709) );
  INV_X1 U12421 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18055) );
  INV_X1 U12422 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17816) );
  AND2_X1 U12423 ( .A1(n13252), .A2(n13251), .ZN(n13466) );
  AND2_X1 U12424 ( .A1(n9700), .A2(n9996), .ZN(n9710) );
  AND2_X1 U12425 ( .A1(n9702), .A2(n10007), .ZN(n9711) );
  INV_X1 U12426 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n9877) );
  INV_X1 U12427 ( .A(n14757), .ZN(n9893) );
  INV_X1 U12428 ( .A(n13818), .ZN(n9982) );
  AND2_X1 U12430 ( .A1(n17187), .A2(n9826), .ZN(n9712) );
  AND2_X1 U12431 ( .A1(n12776), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n13593) );
  INV_X1 U12432 ( .A(n13593), .ZN(n9840) );
  NAND2_X1 U12433 ( .A1(n15345), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9713) );
  INV_X1 U12434 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11477) );
  INV_X1 U12435 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n9935) );
  INV_X1 U12436 ( .A(n17746), .ZN(n9913) );
  INV_X1 U12437 ( .A(n17662), .ZN(n9912) );
  AND2_X1 U12438 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n9714) );
  AND2_X1 U12439 ( .A1(n14528), .A2(n16065), .ZN(n9715) );
  INV_X1 U12440 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n9855) );
  INV_X1 U12441 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n9853) );
  INV_X1 U12442 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n9728) );
  INV_X1 U12443 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n9872) );
  CLKBUF_X1 U12444 ( .A(n18413), .Z(n9716) );
  NOR3_X1 U12445 ( .A1(n18634), .A2(n18330), .A3(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18413) );
  OAI221_X1 U12446 ( .B1(n20283), .B2(n20493), .C1(n20283), .C2(n20267), .A(
        n20556), .ZN(n20285) );
  NOR2_X2 U12447 ( .A1(n20142), .A2(n11630), .ZN(n20636) );
  AOI22_X2 U12448 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20140), .B1(DATAI_26_), 
        .B2(n20100), .ZN(n20623) );
  NOR2_X2 U12449 ( .A1(n20102), .A2(n20101), .ZN(n20140) );
  NOR2_X2 U12450 ( .A1(n20142), .A2(n11635), .ZN(n20618) );
  NOR2_X2 U12451 ( .A1(n12848), .A2(n14068), .ZN(n19593) );
  NAND2_X1 U12452 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19533), .ZN(n14068) );
  AND3_X4 U12453 ( .A1(n10080), .A2(n9717), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10293) );
  NOR2_X2 U12454 ( .A1(n15235), .A2(n11168), .ZN(n15216) );
  INV_X1 U12455 ( .A(n9971), .ZN(n9719) );
  NAND2_X2 U12456 ( .A1(n9749), .A2(n10390), .ZN(n10477) );
  NAND3_X1 U12457 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(P3_EAX_REG_0__SCAN_IN), 
        .A3(P3_EAX_REG_7__SCAN_IN), .ZN(n9725) );
  NOR2_X1 U12458 ( .A1(n17245), .A2(n17292), .ZN(n17241) );
  INV_X1 U12459 ( .A(n17236), .ZN(n17240) );
  INV_X2 U12460 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18786) );
  NAND4_X1 U12462 ( .A1(n11570), .A2(n11572), .A3(n11571), .A4(n13279), .ZN(
        n13094) );
  NAND3_X1 U12463 ( .A1(n9752), .A2(n9750), .A3(n10377), .ZN(n9749) );
  NOR2_X1 U12464 ( .A1(n9751), .A2(n10370), .ZN(n9750) );
  NAND2_X1 U12465 ( .A1(n10375), .A2(n10376), .ZN(n9751) );
  NAND3_X1 U12466 ( .A1(n10367), .A2(n10365), .A3(n10366), .ZN(n9753) );
  NAND2_X1 U12467 ( .A1(n10202), .A2(n10201), .ZN(n10203) );
  NAND2_X1 U12468 ( .A1(n10189), .A2(n10188), .ZN(n10204) );
  NAND2_X2 U12469 ( .A1(n10253), .A2(n10252), .ZN(n10251) );
  NAND2_X1 U12470 ( .A1(n10467), .A2(n13760), .ZN(n9761) );
  NAND2_X1 U12471 ( .A1(n10467), .A2(n9689), .ZN(n9756) );
  NAND2_X1 U12472 ( .A1(n9758), .A2(n14173), .ZN(n9757) );
  INV_X1 U12473 ( .A(n13760), .ZN(n9758) );
  NAND2_X1 U12474 ( .A1(n9761), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9759) );
  NAND2_X1 U12475 ( .A1(n10472), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9760) );
  NOR2_X1 U12476 ( .A1(n10746), .A2(n9766), .ZN(n9762) );
  NAND2_X2 U12477 ( .A1(n10238), .A2(n9762), .ZN(n9763) );
  NAND3_X2 U12478 ( .A1(n9764), .A2(n9765), .A3(n9763), .ZN(n12498) );
  NAND4_X1 U12479 ( .A1(n9764), .A2(n9765), .A3(n9763), .A4(n10247), .ZN(
        n10285) );
  OR2_X2 U12480 ( .A1(n10238), .A2(n9767), .ZN(n9764) );
  NAND2_X1 U12481 ( .A1(n10238), .A2(n10237), .ZN(n10747) );
  NAND2_X1 U12482 ( .A1(n10746), .A2(n9766), .ZN(n9765) );
  INV_X1 U12483 ( .A(n10746), .ZN(n9767) );
  INV_X1 U12484 ( .A(n19810), .ZN(n10683) );
  NAND2_X2 U12485 ( .A1(n9776), .A2(n9775), .ZN(n14059) );
  INV_X1 U12486 ( .A(n10667), .ZN(n9777) );
  NAND2_X2 U12487 ( .A1(n10161), .A2(n10185), .ZN(n10667) );
  INV_X2 U12488 ( .A(n13295), .ZN(n10185) );
  AND2_X4 U12489 ( .A1(n9972), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12677) );
  AND2_X4 U12490 ( .A1(n9972), .A2(n16301), .ZN(n12678) );
  AND2_X2 U12491 ( .A1(n9793), .A2(n11487), .ZN(n11738) );
  AND2_X2 U12492 ( .A1(n9793), .A2(n11486), .ZN(n11593) );
  NAND3_X1 U12493 ( .A1(n9796), .A2(n9794), .A3(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n9803) );
  NAND3_X1 U12494 ( .A1(n13399), .A2(n9795), .A3(n9800), .ZN(n9794) );
  NAND2_X1 U12495 ( .A1(n9797), .A2(n9798), .ZN(n9796) );
  INV_X1 U12496 ( .A(n13399), .ZN(n9797) );
  INV_X1 U12497 ( .A(n13466), .ZN(n9798) );
  OAI211_X1 U12498 ( .C1(n9798), .C2(n13399), .A(n9799), .B(n9800), .ZN(n13465) );
  NAND2_X1 U12499 ( .A1(n13399), .A2(n9801), .ZN(n9799) );
  NOR2_X1 U12500 ( .A1(n13466), .A2(n13397), .ZN(n9801) );
  NAND2_X1 U12501 ( .A1(n9803), .A2(n9802), .ZN(n13627) );
  NAND2_X1 U12502 ( .A1(n9804), .A2(n9798), .ZN(n9802) );
  NAND2_X1 U12503 ( .A1(n9805), .A2(n10033), .ZN(n16008) );
  NAND3_X1 U12504 ( .A1(n14127), .A2(n16014), .A3(n14126), .ZN(n9805) );
  NAND2_X2 U12505 ( .A1(n9806), .A2(n14142), .ZN(n16010) );
  INV_X1 U12506 ( .A(n16008), .ZN(n9806) );
  INV_X2 U12507 ( .A(n13359), .ZN(n11635) );
  NAND3_X1 U12508 ( .A1(n11491), .A2(n11488), .A3(n11489), .ZN(n9808) );
  NAND3_X1 U12509 ( .A1(n11479), .A2(n11490), .A3(n11482), .ZN(n9809) );
  NAND2_X1 U12510 ( .A1(n10048), .A2(n9818), .ZN(n9814) );
  OAI211_X2 U12511 ( .C1(n14426), .C2(n9814), .A(n9813), .B(n9816), .ZN(n9815)
         );
  OR2_X1 U12512 ( .A1(n14426), .A2(n14398), .ZN(n14953) );
  NAND2_X1 U12513 ( .A1(n10048), .A2(n9817), .ZN(n9816) );
  NOR2_X2 U12514 ( .A1(n18786), .A2(n11361), .ZN(n18612) );
  INV_X2 U12515 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11361) );
  NAND3_X1 U12516 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .ZN(n9827) );
  INV_X1 U12517 ( .A(P3_EBX_REG_8__SCAN_IN), .ZN(n9828) );
  OAI21_X1 U12518 ( .B1(n16177), .B2(n19677), .A(n9833), .ZN(P2_U2825) );
  INV_X1 U12519 ( .A(n11247), .ZN(n9838) );
  NAND2_X1 U12520 ( .A1(n12526), .A2(n9842), .ZN(n9841) );
  NAND2_X1 U12521 ( .A1(n12536), .A2(n9846), .ZN(n9844) );
  OAI211_X1 U12522 ( .C1(n12536), .C2(n12718), .A(n9844), .B(n9845), .ZN(
        n15160) );
  OAI22_X1 U12523 ( .A1(n12488), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n19822), 
        .B2(n9789), .ZN(n11225) );
  INV_X1 U12524 ( .A(n11228), .ZN(n9851) );
  NAND2_X1 U12525 ( .A1(n9851), .A2(n9852), .ZN(n11223) );
  OAI21_X2 U12526 ( .B1(n9856), .B2(n9857), .A(n15119), .ZN(n15127) );
  NAND2_X2 U12527 ( .A1(n9857), .A2(n9856), .ZN(n15119) );
  NAND2_X2 U12528 ( .A1(n15131), .A2(n12759), .ZN(n9857) );
  AOI21_X1 U12529 ( .B1(n18876), .B2(n11219), .A(n11247), .ZN(n9858) );
  NAND2_X1 U12530 ( .A1(n11247), .A2(n15287), .ZN(n9859) );
  NAND3_X1 U12531 ( .A1(n11123), .A2(n11234), .A3(n11124), .ZN(n11229) );
  NAND2_X1 U12532 ( .A1(n11190), .A2(n9861), .ZN(n11206) );
  OR2_X2 U12533 ( .A1(n15258), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10602) );
  NAND3_X1 U12534 ( .A1(n15317), .A2(n15597), .A3(n11105), .ZN(n9865) );
  NAND4_X1 U12535 ( .A1(n9868), .A2(n10085), .A3(n10087), .A4(n10086), .ZN(
        n9867) );
  NAND4_X1 U12536 ( .A1(n9870), .A2(n10084), .A3(n10082), .A4(n10081), .ZN(
        n9869) );
  NAND2_X1 U12537 ( .A1(n10537), .A2(n9871), .ZN(n10559) );
  INV_X1 U12538 ( .A(n10505), .ZN(n9880) );
  NAND2_X1 U12539 ( .A1(n9880), .A2(n10506), .ZN(n10521) );
  OR2_X1 U12540 ( .A1(n15437), .A2(n19174), .ZN(n9882) );
  NAND2_X1 U12541 ( .A1(n9886), .A2(n9883), .ZN(n13798) );
  NAND2_X1 U12542 ( .A1(n9888), .A2(n9649), .ZN(n14317) );
  NAND2_X1 U12543 ( .A1(n14756), .A2(n9697), .ZN(n15797) );
  INV_X2 U12544 ( .A(n16805), .ZN(n16845) );
  OAI21_X1 U12545 ( .B1(n17676), .B2(n9934), .A(n17656), .ZN(n12967) );
  NAND2_X1 U12546 ( .A1(n9931), .A2(n9930), .ZN(n17611) );
  NAND2_X1 U12547 ( .A1(n12965), .A2(n17730), .ZN(n9930) );
  NAND3_X1 U12548 ( .A1(n9933), .A2(n12965), .A3(n9932), .ZN(n9931) );
  INV_X1 U12549 ( .A(n17676), .ZN(n9933) );
  AND2_X1 U12550 ( .A1(n9936), .A2(n11705), .ZN(n11708) );
  XNOR2_X2 U12551 ( .A(n9936), .B(n11652), .ZN(n11773) );
  OR2_X2 U12552 ( .A1(n11755), .A2(n11754), .ZN(n11798) );
  NAND2_X1 U12553 ( .A1(n11569), .A2(n9938), .ZN(n11545) );
  NAND2_X1 U12554 ( .A1(n9940), .A2(n9939), .ZN(n13792) );
  INV_X1 U12555 ( .A(n13791), .ZN(n9939) );
  NAND2_X1 U12556 ( .A1(n9687), .A2(n9940), .ZN(n16020) );
  NAND2_X1 U12557 ( .A1(n20371), .A2(n11760), .ZN(n9941) );
  NAND2_X1 U12558 ( .A1(n9941), .A2(n9943), .ZN(n13565) );
  INV_X1 U12559 ( .A(n13565), .ZN(n9942) );
  NAND2_X1 U12560 ( .A1(n9942), .A2(n11778), .ZN(n13562) );
  NAND3_X1 U12561 ( .A1(n11880), .A2(n9618), .A3(n11895), .ZN(n14093) );
  AND3_X2 U12562 ( .A1(n11880), .A2(n9618), .A3(n9696), .ZN(n14094) );
  AND2_X1 U12563 ( .A1(n14623), .A2(n14622), .ZN(n14607) );
  NAND2_X1 U12564 ( .A1(n14623), .A2(n9950), .ZN(n14608) );
  AND2_X2 U12565 ( .A1(n14623), .A2(n9948), .ZN(n14480) );
  XNOR2_X2 U12566 ( .A(n14480), .B(n12320), .ZN(n14599) );
  NAND2_X1 U12567 ( .A1(n14358), .A2(n9692), .ZN(n14709) );
  OAI22_X1 U12568 ( .A1(n14501), .A2(n9956), .B1(n14503), .B2(n14502), .ZN(
        n14521) );
  AND2_X2 U12569 ( .A1(n10717), .A2(n10716), .ZN(n9956) );
  OAI21_X1 U12570 ( .B1(n13700), .B2(n9959), .A(n9957), .ZN(n10714) );
  OAI21_X1 U12571 ( .B1(n13699), .B2(n9959), .A(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n9958) );
  INV_X1 U12572 ( .A(n10710), .ZN(n9959) );
  XNOR2_X2 U12573 ( .A(n10711), .B(n10702), .ZN(n13700) );
  NAND2_X1 U12574 ( .A1(n10723), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9962) );
  NOR2_X1 U12575 ( .A1(n9972), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13953) );
  NOR2_X1 U12576 ( .A1(n13964), .A2(n9972), .ZN(n13965) );
  NAND4_X1 U12577 ( .A1(n10124), .A2(n9974), .A3(n10123), .A4(n10125), .ZN(
        n9973) );
  NAND4_X1 U12578 ( .A1(n10119), .A2(n9976), .A3(n10120), .A4(n10122), .ZN(
        n9975) );
  NAND2_X1 U12579 ( .A1(n10763), .A2(n9643), .ZN(n13658) );
  NAND2_X1 U12580 ( .A1(n15074), .A2(n15135), .ZN(n15137) );
  NAND3_X1 U12581 ( .A1(n10002), .A2(n10001), .A3(n10927), .ZN(n10932) );
  OAI21_X1 U12582 ( .B1(n19222), .B2(n12560), .A(n10010), .ZN(n10374) );
  INV_X1 U12583 ( .A(n12498), .ZN(n13670) );
  AND4_X2 U12584 ( .A1(n9672), .A2(n10602), .A3(n10603), .A4(n10012), .ZN(
        n10624) );
  AND2_X2 U12585 ( .A1(n15239), .A2(n15247), .ZN(n10012) );
  OAI21_X1 U12586 ( .B1(n15268), .B2(n10017), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10016) );
  INV_X1 U12587 ( .A(n10016), .ZN(n10015) );
  NAND2_X1 U12588 ( .A1(n10018), .A2(n10019), .ZN(n15369) );
  NOR2_X4 U12589 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13347) );
  INV_X1 U12590 ( .A(n16013), .ZN(n10031) );
  INV_X1 U12591 ( .A(n14129), .ZN(n10032) );
  INV_X1 U12592 ( .A(n14847), .ZN(n14411) );
  NAND2_X2 U12593 ( .A1(n15962), .A2(n14412), .ZN(n14847) );
  NAND3_X1 U12594 ( .A1(n14412), .A2(n15962), .A3(n14410), .ZN(n10035) );
  NAND2_X1 U12595 ( .A1(n10035), .A2(n10059), .ZN(n14869) );
  NAND2_X1 U12596 ( .A1(n11773), .A2(n20756), .ZN(n10046) );
  NAND3_X1 U12597 ( .A1(n10037), .A2(n9640), .A3(n10036), .ZN(n13249) );
  NAND3_X1 U12598 ( .A1(n10037), .A2(n9671), .A3(n10036), .ZN(n13252) );
  NAND2_X1 U12599 ( .A1(n11773), .A2(n10038), .ZN(n10037) );
  NAND2_X1 U12600 ( .A1(n16010), .A2(n10047), .ZN(n14397) );
  NAND2_X1 U12601 ( .A1(n11195), .A2(n19188), .ZN(n11101) );
  OR2_X1 U12602 ( .A1(n16172), .A2(n19179), .ZN(n10068) );
  NAND2_X1 U12603 ( .A1(n14503), .A2(n14500), .ZN(n10721) );
  OR2_X1 U12604 ( .A1(n15410), .A2(n19004), .ZN(n11275) );
  OAI21_X2 U12605 ( .B1(n14720), .B2(n14726), .A(n14719), .ZN(n15829) );
  MUX2_X2 U12606 ( .A(n14842), .B(n14841), .S(n15987), .Z(n14843) );
  OR2_X1 U12607 ( .A1(n15377), .A2(n16257), .ZN(n15390) );
  AND2_X1 U12608 ( .A1(n14815), .A2(n13417), .ZN(n15947) );
  AND2_X1 U12609 ( .A1(n19069), .A2(n12860), .ZN(n19099) );
  CLKBUF_X1 U12610 ( .A(n13094), .Z(n14582) );
  NAND2_X1 U12611 ( .A1(n10887), .A2(n10886), .ZN(n11039) );
  AND2_X1 U12612 ( .A1(n14418), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14419) );
  INV_X1 U12613 ( .A(n13609), .ZN(n10763) );
  AND3_X1 U12614 ( .A1(n10552), .A2(P2_EBX_REG_21__SCAN_IN), .A3(n12848), .ZN(
        n10553) );
  AND2_X1 U12615 ( .A1(n12848), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10564) );
  AND2_X1 U12616 ( .A1(n12848), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10507) );
  NAND2_X1 U12617 ( .A1(n9594), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10228) );
  AOI21_X1 U12618 ( .B1(n12494), .B2(n11175), .A(n11174), .ZN(n11187) );
  AND2_X1 U12619 ( .A1(n11620), .A2(n13907), .ZN(n14145) );
  INV_X1 U12620 ( .A(n11761), .ZN(n11764) );
  AOI22_X1 U12621 ( .A1(n11513), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12202), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11559) );
  NOR2_X1 U12622 ( .A1(n14569), .A2(n12815), .ZN(n12840) );
  AND2_X1 U12623 ( .A1(n12498), .A2(n12519), .ZN(n10267) );
  OR2_X1 U12624 ( .A1(n10524), .A2(n15378), .ZN(n10050) );
  AND2_X1 U12625 ( .A1(n15945), .A2(n11631), .ZN(n15942) );
  INV_X2 U12626 ( .A(n9651), .ZN(n17125) );
  AND2_X1 U12627 ( .A1(n10570), .A2(n15368), .ZN(n10051) );
  OR2_X1 U12628 ( .A1(n16875), .A2(n13004), .ZN(n10052) );
  INV_X1 U12629 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16339) );
  AND2_X1 U12630 ( .A1(n11874), .A2(n11873), .ZN(n10053) );
  AND3_X1 U12631 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(P3_EBX_REG_16__SCAN_IN), 
        .A3(P3_EBX_REG_17__SCAN_IN), .ZN(n10054) );
  NOR2_X1 U12632 ( .A1(n14146), .A2(n11709), .ZN(n10055) );
  AND2_X1 U12633 ( .A1(n11633), .A2(n11626), .ZN(n10056) );
  AND2_X4 U12634 ( .A1(n14149), .A2(n14148), .ZN(n10059) );
  AND4_X1 U12635 ( .A1(n12901), .A2(n12900), .A3(n12899), .A4(n12898), .ZN(
        n10060) );
  XOR2_X1 U12636 ( .A(n15043), .B(n14926), .Z(n10061) );
  AND3_X1 U12637 ( .A1(n18012), .A2(n17650), .A3(n12963), .ZN(n10062) );
  INV_X1 U12638 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12963) );
  NAND2_X1 U12639 ( .A1(n9938), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11975) );
  INV_X1 U12640 ( .A(n11975), .ZN(n12003) );
  AND2_X1 U12641 ( .A1(n10931), .A2(n10930), .ZN(n10063) );
  AND2_X1 U12642 ( .A1(n11106), .A2(n10570), .ZN(n10064) );
  AND2_X1 U12643 ( .A1(n10212), .A2(n10664), .ZN(n10065) );
  AND2_X1 U12644 ( .A1(n10068), .A2(n11099), .ZN(n10066) );
  OR2_X1 U12645 ( .A1(n11288), .A2(n11287), .ZN(P2_U2824) );
  NAND2_X1 U12646 ( .A1(n15157), .A2(n14046), .ZN(n15124) );
  NAND2_X1 U12647 ( .A1(n11707), .A2(n11706), .ZN(n20149) );
  OR2_X1 U12648 ( .A1(n19692), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n19838) );
  INV_X1 U12649 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n11911) );
  AND2_X1 U12650 ( .A1(n19798), .A2(n10692), .ZN(n10069) );
  INV_X1 U12651 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n13902) );
  INV_X1 U12652 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n16238) );
  INV_X1 U12653 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19784) );
  OR2_X1 U12654 ( .A1(n17656), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10070) );
  AND2_X1 U12655 ( .A1(n10517), .A2(n10946), .ZN(n16257) );
  INV_X1 U12656 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n11202) );
  OR2_X1 U12657 ( .A1(n14395), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10071) );
  AND3_X1 U12658 ( .A1(n13043), .A2(n13042), .A3(n13041), .ZN(n10072) );
  NOR2_X1 U12659 ( .A1(n17823), .A2(n17794), .ZN(n17548) );
  INV_X1 U12660 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19775) );
  INV_X1 U12661 ( .A(n13651), .ZN(n12530) );
  OR2_X1 U12662 ( .A1(n18262), .A2(n18239), .ZN(n18264) );
  AND2_X1 U12663 ( .A1(n12755), .A2(n12775), .ZN(n10074) );
  AND3_X1 U12664 ( .A1(n15296), .A2(n10571), .A3(n10051), .ZN(n10075) );
  INV_X1 U12665 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n13937) );
  INV_X1 U12666 ( .A(n10720), .ZN(n10722) );
  AND2_X1 U12667 ( .A1(n19818), .A2(n10216), .ZN(n10076) );
  INV_X1 U12668 ( .A(n13862), .ZN(n19151) );
  NAND3_X2 U12669 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19764), .A3(n19533), 
        .ZN(n13862) );
  AND2_X2 U12670 ( .A1(n11483), .A2(n11484), .ZN(n11744) );
  AND2_X1 U12671 ( .A1(n11642), .A2(n13280), .ZN(n10078) );
  AND2_X1 U12672 ( .A1(n11631), .A2(n11569), .ZN(n10079) );
  NAND2_X1 U12673 ( .A1(n12353), .A2(n12352), .ZN(n12362) );
  INV_X1 U12674 ( .A(n13470), .ZN(n11709) );
  OR2_X1 U12675 ( .A1(n12362), .A2(n20120), .ZN(n12382) );
  OR2_X1 U12676 ( .A1(n11862), .A2(n11861), .ZN(n14137) );
  INV_X1 U12677 ( .A(n12382), .ZN(n12384) );
  NOR2_X1 U12678 ( .A1(n11620), .A2(n13907), .ZN(n11621) );
  INV_X1 U12679 ( .A(n11640), .ZN(n11622) );
  NAND2_X1 U12680 ( .A1(n10228), .A2(n10227), .ZN(n10229) );
  AND2_X1 U12681 ( .A1(n10663), .A2(n14046), .ZN(n10192) );
  MUX2_X1 U12682 ( .A(n12860), .B(n13295), .S(n14059), .Z(n10164) );
  INV_X1 U12683 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13409) );
  OR2_X1 U12684 ( .A1(n12160), .A2(n14710), .ZN(n12180) );
  OR2_X1 U12685 ( .A1(n11665), .A2(n11664), .ZN(n14151) );
  OR2_X1 U12686 ( .A1(n11818), .A2(n11817), .ZN(n13841) );
  OR2_X1 U12687 ( .A1(n11750), .A2(n11749), .ZN(n13469) );
  OR2_X1 U12688 ( .A1(n11676), .A2(n11675), .ZN(n13471) );
  NAND2_X1 U12689 ( .A1(n10662), .A2(n19830), .ZN(n10197) );
  NAND2_X1 U12690 ( .A1(n12758), .A2(n10074), .ZN(n12759) );
  OR2_X1 U12691 ( .A1(n10332), .A2(n10331), .ZN(n10902) );
  NOR2_X1 U12692 ( .A1(n11359), .A2(n12442), .ZN(n11360) );
  NAND2_X1 U12693 ( .A1(n11651), .A2(n9659), .ZN(n11705) );
  NAND2_X1 U12694 ( .A1(n14472), .A2(n13409), .ZN(n13411) );
  AND2_X1 U12695 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n12219), .ZN(
        n12220) );
  INV_X1 U12696 ( .A(n11969), .ZN(n11970) );
  NAND2_X1 U12697 ( .A1(n9665), .A2(n14145), .ZN(n13847) );
  OAI21_X1 U12698 ( .B1(n10902), .B2(n19809), .A(n10447), .ZN(n10680) );
  INV_X1 U12699 ( .A(n10609), .ZN(n10610) );
  INV_X1 U12700 ( .A(n10197), .ZN(n10198) );
  AND2_X1 U12701 ( .A1(n16258), .A2(n16255), .ZN(n10510) );
  AND2_X1 U12702 ( .A1(n15294), .A2(n10075), .ZN(n15279) );
  AND4_X1 U12703 ( .A1(n10431), .A2(n10430), .A3(n10429), .A4(n10428), .ZN(
        n10441) );
  AOI22_X1 U12704 ( .A1(n12677), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12678), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10132) );
  INV_X1 U12705 ( .A(n10462), .ZN(n10918) );
  OR2_X1 U12706 ( .A1(n12753), .A2(n12507), .ZN(n12511) );
  INV_X1 U12707 ( .A(n12987), .ZN(n18608) );
  INV_X1 U12708 ( .A(n11705), .ZN(n11652) );
  OR2_X1 U12709 ( .A1(n12159), .A2(n14717), .ZN(n14710) );
  NOR2_X1 U12710 ( .A1(n11631), .A2(n20752), .ZN(n12319) );
  NAND2_X1 U12711 ( .A1(n12220), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12265) );
  NOR2_X1 U12712 ( .A1(n12114), .A2(n14900), .ZN(n12177) );
  NAND2_X1 U12713 ( .A1(n11970), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11978) );
  AOI21_X1 U12714 ( .B1(n14135), .B2(n12003), .A(n11879), .ZN(n13876) );
  NAND2_X1 U12715 ( .A1(n14876), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15954) );
  OR2_X1 U12716 ( .A1(n15986), .A2(n14917), .ZN(n14920) );
  INV_X1 U12717 ( .A(n16007), .ZN(n14142) );
  OR2_X1 U12718 ( .A1(n11794), .A2(n11793), .ZN(n13631) );
  AND2_X1 U12719 ( .A1(n20218), .A2(n20602), .ZN(n20220) );
  NOR2_X1 U12720 ( .A1(n20491), .A2(n20490), .ZN(n20594) );
  OAI21_X1 U12721 ( .B1(n15172), .B2(n19001), .A(n11283), .ZN(n11284) );
  NOR2_X1 U12722 ( .A1(n10618), .A2(n10610), .ZN(n11181) );
  AND2_X1 U12723 ( .A1(n12848), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10545) );
  AOI221_X1 U12724 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n10640), 
        .C1(n16339), .C2(n10640), .A(n10639), .ZN(n10684) );
  OR2_X1 U12725 ( .A1(n10979), .A2(n10978), .ZN(n12531) );
  OR2_X1 U12726 ( .A1(n12754), .A2(n12756), .ZN(n12775) );
  AND4_X2 U12727 ( .A1(n10442), .A2(n10441), .A3(n10440), .A4(n10439), .ZN(
        n10733) );
  AOI21_X1 U12728 ( .B1(n13963), .B2(n12510), .A(n12509), .ZN(n13526) );
  AND2_X1 U12729 ( .A1(n10267), .A2(n10276), .ZN(n14019) );
  INV_X1 U12730 ( .A(n10362), .ZN(n19524) );
  INV_X1 U12731 ( .A(n14068), .ZN(n14074) );
  NOR2_X1 U12732 ( .A1(n17536), .A2(n17503), .ZN(n12416) );
  AOI22_X1 U12733 ( .A1(n12966), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B1(
        n17962), .B2(n17730), .ZN(n12965) );
  NOR2_X1 U12734 ( .A1(n13027), .A2(n17762), .ZN(n13029) );
  INV_X1 U12735 ( .A(n17333), .ZN(n13025) );
  NOR4_X1 U12736 ( .A1(n12425), .A2(n12433), .A3(n12435), .A4(n12424), .ZN(
        n12438) );
  AND2_X1 U12737 ( .A1(n14457), .A2(n14456), .ZN(n14721) );
  INV_X1 U12738 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n14687) );
  INV_X1 U12739 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n13992) );
  AND2_X1 U12740 ( .A1(n14369), .A2(n14368), .ZN(n14370) );
  OR2_X1 U12741 ( .A1(n14727), .A2(n14732), .ZN(n14717) );
  INV_X1 U12742 ( .A(n15947), .ZN(n14817) );
  INV_X1 U12743 ( .A(n19971), .ZN(n20031) );
  OR2_X1 U12744 ( .A1(n12224), .A2(n12223), .ZN(n14652) );
  NAND2_X1 U12745 ( .A1(n12177), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12176) );
  NAND2_X1 U12746 ( .A1(n12062), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12114) );
  INV_X1 U12747 ( .A(n11976), .ZN(n11977) );
  OR2_X1 U12748 ( .A1(n11896), .A2(n13992), .ZN(n11912) );
  AND2_X1 U12749 ( .A1(n11848), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11863) );
  AND2_X1 U12750 ( .A1(n13402), .A2(n14579), .ZN(n15750) );
  AND2_X1 U12751 ( .A1(n16151), .A2(n20756), .ZN(n13403) );
  AND2_X1 U12752 ( .A1(n13478), .A2(n13477), .ZN(n14539) );
  NAND2_X1 U12753 ( .A1(n11783), .A2(n11782), .ZN(n20259) );
  AND2_X1 U12754 ( .A1(n12392), .A2(n12391), .ZN(n14589) );
  OR2_X1 U12755 ( .A1(n20217), .A2(n20343), .ZN(n20262) );
  NOR2_X1 U12756 ( .A1(n20106), .A2(n20265), .ZN(n20430) );
  INV_X1 U12757 ( .A(n20371), .ZN(n20372) );
  NOR2_X1 U12758 ( .A1(n20266), .A2(n20265), .ZN(n20556) );
  NAND3_X1 U12759 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20756), .A3(n20104), 
        .ZN(n20142) );
  INV_X1 U12760 ( .A(n16163), .ZN(n16159) );
  INV_X1 U12761 ( .A(n11284), .ZN(n11285) );
  INV_X1 U12762 ( .A(n19809), .ZN(n11252) );
  NAND2_X1 U12763 ( .A1(n19019), .A2(n12510), .ZN(n12506) );
  INV_X1 U12764 ( .A(n19038), .ZN(n15208) );
  INV_X1 U12765 ( .A(n19039), .ZN(n15210) );
  AND2_X1 U12766 ( .A1(n10921), .A2(n10920), .ZN(n19000) );
  OAI21_X1 U12767 ( .B1(n10626), .B2(n12461), .A(n10625), .ZN(n15221) );
  NOR3_X1 U12768 ( .A1(n11109), .A2(n15305), .A3(n15319), .ZN(n11110) );
  AND2_X1 U12769 ( .A1(n13525), .A2(n10002), .ZN(n19777) );
  INV_X1 U12770 ( .A(n19274), .ZN(n19348) );
  OR2_X1 U12771 ( .A1(n19782), .A2(n19787), .ZN(n19193) );
  NAND2_X1 U12772 ( .A1(n19782), .A2(n19787), .ZN(n14047) );
  NAND2_X1 U12773 ( .A1(n15697), .A2(n15700), .ZN(n12985) );
  NOR2_X1 U12774 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16656), .ZN(n16644) );
  NOR2_X1 U12775 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16752), .ZN(n16734) );
  NAND2_X1 U12776 ( .A1(n18806), .A2(n18814), .ZN(n12452) );
  INV_X1 U12777 ( .A(n17188), .ZN(n11396) );
  INV_X1 U12778 ( .A(n15720), .ZN(n17837) );
  NOR2_X1 U12779 ( .A1(n17816), .A2(n12410), .ZN(n12420) );
  INV_X1 U12780 ( .A(n17966), .ZN(n17885) );
  INV_X1 U12781 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16763) );
  INV_X1 U12782 ( .A(n17817), .ZN(n17781) );
  NOR2_X1 U12783 ( .A1(n17502), .A2(n17834), .ZN(n17830) );
  NOR2_X1 U12784 ( .A1(n17698), .A2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n17688) );
  INV_X1 U12785 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18636) );
  NOR2_X1 U12786 ( .A1(n11316), .A2(n11315), .ZN(n18187) );
  INV_X1 U12787 ( .A(n13095), .ZN(n15762) );
  NOR2_X1 U12788 ( .A1(n14589), .A2(n19845), .ZN(n13262) );
  AND2_X1 U12789 ( .A1(n15837), .A2(n13903), .ZN(n19904) );
  NOR2_X1 U12790 ( .A1(n19847), .A2(n15918), .ZN(n19913) );
  AND2_X1 U12791 ( .A1(n15837), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19926) );
  AND2_X1 U12792 ( .A1(n13915), .A2(n13909), .ZN(n19945) );
  INV_X1 U12793 ( .A(n15945), .ZN(n14763) );
  NOR2_X1 U12794 ( .A1(n15952), .A2(n16425), .ZN(n12406) );
  AND2_X1 U12795 ( .A1(n12125), .A2(n12124), .ZN(n14720) );
  INV_X1 U12796 ( .A(n15952), .ZN(n14819) );
  NOR2_X1 U12797 ( .A1(n19950), .A2(n20761), .ZN(n19967) );
  BUF_X1 U12798 ( .A(n14709), .Z(n15857) );
  NAND2_X1 U12799 ( .A1(n12028), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12060) );
  NAND2_X1 U12800 ( .A1(n11929), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11969) );
  AND2_X1 U12801 ( .A1(n16026), .A2(n20090), .ZN(n16021) );
  AND2_X1 U12802 ( .A1(n15750), .A2(n14598), .ZN(n20093) );
  AND2_X1 U12803 ( .A1(n13403), .A2(n20752), .ZN(n16052) );
  AND2_X1 U12804 ( .A1(n15979), .A2(n15978), .ZN(n16071) );
  INV_X1 U12805 ( .A(n14539), .ZN(n15059) );
  NOR2_X1 U12806 ( .A1(n16083), .A2(n15060), .ZN(n16143) );
  AND2_X1 U12807 ( .A1(n13289), .A2(n13270), .ZN(n16144) );
  NOR2_X1 U12808 ( .A1(n20493), .A2(n14589), .ZN(n14561) );
  NAND2_X1 U12809 ( .A1(n20730), .A2(n9620), .ZN(n20217) );
  INV_X1 U12810 ( .A(n20262), .ZN(n20284) );
  INV_X1 U12811 ( .A(n20729), .ZN(n20313) );
  INV_X1 U12812 ( .A(n20361), .ZN(n20366) );
  INV_X1 U12813 ( .A(n20370), .ZN(n20395) );
  INV_X1 U12814 ( .A(n20487), .ZN(n20551) );
  AND2_X1 U12815 ( .A1(n20457), .A2(n20403), .ZN(n20447) );
  OAI22_X1 U12816 ( .A1(n20497), .A2(n20496), .B1(n20549), .B2(n20495), .ZN(
        n20514) );
  INV_X1 U12817 ( .A(n20545), .ZN(n20513) );
  OR2_X1 U12818 ( .A1(n9620), .A2(n20258), .ZN(n20603) );
  INV_X1 U12819 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20663) );
  INV_X1 U12820 ( .A(n20706), .ZN(n20716) );
  AND2_X1 U12821 ( .A1(n10694), .A2(n10693), .ZN(n11113) );
  INV_X1 U12822 ( .A(n16166), .ZN(n16167) );
  OR2_X1 U12823 ( .A1(n19819), .A2(n11261), .ZN(n18978) );
  AND2_X1 U12824 ( .A1(n19819), .A2(n16351), .ZN(n19016) );
  AND2_X1 U12825 ( .A1(n9633), .A2(n14086), .ZN(n14252) );
  INV_X1 U12826 ( .A(n12534), .ZN(n13929) );
  XNOR2_X1 U12827 ( .A(n12736), .B(n12737), .ZN(n15143) );
  NAND2_X1 U12828 ( .A1(n15160), .A2(n15159), .ZN(n15158) );
  AND2_X1 U12829 ( .A1(n14250), .A2(n14249), .ZN(n14383) );
  AND2_X1 U12830 ( .A1(n13301), .A2(n13190), .ZN(n19038) );
  INV_X1 U12831 ( .A(n19069), .ZN(n19098) );
  INV_X1 U12832 ( .A(n13176), .ZN(n13152) );
  AND2_X1 U12833 ( .A1(n13102), .A2(n11264), .ZN(n13112) );
  INV_X1 U12834 ( .A(n19148), .ZN(n16261) );
  AND2_X1 U12835 ( .A1(n19154), .A2(n13310), .ZN(n19141) );
  INV_X1 U12836 ( .A(n13670), .ZN(n16289) );
  INV_X1 U12837 ( .A(n19154), .ZN(n15338) );
  INV_X1 U12838 ( .A(n16203), .ZN(n15466) );
  INV_X1 U12839 ( .A(n19157), .ZN(n19188) );
  INV_X1 U12840 ( .A(n19533), .ZN(n19565) );
  OAI21_X1 U12841 ( .B1(n19200), .B2(n19199), .A(n19198), .ZN(n19218) );
  AND2_X1 U12842 ( .A1(n19076), .A2(n19030), .ZN(n19274) );
  INV_X1 U12843 ( .A(n19244), .ZN(n19267) );
  NOR2_X2 U12844 ( .A1(n19348), .A2(n19487), .ZN(n19343) );
  INV_X1 U12845 ( .A(n19366), .ZN(n19373) );
  NOR2_X1 U12846 ( .A1(n19348), .A2(n19562), .ZN(n19399) );
  INV_X1 U12847 ( .A(n19193), .ZN(n19228) );
  INV_X1 U12848 ( .A(n19447), .ZN(n19453) );
  NOR2_X1 U12849 ( .A1(n19523), .A2(n19487), .ZN(n19508) );
  INV_X1 U12850 ( .A(n19598), .ZN(n19549) );
  INV_X1 U12851 ( .A(n14195), .ZN(n19573) );
  NOR2_X1 U12852 ( .A1(n19523), .A2(n19562), .ZN(n19599) );
  INV_X1 U12853 ( .A(n19561), .ZN(n19630) );
  INV_X1 U12854 ( .A(n19583), .ZN(n19638) );
  AND2_X1 U12855 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10700), .ZN(n19673) );
  NAND2_X1 U12856 ( .A1(n18652), .A2(n18596), .ZN(n17355) );
  NOR2_X1 U12857 ( .A1(n18622), .A2(n12985), .ZN(n18595) );
  NOR2_X1 U12858 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16637), .ZN(n16624) );
  NOR2_X1 U12859 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16702), .ZN(n16685) );
  INV_X1 U12860 ( .A(n12448), .ZN(n16888) );
  NOR2_X1 U12861 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16756), .ZN(n16755) );
  NOR2_X1 U12862 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16799), .ZN(n16772) );
  INV_X1 U12863 ( .A(n16891), .ZN(n16862) );
  INV_X1 U12864 ( .A(n16888), .ZN(n16883) );
  NOR2_X1 U12865 ( .A1(n11385), .A2(n11384), .ZN(n18160) );
  INV_X1 U12866 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17121) );
  INV_X1 U12867 ( .A(n17266), .ZN(n17263) );
  NOR2_X1 U12868 ( .A1(n17211), .A2(n18182), .ZN(n18630) );
  OR3_X1 U12869 ( .A1(n15808), .A2(n18814), .A3(n9732), .ZN(n15809) );
  NOR2_X1 U12870 ( .A1(n17877), .A2(n17626), .ZN(n17540) );
  NAND2_X1 U12871 ( .A1(n17647), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17966) );
  NOR2_X1 U12872 ( .A1(n18006), .A2(n18142), .ZN(n18038) );
  INV_X1 U12873 ( .A(n18043), .ZN(n18058) );
  INV_X1 U12874 ( .A(n18141), .ZN(n18100) );
  INV_X1 U12875 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18773) );
  INV_X1 U12876 ( .A(n18286), .ZN(n18279) );
  INV_X1 U12877 ( .A(n18308), .ZN(n18301) );
  INV_X1 U12878 ( .A(n18329), .ZN(n18322) );
  INV_X1 U12879 ( .A(n18582), .ZN(n18493) );
  NOR2_X1 U12880 ( .A1(n18664), .A2(n18661), .ZN(n18652) );
  NOR2_X1 U12881 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13050), .ZN(n16497)
         );
  INV_X1 U12882 ( .A(U212), .ZN(n20925) );
  NAND2_X1 U12883 ( .A1(n13262), .A2(n15762), .ZN(n19841) );
  INV_X1 U12884 ( .A(n19945), .ZN(n19897) );
  INV_X1 U12885 ( .A(n19913), .ZN(n15929) );
  INV_X1 U12886 ( .A(n19904), .ZN(n15891) );
  AND2_X1 U12887 ( .A1(n15891), .A2(n13905), .ZN(n19949) );
  NAND2_X1 U12888 ( .A1(n15945), .A2(n20141), .ZN(n14761) );
  NAND2_X1 U12889 ( .A1(n14815), .A2(n13416), .ZN(n14828) );
  INV_X1 U12890 ( .A(n19950), .ZN(n19970) );
  INV_X1 U12891 ( .A(n16021), .ZN(n16019) );
  INV_X1 U12892 ( .A(n20093), .ZN(n19850) );
  INV_X1 U12893 ( .A(n16052), .ZN(n16103) );
  INV_X1 U12894 ( .A(n16144), .ZN(n16111) );
  INV_X1 U12895 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20098) );
  OR2_X1 U12896 ( .A1(n20217), .A2(n20487), .ZN(n20175) );
  OR2_X1 U12897 ( .A1(n20217), .A2(n20525), .ZN(n20210) );
  OR2_X1 U12898 ( .A1(n20217), .A2(n20312), .ZN(n20257) );
  NAND2_X1 U12899 ( .A1(n20313), .A2(n20551), .ZN(n20311) );
  OR2_X1 U12900 ( .A1(n20729), .A2(n20525), .ZN(n20336) );
  OR2_X1 U12901 ( .A1(n20729), .A2(n20312), .ZN(n20361) );
  NAND2_X1 U12902 ( .A1(n20457), .A2(n20551), .ZN(n20423) );
  INV_X1 U12903 ( .A(n20447), .ZN(n20455) );
  INV_X1 U12904 ( .A(n20483), .ZN(n20478) );
  NAND2_X1 U12905 ( .A1(n20457), .A2(n20456), .ZN(n20518) );
  OR2_X1 U12906 ( .A1(n20603), .A2(n20487), .ZN(n20545) );
  NAND2_X1 U12907 ( .A1(n20547), .A2(n20546), .ZN(n20657) );
  OR2_X1 U12908 ( .A1(n20660), .A2(n20756), .ZN(n19845) );
  NOR2_X1 U12909 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20663), .ZN(n20750) );
  AND2_X1 U12910 ( .A1(n13102), .A2(n16323), .ZN(n19819) );
  OR2_X1 U12911 ( .A1(n11113), .A2(n11112), .ZN(n13110) );
  NAND2_X1 U12912 ( .A1(n11275), .A2(n11274), .ZN(n11276) );
  INV_X1 U12913 ( .A(n19016), .ZN(n19001) );
  OR2_X1 U12914 ( .A1(n14383), .A2(n14382), .ZN(n16220) );
  INV_X1 U12915 ( .A(n15169), .ZN(n15157) );
  INV_X1 U12916 ( .A(n19071), .ZN(n19107) );
  INV_X1 U12917 ( .A(n19109), .ZN(n19139) );
  OAI21_X1 U12918 ( .B1(n19695), .B2(n13111), .A(n13225), .ZN(n13176) );
  CLKBUF_X1 U12919 ( .A(n13176), .Z(n13224) );
  OR2_X1 U12920 ( .A1(n11148), .A2(n19148), .ZN(n11133) );
  NAND2_X1 U12921 ( .A1(n11132), .A2(n12780), .ZN(n19148) );
  OR2_X1 U12922 ( .A1(n11196), .A2(n19174), .ZN(n11100) );
  OR2_X1 U12923 ( .A1(n11148), .A2(n19174), .ZN(n11149) );
  OR3_X1 U12924 ( .A1(n11088), .A2(n19809), .A3(n19810), .ZN(n19157) );
  OR2_X1 U12925 ( .A1(n11088), .A2(n19806), .ZN(n19174) );
  INV_X1 U12926 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15807) );
  NAND2_X1 U12927 ( .A1(n19228), .A2(n19274), .ZN(n19244) );
  INV_X1 U12928 ( .A(n19241), .ZN(n19254) );
  AOI21_X1 U12929 ( .B1(n14184), .B2(n19764), .A(n14183), .ZN(n19270) );
  AOI21_X1 U12930 ( .B1(n19275), .B2(n19279), .A(n19273), .ZN(n19308) );
  AND3_X1 U12931 ( .A1(n19316), .A2(n19315), .A3(n19533), .ZN(n19347) );
  OR2_X1 U12932 ( .A1(n19312), .A2(n19562), .ZN(n19366) );
  INV_X1 U12933 ( .A(n19399), .ZN(n19407) );
  INV_X1 U12934 ( .A(n19421), .ZN(n19419) );
  NAND2_X1 U12935 ( .A1(n14013), .A2(n19228), .ZN(n19447) );
  NOR2_X1 U12936 ( .A1(n14012), .A2(n14011), .ZN(n15676) );
  INV_X1 U12937 ( .A(n19508), .ZN(n19522) );
  AND2_X1 U12938 ( .A1(n19569), .A2(n19568), .ZN(n19580) );
  INV_X1 U12939 ( .A(n19599), .ZN(n19609) );
  AOI21_X1 U12940 ( .B1(n14109), .B2(n14108), .A(n14107), .ZN(n19636) );
  AND2_X1 U12941 ( .A1(n16354), .A2(n16353), .ZN(n19679) );
  INV_X1 U12942 ( .A(n19761), .ZN(n19680) );
  OR2_X2 U12943 ( .A1(n18603), .A2(n18811), .ZN(n16521) );
  NOR2_X1 U12944 ( .A1(n12456), .A2(n12455), .ZN(n12457) );
  INV_X1 U12945 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17549) );
  INV_X1 U12946 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17685) );
  INV_X1 U12947 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16780) );
  INV_X1 U12948 ( .A(n16876), .ZN(n16875) );
  NOR2_X1 U12949 ( .A1(n16904), .A2(n16903), .ZN(n16930) );
  INV_X1 U12950 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17176) );
  INV_X1 U12951 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17181) );
  INV_X1 U12952 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17198) );
  AND2_X1 U12953 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17301), .ZN(n17304) );
  INV_X1 U12954 ( .A(n16409), .ZN(n17322) );
  NAND2_X1 U12955 ( .A1(n17357), .A2(n18814), .ZN(n17382) );
  NAND2_X1 U12956 ( .A1(n17414), .A2(n17356), .ZN(n17412) );
  INV_X1 U12957 ( .A(n17460), .ZN(n17456) );
  NAND2_X1 U12958 ( .A1(n17936), .A2(n17717), .ZN(n17626) );
  NAND2_X1 U12959 ( .A1(n16409), .A2(n17797), .ZN(n17721) );
  INV_X1 U12960 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n18012) );
  NAND2_X1 U12961 ( .A1(n17632), .A2(n13007), .ZN(n18063) );
  INV_X1 U12962 ( .A(n18125), .ZN(n18142) );
  INV_X1 U12963 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18634) );
  INV_X1 U12964 ( .A(n18578), .ZN(n18496) );
  INV_X1 U12965 ( .A(n18506), .ZN(n18543) );
  INV_X1 U12966 ( .A(n18652), .ZN(n18811) );
  INV_X1 U12967 ( .A(n18760), .ZN(n18672) );
  INV_X1 U12968 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18688) );
  INV_X1 U12969 ( .A(n20927), .ZN(n16472) );
  OR4_X1 U12970 ( .A1(n13064), .A2(n13063), .A3(n13062), .A4(n13061), .ZN(
        P2_U2832) );
  NAND2_X1 U12971 ( .A1(n10073), .A2(n12457), .ZN(P3_U2640) );
  AND2_X4 U12972 ( .A1(n13676), .A2(n10080), .ZN(n12829) );
  AOI22_X1 U12973 ( .A1(n12823), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10084) );
  AOI22_X1 U12974 ( .A1(n12677), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12678), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10083) );
  AND3_X4 U12975 ( .A1(n13968), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n12832) );
  AOI22_X1 U12976 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12832), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10082) );
  AND2_X4 U12977 ( .A1(n13948), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10300) );
  AOI22_X1 U12978 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12686), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10081) );
  AOI22_X1 U12979 ( .A1(n12677), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12678), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10088) );
  AOI22_X1 U12980 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10087) );
  AOI22_X1 U12981 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12832), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10086) );
  AOI22_X1 U12982 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12686), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10085) );
  AOI22_X1 U12983 ( .A1(n12823), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10092) );
  AOI22_X1 U12984 ( .A1(n12677), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12678), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10091) );
  AOI22_X1 U12985 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12832), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10090) );
  AOI22_X1 U12986 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n10089) );
  AOI22_X1 U12987 ( .A1(n12816), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10096) );
  AOI22_X1 U12988 ( .A1(n12677), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12678), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10095) );
  AOI22_X1 U12989 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12832), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10094) );
  AOI22_X1 U12990 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10093) );
  AOI22_X1 U12991 ( .A1(n12832), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10300), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n10101) );
  INV_X2 U12992 ( .A(n10127), .ZN(n12823) );
  AOI22_X1 U12993 ( .A1(n12816), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10100) );
  AOI22_X1 U12994 ( .A1(n12677), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12678), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10099) );
  AOI22_X1 U12995 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n10098) );
  NAND4_X1 U12996 ( .A1(n10101), .A2(n10100), .A3(n10099), .A4(n10098), .ZN(
        n10168) );
  AOI22_X1 U12997 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10105) );
  AOI22_X1 U12998 ( .A1(n12677), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12678), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10104) );
  AOI22_X1 U12999 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12832), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10103) );
  AOI22_X1 U13000 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10102) );
  NAND4_X1 U13001 ( .A1(n10105), .A2(n10104), .A3(n10103), .A4(n10102), .ZN(
        n10167) );
  NAND2_X1 U13002 ( .A1(n10167), .A2(n16304), .ZN(n10106) );
  AOI22_X1 U13003 ( .A1(n12816), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10111) );
  AOI22_X1 U13004 ( .A1(n12677), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12678), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10110) );
  AOI22_X1 U13005 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10109) );
  AOI22_X1 U13006 ( .A1(n12832), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n10300), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10108) );
  AOI22_X1 U13007 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12832), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10116) );
  AOI22_X1 U13008 ( .A1(n12823), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10114) );
  AOI22_X1 U13009 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10113) );
  AND4_X2 U13010 ( .A1(n10448), .A2(n14059), .A3(n12860), .A4(n10185), .ZN(
        n10849) );
  INV_X1 U13011 ( .A(n10849), .ZN(n10853) );
  INV_X1 U13012 ( .A(n12847), .ZN(n10895) );
  AOI22_X1 U13013 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10122) );
  AOI22_X1 U13014 ( .A1(n9598), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12678), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10121) );
  AOI22_X1 U13015 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12832), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10120) );
  AOI22_X1 U13016 ( .A1(n12831), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10119) );
  AOI22_X1 U13017 ( .A1(n12816), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10125) );
  AOI22_X1 U13018 ( .A1(n12831), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10124) );
  AOI22_X1 U13019 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12832), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10123) );
  NAND2_X1 U13020 ( .A1(n10895), .A2(n10885), .ZN(n10851) );
  INV_X1 U13021 ( .A(n10851), .ZN(n10126) );
  INV_X2 U13022 ( .A(n10127), .ZN(n12816) );
  AOI22_X1 U13023 ( .A1(n12823), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10131) );
  AOI22_X1 U13024 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10130) );
  AOI22_X1 U13025 ( .A1(n12832), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10300), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10129) );
  NAND4_X1 U13026 ( .A1(n10132), .A2(n10131), .A3(n10130), .A4(n10129), .ZN(
        n10138) );
  AOI22_X1 U13027 ( .A1(n12677), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12678), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10136) );
  AOI22_X1 U13028 ( .A1(n12823), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10135) );
  AOI22_X1 U13029 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12832), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10134) );
  AOI22_X1 U13030 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10133) );
  NAND4_X1 U13031 ( .A1(n10136), .A2(n10135), .A3(n10134), .A4(n10133), .ZN(
        n10137) );
  MUX2_X2 U13032 ( .A(n10138), .B(n10137), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n19823) );
  NAND2_X1 U13033 ( .A1(n10215), .A2(n10664), .ZN(n10166) );
  AOI22_X1 U13034 ( .A1(n9598), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12678), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10142) );
  AOI22_X1 U13035 ( .A1(n12823), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10141) );
  AOI22_X1 U13036 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12832), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10140) );
  AOI22_X1 U13037 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10139) );
  NAND4_X1 U13038 ( .A1(n10142), .A2(n10141), .A3(n10140), .A4(n10139), .ZN(
        n10143) );
  AOI22_X1 U13039 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12832), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10147) );
  AOI22_X1 U13040 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10146) );
  AOI22_X1 U13041 ( .A1(n12677), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12678), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10145) );
  AOI22_X1 U13042 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10144) );
  NAND4_X1 U13043 ( .A1(n10147), .A2(n10146), .A3(n10145), .A4(n10144), .ZN(
        n10148) );
  INV_X2 U13044 ( .A(n14014), .ZN(n10212) );
  AOI22_X1 U13045 ( .A1(n12677), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12678), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10152) );
  AOI22_X1 U13046 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10151) );
  AOI22_X1 U13047 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12832), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10150) );
  AOI22_X1 U13048 ( .A1(n10300), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10149) );
  AOI22_X1 U13049 ( .A1(n12677), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12678), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10154) );
  AOI22_X1 U13050 ( .A1(n12831), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12817), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10157) );
  AOI22_X1 U13051 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12832), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10156) );
  AOI22_X1 U13052 ( .A1(n12816), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10155) );
  NAND4_X1 U13053 ( .A1(n10158), .A2(n10157), .A3(n10156), .A4(n10155), .ZN(
        n10159) );
  NAND2_X2 U13054 ( .A1(n10160), .A2(n10159), .ZN(n10184) );
  OAI211_X1 U13055 ( .C1(n12847), .C2(n10212), .A(n10184), .B(n10667), .ZN(
        n10165) );
  INV_X2 U13056 ( .A(n10184), .ZN(n10845) );
  NAND4_X1 U13057 ( .A1(n10212), .A2(n14046), .A3(n14059), .A4(n10845), .ZN(
        n10162) );
  NOR2_X2 U13058 ( .A1(n10162), .A2(n10667), .ZN(n10183) );
  INV_X1 U13059 ( .A(n10183), .ZN(n10163) );
  NAND2_X1 U13060 ( .A1(n10166), .A2(n10856), .ZN(n10213) );
  NOR2_X1 U13061 ( .A1(n12847), .A2(n14059), .ZN(n10674) );
  INV_X1 U13062 ( .A(n10674), .ZN(n10211) );
  NAND3_X1 U13063 ( .A1(n10668), .A2(n14059), .A3(n10667), .ZN(n10671) );
  INV_X1 U13064 ( .A(n10167), .ZN(n10171) );
  INV_X1 U13065 ( .A(n10168), .ZN(n10169) );
  OR2_X1 U13066 ( .A1(n10175), .A2(n10169), .ZN(n10170) );
  OAI21_X1 U13067 ( .B1(n10174), .B2(n10171), .A(n10170), .ZN(n10172) );
  NAND3_X1 U13068 ( .A1(n10211), .A2(n10671), .A3(n10172), .ZN(n10177) );
  NAND3_X1 U13069 ( .A1(n10849), .A2(n10175), .A3(n10174), .ZN(n10176) );
  INV_X1 U13070 ( .A(n10662), .ZN(n10180) );
  NAND3_X1 U13071 ( .A1(n19810), .A2(n10184), .A3(n10173), .ZN(n10179) );
  NAND2_X1 U13072 ( .A1(n10180), .A2(n10179), .ZN(n11083) );
  INV_X1 U13073 ( .A(n11083), .ZN(n10181) );
  NAND2_X1 U13074 ( .A1(n10181), .A2(n19830), .ZN(n10219) );
  NAND2_X1 U13075 ( .A1(n10182), .A2(n10219), .ZN(n10231) );
  NAND2_X1 U13076 ( .A1(n10231), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10189) );
  NAND2_X2 U13077 ( .A1(n10183), .A2(n10664), .ZN(n10673) );
  AND3_X1 U13078 ( .A1(n10448), .A2(n10885), .A3(n14046), .ZN(n10877) );
  INV_X1 U13079 ( .A(n10848), .ZN(n10852) );
  NAND4_X1 U13080 ( .A1(n10877), .A2(n10852), .A3(n10664), .A4(n10185), .ZN(
        n10186) );
  NAND2_X1 U13081 ( .A1(n10673), .A2(n10186), .ZN(n10841) );
  NAND2_X1 U13082 ( .A1(n10841), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10195) );
  OAI211_X1 U13083 ( .C1(n19818), .C2(n19793), .A(n10195), .B(n10197), .ZN(
        n10187) );
  INV_X1 U13084 ( .A(n10187), .ZN(n10188) );
  NAND2_X1 U13085 ( .A1(n9723), .A2(n10065), .ZN(n10191) );
  NAND2_X1 U13086 ( .A1(n12847), .A2(n14014), .ZN(n10190) );
  NAND2_X1 U13087 ( .A1(n10191), .A2(n10190), .ZN(n10193) );
  INV_X1 U13088 ( .A(n14059), .ZN(n10663) );
  NAND2_X1 U13089 ( .A1(n10885), .A2(n10664), .ZN(n10847) );
  NAND2_X1 U13090 ( .A1(n10847), .A2(n19809), .ZN(n12844) );
  NAND3_X1 U13091 ( .A1(n10193), .A2(n10192), .A3(n12844), .ZN(n11082) );
  NOR2_X2 U13092 ( .A1(n11082), .A2(n10848), .ZN(n10843) );
  AND2_X2 U13093 ( .A1(n10195), .A2(n10194), .ZN(n10196) );
  NAND2_X2 U13094 ( .A1(n10208), .A2(n10196), .ZN(n10239) );
  NAND2_X1 U13095 ( .A1(n9594), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10202) );
  AND2_X4 U13096 ( .A1(n10198), .A2(n11085), .ZN(n10828) );
  NAND2_X2 U13097 ( .A1(n10199), .A2(n10849), .ZN(n13497) );
  INV_X1 U13099 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n13604) );
  INV_X1 U13100 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13826) );
  AOI21_X1 U13101 ( .B1(n10828), .B2(P2_REIP_REG_1__SCAN_IN), .A(n10200), .ZN(
        n10201) );
  NAND2_X1 U13102 ( .A1(n10204), .A2(n10203), .ZN(n10205) );
  NOR3_X1 U13103 ( .A1(n10848), .A2(n19809), .A3(n19822), .ZN(n10206) );
  INV_X4 U13104 ( .A(n10748), .ZN(n11154) );
  OAI22_X1 U13105 ( .A1(n10231), .A2(n10206), .B1(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n11154), .ZN(n10210) );
  OR2_X1 U13106 ( .A1(n19818), .A2(n19802), .ZN(n10207) );
  AND2_X1 U13107 ( .A1(n10208), .A2(n10207), .ZN(n10209) );
  NAND2_X1 U13108 ( .A1(n10210), .A2(n10209), .ZN(n10246) );
  NAND3_X1 U13109 ( .A1(n10211), .A2(n14046), .A3(n10671), .ZN(n10857) );
  MUX2_X1 U13110 ( .A(n10857), .B(n10853), .S(n10212), .Z(n10214) );
  AOI21_X1 U13111 ( .B1(n10215), .B2(n10214), .A(n10213), .ZN(n10224) );
  INV_X1 U13112 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n10217) );
  NAND2_X1 U13113 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10216) );
  INV_X1 U13114 ( .A(n10218), .ZN(n10221) );
  NAND2_X1 U13115 ( .A1(n10828), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10220) );
  AND3_X1 U13116 ( .A1(n10221), .A2(n10220), .A3(n10219), .ZN(n10223) );
  NAND2_X1 U13117 ( .A1(n10239), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10222) );
  NAND2_X2 U13119 ( .A1(n10246), .A2(n10245), .ZN(n10252) );
  NAND2_X2 U13120 ( .A1(n10251), .A2(n10225), .ZN(n10250) );
  AOI22_X1 U13121 ( .A1(n11154), .A2(P2_EBX_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10226) );
  NAND2_X1 U13122 ( .A1(n10828), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10227) );
  NAND2_X1 U13123 ( .A1(n10231), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10233) );
  AOI21_X1 U13124 ( .B1(n19822), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10232) );
  NAND2_X2 U13125 ( .A1(n10250), .A2(n10248), .ZN(n10238) );
  INV_X1 U13126 ( .A(n10234), .ZN(n10236) );
  NAND2_X1 U13127 ( .A1(n10236), .A2(n10235), .ZN(n10237) );
  BUF_X8 U13128 ( .A(n10239), .Z(n11153) );
  AOI22_X1 U13129 ( .A1(n11154), .A2(P2_EBX_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10241) );
  NAND2_X1 U13130 ( .A1(n10828), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10240) );
  NAND2_X1 U13131 ( .A1(n10241), .A2(n10240), .ZN(n10242) );
  NAND2_X1 U13132 ( .A1(n10231), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10244) );
  OR2_X1 U13133 ( .A1(n19818), .A2(n19775), .ZN(n10243) );
  XNOR2_X2 U13134 ( .A(n10743), .B(n10742), .ZN(n10746) );
  INV_X1 U13135 ( .A(n19019), .ZN(n10247) );
  XNOR2_X2 U13136 ( .A(n10250), .B(n10249), .ZN(n12519) );
  INV_X1 U13137 ( .A(n10252), .ZN(n10254) );
  NAND2_X1 U13138 ( .A1(n10254), .A2(n10256), .ZN(n10255) );
  INV_X1 U13139 ( .A(n13963), .ZN(n15666) );
  INV_X1 U13140 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12612) );
  NOR2_X1 U13141 ( .A1(n14185), .A2(n12612), .ZN(n10264) );
  INV_X1 U13142 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10262) );
  AND2_X1 U13143 ( .A1(n10286), .A2(n10276), .ZN(n10257) );
  NAND2_X1 U13144 ( .A1(n13670), .A2(n10257), .ZN(n19351) );
  INV_X1 U13145 ( .A(n10251), .ZN(n10259) );
  AND2_X1 U13146 ( .A1(n10286), .A2(n10282), .ZN(n10260) );
  NAND2_X1 U13147 ( .A1(n13670), .A2(n10260), .ZN(n13864) );
  INV_X1 U13148 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10261) );
  OAI22_X1 U13149 ( .A1(n10262), .A2(n19351), .B1(n13864), .B2(n10261), .ZN(
        n10263) );
  NOR2_X1 U13150 ( .A1(n10264), .A2(n10263), .ZN(n10266) );
  AOI22_X1 U13151 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n14019), .B1(
        n19491), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10265) );
  NAND2_X1 U13152 ( .A1(n10266), .A2(n10265), .ZN(n10275) );
  NOR2_X1 U13153 ( .A1(n13963), .A2(n19019), .ZN(n10278) );
  AND2_X1 U13154 ( .A1(n13963), .A2(n10247), .ZN(n10283) );
  AOI22_X1 U13155 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19433), .B1(
        n19460), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10273) );
  INV_X1 U13156 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10268) );
  INV_X1 U13157 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10269) );
  NOR2_X1 U13158 ( .A1(n19564), .A2(n10269), .ZN(n10270) );
  NAND2_X1 U13159 ( .A1(n10273), .A2(n10272), .ZN(n10274) );
  NOR2_X1 U13160 ( .A1(n10275), .A2(n10274), .ZN(n10292) );
  AOI21_X1 U13161 ( .B1(n10371), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n12780), .ZN(n10281) );
  AND2_X1 U13162 ( .A1(n12519), .A2(n10276), .ZN(n10277) );
  NAND2_X1 U13163 ( .A1(n13670), .A2(n10277), .ZN(n19222) );
  INV_X1 U13164 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12613) );
  OR2_X1 U13165 ( .A1(n19222), .A2(n12613), .ZN(n10280) );
  INV_X1 U13166 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10279) );
  AOI22_X1 U13167 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n14040), .B1(
        n14102), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10289) );
  NAND2_X1 U13168 ( .A1(n19309), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10288) );
  NAND2_X1 U13169 ( .A1(n19197), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n10287) );
  NAND2_X1 U13170 ( .A1(n10292), .A2(n10291), .ZN(n10334) );
  AND2_X2 U13171 ( .A1(n9598), .A2(n16304), .ZN(n12546) );
  AOI22_X1 U13172 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n12546), .B1(
        n10320), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10297) );
  AND2_X2 U13173 ( .A1(n9601), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10933) );
  AOI22_X1 U13174 ( .A1(n10933), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12551), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10296) );
  AOI22_X1 U13175 ( .A1(n10934), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12545), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10295) );
  CLKBUF_X3 U13176 ( .A(n12699), .Z(n12830) );
  AND2_X2 U13177 ( .A1(n12830), .A2(n16304), .ZN(n12541) );
  AOI22_X1 U13178 ( .A1(n12541), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10294) );
  NAND4_X1 U13179 ( .A1(n10297), .A2(n10296), .A3(n10295), .A4(n10294), .ZN(
        n10308) );
  AND2_X2 U13180 ( .A1(n12816), .A2(n16304), .ZN(n12540) );
  AOI22_X1 U13181 ( .A1(n12540), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12660), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10306) );
  AND2_X2 U13182 ( .A1(n12686), .A2(n16304), .ZN(n12670) );
  NAND2_X1 U13183 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n12679) );
  NOR2_X1 U13184 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n12679), .ZN(
        n10298) );
  NAND2_X1 U13185 ( .A1(n10298), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10339) );
  INV_X1 U13186 ( .A(n10339), .ZN(n10299) );
  AOI22_X1 U13187 ( .A1(n12670), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n10299), .ZN(n10305) );
  NAND3_X1 U13188 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10685) );
  INV_X1 U13189 ( .A(n10685), .ZN(n10301) );
  NAND2_X1 U13190 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10301), .ZN(
        n10340) );
  INV_X1 U13191 ( .A(n10340), .ZN(n10302) );
  AOI22_X1 U13192 ( .A1(n12631), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n10302), .ZN(n10304) );
  AOI22_X1 U13193 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n12552), .B1(
        n12665), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10303) );
  NAND4_X1 U13194 ( .A1(n10306), .A2(n10305), .A3(n10304), .A4(n10303), .ZN(
        n10307) );
  NOR2_X1 U13195 ( .A1(n10308), .A2(n10307), .ZN(n10894) );
  AOI22_X1 U13196 ( .A1(n10933), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10934), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10312) );
  AOI22_X1 U13197 ( .A1(n12540), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12541), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10311) );
  AOI22_X1 U13198 ( .A1(n12551), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10310) );
  AOI22_X1 U13199 ( .A1(n12545), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12546), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10309) );
  NAND4_X1 U13200 ( .A1(n10312), .A2(n10311), .A3(n10310), .A4(n10309), .ZN(
        n10319) );
  AOI22_X1 U13201 ( .A1(n12670), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10317) );
  AOI22_X1 U13202 ( .A1(n12631), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12665), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10316) );
  INV_X1 U13203 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n14085) );
  INV_X1 U13204 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n13296) );
  OAI22_X1 U13205 ( .A1(n10339), .A2(n14085), .B1(n10340), .B2(n13296), .ZN(
        n10313) );
  AOI21_X1 U13206 ( .B1(n10320), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A(
        n10313), .ZN(n10315) );
  NAND2_X1 U13207 ( .A1(n12660), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10314) );
  NAND4_X1 U13208 ( .A1(n10317), .A2(n10316), .A3(n10315), .A4(n10314), .ZN(
        n10318) );
  NAND2_X1 U13209 ( .A1(n10884), .A2(n12780), .ZN(n13234) );
  OR2_X1 U13210 ( .A1(n10894), .A2(n13234), .ZN(n10703) );
  AOI22_X1 U13211 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10320), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10326) );
  AOI22_X1 U13212 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n12665), .B1(
        n12631), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10325) );
  INV_X1 U13213 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10321) );
  INV_X1 U13214 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12520) );
  OAI22_X1 U13215 ( .A1(n10339), .A2(n10321), .B1(n12520), .B2(n10340), .ZN(
        n10322) );
  AOI21_X1 U13216 ( .B1(n12670), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A(
        n10322), .ZN(n10324) );
  NAND2_X1 U13217 ( .A1(n12545), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(
        n10323) );
  NAND4_X1 U13218 ( .A1(n10326), .A2(n10325), .A3(n10324), .A4(n10323), .ZN(
        n10332) );
  AOI22_X1 U13219 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12541), .B1(
        n10934), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10330) );
  AOI22_X1 U13220 ( .A1(n10933), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10329) );
  AOI22_X1 U13221 ( .A1(n12540), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12551), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10328) );
  AOI22_X1 U13222 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12660), .B1(
        n12546), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10327) );
  NAND4_X1 U13223 ( .A1(n10330), .A2(n10329), .A3(n10328), .A4(n10327), .ZN(
        n10331) );
  INV_X1 U13224 ( .A(n10902), .ZN(n10704) );
  NAND2_X1 U13225 ( .A1(n10703), .A2(n10704), .ZN(n10333) );
  AOI22_X1 U13226 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n12540), .B1(
        n10933), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10338) );
  AOI22_X1 U13227 ( .A1(n10934), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10337) );
  AOI22_X1 U13228 ( .A1(n12541), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12551), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10336) );
  AOI22_X1 U13229 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12546), .B1(
        n12545), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10335) );
  NAND4_X1 U13230 ( .A1(n10338), .A2(n10337), .A3(n10336), .A4(n10335), .ZN(
        n10347) );
  AOI22_X1 U13231 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n10320), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10345) );
  AOI22_X1 U13232 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n12665), .B1(
        n12631), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10344) );
  INV_X1 U13233 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11000) );
  OAI22_X1 U13234 ( .A1(n12650), .A2(n19661), .B1(n11000), .B2(n12666), .ZN(
        n10341) );
  AOI21_X1 U13235 ( .B1(n12670), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A(
        n10341), .ZN(n10343) );
  NAND2_X1 U13236 ( .A1(n12660), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10342) );
  NAND4_X1 U13237 ( .A1(n10345), .A2(n10344), .A3(n10343), .A4(n10342), .ZN(
        n10346) );
  AOI22_X1 U13238 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12541), .B1(
        n12540), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10351) );
  AOI22_X1 U13239 ( .A1(n10933), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10350) );
  AOI22_X1 U13240 ( .A1(n10934), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12551), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10349) );
  AOI22_X1 U13241 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12660), .B1(
        n12545), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10348) );
  NAND4_X1 U13242 ( .A1(n10351), .A2(n10350), .A3(n10349), .A4(n10348), .ZN(
        n10360) );
  AOI22_X1 U13243 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10320), .B1(
        n12631), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10358) );
  AOI22_X1 U13244 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12665), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10357) );
  INV_X1 U13245 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10353) );
  INV_X1 U13246 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n10352) );
  OAI22_X1 U13247 ( .A1(n12650), .A2(n10353), .B1(n10352), .B2(n10340), .ZN(
        n10354) );
  AOI21_X1 U13248 ( .B1(n12670), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A(
        n10354), .ZN(n10356) );
  NAND2_X1 U13249 ( .A1(n12546), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10355) );
  NAND4_X1 U13250 ( .A1(n10358), .A2(n10357), .A3(n10356), .A4(n10355), .ZN(
        n10359) );
  AND2_X1 U13251 ( .A1(n10462), .A2(n10702), .ZN(n10361) );
  AOI22_X1 U13252 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19570), .B1(
        n19524), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10367) );
  INV_X1 U13253 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12538) );
  INV_X1 U13254 ( .A(n14102), .ZN(n14105) );
  INV_X1 U13255 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12549) );
  OAI22_X1 U13256 ( .A1(n12538), .A2(n10363), .B1(n14105), .B2(n12549), .ZN(
        n10364) );
  NAND2_X1 U13257 ( .A1(n19309), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10366) );
  NAND2_X1 U13258 ( .A1(n19197), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n10365) );
  INV_X1 U13259 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12547) );
  INV_X1 U13260 ( .A(n19460), .ZN(n19465) );
  INV_X1 U13261 ( .A(n14040), .ZN(n10368) );
  INV_X1 U13262 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14056) );
  OAI22_X1 U13263 ( .A1(n12547), .A2(n19465), .B1(n10368), .B2(n14056), .ZN(
        n10369) );
  INV_X1 U13264 ( .A(n10369), .ZN(n10377) );
  AOI22_X1 U13265 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n14019), .B1(
        n19433), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n10376) );
  INV_X1 U13266 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12559) );
  INV_X1 U13267 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12561) );
  OAI22_X1 U13268 ( .A1(n12559), .A2(n14185), .B1(n19380), .B2(n12561), .ZN(
        n10370) );
  INV_X1 U13269 ( .A(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12560) );
  INV_X1 U13270 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12543) );
  INV_X1 U13271 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10372) );
  INV_X1 U13272 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13871) );
  OAI22_X1 U13273 ( .A1(n10372), .A2(n19351), .B1(n13864), .B2(n13871), .ZN(
        n10373) );
  NOR2_X1 U13274 ( .A1(n10374), .A2(n10373), .ZN(n10375) );
  AOI22_X1 U13275 ( .A1(n10933), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12541), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10381) );
  AOI22_X1 U13276 ( .A1(n10934), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10380) );
  AOI22_X1 U13277 ( .A1(n12540), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12551), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10379) );
  AOI22_X1 U13278 ( .A1(n12546), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12660), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10378) );
  NAND4_X1 U13279 ( .A1(n10381), .A2(n10380), .A3(n10379), .A4(n10378), .ZN(
        n10388) );
  AOI22_X1 U13280 ( .A1(n10320), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12670), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10386) );
  AOI22_X1 U13281 ( .A1(n12631), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12665), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10385) );
  INV_X1 U13282 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13501) );
  OAI22_X1 U13283 ( .A1(n12650), .A2(n14056), .B1(n12666), .B2(n13501), .ZN(
        n10382) );
  AOI21_X1 U13284 ( .B1(n12626), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A(
        n10382), .ZN(n10384) );
  NAND2_X1 U13285 ( .A1(n12545), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n10383) );
  NAND4_X1 U13286 ( .A1(n10386), .A2(n10385), .A3(n10384), .A4(n10383), .ZN(
        n10387) );
  INV_X1 U13287 ( .A(n10922), .ZN(n10389) );
  NAND2_X1 U13288 ( .A1(n10389), .A2(n12780), .ZN(n10390) );
  AOI22_X1 U13289 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19570), .B1(
        n19460), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10399) );
  AOI22_X1 U13290 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19433), .B1(
        n19491), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10398) );
  INV_X1 U13291 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12630) );
  INV_X1 U13292 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10391) );
  OAI22_X1 U13293 ( .A1(n12630), .A2(n19351), .B1(n19277), .B2(n10391), .ZN(
        n10394) );
  INV_X1 U13294 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12636) );
  INV_X1 U13295 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10392) );
  OAI22_X1 U13296 ( .A1(n12636), .A2(n19222), .B1(n13864), .B2(n10392), .ZN(
        n10393) );
  NOR2_X1 U13297 ( .A1(n10394), .A2(n10393), .ZN(n10397) );
  INV_X1 U13298 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n14192) );
  INV_X1 U13299 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12639) );
  OAI22_X1 U13300 ( .A1(n14192), .A2(n14185), .B1(n19380), .B2(n12639), .ZN(
        n10395) );
  INV_X1 U13301 ( .A(n10395), .ZN(n10396) );
  NAND4_X1 U13302 ( .A1(n10399), .A2(n10398), .A3(n10397), .A4(n10396), .ZN(
        n10405) );
  AOI22_X1 U13303 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n14102), .B1(
        n19524), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10403) );
  AOI22_X1 U13304 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n14040), .B1(
        n14019), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10402) );
  NAND2_X1 U13305 ( .A1(n19309), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n10401) );
  NAND2_X1 U13306 ( .A1(n19197), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n10400) );
  NAND4_X1 U13307 ( .A1(n10403), .A2(n10402), .A3(n10401), .A4(n10400), .ZN(
        n10404) );
  INV_X1 U13308 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10406) );
  INV_X1 U13309 ( .A(n10933), .ZN(n12539) );
  INV_X1 U13310 ( .A(n10934), .ZN(n12537) );
  INV_X1 U13311 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12627) );
  OAI22_X1 U13312 ( .A1(n10406), .A2(n12539), .B1(n12537), .B2(n12627), .ZN(
        n10407) );
  INV_X1 U13313 ( .A(n10407), .ZN(n10411) );
  AOI22_X1 U13314 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12541), .B1(
        n12540), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10410) );
  AOI22_X1 U13315 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n12551), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10409) );
  AOI22_X1 U13316 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n12546), .B1(
        n12545), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10408) );
  NAND4_X1 U13317 ( .A1(n10411), .A2(n10410), .A3(n10409), .A4(n10408), .ZN(
        n10419) );
  AOI22_X1 U13318 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12670), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10417) );
  AOI22_X1 U13319 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n12665), .B1(
        n12631), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10416) );
  INV_X1 U13320 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10412) );
  INV_X1 U13321 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11030) );
  OAI22_X1 U13322 ( .A1(n12650), .A2(n10412), .B1(n11030), .B2(n12666), .ZN(
        n10413) );
  AOI21_X1 U13323 ( .B1(n10320), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        n10413), .ZN(n10415) );
  NAND2_X1 U13324 ( .A1(n12660), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n10414) );
  NAND4_X1 U13325 ( .A1(n10417), .A2(n10416), .A3(n10415), .A4(n10414), .ZN(
        n10418) );
  INV_X1 U13326 ( .A(n10929), .ZN(n10420) );
  NAND2_X1 U13327 ( .A1(n10420), .A2(n12780), .ZN(n10421) );
  XNOR2_X2 U13328 ( .A(n10726), .B(n10423), .ZN(n10720) );
  NAND2_X1 U13329 ( .A1(n10933), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10427) );
  NAND2_X1 U13330 ( .A1(n12540), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10426) );
  NAND2_X1 U13331 ( .A1(n10934), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10425) );
  NAND2_X1 U13332 ( .A1(n12631), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10424) );
  NAND2_X1 U13333 ( .A1(n12541), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10431) );
  NAND2_X1 U13334 ( .A1(n12551), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10430) );
  NAND2_X1 U13335 ( .A1(n12545), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10429) );
  NAND2_X1 U13336 ( .A1(n12660), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10428) );
  INV_X1 U13337 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n14051) );
  INV_X1 U13338 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11045) );
  OAI22_X1 U13339 ( .A1(n12650), .A2(n14051), .B1(n11045), .B2(n12666), .ZN(
        n10432) );
  AOI21_X1 U13340 ( .B1(n12670), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A(
        n10432), .ZN(n10434) );
  NAND2_X1 U13341 ( .A1(n12546), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10433) );
  NAND2_X1 U13342 ( .A1(n12552), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10438) );
  NAND2_X1 U13343 ( .A1(n10320), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10437) );
  NAND2_X1 U13344 ( .A1(n12626), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10436) );
  NAND2_X1 U13345 ( .A1(n12665), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10435) );
  NAND2_X1 U13346 ( .A1(n10720), .A2(n10733), .ZN(n10467) );
  XNOR2_X1 U13347 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10647) );
  NAND2_X1 U13348 ( .A1(n19802), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10642) );
  INV_X1 U13349 ( .A(n10642), .ZN(n10443) );
  NAND2_X1 U13350 ( .A1(n10647), .A2(n10443), .ZN(n10445) );
  NAND2_X1 U13351 ( .A1(n19793), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10444) );
  NAND2_X1 U13352 ( .A1(n10445), .A2(n10444), .ZN(n10453) );
  MUX2_X1 U13353 ( .A(n19784), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n10446) );
  XNOR2_X1 U13354 ( .A(n10453), .B(n10446), .ZN(n10659) );
  INV_X1 U13355 ( .A(n10448), .ZN(n10886) );
  NAND2_X1 U13356 ( .A1(n10217), .A2(n13604), .ZN(n10451) );
  MUX2_X1 U13357 ( .A(n10894), .B(n10451), .S(n12848), .Z(n10495) );
  NOR2_X1 U13358 ( .A1(n19809), .A2(n12848), .ZN(n10490) );
  INV_X1 U13359 ( .A(n10702), .ZN(n10911) );
  NAND2_X1 U13360 ( .A1(n10490), .A2(n10911), .ZN(n10460) );
  AND2_X1 U13361 ( .A1(n10886), .A2(n19809), .ZN(n10491) );
  NOR2_X1 U13362 ( .A1(n16301), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10452) );
  NAND2_X1 U13363 ( .A1(n16301), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n10454) );
  MUX2_X1 U13364 ( .A(n19775), .B(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        n16304), .Z(n10456) );
  OR2_X1 U13365 ( .A1(n9669), .A2(n10461), .ZN(n10650) );
  NAND2_X1 U13366 ( .A1(n10491), .A2(n10650), .ZN(n10459) );
  INV_X4 U13367 ( .A(n10886), .ZN(n12848) );
  NAND2_X1 U13368 ( .A1(n12848), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n10458) );
  NAND2_X1 U13369 ( .A1(n10486), .A2(n10484), .ZN(n10500) );
  NAND2_X1 U13370 ( .A1(n10651), .A2(n10491), .ZN(n10464) );
  AOI22_X1 U13371 ( .A1(n10490), .A2(n10918), .B1(n12848), .B2(
        P2_EBX_REG_4__SCAN_IN), .ZN(n10463) );
  NAND2_X1 U13372 ( .A1(n10464), .A2(n10463), .ZN(n10499) );
  NOR2_X2 U13373 ( .A1(n10500), .A2(n10499), .ZN(n10469) );
  INV_X1 U13374 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n10755) );
  MUX2_X1 U13375 ( .A(n10922), .B(n10755), .S(n12848), .Z(n10468) );
  INV_X1 U13376 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13509) );
  MUX2_X1 U13377 ( .A(n10929), .B(n13509), .S(n12848), .Z(n10465) );
  OR2_X1 U13378 ( .A1(n10471), .A2(n10465), .ZN(n10466) );
  NAND2_X1 U13379 ( .A1(n10505), .A2(n10466), .ZN(n13760) );
  INV_X1 U13380 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14173) );
  NOR2_X1 U13381 ( .A1(n10469), .A2(n10468), .ZN(n10470) );
  OR2_X1 U13382 ( .A1(n10471), .A2(n10470), .ZN(n18985) );
  OAI21_X1 U13383 ( .B1(n10718), .B2(n11182), .A(n18985), .ZN(n10472) );
  INV_X1 U13384 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14513) );
  AND2_X1 U13385 ( .A1(n10733), .A2(n14513), .ZN(n10478) );
  INV_X1 U13386 ( .A(n10478), .ZN(n10474) );
  AND2_X1 U13387 ( .A1(n18985), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10479) );
  INV_X1 U13388 ( .A(n10479), .ZN(n10473) );
  MUX2_X1 U13389 ( .A(n10474), .B(n10473), .S(n10477), .Z(n10483) );
  OAI21_X1 U13390 ( .B1(n10733), .B2(n14513), .A(n18985), .ZN(n10476) );
  OAI21_X1 U13391 ( .B1(n18985), .B2(n14513), .A(n10476), .ZN(n10482) );
  MUX2_X1 U13392 ( .A(n10479), .B(n10478), .S(n10477), .Z(n10480) );
  NAND2_X1 U13393 ( .A1(n10480), .A2(n10475), .ZN(n10481) );
  OAI211_X1 U13394 ( .C1(n10483), .C2(n10475), .A(n10482), .B(n10481), .ZN(
        n14504) );
  INV_X1 U13395 ( .A(n10484), .ZN(n10485) );
  XNOR2_X1 U13396 ( .A(n10486), .B(n10485), .ZN(n13771) );
  NOR2_X1 U13397 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13771), .ZN(
        n10498) );
  INV_X1 U13398 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11090) );
  INV_X1 U13399 ( .A(n10486), .ZN(n10489) );
  NAND2_X1 U13400 ( .A1(n10487), .A2(n10495), .ZN(n10488) );
  NAND2_X1 U13401 ( .A1(n10489), .A2(n10488), .ZN(n13689) );
  NOR2_X1 U13402 ( .A1(n11090), .A2(n13689), .ZN(n10497) );
  NAND2_X1 U13403 ( .A1(n10490), .A2(n10884), .ZN(n10493) );
  OAI21_X1 U13404 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19802), .A(
        n10642), .ZN(n10641) );
  INV_X1 U13405 ( .A(n10641), .ZN(n10689) );
  NAND2_X1 U13406 ( .A1(n10491), .A2(n10689), .ZN(n10492) );
  OAI211_X1 U13407 ( .C1(n10217), .C2(n10886), .A(n10493), .B(n10492), .ZN(
        n19021) );
  NAND2_X1 U13408 ( .A1(n19021), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13322) );
  NAND3_X1 U13409 ( .A1(n12848), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n10494) );
  NAND2_X1 U13410 ( .A1(n10495), .A2(n10494), .ZN(n13830) );
  NOR2_X1 U13411 ( .A1(n13322), .A2(n13830), .ZN(n10496) );
  NAND2_X1 U13412 ( .A1(n13322), .A2(n13830), .ZN(n13321) );
  OAI21_X1 U13413 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10496), .A(
        n13321), .ZN(n13339) );
  XOR2_X1 U13414 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n13689), .Z(
        n13338) );
  NOR2_X1 U13415 ( .A1(n13339), .A2(n13338), .ZN(n13337) );
  NOR2_X1 U13416 ( .A1(n10497), .A2(n13337), .ZN(n13704) );
  NAND2_X1 U13417 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13771), .ZN(
        n13703) );
  OAI21_X1 U13418 ( .B1(n10498), .B2(n13704), .A(n13703), .ZN(n19146) );
  XNOR2_X1 U13419 ( .A(n10500), .B(n10499), .ZN(n10501) );
  XNOR2_X1 U13420 ( .A(n10501), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19145) );
  NAND2_X1 U13421 ( .A1(n19146), .A2(n19145), .ZN(n10503) );
  INV_X1 U13422 ( .A(n10501), .ZN(n18998) );
  NAND2_X1 U13423 ( .A1(n18998), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10502) );
  NAND2_X1 U13424 ( .A1(n10503), .A2(n10502), .ZN(n14505) );
  NAND2_X1 U13425 ( .A1(n14504), .A2(n14505), .ZN(n10504) );
  MUX2_X1 U13426 ( .A(n10733), .B(P2_EBX_REG_7__SCAN_IN), .S(n12848), .Z(
        n10509) );
  NAND2_X1 U13427 ( .A1(n10521), .A2(n10507), .ZN(n10508) );
  NAND2_X1 U13428 ( .A1(n10514), .A2(n10508), .ZN(n18965) );
  NOR2_X1 U13429 ( .A1(n18965), .A2(n10733), .ZN(n10516) );
  NAND2_X1 U13430 ( .A1(n10516), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16258) );
  XNOR2_X1 U13431 ( .A(n10505), .B(n10506), .ZN(n18976) );
  NAND2_X1 U13432 ( .A1(n18976), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16255) );
  INV_X1 U13433 ( .A(n18976), .ZN(n10511) );
  NAND2_X1 U13434 ( .A1(n10511), .A2(n14271), .ZN(n16254) );
  NAND2_X1 U13435 ( .A1(n10514), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10512) );
  MUX2_X1 U13436 ( .A(n10512), .B(n10514), .S(n10886), .Z(n10513) );
  INV_X1 U13437 ( .A(n10513), .ZN(n10515) );
  NOR2_X1 U13438 ( .A1(n10515), .A2(n10529), .ZN(n13810) );
  AOI21_X1 U13439 ( .B1(n13810), .B2(n11182), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15387) );
  INV_X1 U13440 ( .A(n15387), .ZN(n10519) );
  INV_X1 U13441 ( .A(n10516), .ZN(n10517) );
  INV_X1 U13442 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10946) );
  INV_X1 U13443 ( .A(n16257), .ZN(n10518) );
  NAND2_X1 U13444 ( .A1(n10519), .A2(n10518), .ZN(n10524) );
  NAND2_X1 U13445 ( .A1(n12848), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10520) );
  MUX2_X1 U13446 ( .A(n10520), .B(P2_EBX_REG_10__SCAN_IN), .S(n10529), .Z(
        n10522) );
  AND2_X1 U13447 ( .A1(n10522), .A2(n10609), .ZN(n18951) );
  AOI21_X1 U13448 ( .B1(n18951), .B2(n11182), .A(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15378) );
  INV_X1 U13449 ( .A(n15378), .ZN(n10523) );
  INV_X1 U13450 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15646) );
  NOR2_X1 U13451 ( .A1(n10733), .A2(n15646), .ZN(n10525) );
  NAND2_X1 U13452 ( .A1(n18951), .A2(n10525), .ZN(n15379) );
  INV_X1 U13453 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n10526) );
  NOR2_X1 U13454 ( .A1(n10733), .A2(n10526), .ZN(n10527) );
  NAND2_X1 U13455 ( .A1(n13810), .A2(n10527), .ZN(n15388) );
  AND2_X1 U13456 ( .A1(n15379), .A2(n15388), .ZN(n10528) );
  INV_X1 U13457 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n13739) );
  INV_X1 U13458 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n13749) );
  NAND2_X2 U13459 ( .A1(n10538), .A2(n10609), .ZN(n10537) );
  INV_X1 U13460 ( .A(n10530), .ZN(n10531) );
  AND3_X1 U13461 ( .A1(n12848), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n10531), .ZN(
        n10532) );
  NOR2_X1 U13462 ( .A1(n10537), .A2(n10532), .ZN(n18941) );
  AND2_X1 U13463 ( .A1(n18941), .A2(n11182), .ZN(n10533) );
  AND2_X1 U13464 ( .A1(n10533), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15635) );
  INV_X1 U13465 ( .A(n10533), .ZN(n10535) );
  INV_X1 U13466 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n10534) );
  NAND2_X1 U13467 ( .A1(n12848), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10536) );
  NAND3_X1 U13468 ( .A1(n12848), .A2(n10538), .A3(P2_EBX_REG_12__SCAN_IN), 
        .ZN(n10539) );
  AND2_X1 U13469 ( .A1(n10541), .A2(n10539), .ZN(n18930) );
  INV_X1 U13470 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15613) );
  NOR2_X1 U13471 ( .A1(n10733), .A2(n15613), .ZN(n10540) );
  NAND2_X1 U13472 ( .A1(n18930), .A2(n10540), .ZN(n15367) );
  NAND2_X1 U13473 ( .A1(n15369), .A2(n15367), .ZN(n15280) );
  AND2_X1 U13474 ( .A1(n12848), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n10543) );
  OAI21_X1 U13475 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(P2_EBX_REG_14__SCAN_IN), 
        .A(n12848), .ZN(n10542) );
  NAND2_X1 U13476 ( .A1(n12848), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10554) );
  OR2_X2 U13477 ( .A1(n10546), .A2(n10545), .ZN(n10548) );
  AOI21_X1 U13478 ( .B1(n10543), .B2(n10548), .A(n10550), .ZN(n15098) );
  INV_X1 U13479 ( .A(n15098), .ZN(n10544) );
  NOR2_X1 U13480 ( .A1(n10733), .A2(n10544), .ZN(n10578) );
  NOR2_X1 U13481 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n10578), .ZN(
        n15305) );
  NAND2_X1 U13482 ( .A1(n10546), .A2(n10545), .ZN(n10547) );
  NAND2_X1 U13483 ( .A1(n10548), .A2(n10547), .ZN(n15107) );
  NOR2_X1 U13484 ( .A1(n10733), .A2(n15107), .ZN(n10579) );
  NOR2_X1 U13485 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n10579), .ZN(
        n15319) );
  NAND2_X1 U13486 ( .A1(n12848), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10549) );
  INV_X1 U13487 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n14384) );
  NAND2_X1 U13488 ( .A1(n10550), .A2(n14384), .ZN(n10552) );
  OAI211_X1 U13489 ( .C1(n10550), .C2(n10549), .A(n10609), .B(n10552), .ZN(
        n18871) );
  OR2_X1 U13490 ( .A1(n18871), .A2(n10733), .ZN(n10584) );
  INV_X1 U13491 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15265) );
  AND2_X1 U13492 ( .A1(n10584), .A2(n15265), .ZN(n11103) );
  OR2_X1 U13493 ( .A1(n15319), .A2(n11103), .ZN(n10551) );
  NOR2_X1 U13494 ( .A1(n15305), .A2(n10551), .ZN(n15294) );
  OR2_X2 U13495 ( .A1(n10552), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10574) );
  INV_X1 U13496 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15501) );
  OAI21_X1 U13497 ( .B1(n18863), .B2(n10733), .A(n15501), .ZN(n15296) );
  INV_X1 U13498 ( .A(n10554), .ZN(n10555) );
  XNOR2_X1 U13499 ( .A(n10556), .B(n10555), .ZN(n18884) );
  NAND2_X1 U13500 ( .A1(n18884), .A2(n11182), .ZN(n10583) );
  INV_X1 U13501 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15549) );
  NAND2_X1 U13502 ( .A1(n10583), .A2(n15549), .ZN(n15332) );
  NAND3_X1 U13503 ( .A1(n10557), .A2(P2_EBX_REG_16__SCAN_IN), .A3(n12848), 
        .ZN(n10558) );
  NAND3_X1 U13504 ( .A1(n10559), .A2(n10609), .A3(n10558), .ZN(n18900) );
  INV_X1 U13505 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15544) );
  OAI21_X1 U13506 ( .B1(n18900), .B2(n10733), .A(n15544), .ZN(n10561) );
  OR2_X1 U13507 ( .A1(n10733), .A2(n15544), .ZN(n10560) );
  NAND2_X1 U13508 ( .A1(n10561), .A2(n15330), .ZN(n15349) );
  INV_X1 U13509 ( .A(n15349), .ZN(n11106) );
  AND2_X1 U13510 ( .A1(n12848), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10563) );
  XNOR2_X1 U13511 ( .A(n10562), .B(n10563), .ZN(n18908) );
  NAND2_X1 U13512 ( .A1(n18908), .A2(n11182), .ZN(n10581) );
  INV_X1 U13513 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15585) );
  NAND2_X1 U13514 ( .A1(n10581), .A2(n15585), .ZN(n15359) );
  INV_X1 U13515 ( .A(n10564), .ZN(n10565) );
  XNOR2_X1 U13516 ( .A(n10541), .B(n10565), .ZN(n18921) );
  NAND2_X1 U13517 ( .A1(n18921), .A2(n11182), .ZN(n10566) );
  INV_X1 U13518 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15596) );
  NAND2_X1 U13519 ( .A1(n10566), .A2(n15596), .ZN(n15598) );
  AND4_X1 U13520 ( .A1(n15332), .A2(n11106), .A3(n15359), .A4(n15598), .ZN(
        n10571) );
  INV_X1 U13521 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n13936) );
  NAND2_X1 U13522 ( .A1(n10562), .A2(n13936), .ZN(n10567) );
  NAND3_X1 U13523 ( .A1(n10567), .A2(P2_EBX_REG_15__SCAN_IN), .A3(n12848), 
        .ZN(n10568) );
  NAND2_X1 U13524 ( .A1(n10568), .A2(n10557), .ZN(n14208) );
  NOR2_X1 U13525 ( .A1(n10733), .A2(n14208), .ZN(n10580) );
  NOR2_X1 U13526 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n10580), .ZN(
        n15564) );
  INV_X1 U13527 ( .A(n15564), .ZN(n10570) );
  INV_X1 U13528 ( .A(n18930), .ZN(n10569) );
  OAI21_X1 U13529 ( .B1(n10569), .B2(n10733), .A(n15613), .ZN(n15368) );
  NAND2_X1 U13530 ( .A1(n12848), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10572) );
  NAND3_X1 U13531 ( .A1(n10574), .A2(P2_EBX_REG_22__SCAN_IN), .A3(n12848), 
        .ZN(n10575) );
  NAND2_X1 U13532 ( .A1(n10593), .A2(n10575), .ZN(n13082) );
  OR2_X1 U13533 ( .A1(n13082), .A2(n10733), .ZN(n10576) );
  INV_X1 U13534 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15493) );
  NAND2_X1 U13535 ( .A1(n10576), .A2(n15493), .ZN(n15284) );
  AND2_X1 U13536 ( .A1(n15279), .A2(n15284), .ZN(n10577) );
  INV_X1 U13537 ( .A(n15284), .ZN(n10590) );
  AND2_X1 U13538 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n10578), .ZN(
        n15306) );
  NAND2_X1 U13539 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n10579), .ZN(
        n15317) );
  AND2_X1 U13540 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n10580), .ZN(
        n15563) );
  NOR2_X1 U13541 ( .A1(n15585), .A2(n10581), .ZN(n15357) );
  NOR2_X1 U13542 ( .A1(n15563), .A2(n15357), .ZN(n11105) );
  NOR2_X1 U13543 ( .A1(n10733), .A2(n15501), .ZN(n10582) );
  NAND2_X1 U13544 ( .A1(n15330), .A2(n9637), .ZN(n11107) );
  INV_X1 U13545 ( .A(n10584), .ZN(n10585) );
  NAND2_X1 U13546 ( .A1(n10585), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11102) );
  NOR2_X1 U13547 ( .A1(n10733), .A2(n15596), .ZN(n10586) );
  NAND2_X1 U13548 ( .A1(n18921), .A2(n10586), .ZN(n15597) );
  NOR2_X1 U13549 ( .A1(n15306), .A2(n10587), .ZN(n15281) );
  OR2_X1 U13550 ( .A1(n10733), .A2(n15493), .ZN(n10588) );
  OR2_X1 U13551 ( .A1(n13082), .A2(n10588), .ZN(n15283) );
  AND2_X1 U13552 ( .A1(n15281), .A2(n15283), .ZN(n10589) );
  OR2_X1 U13553 ( .A1(n10590), .A2(n10589), .ZN(n10591) );
  AND2_X1 U13554 ( .A1(n12848), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10592) );
  OR2_X2 U13555 ( .A1(n10593), .A2(n10592), .ZN(n10598) );
  NAND2_X1 U13556 ( .A1(n10593), .A2(n10592), .ZN(n10594) );
  AND2_X1 U13557 ( .A1(n10598), .A2(n10594), .ZN(n13053) );
  NAND2_X1 U13558 ( .A1(n13053), .A2(n11182), .ZN(n10595) );
  XNOR2_X1 U13559 ( .A(n10595), .B(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n15268) );
  INV_X1 U13560 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15477) );
  NOR2_X1 U13561 ( .A1(n10733), .A2(n15477), .ZN(n10596) );
  NAND2_X1 U13562 ( .A1(n13053), .A2(n10596), .ZN(n10597) );
  NOR2_X2 U13563 ( .A1(n10598), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10608) );
  NAND3_X1 U13564 ( .A1(n10598), .A2(n12848), .A3(P2_EBX_REG_24__SCAN_IN), 
        .ZN(n10599) );
  NAND2_X1 U13565 ( .A1(n10599), .A2(n10609), .ZN(n10600) );
  NOR2_X1 U13566 ( .A1(n10608), .A2(n10600), .ZN(n16202) );
  NAND2_X1 U13567 ( .A1(n16202), .A2(n11182), .ZN(n15256) );
  NAND2_X1 U13568 ( .A1(n10601), .A2(n15256), .ZN(n10603) );
  NAND2_X1 U13569 ( .A1(n12848), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10604) );
  MUX2_X1 U13570 ( .A(n10604), .B(P2_EBX_REG_25__SCAN_IN), .S(n10608), .Z(
        n10605) );
  AND2_X1 U13571 ( .A1(n10605), .A2(n10609), .ZN(n15081) );
  NAND2_X1 U13572 ( .A1(n15081), .A2(n11182), .ZN(n10606) );
  INV_X1 U13573 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15443) );
  NAND2_X1 U13574 ( .A1(n10606), .A2(n15443), .ZN(n15247) );
  INV_X1 U13575 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n10607) );
  NAND2_X1 U13576 ( .A1(n10608), .A2(n10607), .ZN(n10611) );
  NOR2_X2 U13577 ( .A1(n10611), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10618) );
  NAND3_X1 U13578 ( .A1(n12848), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n10611), 
        .ZN(n10612) );
  NAND2_X1 U13579 ( .A1(n11181), .A2(n10612), .ZN(n10614) );
  INV_X1 U13580 ( .A(n10614), .ZN(n16191) );
  INV_X1 U13581 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15434) );
  NOR2_X1 U13582 ( .A1(n10733), .A2(n15434), .ZN(n10613) );
  NAND2_X1 U13583 ( .A1(n16191), .A2(n10613), .ZN(n10623) );
  OAI21_X1 U13584 ( .B1(n10614), .B2(n10733), .A(n15434), .ZN(n10615) );
  NAND2_X1 U13585 ( .A1(n12848), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10617) );
  INV_X1 U13586 ( .A(n10617), .ZN(n10620) );
  INV_X1 U13587 ( .A(n10618), .ZN(n10619) );
  NAND2_X1 U13588 ( .A1(n10620), .A2(n10619), .ZN(n10621) );
  NAND2_X1 U13589 ( .A1(n10629), .A2(n10621), .ZN(n13067) );
  INV_X1 U13590 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15417) );
  NAND2_X1 U13591 ( .A1(n12848), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n10627) );
  XNOR2_X1 U13592 ( .A(n10629), .B(n10627), .ZN(n16178) );
  NAND2_X1 U13593 ( .A1(n16178), .A2(n11182), .ZN(n12461) );
  NOR2_X1 U13594 ( .A1(n10733), .A2(n15443), .ZN(n10622) );
  NAND2_X1 U13595 ( .A1(n15081), .A2(n10622), .ZN(n15246) );
  NAND2_X1 U13596 ( .A1(n15246), .A2(n10623), .ZN(n12458) );
  AOI21_X1 U13597 ( .B1(n10624), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n12458), .ZN(n10625) );
  INV_X1 U13598 ( .A(n10627), .ZN(n10628) );
  NAND2_X1 U13599 ( .A1(n12848), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n10632) );
  XNOR2_X1 U13600 ( .A(n10633), .B(n10632), .ZN(n10631) );
  INV_X1 U13601 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n10630) );
  OAI21_X1 U13602 ( .B1(n10631), .B2(n10733), .A(n10630), .ZN(n15218) );
  NAND2_X1 U13603 ( .A1(n15221), .A2(n15218), .ZN(n11178) );
  INV_X1 U13604 ( .A(n10631), .ZN(n11262) );
  NAND3_X1 U13605 ( .A1(n11262), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n11182), .ZN(n15219) );
  NAND2_X1 U13606 ( .A1(n11178), .A2(n15219), .ZN(n10638) );
  NAND2_X1 U13607 ( .A1(n10633), .A2(n10632), .ZN(n11179) );
  NAND2_X1 U13608 ( .A1(n12848), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10634) );
  XNOR2_X1 U13609 ( .A(n11179), .B(n10634), .ZN(n10635) );
  AOI21_X1 U13610 ( .B1(n10635), .B2(n11182), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11177) );
  INV_X1 U13611 ( .A(n11177), .ZN(n10636) );
  INV_X1 U13612 ( .A(n10635), .ZN(n16170) );
  INV_X1 U13613 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11167) );
  OR3_X1 U13614 ( .A1(n16170), .A2(n10733), .A3(n11167), .ZN(n11176) );
  NAND2_X1 U13615 ( .A1(n10636), .A2(n11176), .ZN(n10637) );
  XNOR2_X1 U13616 ( .A(n10638), .B(n10637), .ZN(n11195) );
  NOR2_X1 U13617 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15807), .ZN(
        n10639) );
  NAND2_X1 U13618 ( .A1(n19829), .A2(n10641), .ZN(n10643) );
  XNOR2_X1 U13619 ( .A(n10647), .B(n10642), .ZN(n10660) );
  NAND2_X1 U13620 ( .A1(n10643), .A2(n10660), .ZN(n10646) );
  INV_X1 U13621 ( .A(n10659), .ZN(n10644) );
  NAND2_X1 U13622 ( .A1(n19829), .A2(n10644), .ZN(n10645) );
  NAND2_X1 U13623 ( .A1(n10646), .A2(n10645), .ZN(n10648) );
  NAND2_X1 U13624 ( .A1(n10647), .A2(n10689), .ZN(n10679) );
  AOI22_X1 U13625 ( .A1(n10648), .A2(n10664), .B1(n11252), .B2(n10679), .ZN(
        n10649) );
  NOR2_X1 U13626 ( .A1(n10684), .A2(n10652), .ZN(n10653) );
  NAND2_X1 U13627 ( .A1(n10684), .A2(n19830), .ZN(n10654) );
  NOR2_X1 U13628 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19691) );
  AOI211_X1 U13629 ( .C1(P2_STATE_REG_1__SCAN_IN), .C2(P2_STATE_REG_2__SCAN_IN), .A(P2_STATE_REG_0__SCAN_IN), .B(n19691), .ZN(n19828) );
  INV_X1 U13630 ( .A(n19828), .ZN(n19687) );
  NAND2_X1 U13631 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19825) );
  INV_X1 U13632 ( .A(n19825), .ZN(n19695) );
  NOR2_X1 U13633 ( .A1(n19687), .A2(n19695), .ZN(n13107) );
  NAND2_X1 U13634 ( .A1(n10845), .A2(n13107), .ZN(n10699) );
  OAI21_X1 U13635 ( .B1(n10655), .B2(n19823), .A(n10663), .ZN(n10656) );
  INV_X1 U13636 ( .A(n10656), .ZN(n10657) );
  NAND2_X1 U13637 ( .A1(n13216), .A2(n10657), .ZN(n10698) );
  INV_X1 U13638 ( .A(n10682), .ZN(n10658) );
  NOR2_X1 U13639 ( .A1(n10659), .A2(n10658), .ZN(n10688) );
  AND2_X1 U13640 ( .A1(n10688), .A2(n10660), .ZN(n10661) );
  NAND2_X1 U13641 ( .A1(n16352), .A2(n13107), .ZN(n10677) );
  NAND2_X1 U13642 ( .A1(n10663), .A2(n12780), .ZN(n10866) );
  NAND2_X1 U13643 ( .A1(n10866), .A2(n10664), .ZN(n10665) );
  NAND2_X1 U13644 ( .A1(n10665), .A2(n14046), .ZN(n10666) );
  NAND2_X1 U13645 ( .A1(n10666), .A2(n10184), .ZN(n10672) );
  NAND2_X1 U13646 ( .A1(n10668), .A2(n10667), .ZN(n10669) );
  NAND2_X1 U13647 ( .A1(n10669), .A2(n14046), .ZN(n10670) );
  AND2_X1 U13648 ( .A1(n12780), .A2(n19823), .ZN(n11256) );
  NAND2_X1 U13649 ( .A1(n10670), .A2(n11256), .ZN(n10858) );
  AND4_X1 U13650 ( .A1(n10672), .A2(n10848), .A3(n10671), .A4(n10858), .ZN(
        n10676) );
  OAI21_X1 U13651 ( .B1(n10674), .B2(n10845), .A(n10673), .ZN(n10675) );
  OAI21_X1 U13652 ( .B1(n16324), .B2(n10677), .A(n10868), .ZN(n13160) );
  MUX2_X1 U13653 ( .A(n16352), .B(n10845), .S(n12780), .Z(n10678) );
  NAND2_X1 U13654 ( .A1(n10678), .A2(n19825), .ZN(n10695) );
  NAND2_X1 U13655 ( .A1(n10680), .A2(n10679), .ZN(n10681) );
  NAND2_X1 U13656 ( .A1(n10682), .A2(n10681), .ZN(n19808) );
  AND2_X1 U13657 ( .A1(n10683), .A2(n11256), .ZN(n10741) );
  INV_X1 U13658 ( .A(n10684), .ZN(n19807) );
  NAND3_X1 U13659 ( .A1(n19808), .A2(n10741), .A3(n19807), .ZN(n10694) );
  NAND2_X1 U13660 ( .A1(n16339), .A2(n10685), .ZN(n13167) );
  OR2_X1 U13661 ( .A1(n12552), .A2(n13167), .ZN(n10687) );
  INV_X1 U13662 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n15806) );
  AND2_X1 U13663 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15806), .ZN(n10686) );
  NAND2_X1 U13664 ( .A1(n10687), .A2(n10686), .ZN(n19798) );
  AOI21_X1 U13665 ( .B1(n10689), .B2(n10688), .A(n16324), .ZN(n10690) );
  INV_X1 U13666 ( .A(n10690), .ZN(n10691) );
  NAND2_X1 U13667 ( .A1(n13937), .A2(n10691), .ZN(n10692) );
  NAND3_X1 U13668 ( .A1(n10683), .A2(n10069), .A3(n11085), .ZN(n10693) );
  OAI21_X1 U13669 ( .B1(n16324), .B2(n10695), .A(n11113), .ZN(n10696) );
  NOR2_X1 U13670 ( .A1(n13160), .A2(n10696), .ZN(n10697) );
  OAI211_X1 U13671 ( .C1(n13216), .C2(n10699), .A(n10698), .B(n10697), .ZN(
        n10701) );
  NAND2_X1 U13672 ( .A1(n13937), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11259) );
  INV_X1 U13673 ( .A(n11259), .ZN(n10700) );
  XOR2_X1 U13674 ( .A(n10704), .B(n10703), .Z(n13342) );
  NAND2_X1 U13675 ( .A1(n13234), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13233) );
  XOR2_X1 U13676 ( .A(n10884), .B(n10894), .Z(n10705) );
  NOR2_X1 U13677 ( .A1(n13233), .A2(n10705), .ZN(n10706) );
  INV_X1 U13678 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13958) );
  XNOR2_X1 U13679 ( .A(n13233), .B(n10705), .ZN(n13325) );
  NOR2_X1 U13680 ( .A1(n13958), .A2(n13325), .ZN(n13324) );
  NOR2_X1 U13681 ( .A1(n10706), .A2(n13324), .ZN(n10707) );
  XOR2_X1 U13682 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n10707), .Z(
        n13341) );
  NOR2_X1 U13683 ( .A1(n13342), .A2(n13341), .ZN(n13340) );
  NOR2_X1 U13684 ( .A1(n10707), .A2(n11090), .ZN(n10708) );
  INV_X1 U13685 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n16299) );
  XNOR2_X1 U13686 ( .A(n10709), .B(n16299), .ZN(n13699) );
  NAND2_X1 U13687 ( .A1(n10709), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10710) );
  OAI21_X1 U13688 ( .B1(n10711), .B2(n10911), .A(n10918), .ZN(n10713) );
  NAND2_X1 U13689 ( .A1(n10713), .A2(n10712), .ZN(n19142) );
  NAND2_X1 U13690 ( .A1(n10714), .A2(n19142), .ZN(n10717) );
  INV_X1 U13691 ( .A(n19144), .ZN(n10715) );
  NAND2_X1 U13692 ( .A1(n10715), .A2(n19161), .ZN(n10716) );
  NAND2_X1 U13693 ( .A1(n10718), .A2(n14513), .ZN(n14499) );
  INV_X1 U13694 ( .A(n10718), .ZN(n10719) );
  NAND2_X1 U13695 ( .A1(n10719), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14500) );
  INV_X1 U13696 ( .A(n14500), .ZN(n14502) );
  NAND2_X1 U13697 ( .A1(n14502), .A2(n10727), .ZN(n10724) );
  XNOR2_X1 U13698 ( .A(n10734), .B(n10733), .ZN(n10729) );
  NAND2_X1 U13699 ( .A1(n14265), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15392) );
  INV_X1 U13700 ( .A(n10729), .ZN(n10730) );
  NAND2_X1 U13701 ( .A1(n10731), .A2(n10730), .ZN(n15391) );
  OR2_X1 U13702 ( .A1(n10733), .A2(n10946), .ZN(n10732) );
  NOR2_X1 U13703 ( .A1(n15613), .A2(n15596), .ZN(n15587) );
  INV_X1 U13704 ( .A(n15587), .ZN(n11093) );
  NOR2_X1 U13705 ( .A1(n11093), .A2(n15585), .ZN(n10738) );
  AND2_X1 U13706 ( .A1(n10738), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10739) );
  AND2_X1 U13707 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n10739), .ZN(
        n15355) );
  AND2_X1 U13708 ( .A1(n15355), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15345) );
  NAND2_X1 U13709 ( .A1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11139) );
  INV_X1 U13710 ( .A(n11139), .ZN(n15475) );
  NAND4_X1 U13711 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A4(n15475), .ZN(n11089) );
  INV_X1 U13712 ( .A(n11089), .ZN(n10740) );
  INV_X1 U13713 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15461) );
  NAND3_X1 U13714 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11168) );
  XNOR2_X1 U13715 ( .A(n15216), .B(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11196) );
  INV_X1 U13716 ( .A(n10741), .ZN(n19806) );
  INV_X1 U13717 ( .A(n10742), .ZN(n10744) );
  AND2_X1 U13718 ( .A1(n10744), .A2(n10743), .ZN(n10745) );
  NAND2_X1 U13719 ( .A1(n11153), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10753) );
  INV_X1 U13720 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n10750) );
  INV_X1 U13721 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n10749) );
  OAI22_X1 U13722 ( .A1(n10826), .A2(n10750), .B1(n13937), .B2(n10749), .ZN(
        n10751) );
  AOI21_X1 U13723 ( .B1(n10828), .B2(P2_REIP_REG_4__SCAN_IN), .A(n10751), .ZN(
        n10752) );
  NAND2_X1 U13724 ( .A1(n10753), .A2(n10752), .ZN(n13598) );
  NAND2_X1 U13725 ( .A1(n11153), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10758) );
  INV_X1 U13726 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10754) );
  OAI22_X1 U13727 ( .A1(n10826), .A2(n10755), .B1(n13937), .B2(n10754), .ZN(
        n10756) );
  AOI21_X1 U13728 ( .B1(n10828), .B2(P2_REIP_REG_5__SCAN_IN), .A(n10756), .ZN(
        n10757) );
  NAND2_X1 U13729 ( .A1(n10758), .A2(n10757), .ZN(n13606) );
  NAND2_X1 U13730 ( .A1(n13607), .A2(n13606), .ZN(n13609) );
  AOI22_X1 U13731 ( .A1(n11154), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10760) );
  NAND2_X1 U13732 ( .A1(n10828), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n10759) );
  NAND2_X1 U13733 ( .A1(n10760), .A2(n10759), .ZN(n10761) );
  AOI21_X1 U13734 ( .B1(n11153), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n10761), .ZN(n13505) );
  AOI22_X1 U13735 ( .A1(n11154), .A2(P2_EBX_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10765) );
  NAND2_X1 U13736 ( .A1(n10828), .A2(P2_REIP_REG_7__SCAN_IN), .ZN(n10764) );
  NAND2_X1 U13737 ( .A1(n10765), .A2(n10764), .ZN(n10766) );
  AOI21_X1 U13738 ( .B1(n11153), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n10766), .ZN(n13587) );
  AOI22_X1 U13739 ( .A1(n11154), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10768) );
  NAND2_X1 U13740 ( .A1(n10828), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10767) );
  NAND2_X1 U13741 ( .A1(n10768), .A2(n10767), .ZN(n10769) );
  AOI21_X1 U13742 ( .B1(n11153), .B2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(
        n10769), .ZN(n13648) );
  NAND2_X1 U13743 ( .A1(n11153), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10772) );
  INV_X1 U13744 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n13806) );
  OAI22_X1 U13745 ( .A1(n10826), .A2(n9877), .B1(n13937), .B2(n13806), .ZN(
        n10770) );
  AOI21_X1 U13746 ( .B1(n10828), .B2(P2_REIP_REG_9__SCAN_IN), .A(n10770), .ZN(
        n10771) );
  NAND2_X1 U13747 ( .A1(n10772), .A2(n10771), .ZN(n13656) );
  AOI22_X1 U13748 ( .A1(n11154), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n10774) );
  NAND2_X1 U13749 ( .A1(n10828), .A2(P2_REIP_REG_10__SCAN_IN), .ZN(n10773) );
  NAND2_X1 U13750 ( .A1(n10774), .A2(n10773), .ZN(n10775) );
  AOI21_X1 U13751 ( .B1(n11153), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n10775), .ZN(n13734) );
  NAND2_X1 U13752 ( .A1(n11153), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10779) );
  INV_X1 U13753 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10776) );
  OAI22_X1 U13754 ( .A1(n10826), .A2(n13749), .B1(n13937), .B2(n10776), .ZN(
        n10777) );
  AOI21_X1 U13755 ( .B1(n10828), .B2(P2_REIP_REG_11__SCAN_IN), .A(n10777), 
        .ZN(n10778) );
  NAND2_X1 U13756 ( .A1(n10779), .A2(n10778), .ZN(n13747) );
  INV_X1 U13757 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n11008) );
  NAND2_X1 U13758 ( .A1(n11154), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10781) );
  NAND2_X1 U13759 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10780) );
  OAI211_X1 U13760 ( .C1(n11157), .C2(n11008), .A(n10781), .B(n10780), .ZN(
        n10782) );
  AOI21_X1 U13761 ( .B1(n11153), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n10782), .ZN(n13818) );
  INV_X1 U13762 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n11011) );
  NAND2_X1 U13763 ( .A1(n11154), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10784) );
  NAND2_X1 U13764 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10783) );
  OAI211_X1 U13765 ( .C1(n11157), .C2(n11011), .A(n10784), .B(n10783), .ZN(
        n10785) );
  AOI21_X1 U13766 ( .B1(n11153), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n10785), .ZN(n13889) );
  INV_X1 U13767 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n10788) );
  NAND2_X1 U13768 ( .A1(n11154), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10787) );
  NAND2_X1 U13769 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10786) );
  OAI211_X1 U13770 ( .C1(n11157), .C2(n10788), .A(n10787), .B(n10786), .ZN(
        n10789) );
  AOI21_X1 U13771 ( .B1(n11153), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n10789), .ZN(n13933) );
  NAND2_X1 U13772 ( .A1(n11153), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10793) );
  INV_X1 U13773 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n10790) );
  OAI22_X1 U13774 ( .A1(n10826), .A2(n10790), .B1(n13937), .B2(n16238), .ZN(
        n10791) );
  AOI21_X1 U13775 ( .B1(n10828), .B2(P2_REIP_REG_15__SCAN_IN), .A(n10791), 
        .ZN(n10792) );
  NAND2_X1 U13776 ( .A1(n10793), .A2(n10792), .ZN(n14030) );
  INV_X1 U13777 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n15350) );
  NAND2_X1 U13778 ( .A1(n11154), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10795) );
  NAND2_X1 U13779 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10794) );
  OAI211_X1 U13780 ( .C1(n11157), .C2(n15350), .A(n10795), .B(n10794), .ZN(
        n10796) );
  AOI21_X1 U13781 ( .B1(n11153), .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n10796), .ZN(n14089) );
  INV_X1 U13782 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19727) );
  NAND2_X1 U13783 ( .A1(n11154), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10798) );
  NAND2_X1 U13784 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10797) );
  OAI211_X1 U13785 ( .C1(n11157), .C2(n19727), .A(n10798), .B(n10797), .ZN(
        n10799) );
  AOI21_X1 U13786 ( .B1(n11153), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n10799), .ZN(n14234) );
  NAND2_X1 U13787 ( .A1(n11153), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10803) );
  INV_X1 U13788 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n10800) );
  INV_X1 U13789 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15324) );
  OAI22_X1 U13790 ( .A1(n10826), .A2(n10800), .B1(n13937), .B2(n15324), .ZN(
        n10801) );
  AOI21_X1 U13791 ( .B1(n10828), .B2(P2_REIP_REG_18__SCAN_IN), .A(n10801), 
        .ZN(n10802) );
  NAND2_X1 U13792 ( .A1(n10803), .A2(n10802), .ZN(n14243) );
  NAND2_X1 U13793 ( .A1(n14244), .A2(n14243), .ZN(n14242) );
  INV_X1 U13794 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n15090) );
  NAND2_X1 U13795 ( .A1(n11154), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n10805) );
  NAND2_X1 U13796 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n10804) );
  OAI211_X1 U13797 ( .C1(n11157), .C2(n15090), .A(n10805), .B(n10804), .ZN(
        n10806) );
  AOI21_X1 U13798 ( .B1(n11153), .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A(
        n10806), .ZN(n14308) );
  INV_X1 U13799 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n11122) );
  NAND2_X1 U13800 ( .A1(n11154), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10808) );
  NAND2_X1 U13801 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10807) );
  OAI211_X1 U13802 ( .C1(n11157), .C2(n11122), .A(n10808), .B(n10807), .ZN(
        n10809) );
  AOI21_X1 U13803 ( .B1(n11153), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n10809), .ZN(n11118) );
  NAND2_X1 U13804 ( .A1(n11153), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10813) );
  INV_X1 U13805 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n10810) );
  INV_X1 U13806 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n18858) );
  OAI22_X1 U13807 ( .A1(n10826), .A2(n10810), .B1(n13937), .B2(n18858), .ZN(
        n10811) );
  AOI21_X1 U13808 ( .B1(n10828), .B2(P2_REIP_REG_21__SCAN_IN), .A(n10811), 
        .ZN(n10812) );
  NAND2_X1 U13809 ( .A1(n10813), .A2(n10812), .ZN(n15166) );
  INV_X1 U13810 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19735) );
  NAND2_X1 U13811 ( .A1(n11153), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10815) );
  AOI22_X1 U13812 ( .A1(n11154), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n10814) );
  OAI211_X1 U13813 ( .C1(n11157), .C2(n19735), .A(n10815), .B(n10814), .ZN(
        n13084) );
  INV_X1 U13814 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19737) );
  NAND2_X1 U13815 ( .A1(n11154), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10817) );
  NAND2_X1 U13816 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n10816) );
  OAI211_X1 U13817 ( .C1(n11157), .C2(n19737), .A(n10817), .B(n10816), .ZN(
        n10818) );
  AOI21_X1 U13818 ( .B1(n11153), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n10818), .ZN(n13057) );
  INV_X1 U13819 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19739) );
  NAND2_X1 U13820 ( .A1(n11154), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10820) );
  NAND2_X1 U13821 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10819) );
  OAI211_X1 U13822 ( .C1(n11157), .C2(n19739), .A(n10820), .B(n10819), .ZN(
        n10821) );
  AOI21_X1 U13823 ( .B1(n11153), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n10821), .ZN(n15151) );
  NAND2_X1 U13824 ( .A1(n11153), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10824) );
  INV_X1 U13825 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15251) );
  OAI22_X1 U13826 ( .A1(n10826), .A2(n10607), .B1(n13937), .B2(n15251), .ZN(
        n10822) );
  AOI21_X1 U13827 ( .B1(n10828), .B2(P2_REIP_REG_25__SCAN_IN), .A(n10822), 
        .ZN(n10823) );
  NAND2_X1 U13828 ( .A1(n10824), .A2(n10823), .ZN(n15076) );
  NAND2_X1 U13829 ( .A1(n11153), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10830) );
  INV_X1 U13830 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n15140) );
  INV_X1 U13831 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10825) );
  OAI22_X1 U13832 ( .A1(n10826), .A2(n15140), .B1(n13937), .B2(n10825), .ZN(
        n10827) );
  AOI21_X1 U13833 ( .B1(n10828), .B2(P2_REIP_REG_26__SCAN_IN), .A(n10827), 
        .ZN(n10829) );
  NAND2_X1 U13834 ( .A1(n10830), .A2(n10829), .ZN(n15135) );
  INV_X1 U13835 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19746) );
  NAND2_X1 U13836 ( .A1(n11154), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10832) );
  NAND2_X1 U13837 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n10831) );
  OAI211_X1 U13838 ( .C1(n11157), .C2(n19746), .A(n10832), .B(n10831), .ZN(
        n10833) );
  AOI21_X1 U13839 ( .B1(n11153), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n10833), .ZN(n13071) );
  INV_X1 U13840 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n12467) );
  NAND2_X1 U13841 ( .A1(n11154), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n10835) );
  NAND2_X1 U13842 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n10834) );
  OAI211_X1 U13843 ( .C1(n11157), .C2(n12467), .A(n10835), .B(n10834), .ZN(
        n10836) );
  AOI21_X1 U13844 ( .B1(n11153), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n10836), .ZN(n12464) );
  INV_X1 U13845 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19748) );
  NAND2_X1 U13846 ( .A1(n11153), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10838) );
  AOI22_X1 U13847 ( .A1(n11154), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n10837) );
  OAI211_X1 U13848 ( .C1(n11157), .C2(n19748), .A(n10838), .B(n10837), .ZN(
        n11251) );
  NAND2_X1 U13849 ( .A1(n12466), .A2(n11251), .ZN(n11250) );
  INV_X1 U13850 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n19752) );
  AOI22_X1 U13851 ( .A1(n11154), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n10839) );
  OAI21_X1 U13852 ( .B1(n11157), .B2(n19752), .A(n10839), .ZN(n10840) );
  AOI21_X1 U13853 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n11153), .A(
        n10840), .ZN(n11151) );
  INV_X1 U13854 ( .A(n10841), .ZN(n10842) );
  NAND2_X1 U13855 ( .A1(n16352), .A2(n19823), .ZN(n11263) );
  NAND2_X1 U13856 ( .A1(n10842), .A2(n11263), .ZN(n13967) );
  AOI21_X1 U13857 ( .B1(n12780), .B2(n13967), .A(n10843), .ZN(n10844) );
  INV_X1 U13858 ( .A(n12844), .ZN(n13106) );
  NAND2_X1 U13859 ( .A1(n10848), .A2(n14059), .ZN(n10846) );
  AOI22_X1 U13860 ( .A1(n13106), .A2(n10846), .B1(n10845), .B2(n19823), .ZN(
        n10855) );
  NOR2_X1 U13861 ( .A1(n10848), .A2(n10847), .ZN(n10850) );
  NAND2_X1 U13862 ( .A1(n10850), .A2(n10849), .ZN(n12842) );
  NAND3_X1 U13863 ( .A1(n10853), .A2(n10852), .A3(n10851), .ZN(n10854) );
  AND4_X1 U13864 ( .A1(n10856), .A2(n10855), .A3(n12842), .A4(n10854), .ZN(
        n10861) );
  NAND2_X1 U13865 ( .A1(n10857), .A2(n10173), .ZN(n13939) );
  NAND2_X1 U13866 ( .A1(n13939), .A2(n10858), .ZN(n10859) );
  NAND2_X1 U13867 ( .A1(n10859), .A2(n14014), .ZN(n10860) );
  NAND2_X1 U13868 ( .A1(n10861), .A2(n10860), .ZN(n13962) );
  INV_X1 U13869 ( .A(n13497), .ZN(n13671) );
  NOR2_X1 U13870 ( .A1(n13962), .A2(n13671), .ZN(n10862) );
  NAND2_X1 U13871 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n19191) );
  INV_X1 U13872 ( .A(n19191), .ZN(n10863) );
  OR2_X1 U13873 ( .A1(n15537), .A2(n10863), .ZN(n10865) );
  INV_X1 U13874 ( .A(n19818), .ZN(n10864) );
  NAND2_X2 U13875 ( .A1(n10864), .A2(n19764), .ZN(n19155) );
  INV_X1 U13876 ( .A(n19155), .ZN(n18902) );
  NAND2_X1 U13877 ( .A1(n11088), .A2(n19155), .ZN(n13227) );
  NAND2_X1 U13878 ( .A1(n10865), .A2(n13227), .ZN(n19182) );
  INV_X1 U13879 ( .A(n10866), .ZN(n10867) );
  NAND2_X1 U13880 ( .A1(n10868), .A2(n10867), .ZN(n16325) );
  NAND3_X1 U13881 ( .A1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10874) );
  NAND2_X1 U13882 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15630) );
  NAND2_X1 U13883 ( .A1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n14506) );
  NAND2_X1 U13884 ( .A1(n11090), .A2(n19191), .ZN(n19169) );
  INV_X1 U13885 ( .A(n15537), .ZN(n10869) );
  NAND2_X1 U13886 ( .A1(n10869), .A2(n11090), .ZN(n19192) );
  OAI211_X1 U13887 ( .C1(n19169), .C2(n19175), .A(n10870), .B(n19192), .ZN(
        n10871) );
  NOR2_X1 U13888 ( .A1(n16299), .A2(n10871), .ZN(n16300) );
  INV_X1 U13889 ( .A(n15534), .ZN(n15626) );
  OR2_X1 U13890 ( .A1(n16300), .A2(n15626), .ZN(n19164) );
  INV_X1 U13891 ( .A(n19164), .ZN(n10872) );
  AOI21_X1 U13892 ( .B1(n14506), .B2(n15534), .A(n10872), .ZN(n14268) );
  NAND2_X1 U13893 ( .A1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16282) );
  OAI21_X1 U13894 ( .B1(n16282), .B2(n14173), .A(n15534), .ZN(n10873) );
  NAND3_X1 U13895 ( .A1(n14268), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(
        n10873), .ZN(n15625) );
  NOR2_X1 U13896 ( .A1(n15630), .A2(n15625), .ZN(n15610) );
  NAND3_X1 U13897 ( .A1(n15610), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n15587), .ZN(n15535) );
  NOR2_X1 U13898 ( .A1(n10874), .A2(n15535), .ZN(n15527) );
  NAND2_X1 U13899 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15527), .ZN(
        n11135) );
  NOR2_X1 U13900 ( .A1(n11089), .A2(n11135), .ZN(n15428) );
  NAND2_X1 U13901 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15429) );
  OR2_X1 U13902 ( .A1(n15461), .A2(n15429), .ZN(n11095) );
  INV_X1 U13903 ( .A(n11095), .ZN(n10875) );
  NAND2_X1 U13904 ( .A1(n15428), .A2(n10875), .ZN(n10876) );
  AND2_X1 U13905 ( .A1(n15534), .A2(n10876), .ZN(n12479) );
  AOI21_X1 U13906 ( .B1(n11168), .B2(n15534), .A(n12479), .ZN(n11170) );
  AOI222_X1 U13907 ( .A1(n11078), .A2(P2_REIP_REG_30__SCAN_IN), .B1(n11160), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .C1(n11161), .C2(
        P2_EAX_REG_30__SCAN_IN), .ZN(n11081) );
  NOR2_X1 U13908 ( .A1(n11164), .A2(n15090), .ZN(n10879) );
  INV_X1 U13909 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15513) );
  INV_X1 U13910 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n14219) );
  OAI22_X1 U13911 ( .A1(n15513), .A2(n10891), .B1(n11059), .B2(n14219), .ZN(
        n10878) );
  OR2_X1 U13912 ( .A1(n10879), .A2(n10878), .ZN(n14218) );
  INV_X1 U13913 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18850) );
  INV_X1 U13914 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13938) );
  NAND2_X1 U13915 ( .A1(n12860), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n10880) );
  OAI211_X1 U13916 ( .C1(n12780), .C2(n13938), .A(n10880), .B(n19794), .ZN(
        n10881) );
  INV_X1 U13917 ( .A(n10881), .ZN(n10882) );
  OAI21_X1 U13918 ( .B1(n11164), .B2(n18850), .A(n10882), .ZN(n13229) );
  NAND2_X1 U13919 ( .A1(n11160), .A2(n12847), .ZN(n10904) );
  NAND2_X1 U13920 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10883) );
  AND2_X1 U13921 ( .A1(n11059), .A2(n10883), .ZN(n10890) );
  AND2_X1 U13922 ( .A1(n10885), .A2(n19794), .ZN(n10887) );
  NAND2_X1 U13923 ( .A1(n10884), .A2(n10888), .ZN(n10889) );
  NAND3_X1 U13924 ( .A1(n10904), .A2(n10890), .A3(n10889), .ZN(n13228) );
  INV_X1 U13925 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19702) );
  NOR2_X1 U13926 ( .A1(n11164), .A2(n19702), .ZN(n10893) );
  INV_X1 U13927 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19137) );
  OAI22_X1 U13928 ( .A1(n13958), .A2(n10891), .B1(n11059), .B2(n19137), .ZN(
        n10892) );
  XNOR2_X1 U13929 ( .A(n13231), .B(n10899), .ZN(n13531) );
  OR2_X1 U13930 ( .A1(n10894), .A2(n11039), .ZN(n10898) );
  NAND2_X1 U13931 ( .A1(n10895), .A2(n14046), .ZN(n10896) );
  MUX2_X1 U13932 ( .A(n10896), .B(n19793), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n10897) );
  NAND2_X1 U13933 ( .A1(n10898), .A2(n10897), .ZN(n13530) );
  NOR2_X1 U13934 ( .A1(n13531), .A2(n13530), .ZN(n10901) );
  NOR2_X1 U13935 ( .A1(n13231), .A2(n10899), .ZN(n10900) );
  NAND2_X1 U13936 ( .A1(n10888), .A2(n10902), .ZN(n10903) );
  OAI211_X1 U13937 ( .C1(n19794), .C2(n19784), .A(n10904), .B(n10903), .ZN(
        n10907) );
  XNOR2_X1 U13938 ( .A(n10908), .B(n10907), .ZN(n13523) );
  INV_X1 U13939 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19704) );
  NOR2_X1 U13940 ( .A1(n11164), .A2(n19704), .ZN(n10906) );
  INV_X1 U13941 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n19135) );
  OAI22_X1 U13942 ( .A1(n11090), .A2(n10891), .B1(n11059), .B2(n19135), .ZN(
        n10905) );
  OR2_X1 U13943 ( .A1(n10906), .A2(n10905), .ZN(n13522) );
  NOR2_X1 U13944 ( .A1(n13523), .A2(n13522), .ZN(n13524) );
  NOR2_X1 U13945 ( .A1(n10908), .A2(n10907), .ZN(n10909) );
  INV_X1 U13946 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n13701) );
  INV_X1 U13947 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n10910) );
  OAI22_X1 U13948 ( .A1(n11039), .A2(n10911), .B1(n11059), .B2(n10910), .ZN(
        n10912) );
  INV_X1 U13949 ( .A(n10912), .ZN(n10915) );
  OAI22_X1 U13950 ( .A1(n10891), .A2(n16299), .B1(n19775), .B2(n19794), .ZN(
        n10913) );
  INV_X1 U13951 ( .A(n10913), .ZN(n10914) );
  OAI211_X1 U13952 ( .C1(n13701), .C2(n11164), .A(n10915), .B(n10914), .ZN(
        n13768) );
  NAND2_X1 U13953 ( .A1(n11161), .A2(P2_EAX_REG_4__SCAN_IN), .ZN(n10917) );
  INV_X1 U13954 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n19161) );
  OR2_X1 U13955 ( .A1(n10891), .A2(n19161), .ZN(n10916) );
  OAI211_X1 U13956 ( .C1(n10918), .C2(n11039), .A(n10917), .B(n10916), .ZN(
        n10919) );
  INV_X1 U13957 ( .A(n10919), .ZN(n10921) );
  NAND2_X1 U13958 ( .A1(n11078), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n10920) );
  AOI22_X1 U13959 ( .A1(n11078), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n11160), 
        .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n10924) );
  AOI22_X1 U13960 ( .A1(n10888), .A2(n10922), .B1(n11161), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n10923) );
  NAND2_X1 U13961 ( .A1(n10924), .A2(n10923), .ZN(n14508) );
  INV_X1 U13962 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19710) );
  NOR2_X1 U13963 ( .A1(n11164), .A2(n19710), .ZN(n10926) );
  INV_X1 U13964 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19128) );
  OAI22_X1 U13965 ( .A1(n10891), .A2(n14173), .B1(n11059), .B2(n19128), .ZN(
        n10925) );
  AND2_X1 U13966 ( .A1(n14508), .A2(n10928), .ZN(n10927) );
  INV_X1 U13967 ( .A(n10928), .ZN(n13755) );
  NAND2_X1 U13968 ( .A1(n10888), .A2(n10929), .ZN(n13754) );
  OR2_X1 U13969 ( .A1(n13755), .A2(n13754), .ZN(n10931) );
  NAND2_X1 U13970 ( .A1(n10888), .A2(n11182), .ZN(n10930) );
  AOI22_X1 U13971 ( .A1(n10933), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12540), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10938) );
  AOI22_X1 U13972 ( .A1(n10934), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12541), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10937) );
  AOI22_X1 U13973 ( .A1(n12551), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10936) );
  AOI22_X1 U13974 ( .A1(n12545), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12660), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10935) );
  NAND4_X1 U13975 ( .A1(n10938), .A2(n10937), .A3(n10936), .A4(n10935), .ZN(
        n10945) );
  AOI22_X1 U13976 ( .A1(n10320), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12670), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10943) );
  AOI22_X1 U13977 ( .A1(n12631), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12665), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10942) );
  INV_X1 U13978 ( .A(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12649) );
  OAI22_X1 U13979 ( .A1(n12650), .A2(n13296), .B1(n12666), .B2(n12649), .ZN(
        n10939) );
  AOI21_X1 U13980 ( .B1(n12626), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A(
        n10939), .ZN(n10941) );
  NAND2_X1 U13981 ( .A1(n12546), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10940) );
  NAND4_X1 U13982 ( .A1(n10943), .A2(n10942), .A3(n10941), .A4(n10940), .ZN(
        n10944) );
  NOR2_X1 U13983 ( .A1(n10945), .A2(n10944), .ZN(n13651) );
  NAND2_X1 U13984 ( .A1(n11161), .A2(P2_EAX_REG_8__SCAN_IN), .ZN(n10948) );
  OR2_X1 U13985 ( .A1(n10891), .A2(n10946), .ZN(n10947) );
  OAI211_X1 U13986 ( .C1(n13651), .C2(n11039), .A(n10948), .B(n10947), .ZN(
        n10949) );
  INV_X1 U13987 ( .A(n10949), .ZN(n10951) );
  NAND2_X1 U13988 ( .A1(n11078), .A2(P2_REIP_REG_8__SCAN_IN), .ZN(n10950) );
  INV_X1 U13989 ( .A(n16277), .ZN(n10954) );
  INV_X1 U13990 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19712) );
  NOR2_X1 U13991 ( .A1(n11164), .A2(n19712), .ZN(n10953) );
  INV_X1 U13992 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n14271) );
  INV_X1 U13993 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19125) );
  OAI22_X1 U13994 ( .A1(n14271), .A2(n10891), .B1(n11059), .B2(n19125), .ZN(
        n10952) );
  OR2_X1 U13995 ( .A1(n10953), .A2(n10952), .ZN(n14274) );
  AND2_X1 U13996 ( .A1(n10954), .A2(n14274), .ZN(n10955) );
  AOI22_X1 U13997 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n10933), .B1(
        n10934), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10959) );
  AOI22_X1 U13998 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n12540), .B1(
        n12541), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10958) );
  AOI22_X1 U13999 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n12551), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10957) );
  AOI22_X1 U14000 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n12545), .B1(
        n12546), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10956) );
  NAND4_X1 U14001 ( .A1(n10959), .A2(n10958), .A3(n10957), .A4(n10956), .ZN(
        n10966) );
  AOI22_X1 U14002 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12670), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10964) );
  AOI22_X1 U14003 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12665), .B1(
        n12631), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10963) );
  INV_X1 U14004 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12507) );
  OAI22_X1 U14005 ( .A1(n10339), .A2(n12507), .B1(n12613), .B2(n12666), .ZN(
        n10960) );
  AOI21_X1 U14006 ( .B1(n10320), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n10960), .ZN(n10962) );
  NAND2_X1 U14007 ( .A1(n12660), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10961) );
  NAND4_X1 U14008 ( .A1(n10964), .A2(n10963), .A3(n10962), .A4(n10961), .ZN(
        n10965) );
  AOI22_X1 U14009 ( .A1(n11078), .A2(P2_REIP_REG_9__SCAN_IN), .B1(n10888), 
        .B2(n13655), .ZN(n10968) );
  AOI22_X1 U14010 ( .A1(n11160), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B1(
        n11161), .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n10967) );
  NAND2_X1 U14011 ( .A1(n10968), .A2(n10967), .ZN(n13803) );
  AOI22_X1 U14012 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n12540), .B1(
        n10933), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10972) );
  AOI22_X1 U14013 ( .A1(n12541), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12631), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10971) );
  AOI22_X1 U14014 ( .A1(n10934), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12551), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10970) );
  AOI22_X1 U14015 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12660), .B1(
        n12546), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10969) );
  NAND4_X1 U14016 ( .A1(n10972), .A2(n10971), .A3(n10970), .A4(n10969), .ZN(
        n10979) );
  AOI22_X1 U14017 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10320), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10977) );
  AOI22_X1 U14018 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12665), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10976) );
  INV_X1 U14019 ( .A(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12599) );
  OAI22_X1 U14020 ( .A1(n12650), .A2(n12520), .B1(n12599), .B2(n12666), .ZN(
        n10973) );
  AOI21_X1 U14021 ( .B1(n12670), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n10973), .ZN(n10975) );
  NAND2_X1 U14022 ( .A1(n12545), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n10974) );
  NAND4_X1 U14023 ( .A1(n10977), .A2(n10976), .A3(n10975), .A4(n10974), .ZN(
        n10978) );
  INV_X1 U14024 ( .A(n12531), .ZN(n13730) );
  NOR2_X1 U14025 ( .A1(n11039), .A2(n13730), .ZN(n10982) );
  INV_X1 U14026 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n10980) );
  OAI22_X1 U14027 ( .A1(n10891), .A2(n15646), .B1(n11059), .B2(n10980), .ZN(
        n10981) );
  AOI211_X1 U14028 ( .C1(P2_REIP_REG_10__SCAN_IN), .C2(n11078), .A(n10982), 
        .B(n10981), .ZN(n15641) );
  AOI22_X1 U14029 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n10933), .B1(
        n10934), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10986) );
  AOI22_X1 U14030 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n12540), .B1(
        n12541), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10985) );
  AOI22_X1 U14031 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n12551), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10984) );
  AOI22_X1 U14032 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n12545), .B1(
        n12546), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10983) );
  NAND4_X1 U14033 ( .A1(n10986), .A2(n10985), .A3(n10984), .A4(n10983), .ZN(
        n10993) );
  AOI22_X1 U14034 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12670), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10991) );
  AOI22_X1 U14035 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12665), .B1(
        n12631), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10990) );
  INV_X1 U14036 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12586) );
  OAI22_X1 U14037 ( .A1(n12650), .A2(n10352), .B1(n12586), .B2(n12666), .ZN(
        n10987) );
  AOI21_X1 U14038 ( .B1(n10320), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n10987), .ZN(n10989) );
  NAND2_X1 U14039 ( .A1(n12660), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n10988) );
  NAND4_X1 U14040 ( .A1(n10991), .A2(n10990), .A3(n10989), .A4(n10988), .ZN(
        n10992) );
  AOI22_X1 U14041 ( .A1(n11078), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n10888), 
        .B2(n13813), .ZN(n10995) );
  AOI22_X1 U14042 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n11160), .B1(
        n11161), .B2(P2_EAX_REG_11__SCAN_IN), .ZN(n10994) );
  NAND2_X1 U14043 ( .A1(n10995), .A2(n10994), .ZN(n15628) );
  AOI22_X1 U14044 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n10933), .B1(
        n10934), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10999) );
  AOI22_X1 U14045 ( .A1(n12540), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n12631), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10998) );
  AOI22_X1 U14046 ( .A1(n12541), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12551), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10997) );
  AOI22_X1 U14047 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12545), .B1(
        n12546), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10996) );
  NAND4_X1 U14048 ( .A1(n10999), .A2(n10998), .A3(n10997), .A4(n10996), .ZN(
        n11007) );
  AOI22_X1 U14049 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10320), .B1(
        n12665), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11005) );
  AOI22_X1 U14050 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n12552), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11004) );
  INV_X1 U14051 ( .A(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12573) );
  OAI22_X1 U14052 ( .A1(n12650), .A2(n11000), .B1(n12573), .B2(n12666), .ZN(
        n11001) );
  AOI21_X1 U14053 ( .B1(n12670), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A(
        n11001), .ZN(n11003) );
  NAND2_X1 U14054 ( .A1(n12660), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11002) );
  NAND4_X1 U14055 ( .A1(n11005), .A2(n11004), .A3(n11003), .A4(n11002), .ZN(
        n11006) );
  OR2_X1 U14056 ( .A1(n11007), .A2(n11006), .ZN(n13815) );
  INV_X1 U14057 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n13132) );
  OAI22_X1 U14058 ( .A1(n15613), .A2(n10891), .B1(n11059), .B2(n13132), .ZN(
        n11010) );
  NOR2_X1 U14059 ( .A1(n11164), .A2(n11008), .ZN(n11009) );
  AOI211_X1 U14060 ( .C1(n10888), .C2(n13815), .A(n11010), .B(n11009), .ZN(
        n15616) );
  OAI22_X1 U14061 ( .A1(n11164), .A2(n11011), .B1(n15596), .B2(n10891), .ZN(
        n11012) );
  INV_X1 U14062 ( .A(n11012), .ZN(n11025) );
  AOI22_X1 U14063 ( .A1(n10933), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n10934), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11016) );
  AOI22_X1 U14064 ( .A1(n12540), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12541), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11015) );
  AOI22_X1 U14065 ( .A1(n12551), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11014) );
  AOI22_X1 U14066 ( .A1(n12545), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12546), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11013) );
  NAND4_X1 U14067 ( .A1(n11016), .A2(n11015), .A3(n11014), .A4(n11013), .ZN(
        n11023) );
  AOI22_X1 U14068 ( .A1(n12670), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11021) );
  AOI22_X1 U14069 ( .A1(n12631), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12665), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11020) );
  OAI22_X1 U14070 ( .A1(n12650), .A2(n13501), .B1(n12666), .B2(n12560), .ZN(
        n11017) );
  AOI21_X1 U14071 ( .B1(n10320), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A(
        n11017), .ZN(n11019) );
  NAND2_X1 U14072 ( .A1(n12660), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11018) );
  NAND4_X1 U14073 ( .A1(n11021), .A2(n11020), .A3(n11019), .A4(n11018), .ZN(
        n11022) );
  OR2_X1 U14074 ( .A1(n11023), .A2(n11022), .ZN(n12534) );
  AOI22_X1 U14075 ( .A1(n10888), .A2(n12534), .B1(n11161), .B2(
        P2_EAX_REG_13__SCAN_IN), .ZN(n11024) );
  NAND2_X1 U14076 ( .A1(n11025), .A2(n11024), .ZN(n15602) );
  AOI22_X1 U14077 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n10934), .B1(
        n10933), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11029) );
  AOI22_X1 U14078 ( .A1(n12541), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12631), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11028) );
  AOI22_X1 U14079 ( .A1(n12540), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12551), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11027) );
  AOI22_X1 U14080 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n12660), .B1(
        n12545), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11026) );
  NAND4_X1 U14081 ( .A1(n11029), .A2(n11028), .A3(n11027), .A4(n11026), .ZN(
        n11037) );
  AOI22_X1 U14082 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n12552), .B1(
        n12665), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11035) );
  AOI22_X1 U14083 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10320), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11034) );
  OAI22_X1 U14084 ( .A1(n12650), .A2(n11030), .B1(n12636), .B2(n12666), .ZN(
        n11031) );
  AOI21_X1 U14085 ( .B1(n12670), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n11031), .ZN(n11033) );
  NAND2_X1 U14086 ( .A1(n12546), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11032) );
  NAND4_X1 U14087 ( .A1(n11035), .A2(n11034), .A3(n11033), .A4(n11032), .ZN(
        n11036) );
  NOR2_X1 U14088 ( .A1(n11037), .A2(n11036), .ZN(n13928) );
  AOI22_X1 U14089 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n11160), .B1(
        n11161), .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n11038) );
  OAI21_X1 U14090 ( .B1(n13928), .B2(n11039), .A(n11038), .ZN(n11040) );
  AOI21_X1 U14091 ( .B1(P2_REIP_REG_14__SCAN_IN), .B2(n11078), .A(n11040), 
        .ZN(n15582) );
  AOI22_X1 U14092 ( .A1(n11078), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n11160), .ZN(n11054) );
  AOI22_X1 U14093 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n10934), .B1(
        n10933), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11044) );
  AOI22_X1 U14094 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n12540), .B1(
        n12541), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11043) );
  AOI22_X1 U14095 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n12551), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11042) );
  AOI22_X1 U14096 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n12546), .B1(
        n12545), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11041) );
  NAND4_X1 U14097 ( .A1(n11044), .A2(n11043), .A3(n11042), .A4(n11041), .ZN(
        n11052) );
  AOI22_X1 U14098 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12670), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11050) );
  AOI22_X1 U14099 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n12665), .B1(
        n12631), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11049) );
  INV_X1 U14100 ( .A(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12668) );
  OAI22_X1 U14101 ( .A1(n12650), .A2(n11045), .B1(n12668), .B2(n12666), .ZN(
        n11046) );
  AOI21_X1 U14102 ( .B1(n10320), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A(
        n11046), .ZN(n11048) );
  NAND2_X1 U14103 ( .A1(n12660), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11047) );
  NAND4_X1 U14104 ( .A1(n11050), .A2(n11049), .A3(n11048), .A4(n11047), .ZN(
        n11051) );
  NOR2_X1 U14105 ( .A1(n11052), .A2(n11051), .ZN(n14029) );
  AOI22_X1 U14106 ( .A1(n10888), .A2(n9848), .B1(n11161), .B2(
        P2_EAX_REG_15__SCAN_IN), .ZN(n11053) );
  NAND2_X1 U14107 ( .A1(n11054), .A2(n11053), .ZN(n14199) );
  NAND2_X1 U14108 ( .A1(n11078), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11058) );
  INV_X1 U14109 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n11055) );
  OAI22_X1 U14110 ( .A1(n15544), .A2(n10891), .B1(n11059), .B2(n11055), .ZN(
        n11056) );
  INV_X1 U14111 ( .A(n11056), .ZN(n11057) );
  INV_X1 U14112 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14228) );
  OAI222_X1 U14113 ( .A1(n19727), .A2(n11164), .B1(n10891), .B2(n15549), .C1(
        n11059), .C2(n14228), .ZN(n14226) );
  AOI222_X1 U14114 ( .A1(P2_REIP_REG_18__SCAN_IN), .A2(n11078), .B1(n11160), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .C1(n11161), .C2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n15101) );
  NAND2_X1 U14115 ( .A1(n14218), .A2(n15100), .ZN(n11137) );
  AOI22_X1 U14116 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n11160), .B1(
        n11161), .B2(P2_EAX_REG_20__SCAN_IN), .ZN(n11061) );
  NAND2_X1 U14117 ( .A1(n11078), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11060) );
  AOI22_X1 U14118 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n11160), .B1(
        n11161), .B2(P2_EAX_REG_21__SCAN_IN), .ZN(n11063) );
  NAND2_X1 U14119 ( .A1(n11078), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11062) );
  NAND2_X1 U14120 ( .A1(n11063), .A2(n11062), .ZN(n14254) );
  AOI22_X1 U14121 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n11160), .B1(
        n11161), .B2(P2_EAX_REG_22__SCAN_IN), .ZN(n11065) );
  NAND2_X1 U14122 ( .A1(n11078), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11064) );
  AND2_X1 U14123 ( .A1(n11065), .A2(n11064), .ZN(n13087) );
  AOI22_X1 U14124 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n11160), .B1(
        n11161), .B2(P2_EAX_REG_23__SCAN_IN), .ZN(n11067) );
  NAND2_X1 U14125 ( .A1(n11078), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11066) );
  AND2_X1 U14126 ( .A1(n11067), .A2(n11066), .ZN(n13059) );
  AOI22_X1 U14127 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n11160), .B1(
        n11161), .B2(P2_EAX_REG_24__SCAN_IN), .ZN(n11069) );
  NAND2_X1 U14128 ( .A1(n11078), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11068) );
  NAND2_X1 U14129 ( .A1(n11069), .A2(n11068), .ZN(n15455) );
  AOI22_X1 U14130 ( .A1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n11160), .B1(
        n11161), .B2(P2_EAX_REG_25__SCAN_IN), .ZN(n11071) );
  NAND2_X1 U14131 ( .A1(n11078), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11070) );
  NAND2_X1 U14132 ( .A1(n11071), .A2(n11070), .ZN(n15079) );
  AOI22_X1 U14133 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n11160), .B1(
        n11161), .B2(P2_EAX_REG_26__SCAN_IN), .ZN(n11073) );
  NAND2_X1 U14134 ( .A1(n11078), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11072) );
  AND2_X1 U14135 ( .A1(n11073), .A2(n11072), .ZN(n15190) );
  AOI22_X1 U14136 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n11160), .B1(
        n11161), .B2(P2_EAX_REG_27__SCAN_IN), .ZN(n11075) );
  NAND2_X1 U14137 ( .A1(n11078), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11074) );
  AND2_X1 U14138 ( .A1(n11075), .A2(n11074), .ZN(n13072) );
  AOI22_X1 U14139 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n11160), .B1(
        n11161), .B2(P2_EAX_REG_28__SCAN_IN), .ZN(n11077) );
  NAND2_X1 U14140 ( .A1(n11078), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11076) );
  AND2_X1 U14141 ( .A1(n11077), .A2(n11076), .ZN(n12474) );
  AOI22_X1 U14142 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n11160), .B1(
        n11161), .B2(P2_EAX_REG_29__SCAN_IN), .ZN(n11080) );
  NAND2_X1 U14143 ( .A1(n11078), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11079) );
  NAND2_X1 U14144 ( .A1(n11080), .A2(n11079), .ZN(n11253) );
  NAND2_X1 U14145 ( .A1(n12476), .A2(n11253), .ZN(n11255) );
  AOI21_X1 U14146 ( .B1(n11081), .B2(n11255), .A(n11166), .ZN(n16173) );
  INV_X1 U14147 ( .A(n11082), .ZN(n11084) );
  NAND2_X1 U14148 ( .A1(n11084), .A2(n11083), .ZN(n16326) );
  NAND2_X1 U14149 ( .A1(n11263), .A2(n10673), .ZN(n16323) );
  NAND2_X1 U14150 ( .A1(n16323), .A2(n11085), .ZN(n11086) );
  AND2_X1 U14151 ( .A1(n16326), .A2(n11086), .ZN(n11087) );
  NOR2_X1 U14152 ( .A1(n19155), .A2(n19752), .ZN(n11192) );
  INV_X1 U14153 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11094) );
  INV_X1 U14154 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15573) );
  INV_X1 U14155 ( .A(n19175), .ZN(n15533) );
  NOR2_X1 U14156 ( .A1(n11090), .A2(n19191), .ZN(n19170) );
  OAI211_X1 U14157 ( .C1(n15533), .C2(n19170), .A(n19169), .B(n15671), .ZN(
        n16298) );
  INV_X1 U14158 ( .A(n14506), .ZN(n11091) );
  INV_X1 U14159 ( .A(n16282), .ZN(n11092) );
  NAND3_X1 U14160 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n15647), .ZN(n15614) );
  NOR2_X1 U14161 ( .A1(n15614), .A2(n11093), .ZN(n15586) );
  NAND2_X1 U14162 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15586), .ZN(
        n15570) );
  NOR3_X1 U14163 ( .A1(n11168), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n12480), .ZN(n11096) );
  AOI211_X1 U14164 ( .C1(n16173), .C2(n16296), .A(n11192), .B(n11096), .ZN(
        n11097) );
  OAI21_X1 U14165 ( .B1(n11170), .B2(n11167), .A(n11097), .ZN(n11098) );
  NAND3_X1 U14166 ( .A1(n11101), .A2(n11100), .A3(n10066), .ZN(P2_U3016) );
  INV_X1 U14167 ( .A(n11102), .ZN(n15292) );
  NOR2_X1 U14168 ( .A1(n15292), .A2(n11103), .ZN(n11111) );
  INV_X1 U14169 ( .A(n15306), .ZN(n11108) );
  NAND2_X1 U14170 ( .A1(n15280), .A2(n15368), .ZN(n15600) );
  INV_X1 U14171 ( .A(n15598), .ZN(n11104) );
  AOI21_X2 U14172 ( .B1(n15600), .B2(n15597), .A(n11104), .ZN(n15358) );
  NAND2_X1 U14173 ( .A1(n15358), .A2(n15359), .ZN(n15566) );
  NAND2_X1 U14174 ( .A1(n11105), .A2(n15566), .ZN(n15346) );
  NAND3_X1 U14175 ( .A1(n11108), .A2(n15317), .A3(n15320), .ZN(n15293) );
  INV_X1 U14176 ( .A(n15293), .ZN(n11109) );
  XOR2_X1 U14177 ( .A(n11111), .B(n11110), .Z(n11147) );
  NAND2_X1 U14178 ( .A1(n19823), .A2(n19673), .ZN(n11112) );
  NAND2_X1 U14179 ( .A1(n16356), .A2(n19822), .ZN(n11117) );
  OAI21_X1 U14180 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(
        P2_STATE2_REG_1__SCAN_IN), .A(n19822), .ZN(n16355) );
  INV_X1 U14181 ( .A(n16355), .ZN(n19824) );
  NOR2_X1 U14182 ( .A1(n19528), .A2(n13937), .ZN(n19799) );
  INV_X1 U14183 ( .A(n19799), .ZN(n11115) );
  NAND2_X1 U14184 ( .A1(n19824), .A2(n11115), .ZN(n11116) );
  AND2_X1 U14185 ( .A1(n9653), .A2(n11118), .ZN(n11120) );
  OR2_X1 U14186 ( .A1(n11120), .A2(n11119), .ZN(n18874) );
  NAND2_X1 U14187 ( .A1(n13937), .A2(n19794), .ZN(n18834) );
  INV_X1 U14188 ( .A(n18834), .ZN(n19763) );
  OR2_X1 U14189 ( .A1(n19764), .A2(n19763), .ZN(n19785) );
  NAND2_X1 U14190 ( .A1(n19785), .A2(n19822), .ZN(n11121) );
  NOR2_X1 U14191 ( .A1(n19155), .A2(n11122), .ZN(n11140) );
  NAND2_X1 U14192 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n11232) );
  NOR2_X1 U14193 ( .A1(n11232), .A2(n16274), .ZN(n11233) );
  AND2_X1 U14194 ( .A1(n11233), .A2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11123) );
  NAND2_X1 U14195 ( .A1(n11227), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n11228) );
  INV_X1 U14196 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n11224) );
  NAND2_X1 U14197 ( .A1(n11222), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11221) );
  INV_X1 U14198 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n15309) );
  NOR2_X1 U14199 ( .A1(n11125), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11126) );
  OR2_X1 U14200 ( .A1(n11190), .A2(n11126), .ZN(n11220) );
  NAND2_X1 U14201 ( .A1(n19822), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12518) );
  INV_X1 U14202 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19382) );
  NAND2_X1 U14203 ( .A1(n19382), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11127) );
  NAND2_X1 U14204 ( .A1(n12518), .A2(n11127), .ZN(n13310) );
  NOR2_X1 U14205 ( .A1(n11220), .A2(n15396), .ZN(n11128) );
  AOI211_X1 U14206 ( .C1(n15338), .C2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n11140), .B(n11128), .ZN(n11129) );
  OAI21_X1 U14207 ( .B1(n13862), .B2(n18874), .A(n11129), .ZN(n11130) );
  AOI21_X1 U14208 ( .B1(n11147), .B2(n11114), .A(n11130), .ZN(n11134) );
  NAND2_X1 U14209 ( .A1(n11131), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15276) );
  INV_X1 U14210 ( .A(n15276), .ZN(n15313) );
  OR2_X1 U14211 ( .A1(n15276), .A2(n15265), .ZN(n15300) );
  OAI21_X1 U14212 ( .B1(n15313), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15300), .ZN(n11148) );
  INV_X1 U14213 ( .A(n13110), .ZN(n11132) );
  NAND2_X1 U14214 ( .A1(n11134), .A2(n11133), .ZN(P2_U2994) );
  NAND2_X1 U14215 ( .A1(n15534), .A2(n11135), .ZN(n15512) );
  INV_X1 U14216 ( .A(n18874), .ZN(n11144) );
  AND2_X1 U14217 ( .A1(n11137), .A2(n11136), .ZN(n11138) );
  OR2_X1 U14218 ( .A1(n11138), .A2(n14255), .ZN(n18873) );
  OAI211_X1 U14219 ( .C1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(n15510), .B(n11139), .ZN(
        n11142) );
  INV_X1 U14220 ( .A(n11140), .ZN(n11141) );
  OAI211_X1 U14221 ( .C1(n19185), .C2(n18873), .A(n11142), .B(n11141), .ZN(
        n11143) );
  AOI21_X1 U14222 ( .B1(n11144), .B2(n16290), .A(n11143), .ZN(n11145) );
  OAI21_X1 U14223 ( .B1(n15265), .B2(n15512), .A(n11145), .ZN(n11146) );
  AOI21_X1 U14224 ( .B1(n11147), .B2(n19188), .A(n11146), .ZN(n11150) );
  NAND2_X1 U14225 ( .A1(n11150), .A2(n11149), .ZN(P2_U3026) );
  INV_X1 U14226 ( .A(n19174), .ZN(n11175) );
  INV_X1 U14227 ( .A(n11151), .ZN(n11152) );
  INV_X1 U14228 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19754) );
  NAND2_X1 U14229 ( .A1(n11153), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11156) );
  AOI22_X1 U14230 ( .A1(n11154), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11155) );
  OAI211_X1 U14231 ( .C1(n11157), .C2(n19754), .A(n11156), .B(n11155), .ZN(
        n11158) );
  NAND2_X1 U14232 ( .A1(n11160), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11163) );
  NAND2_X1 U14233 ( .A1(n11161), .A2(P2_EAX_REG_31__SCAN_IN), .ZN(n11162) );
  OAI211_X1 U14234 ( .C1(n11164), .C2(n19754), .A(n11163), .B(n11162), .ZN(
        n11165) );
  XNOR2_X1 U14235 ( .A(n11166), .B(n11165), .ZN(n15172) );
  NOR2_X1 U14236 ( .A1(n19155), .A2(n19754), .ZN(n12490) );
  INV_X1 U14237 ( .A(n12490), .ZN(n11169) );
  OAI21_X1 U14238 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14269), .A(
        n11170), .ZN(n11171) );
  NAND2_X1 U14239 ( .A1(n11171), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11172) );
  OAI211_X1 U14240 ( .C1(n14392), .C2(n19179), .A(n11173), .B(n11172), .ZN(
        n11174) );
  OAI211_X1 U14241 ( .C1(n11178), .C2(n11177), .A(n11176), .B(n15219), .ZN(
        n11185) );
  NOR2_X1 U14242 ( .A1(n11179), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11180) );
  MUX2_X1 U14243 ( .A(n11181), .B(n11180), .S(n12848), .Z(n11282) );
  NAND2_X1 U14244 ( .A1(n11282), .A2(n11182), .ZN(n11183) );
  XOR2_X1 U14245 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n11183), .Z(
        n11184) );
  XNOR2_X1 U14246 ( .A(n11185), .B(n11184), .ZN(n12493) );
  NAND2_X1 U14247 ( .A1(n12493), .A2(n19188), .ZN(n11186) );
  NAND2_X1 U14248 ( .A1(n11187), .A2(n11186), .ZN(P2_U3015) );
  INV_X1 U14249 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15269) );
  INV_X1 U14250 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n11215) );
  NOR2_X1 U14251 ( .A1(n15269), .A2(n11215), .ZN(n11188) );
  AND2_X1 U14252 ( .A1(n11188), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11189) );
  INV_X1 U14253 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n15231) );
  INV_X1 U14254 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n11203) );
  AND2_X1 U14255 ( .A1(n11204), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11200) );
  XNOR2_X1 U14256 ( .A(n11200), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16166) );
  NOR2_X1 U14257 ( .A1(n16166), .A2(n15396), .ZN(n11191) );
  AOI211_X1 U14258 ( .C1(n15338), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n11192), .B(n11191), .ZN(n11193) );
  OAI21_X1 U14259 ( .B1(n16172), .B2(n13862), .A(n11193), .ZN(n11194) );
  AOI21_X1 U14260 ( .B1(n11195), .B2(n11114), .A(n11194), .ZN(n11198) );
  OR2_X1 U14261 ( .A1(n11196), .A2(n19148), .ZN(n11197) );
  NAND2_X1 U14262 ( .A1(n11198), .A2(n11197), .ZN(P2_U2984) );
  NOR2_X1 U14263 ( .A1(n11204), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11199) );
  OR2_X1 U14264 ( .A1(n11200), .A2(n11199), .ZN(n15222) );
  INV_X1 U14265 ( .A(n15222), .ZN(n11249) );
  AND2_X1 U14266 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11201) );
  INV_X1 U14267 ( .A(n11225), .ZN(n11247) );
  AND2_X1 U14268 ( .A1(n11207), .A2(n11203), .ZN(n11205) );
  OR2_X1 U14269 ( .A1(n11205), .A2(n11204), .ZN(n12468) );
  INV_X1 U14270 ( .A(n12468), .ZN(n16185) );
  INV_X1 U14271 ( .A(n11207), .ZN(n11208) );
  AOI21_X1 U14272 ( .B1(n15231), .B2(n11206), .A(n11208), .ZN(n15229) );
  OR2_X1 U14273 ( .A1(n11212), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11209) );
  NAND2_X1 U14274 ( .A1(n11206), .A2(n11209), .ZN(n15237) );
  INV_X1 U14275 ( .A(n15237), .ZN(n16196) );
  NOR2_X1 U14276 ( .A1(n11210), .A2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n11211) );
  NOR2_X1 U14277 ( .A1(n11213), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n11214) );
  OR2_X1 U14278 ( .A1(n11210), .A2(n11214), .ZN(n15261) );
  INV_X1 U14279 ( .A(n15261), .ZN(n16207) );
  NAND2_X1 U14280 ( .A1(n11190), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n11218) );
  OR2_X1 U14281 ( .A1(n11218), .A2(n11215), .ZN(n11217) );
  AOI21_X1 U14282 ( .B1(n15269), .B2(n11217), .A(n11213), .ZN(n15271) );
  NAND2_X1 U14283 ( .A1(n11218), .A2(n11215), .ZN(n11216) );
  NAND2_X1 U14284 ( .A1(n11217), .A2(n11216), .ZN(n15287) );
  INV_X1 U14285 ( .A(n15287), .ZN(n13081) );
  OAI21_X1 U14286 ( .B1(n11190), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n11218), .ZN(n11219) );
  INV_X1 U14287 ( .A(n11219), .ZN(n18866) );
  INV_X1 U14288 ( .A(n11220), .ZN(n18878) );
  AOI21_X1 U14289 ( .B1(n15309), .B2(n11221), .A(n11125), .ZN(n15312) );
  OAI21_X1 U14290 ( .B1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n11222), .A(
        n11221), .ZN(n15323) );
  INV_X1 U14291 ( .A(n15323), .ZN(n15110) );
  AOI21_X1 U14292 ( .B1(n11224), .B2(n11223), .A(n11222), .ZN(n18893) );
  INV_X1 U14293 ( .A(n18893), .ZN(n18891) );
  OAI21_X1 U14294 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n11226), .A(
        n11244), .ZN(n18913) );
  INV_X1 U14295 ( .A(n18913), .ZN(n11243) );
  OAI21_X1 U14296 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n11227), .A(
        n11228), .ZN(n15371) );
  INV_X1 U14297 ( .A(n15371), .ZN(n18929) );
  AOI21_X1 U14298 ( .B1(n15382), .B2(n11229), .A(n11230), .ZN(n18956) );
  INV_X1 U14299 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16266) );
  AND2_X1 U14300 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n11231), .ZN(
        n11241) );
  AOI21_X1 U14301 ( .B1(n16266), .B2(n11239), .A(n11241), .ZN(n18963) );
  INV_X1 U14302 ( .A(n11234), .ZN(n11236) );
  OR2_X1 U14303 ( .A1(n11236), .A2(n11232), .ZN(n11237) );
  AND2_X1 U14304 ( .A1(n11234), .A2(n11233), .ZN(n11240) );
  AOI21_X1 U14305 ( .B1(n16274), .B2(n11237), .A(n11240), .ZN(n16267) );
  NOR2_X1 U14306 ( .A1(n10749), .A2(n11236), .ZN(n11238) );
  AOI21_X1 U14307 ( .B1(n10749), .B2(n11236), .A(n11238), .ZN(n19140) );
  AOI21_X1 U14308 ( .B1(n13690), .B2(n13826), .A(n11235), .ZN(n13687) );
  AOI22_X1 U14309 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n19822), .ZN(n19035) );
  AOI22_X1 U14310 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n13826), .B2(n19822), .ZN(
        n13832) );
  NAND2_X1 U14311 ( .A1(n19035), .A2(n13832), .ZN(n13831) );
  OAI21_X1 U14312 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11235), .A(
        n11236), .ZN(n13766) );
  OAI21_X1 U14313 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n11238), .A(
        n11237), .ZN(n18990) );
  NOR2_X1 U14314 ( .A1(n16267), .A2(n13752), .ZN(n18973) );
  OAI21_X1 U14315 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n11240), .A(
        n11239), .ZN(n18975) );
  NAND2_X1 U14316 ( .A1(n18973), .A2(n18975), .ZN(n18961) );
  OAI21_X1 U14317 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n11241), .A(
        n11229), .ZN(n15395) );
  INV_X1 U14318 ( .A(n11230), .ZN(n11242) );
  AOI21_X1 U14319 ( .B1(n10776), .B2(n11242), .A(n11227), .ZN(n16246) );
  INV_X1 U14320 ( .A(n16246), .ZN(n18950) );
  NOR2_X1 U14321 ( .A1(n18929), .A2(n18928), .ZN(n18918) );
  AOI21_X1 U14322 ( .B1(n16245), .B2(n11228), .A(n11226), .ZN(n16239) );
  INV_X1 U14323 ( .A(n16239), .ZN(n18919) );
  NAND2_X1 U14324 ( .A1(n18918), .A2(n18919), .ZN(n18911) );
  AOI21_X1 U14325 ( .B1(n16238), .B2(n11244), .A(n11245), .ZN(n16231) );
  INV_X1 U14326 ( .A(n16231), .ZN(n14202) );
  OAI21_X1 U14327 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n11245), .A(
        n11223), .ZN(n11246) );
  INV_X1 U14328 ( .A(n11246), .ZN(n18898) );
  OAI21_X1 U14329 ( .B1(n11247), .B2(n18891), .A(n18890), .ZN(n15109) );
  NOR2_X1 U14330 ( .A1(n15110), .A2(n15109), .ZN(n15108) );
  NOR2_X1 U14331 ( .A1(n11247), .A2(n15108), .ZN(n15095) );
  NOR2_X1 U14332 ( .A1(n15312), .A2(n15095), .ZN(n15094) );
  NOR2_X1 U14333 ( .A1(n11247), .A2(n15094), .ZN(n18877) );
  NOR2_X1 U14335 ( .A1(n11247), .A2(n13051), .ZN(n16205) );
  NOR2_X1 U14338 ( .A1(n11247), .A2(n15084), .ZN(n16195) );
  NOR3_X1 U14339 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(P2_STATEBS16_REG_SCAN_IN), .ZN(n15805) );
  NAND2_X1 U14340 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n15805), .ZN(n19677) );
  AOI211_X1 U14341 ( .C1(n11249), .C2(n11248), .A(n16165), .B(n19677), .ZN(
        n11277) );
  OAI21_X1 U14342 ( .B1(n12466), .B2(n11251), .A(n11250), .ZN(n15410) );
  NAND2_X1 U14343 ( .A1(n19819), .A2(n11252), .ZN(n11258) );
  NAND2_X1 U14344 ( .A1(n19825), .A2(n19382), .ZN(n11266) );
  OR2_X1 U14345 ( .A1(n12476), .A2(n11253), .ZN(n11254) );
  NAND2_X1 U14346 ( .A1(n11255), .A2(n11254), .ZN(n15406) );
  INV_X1 U14347 ( .A(n13107), .ZN(n13155) );
  NOR2_X1 U14348 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n13155), .ZN(n11265) );
  AND2_X1 U14349 ( .A1(n11256), .A2(n11265), .ZN(n16351) );
  NAND2_X1 U14350 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n11266), .ZN(n11257) );
  NOR3_X1 U14351 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n11259), .A3(n19794), 
        .ZN(n16346) );
  INV_X1 U14352 ( .A(n16346), .ZN(n11260) );
  NAND3_X1 U14353 ( .A1(n19677), .A2(n19155), .A3(n11260), .ZN(n11261) );
  AOI22_X1 U14354 ( .A1(n11262), .A2(n19022), .B1(P2_REIP_REG_29__SCAN_IN), 
        .B2(n19017), .ZN(n11272) );
  NAND2_X1 U14355 ( .A1(n18978), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19028) );
  INV_X1 U14356 ( .A(n11263), .ZN(n11264) );
  INV_X1 U14357 ( .A(n11265), .ZN(n11278) );
  NAND2_X1 U14358 ( .A1(n13211), .A2(n11278), .ZN(n11270) );
  INV_X1 U14359 ( .A(n11266), .ZN(n11267) );
  NOR2_X1 U14360 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n11267), .ZN(n11268) );
  NAND2_X1 U14361 ( .A1(n13112), .A2(n11268), .ZN(n11269) );
  NAND2_X2 U14362 ( .A1(n11270), .A2(n11269), .ZN(n19018) );
  AOI22_X1 U14363 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18997), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n19018), .ZN(n11271) );
  OAI211_X1 U14364 ( .C1(n15406), .C2(n19001), .A(n11272), .B(n11271), .ZN(
        n11273) );
  INV_X1 U14365 ( .A(n11273), .ZN(n11274) );
  OR2_X1 U14366 ( .A1(n11277), .A2(n11276), .ZN(P2_U2826) );
  NOR2_X1 U14367 ( .A1(n14392), .A2(n19004), .ZN(n11288) );
  INV_X1 U14368 ( .A(n19677), .ZN(n18993) );
  NAND2_X1 U14369 ( .A1(n19017), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n11280) );
  NAND3_X1 U14370 ( .A1(n13211), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n11278), 
        .ZN(n11279) );
  OAI211_X1 U14371 ( .C1(n19028), .C2(n11202), .A(n11280), .B(n11279), .ZN(
        n11281) );
  AOI21_X1 U14372 ( .B1(n11282), .B2(n19022), .A(n11281), .ZN(n11283) );
  NAND2_X1 U14373 ( .A1(n11286), .A2(n11285), .ZN(n11287) );
  AOI22_X1 U14374 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n17160), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n17125), .ZN(n11305) );
  AOI22_X1 U14375 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n17143), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n17156), .ZN(n11304) );
  NOR2_X2 U14376 ( .A1(n16880), .A2(n11292), .ZN(n11462) );
  AOI22_X1 U14377 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11290) );
  OAI21_X1 U14378 ( .B1(n11441), .B2(n17176), .A(n11290), .ZN(n11302) );
  INV_X2 U14379 ( .A(n12876), .ZN(n17155) );
  AOI22_X1 U14380 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11300) );
  INV_X4 U14381 ( .A(n16958), .ZN(n17020) );
  AOI22_X1 U14382 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11299) );
  AOI22_X1 U14383 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n9606), .B1(n9622), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11298) );
  AOI22_X1 U14384 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n9603), .B1(
        n12941), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11297) );
  NAND4_X1 U14385 ( .A1(n11300), .A2(n11299), .A3(n11298), .A4(n11297), .ZN(
        n11301) );
  AOI211_X1 U14386 ( .C1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .C2(n9602), .A(
        n11302), .B(n11301), .ZN(n11303) );
  AOI22_X1 U14387 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11310) );
  AOI22_X1 U14388 ( .A1(n17052), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11309) );
  AOI22_X1 U14389 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12941), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11308) );
  AOI22_X1 U14390 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11307) );
  NAND4_X1 U14391 ( .A1(n11310), .A2(n11309), .A3(n11308), .A4(n11307), .ZN(
        n11316) );
  AOI22_X1 U14392 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11314) );
  AOI22_X1 U14393 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11313) );
  AOI22_X1 U14394 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11312) );
  AOI22_X1 U14395 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9603), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11311) );
  NAND4_X1 U14396 ( .A1(n11314), .A2(n11313), .A3(n11312), .A4(n11311), .ZN(
        n11315) );
  AOI22_X1 U14397 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9606), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11326) );
  INV_X2 U14398 ( .A(n12876), .ZN(n17137) );
  AOI22_X1 U14399 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9603), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11325) );
  INV_X1 U14400 ( .A(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n20794) );
  AOI22_X1 U14401 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11317) );
  OAI21_X1 U14402 ( .B1(n9652), .B2(n20794), .A(n11317), .ZN(n11323) );
  AOI22_X1 U14403 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9622), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11321) );
  AOI22_X1 U14404 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(n9607), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11320) );
  AOI22_X1 U14405 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17161), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11319) );
  AOI22_X1 U14406 ( .A1(n12941), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11318) );
  NAND4_X1 U14407 ( .A1(n11321), .A2(n11320), .A3(n11319), .A4(n11318), .ZN(
        n11322) );
  AOI211_X1 U14408 ( .C1(n9605), .C2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A(
        n11323), .B(n11322), .ZN(n11324) );
  NAND3_X1 U14409 ( .A1(n11326), .A2(n11325), .A3(n11324), .ZN(n12425) );
  NAND2_X1 U14410 ( .A1(n18187), .A2(n12425), .ZN(n18610) );
  AOI22_X1 U14411 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11337) );
  AOI22_X1 U14412 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11336) );
  INV_X1 U14413 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17196) );
  AOI22_X1 U14414 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(n9603), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11328) );
  OAI21_X1 U14415 ( .B1(n11441), .B2(n17196), .A(n11328), .ZN(n11334) );
  AOI22_X1 U14416 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11332) );
  AOI22_X1 U14417 ( .A1(n17052), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11331) );
  AOI22_X1 U14418 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11330) );
  AOI22_X1 U14419 ( .A1(n12941), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11329) );
  NAND4_X1 U14420 ( .A1(n11332), .A2(n11331), .A3(n11330), .A4(n11329), .ZN(
        n11333) );
  AOI211_X1 U14421 ( .C1(n9605), .C2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A(
        n11334), .B(n11333), .ZN(n11335) );
  NAND3_X1 U14422 ( .A1(n11337), .A2(n11336), .A3(n11335), .ZN(n12990) );
  AOI22_X1 U14423 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11347) );
  AOI22_X1 U14424 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11346) );
  AOI22_X1 U14425 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11338) );
  OAI21_X1 U14426 ( .B1(n11441), .B2(n17181), .A(n11338), .ZN(n11344) );
  AOI22_X1 U14427 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11342) );
  AOI22_X1 U14428 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(n9607), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11341) );
  AOI22_X1 U14429 ( .A1(n9603), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n16916), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11340) );
  AOI22_X1 U14430 ( .A1(n9622), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12941), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11339) );
  NAND4_X1 U14431 ( .A1(n11342), .A2(n11341), .A3(n11340), .A4(n11339), .ZN(
        n11343) );
  AOI211_X1 U14432 ( .C1(n17020), .C2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n11344), .B(n11343), .ZN(n11345) );
  NAND3_X1 U14433 ( .A1(n11347), .A2(n11346), .A3(n11345), .ZN(n12437) );
  NOR2_X1 U14434 ( .A1(n12990), .A2(n18182), .ZN(n15714) );
  INV_X1 U14435 ( .A(n15714), .ZN(n15707) );
  AOI22_X1 U14436 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11358) );
  AOI22_X1 U14437 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11357) );
  AOI22_X1 U14438 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(n9603), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11348) );
  OAI21_X1 U14439 ( .B1(n11441), .B2(n17190), .A(n11348), .ZN(n11355) );
  AOI22_X1 U14440 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11353) );
  AOI22_X1 U14441 ( .A1(n9622), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n9602), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11352) );
  AOI22_X1 U14442 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11351) );
  AOI22_X1 U14443 ( .A1(n12941), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11350) );
  NAND4_X1 U14444 ( .A1(n11353), .A2(n11352), .A3(n11351), .A4(n11350), .ZN(
        n11354) );
  AOI211_X1 U14445 ( .C1(n9597), .C2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A(
        n11355), .B(n11354), .ZN(n11356) );
  NAND3_X1 U14446 ( .A1(n11358), .A2(n11357), .A3(n11356), .ZN(n12433) );
  NAND2_X1 U14447 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18634), .ZN(
        n12442) );
  OAI21_X1 U14448 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18634), .A(
        n12442), .ZN(n12996) );
  OAI22_X1 U14449 ( .A1(n18786), .A2(n18636), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n12443) );
  INV_X1 U14450 ( .A(n12443), .ZN(n11359) );
  NOR2_X1 U14451 ( .A1(n12996), .A2(n11359), .ZN(n11374) );
  OAI22_X1 U14452 ( .A1(n11361), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18641), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11365) );
  NOR2_X1 U14453 ( .A1(n11363), .A2(n18768), .ZN(n11368) );
  NAND2_X1 U14454 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18604), .ZN(
        n11364) );
  AOI22_X1 U14455 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18604), .B1(
        n11363), .B2(n18768), .ZN(n11367) );
  OAI22_X1 U14456 ( .A1(n11368), .A2(n11364), .B1(n11367), .B2(n20792), .ZN(
        n11371) );
  INV_X1 U14457 ( .A(n11371), .ZN(n11373) );
  XNOR2_X1 U14458 ( .A(n11366), .B(n11365), .ZN(n11372) );
  OAI21_X1 U14459 ( .B1(n20792), .B2(n11368), .A(n11367), .ZN(n11369) );
  OAI21_X1 U14460 ( .B1(n18604), .B2(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(
        n11369), .ZN(n11370) );
  INV_X1 U14461 ( .A(n11370), .ZN(n12441) );
  NAND2_X1 U14462 ( .A1(n17211), .A2(n18182), .ZN(n12992) );
  INV_X1 U14463 ( .A(n12433), .ZN(n18173) );
  AOI22_X1 U14464 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11379) );
  AOI22_X1 U14465 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17161), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11378) );
  AOI22_X1 U14466 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11377) );
  AOI22_X1 U14467 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12941), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11376) );
  NAND4_X1 U14468 ( .A1(n11379), .A2(n11378), .A3(n11377), .A4(n11376), .ZN(
        n11385) );
  AOI22_X1 U14469 ( .A1(n17052), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11383) );
  AOI22_X1 U14470 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11382) );
  AOI22_X1 U14471 ( .A1(n9603), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(n9602), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11381) );
  AOI22_X1 U14472 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9605), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11380) );
  NAND4_X1 U14473 ( .A1(n11383), .A2(n11382), .A3(n11381), .A4(n11380), .ZN(
        n11384) );
  AOI22_X1 U14474 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11389) );
  AOI22_X1 U14475 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9605), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11388) );
  AOI22_X1 U14476 ( .A1(n17052), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9603), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11387) );
  AOI22_X1 U14477 ( .A1(n12941), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11386) );
  NAND4_X1 U14478 ( .A1(n11389), .A2(n11388), .A3(n11387), .A4(n11386), .ZN(
        n11395) );
  AOI22_X1 U14479 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11393) );
  AOI22_X1 U14480 ( .A1(n9622), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11392) );
  AOI22_X1 U14481 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11391) );
  AOI22_X1 U14482 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(n9606), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11390) );
  NAND4_X1 U14483 ( .A1(n11393), .A2(n11392), .A3(n11391), .A4(n11390), .ZN(
        n11394) );
  NAND2_X1 U14484 ( .A1(n18773), .A2(P3_STATE2_REG_0__SCAN_IN), .ZN(n18664) );
  INV_X1 U14485 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n16898) );
  INV_X1 U14486 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16897) );
  INV_X1 U14487 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n16896) );
  INV_X1 U14488 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n16894) );
  INV_X1 U14489 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17011) );
  INV_X1 U14490 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16703) );
  INV_X1 U14491 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16724) );
  INV_X1 U14492 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n20839) );
  INV_X1 U14493 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n16849) );
  NAND3_X1 U14494 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17189) );
  NOR2_X1 U14495 ( .A1(n16849), .A2(n17189), .ZN(n17188) );
  INV_X1 U14496 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17119) );
  NOR2_X1 U14497 ( .A1(n16981), .A2(n17292), .ZN(n16982) );
  NAND2_X1 U14498 ( .A1(n16982), .A2(P3_EBX_REG_21__SCAN_IN), .ZN(n16970) );
  NOR2_X1 U14499 ( .A1(n17203), .A2(n16935), .ZN(n16936) );
  INV_X1 U14500 ( .A(n16942), .ZN(n16947) );
  NAND2_X1 U14501 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n16947), .ZN(n11474) );
  AOI22_X1 U14502 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11402) );
  AOI22_X1 U14503 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9603), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11401) );
  AOI22_X1 U14504 ( .A1(n11462), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17137), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11400) );
  AOI22_X1 U14505 ( .A1(n12941), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11399) );
  NAND4_X1 U14506 ( .A1(n11402), .A2(n11401), .A3(n11400), .A4(n11399), .ZN(
        n11409) );
  AOI22_X1 U14507 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(n9607), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11407) );
  AOI22_X1 U14508 ( .A1(n9622), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11406) );
  AOI22_X1 U14509 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11405) );
  AOI22_X1 U14510 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17161), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11404) );
  NAND4_X1 U14511 ( .A1(n11407), .A2(n11406), .A3(n11405), .A4(n11404), .ZN(
        n11408) );
  OR2_X1 U14512 ( .A1(n11409), .A2(n11408), .ZN(n16939) );
  AOI22_X1 U14513 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17161), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11414) );
  AOI22_X1 U14514 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11413) );
  AOI22_X1 U14515 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12941), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11412) );
  AOI22_X1 U14516 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9606), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11411) );
  NAND4_X1 U14517 ( .A1(n11414), .A2(n11413), .A3(n11412), .A4(n11411), .ZN(
        n11420) );
  AOI22_X1 U14518 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11418) );
  AOI22_X1 U14519 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11417) );
  AOI22_X1 U14520 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9603), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11416) );
  AOI22_X1 U14521 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11415) );
  NAND4_X1 U14522 ( .A1(n11418), .A2(n11417), .A3(n11416), .A4(n11415), .ZN(
        n11419) );
  NOR2_X1 U14523 ( .A1(n11420), .A2(n11419), .ZN(n16948) );
  AOI22_X1 U14524 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17161), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11424) );
  AOI22_X1 U14525 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11423) );
  AOI22_X1 U14526 ( .A1(n9603), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12941), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11422) );
  AOI22_X1 U14527 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11421) );
  NAND4_X1 U14528 ( .A1(n11424), .A2(n11423), .A3(n11422), .A4(n11421), .ZN(
        n11430) );
  AOI22_X1 U14529 ( .A1(n17052), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11428) );
  AOI22_X1 U14530 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11427) );
  AOI22_X1 U14531 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11426) );
  AOI22_X1 U14532 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17137), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11425) );
  NAND4_X1 U14533 ( .A1(n11428), .A2(n11427), .A3(n11426), .A4(n11425), .ZN(
        n11429) );
  NOR2_X1 U14534 ( .A1(n11430), .A2(n11429), .ZN(n16956) );
  AOI22_X1 U14535 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11434) );
  AOI22_X1 U14536 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11433) );
  AOI22_X1 U14537 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n17125), .ZN(n11432) );
  AOI22_X1 U14538 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n9607), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n12941), .ZN(n11431) );
  NAND4_X1 U14539 ( .A1(n11434), .A2(n11433), .A3(n11432), .A4(n11431), .ZN(
        n11440) );
  AOI22_X1 U14540 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n9606), .B1(
        P3_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n17143), .ZN(n11438) );
  AOI22_X1 U14541 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n9603), .B1(
        P3_INSTQUEUE_REG_0__7__SCAN_IN), .B2(n9602), .ZN(n11437) );
  AOI22_X1 U14542 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n17156), .B1(
        P3_INSTQUEUE_REG_12__7__SCAN_IN), .B2(n17160), .ZN(n11436) );
  AOI22_X1 U14543 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17161), .B1(
        n9605), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11435) );
  NAND4_X1 U14544 ( .A1(n11438), .A2(n11437), .A3(n11436), .A4(n11435), .ZN(
        n11439) );
  NOR2_X1 U14545 ( .A1(n11440), .A2(n11439), .ZN(n16955) );
  NOR2_X1 U14546 ( .A1(n16956), .A2(n16955), .ZN(n16952) );
  AOI22_X1 U14547 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11451) );
  AOI22_X1 U14548 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11450) );
  AOI22_X1 U14549 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9623), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11442) );
  OAI21_X1 U14550 ( .B1(n16958), .B2(n17198), .A(n11442), .ZN(n11448) );
  AOI22_X1 U14551 ( .A1(n9603), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(n9602), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11446) );
  AOI22_X1 U14552 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(n9605), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11445) );
  AOI22_X1 U14553 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11444) );
  AOI22_X1 U14554 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12941), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11443) );
  NAND4_X1 U14555 ( .A1(n11446), .A2(n11445), .A3(n11444), .A4(n11443), .ZN(
        n11447) );
  AOI211_X1 U14556 ( .C1(n9622), .C2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n11448), .B(n11447), .ZN(n11449) );
  NAND3_X1 U14557 ( .A1(n11451), .A2(n11450), .A3(n11449), .ZN(n16951) );
  NAND2_X1 U14558 ( .A1(n16952), .A2(n16951), .ZN(n16950) );
  NOR2_X1 U14559 ( .A1(n16948), .A2(n16950), .ZN(n16945) );
  AOI22_X1 U14560 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n9607), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11461) );
  AOI22_X1 U14561 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11460) );
  AOI22_X1 U14562 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17161), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11452) );
  OAI21_X1 U14563 ( .B1(n16958), .B2(n17190), .A(n11452), .ZN(n11458) );
  AOI22_X1 U14564 ( .A1(n9603), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11456) );
  AOI22_X1 U14565 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11455) );
  AOI22_X1 U14566 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n9622), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11454) );
  AOI22_X1 U14567 ( .A1(n12941), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11453) );
  NAND4_X1 U14568 ( .A1(n11456), .A2(n11455), .A3(n11454), .A4(n11453), .ZN(
        n11457) );
  AOI211_X1 U14569 ( .C1(n11462), .C2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A(
        n11458), .B(n11457), .ZN(n11459) );
  NAND3_X1 U14570 ( .A1(n11461), .A2(n11460), .A3(n11459), .ZN(n16944) );
  NAND2_X1 U14571 ( .A1(n16945), .A2(n16944), .ZN(n16943) );
  INV_X1 U14572 ( .A(n16943), .ZN(n16940) );
  NAND2_X1 U14573 ( .A1(n16939), .A2(n16940), .ZN(n16938) );
  AOI22_X1 U14574 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11466) );
  AOI22_X1 U14575 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17161), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11465) );
  AOI22_X1 U14576 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n9606), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11464) );
  AOI22_X1 U14577 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12941), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11463) );
  NAND4_X1 U14578 ( .A1(n11466), .A2(n11465), .A3(n11464), .A4(n11463), .ZN(
        n11472) );
  AOI22_X1 U14579 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11470) );
  AOI22_X1 U14580 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11469) );
  AOI22_X1 U14581 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9603), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11468) );
  AOI22_X1 U14582 ( .A1(n17125), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11467) );
  NAND4_X1 U14583 ( .A1(n11470), .A2(n11469), .A3(n11468), .A4(n11467), .ZN(
        n11471) );
  NOR2_X1 U14584 ( .A1(n11472), .A2(n11471), .ZN(n16931) );
  XOR2_X1 U14585 ( .A(n16938), .B(n16931), .Z(n17222) );
  NAND2_X1 U14586 ( .A1(n17203), .A2(n17222), .ZN(n11473) );
  AOI21_X1 U14587 ( .B1(n16936), .B2(P3_EBX_REG_28__SCAN_IN), .A(n11475), .ZN(
        n11476) );
  INV_X1 U14588 ( .A(n11476), .ZN(P3_U2675) );
  NOR2_X2 U14589 ( .A1(n11477), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11484) );
  NOR2_X2 U14590 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n11718), .ZN(
        n11483) );
  NOR2_X2 U14591 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11478), .ZN(
        n11486) );
  AND2_X2 U14592 ( .A1(n11486), .A2(n13347), .ZN(n11658) );
  AOI22_X1 U14593 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11658), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11482) );
  AOI22_X1 U14594 ( .A1(n11593), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11737), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11481) );
  AND2_X2 U14595 ( .A1(n11484), .A2(n13347), .ZN(n11602) );
  NOR2_X4 U14596 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11487) );
  AOI22_X1 U14597 ( .A1(n11602), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11480) );
  AND2_X2 U14598 ( .A1(n11486), .A2(n11483), .ZN(n11513) );
  AOI22_X1 U14599 ( .A1(n11513), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12202), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11479) );
  AND2_X4 U14600 ( .A1(n11483), .A2(n11487), .ZN(n11743) );
  AOI22_X1 U14601 ( .A1(n11743), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12293), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11491) );
  AOI22_X1 U14602 ( .A1(n12278), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11490) );
  AND2_X4 U14603 ( .A1(n11487), .A2(n13377), .ZN(n11659) );
  AOI22_X1 U14604 ( .A1(n11691), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11489) );
  AND3_X2 U14605 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13380) );
  AND2_X2 U14606 ( .A1(n13380), .A2(n14562), .ZN(n12249) );
  AND2_X4 U14607 ( .A1(n13380), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11690) );
  AOI22_X1 U14608 ( .A1(n12249), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11488) );
  NAND2_X1 U14609 ( .A1(n12293), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11496) );
  NAND2_X1 U14610 ( .A1(n11513), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11495) );
  NAND2_X1 U14611 ( .A1(n12278), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11494) );
  NAND2_X1 U14612 ( .A1(n9608), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11493) );
  NAND2_X1 U14613 ( .A1(n11602), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11500) );
  NAND2_X1 U14614 ( .A1(n11691), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11499) );
  NAND2_X1 U14615 ( .A1(n11737), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11498) );
  NAND2_X1 U14616 ( .A1(n11808), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11497) );
  NAND2_X1 U14617 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11504) );
  NAND2_X1 U14618 ( .A1(n11658), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11503) );
  NAND2_X1 U14619 ( .A1(n11743), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11502) );
  NAND2_X1 U14620 ( .A1(n11659), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11501) );
  NAND2_X1 U14621 ( .A1(n11593), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11508) );
  NAND2_X1 U14622 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11507) );
  NAND2_X1 U14623 ( .A1(n11690), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11506) );
  NAND2_X1 U14624 ( .A1(n12249), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11505) );
  NAND4_X4 U14625 ( .A1(n11512), .A2(n11511), .A3(n11510), .A4(n11509), .ZN(
        n11620) );
  NAND2_X1 U14626 ( .A1(n11635), .A2(n11620), .ZN(n11524) );
  AOI22_X1 U14627 ( .A1(n11513), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11737), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11517) );
  AOI22_X1 U14628 ( .A1(n11593), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11516) );
  AOI22_X1 U14629 ( .A1(n9630), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11492), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11515) );
  AOI22_X1 U14630 ( .A1(n12249), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11514) );
  NAND4_X1 U14631 ( .A1(n11517), .A2(n11516), .A3(n11515), .A4(n11514), .ZN(
        n11523) );
  AOI22_X1 U14632 ( .A1(n11602), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11658), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11521) );
  AOI22_X1 U14633 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9624), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11519) );
  AOI22_X1 U14634 ( .A1(n11691), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11518) );
  NAND4_X1 U14635 ( .A1(n11521), .A2(n11520), .A3(n11519), .A4(n11518), .ZN(
        n11522) );
  OR2_X2 U14636 ( .A1(n11523), .A2(n11522), .ZN(n11547) );
  NAND2_X1 U14637 ( .A1(n11524), .A2(n12341), .ZN(n11546) );
  NAND2_X1 U14638 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11528) );
  NAND2_X1 U14639 ( .A1(n11602), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11527) );
  NAND2_X1 U14640 ( .A1(n11658), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11526) );
  NAND2_X1 U14641 ( .A1(n11659), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11525) );
  NAND2_X1 U14642 ( .A1(n9629), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11532) );
  NAND2_X1 U14643 ( .A1(n11513), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11531) );
  NAND2_X1 U14644 ( .A1(n11737), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11530) );
  NAND2_X1 U14645 ( .A1(n11492), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11529) );
  NAND2_X1 U14646 ( .A1(n11691), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11536) );
  NAND2_X1 U14647 ( .A1(n12293), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11535) );
  NAND2_X1 U14648 ( .A1(n9628), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11534) );
  NAND2_X1 U14649 ( .A1(n11808), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11533) );
  NAND2_X1 U14650 ( .A1(n11593), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11540) );
  NAND2_X1 U14651 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11539) );
  NAND2_X1 U14652 ( .A1(n12249), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11538) );
  NAND2_X1 U14653 ( .A1(n11690), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11537) );
  NAND2_X1 U14654 ( .A1(n11546), .A2(n11545), .ZN(n11572) );
  AOI22_X1 U14655 ( .A1(n11602), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11658), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11551) );
  AOI22_X1 U14656 ( .A1(n11691), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12278), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11550) );
  AOI22_X1 U14657 ( .A1(n11593), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9608), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11549) );
  AOI22_X1 U14658 ( .A1(n12249), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11548) );
  NAND4_X1 U14659 ( .A1(n11551), .A2(n11550), .A3(n11549), .A4(n11548), .ZN(
        n11557) );
  AOI22_X1 U14660 ( .A1(n12293), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11513), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n11555) );
  AOI22_X1 U14661 ( .A1(n11737), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11554) );
  AOI22_X1 U14662 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11553) );
  AOI22_X1 U14663 ( .A1(n11743), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11552) );
  NAND4_X1 U14664 ( .A1(n11555), .A2(n11554), .A3(n11553), .A4(n11552), .ZN(
        n11556) );
  AOI22_X1 U14665 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11602), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11562) );
  AOI22_X1 U14666 ( .A1(n11593), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11561) );
  AOI22_X1 U14667 ( .A1(n12278), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11808), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11560) );
  NAND4_X1 U14668 ( .A1(n11562), .A2(n11561), .A3(n11560), .A4(n11559), .ZN(
        n11568) );
  AOI22_X1 U14669 ( .A1(n12293), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11737), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11566) );
  AOI22_X1 U14670 ( .A1(n11691), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11743), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11565) );
  AOI22_X1 U14671 ( .A1(n11658), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11564) );
  AOI22_X1 U14672 ( .A1(n12249), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11563) );
  NAND4_X1 U14673 ( .A1(n11566), .A2(n11565), .A3(n11564), .A4(n11563), .ZN(
        n11567) );
  OR2_X2 U14674 ( .A1(n11568), .A2(n11567), .ZN(n13246) );
  NAND2_X1 U14675 ( .A1(n11634), .A2(n13246), .ZN(n11571) );
  AOI21_X1 U14676 ( .B1(n13400), .B2(n13359), .A(n20141), .ZN(n11570) );
  NAND2_X1 U14677 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11576) );
  NAND2_X1 U14678 ( .A1(n11602), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11575) );
  NAND2_X1 U14679 ( .A1(n11658), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11574) );
  NAND2_X1 U14680 ( .A1(n11659), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11573) );
  NAND2_X1 U14681 ( .A1(n12278), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11580) );
  NAND2_X1 U14682 ( .A1(n11513), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11579) );
  NAND2_X1 U14683 ( .A1(n11737), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11578) );
  NAND2_X1 U14684 ( .A1(n12202), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11577) );
  NAND2_X1 U14685 ( .A1(n11691), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11584) );
  NAND2_X1 U14686 ( .A1(n12293), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11583) );
  NAND2_X1 U14687 ( .A1(n11743), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11582) );
  NAND2_X1 U14688 ( .A1(n11808), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11581) );
  NAND2_X1 U14689 ( .A1(n11593), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11588) );
  NAND2_X1 U14690 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11587) );
  NAND2_X1 U14691 ( .A1(n12249), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11586) );
  NAND2_X1 U14692 ( .A1(n11690), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11585) );
  NAND4_X4 U14693 ( .A1(n11592), .A2(n11591), .A3(n11590), .A4(n11589), .ZN(
        n14596) );
  INV_X1 U14694 ( .A(n13094), .ZN(n11615) );
  NAND2_X1 U14695 ( .A1(n12278), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11597) );
  NAND2_X1 U14696 ( .A1(n11593), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11596) );
  NAND2_X1 U14697 ( .A1(n11738), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11595) );
  NAND2_X1 U14698 ( .A1(n12202), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11594) );
  NAND2_X1 U14699 ( .A1(n11691), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11601) );
  NAND2_X1 U14700 ( .A1(n12293), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11600) );
  NAND2_X1 U14701 ( .A1(n11744), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11599) );
  NAND2_X1 U14702 ( .A1(n11743), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11598) );
  NAND2_X1 U14703 ( .A1(n11658), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11606) );
  NAND2_X1 U14704 ( .A1(n11602), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11605) );
  NAND2_X1 U14705 ( .A1(n11659), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11604) );
  NAND2_X1 U14706 ( .A1(n11808), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11603) );
  NAND2_X1 U14707 ( .A1(n11513), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11610) );
  NAND2_X1 U14708 ( .A1(n11737), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11609) );
  NAND2_X1 U14709 ( .A1(n12249), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11608) );
  NAND2_X1 U14710 ( .A1(n11690), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11607) );
  NAND4_X4 U14711 ( .A1(n11614), .A2(n11613), .A3(n11612), .A4(n11611), .ZN(
        n13907) );
  INV_X4 U14712 ( .A(n13907), .ZN(n20120) );
  NAND2_X1 U14713 ( .A1(n11615), .A2(n20120), .ZN(n12321) );
  AND2_X2 U14714 ( .A1(n11635), .A2(n13246), .ZN(n13395) );
  NOR2_X1 U14715 ( .A1(n12341), .A2(n11569), .ZN(n11616) );
  NAND2_X1 U14716 ( .A1(n11617), .A2(n14467), .ZN(n12348) );
  AND2_X2 U14717 ( .A1(n12321), .A2(n12348), .ZN(n13269) );
  INV_X1 U14718 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n11618) );
  XNOR2_X1 U14719 ( .A(n11618), .B(P1_STATE_REG_1__SCAN_IN), .ZN(n13098) );
  INV_X1 U14720 ( .A(n13098), .ZN(n11619) );
  NOR2_X1 U14721 ( .A1(n13095), .A2(n11619), .ZN(n11623) );
  NOR2_X2 U14722 ( .A1(n13359), .A2(n13246), .ZN(n13426) );
  NAND2_X1 U14723 ( .A1(n12341), .A2(n11631), .ZN(n13260) );
  NOR2_X2 U14724 ( .A1(n13349), .A2(n13260), .ZN(n13283) );
  NOR2_X1 U14725 ( .A1(n11623), .A2(n13283), .ZN(n11624) );
  NAND2_X1 U14726 ( .A1(n13269), .A2(n11624), .ZN(n11625) );
  NAND2_X2 U14727 ( .A1(n11625), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11716) );
  OR2_X1 U14728 ( .A1(n13574), .A2(n13400), .ZN(n11628) );
  NAND2_X2 U14729 ( .A1(n20120), .A2(n14596), .ZN(n14593) );
  OR2_X1 U14730 ( .A1(n14593), .A2(n11626), .ZN(n11627) );
  INV_X1 U14731 ( .A(n13395), .ZN(n11629) );
  INV_X1 U14732 ( .A(n13246), .ZN(n20127) );
  NAND2_X1 U14733 ( .A1(n20127), .A2(n14596), .ZN(n14291) );
  NAND2_X2 U14734 ( .A1(n14291), .A2(n13574), .ZN(n14525) );
  NAND2_X1 U14735 ( .A1(n11629), .A2(n14525), .ZN(n13273) );
  NAND2_X1 U14736 ( .A1(n9667), .A2(n20105), .ZN(n13352) );
  NAND2_X1 U14737 ( .A1(n11630), .A2(n12341), .ZN(n11632) );
  NAND2_X1 U14738 ( .A1(n13254), .A2(n11634), .ZN(n11642) );
  MUX2_X1 U14739 ( .A(n11635), .B(n20120), .S(n20105), .Z(n13280) );
  NAND3_X1 U14740 ( .A1(n9666), .A2(n13352), .A3(n10078), .ZN(n13272) );
  NAND2_X1 U14741 ( .A1(n13272), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11636) );
  MUX2_X1 U14742 ( .A(n13403), .B(n20660), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n11637) );
  INV_X1 U14743 ( .A(n11637), .ZN(n11638) );
  OR2_X1 U14744 ( .A1(n11640), .A2(n12341), .ZN(n11641) );
  NAND2_X1 U14745 ( .A1(n13352), .A2(n11641), .ZN(n13281) );
  INV_X1 U14746 ( .A(n13281), .ZN(n11651) );
  INV_X1 U14747 ( .A(n11642), .ZN(n11643) );
  NAND2_X1 U14748 ( .A1(n11643), .A2(n13907), .ZN(n11650) );
  NAND2_X1 U14749 ( .A1(n20105), .A2(n20120), .ZN(n14588) );
  NAND2_X1 U14750 ( .A1(n11633), .A2(n13246), .ZN(n11646) );
  INV_X1 U14751 ( .A(n11644), .ZN(n11645) );
  OAI211_X1 U14752 ( .C1(n12345), .C2(n14593), .A(P1_STATE2_REG_0__SCAN_IN), 
        .B(n16151), .ZN(n11647) );
  INV_X1 U14753 ( .A(n11647), .ZN(n11648) );
  INV_X1 U14754 ( .A(n14146), .ZN(n11678) );
  AOI22_X1 U14755 ( .A1(n11513), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11657) );
  AOI22_X1 U14757 ( .A1(n11593), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11653), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11656) );
  AOI22_X1 U14758 ( .A1(n12278), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12202), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11655) );
  AOI22_X1 U14759 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11654) );
  NAND4_X1 U14760 ( .A1(n11657), .A2(n11656), .A3(n11655), .A4(n11654), .ZN(
        n11665) );
  AOI22_X1 U14761 ( .A1(n12161), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11663) );
  AOI22_X1 U14762 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11743), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11662) );
  AOI22_X1 U14763 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11661) );
  INV_X1 U14764 ( .A(n11691), .ZN(n13379) );
  AOI22_X1 U14765 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11660) );
  NAND4_X1 U14766 ( .A1(n11663), .A2(n11662), .A3(n11661), .A4(n11660), .ZN(
        n11664) );
  AOI22_X1 U14767 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12278), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11670) );
  BUF_X1 U14768 ( .A(n11737), .Z(n11666) );
  AOI22_X1 U14769 ( .A1(n11593), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11669) );
  AOI22_X1 U14770 ( .A1(n11602), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11743), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11668) );
  AOI22_X1 U14771 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11667) );
  NAND4_X1 U14772 ( .A1(n11670), .A2(n11669), .A3(n11668), .A4(n11667), .ZN(
        n11676) );
  AOI22_X1 U14773 ( .A1(n12233), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11653), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11674) );
  AOI22_X1 U14774 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11673) );
  AOI22_X1 U14775 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11672) );
  AOI22_X1 U14776 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12202), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11671) );
  NAND4_X1 U14777 ( .A1(n11674), .A2(n11673), .A3(n11672), .A4(n11671), .ZN(
        n11675) );
  XNOR2_X1 U14778 ( .A(n11683), .B(n13471), .ZN(n11677) );
  NAND2_X1 U14779 ( .A1(n11678), .A2(n11677), .ZN(n11679) );
  INV_X1 U14780 ( .A(n13471), .ZN(n11682) );
  NAND2_X1 U14781 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11681) );
  AOI21_X1 U14782 ( .B1(n11626), .B2(n14151), .A(n20756), .ZN(n11680) );
  OAI211_X1 U14783 ( .C1(n11682), .C2(n14596), .A(n11681), .B(n11680), .ZN(
        n11770) );
  NAND2_X1 U14784 ( .A1(n11771), .A2(n11770), .ZN(n11685) );
  NAND2_X1 U14785 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11700) );
  OR2_X1 U14786 ( .A1(n14146), .A2(n14151), .ZN(n11699) );
  AOI22_X1 U14787 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12278), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11689) );
  AOI22_X1 U14788 ( .A1(n11593), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11653), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11688) );
  AOI22_X1 U14789 ( .A1(n12161), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11743), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11687) );
  AOI22_X1 U14790 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11686) );
  NAND4_X1 U14791 ( .A1(n11689), .A2(n11688), .A3(n11687), .A4(n11686), .ZN(
        n11697) );
  AOI22_X1 U14792 ( .A1(n12233), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U14793 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U14794 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U14795 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12202), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11692) );
  NAND4_X1 U14796 ( .A1(n11695), .A2(n11694), .A3(n11693), .A4(n11692), .ZN(
        n11696) );
  OR2_X1 U14797 ( .A1(n11784), .A2(n11709), .ZN(n11698) );
  NAND2_X1 U14798 ( .A1(n11722), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11703) );
  NAND2_X1 U14799 ( .A1(n20424), .A2(n20519), .ZN(n11701) );
  NAND2_X1 U14800 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11726) );
  AND2_X1 U14801 ( .A1(n11701), .A2(n11726), .ZN(n20428) );
  AND2_X1 U14802 ( .A1(n20660), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11717) );
  AOI21_X1 U14803 ( .B1(n13403), .B2(n20428), .A(n11717), .ZN(n11702) );
  XNOR2_X2 U14804 ( .A(n11704), .B(n11716), .ZN(n20214) );
  INV_X1 U14805 ( .A(n20214), .ZN(n11707) );
  INV_X1 U14806 ( .A(n11708), .ZN(n11706) );
  NAND2_X2 U14807 ( .A1(n20214), .A2(n11708), .ZN(n11735) );
  INV_X1 U14808 ( .A(n13348), .ZN(n11710) );
  AOI21_X2 U14809 ( .B1(n11710), .B2(n20756), .A(n10055), .ZN(n13394) );
  NAND2_X1 U14810 ( .A1(n11761), .A2(n13394), .ZN(n11715) );
  INV_X1 U14811 ( .A(n11711), .ZN(n11712) );
  NAND2_X1 U14812 ( .A1(n11715), .A2(n11714), .ZN(n11754) );
  INV_X1 U14813 ( .A(n11716), .ZN(n11721) );
  INV_X1 U14814 ( .A(n11717), .ZN(n11719) );
  NAND2_X1 U14815 ( .A1(n11719), .A2(n11718), .ZN(n11720) );
  NAND2_X1 U14816 ( .A1(n11721), .A2(n11720), .ZN(n11733) );
  NAND2_X1 U14817 ( .A1(n11735), .A2(n11733), .ZN(n11729) );
  NAND2_X1 U14818 ( .A1(n11722), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11724) );
  NAND2_X1 U14819 ( .A1(n20660), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11723) );
  INV_X1 U14820 ( .A(n11726), .ZN(n11725) );
  NAND2_X1 U14821 ( .A1(n11725), .A2(n20488), .ZN(n20458) );
  NAND2_X1 U14822 ( .A1(n11726), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11727) );
  NAND2_X1 U14823 ( .A1(n20458), .A2(n11727), .ZN(n20114) );
  AND2_X1 U14824 ( .A1(n13403), .A2(n20114), .ZN(n11731) );
  NAND2_X1 U14825 ( .A1(n11729), .A2(n11728), .ZN(n11780) );
  INV_X1 U14826 ( .A(n11730), .ZN(n11734) );
  INV_X1 U14827 ( .A(n11731), .ZN(n11732) );
  NAND4_X1 U14828 ( .A1(n11735), .A2(n11734), .A3(n11733), .A4(n11732), .ZN(
        n11736) );
  NAND2_X1 U14829 ( .A1(n11780), .A2(n11736), .ZN(n13421) );
  AOI22_X1 U14830 ( .A1(n12233), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11742) );
  AOI22_X1 U14831 ( .A1(n11593), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11653), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11741) );
  AOI22_X1 U14832 ( .A1(n12278), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12202), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11740) );
  AOI22_X1 U14833 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11739) );
  NAND4_X1 U14834 ( .A1(n11742), .A2(n11741), .A3(n11740), .A4(n11739), .ZN(
        n11750) );
  AOI22_X1 U14835 ( .A1(n12161), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11748) );
  AOI22_X1 U14836 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11743), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11747) );
  AOI22_X1 U14837 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11746) );
  INV_X2 U14838 ( .A(n13379), .ZN(n12294) );
  AOI22_X1 U14839 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11745) );
  NAND4_X1 U14840 ( .A1(n11748), .A2(n11747), .A3(n11746), .A4(n11745), .ZN(
        n11749) );
  NAND2_X1 U14841 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11751) );
  OAI21_X1 U14842 ( .B1(n11784), .B2(n13468), .A(n11751), .ZN(n11752) );
  NAND2_X1 U14843 ( .A1(n11755), .A2(n11754), .ZN(n11756) );
  INV_X1 U14844 ( .A(n13260), .ZN(n13415) );
  NAND2_X1 U14845 ( .A1(n13415), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n11831) );
  XNOR2_X1 U14846 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13919) );
  AOI21_X1 U14847 ( .B1(n12290), .B2(n13919), .A(n12318), .ZN(n11758) );
  NAND2_X1 U14848 ( .A1(n12319), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11757) );
  OAI211_X1 U14849 ( .C1(n11831), .C2(n11478), .A(n11758), .B(n11757), .ZN(
        n11759) );
  INV_X1 U14850 ( .A(n11759), .ZN(n11760) );
  NAND2_X1 U14851 ( .A1(n12318), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11779) );
  NAND2_X1 U14852 ( .A1(n9593), .A2(n12003), .ZN(n11769) );
  AOI22_X1 U14853 ( .A1(n12319), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20752), .ZN(n11767) );
  INV_X1 U14854 ( .A(n11831), .ZN(n11765) );
  NAND2_X1 U14855 ( .A1(n11765), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11766) );
  AND2_X1 U14856 ( .A1(n11767), .A2(n11766), .ZN(n11768) );
  NAND2_X1 U14857 ( .A1(n11769), .A2(n11768), .ZN(n13393) );
  NAND2_X1 U14858 ( .A1(n13249), .A2(n9938), .ZN(n11772) );
  NAND2_X1 U14859 ( .A1(n11772), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13316) );
  NAND2_X1 U14860 ( .A1(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n20752), .ZN(
        n11775) );
  NAND2_X1 U14861 ( .A1(n12319), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n11774) );
  OAI211_X1 U14862 ( .C1(n11831), .C2(n14562), .A(n11775), .B(n11774), .ZN(
        n11776) );
  AOI21_X1 U14863 ( .B1(n9621), .B2(n12003), .A(n11776), .ZN(n13317) );
  OR2_X1 U14864 ( .A1(n13316), .A2(n13317), .ZN(n13318) );
  NAND2_X1 U14865 ( .A1(n13317), .A2(n12290), .ZN(n11777) );
  NAND2_X1 U14866 ( .A1(n13318), .A2(n11777), .ZN(n13392) );
  INV_X1 U14867 ( .A(n13564), .ZN(n11778) );
  NAND2_X1 U14868 ( .A1(n11722), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11783) );
  NAND3_X1 U14869 ( .A1(n20738), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20345) );
  INV_X1 U14870 ( .A(n20365), .ZN(n11781) );
  NAND3_X1 U14871 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20604) );
  AOI21_X1 U14872 ( .B1(n20738), .B2(n11781), .A(n20648), .ZN(n20373) );
  AOI22_X1 U14873 ( .A1(n13403), .A2(n20373), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20660), .ZN(n11782) );
  AOI22_X1 U14874 ( .A1(n12233), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11788) );
  AOI22_X1 U14875 ( .A1(n11593), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11653), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U14876 ( .A1(n12278), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12202), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11786) );
  AOI22_X1 U14877 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11785) );
  NAND4_X1 U14878 ( .A1(n11788), .A2(n11787), .A3(n11786), .A4(n11785), .ZN(
        n11794) );
  AOI22_X1 U14879 ( .A1(n12161), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11792) );
  INV_X1 U14880 ( .A(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n20811) );
  AOI22_X1 U14881 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11743), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11791) );
  AOI22_X1 U14882 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11790) );
  AOI22_X1 U14883 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11789) );
  NAND4_X1 U14884 ( .A1(n11792), .A2(n11791), .A3(n11790), .A4(n11789), .ZN(
        n11793) );
  AOI22_X1 U14885 ( .A1(n12357), .A2(n13631), .B1(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n12385), .ZN(n11795) );
  NAND2_X1 U14886 ( .A1(n11798), .A2(n20258), .ZN(n11799) );
  INV_X1 U14887 ( .A(n11801), .ZN(n11802) );
  INV_X1 U14888 ( .A(n11825), .ZN(n11826) );
  OAI21_X1 U14889 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n11802), .A(
        n11826), .ZN(n19925) );
  AOI22_X1 U14890 ( .A1(n12290), .A2(n19925), .B1(n12318), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n11804) );
  NAND2_X1 U14891 ( .A1(n12311), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n11803) );
  OAI211_X1 U14892 ( .C1(n11831), .C2(n11477), .A(n11804), .B(n11803), .ZN(
        n11805) );
  INV_X1 U14893 ( .A(n11805), .ZN(n11806) );
  OAI21_X1 U14894 ( .B1(n20730), .B2(n11975), .A(n11806), .ZN(n13571) );
  AOI22_X1 U14895 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12161), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11812) );
  AOI22_X1 U14896 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n9631), .B1(
        n11653), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11811) );
  AOI22_X1 U14897 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12294), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11810) );
  AOI22_X1 U14898 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n11690), .B1(
        n12249), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11809) );
  NAND4_X1 U14899 ( .A1(n11812), .A2(n11811), .A3(n11810), .A4(n11809), .ZN(
        n11818) );
  AOI22_X1 U14900 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n12228), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11816) );
  AOI22_X1 U14901 ( .A1(n12278), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11743), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11815) );
  AOI22_X1 U14902 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11814) );
  AOI22_X1 U14903 ( .A1(n12233), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12202), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11813) );
  NAND4_X1 U14904 ( .A1(n11816), .A2(n11815), .A3(n11814), .A4(n11813), .ZN(
        n11817) );
  NAND2_X1 U14905 ( .A1(n12357), .A2(n13841), .ZN(n11820) );
  NAND2_X1 U14906 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11819) );
  NAND2_X1 U14907 ( .A1(n11820), .A2(n11819), .ZN(n11822) );
  NAND2_X1 U14908 ( .A1(n11807), .A2(n9947), .ZN(n11823) );
  NAND2_X1 U14909 ( .A1(n11846), .A2(n11823), .ZN(n13717) );
  INV_X1 U14910 ( .A(n13717), .ZN(n11824) );
  NAND2_X1 U14911 ( .A1(n11824), .A2(n12003), .ZN(n11834) );
  INV_X1 U14912 ( .A(n11848), .ZN(n11828) );
  INV_X1 U14913 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n20800) );
  NAND2_X1 U14914 ( .A1(n20800), .A2(n11826), .ZN(n11827) );
  NAND2_X1 U14915 ( .A1(n11828), .A2(n11827), .ZN(n14691) );
  INV_X1 U14916 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20753) );
  OAI21_X1 U14917 ( .B1(n20753), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20752), .ZN(n11830) );
  NAND2_X1 U14918 ( .A1(n12311), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n11829) );
  OAI211_X1 U14919 ( .C1(n11831), .C2(n16154), .A(n11830), .B(n11829), .ZN(
        n11832) );
  OAI21_X1 U14920 ( .B1(n12317), .B2(n14691), .A(n11832), .ZN(n11833) );
  AOI22_X1 U14921 ( .A1(n12233), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11838) );
  AOI22_X1 U14922 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11653), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U14923 ( .A1(n9630), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12202), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11836) );
  AOI22_X1 U14924 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11835) );
  NAND4_X1 U14925 ( .A1(n11838), .A2(n11837), .A3(n11836), .A4(n11835), .ZN(
        n11844) );
  AOI22_X1 U14926 ( .A1(n12161), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11842) );
  AOI22_X1 U14927 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11743), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11841) );
  AOI22_X1 U14928 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11840) );
  INV_X1 U14929 ( .A(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n20877) );
  AOI22_X1 U14930 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11839) );
  NAND4_X1 U14931 ( .A1(n11842), .A2(n11841), .A3(n11840), .A4(n11839), .ZN(
        n11843) );
  AOI22_X1 U14932 ( .A1(n12357), .A2(n13844), .B1(
        P1_INSTQUEUE_REG_0__5__SCAN_IN), .B2(n12385), .ZN(n11845) );
  NAND2_X1 U14933 ( .A1(n11846), .A2(n11845), .ZN(n11847) );
  NOR2_X1 U14934 ( .A1(n11848), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11849) );
  NOR2_X1 U14935 ( .A1(n11863), .A2(n11849), .ZN(n19914) );
  INV_X1 U14936 ( .A(n12318), .ZN(n11954) );
  INV_X1 U14937 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16027) );
  OAI22_X1 U14938 ( .A1(n19914), .A2(n12317), .B1(n11954), .B2(n16027), .ZN(
        n11850) );
  AOI21_X1 U14939 ( .B1(n12311), .B2(P1_EAX_REG_5__SCAN_IN), .A(n11850), .ZN(
        n11851) );
  NAND2_X1 U14940 ( .A1(n11852), .A2(n11851), .ZN(n13725) );
  INV_X1 U14941 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n11870) );
  AOI22_X1 U14942 ( .A1(n12161), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11856) );
  AOI22_X1 U14943 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11855) );
  AOI22_X1 U14944 ( .A1(n12233), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11743), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11854) );
  AOI22_X1 U14945 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11853) );
  NAND4_X1 U14946 ( .A1(n11856), .A2(n11855), .A3(n11854), .A4(n11853), .ZN(
        n11862) );
  AOI22_X1 U14947 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12278), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11860) );
  AOI22_X1 U14948 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11859) );
  AOI22_X1 U14949 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11858) );
  AOI22_X1 U14950 ( .A1(n11653), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n12202), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11857) );
  NAND4_X1 U14951 ( .A1(n11860), .A2(n11859), .A3(n11858), .A4(n11857), .ZN(
        n11861) );
  AOI22_X1 U14952 ( .A1(n12357), .A2(n14137), .B1(n12385), .B2(
        P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11872) );
  NAND2_X1 U14953 ( .A1(n11871), .A2(n11872), .ZN(n14130) );
  NAND2_X1 U14954 ( .A1(n14130), .A2(n12003), .ZN(n11869) );
  INV_X1 U14955 ( .A(n11876), .ZN(n11867) );
  INV_X1 U14956 ( .A(n11863), .ZN(n11865) );
  INV_X1 U14957 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11864) );
  NAND2_X1 U14958 ( .A1(n11865), .A2(n11864), .ZN(n11866) );
  NAND2_X1 U14959 ( .A1(n11867), .A2(n11866), .ZN(n19910) );
  AOI22_X1 U14960 ( .A1(n19910), .A2(n13895), .B1(n12318), .B2(
        P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n11868) );
  OAI211_X1 U14961 ( .C1(n12043), .C2(n11870), .A(n11869), .B(n11868), .ZN(
        n13791) );
  NAND2_X1 U14962 ( .A1(n12357), .A2(n14151), .ZN(n11874) );
  NAND2_X1 U14963 ( .A1(n12385), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n11873) );
  INV_X1 U14964 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n11878) );
  OAI21_X1 U14965 ( .B1(n11876), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n11896), .ZN(n19885) );
  AOI22_X1 U14966 ( .A1(n19885), .A2(n13895), .B1(n12318), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n11877) );
  OAI21_X1 U14967 ( .B1(n12043), .B2(n11878), .A(n11877), .ZN(n11879) );
  AOI22_X1 U14968 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12161), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11884) );
  AOI22_X1 U14969 ( .A1(n12233), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11653), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11883) );
  AOI22_X1 U14970 ( .A1(n9628), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11882) );
  AOI22_X1 U14971 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12202), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11881) );
  NAND4_X1 U14972 ( .A1(n11884), .A2(n11883), .A3(n11882), .A4(n11881), .ZN(
        n11890) );
  AOI22_X1 U14973 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9629), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11888) );
  AOI22_X1 U14974 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11887) );
  AOI22_X1 U14975 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11886) );
  AOI22_X1 U14976 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11885) );
  NAND4_X1 U14977 ( .A1(n11888), .A2(n11887), .A3(n11886), .A4(n11885), .ZN(
        n11889) );
  OAI21_X1 U14978 ( .B1(n11890), .B2(n11889), .A(n12003), .ZN(n11894) );
  NAND2_X1 U14979 ( .A1(n12311), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n11893) );
  INV_X1 U14980 ( .A(n11896), .ZN(n11891) );
  XNOR2_X1 U14981 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n11891), .ZN(
        n14155) );
  AOI22_X1 U14982 ( .A1(n13895), .A2(n14155), .B1(n12318), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n11892) );
  XOR2_X1 U14983 ( .A(n11911), .B(n11912), .Z(n14434) );
  INV_X1 U14984 ( .A(n14434), .ZN(n19871) );
  AOI22_X1 U14985 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11900) );
  AOI22_X1 U14986 ( .A1(n12233), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11737), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11899) );
  AOI22_X1 U14987 ( .A1(n9630), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11898) );
  AOI22_X1 U14988 ( .A1(n12161), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11897) );
  NAND4_X1 U14989 ( .A1(n11900), .A2(n11899), .A3(n11898), .A4(n11897), .ZN(
        n11906) );
  AOI22_X1 U14990 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11653), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11904) );
  AOI22_X1 U14991 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11903) );
  AOI22_X1 U14992 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11902) );
  AOI22_X1 U14993 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12202), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11901) );
  NAND4_X1 U14994 ( .A1(n11904), .A2(n11903), .A3(n11902), .A4(n11901), .ZN(
        n11905) );
  OAI21_X1 U14995 ( .B1(n11906), .B2(n11905), .A(n12003), .ZN(n11909) );
  NAND2_X1 U14996 ( .A1(n12311), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n11908) );
  NAND2_X1 U14997 ( .A1(n12318), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11907) );
  NAND3_X1 U14998 ( .A1(n11909), .A2(n11908), .A3(n11907), .ZN(n11910) );
  INV_X1 U14999 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n14957) );
  XNOR2_X1 U15000 ( .A(n11928), .B(n14957), .ZN(n15926) );
  OR2_X1 U15001 ( .A1(n15926), .A2(n12317), .ZN(n11927) );
  AOI22_X1 U15002 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9629), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11916) );
  AOI22_X1 U15003 ( .A1(n12233), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11737), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11915) );
  AOI22_X1 U15004 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11653), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11914) );
  AOI22_X1 U15005 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9624), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11913) );
  NAND4_X1 U15006 ( .A1(n11916), .A2(n11915), .A3(n11914), .A4(n11913), .ZN(
        n11922) );
  AOI22_X1 U15007 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11920) );
  AOI22_X1 U15008 ( .A1(n12161), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11919) );
  AOI22_X1 U15009 ( .A1(n11743), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12202), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11918) );
  AOI22_X1 U15010 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11917) );
  NAND4_X1 U15011 ( .A1(n11920), .A2(n11919), .A3(n11918), .A4(n11917), .ZN(
        n11921) );
  OAI21_X1 U15012 ( .B1(n11922), .B2(n11921), .A(n12003), .ZN(n11925) );
  NAND2_X1 U15013 ( .A1(n12319), .A2(P1_EAX_REG_10__SCAN_IN), .ZN(n11924) );
  NAND2_X1 U15014 ( .A1(n12318), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n11923) );
  AND3_X1 U15015 ( .A1(n11925), .A2(n11924), .A3(n11923), .ZN(n11926) );
  NAND2_X1 U15016 ( .A1(n11927), .A2(n11926), .ZN(n14160) );
  NAND2_X1 U15017 ( .A1(n14094), .A2(n14160), .ZN(n14161) );
  NAND2_X1 U15018 ( .A1(n12319), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n11931) );
  OAI21_X1 U15019 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n11929), .A(
        n11969), .ZN(n16006) );
  AOI22_X1 U15020 ( .A1(n12290), .A2(n16006), .B1(n12318), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n11930) );
  NAND2_X1 U15021 ( .A1(n11931), .A2(n11930), .ZN(n14677) );
  AOI22_X1 U15022 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9629), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11935) );
  AOI22_X1 U15023 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11653), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11934) );
  AOI22_X1 U15024 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11933) );
  AOI22_X1 U15025 ( .A1(n11666), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9608), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11932) );
  NAND4_X1 U15026 ( .A1(n11935), .A2(n11934), .A3(n11933), .A4(n11932), .ZN(
        n11941) );
  AOI22_X1 U15027 ( .A1(n12233), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11939) );
  AOI22_X1 U15028 ( .A1(n12161), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11938) );
  AOI22_X1 U15029 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11937) );
  AOI22_X1 U15030 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11936) );
  NAND4_X1 U15031 ( .A1(n11939), .A2(n11938), .A3(n11937), .A4(n11936), .ZN(
        n11940) );
  OR2_X1 U15032 ( .A1(n11941), .A2(n11940), .ZN(n11942) );
  AND2_X1 U15033 ( .A1(n12003), .A2(n11942), .ZN(n14313) );
  AOI22_X1 U15034 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12233), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11946) );
  AOI22_X1 U15035 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11653), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11945) );
  AOI22_X1 U15036 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12161), .B1(
        n9624), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11944) );
  AOI22_X1 U15037 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n9627), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11943) );
  NAND4_X1 U15038 ( .A1(n11946), .A2(n11945), .A3(n11944), .A4(n11943), .ZN(
        n11952) );
  AOI22_X1 U15039 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11950) );
  AOI22_X1 U15040 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12278), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11949) );
  AOI22_X1 U15041 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12202), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11948) );
  AOI22_X1 U15042 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12295), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11947) );
  NAND4_X1 U15043 ( .A1(n11950), .A2(n11949), .A3(n11948), .A4(n11947), .ZN(
        n11951) );
  NOR2_X1 U15044 ( .A1(n11952), .A2(n11951), .ZN(n11958) );
  XNOR2_X1 U15045 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n11969), .ZN(
        n15999) );
  INV_X1 U15046 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n11953) );
  OAI22_X1 U15047 ( .A1(n15999), .A2(n12317), .B1(n11954), .B2(n11953), .ZN(
        n11955) );
  INV_X1 U15048 ( .A(n11955), .ZN(n11957) );
  NAND2_X1 U15049 ( .A1(n12311), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n11956) );
  OAI211_X1 U15050 ( .C1(n11975), .C2(n11958), .A(n11957), .B(n11956), .ZN(
        n14679) );
  AOI22_X1 U15051 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11962) );
  AOI22_X1 U15052 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9629), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11961) );
  AOI22_X1 U15053 ( .A1(n11737), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11960) );
  AOI22_X1 U15054 ( .A1(n12161), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11959) );
  NAND4_X1 U15055 ( .A1(n11962), .A2(n11961), .A3(n11960), .A4(n11959), .ZN(
        n11968) );
  AOI22_X1 U15056 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12233), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11966) );
  AOI22_X1 U15057 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11965) );
  AOI22_X1 U15058 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11964) );
  AOI22_X1 U15059 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9608), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11963) );
  NAND4_X1 U15060 ( .A1(n11966), .A2(n11965), .A3(n11964), .A4(n11963), .ZN(
        n11967) );
  NOR2_X1 U15061 ( .A1(n11968), .A2(n11967), .ZN(n11974) );
  INV_X1 U15062 ( .A(n11978), .ZN(n11971) );
  XNOR2_X1 U15063 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n11971), .ZN(
        n14948) );
  AOI22_X1 U15064 ( .A1(n13895), .A2(n14948), .B1(n12318), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n11973) );
  NAND2_X1 U15065 ( .A1(n12311), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n11972) );
  OAI211_X1 U15066 ( .C1(n11975), .C2(n11974), .A(n11973), .B(n11972), .ZN(
        n14681) );
  OAI211_X1 U15067 ( .C1(n14677), .C2(n14313), .A(n14679), .B(n14681), .ZN(
        n11976) );
  XOR2_X1 U15068 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B(n11994), .Z(
        n15990) );
  INV_X1 U15069 ( .A(n15990), .ZN(n11993) );
  AOI22_X1 U15070 ( .A1(n12161), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11982) );
  AOI22_X1 U15071 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9630), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11981) );
  AOI22_X1 U15072 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11980) );
  AOI22_X1 U15073 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11492), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11979) );
  NAND4_X1 U15074 ( .A1(n11982), .A2(n11981), .A3(n11980), .A4(n11979), .ZN(
        n11988) );
  AOI22_X1 U15075 ( .A1(n11666), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11653), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11986) );
  AOI22_X1 U15076 ( .A1(n12233), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11743), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11985) );
  AOI22_X1 U15077 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11984) );
  AOI22_X1 U15078 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11983) );
  NAND4_X1 U15079 ( .A1(n11986), .A2(n11985), .A3(n11984), .A4(n11983), .ZN(
        n11987) );
  OAI21_X1 U15080 ( .B1(n11988), .B2(n11987), .A(n12003), .ZN(n11991) );
  NAND2_X1 U15081 ( .A1(n12311), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n11990) );
  NAND2_X1 U15082 ( .A1(n12318), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11989) );
  NAND3_X1 U15083 ( .A1(n11991), .A2(n11990), .A3(n11989), .ZN(n11992) );
  AOI21_X1 U15084 ( .B1(n11993), .B2(n13895), .A(n11992), .ZN(n14285) );
  NOR2_X2 U15085 ( .A1(n14680), .A2(n14285), .ZN(n14327) );
  XNOR2_X1 U15086 ( .A(n12027), .B(n12026), .ZN(n14935) );
  NAND2_X1 U15087 ( .A1(n14935), .A2(n12290), .ZN(n12010) );
  AOI22_X1 U15088 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11998) );
  AOI22_X1 U15089 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11743), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11997) );
  AOI22_X1 U15090 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11996) );
  AOI22_X1 U15091 ( .A1(n12233), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11492), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11995) );
  NAND4_X1 U15092 ( .A1(n11998), .A2(n11997), .A3(n11996), .A4(n11995), .ZN(
        n12005) );
  AOI22_X1 U15093 ( .A1(n12161), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12002) );
  AOI22_X1 U15094 ( .A1(n9629), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12001) );
  AOI22_X1 U15095 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9624), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12000) );
  AOI22_X1 U15096 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11999) );
  NAND4_X1 U15097 ( .A1(n12002), .A2(n12001), .A3(n12000), .A4(n11999), .ZN(
        n12004) );
  OAI21_X1 U15098 ( .B1(n12005), .B2(n12004), .A(n12003), .ZN(n12008) );
  NAND2_X1 U15099 ( .A1(n12311), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12007) );
  NAND2_X1 U15100 ( .A1(n12318), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12006) );
  AND3_X1 U15101 ( .A1(n12008), .A2(n12007), .A3(n12006), .ZN(n12009) );
  NAND2_X1 U15102 ( .A1(n12010), .A2(n12009), .ZN(n14326) );
  AND2_X2 U15103 ( .A1(n14327), .A2(n14326), .ZN(n14358) );
  INV_X1 U15104 ( .A(n11634), .ZN(n12011) );
  AOI22_X1 U15105 ( .A1(n12161), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12015) );
  AOI22_X1 U15106 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12014) );
  AOI22_X1 U15107 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12013) );
  AOI22_X1 U15108 ( .A1(n12233), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12012) );
  NAND4_X1 U15109 ( .A1(n12015), .A2(n12014), .A3(n12013), .A4(n12012), .ZN(
        n12021) );
  AOI22_X1 U15110 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9630), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12019) );
  AOI22_X1 U15111 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U15112 ( .A1(n11666), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9608), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12017) );
  AOI22_X1 U15113 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12016) );
  NAND4_X1 U15114 ( .A1(n12019), .A2(n12018), .A3(n12017), .A4(n12016), .ZN(
        n12020) );
  NOR2_X1 U15115 ( .A1(n12021), .A2(n12020), .ZN(n12025) );
  NAND2_X1 U15116 ( .A1(n20752), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12022) );
  NAND2_X1 U15117 ( .A1(n12317), .A2(n12022), .ZN(n12023) );
  AOI21_X1 U15118 ( .B1(n12311), .B2(P1_EAX_REG_16__SCAN_IN), .A(n12023), .ZN(
        n12024) );
  OAI21_X1 U15119 ( .B1(n12314), .B2(n12025), .A(n12024), .ZN(n12030) );
  OAI21_X1 U15120 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12028), .A(
        n12060), .ZN(n15984) );
  OR2_X1 U15121 ( .A1(n12317), .A2(n15984), .ZN(n12029) );
  AOI22_X1 U15122 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12233), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12034) );
  AOI22_X1 U15123 ( .A1(n12161), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12033) );
  AOI22_X1 U15124 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12032) );
  AOI22_X1 U15125 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12031) );
  NAND4_X1 U15126 ( .A1(n12034), .A2(n12033), .A3(n12032), .A4(n12031), .ZN(
        n12040) );
  AOI22_X1 U15127 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11653), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12038) );
  AOI22_X1 U15128 ( .A1(n9629), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11743), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12037) );
  AOI22_X1 U15129 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9624), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12036) );
  AOI22_X1 U15130 ( .A1(n11737), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9608), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12035) );
  NAND4_X1 U15131 ( .A1(n12038), .A2(n12037), .A3(n12036), .A4(n12035), .ZN(
        n12039) );
  OR2_X1 U15132 ( .A1(n12040), .A2(n12039), .ZN(n12045) );
  INV_X1 U15133 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n14816) );
  INV_X1 U15134 ( .A(n12060), .ZN(n12041) );
  XNOR2_X1 U15135 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12041), .ZN(
        n15890) );
  AOI22_X1 U15136 ( .A1(n12290), .A2(n15890), .B1(n12318), .B2(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12042) );
  OAI21_X1 U15137 ( .B1(n12043), .B2(n14816), .A(n12042), .ZN(n12044) );
  AOI21_X1 U15138 ( .B1(n12287), .B2(n12045), .A(n12044), .ZN(n14753) );
  AOI22_X1 U15139 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12049) );
  AOI22_X1 U15140 ( .A1(n12233), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9629), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12048) );
  AOI22_X1 U15141 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11653), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12047) );
  AOI22_X1 U15142 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12046) );
  NAND4_X1 U15143 ( .A1(n12049), .A2(n12048), .A3(n12047), .A4(n12046), .ZN(
        n12055) );
  AOI22_X1 U15144 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9627), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12053) );
  AOI22_X1 U15145 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12052) );
  AOI22_X1 U15146 ( .A1(n12161), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12051) );
  AOI22_X1 U15147 ( .A1(n11666), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11492), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12050) );
  NAND4_X1 U15148 ( .A1(n12053), .A2(n12052), .A3(n12051), .A4(n12050), .ZN(
        n12054) );
  NOR2_X1 U15149 ( .A1(n12055), .A2(n12054), .ZN(n12059) );
  NAND2_X1 U15150 ( .A1(n20752), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12056) );
  NAND2_X1 U15151 ( .A1(n12317), .A2(n12056), .ZN(n12057) );
  AOI21_X1 U15152 ( .B1(n12311), .B2(P1_EAX_REG_18__SCAN_IN), .A(n12057), .ZN(
        n12058) );
  OAI21_X1 U15153 ( .B1(n12314), .B2(n12059), .A(n12058), .ZN(n12065) );
  INV_X1 U15154 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14908) );
  INV_X1 U15155 ( .A(n12062), .ZN(n12061) );
  NAND2_X1 U15156 ( .A1(n14908), .A2(n12061), .ZN(n12063) );
  AND2_X1 U15157 ( .A1(n12063), .A2(n12114), .ZN(n15886) );
  NAND2_X1 U15158 ( .A1(n15886), .A2(n12290), .ZN(n12064) );
  NAND2_X1 U15159 ( .A1(n12065), .A2(n12064), .ZN(n14747) );
  AOI22_X1 U15160 ( .A1(n12161), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U15161 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12068) );
  AOI22_X1 U15162 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12067) );
  AOI22_X1 U15163 ( .A1(n11743), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11492), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12066) );
  NAND4_X1 U15164 ( .A1(n12069), .A2(n12068), .A3(n12067), .A4(n12066), .ZN(
        n12075) );
  AOI22_X1 U15165 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9630), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12073) );
  AOI22_X1 U15166 ( .A1(n12233), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11653), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12072) );
  AOI22_X1 U15167 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12071) );
  AOI22_X1 U15168 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12070) );
  NAND4_X1 U15169 ( .A1(n12073), .A2(n12072), .A3(n12071), .A4(n12070), .ZN(
        n12074) );
  NOR2_X1 U15170 ( .A1(n12075), .A2(n12074), .ZN(n12078) );
  AOI21_X1 U15171 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n14900), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12076) );
  AOI21_X1 U15172 ( .B1(n12311), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12076), .ZN(
        n12077) );
  OAI21_X1 U15173 ( .B1(n12314), .B2(n12078), .A(n12077), .ZN(n12080) );
  XNOR2_X1 U15174 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B(n12114), .ZN(
        n15867) );
  NAND2_X1 U15175 ( .A1(n12290), .A2(n15867), .ZN(n12079) );
  AOI22_X1 U15176 ( .A1(n12161), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12084) );
  AOI22_X1 U15177 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12083) );
  AOI22_X1 U15178 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12082) );
  AOI22_X1 U15179 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12081) );
  NAND4_X1 U15180 ( .A1(n12084), .A2(n12083), .A3(n12082), .A4(n12081), .ZN(
        n12090) );
  AOI22_X1 U15181 ( .A1(n12233), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11737), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12088) );
  AOI22_X1 U15182 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11653), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12087) );
  AOI22_X1 U15183 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11743), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12086) );
  AOI22_X1 U15184 ( .A1(n12278), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9608), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12085) );
  NAND4_X1 U15185 ( .A1(n12088), .A2(n12087), .A3(n12086), .A4(n12085), .ZN(
        n12089) );
  NOR2_X1 U15186 ( .A1(n12090), .A2(n12089), .ZN(n12120) );
  AOI22_X1 U15187 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12094) );
  AOI22_X1 U15188 ( .A1(n11513), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11653), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12093) );
  AOI22_X1 U15189 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9608), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12092) );
  AOI22_X1 U15190 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12091) );
  NAND4_X1 U15191 ( .A1(n12094), .A2(n12093), .A3(n12092), .A4(n12091), .ZN(
        n12100) );
  AOI22_X1 U15192 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9629), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12098) );
  AOI22_X1 U15193 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12097) );
  AOI22_X1 U15194 ( .A1(n12161), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12096) );
  AOI22_X1 U15195 ( .A1(n9628), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12095) );
  NAND4_X1 U15196 ( .A1(n12098), .A2(n12097), .A3(n12096), .A4(n12095), .ZN(
        n12099) );
  NOR2_X1 U15197 ( .A1(n12100), .A2(n12099), .ZN(n12119) );
  NOR2_X1 U15198 ( .A1(n12120), .A2(n12119), .ZN(n12183) );
  AOI22_X1 U15199 ( .A1(n11513), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12104) );
  AOI22_X1 U15200 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11653), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12103) );
  AOI22_X1 U15201 ( .A1(n9629), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(n9608), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U15202 ( .A1(n12249), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12101) );
  NAND4_X1 U15203 ( .A1(n12104), .A2(n12103), .A3(n12102), .A4(n12101), .ZN(
        n12110) );
  AOI22_X1 U15204 ( .A1(n12161), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12108) );
  AOI22_X1 U15205 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11743), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12107) );
  AOI22_X1 U15206 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12106) );
  AOI22_X1 U15207 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12105) );
  NAND4_X1 U15208 ( .A1(n12108), .A2(n12107), .A3(n12106), .A4(n12105), .ZN(
        n12109) );
  OR2_X1 U15209 ( .A1(n12110), .A2(n12109), .ZN(n12182) );
  INV_X1 U15210 ( .A(n12182), .ZN(n12111) );
  XNOR2_X1 U15211 ( .A(n12183), .B(n12111), .ZN(n12112) );
  NAND2_X1 U15212 ( .A1(n12112), .A2(n12287), .ZN(n12118) );
  INV_X1 U15213 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n15814) );
  AOI21_X1 U15214 ( .B1(n15814), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12113) );
  AOI21_X1 U15215 ( .B1(n12311), .B2(P1_EAX_REG_24__SCAN_IN), .A(n12113), .ZN(
        n12117) );
  INV_X1 U15216 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15823) );
  OAI21_X1 U15217 ( .B1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n12115), .A(
        n12218), .ZN(n15960) );
  NOR2_X1 U15218 ( .A1(n12317), .A2(n15960), .ZN(n12116) );
  AOI21_X1 U15219 ( .B1(n12118), .B2(n12117), .A(n12116), .ZN(n14711) );
  INV_X1 U15220 ( .A(n14711), .ZN(n12160) );
  XNOR2_X1 U15221 ( .A(n12120), .B(n12119), .ZN(n12123) );
  OAI21_X1 U15222 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n15823), .A(n12317), 
        .ZN(n12121) );
  AOI21_X1 U15223 ( .B1(n12311), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12121), .ZN(
        n12122) );
  OAI21_X1 U15224 ( .B1(n12123), .B2(n12314), .A(n12122), .ZN(n12125) );
  XNOR2_X1 U15225 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B(n12140), .ZN(
        n15832) );
  NAND2_X1 U15226 ( .A1(n15832), .A2(n12290), .ZN(n12124) );
  INV_X1 U15227 ( .A(n14720), .ZN(n12159) );
  AOI22_X1 U15228 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12129) );
  AOI22_X1 U15229 ( .A1(n11593), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12128) );
  AOI22_X1 U15230 ( .A1(n9630), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11743), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12127) );
  AOI22_X1 U15231 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12126) );
  NAND4_X1 U15232 ( .A1(n12129), .A2(n12128), .A3(n12127), .A4(n12126), .ZN(
        n12135) );
  AOI22_X1 U15233 ( .A1(n12233), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11653), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12133) );
  AOI22_X1 U15234 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12132) );
  AOI22_X1 U15235 ( .A1(n12161), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12131) );
  AOI22_X1 U15236 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9608), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12130) );
  NAND4_X1 U15237 ( .A1(n12133), .A2(n12132), .A3(n12131), .A4(n12130), .ZN(
        n12134) );
  NOR2_X1 U15238 ( .A1(n12135), .A2(n12134), .ZN(n12139) );
  NAND2_X1 U15239 ( .A1(n20752), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12136) );
  NAND2_X1 U15240 ( .A1(n12317), .A2(n12136), .ZN(n12137) );
  AOI21_X1 U15241 ( .B1(n12311), .B2(P1_EAX_REG_22__SCAN_IN), .A(n12137), .ZN(
        n12138) );
  OAI21_X1 U15242 ( .B1(n12314), .B2(n12139), .A(n12138), .ZN(n12143) );
  OAI21_X1 U15243 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12141), .A(
        n12140), .ZN(n15967) );
  OR2_X1 U15244 ( .A1(n12317), .A2(n15967), .ZN(n12142) );
  NAND2_X1 U15245 ( .A1(n12143), .A2(n12142), .ZN(n14727) );
  AOI22_X1 U15246 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12147) );
  AOI22_X1 U15247 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11653), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12146) );
  AOI22_X1 U15248 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12145) );
  AOI22_X1 U15249 ( .A1(n12233), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9608), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12144) );
  NAND4_X1 U15250 ( .A1(n12147), .A2(n12146), .A3(n12145), .A4(n12144), .ZN(
        n12153) );
  AOI22_X1 U15251 ( .A1(n12278), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12151) );
  AOI22_X1 U15252 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12150) );
  AOI22_X1 U15253 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12149) );
  AOI22_X1 U15254 ( .A1(n12161), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12148) );
  NAND4_X1 U15255 ( .A1(n12151), .A2(n12150), .A3(n12149), .A4(n12148), .ZN(
        n12152) );
  NOR2_X1 U15256 ( .A1(n12153), .A2(n12152), .ZN(n12156) );
  AOI21_X1 U15257 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15845), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12154) );
  AOI21_X1 U15258 ( .B1(n12311), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12154), .ZN(
        n12155) );
  OAI21_X1 U15259 ( .B1(n12314), .B2(n12156), .A(n12155), .ZN(n12158) );
  XNOR2_X1 U15260 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n12176), .ZN(
        n15844) );
  NAND2_X1 U15261 ( .A1(n15844), .A2(n12290), .ZN(n12157) );
  NAND2_X1 U15262 ( .A1(n12158), .A2(n12157), .ZN(n14732) );
  AOI22_X1 U15263 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12228), .B1(
        n12233), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12165) );
  AOI22_X1 U15264 ( .A1(n12161), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12164) );
  AOI22_X1 U15265 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12163) );
  AOI22_X1 U15266 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11492), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12162) );
  NAND4_X1 U15267 ( .A1(n12165), .A2(n12164), .A3(n12163), .A4(n12162), .ZN(
        n12171) );
  AOI22_X1 U15268 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12294), .B1(
        n12278), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12169) );
  AOI22_X1 U15269 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n11738), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12168) );
  AOI22_X1 U15270 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9624), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12167) );
  AOI22_X1 U15271 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n11690), .B1(
        n12249), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12166) );
  NAND4_X1 U15272 ( .A1(n12169), .A2(n12168), .A3(n12167), .A4(n12166), .ZN(
        n12170) );
  NOR2_X1 U15273 ( .A1(n12171), .A2(n12170), .ZN(n12175) );
  OAI21_X1 U15274 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20753), .A(
        n20752), .ZN(n12172) );
  INV_X1 U15275 ( .A(n12172), .ZN(n12173) );
  AOI21_X1 U15276 ( .B1(n12311), .B2(P1_EAX_REG_20__SCAN_IN), .A(n12173), .ZN(
        n12174) );
  OAI21_X1 U15277 ( .B1(n12314), .B2(n12175), .A(n12174), .ZN(n12179) );
  OAI21_X1 U15278 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12177), .A(
        n12176), .ZN(n15853) );
  INV_X1 U15279 ( .A(n15853), .ZN(n15968) );
  NAND2_X1 U15280 ( .A1(n15968), .A2(n12290), .ZN(n12178) );
  NAND2_X1 U15281 ( .A1(n12179), .A2(n12178), .ZN(n15858) );
  NAND2_X1 U15282 ( .A1(n12183), .A2(n12182), .ZN(n12200) );
  AOI22_X1 U15283 ( .A1(n11513), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11666), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12187) );
  AOI22_X1 U15284 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12186) );
  AOI22_X1 U15285 ( .A1(n12249), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12185) );
  AOI22_X1 U15286 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9624), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12184) );
  NAND4_X1 U15287 ( .A1(n12187), .A2(n12186), .A3(n12185), .A4(n12184), .ZN(
        n12193) );
  AOI22_X1 U15288 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12161), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12191) );
  AOI22_X1 U15289 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12190) );
  AOI22_X1 U15290 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U15291 ( .A1(n12278), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9608), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12188) );
  NAND4_X1 U15292 ( .A1(n12191), .A2(n12190), .A3(n12189), .A4(n12188), .ZN(
        n12192) );
  NOR2_X1 U15293 ( .A1(n12193), .A2(n12192), .ZN(n12201) );
  XOR2_X1 U15294 ( .A(n12200), .B(n12201), .Z(n12194) );
  NAND2_X1 U15295 ( .A1(n12194), .A2(n12287), .ZN(n12199) );
  NAND2_X1 U15296 ( .A1(n20752), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12195) );
  NAND2_X1 U15297 ( .A1(n12317), .A2(n12195), .ZN(n12196) );
  AOI21_X1 U15298 ( .B1(n12311), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12196), .ZN(
        n12198) );
  XNOR2_X1 U15299 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B(n12218), .ZN(
        n14882) );
  AOI21_X1 U15300 ( .B1(n12199), .B2(n12198), .A(n12197), .ZN(n14663) );
  NAND2_X1 U15301 ( .A1(n14662), .A2(n14663), .ZN(n14650) );
  NOR2_X1 U15302 ( .A1(n12201), .A2(n12200), .ZN(n12227) );
  AOI22_X1 U15303 ( .A1(n11513), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11737), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12206) );
  AOI22_X1 U15304 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12205) );
  AOI22_X1 U15305 ( .A1(n9629), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11492), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12204) );
  AOI22_X1 U15306 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12203) );
  NAND4_X1 U15307 ( .A1(n12206), .A2(n12205), .A3(n12204), .A4(n12203), .ZN(
        n12213) );
  AOI22_X1 U15308 ( .A1(n11602), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12211) );
  AOI22_X1 U15309 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11743), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U15310 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12209) );
  AOI22_X1 U15311 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12208) );
  NAND4_X1 U15312 ( .A1(n12211), .A2(n12210), .A3(n12209), .A4(n12208), .ZN(
        n12212) );
  OR2_X1 U15313 ( .A1(n12213), .A2(n12212), .ZN(n12226) );
  INV_X1 U15314 ( .A(n12226), .ZN(n12214) );
  XNOR2_X1 U15315 ( .A(n12227), .B(n12214), .ZN(n12217) );
  INV_X1 U15316 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14653) );
  NAND2_X1 U15317 ( .A1(n12311), .A2(P1_EAX_REG_26__SCAN_IN), .ZN(n12215) );
  OAI211_X1 U15318 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n14653), .A(n12215), 
        .B(n12317), .ZN(n12216) );
  AOI21_X1 U15319 ( .B1(n12217), .B2(n12287), .A(n12216), .ZN(n12224) );
  INV_X1 U15320 ( .A(n12218), .ZN(n12219) );
  INV_X1 U15321 ( .A(n12220), .ZN(n12221) );
  NAND2_X1 U15322 ( .A1(n12221), .A2(n14653), .ZN(n12222) );
  NAND2_X1 U15323 ( .A1(n12265), .A2(n12222), .ZN(n14872) );
  NOR2_X1 U15324 ( .A1(n14872), .A2(n12317), .ZN(n12223) );
  NOR2_X2 U15325 ( .A1(n14650), .A2(n14652), .ZN(n12225) );
  INV_X1 U15326 ( .A(n12225), .ZN(n14636) );
  NAND2_X1 U15327 ( .A1(n12227), .A2(n12226), .ZN(n12247) );
  AOI22_X1 U15328 ( .A1(n11602), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12232) );
  AOI22_X1 U15329 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12228), .B1(
        n11653), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12231) );
  AOI22_X1 U15330 ( .A1(n11743), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11492), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12230) );
  AOI22_X1 U15331 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n11690), .B1(
        n12249), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12229) );
  NAND4_X1 U15332 ( .A1(n12232), .A2(n12231), .A3(n12230), .A4(n12229), .ZN(
        n12239) );
  AOI22_X1 U15333 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9629), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12237) );
  AOI22_X1 U15334 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12233), .B1(
        n11737), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12236) );
  AOI22_X1 U15335 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12235) );
  AOI22_X1 U15336 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n12300), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12234) );
  NAND4_X1 U15337 ( .A1(n12237), .A2(n12236), .A3(n12235), .A4(n12234), .ZN(
        n12238) );
  NOR2_X1 U15338 ( .A1(n12239), .A2(n12238), .ZN(n12248) );
  XOR2_X1 U15339 ( .A(n12247), .B(n12248), .Z(n12240) );
  NAND2_X1 U15340 ( .A1(n12240), .A2(n12287), .ZN(n12244) );
  NAND2_X1 U15341 ( .A1(n20752), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12241) );
  NAND2_X1 U15342 ( .A1(n12317), .A2(n12241), .ZN(n12242) );
  AOI21_X1 U15343 ( .B1(n12311), .B2(P1_EAX_REG_27__SCAN_IN), .A(n12242), .ZN(
        n12243) );
  NAND2_X1 U15344 ( .A1(n12244), .A2(n12243), .ZN(n12246) );
  XNOR2_X1 U15345 ( .A(n12265), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14862) );
  NAND2_X1 U15346 ( .A1(n14862), .A2(n13895), .ZN(n12245) );
  NAND2_X1 U15347 ( .A1(n12246), .A2(n12245), .ZN(n14637) );
  NOR2_X1 U15348 ( .A1(n12248), .A2(n12247), .ZN(n12273) );
  AOI22_X1 U15349 ( .A1(n11513), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11737), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U15350 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12252) );
  AOI22_X1 U15351 ( .A1(n9629), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11492), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12251) );
  AOI22_X1 U15352 ( .A1(n12249), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12250) );
  NAND4_X1 U15353 ( .A1(n12253), .A2(n12252), .A3(n12251), .A4(n12250), .ZN(
        n12260) );
  AOI22_X1 U15354 ( .A1(n11602), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12258) );
  AOI22_X1 U15355 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9627), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12257) );
  AOI22_X1 U15356 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12256) );
  AOI22_X1 U15357 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12255) );
  NAND4_X1 U15358 ( .A1(n12258), .A2(n12257), .A3(n12256), .A4(n12255), .ZN(
        n12259) );
  OR2_X1 U15359 ( .A1(n12260), .A2(n12259), .ZN(n12272) );
  INV_X1 U15360 ( .A(n12272), .ZN(n12261) );
  XNOR2_X1 U15361 ( .A(n12273), .B(n12261), .ZN(n12262) );
  NAND2_X1 U15362 ( .A1(n12262), .A2(n12287), .ZN(n12271) );
  NAND2_X1 U15363 ( .A1(n20752), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12263) );
  NAND2_X1 U15364 ( .A1(n12317), .A2(n12263), .ZN(n12264) );
  AOI21_X1 U15365 ( .B1(n12311), .B2(P1_EAX_REG_28__SCAN_IN), .A(n12264), .ZN(
        n12270) );
  INV_X1 U15366 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14864) );
  NAND2_X1 U15367 ( .A1(n12266), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12291) );
  INV_X1 U15368 ( .A(n12266), .ZN(n12267) );
  INV_X1 U15369 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14626) );
  NAND2_X1 U15370 ( .A1(n12267), .A2(n14626), .ZN(n12268) );
  NAND2_X1 U15371 ( .A1(n12291), .A2(n12268), .ZN(n14855) );
  NOR2_X1 U15372 ( .A1(n14855), .A2(n12317), .ZN(n12269) );
  AOI21_X1 U15373 ( .B1(n12271), .B2(n12270), .A(n12269), .ZN(n14622) );
  XNOR2_X1 U15374 ( .A(n12291), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14839) );
  NAND2_X1 U15375 ( .A1(n12273), .A2(n12272), .ZN(n12307) );
  AOI22_X1 U15376 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12300), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12277) );
  AOI22_X1 U15377 ( .A1(n11602), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12276) );
  AOI22_X1 U15378 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9627), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12275) );
  AOI22_X1 U15379 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12274) );
  NAND4_X1 U15380 ( .A1(n12277), .A2(n12276), .A3(n12275), .A4(n12274), .ZN(
        n12284) );
  AOI22_X1 U15381 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12278), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12282) );
  AOI22_X1 U15382 ( .A1(n11666), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11653), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12281) );
  AOI22_X1 U15383 ( .A1(n12207), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11659), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12280) );
  AOI22_X1 U15384 ( .A1(n11513), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11492), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12279) );
  NAND4_X1 U15385 ( .A1(n12282), .A2(n12281), .A3(n12280), .A4(n12279), .ZN(
        n12283) );
  NOR2_X1 U15386 ( .A1(n12284), .A2(n12283), .ZN(n12308) );
  XOR2_X1 U15387 ( .A(n12307), .B(n12308), .Z(n12288) );
  INV_X1 U15388 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14837) );
  NAND2_X1 U15389 ( .A1(n12311), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n12285) );
  OAI211_X1 U15390 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n14837), .A(n12285), 
        .B(n12317), .ZN(n12286) );
  AOI21_X1 U15391 ( .B1(n12288), .B2(n12287), .A(n12286), .ZN(n12289) );
  AOI21_X1 U15392 ( .B1(n12290), .B2(n14839), .A(n12289), .ZN(n14609) );
  INV_X1 U15393 ( .A(n12291), .ZN(n12292) );
  XNOR2_X1 U15394 ( .A(n13899), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14833) );
  AOI22_X1 U15395 ( .A1(n12254), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12161), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12299) );
  AOI22_X1 U15396 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12233), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U15397 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12297) );
  AOI22_X1 U15398 ( .A1(n12295), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11690), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12296) );
  NAND4_X1 U15399 ( .A1(n12299), .A2(n12298), .A3(n12297), .A4(n12296), .ZN(
        n12306) );
  AOI22_X1 U15400 ( .A1(n12228), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11738), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12304) );
  AOI22_X1 U15401 ( .A1(n12300), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9624), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12303) );
  AOI22_X1 U15402 ( .A1(n9630), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12207), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12302) );
  AOI22_X1 U15403 ( .A1(n11666), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11492), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12301) );
  NAND4_X1 U15404 ( .A1(n12304), .A2(n12303), .A3(n12302), .A4(n12301), .ZN(
        n12305) );
  NOR2_X1 U15405 ( .A1(n12306), .A2(n12305), .ZN(n12310) );
  NOR2_X1 U15406 ( .A1(n12308), .A2(n12307), .ZN(n12309) );
  XOR2_X1 U15407 ( .A(n12310), .B(n12309), .Z(n12315) );
  AOI21_X1 U15408 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20752), .A(
        n13895), .ZN(n12313) );
  NAND2_X1 U15409 ( .A1(n12311), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n12312) );
  OAI211_X1 U15410 ( .C1(n12315), .C2(n12314), .A(n12313), .B(n12312), .ZN(
        n12316) );
  OAI21_X1 U15411 ( .B1(n12317), .B2(n14833), .A(n12316), .ZN(n14481) );
  AOI22_X1 U15412 ( .A1(n12319), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12318), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12320) );
  INV_X1 U15413 ( .A(n12321), .ZN(n12340) );
  XNOR2_X1 U15414 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n12336) );
  NAND2_X1 U15415 ( .A1(n20519), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n12355) );
  NAND2_X1 U15416 ( .A1(n12336), .A2(n12337), .ZN(n12323) );
  NAND2_X1 U15417 ( .A1(n20424), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12322) );
  NAND2_X1 U15418 ( .A1(n12323), .A2(n12322), .ZN(n12335) );
  XNOR2_X1 U15419 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n12334) );
  NAND2_X1 U15420 ( .A1(n12335), .A2(n12334), .ZN(n12325) );
  NAND2_X1 U15421 ( .A1(n20488), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12324) );
  NAND2_X1 U15422 ( .A1(n12325), .A2(n12324), .ZN(n12333) );
  XNOR2_X1 U15423 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12332) );
  NAND2_X1 U15424 ( .A1(n12333), .A2(n12332), .ZN(n12327) );
  NAND2_X1 U15425 ( .A1(n20738), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12326) );
  NOR2_X1 U15426 ( .A1(n16154), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n12328) );
  XNOR2_X1 U15427 ( .A(n12333), .B(n12332), .ZN(n12376) );
  XNOR2_X1 U15428 ( .A(n12335), .B(n12334), .ZN(n12370) );
  XNOR2_X1 U15429 ( .A(n12337), .B(n12336), .ZN(n12363) );
  NOR4_X1 U15430 ( .A1(n12383), .A2(n12376), .A3(n12370), .A4(n12363), .ZN(
        n12338) );
  NOR2_X1 U15431 ( .A1(n12351), .A2(n12338), .ZN(n14581) );
  NAND2_X1 U15432 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n20760) );
  AND2_X1 U15433 ( .A1(n14581), .A2(n20760), .ZN(n12339) );
  NAND2_X1 U15434 ( .A1(n12340), .A2(n12339), .ZN(n13363) );
  INV_X1 U15435 ( .A(n13349), .ZN(n12342) );
  AND3_X1 U15436 ( .A1(n20141), .A2(n11626), .A3(n12341), .ZN(n13313) );
  NAND2_X1 U15437 ( .A1(n12342), .A2(n13313), .ZN(n12343) );
  NAND2_X1 U15438 ( .A1(n13363), .A2(n12343), .ZN(n12344) );
  NAND2_X1 U15439 ( .A1(n12344), .A2(n14598), .ZN(n12394) );
  OR2_X1 U15440 ( .A1(n11633), .A2(n11569), .ZN(n12346) );
  AND2_X1 U15441 ( .A1(n12346), .A2(n12345), .ZN(n13274) );
  NAND2_X1 U15442 ( .A1(n11634), .A2(n20105), .ZN(n12347) );
  NAND3_X1 U15443 ( .A1(n13274), .A2(n13395), .A3(n12347), .ZN(n13401) );
  INV_X1 U15444 ( .A(n13401), .ZN(n13266) );
  INV_X1 U15445 ( .A(n14588), .ZN(n13904) );
  NAND2_X1 U15446 ( .A1(n13266), .A2(n13904), .ZN(n13373) );
  INV_X1 U15447 ( .A(n20760), .ZN(n20674) );
  OR2_X1 U15448 ( .A1(n12348), .A2(n20674), .ZN(n12349) );
  NAND2_X1 U15449 ( .A1(n13373), .A2(n12349), .ZN(n13367) );
  INV_X1 U15450 ( .A(n12351), .ZN(n12350) );
  NAND2_X1 U15451 ( .A1(n12351), .A2(n12357), .ZN(n12390) );
  INV_X1 U15452 ( .A(n12385), .ZN(n12375) );
  NAND2_X1 U15453 ( .A1(n12357), .A2(n13907), .ZN(n12353) );
  NAND2_X1 U15454 ( .A1(n11630), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12352) );
  NOR2_X1 U15455 ( .A1(n12363), .A2(n12362), .ZN(n12361) );
  NAND2_X1 U15456 ( .A1(n11630), .A2(n14596), .ZN(n12354) );
  NAND2_X1 U15457 ( .A1(n12354), .A2(n20120), .ZN(n12371) );
  OAI21_X1 U15458 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20519), .A(
        n12355), .ZN(n12358) );
  INV_X1 U15459 ( .A(n12358), .ZN(n12356) );
  OAI211_X1 U15460 ( .C1(n20105), .C2(n13400), .A(n12371), .B(n12356), .ZN(
        n12360) );
  INV_X1 U15461 ( .A(n12357), .ZN(n12372) );
  OAI21_X1 U15462 ( .B1(n12372), .B2(n12358), .A(n12377), .ZN(n12359) );
  NAND2_X1 U15463 ( .A1(n12360), .A2(n12359), .ZN(n12364) );
  NAND2_X1 U15464 ( .A1(n12361), .A2(n12364), .ZN(n12369) );
  INV_X1 U15465 ( .A(n12362), .ZN(n12365) );
  OAI211_X1 U15466 ( .C1(n12365), .C2(n12364), .A(n12363), .B(n12382), .ZN(
        n12368) );
  NAND2_X1 U15467 ( .A1(n12385), .A2(n12370), .ZN(n12366) );
  OAI211_X1 U15468 ( .C1(n12372), .C2(n12370), .A(n12366), .B(n12371), .ZN(
        n12367) );
  NAND3_X1 U15469 ( .A1(n12369), .A2(n12368), .A3(n12367), .ZN(n12374) );
  AOI22_X1 U15470 ( .A1(n12375), .A2(n12376), .B1(n12374), .B2(n12373), .ZN(
        n12381) );
  INV_X1 U15471 ( .A(n12376), .ZN(n12378) );
  NOR2_X1 U15472 ( .A1(n12378), .A2(n12377), .ZN(n12380) );
  INV_X1 U15473 ( .A(n12383), .ZN(n12379) );
  OAI22_X1 U15474 ( .A1(n12381), .A2(n12380), .B1(n12385), .B2(n12379), .ZN(
        n12387) );
  NAND3_X1 U15475 ( .A1(n12385), .A2(n12384), .A3(n12383), .ZN(n12386) );
  NAND2_X1 U15476 ( .A1(n12387), .A2(n12386), .ZN(n12388) );
  NAND2_X1 U15477 ( .A1(n12390), .A2(n12389), .ZN(n12391) );
  NAND2_X1 U15478 ( .A1(n13367), .A2(n13262), .ZN(n12393) );
  NAND3_X1 U15479 ( .A1(n14599), .A2(n14815), .A3(n20141), .ZN(n12409) );
  NOR4_X1 U15480 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(
        P1_ADDRESS_REG_15__SCAN_IN), .A3(P1_ADDRESS_REG_14__SCAN_IN), .A4(
        P1_ADDRESS_REG_13__SCAN_IN), .ZN(n12398) );
  NOR4_X1 U15481 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(
        P1_ADDRESS_REG_19__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_18__SCAN_IN), .ZN(n12397) );
  NOR4_X1 U15482 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(
        P1_ADDRESS_REG_7__SCAN_IN), .A3(P1_ADDRESS_REG_6__SCAN_IN), .A4(
        P1_ADDRESS_REG_5__SCAN_IN), .ZN(n12396) );
  NOR4_X1 U15483 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_11__SCAN_IN), .A4(
        P1_ADDRESS_REG_10__SCAN_IN), .ZN(n12395) );
  AND4_X1 U15484 ( .A1(n12398), .A2(n12397), .A3(n12396), .A4(n12395), .ZN(
        n12403) );
  NOR4_X1 U15485 ( .A1(P1_ADDRESS_REG_4__SCAN_IN), .A2(
        P1_ADDRESS_REG_3__SCAN_IN), .A3(P1_ADDRESS_REG_0__SCAN_IN), .A4(
        P1_ADDRESS_REG_2__SCAN_IN), .ZN(n12401) );
  NOR4_X1 U15486 ( .A1(P1_ADDRESS_REG_24__SCAN_IN), .A2(
        P1_ADDRESS_REG_23__SCAN_IN), .A3(P1_ADDRESS_REG_22__SCAN_IN), .A4(
        P1_ADDRESS_REG_21__SCAN_IN), .ZN(n12400) );
  NOR4_X1 U15487 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(
        P1_ADDRESS_REG_27__SCAN_IN), .A3(P1_ADDRESS_REG_26__SCAN_IN), .A4(
        P1_ADDRESS_REG_25__SCAN_IN), .ZN(n12399) );
  INV_X1 U15488 ( .A(P1_ADDRESS_REG_1__SCAN_IN), .ZN(n20681) );
  AND4_X1 U15489 ( .A1(n12401), .A2(n12400), .A3(n12399), .A4(n20681), .ZN(
        n12402) );
  NAND2_X1 U15490 ( .A1(n12403), .A2(n12402), .ZN(n12404) );
  INV_X1 U15491 ( .A(n20099), .ZN(n20101) );
  AOI22_X1 U15492 ( .A1(n15948), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n15946), .ZN(n12405) );
  INV_X1 U15493 ( .A(n12405), .ZN(n12407) );
  NAND2_X1 U15494 ( .A1(n13418), .A2(n20099), .ZN(n15952) );
  INV_X1 U15495 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16425) );
  NOR2_X1 U15496 ( .A1(n12407), .A2(n12406), .ZN(n12408) );
  NAND2_X1 U15497 ( .A1(n12409), .A2(n12408), .ZN(P1_U2873) );
  INV_X1 U15498 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16540) );
  INV_X1 U15499 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16550) );
  NAND2_X1 U15500 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16764) );
  NOR3_X1 U15501 ( .A1(n16764), .A2(n16763), .A3(n17685), .ZN(n16721) );
  NAND2_X1 U15502 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17662) );
  NAND2_X1 U15503 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17619) );
  NAND2_X1 U15504 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17586) );
  INV_X1 U15505 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17564) );
  NOR2_X1 U15506 ( .A1(n17564), .A2(n17549), .ZN(n17545) );
  INV_X1 U15507 ( .A(n17545), .ZN(n12411) );
  NAND2_X1 U15508 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17534), .ZN(
        n17504) );
  NAND2_X1 U15509 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17505) );
  NAND2_X1 U15510 ( .A1(n17494), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17467) );
  NAND2_X1 U15511 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17468) );
  XNOR2_X1 U15512 ( .A(n16540), .B(n12421), .ZN(n16539) );
  AOI21_X1 U15513 ( .B1(n16550), .B2(n12412), .A(n12421), .ZN(n16549) );
  INV_X1 U15514 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17487) );
  INV_X1 U15515 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17507) );
  INV_X1 U15516 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17536) );
  INV_X1 U15517 ( .A(n12420), .ZN(n12419) );
  NOR2_X1 U15518 ( .A1(n12411), .A2(n12419), .ZN(n12417) );
  INV_X1 U15519 ( .A(n12417), .ZN(n17503) );
  NAND2_X1 U15520 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n12416), .ZN(
        n12415) );
  NAND2_X1 U15521 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n17464), .ZN(
        n12414) );
  NOR2_X1 U15522 ( .A1(n17487), .A2(n12414), .ZN(n12413) );
  OAI21_X1 U15523 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n12413), .A(
        n12412), .ZN(n17471) );
  INV_X1 U15524 ( .A(n17471), .ZN(n16564) );
  AOI21_X1 U15525 ( .B1(n17487), .B2(n12414), .A(n12413), .ZN(n17483) );
  OAI21_X1 U15526 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17464), .A(
        n12414), .ZN(n17497) );
  INV_X1 U15527 ( .A(n17497), .ZN(n16584) );
  AOI21_X1 U15528 ( .B1(n17507), .B2(n12415), .A(n17464), .ZN(n17509) );
  OAI21_X1 U15529 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n12416), .A(
        n12415), .ZN(n17519) );
  INV_X1 U15530 ( .A(n17519), .ZN(n16609) );
  AOI21_X1 U15531 ( .B1(n17536), .B2(n17503), .A(n12416), .ZN(n17532) );
  NAND2_X1 U15532 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12420), .ZN(
        n12418) );
  AOI21_X1 U15533 ( .B1(n17549), .B2(n12418), .A(n12417), .ZN(n17552) );
  AOI22_X1 U15534 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n12420), .B1(
        n12419), .B2(n17564), .ZN(n17567) );
  NAND2_X1 U15535 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n9677), .ZN(
        n17546) );
  AOI21_X1 U15536 ( .B1(n9903), .B2(n17546), .A(n12420), .ZN(n17578) );
  NAND2_X1 U15537 ( .A1(n12421), .A2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12422) );
  INV_X1 U15538 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13004) );
  INV_X1 U15539 ( .A(n17619), .ZN(n12423) );
  NOR2_X1 U15540 ( .A1(n17816), .A2(n17618), .ZN(n17617) );
  NAND2_X1 U15541 ( .A1(n12423), .A2(n17617), .ZN(n16690) );
  NOR2_X1 U15542 ( .A1(n9902), .A2(n16690), .ZN(n17584) );
  NAND2_X1 U15543 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17584), .ZN(
        n16666) );
  INV_X1 U15544 ( .A(n16666), .ZN(n16653) );
  NAND2_X1 U15545 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17617), .ZN(
        n16699) );
  NOR2_X1 U15546 ( .A1(n16699), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16693) );
  NOR2_X1 U15547 ( .A1(n17578), .A2(n16647), .ZN(n16646) );
  NOR2_X1 U15548 ( .A1(n16646), .A2(n16845), .ZN(n16636) );
  NOR2_X1 U15549 ( .A1(n17567), .A2(n16636), .ZN(n16635) );
  NOR2_X1 U15550 ( .A1(n16635), .A2(n16845), .ZN(n16630) );
  NOR2_X1 U15551 ( .A1(n17552), .A2(n16630), .ZN(n16629) );
  NOR2_X1 U15552 ( .A1(n16629), .A2(n16845), .ZN(n16616) );
  NOR2_X1 U15553 ( .A1(n17532), .A2(n16616), .ZN(n16615) );
  NOR2_X1 U15554 ( .A1(n16615), .A2(n16845), .ZN(n16608) );
  NOR2_X1 U15555 ( .A1(n16609), .A2(n16608), .ZN(n16607) );
  NOR2_X1 U15556 ( .A1(n16607), .A2(n16845), .ZN(n16597) );
  NOR2_X1 U15557 ( .A1(n17509), .A2(n16597), .ZN(n16596) );
  NOR2_X1 U15558 ( .A1(n16596), .A2(n16845), .ZN(n16583) );
  NOR2_X1 U15559 ( .A1(n16584), .A2(n16583), .ZN(n16582) );
  NOR2_X1 U15560 ( .A1(n16582), .A2(n16845), .ZN(n16571) );
  NOR2_X1 U15561 ( .A1(n17483), .A2(n16571), .ZN(n16572) );
  NOR2_X1 U15562 ( .A1(n16572), .A2(n16845), .ZN(n16563) );
  NOR2_X1 U15563 ( .A1(n16564), .A2(n16563), .ZN(n16562) );
  NOR2_X1 U15564 ( .A1(n16562), .A2(n16845), .ZN(n16547) );
  NOR2_X1 U15565 ( .A1(n16548), .A2(n16845), .ZN(n16538) );
  INV_X1 U15566 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n14386) );
  INV_X1 U15567 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18813) );
  NAND4_X1 U15568 ( .A1(n18661), .A2(n14386), .A3(n18813), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n18667) );
  NOR2_X1 U15569 ( .A1(n16845), .A2(n18667), .ZN(n16877) );
  INV_X1 U15570 ( .A(n16877), .ZN(n16689) );
  NAND2_X1 U15571 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .ZN(n12444) );
  INV_X2 U15572 ( .A(n18823), .ZN(n18822) );
  NAND2_X2 U15573 ( .A1(n18822), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18752) );
  OAI211_X1 U15574 ( .C1(P3_STATE_REG_1__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18688), .B(n18752), .ZN(n18812) );
  NAND2_X1 U15575 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18815) );
  INV_X1 U15576 ( .A(n18815), .ZN(n18681) );
  AOI211_X1 U15577 ( .C1(n18812), .C2(n18164), .A(n18681), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n12447) );
  INV_X1 U15578 ( .A(n12447), .ZN(n18653) );
  NAND2_X1 U15579 ( .A1(n18160), .A2(n17292), .ZN(n12435) );
  NOR2_X1 U15580 ( .A1(n18187), .A2(n18182), .ZN(n12427) );
  INV_X1 U15581 ( .A(n12427), .ZN(n12424) );
  NAND3_X1 U15582 ( .A1(n18169), .A2(n18610), .A3(n12992), .ZN(n12431) );
  INV_X1 U15583 ( .A(n12425), .ZN(n18178) );
  NOR2_X1 U15584 ( .A1(n18193), .A2(n12427), .ZN(n12428) );
  OAI22_X1 U15585 ( .A1(n18178), .A2(n12428), .B1(n12427), .B2(n12426), .ZN(
        n12429) );
  AOI21_X1 U15586 ( .B1(n18173), .B2(n12435), .A(n12429), .ZN(n12430) );
  OAI21_X1 U15587 ( .B1(n18814), .B2(n12431), .A(n12430), .ZN(n15694) );
  NOR2_X1 U15588 ( .A1(n9732), .A2(n18160), .ZN(n12988) );
  OAI21_X1 U15589 ( .B1(n18193), .B2(n18630), .A(n12988), .ZN(n12432) );
  INV_X1 U15590 ( .A(n12432), .ZN(n15693) );
  AOI211_X1 U15591 ( .C1(n12433), .C2(n12436), .A(n15694), .B(n15693), .ZN(
        n12984) );
  NAND2_X1 U15592 ( .A1(n12438), .A2(n12984), .ZN(n12982) );
  NOR2_X1 U15593 ( .A1(n12435), .A2(n12434), .ZN(n12439) );
  NAND2_X1 U15594 ( .A1(n12438), .A2(n12990), .ZN(n15696) );
  NAND2_X1 U15595 ( .A1(n15697), .A2(n15696), .ZN(n16520) );
  INV_X2 U15596 ( .A(n12983), .ZN(n18619) );
  NAND2_X1 U15597 ( .A1(n12443), .A2(n12442), .ZN(n12440) );
  OAI211_X1 U15598 ( .C1(n12443), .C2(n12442), .A(n12441), .B(n12440), .ZN(
        n12998) );
  NAND2_X1 U15599 ( .A1(n18773), .A2(n18763), .ZN(n18825) );
  OR3_X2 U15600 ( .A1(n18825), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18141) );
  INV_X1 U15601 ( .A(n18806), .ZN(n18827) );
  NAND2_X1 U15602 ( .A1(n18661), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18533) );
  OR2_X1 U15603 ( .A1(n18664), .A2(n18533), .ZN(n18658) );
  NOR2_X1 U15604 ( .A1(n16843), .A2(n16862), .ZN(n16627) );
  INV_X1 U15605 ( .A(n16627), .ZN(n16889) );
  INV_X1 U15606 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18743) );
  INV_X1 U15607 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18741) );
  INV_X1 U15608 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18739) );
  INV_X1 U15609 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18734) );
  INV_X1 U15610 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18712) );
  INV_X1 U15611 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18705) );
  INV_X1 U15612 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18700) );
  INV_X1 U15613 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18696) );
  NAND3_X1 U15614 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16834) );
  NOR2_X1 U15615 ( .A1(n18696), .A2(n16834), .ZN(n16823) );
  NAND2_X1 U15616 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16823), .ZN(n16822) );
  NOR2_X1 U15617 ( .A1(n18700), .A2(n16822), .ZN(n16794) );
  NAND2_X1 U15618 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n16794), .ZN(n16787) );
  NOR2_X1 U15619 ( .A1(n18705), .A2(n16787), .ZN(n16745) );
  NAND4_X1 U15620 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16745), .A3(
        P3_REIP_REG_10__SCAN_IN), .A4(P3_REIP_REG_9__SCAN_IN), .ZN(n16744) );
  NOR2_X1 U15621 ( .A1(n18712), .A2(n16744), .ZN(n16709) );
  NAND3_X1 U15622 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n16709), .ZN(n16626) );
  INV_X1 U15623 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18729) );
  NAND3_X1 U15624 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_16__SCAN_IN), 
        .A3(P3_REIP_REG_15__SCAN_IN), .ZN(n16660) );
  NAND2_X1 U15625 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16661) );
  NOR3_X1 U15626 ( .A1(n18729), .A2(n16660), .A3(n16661), .ZN(n16628) );
  NAND3_X1 U15627 ( .A1(n16628), .A2(P3_REIP_REG_22__SCAN_IN), .A3(
        P3_REIP_REG_21__SCAN_IN), .ZN(n16614) );
  NOR3_X1 U15628 ( .A1(n18734), .A2(n16626), .A3(n16614), .ZN(n16605) );
  NAND2_X1 U15629 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16605), .ZN(n16579) );
  NOR3_X1 U15630 ( .A1(n18741), .A2(n18739), .A3(n16579), .ZN(n12445) );
  OAI21_X1 U15631 ( .B1(n12445), .B2(n16879), .A(n16891), .ZN(n16560) );
  AOI221_X1 U15632 ( .B1(n12444), .B2(n16889), .C1(n18743), .C2(n16889), .A(
        n16560), .ZN(n16558) );
  NAND2_X1 U15633 ( .A1(n16843), .A2(n12445), .ZN(n16573) );
  NOR2_X1 U15634 ( .A1(n18743), .A2(n16573), .ZN(n16559) );
  NAND3_X1 U15635 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(n16559), .ZN(n12449) );
  NOR2_X1 U15636 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n12449), .ZN(n16542) );
  INV_X1 U15637 ( .A(n16542), .ZN(n12446) );
  INV_X1 U15638 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18749) );
  AOI21_X1 U15639 ( .B1(n16558), .B2(n12446), .A(n18749), .ZN(n12456) );
  AOI211_X1 U15640 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n9732), .A(n12447), .B(
        n12452), .ZN(n12448) );
  INV_X1 U15641 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18751) );
  NOR3_X1 U15642 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18751), .A3(n12449), 
        .ZN(n12450) );
  AOI21_X1 U15643 ( .B1(n16883), .B2(P3_EBX_REG_31__SCAN_IN), .A(n12450), .ZN(
        n12454) );
  NAND2_X1 U15644 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n9732), .ZN(n12451) );
  AOI211_X4 U15645 ( .C1(n18813), .C2(n18815), .A(n12452), .B(n12451), .ZN(
        n16848) );
  NOR3_X1 U15646 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16858) );
  NAND2_X1 U15647 ( .A1(n16858), .A2(n16849), .ZN(n16847) );
  NOR2_X1 U15648 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16847), .ZN(n16833) );
  INV_X1 U15649 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16821) );
  NAND2_X1 U15650 ( .A1(n16833), .A2(n16821), .ZN(n16820) );
  NAND2_X1 U15651 ( .A1(n16806), .A2(n17121), .ZN(n16799) );
  NAND2_X1 U15652 ( .A1(n16772), .A2(n16780), .ZN(n16756) );
  NAND2_X1 U15653 ( .A1(n16755), .A2(n17119), .ZN(n16752) );
  NAND2_X1 U15654 ( .A1(n16734), .A2(n16724), .ZN(n16723) );
  NAND2_X1 U15655 ( .A1(n16715), .A2(n16703), .ZN(n16702) );
  INV_X1 U15656 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16681) );
  NAND2_X1 U15657 ( .A1(n16685), .A2(n16681), .ZN(n16680) );
  NAND2_X1 U15658 ( .A1(n16664), .A2(n17011), .ZN(n16656) );
  INV_X1 U15659 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n20795) );
  NAND2_X1 U15660 ( .A1(n16644), .A2(n20795), .ZN(n16637) );
  INV_X1 U15661 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16895) );
  NAND2_X1 U15662 ( .A1(n16624), .A2(n16895), .ZN(n16621) );
  NOR2_X1 U15663 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16621), .ZN(n16594) );
  INV_X1 U15664 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16600) );
  NAND2_X1 U15665 ( .A1(n16594), .A2(n16600), .ZN(n16581) );
  NOR2_X1 U15666 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16581), .ZN(n16580) );
  NAND2_X1 U15667 ( .A1(n16580), .A2(n16897), .ZN(n16576) );
  NOR2_X1 U15668 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16576), .ZN(n16561) );
  INV_X1 U15669 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16934) );
  NAND2_X1 U15670 ( .A1(n16561), .A2(n16934), .ZN(n16537) );
  NOR2_X1 U15671 ( .A1(n16887), .A2(n16537), .ZN(n16544) );
  INV_X1 U15672 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16904) );
  NAND2_X1 U15673 ( .A1(n16544), .A2(n16904), .ZN(n12453) );
  NAND3_X1 U15674 ( .A1(n12454), .A2(n12453), .A3(n10052), .ZN(n12455) );
  OAI22_X1 U15675 ( .A1(n15227), .A2(n15417), .B1(n12460), .B2(n12459), .ZN(
        n12463) );
  XOR2_X1 U15676 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n12461), .Z(
        n12462) );
  XNOR2_X1 U15677 ( .A(n12463), .B(n12462), .ZN(n12484) );
  AND2_X1 U15678 ( .A1(n13069), .A2(n12464), .ZN(n12465) );
  OR2_X1 U15679 ( .A1(n12466), .A2(n12465), .ZN(n16181) );
  NOR2_X1 U15680 ( .A1(n19155), .A2(n12467), .ZN(n12478) );
  NOR2_X1 U15681 ( .A1(n12468), .A2(n15396), .ZN(n12469) );
  AOI211_X1 U15682 ( .C1(n15338), .C2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n12478), .B(n12469), .ZN(n12470) );
  OAI21_X1 U15683 ( .B1(n13862), .B2(n16181), .A(n12470), .ZN(n12471) );
  AOI21_X1 U15684 ( .B1(n12484), .B2(n11114), .A(n12471), .ZN(n12473) );
  XNOR2_X1 U15685 ( .A(n15228), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12485) );
  OR2_X1 U15686 ( .A1(n12485), .A2(n19148), .ZN(n12472) );
  NAND2_X1 U15687 ( .A1(n12473), .A2(n12472), .ZN(P2_U2986) );
  AND2_X1 U15688 ( .A1(n13074), .A2(n12474), .ZN(n12475) );
  NOR2_X1 U15689 ( .A1(n12476), .A2(n12475), .ZN(n16179) );
  NOR3_X1 U15690 ( .A1(n15417), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n12480), .ZN(n12477) );
  AOI211_X1 U15691 ( .C1(n16179), .C2(n16296), .A(n12478), .B(n12477), .ZN(
        n12482) );
  INV_X1 U15692 ( .A(n12479), .ZN(n15418) );
  INV_X1 U15693 ( .A(n12480), .ZN(n15402) );
  NAND2_X1 U15694 ( .A1(n15417), .A2(n15402), .ZN(n15419) );
  NAND2_X1 U15695 ( .A1(n15418), .A2(n15419), .ZN(n15408) );
  NAND2_X1 U15696 ( .A1(n15408), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12481) );
  OAI211_X1 U15697 ( .C1(n16181), .C2(n19179), .A(n12482), .B(n12481), .ZN(
        n12483) );
  AOI21_X1 U15698 ( .B1(n12484), .B2(n19188), .A(n12483), .ZN(n12487) );
  NAND2_X1 U15699 ( .A1(n12487), .A2(n12486), .ZN(P2_U3018) );
  NOR2_X1 U15700 ( .A1(n12488), .A2(n15396), .ZN(n12489) );
  AOI211_X1 U15701 ( .C1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(n15338), .A(
        n12490), .B(n12489), .ZN(n12491) );
  OAI21_X1 U15702 ( .B1(n14392), .B2(n13862), .A(n12491), .ZN(n12492) );
  AOI21_X1 U15703 ( .B1(n12493), .B2(n11114), .A(n12492), .ZN(n12496) );
  NAND2_X1 U15704 ( .A1(n12496), .A2(n12495), .ZN(P2_U2983) );
  NAND2_X1 U15705 ( .A1(n12498), .A2(n12510), .ZN(n12502) );
  AND2_X1 U15706 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19490) );
  NAND2_X1 U15707 ( .A1(n19490), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n14038) );
  NAND2_X1 U15708 ( .A1(n14038), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12499) );
  NAND3_X1 U15709 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A3(n19775), .ZN(n19378) );
  INV_X1 U15710 ( .A(n19378), .ZN(n13866) );
  NAND2_X1 U15711 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13866), .ZN(
        n19429) );
  NAND2_X1 U15712 ( .A1(n12499), .A2(n19429), .ZN(n12500) );
  AND2_X1 U15713 ( .A1(n12500), .A2(n19764), .ZN(n19525) );
  AOI21_X1 U15714 ( .B1(n12516), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19525), .ZN(n12501) );
  NAND2_X1 U15715 ( .A1(n12527), .A2(n12503), .ZN(n13594) );
  OAI21_X1 U15716 ( .B1(n12503), .B2(n12527), .A(n13594), .ZN(n12504) );
  INV_X1 U15717 ( .A(n12504), .ZN(n13510) );
  AOI22_X1 U15718 ( .A1(n12516), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19764), .B2(n19802), .ZN(n12505) );
  XNOR2_X1 U15719 ( .A(n13299), .B(n12511), .ZN(n13527) );
  NAND2_X1 U15720 ( .A1(n12516), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12508) );
  NAND2_X1 U15721 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19793), .ZN(
        n19223) );
  NAND2_X1 U15722 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19802), .ZN(
        n19459) );
  NAND2_X1 U15723 ( .A1(n19223), .A2(n19459), .ZN(n19310) );
  NAND2_X1 U15724 ( .A1(n19764), .A2(n19310), .ZN(n19462) );
  NAND2_X1 U15725 ( .A1(n12508), .A2(n19462), .ZN(n12509) );
  NAND2_X1 U15726 ( .A1(n13527), .A2(n13526), .ZN(n13529) );
  INV_X1 U15727 ( .A(n13299), .ZN(n13941) );
  NAND2_X1 U15728 ( .A1(n13941), .A2(n12511), .ZN(n12512) );
  INV_X1 U15729 ( .A(n19764), .ZN(n19771) );
  INV_X1 U15730 ( .A(n19490), .ZN(n12513) );
  NAND2_X1 U15731 ( .A1(n12513), .A2(n19784), .ZN(n12514) );
  NAND2_X1 U15732 ( .A1(n14038), .A2(n12514), .ZN(n19311) );
  NOR2_X1 U15733 ( .A1(n19771), .A2(n19311), .ZN(n12515) );
  AOI21_X1 U15734 ( .B1(n12516), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12515), .ZN(n12517) );
  OAI21_X2 U15735 ( .B1(n12519), .B2(n12518), .A(n12517), .ZN(n12523) );
  NAND2_X1 U15736 ( .A1(n13517), .A2(n13516), .ZN(n13521) );
  INV_X1 U15737 ( .A(n12521), .ZN(n12522) );
  NAND2_X1 U15738 ( .A1(n12523), .A2(n12522), .ZN(n12524) );
  NAND2_X1 U15739 ( .A1(n13510), .A2(n13511), .ZN(n12526) );
  NAND2_X1 U15740 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n10185), .ZN(
        n12525) );
  NAND2_X1 U15741 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12529) );
  NAND2_X1 U15742 ( .A1(n13655), .A2(n12531), .ZN(n12532) );
  AND2_X1 U15743 ( .A1(n13813), .A2(n13815), .ZN(n12533) );
  NAND2_X1 U15744 ( .A1(n13729), .A2(n12533), .ZN(n13814) );
  OAI22_X1 U15745 ( .A1(n12539), .A2(n12538), .B1(n12537), .B2(n14056), .ZN(
        n12558) );
  INV_X1 U15746 ( .A(n12540), .ZN(n12544) );
  INV_X1 U15747 ( .A(n12541), .ZN(n12542) );
  OAI22_X1 U15748 ( .A1(n12544), .A2(n12543), .B1(n12542), .B2(n13871), .ZN(
        n12557) );
  INV_X1 U15749 ( .A(n12545), .ZN(n12550) );
  INV_X1 U15750 ( .A(n12546), .ZN(n12548) );
  OAI22_X1 U15751 ( .A1(n12550), .A2(n12549), .B1(n12548), .B2(n12547), .ZN(
        n12556) );
  INV_X1 U15752 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12554) );
  INV_X1 U15753 ( .A(n12552), .ZN(n12553) );
  OAI22_X1 U15754 ( .A1(n9612), .A2(n12554), .B1(n12553), .B2(n13501), .ZN(
        n12555) );
  NOR4_X1 U15755 ( .A1(n12558), .A2(n12557), .A3(n12556), .A4(n12555), .ZN(
        n12567) );
  OAI22_X1 U15756 ( .A1(n12650), .A2(n12560), .B1(n12666), .B2(n12559), .ZN(
        n12563) );
  INV_X1 U15757 ( .A(n12660), .ZN(n12640) );
  NOR2_X1 U15758 ( .A1(n12640), .A2(n12561), .ZN(n12562) );
  AOI211_X1 U15759 ( .C1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .C2(n10320), .A(
        n12563), .B(n12562), .ZN(n12566) );
  AOI22_X1 U15760 ( .A1(n12670), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12565) );
  AOI22_X1 U15761 ( .A1(n12631), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12665), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12564) );
  NAND4_X1 U15762 ( .A1(n12567), .A2(n12566), .A3(n12565), .A4(n12564), .ZN(
        n14253) );
  AOI22_X1 U15763 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10933), .B1(
        n10934), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12571) );
  AOI22_X1 U15764 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12540), .B1(
        n12541), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12570) );
  AOI22_X1 U15765 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12551), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12569) );
  AOI22_X1 U15766 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n12546), .B1(
        n12545), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12568) );
  NAND4_X1 U15767 ( .A1(n12571), .A2(n12570), .A3(n12569), .A4(n12568), .ZN(
        n12580) );
  AOI22_X1 U15768 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12670), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12578) );
  AOI22_X1 U15769 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12665), .B1(
        n12631), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12577) );
  INV_X1 U15770 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12572) );
  OAI22_X1 U15771 ( .A1(n12650), .A2(n12573), .B1(n12572), .B2(n12666), .ZN(
        n12574) );
  AOI21_X1 U15772 ( .B1(n10320), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A(
        n12574), .ZN(n12576) );
  NAND2_X1 U15773 ( .A1(n12660), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12575) );
  NAND4_X1 U15774 ( .A1(n12578), .A2(n12577), .A3(n12576), .A4(n12575), .ZN(
        n12579) );
  OR2_X1 U15775 ( .A1(n12580), .A2(n12579), .ZN(n14380) );
  INV_X1 U15776 ( .A(n14380), .ZN(n12607) );
  AOI22_X1 U15777 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n10933), .B1(
        n10934), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12584) );
  AOI22_X1 U15778 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n12540), .B1(
        n12541), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12583) );
  AOI22_X1 U15779 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n12551), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12582) );
  AOI22_X1 U15780 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n12546), .B1(
        n12545), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12581) );
  NAND4_X1 U15781 ( .A1(n12584), .A2(n12583), .A3(n12582), .A4(n12581), .ZN(
        n12593) );
  AOI22_X1 U15782 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n12670), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12591) );
  AOI22_X1 U15783 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n12665), .B1(
        n12631), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12590) );
  INV_X1 U15784 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12585) );
  OAI22_X1 U15785 ( .A1(n12650), .A2(n12586), .B1(n12585), .B2(n12666), .ZN(
        n12587) );
  AOI21_X1 U15786 ( .B1(n10320), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A(
        n12587), .ZN(n12589) );
  NAND2_X1 U15787 ( .A1(n12660), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12588) );
  NAND4_X1 U15788 ( .A1(n12591), .A2(n12590), .A3(n12589), .A4(n12588), .ZN(
        n12592) );
  NOR2_X1 U15789 ( .A1(n12593), .A2(n12592), .ZN(n14214) );
  AOI22_X1 U15790 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n10933), .B1(
        n10934), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12597) );
  AOI22_X1 U15791 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n12540), .B1(
        n12541), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12596) );
  AOI22_X1 U15792 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n12551), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12595) );
  AOI22_X1 U15793 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n12546), .B1(
        n12545), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12594) );
  NAND4_X1 U15794 ( .A1(n12597), .A2(n12596), .A3(n12595), .A4(n12594), .ZN(
        n12606) );
  AOI22_X1 U15795 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n12670), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12604) );
  AOI22_X1 U15796 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n12665), .B1(
        n12631), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12603) );
  INV_X1 U15797 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12598) );
  OAI22_X1 U15798 ( .A1(n12650), .A2(n12599), .B1(n12598), .B2(n12666), .ZN(
        n12600) );
  AOI21_X1 U15799 ( .B1(n10320), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A(
        n12600), .ZN(n12602) );
  NAND2_X1 U15800 ( .A1(n12660), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n12601) );
  NAND4_X1 U15801 ( .A1(n12604), .A2(n12603), .A3(n12602), .A4(n12601), .ZN(
        n12605) );
  NOR2_X1 U15802 ( .A1(n12606), .A2(n12605), .ZN(n14241) );
  OR2_X1 U15803 ( .A1(n14214), .A2(n14241), .ZN(n14215) );
  NOR2_X1 U15804 ( .A1(n12607), .A2(n14215), .ZN(n14249) );
  AND2_X1 U15805 ( .A1(n14253), .A2(n14249), .ZN(n12621) );
  AOI22_X1 U15806 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n10933), .B1(
        n10934), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12611) );
  AOI22_X1 U15807 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n12540), .B1(
        n12541), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12610) );
  AOI22_X1 U15808 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n12551), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12609) );
  AOI22_X1 U15809 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n12546), .B1(
        n12545), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12608) );
  NAND4_X1 U15810 ( .A1(n12611), .A2(n12610), .A3(n12609), .A4(n12608), .ZN(
        n12620) );
  AOI22_X1 U15811 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n12670), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12618) );
  AOI22_X1 U15812 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n12665), .B1(
        n12631), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12617) );
  OAI22_X1 U15813 ( .A1(n10339), .A2(n12613), .B1(n12612), .B2(n12666), .ZN(
        n12614) );
  AOI21_X1 U15814 ( .B1(n10320), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A(
        n12614), .ZN(n12616) );
  NAND2_X1 U15815 ( .A1(n12660), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12615) );
  NAND4_X1 U15816 ( .A1(n12618), .A2(n12617), .A3(n12616), .A4(n12615), .ZN(
        n12619) );
  OR2_X1 U15817 ( .A1(n12620), .A2(n12619), .ZN(n14248) );
  AND2_X1 U15818 ( .A1(n12621), .A2(n14248), .ZN(n14251) );
  AOI22_X1 U15819 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10933), .B1(
        n10934), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12625) );
  AOI22_X1 U15820 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n12540), .B1(
        n12541), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12624) );
  AOI22_X1 U15821 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n12551), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12623) );
  AOI22_X1 U15822 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n12545), .B1(
        n12546), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12622) );
  NAND4_X1 U15823 ( .A1(n12625), .A2(n12624), .A3(n12623), .A4(n12622), .ZN(
        n12644) );
  INV_X1 U15824 ( .A(n12670), .ZN(n12629) );
  INV_X1 U15825 ( .A(n12626), .ZN(n12628) );
  OAI22_X1 U15826 ( .A1(n12630), .A2(n12629), .B1(n12628), .B2(n12627), .ZN(
        n12643) );
  INV_X1 U15827 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12635) );
  INV_X1 U15828 ( .A(n12631), .ZN(n12634) );
  INV_X1 U15829 ( .A(n12665), .ZN(n12633) );
  INV_X1 U15830 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12632) );
  OAI22_X1 U15831 ( .A1(n12635), .A2(n12634), .B1(n12633), .B2(n12632), .ZN(
        n12642) );
  OAI22_X1 U15832 ( .A1(n10339), .A2(n12636), .B1(n14192), .B2(n12666), .ZN(
        n12637) );
  AOI21_X1 U15833 ( .B1(n10320), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n12637), .ZN(n12638) );
  OAI21_X1 U15834 ( .B1(n12640), .B2(n12639), .A(n12638), .ZN(n12641) );
  OR4_X1 U15835 ( .A1(n12644), .A2(n12643), .A3(n12642), .A4(n12641), .ZN(
        n14338) );
  AND2_X1 U15836 ( .A1(n14251), .A2(n14338), .ZN(n12658) );
  AOI22_X1 U15837 ( .A1(n10933), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n10934), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12648) );
  AOI22_X1 U15838 ( .A1(n12540), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12541), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12647) );
  AOI22_X1 U15839 ( .A1(n12551), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12646) );
  AOI22_X1 U15840 ( .A1(n12545), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12546), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12645) );
  NAND4_X1 U15841 ( .A1(n12648), .A2(n12647), .A3(n12646), .A4(n12645), .ZN(
        n12657) );
  AOI22_X1 U15842 ( .A1(n12670), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12655) );
  AOI22_X1 U15843 ( .A1(n12631), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12665), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12654) );
  INV_X1 U15844 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14198) );
  OAI22_X1 U15845 ( .A1(n12650), .A2(n12649), .B1(n10340), .B2(n14198), .ZN(
        n12651) );
  AOI21_X1 U15846 ( .B1(n10320), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A(
        n12651), .ZN(n12653) );
  NAND2_X1 U15847 ( .A1(n12660), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12652) );
  NAND4_X1 U15848 ( .A1(n12655), .A2(n12654), .A3(n12653), .A4(n12652), .ZN(
        n12656) );
  OR2_X1 U15849 ( .A1(n12657), .A2(n12656), .ZN(n14086) );
  AND2_X1 U15850 ( .A1(n12658), .A2(n14086), .ZN(n12659) );
  AOI22_X1 U15851 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n12541), .B1(
        n10934), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12664) );
  AOI22_X1 U15852 ( .A1(n10933), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12552), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12663) );
  AOI22_X1 U15853 ( .A1(n12540), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n12551), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12662) );
  AOI22_X1 U15854 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n12660), .B1(
        n12546), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12661) );
  NAND4_X1 U15855 ( .A1(n12664), .A2(n12663), .A3(n12662), .A4(n12661), .ZN(
        n12676) );
  AOI22_X1 U15856 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n10320), .B1(
        n12626), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12674) );
  AOI22_X1 U15857 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n12665), .B1(
        n12631), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12673) );
  INV_X1 U15858 ( .A(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12667) );
  OAI22_X1 U15859 ( .A1(n10339), .A2(n12668), .B1(n12667), .B2(n12666), .ZN(
        n12669) );
  AOI21_X1 U15860 ( .B1(n12670), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A(
        n12669), .ZN(n12672) );
  NAND2_X1 U15861 ( .A1(n12545), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n12671) );
  NAND4_X1 U15862 ( .A1(n12674), .A2(n12673), .A3(n12672), .A4(n12671), .ZN(
        n12675) );
  NOR2_X1 U15863 ( .A1(n12676), .A2(n12675), .ZN(n12696) );
  INV_X1 U15864 ( .A(n12696), .ZN(n12695) );
  AOI22_X1 U15865 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12823), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12685) );
  AOI22_X1 U15866 ( .A1(n12832), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12831), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12684) );
  AOI22_X1 U15867 ( .A1(n9598), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12683) );
  INV_X1 U15868 ( .A(n12678), .ZN(n12822) );
  INV_X1 U15869 ( .A(n12822), .ZN(n12824) );
  NAND2_X1 U15870 ( .A1(n12824), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n12681) );
  NAND2_X1 U15871 ( .A1(n12686), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12680) );
  OAI21_X1 U15872 ( .B1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(n12679), .ZN(n12825) );
  AND3_X1 U15873 ( .A1(n12681), .A2(n12680), .A3(n12825), .ZN(n12682) );
  NAND4_X1 U15874 ( .A1(n12685), .A2(n12684), .A3(n12683), .A4(n12682), .ZN(
        n12694) );
  AOI22_X1 U15875 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12692) );
  AOI22_X1 U15876 ( .A1(n12816), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12677), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12691) );
  NAND2_X1 U15877 ( .A1(n12824), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n12688) );
  NAND2_X1 U15878 ( .A1(n12686), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12687) );
  INV_X1 U15879 ( .A(n12825), .ZN(n12803) );
  AND3_X1 U15880 ( .A1(n12688), .A2(n12687), .A3(n12803), .ZN(n12690) );
  AOI22_X1 U15881 ( .A1(n12832), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10300), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12689) );
  NAND4_X1 U15882 ( .A1(n12692), .A2(n12691), .A3(n12690), .A4(n12689), .ZN(
        n12693) );
  NAND2_X1 U15883 ( .A1(n12694), .A2(n12693), .ZN(n12698) );
  INV_X1 U15884 ( .A(n12698), .ZN(n12716) );
  NAND2_X1 U15885 ( .A1(n12695), .A2(n12716), .ZN(n12714) );
  OAI21_X1 U15886 ( .B1(n12780), .B2(n12698), .A(n12696), .ZN(n12697) );
  OAI21_X1 U15887 ( .B1(n12714), .B2(n12780), .A(n12697), .ZN(n12718) );
  NOR2_X1 U15888 ( .A1(n10173), .A2(n12698), .ZN(n15159) );
  NAND2_X1 U15889 ( .A1(n15158), .A2(n10057), .ZN(n15146) );
  AOI22_X1 U15890 ( .A1(n12699), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12705) );
  AOI22_X1 U15891 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12677), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12704) );
  NAND2_X1 U15892 ( .A1(n12824), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n12701) );
  NAND2_X1 U15893 ( .A1(n10293), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n12700) );
  AND3_X1 U15894 ( .A1(n12701), .A2(n12700), .A3(n12825), .ZN(n12703) );
  AOI22_X1 U15895 ( .A1(n12832), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12831), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12702) );
  NAND4_X1 U15896 ( .A1(n12705), .A2(n12704), .A3(n12703), .A4(n12702), .ZN(
        n12713) );
  AOI22_X1 U15897 ( .A1(n12823), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9598), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12711) );
  AOI22_X1 U15898 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12710) );
  NAND2_X1 U15899 ( .A1(n12824), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n12707) );
  NAND2_X1 U15900 ( .A1(n10293), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n12706) );
  AND3_X1 U15901 ( .A1(n12707), .A2(n12706), .A3(n12803), .ZN(n12709) );
  AOI22_X1 U15902 ( .A1(n12832), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12831), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12708) );
  NAND4_X1 U15903 ( .A1(n12711), .A2(n12710), .A3(n12709), .A4(n12708), .ZN(
        n12712) );
  NAND2_X1 U15904 ( .A1(n12713), .A2(n12712), .ZN(n12715) );
  NOR2_X1 U15905 ( .A1(n12714), .A2(n12715), .ZN(n12733) );
  AOI211_X1 U15906 ( .C1(n12715), .C2(n12714), .A(n12753), .B(n12733), .ZN(
        n15147) );
  NAND2_X1 U15907 ( .A1(n15146), .A2(n15147), .ZN(n15145) );
  NOR2_X1 U15908 ( .A1(n10173), .A2(n12715), .ZN(n15148) );
  NAND2_X1 U15909 ( .A1(n15148), .A2(n12716), .ZN(n12717) );
  AOI22_X1 U15910 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12724) );
  AOI22_X1 U15911 ( .A1(n12816), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12677), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12723) );
  NAND2_X1 U15912 ( .A1(n12824), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n12720) );
  NAND2_X1 U15913 ( .A1(n10293), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n12719) );
  AND3_X1 U15914 ( .A1(n12720), .A2(n12719), .A3(n12825), .ZN(n12722) );
  AOI22_X1 U15915 ( .A1(n12832), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12831), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12721) );
  NAND4_X1 U15916 ( .A1(n12724), .A2(n12723), .A3(n12722), .A4(n12721), .ZN(
        n12732) );
  AOI22_X1 U15917 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12677), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12730) );
  AOI22_X1 U15918 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12729) );
  NAND2_X1 U15919 ( .A1(n12824), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(
        n12726) );
  NAND2_X1 U15920 ( .A1(n10293), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n12725) );
  AND3_X1 U15921 ( .A1(n12726), .A2(n12725), .A3(n12803), .ZN(n12728) );
  AOI22_X1 U15922 ( .A1(n12832), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12831), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n12727) );
  NAND4_X1 U15923 ( .A1(n12730), .A2(n12729), .A3(n12728), .A4(n12727), .ZN(
        n12731) );
  AND2_X1 U15924 ( .A1(n12732), .A2(n12731), .ZN(n12734) );
  NAND2_X1 U15925 ( .A1(n12733), .A2(n12734), .ZN(n12754) );
  OAI211_X1 U15926 ( .C1(n12733), .C2(n12734), .A(n12754), .B(n12776), .ZN(
        n12737) );
  INV_X1 U15927 ( .A(n12734), .ZN(n12735) );
  NOR2_X1 U15928 ( .A1(n10173), .A2(n12735), .ZN(n15142) );
  NAND2_X1 U15929 ( .A1(n15143), .A2(n15142), .ZN(n15141) );
  INV_X1 U15930 ( .A(n12736), .ZN(n12738) );
  NAND2_X1 U15931 ( .A1(n15141), .A2(n10058), .ZN(n12758) );
  AOI22_X1 U15932 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12744) );
  AOI22_X1 U15933 ( .A1(n12823), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12677), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12743) );
  NAND2_X1 U15934 ( .A1(n12824), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(
        n12740) );
  NAND2_X1 U15935 ( .A1(n10293), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n12739) );
  AND3_X1 U15936 ( .A1(n12740), .A2(n12739), .A3(n12825), .ZN(n12742) );
  AOI22_X1 U15937 ( .A1(n12832), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12831), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12741) );
  NAND4_X1 U15938 ( .A1(n12744), .A2(n12743), .A3(n12742), .A4(n12741), .ZN(
        n12752) );
  AOI22_X1 U15939 ( .A1(n12823), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9598), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12750) );
  AOI22_X1 U15940 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12749) );
  NAND2_X1 U15941 ( .A1(n12824), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n12746) );
  NAND2_X1 U15942 ( .A1(n10293), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n12745) );
  AND3_X1 U15943 ( .A1(n12746), .A2(n12745), .A3(n12803), .ZN(n12748) );
  AOI22_X1 U15944 ( .A1(n12832), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12831), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12747) );
  NAND4_X1 U15945 ( .A1(n12750), .A2(n12749), .A3(n12748), .A4(n12747), .ZN(
        n12751) );
  NAND2_X1 U15946 ( .A1(n12752), .A2(n12751), .ZN(n12756) );
  AOI21_X1 U15947 ( .B1(n12754), .B2(n12756), .A(n12753), .ZN(n12755) );
  XNOR2_X1 U15948 ( .A(n12758), .B(n10074), .ZN(n15134) );
  INV_X1 U15949 ( .A(n12756), .ZN(n12757) );
  NAND2_X1 U15950 ( .A1(n12780), .A2(n12757), .ZN(n15133) );
  AOI22_X1 U15951 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12765) );
  AOI22_X1 U15952 ( .A1(n12816), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12677), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12764) );
  NAND2_X1 U15953 ( .A1(n12824), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n12761) );
  NAND2_X1 U15954 ( .A1(n10293), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n12760) );
  AND3_X1 U15955 ( .A1(n12761), .A2(n12760), .A3(n12825), .ZN(n12763) );
  AOI22_X1 U15956 ( .A1(n12832), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12831), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12762) );
  NAND4_X1 U15957 ( .A1(n12765), .A2(n12764), .A3(n12763), .A4(n12762), .ZN(
        n12773) );
  AOI22_X1 U15958 ( .A1(n12823), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12677), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12771) );
  AOI22_X1 U15959 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12770) );
  NAND2_X1 U15960 ( .A1(n12824), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n12767) );
  NAND2_X1 U15961 ( .A1(n10293), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12766) );
  AND3_X1 U15962 ( .A1(n12767), .A2(n12766), .A3(n12803), .ZN(n12769) );
  AOI22_X1 U15963 ( .A1(n12832), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12831), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12768) );
  NAND4_X1 U15964 ( .A1(n12771), .A2(n12770), .A3(n12769), .A4(n12768), .ZN(
        n12772) );
  NAND2_X1 U15965 ( .A1(n12773), .A2(n12772), .ZN(n12774) );
  INV_X1 U15966 ( .A(n12774), .ZN(n12779) );
  INV_X1 U15967 ( .A(n12775), .ZN(n12777) );
  OR2_X1 U15968 ( .A1(n12775), .A2(n12774), .ZN(n15118) );
  OAI211_X1 U15969 ( .C1(n12779), .C2(n12777), .A(n15118), .B(n12776), .ZN(
        n12778) );
  NAND2_X1 U15970 ( .A1(n12780), .A2(n12779), .ZN(n15126) );
  AOI22_X1 U15971 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12786) );
  AOI22_X1 U15972 ( .A1(n12816), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12677), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12785) );
  NAND2_X1 U15973 ( .A1(n12824), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n12782) );
  NAND2_X1 U15974 ( .A1(n10293), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n12781) );
  AND3_X1 U15975 ( .A1(n12782), .A2(n12781), .A3(n12825), .ZN(n12784) );
  AOI22_X1 U15976 ( .A1(n12832), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n12831), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12783) );
  NAND4_X1 U15977 ( .A1(n12786), .A2(n12785), .A3(n12784), .A4(n12783), .ZN(
        n12794) );
  AOI22_X1 U15978 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12677), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12792) );
  AOI22_X1 U15979 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12791) );
  NAND2_X1 U15980 ( .A1(n12824), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n12788) );
  NAND2_X1 U15981 ( .A1(n10293), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n12787) );
  AND3_X1 U15982 ( .A1(n12788), .A2(n12787), .A3(n12803), .ZN(n12790) );
  AOI22_X1 U15983 ( .A1(n12832), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12831), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12789) );
  NAND4_X1 U15984 ( .A1(n12792), .A2(n12791), .A3(n12790), .A4(n12789), .ZN(
        n12793) );
  AND2_X1 U15985 ( .A1(n12794), .A2(n12793), .ZN(n15120) );
  NAND2_X1 U15986 ( .A1(n10173), .A2(n15120), .ZN(n12796) );
  NOR2_X1 U15987 ( .A1(n15118), .A2(n12796), .ZN(n12813) );
  AOI22_X1 U15988 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12677), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12802) );
  AOI22_X1 U15989 ( .A1(n12816), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12801) );
  NAND2_X1 U15990 ( .A1(n12824), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n12798) );
  NAND2_X1 U15991 ( .A1(n10293), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n12797) );
  AND3_X1 U15992 ( .A1(n12798), .A2(n12797), .A3(n12825), .ZN(n12800) );
  AOI22_X1 U15993 ( .A1(n12832), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12831), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12799) );
  NAND4_X1 U15994 ( .A1(n12802), .A2(n12801), .A3(n12800), .A4(n12799), .ZN(
        n12811) );
  AOI22_X1 U15995 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12677), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12809) );
  AOI22_X1 U15996 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12808) );
  NAND2_X1 U15997 ( .A1(n12824), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n12805) );
  NAND2_X1 U15998 ( .A1(n12832), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12804) );
  AND3_X1 U15999 ( .A1(n12805), .A2(n12804), .A3(n12803), .ZN(n12807) );
  AOI22_X1 U16000 ( .A1(n12831), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12806) );
  NAND4_X1 U16001 ( .A1(n12809), .A2(n12808), .A3(n12807), .A4(n12806), .ZN(
        n12810) );
  AND2_X1 U16002 ( .A1(n12811), .A2(n12810), .ZN(n12812) );
  NAND2_X1 U16003 ( .A1(n12813), .A2(n12812), .ZN(n12814) );
  OAI21_X1 U16004 ( .B1(n12813), .B2(n12812), .A(n12814), .ZN(n14570) );
  INV_X1 U16005 ( .A(n12814), .ZN(n12815) );
  AOI22_X1 U16006 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12816), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12819) );
  AOI22_X1 U16007 ( .A1(n12832), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10293), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12818) );
  NAND2_X1 U16008 ( .A1(n12819), .A2(n12818), .ZN(n12838) );
  AOI22_X1 U16009 ( .A1(n12677), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12821) );
  AOI21_X1 U16010 ( .B1(n12831), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A(
        n12825), .ZN(n12820) );
  OAI211_X1 U16011 ( .C1(n12822), .C2(n14051), .A(n12821), .B(n12820), .ZN(
        n12837) );
  AOI22_X1 U16012 ( .A1(n9601), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12677), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12828) );
  NAND2_X1 U16013 ( .A1(n10293), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n12827) );
  NAND2_X1 U16014 ( .A1(n12824), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n12826) );
  NAND4_X1 U16015 ( .A1(n12828), .A2(n12827), .A3(n12826), .A4(n12825), .ZN(
        n12836) );
  AOI22_X1 U16016 ( .A1(n12830), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n12829), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12834) );
  AOI22_X1 U16017 ( .A1(n12832), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12831), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12833) );
  NAND2_X1 U16018 ( .A1(n12834), .A2(n12833), .ZN(n12835) );
  OAI22_X1 U16019 ( .A1(n12838), .A2(n12837), .B1(n12836), .B2(n12835), .ZN(
        n12839) );
  XNOR2_X1 U16020 ( .A(n12840), .B(n12839), .ZN(n14568) );
  INV_X1 U16021 ( .A(n16325), .ZN(n12841) );
  NAND2_X1 U16022 ( .A1(n16328), .A2(n12841), .ZN(n13161) );
  NAND2_X1 U16023 ( .A1(n13161), .A2(n12842), .ZN(n12843) );
  AND2_X1 U16024 ( .A1(n12844), .A2(n19825), .ZN(n13157) );
  NAND2_X1 U16025 ( .A1(n19819), .A2(n13157), .ZN(n12845) );
  AND2_X1 U16026 ( .A1(n14046), .A2(n12848), .ZN(n12849) );
  NOR4_X1 U16027 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_6__SCAN_IN), .A4(
        P2_ADDRESS_REG_5__SCAN_IN), .ZN(n12853) );
  NOR4_X1 U16028 ( .A1(P2_ADDRESS_REG_14__SCAN_IN), .A2(
        P2_ADDRESS_REG_13__SCAN_IN), .A3(P2_ADDRESS_REG_8__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n12852) );
  NOR4_X1 U16029 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_16__SCAN_IN), .A3(P2_ADDRESS_REG_19__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n12851) );
  NOR4_X1 U16030 ( .A1(P2_ADDRESS_REG_2__SCAN_IN), .A2(
        P2_ADDRESS_REG_10__SCAN_IN), .A3(P2_ADDRESS_REG_1__SCAN_IN), .A4(
        P2_ADDRESS_REG_0__SCAN_IN), .ZN(n12850) );
  NAND4_X1 U16031 ( .A1(n12853), .A2(n12852), .A3(n12851), .A4(n12850), .ZN(
        n12858) );
  NOR4_X1 U16032 ( .A1(P2_ADDRESS_REG_3__SCAN_IN), .A2(
        P2_ADDRESS_REG_4__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_27__SCAN_IN), .ZN(n12856) );
  NOR4_X1 U16033 ( .A1(P2_ADDRESS_REG_22__SCAN_IN), .A2(
        P2_ADDRESS_REG_21__SCAN_IN), .A3(P2_ADDRESS_REG_18__SCAN_IN), .A4(
        P2_ADDRESS_REG_17__SCAN_IN), .ZN(n12855) );
  NOR4_X1 U16034 ( .A1(P2_ADDRESS_REG_26__SCAN_IN), .A2(
        P2_ADDRESS_REG_25__SCAN_IN), .A3(P2_ADDRESS_REG_24__SCAN_IN), .A4(
        P2_ADDRESS_REG_23__SCAN_IN), .ZN(n12854) );
  INV_X1 U16035 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19719) );
  NAND4_X1 U16036 ( .A1(n12856), .A2(n12855), .A3(n12854), .A4(n19719), .ZN(
        n12857) );
  AOI22_X1 U16037 ( .A1(n13863), .A2(BUF1_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n13861), .ZN(n19049) );
  INV_X1 U16038 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n13442) );
  OAI22_X1 U16039 ( .A1(n15206), .A2(n19049), .B1(n19069), .B2(n13442), .ZN(
        n12859) );
  AOI21_X1 U16040 ( .B1(n16173), .B2(n19099), .A(n12859), .ZN(n12863) );
  NOR2_X1 U16041 ( .A1(n12860), .A2(n13295), .ZN(n12861) );
  AOI22_X1 U16042 ( .A1(n19039), .A2(BUF1_REG_30__SCAN_IN), .B1(n19038), .B2(
        BUF2_REG_30__SCAN_IN), .ZN(n12862) );
  AND2_X1 U16043 ( .A1(n12863), .A2(n12862), .ZN(n12864) );
  OAI21_X1 U16044 ( .B1(n14568), .B2(n19103), .A(n12864), .ZN(P2_U2889) );
  AOI22_X1 U16045 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9605), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12874) );
  AOI22_X1 U16046 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9597), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12873) );
  AOI22_X1 U16047 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12865) );
  OAI21_X1 U16048 ( .B1(n9651), .B2(n17176), .A(n12865), .ZN(n12871) );
  AOI22_X1 U16049 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12869) );
  AOI22_X1 U16050 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9606), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12868) );
  AOI22_X1 U16051 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17161), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12867) );
  AOI22_X1 U16052 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9603), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12866) );
  NAND4_X1 U16053 ( .A1(n12869), .A2(n12868), .A3(n12867), .A4(n12866), .ZN(
        n12870) );
  AOI211_X1 U16054 ( .C1(n12941), .C2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A(
        n12871), .B(n12870), .ZN(n12872) );
  AOI22_X1 U16055 ( .A1(n9603), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12885) );
  AOI22_X1 U16056 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12884) );
  INV_X1 U16057 ( .A(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n20906) );
  AOI22_X1 U16058 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12875) );
  OAI21_X1 U16059 ( .B1(n12876), .B2(n20906), .A(n12875), .ZN(n12882) );
  AOI22_X1 U16060 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12880) );
  AOI22_X1 U16061 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12879) );
  AOI22_X1 U16062 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9606), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12878) );
  AOI22_X1 U16063 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12941), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12877) );
  NAND4_X1 U16064 ( .A1(n12880), .A2(n12879), .A3(n12878), .A4(n12877), .ZN(
        n12881) );
  AOI211_X1 U16065 ( .C1(n9597), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n12882), .B(n12881), .ZN(n12883) );
  NAND3_X1 U16066 ( .A1(n12885), .A2(n12884), .A3(n12883), .ZN(n13010) );
  AOI22_X1 U16067 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12895) );
  AOI22_X1 U16068 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9606), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12894) );
  AOI22_X1 U16069 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9623), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12886) );
  OAI21_X1 U16070 ( .B1(n9651), .B2(n17190), .A(n12886), .ZN(n12892) );
  AOI22_X1 U16071 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12890) );
  AOI22_X1 U16072 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12889) );
  AOI22_X1 U16073 ( .A1(n9603), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12888) );
  AOI22_X1 U16074 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12941), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12887) );
  NAND4_X1 U16075 ( .A1(n12890), .A2(n12889), .A3(n12888), .A4(n12887), .ZN(
        n12891) );
  AOI211_X1 U16076 ( .C1(n17020), .C2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n12892), .B(n12891), .ZN(n12893) );
  NAND3_X1 U16077 ( .A1(n12895), .A2(n12894), .A3(n12893), .ZN(n13013) );
  AOI22_X1 U16078 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12905) );
  AOI22_X1 U16079 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9623), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12904) );
  INV_X1 U16080 ( .A(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12903) );
  AOI22_X1 U16081 ( .A1(n11403), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11349), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12896) );
  OAI21_X1 U16082 ( .B1(n9651), .B2(n17198), .A(n12896), .ZN(n12897) );
  INV_X1 U16083 ( .A(n12897), .ZN(n12902) );
  AOI22_X1 U16084 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9596), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12901) );
  AOI22_X1 U16085 ( .A1(n11327), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9603), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12900) );
  AOI22_X1 U16086 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12899) );
  AOI22_X1 U16087 ( .A1(n12941), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12898) );
  AOI22_X1 U16088 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12909) );
  AOI22_X1 U16089 ( .A1(n9603), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12908) );
  AOI22_X1 U16090 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(n9607), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12907) );
  AOI22_X1 U16091 ( .A1(n12941), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12906) );
  NAND4_X1 U16092 ( .A1(n12909), .A2(n12908), .A3(n12907), .A4(n12906), .ZN(
        n12915) );
  AOI22_X1 U16093 ( .A1(n9622), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12913) );
  AOI22_X1 U16094 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17137), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12912) );
  AOI22_X1 U16095 ( .A1(n17154), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9623), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12911) );
  AOI22_X1 U16096 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12910) );
  NAND4_X1 U16097 ( .A1(n12913), .A2(n12912), .A3(n12911), .A4(n12910), .ZN(
        n12914) );
  NAND2_X1 U16098 ( .A1(n17346), .A2(n13015), .ZN(n12939) );
  AOI22_X1 U16099 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17161), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12919) );
  AOI22_X1 U16100 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12918) );
  AOI22_X1 U16101 ( .A1(n9603), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n9602), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12917) );
  AOI22_X1 U16102 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n12941), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12916) );
  NAND4_X1 U16103 ( .A1(n12919), .A2(n12918), .A3(n12917), .A4(n12916), .ZN(
        n12925) );
  AOI22_X1 U16104 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12923) );
  AOI22_X1 U16105 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17156), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12922) );
  AOI22_X1 U16106 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17124), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12921) );
  AOI22_X1 U16107 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12920) );
  NAND4_X1 U16108 ( .A1(n12923), .A2(n12922), .A3(n12921), .A4(n12920), .ZN(
        n12924) );
  AOI22_X1 U16109 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12929) );
  AOI22_X1 U16110 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17137), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12928) );
  AOI22_X1 U16111 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(n9603), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12927) );
  AOI22_X1 U16112 ( .A1(n12941), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12926) );
  NAND4_X1 U16113 ( .A1(n12929), .A2(n12928), .A3(n12927), .A4(n12926), .ZN(
        n12935) );
  AOI22_X1 U16114 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12933) );
  AOI22_X1 U16115 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12932) );
  AOI22_X1 U16116 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9605), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12931) );
  AOI22_X1 U16117 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17161), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12930) );
  NAND4_X1 U16118 ( .A1(n12933), .A2(n12932), .A3(n12931), .A4(n12930), .ZN(
        n12934) );
  INV_X1 U16119 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18086) );
  XOR2_X1 U16120 ( .A(n12936), .B(n17329), .Z(n17760) );
  XOR2_X1 U16121 ( .A(n12937), .B(n13025), .Z(n12938) );
  NAND2_X1 U16122 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n12938), .ZN(
        n12955) );
  XOR2_X1 U16123 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B(n12938), .Z(
        n17774) );
  INV_X1 U16124 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n15717) );
  XOR2_X1 U16125 ( .A(n12939), .B(n17336), .Z(n17791) );
  AOI22_X1 U16126 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(n9623), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12950) );
  AOI22_X1 U16127 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12949) );
  INV_X1 U16128 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17158) );
  AOI22_X1 U16129 ( .A1(n9603), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12940) );
  OAI21_X1 U16130 ( .B1(n9651), .B2(n17158), .A(n12940), .ZN(n12947) );
  AOI22_X1 U16131 ( .A1(n9622), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12945) );
  AOI22_X1 U16132 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12944) );
  AOI22_X1 U16133 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12941), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12943) );
  AOI22_X1 U16134 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12942) );
  NAND4_X1 U16135 ( .A1(n12945), .A2(n12944), .A3(n12943), .A4(n12942), .ZN(
        n12946) );
  AOI211_X1 U16136 ( .C1(n9607), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n12947), .B(n12946), .ZN(n12948) );
  INV_X1 U16137 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18790) );
  NOR2_X1 U16138 ( .A1(n17821), .A2(n18790), .ZN(n17820) );
  NAND2_X1 U16139 ( .A1(n17820), .A2(n17813), .ZN(n17812) );
  INV_X1 U16140 ( .A(n17346), .ZN(n13019) );
  NAND2_X1 U16141 ( .A1(n13019), .A2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n12951) );
  NAND2_X1 U16142 ( .A1(n17812), .A2(n12951), .ZN(n17805) );
  XNOR2_X1 U16143 ( .A(n17346), .B(n13015), .ZN(n12952) );
  INV_X1 U16144 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13016) );
  NAND2_X1 U16145 ( .A1(n17805), .A2(n17806), .ZN(n17804) );
  OR2_X1 U16146 ( .A1(n13016), .A2(n12952), .ZN(n12953) );
  NAND2_X1 U16147 ( .A1(n17804), .A2(n12953), .ZN(n17790) );
  NAND2_X1 U16148 ( .A1(n17791), .A2(n17790), .ZN(n12954) );
  NOR2_X1 U16149 ( .A1(n17791), .A2(n17790), .ZN(n17789) );
  AOI21_X1 U16150 ( .B1(n15717), .B2(n12954), .A(n17789), .ZN(n17773) );
  NAND2_X1 U16151 ( .A1(n17774), .A2(n17773), .ZN(n17772) );
  XOR2_X1 U16152 ( .A(n12957), .B(n12956), .Z(n12958) );
  XOR2_X1 U16153 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n12958), .Z(
        n17751) );
  NAND2_X1 U16154 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n12958), .ZN(
        n12959) );
  AOI21_X1 U16155 ( .B1(n17322), .B2(n12960), .A(n17730), .ZN(n12962) );
  NAND2_X1 U16156 ( .A1(n17740), .A2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17739) );
  INV_X1 U16157 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18037) );
  INV_X1 U16158 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17693) );
  INV_X1 U16159 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17650) );
  NOR2_X2 U16160 ( .A1(n12964), .A2(n18055), .ZN(n17653) );
  NAND2_X1 U16161 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17692) );
  INV_X1 U16162 ( .A(n17692), .ZN(n18019) );
  NAND2_X1 U16163 ( .A1(n18019), .A2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n18005) );
  INV_X1 U16164 ( .A(n18005), .ZN(n17679) );
  NAND3_X1 U16165 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n17679), .A3(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17633) );
  NOR2_X1 U16166 ( .A1(n18012), .A2(n17633), .ZN(n17965) );
  NAND2_X1 U16167 ( .A1(n17965), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17831) );
  NAND2_X1 U16168 ( .A1(n17653), .A2(n17936), .ZN(n12966) );
  INV_X1 U16169 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17962) );
  INV_X1 U16170 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17947) );
  NAND2_X1 U16171 ( .A1(n17611), .A2(n17947), .ZN(n17610) );
  NAND2_X2 U16172 ( .A1(n17610), .A2(n17656), .ZN(n17573) );
  NAND2_X1 U16173 ( .A1(n12967), .A2(n12966), .ZN(n17615) );
  INV_X1 U16174 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17870) );
  NOR2_X1 U16175 ( .A1(n17962), .A2(n17947), .ZN(n17939) );
  INV_X1 U16176 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n20891) );
  INV_X1 U16177 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17932) );
  NOR2_X1 U16178 ( .A1(n20891), .A2(n17932), .ZN(n17568) );
  NAND3_X1 U16179 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n17568), .ZN(n17553) );
  INV_X1 U16180 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17892) );
  NOR2_X1 U16181 ( .A1(n17553), .A2(n17892), .ZN(n12972) );
  NAND2_X1 U16182 ( .A1(n17939), .A2(n12972), .ZN(n17877) );
  NOR2_X1 U16183 ( .A1(n17870), .A2(n17877), .ZN(n17524) );
  NOR2_X1 U16184 ( .A1(n17730), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17600) );
  NAND2_X1 U16185 ( .A1(n17600), .A2(n17932), .ZN(n12968) );
  NOR2_X1 U16186 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n12968), .ZN(
        n17561) );
  INV_X1 U16187 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17906) );
  NAND2_X1 U16188 ( .A1(n17561), .A2(n17906), .ZN(n17543) );
  NOR3_X1 U16189 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(n17543), .ZN(n12969) );
  INV_X1 U16190 ( .A(n12970), .ZN(n12971) );
  NOR2_X2 U16191 ( .A1(n17518), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n17517) );
  NAND2_X1 U16192 ( .A1(n17939), .A2(n17615), .ZN(n17559) );
  NAND2_X1 U16193 ( .A1(n17573), .A2(n17559), .ZN(n17560) );
  NAND2_X1 U16194 ( .A1(n12972), .A2(n17560), .ZN(n17528) );
  NOR3_X1 U16195 ( .A1(n17517), .A2(n17528), .A3(n17870), .ZN(n12974) );
  INV_X1 U16196 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17854) );
  INV_X1 U16197 ( .A(n17517), .ZN(n17513) );
  NAND2_X1 U16198 ( .A1(n17656), .A2(n17513), .ZN(n12973) );
  OAI211_X1 U16199 ( .C1(n12974), .C2(n17854), .A(n12973), .B(n10070), .ZN(
        n17493) );
  NOR2_X1 U16200 ( .A1(n12974), .A2(n17656), .ZN(n17512) );
  NAND2_X1 U16201 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17834) );
  INV_X1 U16202 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17466) );
  NOR2_X2 U16203 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15728), .ZN(
        n12977) );
  NAND2_X1 U16204 ( .A1(n12977), .A2(n17656), .ZN(n15777) );
  INV_X1 U16205 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15782) );
  NAND2_X1 U16206 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n15782), .ZN(
        n16393) );
  INV_X1 U16207 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17829) );
  NOR2_X1 U16208 ( .A1(n17829), .A2(n17466), .ZN(n15721) );
  INV_X1 U16209 ( .A(n15721), .ZN(n15719) );
  INV_X1 U16210 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16383) );
  NOR2_X1 U16211 ( .A1(n15719), .A2(n16383), .ZN(n16392) );
  NAND2_X1 U16212 ( .A1(n12975), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17480) );
  NOR2_X2 U16213 ( .A1(n17656), .A2(n17480), .ZN(n16413) );
  NAND2_X1 U16214 ( .A1(n16392), .A2(n16413), .ZN(n15776) );
  INV_X1 U16215 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18772) );
  NAND2_X1 U16216 ( .A1(n18772), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12976) );
  OAI211_X1 U16217 ( .C1(n17730), .C2(n12977), .A(n15776), .B(n12976), .ZN(
        n12978) );
  AOI21_X1 U16218 ( .B1(n17730), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n18772), .ZN(n12980) );
  AND2_X1 U16219 ( .A1(n17730), .A2(n18772), .ZN(n12979) );
  NOR2_X1 U16220 ( .A1(n12980), .A2(n12979), .ZN(n12981) );
  NAND2_X1 U16221 ( .A1(n9732), .A2(n12991), .ZN(n12986) );
  OAI21_X1 U16222 ( .B1(n12986), .B2(n12985), .A(n12984), .ZN(n12987) );
  NOR2_X1 U16223 ( .A1(n12989), .A2(n12988), .ZN(n18826) );
  NOR2_X1 U16224 ( .A1(n18164), .A2(n12990), .ZN(n15709) );
  NAND2_X1 U16225 ( .A1(n15709), .A2(n17211), .ZN(n15711) );
  INV_X1 U16226 ( .A(n12992), .ZN(n12994) );
  NOR2_X1 U16227 ( .A1(n12994), .A2(n12993), .ZN(n12995) );
  OAI211_X1 U16228 ( .C1(n18178), .C2(n18630), .A(n9832), .B(n12995), .ZN(
        n15695) );
  INV_X1 U16229 ( .A(n12996), .ZN(n12999) );
  OAI21_X1 U16230 ( .B1(n12999), .B2(n12998), .A(n12997), .ZN(n18599) );
  NOR2_X2 U16231 ( .A1(n16521), .A2(n18164), .ZN(n17797) );
  NAND2_X1 U16232 ( .A1(n16399), .A2(n17731), .ZN(n13044) );
  OAI21_X1 U16233 ( .B1(n18773), .B2(n18661), .A(n18763), .ZN(n18149) );
  OAI21_X4 U16234 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18149), .A(n16521), 
        .ZN(n17822) );
  NAND3_X2 U16235 ( .A1(n18813), .A2(n17822), .A3(P3_STATE2_REG_1__SCAN_IN), 
        .ZN(n17666) );
  NOR2_X1 U16236 ( .A1(n18749), .A2(n18141), .ZN(n16396) );
  NAND2_X1 U16237 ( .A1(n13000), .A2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13001) );
  NAND2_X1 U16238 ( .A1(n14386), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17823) );
  NAND2_X1 U16239 ( .A1(n18604), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18775) );
  OAI221_X1 U16240 ( .B1(n18661), .B2(P3_STATE2_REG_1__SCAN_IN), .C1(
        P3_STATE2_REG_2__SCAN_IN), .C2(n18773), .A(n18775), .ZN(n18158) );
  NAND3_X1 U16241 ( .A1(n18661), .A2(n18763), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18239) );
  OR2_X1 U16242 ( .A1(n13001), .A2(n17661), .ZN(n16369) );
  XNOR2_X1 U16243 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n13005) );
  INV_X1 U16244 ( .A(n17548), .ZN(n17577) );
  NOR2_X1 U16245 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17577), .ZN(
        n16387) );
  NAND2_X1 U16246 ( .A1(n18539), .A2(n13001), .ZN(n13002) );
  OAI211_X1 U16247 ( .C1(n13003), .C2(n17823), .A(n17822), .B(n13002), .ZN(
        n16380) );
  NOR2_X1 U16248 ( .A1(n16387), .A2(n16380), .ZN(n16368) );
  OAI22_X1 U16249 ( .A1(n16369), .A2(n13005), .B1(n16368), .B2(n13004), .ZN(
        n13006) );
  AOI211_X1 U16250 ( .C1(n17675), .C2(n16805), .A(n16396), .B(n13006), .ZN(
        n13043) );
  INV_X1 U16251 ( .A(n17653), .ZN(n17632) );
  AND2_X1 U16252 ( .A1(n17524), .A2(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15718) );
  NAND2_X1 U16253 ( .A1(n17885), .A2(n15718), .ZN(n17511) );
  NOR2_X1 U16254 ( .A1(n17854), .A2(n17511), .ZN(n17510) );
  NAND2_X1 U16255 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17510), .ZN(
        n15720) );
  NAND2_X1 U16256 ( .A1(n17837), .A2(n16392), .ZN(n16386) );
  INV_X1 U16257 ( .A(n16386), .ZN(n16372) );
  NAND2_X1 U16258 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16372), .ZN(
        n13008) );
  XOR2_X1 U16259 ( .A(n18772), .B(n13008), .Z(n16400) );
  NAND2_X1 U16260 ( .A1(n16400), .A2(n17690), .ZN(n13042) );
  NAND2_X1 U16261 ( .A1(n17346), .A2(n15811), .ZN(n13014) );
  NAND2_X1 U16262 ( .A1(n17341), .A2(n13014), .ZN(n13012) );
  AND2_X1 U16263 ( .A1(n13013), .A2(n13012), .ZN(n13024) );
  NAND2_X1 U16264 ( .A1(n13009), .A2(n13010), .ZN(n13028) );
  NOR2_X1 U16265 ( .A1(n17326), .A2(n13028), .ZN(n13032) );
  NAND2_X1 U16266 ( .A1(n13032), .A2(n16409), .ZN(n13033) );
  XOR2_X1 U16267 ( .A(n13010), .B(n13009), .Z(n13011) );
  AND2_X1 U16268 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13011), .ZN(
        n13027) );
  XOR2_X1 U16269 ( .A(n18086), .B(n13011), .Z(n17764) );
  XNOR2_X1 U16270 ( .A(n13013), .B(n13012), .ZN(n13022) );
  NOR2_X1 U16271 ( .A1(n15717), .A2(n13022), .ZN(n13023) );
  XNOR2_X1 U16272 ( .A(n13015), .B(n13014), .ZN(n13017) );
  NOR2_X1 U16273 ( .A1(n13017), .A2(n13016), .ZN(n13021) );
  XOR2_X1 U16274 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n13017), .Z(
        n17803) );
  NOR2_X1 U16275 ( .A1(n13019), .A2(n18790), .ZN(n13020) );
  NAND3_X1 U16276 ( .A1(n17821), .A2(n13019), .A3(n18790), .ZN(n13018) );
  OAI221_X1 U16277 ( .B1(n13020), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n17821), .C2(n13019), .A(n13018), .ZN(n17802) );
  NOR2_X1 U16278 ( .A1(n17803), .A2(n17802), .ZN(n17801) );
  NOR2_X1 U16279 ( .A1(n13021), .A2(n17801), .ZN(n17788) );
  XOR2_X1 U16280 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n13022), .Z(
        n17787) );
  NOR2_X1 U16281 ( .A1(n17788), .A2(n17787), .ZN(n17786) );
  NOR2_X1 U16282 ( .A1(n13023), .A2(n17786), .ZN(n17776) );
  XNOR2_X1 U16283 ( .A(n13025), .B(n13024), .ZN(n17777) );
  NOR2_X1 U16284 ( .A1(n17776), .A2(n17777), .ZN(n13026) );
  NAND2_X1 U16285 ( .A1(n17776), .A2(n17777), .ZN(n17775) );
  OAI21_X1 U16286 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n13026), .A(
        n17775), .ZN(n17763) );
  NOR2_X1 U16287 ( .A1(n17764), .A2(n17763), .ZN(n17762) );
  XNOR2_X1 U16288 ( .A(n17326), .B(n13028), .ZN(n13030) );
  NOR2_X1 U16289 ( .A1(n13029), .A2(n13030), .ZN(n13031) );
  INV_X1 U16290 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18077) );
  XNOR2_X1 U16291 ( .A(n13030), .B(n13029), .ZN(n17748) );
  NOR2_X1 U16292 ( .A1(n18077), .A2(n17748), .ZN(n17747) );
  NOR2_X1 U16293 ( .A1(n13031), .A2(n17747), .ZN(n13034) );
  XOR2_X1 U16294 ( .A(n17322), .B(n13032), .Z(n13035) );
  NAND2_X1 U16295 ( .A1(n13034), .A2(n13035), .ZN(n17736) );
  NAND2_X1 U16296 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17736), .ZN(
        n13037) );
  NOR2_X1 U16297 ( .A1(n13033), .A2(n13037), .ZN(n13039) );
  INV_X1 U16298 ( .A(n13033), .ZN(n13038) );
  OR2_X1 U16299 ( .A1(n13035), .A2(n13034), .ZN(n17737) );
  OAI21_X1 U16300 ( .B1(n13038), .B2(n13037), .A(n17737), .ZN(n13036) );
  AOI21_X1 U16301 ( .B1(n13038), .B2(n13037), .A(n13036), .ZN(n17728) );
  NAND2_X1 U16302 ( .A1(n15718), .A2(n17971), .ZN(n17502) );
  NAND3_X1 U16303 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n17830), .A3(
        n16392), .ZN(n13040) );
  XNOR2_X1 U16304 ( .A(n18772), .B(n13040), .ZN(n16402) );
  NOR2_X4 U16305 ( .A1(n9732), .A2(n16521), .ZN(n17815) );
  OR2_X1 U16306 ( .A1(n16402), .A2(n17827), .ZN(n13041) );
  NAND2_X1 U16307 ( .A1(n13044), .A2(n10072), .ZN(P3_U2799) );
  NOR2_X1 U16308 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13046) );
  NOR4_X1 U16309 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13045) );
  NAND4_X1 U16310 ( .A1(n13046), .A2(P2_W_R_N_REG_SCAN_IN), .A3(
        P2_M_IO_N_REG_SCAN_IN), .A4(n13045), .ZN(n13050) );
  NOR4_X1 U16311 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(P1_BE_N_REG_1__SCAN_IN), .A4(P1_BE_N_REG_3__SCAN_IN), .ZN(n13049)
         );
  NAND2_X1 U16312 ( .A1(P1_M_IO_N_REG_SCAN_IN), .A2(P1_W_R_N_REG_SCAN_IN), 
        .ZN(n13047) );
  NOR3_X1 U16313 ( .A1(P1_D_C_N_REG_SCAN_IN), .A2(P1_ADS_N_REG_SCAN_IN), .A3(
        n13047), .ZN(n13048) );
  NAND3_X1 U16314 ( .A1(n20099), .A2(n13049), .A3(n13048), .ZN(U214) );
  NOR2_X1 U16315 ( .A1(n13861), .A2(n13050), .ZN(n16424) );
  NAND2_X1 U16316 ( .A1(n16424), .A2(U214), .ZN(U212) );
  AOI211_X1 U16317 ( .C1(n15271), .C2(n13052), .A(n13051), .B(n19677), .ZN(
        n13064) );
  INV_X1 U16318 ( .A(n13053), .ZN(n13054) );
  OAI22_X1 U16319 ( .A1(n13054), .A2(n18984), .B1(n19737), .B2(n18978), .ZN(
        n13063) );
  INV_X1 U16320 ( .A(n19018), .ZN(n19002) );
  INV_X1 U16321 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n13055) );
  OAI22_X1 U16322 ( .A1(n19002), .A2(n13055), .B1(n15269), .B2(n19028), .ZN(
        n13062) );
  INV_X1 U16323 ( .A(n13056), .ZN(n13058) );
  OAI21_X1 U16324 ( .B1(n13058), .B2(n9985), .A(n15152), .ZN(n15470) );
  AND2_X1 U16325 ( .A1(n13089), .A2(n13059), .ZN(n13060) );
  OR2_X1 U16326 ( .A1(n13060), .A2(n15456), .ZN(n15474) );
  OAI22_X1 U16327 ( .A1(n15470), .A2(n19004), .B1(n15474), .B2(n19001), .ZN(
        n13061) );
  AOI211_X1 U16328 ( .C1(n15229), .C2(n13066), .A(n13065), .B(n19677), .ZN(
        n13079) );
  OAI22_X1 U16329 ( .A1(n13067), .A2(n18984), .B1(n19746), .B2(n18978), .ZN(
        n13078) );
  INV_X1 U16330 ( .A(P2_EBX_REG_27__SCAN_IN), .ZN(n13068) );
  OAI22_X1 U16331 ( .A1(n19002), .A2(n13068), .B1(n15231), .B2(n19028), .ZN(
        n13077) );
  INV_X1 U16332 ( .A(n13069), .ZN(n13070) );
  AOI21_X1 U16333 ( .B1(n13071), .B2(n15137), .A(n13070), .ZN(n15424) );
  INV_X1 U16334 ( .A(n15424), .ZN(n13075) );
  NAND2_X1 U16335 ( .A1(n15192), .A2(n13072), .ZN(n13073) );
  NAND2_X1 U16336 ( .A1(n13074), .A2(n13073), .ZN(n15421) );
  OAI22_X1 U16337 ( .A1(n13075), .A2(n19004), .B1(n15421), .B2(n19001), .ZN(
        n13076) );
  AOI211_X1 U16338 ( .C1(n13081), .C2(n9858), .A(n13080), .B(n19677), .ZN(
        n13093) );
  OAI22_X1 U16339 ( .A1(n13082), .A2(n18984), .B1(n19735), .B2(n18978), .ZN(
        n13092) );
  AOI22_X1 U16340 ( .A1(n19018), .A2(P2_EBX_REG_22__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n18997), .ZN(n13083) );
  INV_X1 U16341 ( .A(n13083), .ZN(n13091) );
  OR2_X1 U16342 ( .A1(n15168), .A2(n13084), .ZN(n13085) );
  NAND2_X1 U16343 ( .A1(n13056), .A2(n13085), .ZN(n15485) );
  NAND2_X1 U16344 ( .A1(n13086), .A2(n13087), .ZN(n13088) );
  NAND2_X1 U16345 ( .A1(n13089), .A2(n13088), .ZN(n15489) );
  OAI22_X1 U16346 ( .A1(n15485), .A2(n19004), .B1(n15489), .B2(n19001), .ZN(
        n13090) );
  OR4_X1 U16347 ( .A1(n13093), .A2(n13092), .A3(n13091), .A4(n13090), .ZN(
        P2_U2833) );
  NOR2_X1 U16348 ( .A1(n14582), .A2(n20120), .ZN(n15732) );
  NAND2_X1 U16349 ( .A1(n15762), .A2(n20120), .ZN(n13284) );
  INV_X1 U16350 ( .A(n13284), .ZN(n13096) );
  OR2_X1 U16351 ( .A1(n15732), .A2(n13096), .ZN(n13100) );
  INV_X1 U16352 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n13097) );
  NAND2_X1 U16353 ( .A1(n13098), .A2(n13097), .ZN(n15788) );
  INV_X1 U16354 ( .A(n15788), .ZN(n14592) );
  AND2_X1 U16355 ( .A1(n13262), .A2(n14592), .ZN(n13099) );
  AND2_X1 U16356 ( .A1(n13100), .A2(n13099), .ZN(n19950) );
  NAND2_X1 U16357 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16163) );
  NOR2_X1 U16358 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16163), .ZN(n19968) );
  AND2_X1 U16359 ( .A1(n19962), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  INV_X1 U16360 ( .A(n10673), .ZN(n13101) );
  NAND2_X1 U16361 ( .A1(n13102), .A2(n13101), .ZN(n19005) );
  INV_X1 U16362 ( .A(n19005), .ZN(n19029) );
  INV_X1 U16363 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13103) );
  INV_X1 U16364 ( .A(n13112), .ZN(n13111) );
  NAND2_X1 U16365 ( .A1(n19764), .A2(n13937), .ZN(n13104) );
  OAI211_X1 U16366 ( .C1(n19029), .C2(n13103), .A(n13111), .B(n13104), .ZN(
        P2_U2814) );
  NOR2_X1 U16367 ( .A1(n19819), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n13105)
         );
  AOI22_X1 U16368 ( .A1(n19819), .A2(n13106), .B1(n13105), .B2(n13104), .ZN(
        P2_U3612) );
  NOR2_X1 U16369 ( .A1(n13157), .A2(n13107), .ZN(n13108) );
  NAND2_X1 U16370 ( .A1(n16323), .A2(n13108), .ZN(n13109) );
  NOR2_X1 U16371 ( .A1(n16324), .A2(n13109), .ZN(n16333) );
  NOR2_X1 U16372 ( .A1(n16333), .A2(n16361), .ZN(n19805) );
  OAI21_X1 U16373 ( .B1(n19805), .B2(n15806), .A(n13110), .ZN(P2_U2819) );
  INV_X1 U16374 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n13114) );
  NAND3_X1 U16375 ( .A1(n13112), .A2(n10173), .A3(n19825), .ZN(n13226) );
  AOI22_X1 U16376 ( .A1(n13863), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n13190), .ZN(n19097) );
  NOR2_X1 U16377 ( .A1(n13226), .A2(n19097), .ZN(n13199) );
  AOI21_X1 U16378 ( .B1(P2_EAX_REG_3__SCAN_IN), .B2(n13211), .A(n13199), .ZN(
        n13113) );
  OAI21_X1 U16379 ( .B1(n13176), .B2(n13114), .A(n13113), .ZN(P2_U2970) );
  INV_X1 U16380 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n13116) );
  AOI22_X1 U16381 ( .A1(n13863), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n13190), .ZN(n19065) );
  NOR2_X1 U16382 ( .A1(n13226), .A2(n19065), .ZN(n13187) );
  AOI21_X1 U16383 ( .B1(n13211), .B2(P2_EAX_REG_7__SCAN_IN), .A(n13187), .ZN(
        n13115) );
  OAI21_X1 U16384 ( .B1(n13176), .B2(n13116), .A(n13115), .ZN(P2_U2974) );
  INV_X1 U16385 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n13118) );
  OAI22_X1 U16386 ( .A1(n13190), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n13863), .ZN(n13537) );
  NOR2_X1 U16387 ( .A1(n13226), .A2(n13537), .ZN(n13193) );
  AOI21_X1 U16388 ( .B1(P2_EAX_REG_2__SCAN_IN), .B2(n13211), .A(n13193), .ZN(
        n13117) );
  OAI21_X1 U16389 ( .B1(n13176), .B2(n13118), .A(n13117), .ZN(P2_U2969) );
  INV_X1 U16390 ( .A(P2_LWORD_REG_14__SCAN_IN), .ZN(n13121) );
  INV_X1 U16391 ( .A(n13226), .ZN(n13148) );
  INV_X1 U16392 ( .A(n19049), .ZN(n13119) );
  NAND2_X1 U16393 ( .A1(n13148), .A2(n13119), .ZN(n13142) );
  NAND2_X1 U16394 ( .A1(n13211), .A2(P2_EAX_REG_14__SCAN_IN), .ZN(n13120) );
  OAI211_X1 U16395 ( .C1(n13176), .C2(n13121), .A(n13142), .B(n13120), .ZN(
        P2_U2981) );
  INV_X1 U16396 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n13123) );
  OAI22_X1 U16397 ( .A1(n13190), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n13863), .ZN(n13302) );
  INV_X1 U16398 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13122) );
  OAI222_X1 U16399 ( .A1(n13123), .A2(n13176), .B1(n13226), .B2(n13302), .C1(
        n13225), .C2(n13122), .ZN(P2_U2967) );
  INV_X1 U16400 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14572) );
  NAND2_X1 U16401 ( .A1(n13152), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13128) );
  INV_X1 U16402 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n13124) );
  OR2_X1 U16403 ( .A1(n13190), .A2(n13124), .ZN(n13126) );
  NAND2_X1 U16404 ( .A1(n13861), .A2(BUF2_REG_13__SCAN_IN), .ZN(n13125) );
  AND2_X1 U16405 ( .A1(n13126), .A2(n13125), .ZN(n19051) );
  INV_X1 U16406 ( .A(n19051), .ZN(n13127) );
  NAND2_X1 U16407 ( .A1(n13148), .A2(n13127), .ZN(n13203) );
  OAI211_X1 U16408 ( .C1(n13225), .C2(n14572), .A(n13128), .B(n13203), .ZN(
        P2_U2965) );
  NAND2_X1 U16409 ( .A1(n13152), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n13129) );
  MUX2_X1 U16410 ( .A(BUF1_REG_10__SCAN_IN), .B(BUF2_REG_10__SCAN_IN), .S(
        n13861), .Z(n19057) );
  NAND2_X1 U16411 ( .A1(n13148), .A2(n19057), .ZN(n13150) );
  OAI211_X1 U16412 ( .C1(n10980), .C2(n13225), .A(n13129), .B(n13150), .ZN(
        P2_U2977) );
  NAND2_X1 U16413 ( .A1(n13152), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n13131) );
  AOI22_X1 U16414 ( .A1(n13863), .A2(BUF1_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n13190), .ZN(n19053) );
  INV_X1 U16415 ( .A(n19053), .ZN(n13130) );
  NAND2_X1 U16416 ( .A1(n13148), .A2(n13130), .ZN(n13133) );
  OAI211_X1 U16417 ( .C1(n13225), .C2(n13132), .A(n13131), .B(n13133), .ZN(
        P2_U2979) );
  INV_X1 U16418 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n15176) );
  NAND2_X1 U16419 ( .A1(n13152), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13134) );
  OAI211_X1 U16420 ( .C1(n13225), .C2(n15176), .A(n13134), .B(n13133), .ZN(
        P2_U2964) );
  INV_X1 U16421 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n15181) );
  NAND2_X1 U16422 ( .A1(n13152), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13138) );
  INV_X1 U16423 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n14321) );
  OR2_X1 U16424 ( .A1(n13190), .A2(n14321), .ZN(n13136) );
  NAND2_X1 U16425 ( .A1(n13861), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13135) );
  AND2_X1 U16426 ( .A1(n13136), .A2(n13135), .ZN(n19055) );
  INV_X1 U16427 ( .A(n19055), .ZN(n13137) );
  NAND2_X1 U16428 ( .A1(n13148), .A2(n13137), .ZN(n13209) );
  OAI211_X1 U16429 ( .C1(n13225), .C2(n15181), .A(n13138), .B(n13209), .ZN(
        P2_U2963) );
  NAND2_X1 U16430 ( .A1(n13152), .A2(P2_UWORD_REG_1__SCAN_IN), .ZN(n13140) );
  AOI22_X1 U16431 ( .A1(n13863), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n13861), .ZN(n19108) );
  INV_X1 U16432 ( .A(n19108), .ZN(n13139) );
  NAND2_X1 U16433 ( .A1(n13148), .A2(n13139), .ZN(n13213) );
  OAI211_X1 U16434 ( .C1(n13225), .C2(n14228), .A(n13140), .B(n13213), .ZN(
        P2_U2953) );
  INV_X1 U16435 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n13447) );
  NAND2_X1 U16436 ( .A1(n13152), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13141) );
  INV_X1 U16437 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16461) );
  INV_X1 U16438 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17444) );
  AOI22_X1 U16439 ( .A1(n13863), .A2(n16461), .B1(n17444), .B2(n13861), .ZN(
        n19062) );
  NAND2_X1 U16440 ( .A1(n13148), .A2(n19062), .ZN(n13153) );
  OAI211_X1 U16441 ( .C1(n13447), .C2(n13225), .A(n13141), .B(n13153), .ZN(
        P2_U2960) );
  NAND2_X1 U16442 ( .A1(n13152), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13143) );
  OAI211_X1 U16443 ( .C1(n13225), .C2(n13442), .A(n13143), .B(n13142), .ZN(
        P2_U2966) );
  INV_X1 U16444 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n15197) );
  NAND2_X1 U16445 ( .A1(n13152), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13149) );
  INV_X1 U16446 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n13144) );
  OR2_X1 U16447 ( .A1(n13861), .A2(n13144), .ZN(n13146) );
  NAND2_X1 U16448 ( .A1(n13861), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13145) );
  AND2_X1 U16449 ( .A1(n13146), .A2(n13145), .ZN(n19060) );
  INV_X1 U16450 ( .A(n19060), .ZN(n13147) );
  NAND2_X1 U16451 ( .A1(n13148), .A2(n13147), .ZN(n13206) );
  OAI211_X1 U16452 ( .C1(n13225), .C2(n15197), .A(n13149), .B(n13206), .ZN(
        P2_U2961) );
  INV_X1 U16453 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n13222) );
  NAND2_X1 U16454 ( .A1(n13152), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13151) );
  OAI211_X1 U16455 ( .C1(n13222), .C2(n13225), .A(n13151), .B(n13150), .ZN(
        P2_U2962) );
  INV_X1 U16456 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19123) );
  NAND2_X1 U16457 ( .A1(n13152), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13154) );
  OAI211_X1 U16458 ( .C1(n19123), .C2(n13225), .A(n13154), .B(n13153), .ZN(
        P2_U2975) );
  OR2_X1 U16459 ( .A1(n10673), .A2(n13155), .ZN(n13156) );
  OR2_X1 U16460 ( .A1(n13216), .A2(n13156), .ZN(n13163) );
  NAND2_X1 U16461 ( .A1(n16323), .A2(n13157), .ZN(n13158) );
  NOR2_X1 U16462 ( .A1(n16324), .A2(n13158), .ZN(n13159) );
  NOR2_X1 U16463 ( .A1(n13160), .A2(n13159), .ZN(n13162) );
  OR2_X1 U16464 ( .A1(n16328), .A2(n16326), .ZN(n13498) );
  NAND4_X1 U16465 ( .A1(n13163), .A2(n13162), .A3(n13498), .A4(n13161), .ZN(
        n16340) );
  NAND2_X1 U16466 ( .A1(n16340), .A2(n19673), .ZN(n13166) );
  NAND2_X1 U16467 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19799), .ZN(n16363) );
  NOR2_X1 U16468 ( .A1(n15806), .A2(n16363), .ZN(n13164) );
  AOI21_X1 U16469 ( .B1(n19822), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n13164), 
        .ZN(n13165) );
  INV_X1 U16470 ( .A(n13975), .ZN(n13170) );
  INV_X1 U16471 ( .A(n13167), .ZN(n13168) );
  NOR2_X1 U16472 ( .A1(n10673), .A2(n13168), .ZN(n16334) );
  NAND4_X1 U16473 ( .A1(n13170), .A2(n19829), .A3(n16334), .A4(n19763), .ZN(
        n13169) );
  OAI21_X1 U16474 ( .B1(n16339), .B2(n13170), .A(n13169), .ZN(P2_U3595) );
  INV_X1 U16475 ( .A(n14581), .ZN(n13171) );
  NOR2_X1 U16476 ( .A1(n14582), .A2(n13171), .ZN(n14587) );
  NAND2_X1 U16477 ( .A1(n14587), .A2(n14598), .ZN(n19840) );
  INV_X1 U16478 ( .A(n20758), .ZN(n13174) );
  NOR2_X2 U16479 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20602) );
  NAND2_X1 U16480 ( .A1(n13902), .A2(n20602), .ZN(n19847) );
  INV_X1 U16481 ( .A(n19847), .ZN(n13172) );
  OAI21_X1 U16482 ( .B1(P1_READREQUEST_REG_SCAN_IN), .B2(n13172), .A(n13174), 
        .ZN(n13173) );
  OAI21_X1 U16483 ( .B1(n13175), .B2(n13174), .A(n13173), .ZN(P1_U3487) );
  INV_X1 U16484 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n13178) );
  AOI22_X1 U16485 ( .A1(n13863), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n13190), .ZN(n19068) );
  NOR2_X1 U16486 ( .A1(n13226), .A2(n19068), .ZN(n13181) );
  AOI21_X1 U16487 ( .B1(n13211), .B2(P2_EAX_REG_6__SCAN_IN), .A(n13181), .ZN(
        n13177) );
  OAI21_X1 U16488 ( .B1(n13224), .B2(n13178), .A(n13177), .ZN(P2_U2973) );
  INV_X1 U16489 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n13180) );
  OAI22_X1 U16490 ( .A1(n13861), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n13863), .ZN(n19090) );
  NOR2_X1 U16491 ( .A1(n13226), .A2(n19090), .ZN(n13184) );
  AOI21_X1 U16492 ( .B1(n13211), .B2(P2_EAX_REG_20__SCAN_IN), .A(n13184), .ZN(
        n13179) );
  OAI21_X1 U16493 ( .B1(n13224), .B2(n13180), .A(n13179), .ZN(P2_U2956) );
  INV_X1 U16494 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n13183) );
  AOI21_X1 U16495 ( .B1(n13211), .B2(P2_EAX_REG_22__SCAN_IN), .A(n13181), .ZN(
        n13182) );
  OAI21_X1 U16496 ( .B1(n13224), .B2(n13183), .A(n13182), .ZN(P2_U2958) );
  INV_X1 U16497 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n13186) );
  AOI21_X1 U16498 ( .B1(P2_EAX_REG_4__SCAN_IN), .B2(n13211), .A(n13184), .ZN(
        n13185) );
  OAI21_X1 U16499 ( .B1(n13224), .B2(n13186), .A(n13185), .ZN(P2_U2971) );
  INV_X1 U16500 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n13189) );
  AOI21_X1 U16501 ( .B1(n13211), .B2(P2_EAX_REG_23__SCAN_IN), .A(n13187), .ZN(
        n13188) );
  OAI21_X1 U16502 ( .B1(n13224), .B2(n13189), .A(n13188), .ZN(P2_U2959) );
  INV_X1 U16503 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n13192) );
  AOI22_X1 U16504 ( .A1(n13863), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n13190), .ZN(n14258) );
  NOR2_X1 U16505 ( .A1(n13226), .A2(n14258), .ZN(n13196) );
  AOI21_X1 U16506 ( .B1(n13211), .B2(P2_EAX_REG_5__SCAN_IN), .A(n13196), .ZN(
        n13191) );
  OAI21_X1 U16507 ( .B1(n13224), .B2(n13192), .A(n13191), .ZN(P2_U2972) );
  INV_X1 U16508 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n13195) );
  AOI21_X1 U16509 ( .B1(n13211), .B2(P2_EAX_REG_18__SCAN_IN), .A(n13193), .ZN(
        n13194) );
  OAI21_X1 U16510 ( .B1(n13224), .B2(n13195), .A(n13194), .ZN(P2_U2954) );
  INV_X1 U16511 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n13198) );
  AOI21_X1 U16512 ( .B1(n13211), .B2(P2_EAX_REG_21__SCAN_IN), .A(n13196), .ZN(
        n13197) );
  OAI21_X1 U16513 ( .B1(n13224), .B2(n13198), .A(n13197), .ZN(P2_U2957) );
  INV_X1 U16514 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n13201) );
  AOI21_X1 U16515 ( .B1(n13211), .B2(P2_EAX_REG_19__SCAN_IN), .A(n13199), .ZN(
        n13200) );
  OAI21_X1 U16516 ( .B1(n13224), .B2(n13201), .A(n13200), .ZN(P2_U2955) );
  INV_X1 U16517 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n13204) );
  NAND2_X1 U16518 ( .A1(n13211), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n13202) );
  OAI211_X1 U16519 ( .C1(n13224), .C2(n13204), .A(n13203), .B(n13202), .ZN(
        P2_U2980) );
  INV_X1 U16520 ( .A(P2_LWORD_REG_9__SCAN_IN), .ZN(n13207) );
  NAND2_X1 U16521 ( .A1(n13211), .A2(P2_EAX_REG_9__SCAN_IN), .ZN(n13205) );
  OAI211_X1 U16522 ( .C1(n13224), .C2(n13207), .A(n13206), .B(n13205), .ZN(
        P2_U2976) );
  INV_X1 U16523 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n13210) );
  NAND2_X1 U16524 ( .A1(n13211), .A2(P2_EAX_REG_11__SCAN_IN), .ZN(n13208) );
  OAI211_X1 U16525 ( .C1(n13224), .C2(n13210), .A(n13209), .B(n13208), .ZN(
        P2_U2978) );
  INV_X1 U16526 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n13214) );
  NAND2_X1 U16527 ( .A1(n13211), .A2(P2_EAX_REG_1__SCAN_IN), .ZN(n13212) );
  OAI211_X1 U16528 ( .C1(n13224), .C2(n13214), .A(n13213), .B(n13212), .ZN(
        P2_U2968) );
  OR2_X1 U16529 ( .A1(n10673), .A2(n16361), .ZN(n13215) );
  OAI21_X1 U16530 ( .B1(n13216), .B2(n13215), .A(n13225), .ZN(n13217) );
  NAND2_X1 U16531 ( .A1(n19109), .A2(n19830), .ZN(n13454) );
  AND2_X2 U16532 ( .A1(n19822), .A2(n19799), .ZN(n19821) );
  NOR2_X4 U16533 ( .A1(n19109), .A2(n19821), .ZN(n19126) );
  AOI22_X1 U16534 ( .A1(n19821), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n13218) );
  OAI21_X1 U16535 ( .B1(n15197), .B2(n13454), .A(n13218), .ZN(P2_U2926) );
  AOI22_X1 U16536 ( .A1(n19821), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n13219) );
  OAI21_X1 U16537 ( .B1(n14572), .B2(n13454), .A(n13219), .ZN(P2_U2922) );
  AOI22_X1 U16538 ( .A1(n19821), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n13220) );
  OAI21_X1 U16539 ( .B1(n15176), .B2(n13454), .A(n13220), .ZN(P2_U2923) );
  AOI22_X1 U16540 ( .A1(n19821), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n13221) );
  OAI21_X1 U16541 ( .B1(n13222), .B2(n13454), .A(n13221), .ZN(P2_U2925) );
  INV_X1 U16542 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n20881) );
  AOI22_X1 U16543 ( .A1(n13863), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n13861), .ZN(n19047) );
  INV_X1 U16544 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n19111) );
  OAI222_X1 U16545 ( .A1(n13224), .A2(n20881), .B1(n13226), .B2(n19047), .C1(
        n13225), .C2(n19111), .ZN(P2_U2982) );
  INV_X1 U16546 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n13223) );
  OAI222_X1 U16547 ( .A1(n13226), .A2(n13302), .B1(n13225), .B2(n11055), .C1(
        n13224), .C2(n13223), .ZN(P2_U2952) );
  INV_X1 U16548 ( .A(n13227), .ZN(n15669) );
  AND2_X1 U16549 ( .A1(n18902), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13308) );
  NOR2_X1 U16550 ( .A1(n13229), .A2(n13228), .ZN(n13230) );
  OR2_X1 U16551 ( .A1(n13231), .A2(n13230), .ZN(n19014) );
  OAI22_X1 U16552 ( .A1(n10247), .A2(n19179), .B1(n19185), .B2(n19014), .ZN(
        n13232) );
  AOI211_X1 U16553 ( .C1(n15669), .C2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13308), .B(n13232), .ZN(n13238) );
  OAI21_X1 U16554 ( .B1(n13234), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13233), .ZN(n13306) );
  OR2_X1 U16555 ( .A1(n19021), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13235) );
  NAND2_X1 U16556 ( .A1(n13322), .A2(n13235), .ZN(n13305) );
  OAI22_X1 U16557 ( .A1(n19174), .A2(n13306), .B1(n19157), .B2(n13305), .ZN(
        n13236) );
  AOI21_X1 U16558 ( .B1(n13938), .B2(n15671), .A(n13236), .ZN(n13237) );
  NAND2_X1 U16559 ( .A1(n13238), .A2(n13237), .ZN(P2_U3046) );
  INV_X1 U16560 ( .A(n19841), .ZN(n13239) );
  NAND2_X2 U16561 ( .A1(n13239), .A2(n20120), .ZN(n20088) );
  INV_X1 U16562 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n13245) );
  INV_X1 U16563 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13244) );
  AND2_X1 U16564 ( .A1(n14593), .A2(n20674), .ZN(n13240) );
  NOR2_X1 U16565 ( .A1(n19841), .A2(n13240), .ZN(n19973) );
  NAND2_X1 U16566 ( .A1(n13907), .A2(n20760), .ZN(n13241) );
  OR2_X1 U16567 ( .A1(n19841), .A2(n13241), .ZN(n19971) );
  INV_X1 U16568 ( .A(DATAI_15_), .ZN(n13243) );
  INV_X1 U16569 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13242) );
  MUX2_X1 U16570 ( .A(n13243), .B(n13242), .S(n20099), .Z(n14378) );
  OAI222_X1 U16571 ( .A1(n20088), .A2(n13245), .B1(n13244), .B2(n19973), .C1(
        n19971), .C2(n14378), .ZN(P1_U2967) );
  INV_X1 U16572 ( .A(n14145), .ZN(n13716) );
  OR2_X1 U16573 ( .A1(n13249), .A2(n13716), .ZN(n13248) );
  NAND2_X1 U16574 ( .A1(n20105), .A2(n13246), .ZN(n13473) );
  OAI21_X1 U16575 ( .B1(n14593), .B2(n13471), .A(n13473), .ZN(n13247) );
  INV_X1 U16576 ( .A(n13247), .ZN(n13250) );
  AND2_X1 U16577 ( .A1(n13248), .A2(n13250), .ZN(n13253) );
  INV_X1 U16578 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n15018) );
  OR2_X1 U16579 ( .A1(n15018), .A2(n13250), .ZN(n13251) );
  AOI21_X1 U16580 ( .B1(n13253), .B2(n15018), .A(n9798), .ZN(n20094) );
  INV_X1 U16581 ( .A(n20094), .ZN(n13293) );
  OR2_X1 U16582 ( .A1(n11633), .A2(n20120), .ZN(n13271) );
  AND3_X1 U16583 ( .A1(n13254), .A2(n14596), .A3(n13271), .ZN(n13276) );
  OAI21_X1 U16584 ( .B1(n13401), .B2(n13276), .A(n14582), .ZN(n13361) );
  NAND2_X1 U16585 ( .A1(n13907), .A2(n15788), .ZN(n14595) );
  NAND4_X1 U16586 ( .A1(n14581), .A2(n13359), .A3(n20760), .A4(n14595), .ZN(
        n13257) );
  NOR2_X1 U16587 ( .A1(n11634), .A2(n20120), .ZN(n13255) );
  NAND2_X1 U16588 ( .A1(n14589), .A2(n13255), .ZN(n13256) );
  NAND3_X1 U16589 ( .A1(n13361), .A2(n13257), .A3(n13256), .ZN(n13258) );
  NAND2_X1 U16590 ( .A1(n13258), .A2(n14598), .ZN(n13264) );
  OAI21_X1 U16591 ( .B1(n13907), .B2(n14592), .A(n20760), .ZN(n13911) );
  OAI211_X1 U16592 ( .C1(n13259), .C2(n13911), .A(n14596), .B(n13260), .ZN(
        n13261) );
  NAND3_X1 U16593 ( .A1(n13262), .A2(n11635), .A3(n13261), .ZN(n13263) );
  NAND2_X1 U16594 ( .A1(n14588), .A2(n13400), .ZN(n13265) );
  NAND2_X1 U16595 ( .A1(n13266), .A2(n13265), .ZN(n14580) );
  NAND2_X1 U16596 ( .A1(n13283), .A2(n11569), .ZN(n13267) );
  AND2_X1 U16597 ( .A1(n14580), .A2(n13267), .ZN(n13268) );
  NAND2_X1 U16598 ( .A1(n13269), .A2(n13268), .ZN(n13270) );
  NOR2_X1 U16599 ( .A1(n13272), .A2(n13271), .ZN(n14578) );
  OAI21_X1 U16600 ( .B1(n13274), .B2(n14522), .A(n13273), .ZN(n13275) );
  INV_X1 U16601 ( .A(n13275), .ZN(n13278) );
  INV_X1 U16602 ( .A(n13276), .ZN(n13277) );
  OAI211_X1 U16603 ( .C1(n13280), .C2(n13279), .A(n13278), .B(n13277), .ZN(
        n13351) );
  OR2_X1 U16604 ( .A1(n13281), .A2(n13351), .ZN(n13282) );
  NAND2_X1 U16605 ( .A1(n13289), .A2(n13282), .ZN(n15019) );
  NAND2_X1 U16606 ( .A1(n15055), .A2(n15019), .ZN(n14547) );
  NAND2_X1 U16607 ( .A1(n13283), .A2(n11626), .ZN(n13285) );
  NAND2_X1 U16608 ( .A1(n13285), .A2(n13284), .ZN(n13286) );
  NOR2_X1 U16609 ( .A1(n14525), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13288) );
  INV_X1 U16610 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13287) );
  OAI22_X1 U16611 ( .A1(n13781), .A2(n13287), .B1(n14522), .B2(
        P1_EBX_REG_0__SCAN_IN), .ZN(n13414) );
  OR2_X1 U16612 ( .A1(n13288), .A2(n13414), .ZN(n19942) );
  NAND2_X1 U16613 ( .A1(n16052), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n20095) );
  OAI21_X1 U16614 ( .B1(n16068), .B2(n19942), .A(n20095), .ZN(n13291) );
  OR2_X1 U16615 ( .A1(n13289), .A2(n16141), .ZN(n13477) );
  NAND2_X1 U16616 ( .A1(n13289), .A2(n15732), .ZN(n15794) );
  AOI21_X1 U16617 ( .B1(n13477), .B2(n15794), .A(n15018), .ZN(n13290) );
  AOI211_X1 U16618 ( .C1(n15018), .C2(n14547), .A(n13291), .B(n13290), .ZN(
        n13292) );
  OAI21_X1 U16619 ( .B1(n13293), .B2(n16111), .A(n13292), .ZN(P1_U3031) );
  INV_X1 U16620 ( .A(n19099), .ZN(n19046) );
  AND2_X1 U16621 ( .A1(n19794), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n13294) );
  OAI211_X1 U16622 ( .C1(n19829), .C2(n13296), .A(n13295), .B(n13294), .ZN(
        n13297) );
  INV_X1 U16623 ( .A(n13297), .ZN(n13298) );
  NOR2_X1 U16624 ( .A1(n19796), .A2(n19014), .ZN(n19102) );
  AOI211_X1 U16625 ( .C1(n19796), .C2(n19014), .A(n19102), .B(n19103), .ZN(
        n13300) );
  AOI21_X1 U16626 ( .B1(P2_EAX_REG_0__SCAN_IN), .B2(n19098), .A(n13300), .ZN(
        n13304) );
  INV_X1 U16627 ( .A(n15206), .ZN(n19037) );
  INV_X1 U16628 ( .A(n13302), .ZN(n19036) );
  NAND2_X1 U16629 ( .A1(n19071), .A2(n19036), .ZN(n13303) );
  OAI211_X1 U16630 ( .C1(n19014), .C2(n19046), .A(n13304), .B(n13303), .ZN(
        P2_U2919) );
  INV_X1 U16631 ( .A(n13305), .ZN(n13309) );
  NOR2_X1 U16632 ( .A1(n19148), .A2(n13306), .ZN(n13307) );
  AOI211_X1 U16633 ( .C1(n11114), .C2(n13309), .A(n13308), .B(n13307), .ZN(
        n13312) );
  OAI21_X1 U16634 ( .B1(n15338), .B2(n13310), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13311) );
  OAI211_X1 U16635 ( .C1(n13862), .C2(n10247), .A(n13312), .B(n13311), .ZN(
        P2_U3014) );
  NAND2_X1 U16636 ( .A1(n14578), .A2(n14589), .ZN(n13370) );
  NAND4_X1 U16637 ( .A1(n13313), .A2(n11630), .A3(n13426), .A4(n14467), .ZN(
        n13314) );
  NAND2_X1 U16638 ( .A1(n13370), .A2(n13314), .ZN(n13315) );
  INV_X1 U16639 ( .A(n13316), .ZN(n13320) );
  INV_X1 U16640 ( .A(n13317), .ZN(n13319) );
  OAI21_X1 U16641 ( .B1(n13320), .B2(n13319), .A(n13318), .ZN(n20097) );
  INV_X2 U16642 ( .A(n15942), .ZN(n14750) );
  OAI222_X1 U16643 ( .A1(n19942), .A2(n14761), .B1(n13287), .B2(n15945), .C1(
        n20097), .C2(n14750), .ZN(P1_U2872) );
  OAI21_X1 U16644 ( .B1(n13830), .B2(n13322), .A(n13321), .ZN(n13323) );
  XNOR2_X1 U16645 ( .A(n13323), .B(n13958), .ZN(n15665) );
  AOI21_X1 U16646 ( .B1(n13958), .B2(n13325), .A(n13324), .ZN(n15670) );
  AND2_X1 U16647 ( .A1(n18902), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n15668) );
  NOR2_X1 U16648 ( .A1(n19154), .A2(n13826), .ZN(n13326) );
  AOI211_X1 U16649 ( .C1(n16261), .C2(n15670), .A(n15668), .B(n13326), .ZN(
        n13327) );
  OAI21_X1 U16650 ( .B1(n15396), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n13327), .ZN(n13328) );
  AOI21_X1 U16651 ( .B1(n19151), .B2(n13963), .A(n13328), .ZN(n13329) );
  OAI21_X1 U16652 ( .B1(n19147), .B2(n15665), .A(n13329), .ZN(P2_U3013) );
  INV_X1 U16653 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n20011) );
  NAND2_X1 U16654 ( .A1(n19950), .A2(n14596), .ZN(n13624) );
  AOI22_X1 U16655 ( .A1(n20761), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n19967), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13330) );
  OAI21_X1 U16656 ( .B1(n20011), .B2(n13624), .A(n13330), .ZN(P1_U2911) );
  INV_X1 U16657 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n20025) );
  AOI22_X1 U16658 ( .A1(n20761), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n19967), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13331) );
  OAI21_X1 U16659 ( .B1(n20025), .B2(n13624), .A(n13331), .ZN(P1_U2908) );
  INV_X1 U16660 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n20029) );
  AOI22_X1 U16661 ( .A1(n20761), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n19967), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13332) );
  OAI21_X1 U16662 ( .B1(n20029), .B2(n13624), .A(n13332), .ZN(P1_U2907) );
  INV_X1 U16663 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n20021) );
  AOI22_X1 U16664 ( .A1(n20761), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n19967), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13333) );
  OAI21_X1 U16665 ( .B1(n20021), .B2(n13624), .A(n13333), .ZN(P1_U2909) );
  INV_X1 U16666 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n20016) );
  AOI22_X1 U16667 ( .A1(n20761), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n19967), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13334) );
  OAI21_X1 U16668 ( .B1(n20016), .B2(n13624), .A(n13334), .ZN(P1_U2910) );
  INV_X1 U16669 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n20007) );
  AOI22_X1 U16670 ( .A1(n20761), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n19967), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13335) );
  OAI21_X1 U16671 ( .B1(n20007), .B2(n13624), .A(n13335), .ZN(P1_U2912) );
  INV_X1 U16672 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n20034) );
  AOI22_X1 U16673 ( .A1(n20761), .A2(P1_UWORD_REG_14__SCAN_IN), .B1(n19967), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n13336) );
  OAI21_X1 U16674 ( .B1(n20034), .B2(n13624), .A(n13336), .ZN(P1_U2906) );
  AOI21_X1 U16675 ( .B1(n13339), .B2(n13338), .A(n13337), .ZN(n19187) );
  AOI21_X1 U16676 ( .B1(n13342), .B2(n13341), .A(n13340), .ZN(n19172) );
  AOI22_X1 U16677 ( .A1(n19187), .A2(n11114), .B1(n16261), .B2(n19172), .ZN(
        n13343) );
  OR2_X1 U16678 ( .A1(n19155), .A2(n19704), .ZN(n19177) );
  OAI211_X1 U16679 ( .C1(n19154), .C2(n13690), .A(n13343), .B(n19177), .ZN(
        n13346) );
  INV_X1 U16680 ( .A(n13687), .ZN(n13344) );
  OAI22_X1 U16681 ( .A1(n19178), .A2(n13862), .B1(n15396), .B2(n13344), .ZN(
        n13345) );
  OR2_X1 U16682 ( .A1(n13346), .A2(n13345), .ZN(P2_U3012) );
  INV_X1 U16683 ( .A(n13347), .ZN(n13546) );
  INV_X1 U16684 ( .A(n13377), .ZN(n13375) );
  NAND2_X1 U16685 ( .A1(n13546), .A2(n13375), .ZN(n13354) );
  INV_X1 U16686 ( .A(n13354), .ZN(n13358) );
  INV_X1 U16687 ( .A(n13348), .ZN(n20553) );
  NAND2_X1 U16688 ( .A1(n13349), .A2(n13259), .ZN(n13350) );
  NOR2_X1 U16689 ( .A1(n13351), .A2(n13350), .ZN(n13353) );
  AND3_X1 U16690 ( .A1(n13353), .A2(n13352), .A3(n12321), .ZN(n13427) );
  INV_X1 U16691 ( .A(n13427), .ZN(n14558) );
  INV_X1 U16692 ( .A(n15732), .ZN(n13431) );
  OAI22_X1 U16693 ( .A1(n13431), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n13354), .B2(n11634), .ZN(n13355) );
  AOI21_X1 U16694 ( .B1(n20553), .B2(n14558), .A(n13355), .ZN(n15735) );
  INV_X1 U16695 ( .A(n16151), .ZN(n13356) );
  INV_X1 U16696 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13633) );
  INV_X1 U16697 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14537) );
  AOI22_X1 U16698 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n13633), .B2(n14537), .ZN(
        n13437) );
  NOR2_X1 U16699 ( .A1(n13902), .A2(n15018), .ZN(n13436) );
  INV_X1 U16700 ( .A(n13436), .ZN(n14560) );
  OAI22_X1 U16701 ( .A1(n15735), .A2(n13356), .B1(n13437), .B2(n14560), .ZN(
        n13357) );
  AOI21_X1 U16702 ( .B1(n14561), .B2(n13358), .A(n13357), .ZN(n13372) );
  NAND2_X1 U16703 ( .A1(n20105), .A2(n13907), .ZN(n13920) );
  OR2_X1 U16704 ( .A1(n13920), .A2(n13359), .ZN(n13360) );
  AND2_X1 U16705 ( .A1(n13361), .A2(n13360), .ZN(n13362) );
  AND2_X1 U16706 ( .A1(n13363), .A2(n13362), .ZN(n13369) );
  NOR2_X1 U16707 ( .A1(n15788), .A2(n20674), .ZN(n13366) );
  NAND2_X1 U16708 ( .A1(n13373), .A2(n13259), .ZN(n13364) );
  OR2_X1 U16709 ( .A1(n13364), .A2(n15732), .ZN(n13365) );
  OAI211_X1 U16710 ( .C1(n13367), .C2(n13366), .A(n13365), .B(n14579), .ZN(
        n13368) );
  NAND2_X1 U16711 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16159), .ZN(n13554) );
  INV_X1 U16712 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19851) );
  OAI22_X1 U16713 ( .A1(n13550), .A2(n19845), .B1(n13554), .B2(n19851), .ZN(
        n16150) );
  AOI21_X1 U16714 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20756), .A(n16150), 
        .ZN(n14564) );
  NAND2_X1 U16715 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n14564), .ZN(
        n13371) );
  OAI21_X1 U16716 ( .B1(n13372), .B2(n14564), .A(n13371), .ZN(P1_U3473) );
  NAND2_X1 U16717 ( .A1(n20735), .A2(n14558), .ZN(n13387) );
  INV_X1 U16718 ( .A(n13373), .ZN(n13374) );
  OR2_X1 U16719 ( .A1(n14578), .A2(n13374), .ZN(n13424) );
  NAND2_X1 U16720 ( .A1(n13375), .A2(n11478), .ZN(n13423) );
  XNOR2_X1 U16721 ( .A(n13423), .B(n11477), .ZN(n13376) );
  NAND2_X1 U16722 ( .A1(n13424), .A2(n13376), .ZN(n13386) );
  NAND2_X1 U16723 ( .A1(n13377), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13422) );
  NAND2_X1 U16724 ( .A1(n13422), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13378) );
  NAND2_X1 U16725 ( .A1(n13379), .A2(n13378), .ZN(n13388) );
  NAND3_X1 U16726 ( .A1(n13427), .A2(n13426), .A3(n13388), .ZN(n13385) );
  INV_X1 U16727 ( .A(n13380), .ZN(n13383) );
  NAND2_X1 U16728 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13381) );
  NAND2_X1 U16729 ( .A1(n11477), .A2(n13381), .ZN(n13382) );
  NAND3_X1 U16730 ( .A1(n15732), .A2(n13383), .A3(n13382), .ZN(n13384) );
  NAND4_X1 U16731 ( .A1(n13387), .A2(n13386), .A3(n13385), .A4(n13384), .ZN(
        n13542) );
  AOI22_X1 U16732 ( .A1(n13542), .A2(n16151), .B1(n14561), .B2(n13388), .ZN(
        n13390) );
  NAND2_X1 U16733 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n14564), .ZN(
        n13389) );
  OAI21_X1 U16734 ( .B1(n13390), .B2(n14564), .A(n13389), .ZN(P1_U3469) );
  NAND3_X1 U16735 ( .A1(n20756), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16157) );
  INV_X1 U16736 ( .A(n16157), .ZN(n13391) );
  OAI21_X1 U16737 ( .B1(n13393), .B2(n13392), .A(n13564), .ZN(n14009) );
  NAND2_X1 U16738 ( .A1(n13394), .A2(n13907), .ZN(n13399) );
  XNOR2_X1 U16739 ( .A(n13471), .B(n13470), .ZN(n13396) );
  OAI211_X1 U16740 ( .C1(n13396), .C2(n14593), .A(n13395), .B(n11620), .ZN(
        n13397) );
  INV_X1 U16741 ( .A(n13397), .ZN(n13398) );
  XOR2_X1 U16742 ( .A(n13465), .B(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n13463) );
  NOR2_X1 U16743 ( .A1(n13401), .A2(n13400), .ZN(n13402) );
  NAND2_X1 U16744 ( .A1(n13463), .A2(n20093), .ZN(n13408) );
  OR2_X1 U16745 ( .A1(n13403), .A2(n20602), .ZN(n20759) );
  AND2_X1 U16746 ( .A1(n20759), .A2(n20756), .ZN(n13404) );
  NAND2_X1 U16747 ( .A1(n20756), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15763) );
  NAND2_X1 U16748 ( .A1(n20753), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13405) );
  NAND2_X1 U16749 ( .A1(n15763), .A2(n13405), .ZN(n20090) );
  INV_X1 U16750 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14003) );
  NAND2_X1 U16751 ( .A1(n16052), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n13456) );
  OAI21_X1 U16752 ( .B1(n16026), .B2(n14003), .A(n13456), .ZN(n13406) );
  AOI21_X1 U16753 ( .B1(n16021), .B2(n14003), .A(n13406), .ZN(n13407) );
  OAI211_X1 U16754 ( .C1(n20102), .C2(n14009), .A(n13408), .B(n13407), .ZN(
        P1_U2998) );
  NAND2_X1 U16755 ( .A1(n14522), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n13410) );
  OR2_X1 U16756 ( .A1(n14525), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13412) );
  NAND2_X1 U16757 ( .A1(n13413), .A2(n13412), .ZN(n13482) );
  XNOR2_X1 U16758 ( .A(n13482), .B(n13414), .ZN(n13483) );
  INV_X1 U16759 ( .A(n14467), .ZN(n14524) );
  XNOR2_X1 U16760 ( .A(n13483), .B(n14524), .ZN(n14006) );
  OAI222_X1 U16761 ( .A1(n14009), .A2(n14750), .B1(n13409), .B2(n15945), .C1(
        n14006), .C2(n14761), .ZN(P1_U2871) );
  NOR2_X1 U16762 ( .A1(n13417), .A2(n13415), .ZN(n13416) );
  NAND2_X1 U16763 ( .A1(n20101), .A2(DATAI_1_), .ZN(n13420) );
  NAND2_X1 U16764 ( .A1(n20099), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13419) );
  AND2_X1 U16765 ( .A1(n13420), .A2(n13419), .ZN(n20121) );
  INV_X1 U16766 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20042) );
  OAI222_X1 U16767 ( .A1(n14009), .A2(n14828), .B1(n14379), .B2(n20121), .C1(
        n14815), .C2(n20042), .ZN(P1_U2903) );
  OR2_X1 U16768 ( .A1(n20491), .A2(n13427), .ZN(n13434) );
  XNOR2_X1 U16769 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13430) );
  NAND2_X1 U16770 ( .A1(n13423), .A2(n13422), .ZN(n13425) );
  NAND2_X1 U16771 ( .A1(n13424), .A2(n13425), .ZN(n13429) );
  INV_X1 U16772 ( .A(n13425), .ZN(n13435) );
  NAND3_X1 U16773 ( .A1(n13427), .A2(n13426), .A3(n13435), .ZN(n13428) );
  OAI211_X1 U16774 ( .C1(n13431), .C2(n13430), .A(n13429), .B(n13428), .ZN(
        n13432) );
  INV_X1 U16775 ( .A(n13432), .ZN(n13433) );
  NAND2_X1 U16776 ( .A1(n13434), .A2(n13433), .ZN(n13543) );
  AOI222_X1 U16777 ( .A1(n13543), .A2(n16151), .B1(n13437), .B2(n13436), .C1(
        n13435), .C2(n14561), .ZN(n13438) );
  INV_X1 U16778 ( .A(n14564), .ZN(n16155) );
  MUX2_X1 U16779 ( .A(n11478), .B(n13438), .S(n16155), .Z(n13439) );
  INV_X1 U16780 ( .A(n13439), .ZN(P1_U3472) );
  INV_X1 U16781 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n14257) );
  AOI22_X1 U16782 ( .A1(n19821), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n13440) );
  OAI21_X1 U16783 ( .B1(n14257), .B2(n13454), .A(n13440), .ZN(P2_U2930) );
  AOI22_X1 U16784 ( .A1(n19821), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .ZN(n13441) );
  OAI21_X1 U16785 ( .B1(n13442), .B2(n13454), .A(n13441), .ZN(P2_U2921) );
  INV_X1 U16786 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n15205) );
  AOI22_X1 U16787 ( .A1(n19821), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n13443) );
  OAI21_X1 U16788 ( .B1(n15205), .B2(n13454), .A(n13443), .ZN(P2_U2928) );
  INV_X1 U16789 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14340) );
  AOI22_X1 U16790 ( .A1(n19821), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n13444) );
  OAI21_X1 U16791 ( .B1(n14340), .B2(n13454), .A(n13444), .ZN(P2_U2929) );
  AOI22_X1 U16792 ( .A1(n19821), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n13445) );
  OAI21_X1 U16793 ( .B1(n15181), .B2(n13454), .A(n13445), .ZN(P2_U2924) );
  AOI22_X1 U16794 ( .A1(n19821), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n13446) );
  OAI21_X1 U16795 ( .B1(n13447), .B2(n13454), .A(n13446), .ZN(P2_U2927) );
  INV_X1 U16796 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n13449) );
  AOI22_X1 U16797 ( .A1(n19821), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n13448) );
  OAI21_X1 U16798 ( .B1(n13449), .B2(n13454), .A(n13448), .ZN(P2_U2931) );
  AOI22_X1 U16799 ( .A1(n19821), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n13450) );
  OAI21_X1 U16800 ( .B1(n11055), .B2(n13454), .A(n13450), .ZN(P2_U2935) );
  AOI22_X1 U16801 ( .A1(n19821), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n13451) );
  OAI21_X1 U16802 ( .B1(n14228), .B2(n13454), .A(n13451), .ZN(P2_U2934) );
  AOI22_X1 U16803 ( .A1(n19821), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n13452) );
  OAI21_X1 U16804 ( .B1(n14219), .B2(n13454), .A(n13452), .ZN(P2_U2932) );
  INV_X1 U16805 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n13455) );
  AOI22_X1 U16806 ( .A1(n19821), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n13453) );
  OAI21_X1 U16807 ( .B1(n13455), .B2(n13454), .A(n13453), .ZN(P2_U2933) );
  OAI21_X1 U16808 ( .B1(n16068), .B2(n14006), .A(n13456), .ZN(n13462) );
  AND2_X1 U16809 ( .A1(n15018), .A2(n15794), .ZN(n13479) );
  NOR2_X1 U16810 ( .A1(n16131), .A2(n13479), .ZN(n13460) );
  INV_X1 U16811 ( .A(n13477), .ZN(n13457) );
  AOI21_X1 U16812 ( .B1(n15018), .B2(n14547), .A(n13457), .ZN(n13458) );
  INV_X1 U16813 ( .A(n13458), .ZN(n13459) );
  MUX2_X1 U16814 ( .A(n13460), .B(n13459), .S(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(n13461) );
  AOI211_X1 U16815 ( .C1(n16144), .C2(n13463), .A(n13462), .B(n13461), .ZN(
        n13464) );
  INV_X1 U16816 ( .A(n13464), .ZN(P1_U3030) );
  INV_X1 U16817 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n13634) );
  INV_X1 U16818 ( .A(n14593), .ZN(n20754) );
  NAND2_X1 U16819 ( .A1(n13471), .A2(n13470), .ZN(n13467) );
  NAND2_X1 U16820 ( .A1(n13468), .A2(n13467), .ZN(n13630) );
  NAND3_X1 U16821 ( .A1(n13471), .A2(n13470), .A3(n13469), .ZN(n13472) );
  NAND2_X1 U16822 ( .A1(n13630), .A2(n13472), .ZN(n13475) );
  INV_X1 U16823 ( .A(n13473), .ZN(n13474) );
  AOI21_X1 U16824 ( .B1(n20754), .B2(n13475), .A(n13474), .ZN(n13476) );
  OAI21_X1 U16825 ( .B1(n20371), .B2(n13716), .A(n13476), .ZN(n13625) );
  XNOR2_X1 U16826 ( .A(n13626), .B(n13625), .ZN(n13569) );
  OR2_X1 U16827 ( .A1(n15019), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13478) );
  OAI21_X1 U16828 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n15057), .A(
        n14539), .ZN(n13481) );
  NOR2_X1 U16829 ( .A1(n15057), .A2(n13479), .ZN(n14535) );
  INV_X1 U16830 ( .A(n14535), .ZN(n16127) );
  OAI21_X1 U16831 ( .B1(n13633), .B2(n16127), .A(n13634), .ZN(n13480) );
  OAI21_X1 U16832 ( .B1(n13634), .B2(n13481), .A(n13480), .ZN(n13496) );
  AOI21_X1 U16833 ( .B1(n13483), .B2(n14467), .A(n13482), .ZN(n13487) );
  INV_X1 U16834 ( .A(n13487), .ZN(n13490) );
  MUX2_X1 U16835 ( .A(n14472), .B(n14522), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n13485) );
  OR2_X1 U16836 ( .A1(n14525), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13484) );
  NAND2_X1 U16837 ( .A1(n13485), .A2(n13484), .ZN(n13489) );
  INV_X1 U16838 ( .A(n13489), .ZN(n13486) );
  NAND2_X1 U16839 ( .A1(n13487), .A2(n13486), .ZN(n13582) );
  AOI21_X1 U16840 ( .B1(n13490), .B2(n13489), .A(n13488), .ZN(n13925) );
  AND2_X1 U16841 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n13492) );
  OAI21_X1 U16842 ( .B1(n15018), .B2(n13633), .A(n13634), .ZN(n13848) );
  INV_X1 U16843 ( .A(n13848), .ZN(n13491) );
  AOI21_X1 U16844 ( .B1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n13492), .A(
        n13491), .ZN(n13493) );
  INV_X1 U16845 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n20682) );
  OAI22_X1 U16846 ( .A1(n15055), .A2(n13493), .B1(n20682), .B2(n16103), .ZN(
        n13494) );
  AOI21_X1 U16847 ( .B1(n13925), .B2(n16142), .A(n13494), .ZN(n13495) );
  OAI211_X1 U16848 ( .C1(n16111), .C2(n13569), .A(n13496), .B(n13495), .ZN(
        P1_U3029) );
  NAND2_X1 U16849 ( .A1(n13498), .A2(n13497), .ZN(n13499) );
  NOR2_X1 U16850 ( .A1(n13500), .A2(n13501), .ZN(n13504) );
  INV_X1 U16851 ( .A(n13502), .ZN(n13503) );
  OAI211_X1 U16852 ( .C1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .C2(n13504), .A(
        n13503), .B(n15150), .ZN(n13508) );
  NAND2_X1 U16853 ( .A1(n13609), .A2(n13505), .ZN(n13506) );
  AND2_X1 U16854 ( .A1(n13588), .A2(n13506), .ZN(n16271) );
  NAND2_X1 U16855 ( .A1(n16271), .A2(n15157), .ZN(n13507) );
  OAI211_X1 U16856 ( .C1(n15157), .C2(n13509), .A(n13508), .B(n13507), .ZN(
        P2_U2881) );
  INV_X1 U16857 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n13512) );
  MUX2_X1 U16858 ( .A(n13512), .B(n13670), .S(n15157), .Z(n13513) );
  OAI21_X1 U16859 ( .B1(n19076), .B2(n15124), .A(n13513), .ZN(P2_U2884) );
  NAND2_X1 U16860 ( .A1(n20101), .A2(DATAI_0_), .ZN(n13515) );
  NAND2_X1 U16861 ( .A1(n20099), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13514) );
  AND2_X1 U16862 ( .A1(n13515), .A2(n13514), .ZN(n20112) );
  INV_X1 U16863 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20038) );
  OAI222_X1 U16864 ( .A1(n20097), .A2(n14814), .B1(n14379), .B2(n20112), .C1(
        n14815), .C2(n20038), .ZN(P1_U2904) );
  INV_X1 U16865 ( .A(n13516), .ZN(n13519) );
  INV_X1 U16866 ( .A(n13517), .ZN(n13518) );
  NAND2_X1 U16867 ( .A1(n13519), .A2(n13518), .ZN(n13520) );
  NAND2_X1 U16868 ( .A1(n13523), .A2(n13522), .ZN(n13525) );
  INV_X1 U16869 ( .A(n19777), .ZN(n13695) );
  XNOR2_X1 U16870 ( .A(n19782), .B(n13695), .ZN(n13536) );
  XNOR2_X1 U16871 ( .A(n13531), .B(n13530), .ZN(n19791) );
  INV_X1 U16872 ( .A(n19791), .ZN(n13532) );
  NAND2_X1 U16873 ( .A1(n14180), .A2(n13532), .ZN(n13533) );
  OAI21_X1 U16874 ( .B1(n14180), .B2(n13532), .A(n13533), .ZN(n19101) );
  NOR2_X1 U16875 ( .A1(n19101), .A2(n19102), .ZN(n19100) );
  INV_X1 U16876 ( .A(n13533), .ZN(n13534) );
  NOR2_X1 U16877 ( .A1(n19100), .A2(n13534), .ZN(n13535) );
  NOR2_X1 U16878 ( .A1(n13535), .A2(n13536), .ZN(n19073) );
  AOI21_X1 U16879 ( .B1(n13536), .B2(n13535), .A(n19073), .ZN(n13540) );
  INV_X1 U16880 ( .A(n13537), .ZN(n16225) );
  AOI22_X1 U16881 ( .A1(n19071), .A2(n16225), .B1(n19098), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n13539) );
  NAND2_X1 U16882 ( .A1(n13695), .A2(n19099), .ZN(n13538) );
  OAI211_X1 U16883 ( .C1(n13540), .C2(n19103), .A(n13539), .B(n13538), .ZN(
        P2_U2917) );
  MUX2_X1 U16884 ( .A(n10247), .B(n10217), .S(n15169), .Z(n13541) );
  OAI21_X1 U16885 ( .B1(n15124), .B2(n19796), .A(n13541), .ZN(P2_U2887) );
  MUX2_X1 U16886 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n13542), .S(
        n15737), .Z(n15745) );
  AND2_X1 U16887 ( .A1(n19851), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13552) );
  AOI22_X1 U16888 ( .A1(n13902), .A2(n15745), .B1(n13552), .B2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n15748) );
  MUX2_X1 U16889 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n13543), .S(
        n15737), .Z(n15741) );
  NAND2_X1 U16890 ( .A1(n15741), .A2(n13902), .ZN(n13545) );
  NAND2_X1 U16891 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n13552), .ZN(
        n13544) );
  NAND2_X1 U16892 ( .A1(n13545), .A2(n13544), .ZN(n15757) );
  NAND2_X1 U16893 ( .A1(n15757), .A2(n13546), .ZN(n13547) );
  OR2_X1 U16894 ( .A1(n15748), .A2(n13547), .ZN(n13553) );
  INV_X1 U16895 ( .A(n20259), .ZN(n20490) );
  OR2_X1 U16896 ( .A1(n11780), .A2(n20490), .ZN(n13548) );
  XNOR2_X1 U16897 ( .A(n13548), .B(n16154), .ZN(n14695) );
  NOR2_X1 U16898 ( .A1(n14695), .A2(n12321), .ZN(n16152) );
  OAI21_X1 U16899 ( .B1(n16152), .B2(n13550), .A(n13902), .ZN(n13549) );
  AOI21_X1 U16900 ( .B1(n13550), .B2(n16154), .A(n13549), .ZN(n13551) );
  AOI21_X1 U16901 ( .B1(n13552), .B2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n13551), .ZN(n15753) );
  NAND2_X1 U16902 ( .A1(n13553), .A2(n15753), .ZN(n13558) );
  INV_X1 U16903 ( .A(n13554), .ZN(n13555) );
  OAI21_X1 U16904 ( .B1(n13558), .B2(P1_FLUSH_REG_SCAN_IN), .A(n13555), .ZN(
        n13557) );
  NAND2_X1 U16905 ( .A1(n20752), .A2(n13902), .ZN(n20755) );
  INV_X1 U16906 ( .A(n20755), .ZN(n13556) );
  NAND2_X1 U16907 ( .A1(n13557), .A2(n20265), .ZN(n20736) );
  NOR2_X1 U16908 ( .A1(n13558), .A2(n16163), .ZN(n15770) );
  INV_X1 U16909 ( .A(n9621), .ZN(n13559) );
  NAND2_X1 U16910 ( .A1(n20493), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n20734) );
  INV_X1 U16911 ( .A(n20734), .ZN(n15071) );
  OAI22_X1 U16912 ( .A1(n13249), .A2(n20728), .B1(n13559), .B2(n15071), .ZN(
        n13560) );
  OAI21_X1 U16913 ( .B1(n15770), .B2(n13560), .A(n20736), .ZN(n13561) );
  OAI21_X1 U16914 ( .B1(n20736), .B2(n20519), .A(n13561), .ZN(P1_U3478) );
  INV_X1 U16915 ( .A(n13562), .ZN(n13563) );
  AOI21_X1 U16916 ( .B1(n13565), .B2(n13564), .A(n13563), .ZN(n13585) );
  AOI22_X1 U16917 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n16141), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n13566) );
  OAI21_X1 U16918 ( .B1(n16019), .B2(n13919), .A(n13566), .ZN(n13567) );
  AOI21_X1 U16919 ( .B1(n13585), .B2(n16022), .A(n13567), .ZN(n13568) );
  OAI21_X1 U16920 ( .B1(n19850), .B2(n13569), .A(n13568), .ZN(P1_U2997) );
  OR2_X1 U16921 ( .A1(n13572), .A2(n13571), .ZN(n13573) );
  NAND2_X1 U16922 ( .A1(n13570), .A2(n13573), .ZN(n19932) );
  INV_X1 U16923 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n13575) );
  NAND2_X1 U16924 ( .A1(n14466), .A2(n13575), .ZN(n13579) );
  INV_X1 U16925 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13720) );
  NAND2_X1 U16926 ( .A1(n13781), .A2(n13720), .ZN(n13577) );
  NAND2_X1 U16927 ( .A1(n14467), .A2(n13575), .ZN(n13576) );
  NAND3_X1 U16928 ( .A1(n13577), .A2(n14522), .A3(n13576), .ZN(n13578) );
  AND2_X1 U16929 ( .A1(n13579), .A2(n13578), .ZN(n13581) );
  NAND2_X1 U16930 ( .A1(n13582), .A2(n13581), .ZN(n13583) );
  AND2_X1 U16931 ( .A1(n13645), .A2(n13583), .ZN(n19930) );
  AOI22_X1 U16932 ( .A1(n15941), .A2(n19930), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n14763), .ZN(n13584) );
  OAI21_X1 U16933 ( .B1(n19932), .B2(n14750), .A(n13584), .ZN(P1_U2869) );
  INV_X1 U16934 ( .A(n13585), .ZN(n13927) );
  AOI22_X1 U16935 ( .A1(n15941), .A2(n13925), .B1(P1_EBX_REG_2__SCAN_IN), .B2(
        n14763), .ZN(n13586) );
  OAI21_X1 U16936 ( .B1(n13927), .B2(n14750), .A(n13586), .ZN(P1_U2870) );
  XNOR2_X1 U16937 ( .A(n13502), .B(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13592) );
  NAND2_X1 U16938 ( .A1(n13588), .A2(n13587), .ZN(n13589) );
  NAND2_X1 U16939 ( .A1(n13649), .A2(n13589), .ZN(n18979) );
  INV_X1 U16940 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13590) );
  MUX2_X1 U16941 ( .A(n18979), .B(n13590), .S(n15169), .Z(n13591) );
  OAI21_X1 U16942 ( .B1(n13592), .B2(n15124), .A(n13591), .ZN(P2_U2880) );
  NAND2_X1 U16943 ( .A1(n13594), .A2(n9840), .ZN(n13595) );
  OR2_X1 U16944 ( .A1(n13596), .A2(n13595), .ZN(n13597) );
  NAND2_X1 U16945 ( .A1(n13500), .A2(n13597), .ZN(n19084) );
  NOR2_X1 U16946 ( .A1(n13599), .A2(n13598), .ZN(n13600) );
  OR2_X1 U16947 ( .A1(n13607), .A2(n13600), .ZN(n19163) );
  MUX2_X1 U16948 ( .A(n10750), .B(n19163), .S(n15157), .Z(n13601) );
  OAI21_X1 U16949 ( .B1(n19084), .B2(n15124), .A(n13601), .ZN(P2_U2883) );
  INV_X1 U16950 ( .A(n19782), .ZN(n19074) );
  INV_X1 U16951 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n13602) );
  MUX2_X1 U16952 ( .A(n19178), .B(n13602), .S(n15169), .Z(n13603) );
  OAI21_X1 U16953 ( .B1(n19074), .B2(n15124), .A(n13603), .ZN(P2_U2885) );
  MUX2_X1 U16954 ( .A(n15666), .B(n13604), .S(n15169), .Z(n13605) );
  OAI21_X1 U16955 ( .B1(n14180), .B2(n15124), .A(n13605), .ZN(P2_U2886) );
  XOR2_X1 U16956 ( .A(n13500), .B(P2_INSTQUEUE_REG_0__5__SCAN_IN), .Z(n13611)
         );
  OR2_X1 U16957 ( .A1(n13607), .A2(n13606), .ZN(n13608) );
  NAND2_X1 U16958 ( .A1(n13609), .A2(n13608), .ZN(n18991) );
  MUX2_X1 U16959 ( .A(n10755), .B(n18991), .S(n15157), .Z(n13610) );
  OAI21_X1 U16960 ( .B1(n13611), .B2(n15124), .A(n13610), .ZN(P2_U2882) );
  NAND2_X1 U16961 ( .A1(n20101), .A2(DATAI_2_), .ZN(n13613) );
  NAND2_X1 U16962 ( .A1(n20099), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13612) );
  AND2_X1 U16963 ( .A1(n13613), .A2(n13612), .ZN(n20124) );
  INV_X1 U16964 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20866) );
  OAI222_X1 U16965 ( .A1(n13927), .A2(n14828), .B1(n14379), .B2(n20124), .C1(
        n20866), .C2(n14815), .ZN(P1_U2902) );
  NAND2_X1 U16966 ( .A1(n20101), .A2(DATAI_3_), .ZN(n13615) );
  NAND2_X1 U16967 ( .A1(n20099), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13614) );
  AND2_X1 U16968 ( .A1(n13615), .A2(n13614), .ZN(n20128) );
  INV_X1 U16969 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20049) );
  OAI222_X1 U16970 ( .A1(n19932), .A2(n14814), .B1(n14379), .B2(n20128), .C1(
        n14815), .C2(n20049), .ZN(P1_U2901) );
  INV_X1 U16971 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n19976) );
  AOI22_X1 U16972 ( .A1(n19968), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(n19962), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13616) );
  OAI21_X1 U16973 ( .B1(n19976), .B2(n13624), .A(n13616), .ZN(P1_U2920) );
  AOI22_X1 U16974 ( .A1(n19968), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n19962), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13617) );
  OAI21_X1 U16975 ( .B1(n14816), .B2(n13624), .A(n13617), .ZN(P1_U2919) );
  INV_X1 U16976 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n19991) );
  AOI22_X1 U16977 ( .A1(n20761), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n19962), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13618) );
  OAI21_X1 U16978 ( .B1(n19991), .B2(n13624), .A(n13618), .ZN(P1_U2916) );
  INV_X1 U16979 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n19999) );
  AOI22_X1 U16980 ( .A1(n20761), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n19962), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13619) );
  OAI21_X1 U16981 ( .B1(n19999), .B2(n13624), .A(n13619), .ZN(P1_U2914) );
  INV_X1 U16982 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n19983) );
  AOI22_X1 U16983 ( .A1(n20761), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n19962), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13620) );
  OAI21_X1 U16984 ( .B1(n19983), .B2(n13624), .A(n13620), .ZN(P1_U2918) );
  INV_X1 U16985 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n19995) );
  AOI22_X1 U16986 ( .A1(n20761), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n19962), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13621) );
  OAI21_X1 U16987 ( .B1(n19995), .B2(n13624), .A(n13621), .ZN(P1_U2915) );
  INV_X1 U16988 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n20807) );
  AOI22_X1 U16989 ( .A1(n20761), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n19962), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13622) );
  OAI21_X1 U16990 ( .B1(n20807), .B2(n13624), .A(n13622), .ZN(P1_U2913) );
  INV_X1 U16991 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n19987) );
  AOI22_X1 U16992 ( .A1(n20761), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n19962), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13623) );
  OAI21_X1 U16993 ( .B1(n19987), .B2(n13624), .A(n13623), .ZN(P1_U2917) );
  NAND2_X1 U16994 ( .A1(n13626), .A2(n13625), .ZN(n13629) );
  NAND2_X1 U16995 ( .A1(n13627), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13628) );
  NAND2_X1 U16996 ( .A1(n13630), .A2(n13631), .ZN(n13843) );
  OAI211_X1 U16997 ( .C1(n13631), .C2(n13630), .A(n13843), .B(n20754), .ZN(
        n13632) );
  OAI21_X1 U16998 ( .B1(n20730), .B2(n13716), .A(n13632), .ZN(n13709) );
  XNOR2_X1 U16999 ( .A(n13710), .B(n13709), .ZN(n13669) );
  INV_X1 U17000 ( .A(n15057), .ZN(n14542) );
  NOR2_X1 U17001 ( .A1(n13634), .A2(n13633), .ZN(n13850) );
  INV_X1 U17002 ( .A(n13850), .ZN(n14533) );
  AOI21_X1 U17003 ( .B1(n14542), .B2(n14533), .A(n15059), .ZN(n14427) );
  OAI21_X1 U17004 ( .B1(n15055), .B2(n13848), .A(n14427), .ZN(n13718) );
  OAI21_X1 U17005 ( .B1(n14533), .B2(n16127), .A(n15055), .ZN(n14429) );
  NAND2_X1 U17006 ( .A1(n13848), .A2(n14429), .ZN(n13852) );
  NAND2_X1 U17007 ( .A1(n19930), .A2(n16142), .ZN(n13635) );
  NAND2_X1 U17008 ( .A1(n16052), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n13665) );
  OAI211_X1 U17009 ( .C1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .C2(n13852), .A(
        n13635), .B(n13665), .ZN(n13636) );
  AOI21_X1 U17010 ( .B1(n13718), .B2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n13636), .ZN(n13637) );
  OAI21_X1 U17011 ( .B1(n13669), .B2(n16111), .A(n13637), .ZN(P1_U3028) );
  AND2_X1 U17012 ( .A1(n13570), .A2(n13638), .ZN(n13640) );
  OR2_X1 U17013 ( .A1(n13640), .A2(n13639), .ZN(n14701) );
  INV_X1 U17014 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13721) );
  INV_X1 U17015 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13641) );
  NAND2_X1 U17016 ( .A1(n14467), .A2(n13641), .ZN(n13642) );
  OAI211_X1 U17017 ( .C1(n14475), .C2(n13721), .A(n13642), .B(n13781), .ZN(
        n13643) );
  OAI21_X1 U17018 ( .B1(n14472), .B2(P1_EBX_REG_4__SCAN_IN), .A(n13643), .ZN(
        n13644) );
  AND2_X1 U17019 ( .A1(n13645), .A2(n13644), .ZN(n13646) );
  NOR2_X1 U17020 ( .A1(n13787), .A2(n13646), .ZN(n14698) );
  AOI22_X1 U17021 ( .A1(n15941), .A2(n14698), .B1(P1_EBX_REG_4__SCAN_IN), .B2(
        n14763), .ZN(n13647) );
  OAI21_X1 U17022 ( .B1(n14701), .B2(n14750), .A(n13647), .ZN(P1_U2868) );
  AND2_X1 U17023 ( .A1(n13649), .A2(n13648), .ZN(n13650) );
  OR2_X1 U17024 ( .A1(n13650), .A2(n13657), .ZN(n18968) );
  OAI211_X1 U17025 ( .C1(n10077), .C2(n12530), .A(n15150), .B(n13652), .ZN(
        n13654) );
  NAND2_X1 U17026 ( .A1(n15169), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13653) );
  OAI211_X1 U17027 ( .C1(n18968), .C2(n15169), .A(n13654), .B(n13653), .ZN(
        P2_U2879) );
  INV_X1 U17028 ( .A(n13655), .ZN(n13731) );
  XNOR2_X1 U17029 ( .A(n13652), .B(n13731), .ZN(n13661) );
  OR2_X1 U17030 ( .A1(n13657), .A2(n13656), .ZN(n13659) );
  NAND2_X1 U17031 ( .A1(n13659), .A2(n13658), .ZN(n15659) );
  MUX2_X1 U17032 ( .A(n15659), .B(n9877), .S(n15169), .Z(n13660) );
  OAI21_X1 U17033 ( .B1(n13661), .B2(n15124), .A(n13660), .ZN(P2_U2878) );
  NAND2_X1 U17034 ( .A1(n20101), .A2(DATAI_4_), .ZN(n13663) );
  NAND2_X1 U17035 ( .A1(n20099), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13662) );
  AND2_X1 U17036 ( .A1(n13663), .A2(n13662), .ZN(n20131) );
  INV_X1 U17037 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20053) );
  OAI222_X1 U17038 ( .A1(n14701), .A2(n14814), .B1(n14379), .B2(n20131), .C1(
        n20053), .C2(n14815), .ZN(P1_U2900) );
  INV_X1 U17039 ( .A(n19932), .ZN(n13667) );
  NAND2_X1 U17040 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13664) );
  OAI211_X1 U17041 ( .C1(n16019), .C2(n19925), .A(n13665), .B(n13664), .ZN(
        n13666) );
  AOI21_X1 U17042 ( .B1(n13667), .B2(n16022), .A(n13666), .ZN(n13668) );
  OAI21_X1 U17043 ( .B1(n13669), .B2(n19850), .A(n13668), .ZN(P1_U2996) );
  INV_X1 U17044 ( .A(n19076), .ZN(n19766) );
  NAND2_X1 U17045 ( .A1(n16289), .A2(n13962), .ZN(n13683) );
  NAND2_X1 U17046 ( .A1(n16325), .A2(n16326), .ZN(n13947) );
  NAND2_X1 U17047 ( .A1(n13947), .A2(n13953), .ZN(n13674) );
  OR2_X1 U17048 ( .A1(n10843), .A2(n13671), .ZN(n13672) );
  NAND2_X1 U17049 ( .A1(n13672), .A2(n9599), .ZN(n13952) );
  INV_X1 U17050 ( .A(n13676), .ZN(n13673) );
  NAND2_X1 U17051 ( .A1(n13967), .A2(n13673), .ZN(n13949) );
  NAND3_X1 U17052 ( .A1(n13674), .A2(n13952), .A3(n13949), .ZN(n13680) );
  INV_X1 U17053 ( .A(n13953), .ZN(n13675) );
  NAND2_X1 U17054 ( .A1(n13947), .A2(n13675), .ZN(n13678) );
  AOI21_X1 U17055 ( .B1(n13967), .B2(n13676), .A(n9598), .ZN(n13677) );
  NAND2_X1 U17056 ( .A1(n13678), .A2(n13677), .ZN(n13679) );
  MUX2_X1 U17057 ( .A(n13680), .B(n13679), .S(n16304), .Z(n13681) );
  INV_X1 U17058 ( .A(n13681), .ZN(n13682) );
  NAND2_X1 U17059 ( .A1(n13683), .A2(n13682), .ZN(n16303) );
  AOI22_X1 U17060 ( .A1(n19766), .A2(n16356), .B1(n19763), .B2(n16303), .ZN(
        n13685) );
  NAND2_X1 U17061 ( .A1(n13975), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13684) );
  OAI21_X1 U17062 ( .B1(n13685), .B2(n13975), .A(n13684), .ZN(P2_U3596) );
  NAND2_X1 U17063 ( .A1(n9838), .A2(n13831), .ZN(n13686) );
  XNOR2_X1 U17064 ( .A(n13687), .B(n13686), .ZN(n13688) );
  NAND2_X1 U17065 ( .A1(n13688), .A2(n18993), .ZN(n13697) );
  NOR2_X1 U17066 ( .A1(n18984), .A2(n13689), .ZN(n13692) );
  OAI22_X1 U17067 ( .A1(n13690), .A2(n19028), .B1(n19704), .B2(n18978), .ZN(
        n13691) );
  AOI211_X1 U17068 ( .C1(P2_EBX_REG_2__SCAN_IN), .C2(n19018), .A(n13692), .B(
        n13691), .ZN(n13693) );
  OAI21_X1 U17069 ( .B1(n19178), .B2(n19004), .A(n13693), .ZN(n13694) );
  AOI21_X1 U17070 ( .B1(n19016), .B2(n13695), .A(n13694), .ZN(n13696) );
  OAI211_X1 U17071 ( .C1(n19005), .C2(n19074), .A(n13697), .B(n13696), .ZN(
        P2_U2853) );
  OAI21_X1 U17072 ( .B1(n13700), .B2(n13699), .A(n13698), .ZN(n16293) );
  NOR2_X1 U17073 ( .A1(n19155), .A2(n13701), .ZN(n16288) );
  AOI21_X1 U17074 ( .B1(n15338), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A(
        n16288), .ZN(n13702) );
  OAI21_X1 U17075 ( .B1(n15396), .B2(n13766), .A(n13702), .ZN(n13707) );
  OAI21_X1 U17076 ( .B1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n13771), .A(
        n13703), .ZN(n13705) );
  XNOR2_X1 U17077 ( .A(n13705), .B(n13704), .ZN(n16292) );
  NOR2_X1 U17078 ( .A1(n16292), .A2(n19147), .ZN(n13706) );
  AOI211_X1 U17079 ( .C1(n19151), .C2(n16289), .A(n13707), .B(n13706), .ZN(
        n13708) );
  OAI21_X1 U17080 ( .B1(n16293), .B2(n19148), .A(n13708), .ZN(P2_U3011) );
  NAND2_X1 U17081 ( .A1(n13710), .A2(n13709), .ZN(n13713) );
  NAND2_X1 U17082 ( .A1(n13711), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13712) );
  NAND2_X1 U17083 ( .A1(n13713), .A2(n13712), .ZN(n13837) );
  XNOR2_X1 U17084 ( .A(n13843), .B(n13841), .ZN(n13714) );
  NAND2_X1 U17085 ( .A1(n13714), .A2(n20754), .ZN(n13715) );
  XNOR2_X1 U17086 ( .A(n13838), .B(n13721), .ZN(n13836) );
  XNOR2_X1 U17087 ( .A(n13837), .B(n13836), .ZN(n13745) );
  NAND2_X1 U17088 ( .A1(n16052), .A2(P1_REIP_REG_4__SCAN_IN), .ZN(n13741) );
  NAND2_X1 U17089 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n13718), .ZN(
        n13719) );
  NAND2_X1 U17090 ( .A1(n13741), .A2(n13719), .ZN(n13723) );
  NOR2_X1 U17091 ( .A1(n13721), .A2(n13720), .ZN(n14531) );
  AOI211_X1 U17092 ( .C1(n13721), .C2(n13720), .A(n14531), .B(n13852), .ZN(
        n13722) );
  AOI211_X1 U17093 ( .C1(n16142), .C2(n14698), .A(n13723), .B(n13722), .ZN(
        n13724) );
  OAI21_X1 U17094 ( .B1(n16111), .B2(n13745), .A(n13724), .ZN(P1_U3027) );
  NAND2_X1 U17095 ( .A1(n20101), .A2(DATAI_5_), .ZN(n13727) );
  NAND2_X1 U17096 ( .A1(n20099), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13726) );
  AND2_X1 U17097 ( .A1(n13727), .A2(n13726), .ZN(n20134) );
  INV_X1 U17098 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n13728) );
  OAI222_X1 U17099 ( .A1(n16020), .A2(n14814), .B1(n20134), .B2(n14379), .C1(
        n13728), .C2(n14815), .ZN(P1_U2899) );
  INV_X1 U17100 ( .A(n13729), .ZN(n13733) );
  OAI21_X1 U17101 ( .B1(n13652), .B2(n13731), .A(n13730), .ZN(n13732) );
  NAND3_X1 U17102 ( .A1(n13733), .A2(n15150), .A3(n13732), .ZN(n13738) );
  NAND2_X1 U17103 ( .A1(n13734), .A2(n13658), .ZN(n13736) );
  INV_X1 U17104 ( .A(n13746), .ZN(n13735) );
  NAND2_X1 U17105 ( .A1(n13736), .A2(n13735), .ZN(n15644) );
  INV_X1 U17106 ( .A(n15644), .ZN(n18957) );
  NAND2_X1 U17107 ( .A1(n15157), .A2(n18957), .ZN(n13737) );
  OAI211_X1 U17108 ( .C1(n15157), .C2(n13739), .A(n13738), .B(n13737), .ZN(
        P2_U2877) );
  INV_X1 U17109 ( .A(n14701), .ZN(n13743) );
  NAND2_X1 U17110 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13740) );
  OAI211_X1 U17111 ( .C1(n16019), .C2(n14691), .A(n13741), .B(n13740), .ZN(
        n13742) );
  AOI21_X1 U17112 ( .B1(n13743), .B2(n16022), .A(n13742), .ZN(n13744) );
  OAI21_X1 U17113 ( .B1(n13745), .B2(n19850), .A(n13744), .ZN(P1_U2995) );
  XNOR2_X1 U17114 ( .A(n9610), .B(n13813), .ZN(n13751) );
  OR2_X1 U17115 ( .A1(n13747), .A2(n13746), .ZN(n13748) );
  NAND2_X1 U17116 ( .A1(n13817), .A2(n13748), .ZN(n18939) );
  MUX2_X1 U17117 ( .A(n18939), .B(n13749), .S(n15169), .Z(n13750) );
  OAI21_X1 U17118 ( .B1(n13751), .B2(n15124), .A(n13750), .ZN(P2_U2876) );
  INV_X1 U17119 ( .A(n16271), .ZN(n13764) );
  NAND2_X1 U17120 ( .A1(n9838), .A2(n13752), .ZN(n13753) );
  XNOR2_X1 U17121 ( .A(n16267), .B(n13753), .ZN(n13757) );
  NAND2_X1 U17122 ( .A1(n9705), .A2(n14508), .ZN(n14507) );
  NAND2_X1 U17123 ( .A1(n14507), .A2(n13754), .ZN(n13756) );
  XNOR2_X1 U17124 ( .A(n13756), .B(n13755), .ZN(n19067) );
  AOI22_X1 U17125 ( .A1(n18993), .A2(n13757), .B1(n19016), .B2(n19067), .ZN(
        n13763) );
  OAI21_X1 U17126 ( .B1(n19710), .B2(n18978), .A(n19155), .ZN(n13758) );
  AOI21_X1 U17127 ( .B1(n18997), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n13758), .ZN(n13759) );
  OAI21_X1 U17128 ( .B1(n18984), .B2(n13760), .A(n13759), .ZN(n13761) );
  AOI21_X1 U17129 ( .B1(P2_EBX_REG_6__SCAN_IN), .B2(n19018), .A(n13761), .ZN(
        n13762) );
  OAI211_X1 U17130 ( .C1(n19004), .C2(n13764), .A(n13763), .B(n13762), .ZN(
        P2_U2849) );
  NOR2_X1 U17131 ( .A1(n11247), .A2(n13765), .ZN(n13767) );
  XNOR2_X1 U17132 ( .A(n13767), .B(n13766), .ZN(n13779) );
  NOR2_X1 U17133 ( .A1(n19076), .A2(n19005), .ZN(n13778) );
  OR2_X1 U17134 ( .A1(n13769), .A2(n13768), .ZN(n13770) );
  NAND2_X1 U17135 ( .A1(n13770), .A2(n18999), .ZN(n19075) );
  INV_X1 U17136 ( .A(n13771), .ZN(n13774) );
  NAND2_X1 U17137 ( .A1(n19018), .A2(P2_EBX_REG_3__SCAN_IN), .ZN(n13773) );
  AOI22_X1 U17138 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n18997), .B1(
        P2_REIP_REG_3__SCAN_IN), .B2(n19017), .ZN(n13772) );
  OAI211_X1 U17139 ( .C1(n18984), .C2(n13774), .A(n13773), .B(n13772), .ZN(
        n13775) );
  AOI21_X1 U17140 ( .B1(n16289), .B2(n19020), .A(n13775), .ZN(n13776) );
  OAI21_X1 U17141 ( .B1(n19075), .B2(n19001), .A(n13776), .ZN(n13777) );
  AOI211_X1 U17142 ( .C1(n13779), .C2(n18993), .A(n13778), .B(n13777), .ZN(
        n13780) );
  INV_X1 U17143 ( .A(n13780), .ZN(P2_U2852) );
  NAND2_X1 U17144 ( .A1(n14522), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13782) );
  NAND2_X1 U17145 ( .A1(n13781), .A2(n13782), .ZN(n13784) );
  INV_X1 U17146 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n13789) );
  NAND2_X1 U17147 ( .A1(n14467), .A2(n13789), .ZN(n13783) );
  NAND2_X1 U17148 ( .A1(n13784), .A2(n13783), .ZN(n13785) );
  OAI21_X1 U17149 ( .B1(n14474), .B2(P1_EBX_REG_5__SCAN_IN), .A(n13785), .ZN(
        n13786) );
  OR2_X1 U17150 ( .A1(n13787), .A2(n13786), .ZN(n13788) );
  NAND2_X1 U17151 ( .A1(n13798), .A2(n13788), .ZN(n19911) );
  OAI222_X1 U17152 ( .A1(n19911), .A2(n14761), .B1(n13789), .B2(n15945), .C1(
        n16020), .C2(n14750), .ZN(P1_U2867) );
  AND2_X1 U17153 ( .A1(n13790), .A2(n13792), .ZN(n19905) );
  INV_X1 U17154 ( .A(n19905), .ZN(n13825) );
  INV_X1 U17155 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n19896) );
  NAND2_X1 U17156 ( .A1(n14467), .A2(n19896), .ZN(n13794) );
  NAND2_X1 U17157 ( .A1(n14522), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13793) );
  NAND3_X1 U17158 ( .A1(n13794), .A2(n13781), .A3(n13793), .ZN(n13795) );
  OAI21_X1 U17159 ( .B1(n14472), .B2(P1_EBX_REG_6__SCAN_IN), .A(n13795), .ZN(
        n13799) );
  AOI21_X1 U17160 ( .B1(n13799), .B2(n13798), .A(n9888), .ZN(n19894) );
  AOI22_X1 U17161 ( .A1(n19894), .A2(n15941), .B1(P1_EBX_REG_6__SCAN_IN), .B2(
        n14763), .ZN(n13800) );
  OAI21_X1 U17162 ( .B1(n13825), .B2(n14750), .A(n13800), .ZN(P1_U2866) );
  NOR2_X1 U17163 ( .A1(n11247), .A2(n13801), .ZN(n13802) );
  XNOR2_X1 U17164 ( .A(n13802), .B(n15395), .ZN(n13805) );
  XNOR2_X1 U17165 ( .A(n16275), .B(n13803), .ZN(n19061) );
  INV_X1 U17166 ( .A(n19061), .ZN(n13804) );
  AOI22_X1 U17167 ( .A1(n18993), .A2(n13805), .B1(n19016), .B2(n13804), .ZN(
        n13812) );
  OAI21_X1 U17168 ( .B1(n19028), .B2(n13806), .A(n19155), .ZN(n13807) );
  AOI21_X1 U17169 ( .B1(n19017), .B2(P2_REIP_REG_9__SCAN_IN), .A(n13807), .ZN(
        n13808) );
  OAI21_X1 U17170 ( .B1(n19002), .B2(n9877), .A(n13808), .ZN(n13809) );
  AOI21_X1 U17171 ( .B1(n13810), .B2(n19022), .A(n13809), .ZN(n13811) );
  OAI211_X1 U17172 ( .C1(n19004), .C2(n15659), .A(n13812), .B(n13811), .ZN(
        P2_U2846) );
  INV_X1 U17173 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n13822) );
  AND2_X1 U17174 ( .A1(n9610), .A2(n13813), .ZN(n13816) );
  OAI211_X1 U17175 ( .C1(n13816), .C2(n13815), .A(n15150), .B(n13814), .ZN(
        n13821) );
  INV_X1 U17176 ( .A(n13817), .ZN(n13819) );
  OAI21_X1 U17177 ( .B1(n13819), .B2(n9982), .A(n13888), .ZN(n15617) );
  INV_X1 U17178 ( .A(n15617), .ZN(n18933) );
  NAND2_X1 U17179 ( .A1(n15157), .A2(n18933), .ZN(n13820) );
  OAI211_X1 U17180 ( .C1(n15157), .C2(n13822), .A(n13821), .B(n13820), .ZN(
        P2_U2875) );
  NAND2_X1 U17181 ( .A1(n20101), .A2(DATAI_6_), .ZN(n13824) );
  NAND2_X1 U17182 ( .A1(n20099), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13823) );
  AND2_X1 U17183 ( .A1(n13824), .A2(n13823), .ZN(n20137) );
  OAI222_X1 U17184 ( .A1(n13825), .A2(n14814), .B1(n20137), .B2(n14379), .C1(
        n14815), .C2(n11870), .ZN(P1_U2898) );
  AOI22_X1 U17185 ( .A1(P2_EBX_REG_1__SCAN_IN), .A2(n19018), .B1(n19020), .B2(
        n13963), .ZN(n13829) );
  OAI22_X1 U17186 ( .A1(n13826), .A2(n19028), .B1(n19702), .B2(n18978), .ZN(
        n13827) );
  AOI21_X1 U17187 ( .B1(n19016), .B2(n19791), .A(n13827), .ZN(n13828) );
  OAI211_X1 U17188 ( .C1(n18984), .C2(n13830), .A(n13829), .B(n13828), .ZN(
        n13834) );
  NAND2_X1 U17189 ( .A1(n18993), .A2(n11247), .ZN(n19027) );
  OAI211_X1 U17190 ( .C1(n19035), .C2(n13832), .A(n9838), .B(n13831), .ZN(
        n13957) );
  OAI22_X1 U17191 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n19027), .B1(
        n13957), .B2(n19677), .ZN(n13833) );
  AOI211_X1 U17192 ( .C1(n19029), .C2(n19787), .A(n13834), .B(n13833), .ZN(
        n13835) );
  INV_X1 U17193 ( .A(n13835), .ZN(P2_U2854) );
  NAND2_X1 U17194 ( .A1(n13837), .A2(n13836), .ZN(n13840) );
  NAND2_X1 U17195 ( .A1(n13838), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13839) );
  INV_X1 U17196 ( .A(n13841), .ZN(n13842) );
  NOR2_X1 U17197 ( .A1(n13843), .A2(n13842), .ZN(n13845) );
  NAND2_X1 U17198 ( .A1(n13845), .A2(n13844), .ZN(n14136) );
  OAI211_X1 U17199 ( .C1(n13845), .C2(n13844), .A(n14136), .B(n20754), .ZN(
        n13846) );
  NAND2_X1 U17200 ( .A1(n13847), .A2(n13846), .ZN(n14128) );
  INV_X1 U17201 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13851) );
  XNOR2_X1 U17202 ( .A(n14128), .B(n13851), .ZN(n14126) );
  XOR2_X1 U17203 ( .A(n14127), .B(n14126), .Z(n16023) );
  INV_X1 U17204 ( .A(n16023), .ZN(n13856) );
  INV_X1 U17205 ( .A(n15055), .ZN(n15061) );
  NAND3_X1 U17206 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14531), .A3(
        n13848), .ZN(n15060) );
  AOI21_X1 U17207 ( .B1(n15061), .B2(n15060), .A(n15059), .ZN(n13849) );
  OAI221_X1 U17208 ( .B1(n15057), .B2(n14531), .C1(n15057), .C2(n13850), .A(
        n13849), .ZN(n16129) );
  NOR2_X1 U17209 ( .A1(n19911), .A2(n16068), .ZN(n13854) );
  NAND2_X1 U17210 ( .A1(n13851), .A2(n14531), .ZN(n16128) );
  NAND2_X1 U17211 ( .A1(n16052), .A2(P1_REIP_REG_5__SCAN_IN), .ZN(n16024) );
  OAI21_X1 U17212 ( .B1(n16128), .B2(n13852), .A(n16024), .ZN(n13853) );
  AOI211_X1 U17213 ( .C1(n16129), .C2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n13854), .B(n13853), .ZN(n13855) );
  OAI21_X1 U17214 ( .B1(n13856), .B2(n16111), .A(n13855), .ZN(P1_U3026) );
  NAND2_X1 U17215 ( .A1(n19076), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19227) );
  OR2_X1 U17216 ( .A1(n19227), .A2(n14047), .ZN(n19772) );
  NAND2_X1 U17217 ( .A1(n19772), .A2(n19378), .ZN(n13860) );
  OR2_X1 U17218 ( .A1(n13864), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n13858) );
  INV_X1 U17219 ( .A(n19429), .ZN(n19432) );
  NOR2_X1 U17220 ( .A1(n19764), .A2(n19432), .ZN(n13857) );
  AOI21_X1 U17221 ( .B1(n13858), .B2(n13857), .A(n19565), .ZN(n13859) );
  NAND2_X1 U17222 ( .A1(n13860), .A2(n13859), .ZN(n19416) );
  INV_X1 U17223 ( .A(n19416), .ZN(n19425) );
  INV_X1 U17224 ( .A(n14047), .ZN(n14037) );
  AOI22_X1 U17225 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n14073), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n14072), .ZN(n19552) );
  AOI22_X1 U17226 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n14073), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n14072), .ZN(n19598) );
  AOI22_X1 U17227 ( .A1(n19444), .A2(n19595), .B1(n19421), .B2(n19549), .ZN(
        n13870) );
  INV_X1 U17228 ( .A(n14258), .ZN(n19072) );
  NAND2_X1 U17229 ( .A1(n19072), .A2(n19533), .ZN(n19298) );
  NAND2_X1 U17230 ( .A1(n13864), .A2(n19429), .ZN(n13865) );
  NAND2_X1 U17231 ( .A1(n13865), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n13868) );
  NAND2_X1 U17232 ( .A1(n19764), .A2(n13866), .ZN(n13867) );
  NAND2_X1 U17233 ( .A1(n13868), .A2(n13867), .ZN(n19420) );
  AOI22_X1 U17234 ( .A1(n19594), .A2(n19420), .B1(n19432), .B2(n19593), .ZN(
        n13869) );
  OAI211_X1 U17235 ( .C1(n19425), .C2(n13871), .A(n13870), .B(n13869), .ZN(
        P2_U3109) );
  INV_X1 U17236 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13874) );
  AOI22_X1 U17237 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n14073), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n14072), .ZN(n19537) );
  INV_X1 U17238 ( .A(n19537), .ZN(n19575) );
  INV_X1 U17239 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18154) );
  INV_X1 U17240 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16437) );
  OAI22_X2 U17241 ( .A1(n18154), .A2(n14057), .B1(n16437), .B2(n14058), .ZN(
        n19576) );
  AOI22_X1 U17242 ( .A1(n19444), .A2(n19575), .B1(n19421), .B2(n19576), .ZN(
        n13873) );
  NAND2_X1 U17243 ( .A1(n19036), .A2(n19533), .ZN(n19283) );
  NAND2_X1 U17244 ( .A1(n19823), .A2(n14074), .ZN(n14195) );
  AOI22_X1 U17245 ( .A1(n19420), .A2(n19574), .B1(n19432), .B2(n19573), .ZN(
        n13872) );
  OAI211_X1 U17246 ( .C1(n19425), .C2(n13874), .A(n13873), .B(n13872), .ZN(
        P2_U3104) );
  NAND2_X1 U17247 ( .A1(n13790), .A2(n13876), .ZN(n13877) );
  AND2_X1 U17248 ( .A1(n13875), .A2(n13877), .ZN(n19888) );
  INV_X1 U17249 ( .A(n19888), .ZN(n13886) );
  NAND2_X1 U17250 ( .A1(n14522), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13878) );
  NAND2_X1 U17251 ( .A1(n13781), .A2(n13878), .ZN(n13881) );
  INV_X1 U17252 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13879) );
  NAND2_X1 U17253 ( .A1(n14467), .A2(n13879), .ZN(n13880) );
  NAND2_X1 U17254 ( .A1(n13881), .A2(n13880), .ZN(n13882) );
  OAI21_X1 U17255 ( .B1(n14474), .B2(P1_EBX_REG_7__SCAN_IN), .A(n13882), .ZN(
        n13983) );
  XNOR2_X1 U17256 ( .A(n13986), .B(n13983), .ZN(n19887) );
  AOI22_X1 U17257 ( .A1(n19887), .A2(n15941), .B1(P1_EBX_REG_7__SCAN_IN), .B2(
        n14763), .ZN(n13883) );
  OAI21_X1 U17258 ( .B1(n13886), .B2(n14750), .A(n13883), .ZN(P1_U2865) );
  NAND2_X1 U17259 ( .A1(n20101), .A2(DATAI_7_), .ZN(n13885) );
  NAND2_X1 U17260 ( .A1(n20099), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13884) );
  AND2_X1 U17261 ( .A1(n13885), .A2(n13884), .ZN(n20144) );
  OAI222_X1 U17262 ( .A1(n13886), .A2(n14828), .B1(n20144), .B2(n14379), .C1(
        n14815), .C2(n11878), .ZN(P1_U2897) );
  XNOR2_X1 U17263 ( .A(n13814), .B(n13929), .ZN(n13892) );
  INV_X1 U17264 ( .A(n13932), .ZN(n13887) );
  AOI21_X1 U17265 ( .B1(n13889), .B2(n13888), .A(n13887), .ZN(n16240) );
  INV_X1 U17266 ( .A(n16240), .ZN(n18923) );
  INV_X1 U17267 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n13890) );
  MUX2_X1 U17268 ( .A(n18923), .B(n13890), .S(n15169), .Z(n13891) );
  OAI21_X1 U17269 ( .B1(n13892), .B2(n15124), .A(n13891), .ZN(P2_U2874) );
  NOR2_X1 U17270 ( .A1(n20493), .A2(n20755), .ZN(n15769) );
  INV_X1 U17271 ( .A(n15769), .ZN(n13893) );
  NOR2_X1 U17272 ( .A1(n13893), .A2(n20756), .ZN(n13898) );
  AND2_X1 U17273 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20756), .ZN(n13894) );
  AND2_X1 U17274 ( .A1(n13895), .A2(n13894), .ZN(n13896) );
  NAND2_X1 U17275 ( .A1(n13899), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13901) );
  INV_X1 U17276 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n13900) );
  XNOR2_X1 U17277 ( .A(n13901), .B(n13900), .ZN(n14422) );
  NOR2_X1 U17278 ( .A1(n14422), .A2(n13902), .ZN(n13903) );
  INV_X1 U17279 ( .A(n13906), .ZN(n13922) );
  NAND2_X1 U17280 ( .A1(n13922), .A2(n13904), .ZN(n13905) );
  NOR2_X1 U17281 ( .A1(n13906), .A2(n20105), .ZN(n13915) );
  NAND2_X1 U17282 ( .A1(n13907), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13912) );
  AND2_X1 U17283 ( .A1(n20760), .A2(n20753), .ZN(n13908) );
  NOR2_X1 U17284 ( .A1(n13912), .A2(n13908), .ZN(n13909) );
  AND2_X1 U17285 ( .A1(n14422), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13910) );
  OR2_X1 U17286 ( .A1(n13911), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13914) );
  AND2_X1 U17287 ( .A1(n13914), .A2(n13912), .ZN(n13913) );
  NAND2_X1 U17288 ( .A1(n19938), .A2(P1_EBX_REG_2__SCAN_IN), .ZN(n13918) );
  INV_X1 U17289 ( .A(n13914), .ZN(n15761) );
  NAND2_X1 U17290 ( .A1(n19881), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n19929) );
  INV_X1 U17291 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20740) );
  AOI21_X1 U17292 ( .B1(n19881), .B2(n20740), .A(n15918), .ZN(n19937) );
  OAI22_X1 U17293 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n19929), .B1(n20682), 
        .B2(n19937), .ZN(n13916) );
  AOI21_X1 U17294 ( .B1(n19926), .B2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n13916), .ZN(n13917) );
  OAI211_X1 U17295 ( .C1(n19940), .C2(n13919), .A(n13918), .B(n13917), .ZN(
        n13924) );
  INV_X1 U17296 ( .A(n13920), .ZN(n13921) );
  NAND2_X1 U17297 ( .A1(n13922), .A2(n13921), .ZN(n14694) );
  NOR2_X1 U17298 ( .A1(n20491), .A2(n14694), .ZN(n13923) );
  AOI211_X1 U17299 ( .C1(n13925), .C2(n19945), .A(n13924), .B(n13923), .ZN(
        n13926) );
  OAI21_X1 U17300 ( .B1(n13927), .B2(n19949), .A(n13926), .ZN(P1_U2838) );
  OAI21_X1 U17301 ( .B1(n13814), .B2(n13929), .A(n13928), .ZN(n13931) );
  NAND3_X1 U17302 ( .A1(n13931), .A2(n15150), .A3(n13930), .ZN(n13935) );
  AOI21_X1 U17303 ( .B1(n13933), .B2(n13932), .A(n14031), .ZN(n18914) );
  NAND2_X1 U17304 ( .A1(n15157), .A2(n18914), .ZN(n13934) );
  OAI211_X1 U17305 ( .C1(n15157), .C2(n13936), .A(n13935), .B(n13934), .ZN(
        P2_U2873) );
  AOI221_X1 U17306 ( .B1(n19035), .B2(n9838), .C1(n13938), .C2(n11247), .A(
        n13937), .ZN(n13972) );
  INV_X1 U17307 ( .A(n13972), .ZN(n13943) );
  NAND2_X1 U17308 ( .A1(n13939), .A2(n11082), .ZN(n13966) );
  MUX2_X1 U17309 ( .A(n13966), .B(n13967), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n13940) );
  AOI21_X1 U17310 ( .B1(n19019), .B2(n13962), .A(n13940), .ZN(n16308) );
  OAI21_X1 U17311 ( .B1(n16308), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n13937), 
        .ZN(n13942) );
  AOI22_X1 U17312 ( .A1(n13943), .A2(n13942), .B1(n13941), .B2(n16356), .ZN(
        n13945) );
  NAND2_X1 U17313 ( .A1(n13975), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13944) );
  OAI21_X1 U17314 ( .B1(n13945), .B2(n13975), .A(n13944), .ZN(P2_U3601) );
  INV_X1 U17315 ( .A(n13962), .ZN(n13946) );
  OR2_X1 U17316 ( .A1(n19178), .A2(n13946), .ZN(n13956) );
  OAI21_X1 U17317 ( .B1(n12677), .B2(n13953), .A(n13947), .ZN(n13951) );
  OR2_X1 U17318 ( .A1(n13949), .A2(n13948), .ZN(n13950) );
  OAI211_X1 U17319 ( .C1(n13953), .C2(n13952), .A(n13951), .B(n13950), .ZN(
        n13954) );
  INV_X1 U17320 ( .A(n13954), .ZN(n13955) );
  NAND2_X1 U17321 ( .A1(n13956), .A2(n13955), .ZN(n16314) );
  OAI21_X1 U17322 ( .B1(n9838), .B2(n13958), .A(n13957), .ZN(n13971) );
  AOI222_X1 U17323 ( .A1(n16314), .A2(n19763), .B1(n13972), .B2(n13971), .C1(
        n16356), .C2(n19782), .ZN(n13961) );
  NAND2_X1 U17324 ( .A1(n13975), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13960) );
  OAI21_X1 U17325 ( .B1(n13961), .B2(n13975), .A(n13960), .ZN(P2_U3599) );
  NAND2_X1 U17326 ( .A1(n13963), .A2(n13962), .ZN(n13970) );
  AOI22_X1 U17327 ( .A1(n13968), .A2(n13967), .B1(n13966), .B2(n13965), .ZN(
        n13969) );
  NAND2_X1 U17328 ( .A1(n13970), .A2(n13969), .ZN(n16311) );
  INV_X1 U17329 ( .A(n13971), .ZN(n13973) );
  AOI222_X1 U17330 ( .A1(n19763), .A2(n16311), .B1(n13973), .B2(n13972), .C1(
        n19787), .C2(n16356), .ZN(n13976) );
  NAND2_X1 U17331 ( .A1(n13975), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13974) );
  OAI21_X1 U17332 ( .B1(n13976), .B2(n13975), .A(n13974), .ZN(P2_U3600) );
  NAND2_X1 U17333 ( .A1(n13875), .A2(n13977), .ZN(n13978) );
  NAND2_X1 U17334 ( .A1(n14093), .A2(n13978), .ZN(n14159) );
  INV_X1 U17335 ( .A(n14472), .ZN(n14366) );
  INV_X1 U17336 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n20808) );
  NAND2_X1 U17337 ( .A1(n14366), .A2(n20808), .ZN(n13982) );
  INV_X1 U17338 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n13980) );
  NAND2_X1 U17339 ( .A1(n14467), .A2(n20808), .ZN(n13979) );
  OAI211_X1 U17340 ( .C1(n14475), .C2(n13980), .A(n13979), .B(n13781), .ZN(
        n13981) );
  AOI21_X1 U17341 ( .B1(n9888), .B2(n13983), .A(n13984), .ZN(n13987) );
  NAND2_X1 U17342 ( .A1(n13984), .A2(n13983), .ZN(n13985) );
  OR2_X1 U17343 ( .A1(n13987), .A2(n14124), .ZN(n13990) );
  OAI22_X1 U17344 ( .A1(n13990), .A2(n14761), .B1(n20808), .B2(n15945), .ZN(
        n13988) );
  INV_X1 U17345 ( .A(n13988), .ZN(n13989) );
  OAI21_X1 U17346 ( .B1(n14159), .B2(n14750), .A(n13989), .ZN(P1_U2864) );
  INV_X1 U17347 ( .A(n14155), .ZN(n13999) );
  INV_X1 U17348 ( .A(n13990), .ZN(n16126) );
  AOI22_X1 U17349 ( .A1(n19945), .A2(n16126), .B1(n19938), .B2(
        P1_EBX_REG_8__SCAN_IN), .ZN(n13991) );
  OAI211_X1 U17350 ( .C1(n19941), .C2(n13992), .A(n13991), .B(n15929), .ZN(
        n13998) );
  NAND3_X1 U17351 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(P1_REIP_REG_6__SCAN_IN), 
        .A3(P1_REIP_REG_5__SCAN_IN), .ZN(n13994) );
  NAND3_X1 U17352 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n13993) );
  NOR2_X1 U17353 ( .A1(n15911), .A2(n13993), .ZN(n14697) );
  NAND2_X1 U17354 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(n14697), .ZN(n19924) );
  NOR2_X1 U17355 ( .A1(n13994), .A2(n19924), .ZN(n13996) );
  NAND4_X1 U17356 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(P1_REIP_REG_6__SCAN_IN), .A4(P1_REIP_REG_5__SCAN_IN), .ZN(n19869)
         );
  INV_X1 U17357 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20683) );
  INV_X1 U17358 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20684) );
  NOR4_X1 U17359 ( .A1(n20683), .A2(n20740), .A3(n20684), .A4(n20682), .ZN(
        n14346) );
  OAI21_X1 U17360 ( .B1(n15911), .B2(n14346), .A(n15837), .ZN(n19919) );
  AOI21_X1 U17361 ( .B1(n19881), .B2(n19869), .A(n19919), .ZN(n19880) );
  INV_X1 U17362 ( .A(n19880), .ZN(n13995) );
  MUX2_X1 U17363 ( .A(n13996), .B(n13995), .S(P1_REIP_REG_8__SCAN_IN), .Z(
        n13997) );
  AOI211_X1 U17364 ( .C1(n19927), .C2(n13999), .A(n13998), .B(n13997), .ZN(
        n14000) );
  OAI21_X1 U17365 ( .B1(n15891), .B2(n14159), .A(n14000), .ZN(P1_U2832) );
  INV_X1 U17366 ( .A(n14694), .ZN(n19943) );
  NAND2_X1 U17367 ( .A1(n19938), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n14002) );
  AOI22_X1 U17368 ( .A1(n19927), .A2(n14003), .B1(n15918), .B2(
        P1_REIP_REG_1__SCAN_IN), .ZN(n14001) );
  OAI211_X1 U17369 ( .C1(n19941), .C2(n14003), .A(n14002), .B(n14001), .ZN(
        n14004) );
  AOI21_X1 U17370 ( .B1(n19881), .B2(n20740), .A(n14004), .ZN(n14005) );
  OAI21_X1 U17371 ( .B1(n19897), .B2(n14006), .A(n14005), .ZN(n14007) );
  AOI21_X1 U17372 ( .B1(n20553), .B2(n19943), .A(n14007), .ZN(n14008) );
  OAI21_X1 U17373 ( .B1(n14009), .B2(n19949), .A(n14008), .ZN(P1_U2839) );
  NAND2_X1 U17374 ( .A1(n19784), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19489) );
  NOR2_X1 U17375 ( .A1(n19489), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n14017) );
  INV_X1 U17376 ( .A(n14017), .ZN(n19426) );
  OR2_X1 U17377 ( .A1(n19076), .A2(n19382), .ZN(n19563) );
  OAI21_X1 U17378 ( .B1(n19563), .B2(n19193), .A(n19764), .ZN(n14018) );
  NOR2_X1 U17379 ( .A1(n19426), .A2(n14018), .ZN(n14012) );
  INV_X1 U17380 ( .A(n14019), .ZN(n14010) );
  NOR2_X1 U17381 ( .A1(n19223), .A2(n19489), .ZN(n19463) );
  INV_X1 U17382 ( .A(n19463), .ZN(n15682) );
  AOI21_X1 U17383 ( .B1(n14010), .B2(n15682), .A(n19528), .ZN(n14011) );
  NOR2_X2 U17384 ( .A1(n19097), .A2(n19565), .ZN(n19650) );
  INV_X1 U17385 ( .A(n19650), .ZN(n19292) );
  INV_X1 U17386 ( .A(n19523), .ZN(n14013) );
  AOI22_X1 U17387 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n14072), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n14073), .ZN(n19589) );
  AOI22_X1 U17388 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n14073), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n14072), .ZN(n19546) );
  NOR2_X2 U17389 ( .A1(n19488), .A2(n19193), .ZN(n19483) );
  INV_X1 U17390 ( .A(n19483), .ZN(n14015) );
  NAND2_X1 U17391 ( .A1(n14014), .A2(n14074), .ZN(n19207) );
  OAI22_X1 U17392 ( .A1(n19546), .A2(n14015), .B1(n15682), .B2(n19207), .ZN(
        n14016) );
  AOI21_X1 U17393 ( .B1(n19453), .B2(n19651), .A(n14016), .ZN(n14025) );
  OR2_X1 U17394 ( .A1(n14018), .A2(n14017), .ZN(n14023) );
  NAND2_X1 U17395 ( .A1(n14019), .A2(n19794), .ZN(n14021) );
  NOR2_X1 U17396 ( .A1(n19764), .A2(n19463), .ZN(n14020) );
  AOI21_X1 U17397 ( .B1(n14021), .B2(n14020), .A(n19565), .ZN(n14022) );
  NAND2_X1 U17398 ( .A1(n14023), .A2(n14022), .ZN(n15684) );
  NAND2_X1 U17399 ( .A1(n15684), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n14024) );
  OAI211_X1 U17400 ( .C1(n15676), .C2(n19292), .A(n14025), .B(n14024), .ZN(
        P2_U3123) );
  NAND2_X1 U17401 ( .A1(n20101), .A2(DATAI_8_), .ZN(n14027) );
  NAND2_X1 U17402 ( .A1(n20099), .A2(BUF1_REG_8__SCAN_IN), .ZN(n14026) );
  AND2_X1 U17403 ( .A1(n14027), .A2(n14026), .ZN(n20003) );
  INV_X1 U17404 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n14028) );
  OAI222_X1 U17405 ( .A1(n14159), .A2(n14814), .B1(n20003), .B2(n14379), .C1(
        n14028), .C2(n14815), .ZN(P1_U2896) );
  XNOR2_X1 U17406 ( .A(n13930), .B(n14029), .ZN(n14036) );
  OR2_X1 U17407 ( .A1(n14031), .A2(n14030), .ZN(n14033) );
  AND2_X1 U17408 ( .A1(n14033), .A2(n14032), .ZN(n16234) );
  NOR2_X1 U17409 ( .A1(n15157), .A2(n10790), .ZN(n14034) );
  AOI21_X1 U17410 ( .B1(n16234), .B2(n15157), .A(n14034), .ZN(n14035) );
  OAI21_X1 U17411 ( .B1(n14036), .B2(n15124), .A(n14035), .ZN(P2_U2872) );
  INV_X1 U17412 ( .A(n19563), .ZN(n19495) );
  NAND2_X1 U17413 ( .A1(n19495), .A2(n14037), .ZN(n14042) );
  NAND3_X1 U17414 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n14101) );
  NOR2_X1 U17415 ( .A1(n14038), .A2(n19775), .ZN(n19662) );
  OR2_X1 U17416 ( .A1(n19662), .A2(n19528), .ZN(n14039) );
  OAI21_X1 U17417 ( .B1(n19662), .B2(n19794), .A(n19533), .ZN(n14041) );
  AOI211_X2 U17418 ( .C1(n14042), .C2(n14101), .A(n14045), .B(n14041), .ZN(
        n19672) );
  INV_X1 U17419 ( .A(n14101), .ZN(n14043) );
  AOI21_X1 U17420 ( .B1(n19794), .B2(n14043), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14044) );
  NOR2_X2 U17421 ( .A1(n19065), .A2(n19565), .ZN(n19632) );
  NAND2_X1 U17422 ( .A1(n14046), .A2(n14074), .ZN(n19216) );
  INV_X1 U17423 ( .A(n19662), .ZN(n14082) );
  AOI22_X1 U17424 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n14073), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n14072), .ZN(n19561) );
  NOR2_X2 U17425 ( .A1(n19523), .A2(n14047), .ZN(n19667) );
  INV_X1 U17426 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n16506) );
  OAI22_X2 U17427 ( .A1(n16425), .A2(n14058), .B1(n16506), .B2(n14057), .ZN(
        n19629) );
  AOI22_X1 U17428 ( .A1(n19669), .A2(n19630), .B1(n19667), .B2(n19629), .ZN(
        n14048) );
  OAI21_X1 U17429 ( .B1(n19216), .B2(n14082), .A(n14048), .ZN(n14049) );
  AOI21_X1 U17430 ( .B1(n19665), .B2(n19632), .A(n14049), .ZN(n14050) );
  OAI21_X1 U17431 ( .B1(n19672), .B2(n14051), .A(n14050), .ZN(P2_U3175) );
  INV_X1 U17432 ( .A(n19593), .ZN(n14053) );
  AOI22_X1 U17433 ( .A1(n19669), .A2(n19595), .B1(n19667), .B2(n19549), .ZN(
        n14052) );
  OAI21_X1 U17434 ( .B1(n14053), .B2(n14082), .A(n14052), .ZN(n14054) );
  AOI21_X1 U17435 ( .B1(n19665), .B2(n19594), .A(n14054), .ZN(n14055) );
  OAI21_X1 U17436 ( .B1(n19672), .B2(n14056), .A(n14055), .ZN(P2_U3173) );
  INV_X1 U17437 ( .A(n19090), .ZN(n16219) );
  NAND2_X1 U17438 ( .A1(n16219), .A2(n19533), .ZN(n19295) );
  INV_X1 U17439 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16431) );
  INV_X1 U17440 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n18176) );
  OAI22_X2 U17441 ( .A1(n16431), .A2(n14058), .B1(n18176), .B2(n14057), .ZN(
        n19658) );
  INV_X1 U17442 ( .A(n19658), .ZN(n14061) );
  AOI22_X1 U17443 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n14073), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n14072), .ZN(n19592) );
  INV_X1 U17444 ( .A(n19592), .ZN(n19657) );
  NOR2_X2 U17445 ( .A1(n14059), .A2(n14068), .ZN(n19655) );
  AOI22_X1 U17446 ( .A1(n19657), .A2(n19483), .B1(n19463), .B2(n19655), .ZN(
        n14060) );
  OAI21_X1 U17447 ( .B1(n14061), .B2(n19447), .A(n14060), .ZN(n14062) );
  AOI21_X1 U17448 ( .B1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B2(n15684), .A(
        n14062), .ZN(n14063) );
  OAI21_X1 U17449 ( .B1(n15676), .B2(n19295), .A(n14063), .ZN(P2_U3124) );
  NOR2_X2 U17450 ( .A1(n19108), .A2(n19565), .ZN(n19637) );
  INV_X1 U17451 ( .A(n19637), .ZN(n19286) );
  AOI22_X1 U17452 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n14073), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n14072), .ZN(n19583) );
  AOI22_X1 U17453 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n14073), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n14072), .ZN(n19540) );
  AOI22_X1 U17454 ( .A1(n19639), .A2(n19483), .B1(n19463), .B2(n14064), .ZN(
        n14065) );
  OAI21_X1 U17455 ( .B1(n19447), .B2(n19583), .A(n14065), .ZN(n14066) );
  AOI21_X1 U17456 ( .B1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n15684), .A(
        n14066), .ZN(n14067) );
  OAI21_X1 U17457 ( .B1(n15676), .B2(n19286), .A(n14067), .ZN(P2_U3121) );
  NAND2_X1 U17458 ( .A1(n16225), .A2(n19533), .ZN(n19289) );
  AOI22_X1 U17459 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n14073), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n14072), .ZN(n19586) );
  AOI22_X1 U17460 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n14073), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n14072), .ZN(n19543) );
  NOR2_X2 U17461 ( .A1(n10184), .A2(n14068), .ZN(n19643) );
  AOI22_X1 U17462 ( .A1(n19646), .A2(n19483), .B1(n19463), .B2(n19643), .ZN(
        n14069) );
  OAI21_X1 U17463 ( .B1(n19447), .B2(n19586), .A(n14069), .ZN(n14070) );
  AOI21_X1 U17464 ( .B1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B2(n15684), .A(
        n14070), .ZN(n14071) );
  OAI21_X1 U17465 ( .B1(n15676), .B2(n19289), .A(n14071), .ZN(P2_U3122) );
  NOR2_X2 U17466 ( .A1(n19068), .A2(n19565), .ZN(n19664) );
  INV_X1 U17467 ( .A(n19664), .ZN(n19301) );
  AOI22_X1 U17468 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n14073), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n14072), .ZN(n19516) );
  AOI22_X1 U17469 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n14073), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n14072), .ZN(n19603) );
  NAND2_X1 U17470 ( .A1(n10185), .A2(n14074), .ZN(n14189) );
  AOI22_X1 U17471 ( .A1(n19668), .A2(n19483), .B1(n19663), .B2(n19463), .ZN(
        n14075) );
  OAI21_X1 U17472 ( .B1(n19447), .B2(n19516), .A(n14075), .ZN(n14076) );
  AOI21_X1 U17473 ( .B1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B2(n15684), .A(
        n14076), .ZN(n14077) );
  OAI21_X1 U17474 ( .B1(n15676), .B2(n19301), .A(n14077), .ZN(P2_U3126) );
  AOI22_X1 U17475 ( .A1(n19595), .A2(n19483), .B1(n19463), .B2(n19593), .ZN(
        n14078) );
  OAI21_X1 U17476 ( .B1(n19598), .B2(n19447), .A(n14078), .ZN(n14079) );
  AOI21_X1 U17477 ( .B1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B2(n15684), .A(
        n14079), .ZN(n14080) );
  OAI21_X1 U17478 ( .B1(n15676), .B2(n19298), .A(n14080), .ZN(P2_U3125) );
  AOI22_X1 U17479 ( .A1(n19667), .A2(n19576), .B1(n19669), .B2(n19575), .ZN(
        n14081) );
  OAI21_X1 U17480 ( .B1(n14195), .B2(n14082), .A(n14081), .ZN(n14083) );
  AOI21_X1 U17481 ( .B1(n19665), .B2(n19574), .A(n14083), .ZN(n14084) );
  OAI21_X1 U17482 ( .B1(n19672), .B2(n14085), .A(n14084), .ZN(P2_U3168) );
  NOR2_X1 U17483 ( .A1(n9633), .A2(n14086), .ZN(n14087) );
  OR2_X1 U17484 ( .A1(n14252), .A2(n14087), .ZN(n19040) );
  NAND2_X1 U17485 ( .A1(n14032), .A2(n14089), .ZN(n14090) );
  NAND2_X1 U17486 ( .A1(n14088), .A2(n14090), .ZN(n18903) );
  MUX2_X1 U17487 ( .A(n18903), .B(n9872), .S(n15169), .Z(n14091) );
  OAI21_X1 U17488 ( .B1(n19040), .B2(n15124), .A(n14091), .ZN(P2_U2871) );
  AND2_X1 U17489 ( .A1(n14093), .A2(n14092), .ZN(n14096) );
  OR2_X1 U17490 ( .A1(n14096), .A2(n14095), .ZN(n19868) );
  INV_X1 U17491 ( .A(DATAI_9_), .ZN(n14098) );
  NAND2_X1 U17492 ( .A1(n20099), .A2(BUF1_REG_9__SCAN_IN), .ZN(n14097) );
  OAI21_X1 U17493 ( .B1(n20099), .B2(n14098), .A(n14097), .ZN(n20008) );
  AOI22_X1 U17494 ( .A1(n14826), .A2(n20008), .B1(P1_EAX_REG_9__SCAN_IN), .B2(
        n15946), .ZN(n14099) );
  OAI21_X1 U17495 ( .B1(n19868), .B2(n14828), .A(n14099), .ZN(P1_U2895) );
  NOR2_X2 U17496 ( .A1(n19488), .A2(n19562), .ZN(n19628) );
  OAI21_X1 U17497 ( .B1(n19628), .B2(n19667), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n14100) );
  NAND2_X1 U17498 ( .A1(n14100), .A2(n19764), .ZN(n14104) );
  NOR2_X1 U17499 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n14101), .ZN(
        n19626) );
  NAND3_X1 U17500 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19793), .ZN(n19572) );
  NOR2_X1 U17501 ( .A1(n19802), .A2(n19572), .ZN(n19604) );
  NOR2_X1 U17502 ( .A1(n19626), .A2(n19604), .ZN(n14108) );
  OAI21_X1 U17503 ( .B1(n14102), .B2(n19626), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14103) );
  INV_X1 U17504 ( .A(n19631), .ZN(n14118) );
  INV_X1 U17505 ( .A(n14104), .ZN(n14109) );
  AOI21_X1 U17506 ( .B1(n14105), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n14106) );
  OAI21_X1 U17507 ( .B1(n14106), .B2(n19626), .A(n19533), .ZN(n14107) );
  INV_X1 U17508 ( .A(n19636), .ZN(n14116) );
  INV_X1 U17509 ( .A(n19576), .ZN(n14111) );
  INV_X1 U17510 ( .A(n19628), .ZN(n19602) );
  AOI22_X1 U17511 ( .A1(n19575), .A2(n19667), .B1(n19573), .B2(n19626), .ZN(
        n14110) );
  OAI21_X1 U17512 ( .B1(n14111), .B2(n19602), .A(n14110), .ZN(n14112) );
  AOI21_X1 U17513 ( .B1(n14116), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A(
        n14112), .ZN(n14113) );
  OAI21_X1 U17514 ( .B1(n19283), .B2(n14118), .A(n14113), .ZN(P2_U3160) );
  AOI22_X1 U17515 ( .A1(n19595), .A2(n19667), .B1(n19593), .B2(n19626), .ZN(
        n14114) );
  OAI21_X1 U17516 ( .B1(n19598), .B2(n19602), .A(n14114), .ZN(n14115) );
  AOI21_X1 U17517 ( .B1(n14116), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A(
        n14115), .ZN(n14117) );
  OAI21_X1 U17518 ( .B1(n19298), .B2(n14118), .A(n14117), .ZN(P2_U3165) );
  INV_X1 U17519 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n14125) );
  NAND2_X1 U17520 ( .A1(n14522), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14119) );
  NAND2_X1 U17521 ( .A1(n13781), .A2(n14119), .ZN(n14121) );
  NAND2_X1 U17522 ( .A1(n14467), .A2(n14125), .ZN(n14120) );
  NAND2_X1 U17523 ( .A1(n14121), .A2(n14120), .ZN(n14122) );
  OAI21_X1 U17524 ( .B1(n14474), .B2(P1_EBX_REG_9__SCAN_IN), .A(n14122), .ZN(
        n14123) );
  OAI21_X1 U17525 ( .B1(n14124), .B2(n14123), .A(n14166), .ZN(n19874) );
  OAI222_X1 U17526 ( .A1(n19868), .A2(n14750), .B1(n14125), .B2(n15945), .C1(
        n19874), .C2(n14761), .ZN(P1_U2863) );
  NAND2_X1 U17527 ( .A1(n14128), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n14129) );
  NAND3_X1 U17528 ( .A1(n14149), .A2(n14130), .A3(n14145), .ZN(n14133) );
  XNOR2_X1 U17529 ( .A(n14136), .B(n14137), .ZN(n14131) );
  NAND2_X1 U17530 ( .A1(n14131), .A2(n20754), .ZN(n14132) );
  NAND2_X1 U17531 ( .A1(n14133), .A2(n14132), .ZN(n14134) );
  NAND2_X1 U17532 ( .A1(n14134), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16013) );
  NAND2_X1 U17533 ( .A1(n14135), .A2(n14145), .ZN(n14141) );
  INV_X1 U17534 ( .A(n14136), .ZN(n14138) );
  NAND2_X1 U17535 ( .A1(n14138), .A2(n14137), .ZN(n14150) );
  XNOR2_X1 U17536 ( .A(n14150), .B(n14151), .ZN(n14139) );
  NAND2_X1 U17537 ( .A1(n14139), .A2(n20754), .ZN(n14140) );
  NAND2_X1 U17538 ( .A1(n14141), .A2(n14140), .ZN(n14143) );
  XNOR2_X1 U17539 ( .A(n14143), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16007) );
  OR2_X1 U17540 ( .A1(n14143), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14144) );
  NAND2_X1 U17541 ( .A1(n14145), .A2(n14151), .ZN(n14147) );
  NOR2_X1 U17542 ( .A1(n14147), .A2(n14146), .ZN(n14148) );
  INV_X1 U17543 ( .A(n14150), .ZN(n14152) );
  NAND3_X1 U17544 ( .A1(n14152), .A2(n20754), .A3(n14151), .ZN(n14153) );
  NAND2_X1 U17545 ( .A1(n9626), .A2(n14153), .ZN(n14395) );
  XOR2_X1 U17546 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n14395), .Z(
        n14154) );
  XNOR2_X1 U17547 ( .A(n14394), .B(n14154), .ZN(n16132) );
  NAND2_X1 U17548 ( .A1(n16132), .A2(n20093), .ZN(n14158) );
  AND2_X1 U17549 ( .A1(n16141), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n16125) );
  NOR2_X1 U17550 ( .A1(n16019), .A2(n14155), .ZN(n14156) );
  AOI211_X1 U17551 ( .C1(n20091), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16125), .B(n14156), .ZN(n14157) );
  OAI211_X1 U17552 ( .C1(n20102), .C2(n14159), .A(n14158), .B(n14157), .ZN(
        P1_U2991) );
  INV_X1 U17553 ( .A(n14160), .ZN(n14163) );
  INV_X1 U17554 ( .A(n14095), .ZN(n14162) );
  INV_X1 U17555 ( .A(n14161), .ZN(n14678) );
  AOI21_X1 U17556 ( .B1(n14163), .B2(n14162), .A(n14678), .ZN(n15933) );
  INV_X1 U17557 ( .A(n15933), .ZN(n14960) );
  MUX2_X1 U17558 ( .A(n14472), .B(n14522), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n14164) );
  OAI21_X1 U17559 ( .B1(n14525), .B2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n14164), .ZN(n14167) );
  INV_X1 U17560 ( .A(n14317), .ZN(n14165) );
  AOI21_X1 U17561 ( .B1(n14167), .B2(n14166), .A(n14165), .ZN(n16115) );
  AOI22_X1 U17562 ( .A1(n16115), .A2(n15941), .B1(P1_EBX_REG_10__SCAN_IN), 
        .B2(n14763), .ZN(n14168) );
  OAI21_X1 U17563 ( .B1(n14960), .B2(n14750), .A(n14168), .ZN(P1_U2862) );
  XNOR2_X1 U17564 ( .A(n14169), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n16269) );
  XNOR2_X1 U17565 ( .A(n14171), .B(n14170), .ZN(n16268) );
  AOI22_X1 U17566 ( .A1(n19067), .A2(n16296), .B1(n16290), .B2(n16271), .ZN(
        n14177) );
  NAND2_X1 U17567 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n18902), .ZN(n14172) );
  OAI221_X1 U17568 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n14174), .C1(
        n14173), .C2(n14268), .A(n14172), .ZN(n14175) );
  INV_X1 U17569 ( .A(n14175), .ZN(n14176) );
  OAI211_X1 U17570 ( .C1(n16268), .C2(n19157), .A(n14177), .B(n14176), .ZN(
        n14178) );
  INV_X1 U17571 ( .A(n14178), .ZN(n14179) );
  OAI21_X1 U17572 ( .B1(n16269), .B2(n19174), .A(n14179), .ZN(P2_U3040) );
  NOR2_X2 U17573 ( .A1(n19487), .A2(n19312), .ZN(n19303) );
  NAND2_X1 U17574 ( .A1(n19775), .A2(n19784), .ZN(n19271) );
  NOR2_X1 U17575 ( .A1(n19462), .A2(n19271), .ZN(n14181) );
  AOI221_X1 U17576 ( .B1(n19267), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19303), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n14181), .ZN(n14184) );
  AOI21_X1 U17577 ( .B1(n14185), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n14182) );
  NOR2_X1 U17578 ( .A1(n19459), .A2(n19271), .ZN(n19265) );
  OAI21_X1 U17579 ( .B1(n14182), .B2(n19265), .A(n19533), .ZN(n14183) );
  INV_X1 U17580 ( .A(n14185), .ZN(n14186) );
  OAI21_X1 U17581 ( .B1(n14186), .B2(n19265), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n14187) );
  OAI21_X1 U17582 ( .B1(n19271), .B2(n19462), .A(n14187), .ZN(n19266) );
  INV_X1 U17583 ( .A(n19265), .ZN(n14194) );
  AOI22_X1 U17584 ( .A1(n19303), .A2(n19668), .B1(n19267), .B2(n19666), .ZN(
        n14188) );
  OAI21_X1 U17585 ( .B1(n14189), .B2(n14194), .A(n14188), .ZN(n14190) );
  AOI21_X1 U17586 ( .B1(n19266), .B2(n19664), .A(n14190), .ZN(n14191) );
  OAI21_X1 U17587 ( .B1(n19270), .B2(n14192), .A(n14191), .ZN(P2_U3070) );
  AOI22_X1 U17588 ( .A1(n19267), .A2(n19576), .B1(n19303), .B2(n19575), .ZN(
        n14193) );
  OAI21_X1 U17589 ( .B1(n14195), .B2(n14194), .A(n14193), .ZN(n14196) );
  AOI21_X1 U17590 ( .B1(n19266), .B2(n19574), .A(n14196), .ZN(n14197) );
  OAI21_X1 U17591 ( .B1(n19270), .B2(n14198), .A(n14197), .ZN(P2_U3064) );
  XNOR2_X1 U17592 ( .A(n14200), .B(n14199), .ZN(n19048) );
  INV_X1 U17593 ( .A(n19048), .ZN(n15576) );
  OAI22_X1 U17594 ( .A1(n19002), .A2(n10790), .B1(n14202), .B2(n19027), .ZN(
        n14210) );
  NAND2_X1 U17595 ( .A1(n9838), .A2(n18993), .ZN(n19034) );
  INV_X1 U17596 ( .A(n19034), .ZN(n14201) );
  OAI211_X1 U17597 ( .C1(n14203), .C2(n14202), .A(n14201), .B(n18896), .ZN(
        n14207) );
  AOI22_X1 U17598 ( .A1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n18997), .B1(
        P2_REIP_REG_15__SCAN_IN), .B2(n19017), .ZN(n14204) );
  NAND2_X1 U17599 ( .A1(n19155), .A2(n14204), .ZN(n14205) );
  AOI21_X1 U17600 ( .B1(n16234), .B2(n19020), .A(n14205), .ZN(n14206) );
  OAI211_X1 U17601 ( .C1(n18984), .C2(n14208), .A(n14207), .B(n14206), .ZN(
        n14209) );
  AOI211_X1 U17602 ( .C1(n19016), .C2(n15576), .A(n14210), .B(n14209), .ZN(
        n14211) );
  INV_X1 U17603 ( .A(n14211), .ZN(P2_U2840) );
  INV_X1 U17604 ( .A(DATAI_10_), .ZN(n14212) );
  INV_X1 U17605 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n16458) );
  MUX2_X1 U17606 ( .A(n14212), .B(n16458), .S(n20099), .Z(n20012) );
  INV_X1 U17607 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n14213) );
  OAI222_X1 U17608 ( .A1(n14960), .A2(n14814), .B1(n20012), .B2(n14379), .C1(
        n14213), .C2(n14815), .ZN(P1_U2894) );
  NAND2_X1 U17609 ( .A1(n14252), .A2(n14248), .ZN(n14240) );
  NOR2_X1 U17610 ( .A1(n14240), .A2(n14241), .ZN(n14239) );
  INV_X1 U17611 ( .A(n14214), .ZN(n14217) );
  NOR2_X1 U17612 ( .A1(n14240), .A2(n14215), .ZN(n14381) );
  INV_X1 U17613 ( .A(n14381), .ZN(n14216) );
  OAI21_X1 U17614 ( .B1(n14239), .B2(n14217), .A(n14216), .ZN(n14312) );
  XNOR2_X1 U17615 ( .A(n14218), .B(n15100), .ZN(n15515) );
  INV_X1 U17616 ( .A(n15515), .ZN(n14224) );
  OAI22_X1 U17617 ( .A1(n15206), .A2(n19097), .B1(n14219), .B2(n19069), .ZN(
        n14223) );
  INV_X1 U17618 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n14221) );
  INV_X1 U17619 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n14220) );
  OAI22_X1 U17620 ( .A1(n15210), .A2(n14221), .B1(n15208), .B2(n14220), .ZN(
        n14222) );
  AOI211_X1 U17621 ( .C1(n19099), .C2(n14224), .A(n14223), .B(n14222), .ZN(
        n14225) );
  OAI21_X1 U17622 ( .B1(n14312), .B2(n19103), .A(n14225), .ZN(P2_U2900) );
  OAI21_X1 U17623 ( .B1(n15555), .B2(n14226), .A(n15102), .ZN(n18887) );
  INV_X1 U17624 ( .A(n18887), .ZN(n15547) );
  OR2_X1 U17625 ( .A1(n14252), .A2(n14248), .ZN(n14227) );
  NAND2_X1 U17626 ( .A1(n14240), .A2(n14227), .ZN(n14238) );
  OAI22_X1 U17627 ( .A1(n15206), .A2(n19108), .B1(n19069), .B2(n14228), .ZN(
        n14229) );
  AOI21_X1 U17628 ( .B1(n19039), .B2(BUF1_REG_17__SCAN_IN), .A(n14229), .ZN(
        n14231) );
  NAND2_X1 U17629 ( .A1(n19038), .A2(BUF2_REG_17__SCAN_IN), .ZN(n14230) );
  OAI211_X1 U17630 ( .C1(n14238), .C2(n19103), .A(n14231), .B(n14230), .ZN(
        n14232) );
  AOI21_X1 U17631 ( .B1(n15547), .B2(n19099), .A(n14232), .ZN(n14233) );
  INV_X1 U17632 ( .A(n14233), .ZN(P2_U2902) );
  AND2_X1 U17633 ( .A1(n14088), .A2(n14234), .ZN(n14235) );
  NOR2_X1 U17634 ( .A1(n14244), .A2(n14235), .ZN(n15539) );
  INV_X1 U17635 ( .A(n15539), .ZN(n18886) );
  NOR2_X1 U17636 ( .A1(n18886), .A2(n15169), .ZN(n14236) );
  AOI21_X1 U17637 ( .B1(P2_EBX_REG_17__SCAN_IN), .B2(n15169), .A(n14236), .ZN(
        n14237) );
  OAI21_X1 U17638 ( .B1(n14238), .B2(n15124), .A(n14237), .ZN(P2_U2870) );
  AOI21_X1 U17639 ( .B1(n14241), .B2(n14240), .A(n14239), .ZN(n16226) );
  NAND2_X1 U17640 ( .A1(n16226), .A2(n15150), .ZN(n14247) );
  OR2_X1 U17641 ( .A1(n14244), .A2(n14243), .ZN(n14245) );
  NAND2_X1 U17642 ( .A1(n14242), .A2(n14245), .ZN(n15325) );
  INV_X1 U17643 ( .A(n15325), .ZN(n15524) );
  NAND2_X1 U17644 ( .A1(n15524), .A2(n15157), .ZN(n14246) );
  OAI211_X1 U17645 ( .C1(n15157), .C2(n10800), .A(n14247), .B(n14246), .ZN(
        P2_U2869) );
  AND2_X1 U17646 ( .A1(n14252), .A2(n14248), .ZN(n14250) );
  NAND2_X1 U17647 ( .A1(n14252), .A2(n14251), .ZN(n14337) );
  OAI21_X1 U17648 ( .B1(n14383), .B2(n14253), .A(n14337), .ZN(n15171) );
  OR2_X1 U17649 ( .A1(n14255), .A2(n14254), .ZN(n14256) );
  NAND2_X1 U17650 ( .A1(n13086), .A2(n14256), .ZN(n18870) );
  INV_X1 U17651 ( .A(n18870), .ZN(n14263) );
  OAI22_X1 U17652 ( .A1(n15206), .A2(n14258), .B1(n14257), .B2(n19069), .ZN(
        n14262) );
  INV_X1 U17653 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n14260) );
  INV_X1 U17654 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n14259) );
  OAI22_X1 U17655 ( .A1(n15210), .A2(n14260), .B1(n15208), .B2(n14259), .ZN(
        n14261) );
  AOI211_X1 U17656 ( .C1(n19099), .C2(n14263), .A(n14262), .B(n14261), .ZN(
        n14264) );
  OAI21_X1 U17657 ( .B1(n15171), .B2(n19103), .A(n14264), .ZN(P2_U2898) );
  XNOR2_X1 U17658 ( .A(n14265), .B(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n14284) );
  NAND2_X1 U17659 ( .A1(n16254), .A2(n16255), .ZN(n14267) );
  XOR2_X1 U17660 ( .A(n14267), .B(n14266), .Z(n14282) );
  OAI21_X1 U17661 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n14269), .A(
        n14268), .ZN(n16278) );
  NOR2_X1 U17662 ( .A1(n19712), .A2(n19155), .ZN(n14270) );
  AOI221_X1 U17663 ( .B1(n16283), .B2(n14271), .C1(n16278), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n14270), .ZN(n14272) );
  INV_X1 U17664 ( .A(n14272), .ZN(n14277) );
  OR2_X1 U17665 ( .A1(n14273), .A2(n14274), .ZN(n14275) );
  NAND2_X1 U17666 ( .A1(n14274), .A2(n14273), .ZN(n16276) );
  NAND2_X1 U17667 ( .A1(n14275), .A2(n16276), .ZN(n19066) );
  OAI22_X1 U17668 ( .A1(n19066), .A2(n19185), .B1(n19179), .B2(n18979), .ZN(
        n14276) );
  AOI211_X1 U17669 ( .C1(n14282), .C2(n19188), .A(n14277), .B(n14276), .ZN(
        n14278) );
  OAI21_X1 U17670 ( .B1(n14284), .B2(n19174), .A(n14278), .ZN(P2_U3039) );
  OAI22_X1 U17671 ( .A1(n19712), .A2(n19155), .B1(n15396), .B2(n18975), .ZN(
        n14279) );
  AOI21_X1 U17672 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n15338), .A(
        n14279), .ZN(n14280) );
  OAI21_X1 U17673 ( .B1(n13862), .B2(n18979), .A(n14280), .ZN(n14281) );
  AOI21_X1 U17674 ( .B1(n14282), .B2(n11114), .A(n14281), .ZN(n14283) );
  OAI21_X1 U17675 ( .B1(n14284), .B2(n19148), .A(n14283), .ZN(P2_U3007) );
  AND2_X1 U17676 ( .A1(n14680), .A2(n14285), .ZN(n14286) );
  NOR2_X1 U17677 ( .A1(n14327), .A2(n14286), .ZN(n15991) );
  INV_X1 U17678 ( .A(n15991), .ZN(n14307) );
  INV_X1 U17679 ( .A(DATAI_14_), .ZN(n14288) );
  NAND2_X1 U17680 ( .A1(n20099), .A2(BUF1_REG_14__SCAN_IN), .ZN(n14287) );
  OAI21_X1 U17681 ( .B1(n20099), .B2(n14288), .A(n14287), .ZN(n20030) );
  AOI22_X1 U17682 ( .A1(n14826), .A2(n20030), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n15946), .ZN(n14289) );
  OAI21_X1 U17683 ( .B1(n14307), .B2(n14828), .A(n14289), .ZN(P1_U2890) );
  INV_X1 U17684 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n15919) );
  NAND2_X1 U17685 ( .A1(n14466), .A2(n15919), .ZN(n14295) );
  INV_X1 U17686 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14290) );
  NAND2_X1 U17687 ( .A1(n14291), .A2(n14290), .ZN(n14293) );
  NAND2_X1 U17688 ( .A1(n14467), .A2(n15919), .ZN(n14292) );
  NAND3_X1 U17689 ( .A1(n14293), .A2(n14522), .A3(n14292), .ZN(n14294) );
  INV_X1 U17690 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15944) );
  NAND2_X1 U17691 ( .A1(n14467), .A2(n15944), .ZN(n14297) );
  NAND2_X1 U17692 ( .A1(n14522), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n14296) );
  NAND3_X1 U17693 ( .A1(n14297), .A2(n13781), .A3(n14296), .ZN(n14298) );
  OAI21_X1 U17694 ( .B1(n14472), .B2(P1_EBX_REG_12__SCAN_IN), .A(n14298), .ZN(
        n15907) );
  INV_X1 U17695 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16098) );
  NAND2_X1 U17696 ( .A1(n13781), .A2(n16098), .ZN(n14301) );
  INV_X1 U17697 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14299) );
  NAND2_X1 U17698 ( .A1(n14467), .A2(n14299), .ZN(n14300) );
  NAND3_X1 U17699 ( .A1(n14301), .A2(n14522), .A3(n14300), .ZN(n14302) );
  OAI21_X1 U17700 ( .B1(n14474), .B2(P1_EBX_REG_13__SCAN_IN), .A(n14302), .ZN(
        n14683) );
  MUX2_X1 U17701 ( .A(n14472), .B(n14522), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n14303) );
  OAI21_X1 U17702 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n14525), .A(
        n14303), .ZN(n14304) );
  NAND2_X1 U17703 ( .A1(n14682), .A2(n14304), .ZN(n14305) );
  AND2_X1 U17704 ( .A1(n14333), .A2(n14305), .ZN(n16086) );
  AOI22_X1 U17705 ( .A1(n16086), .A2(n15941), .B1(P1_EBX_REG_14__SCAN_IN), 
        .B2(n14763), .ZN(n14306) );
  OAI21_X1 U17706 ( .B1(n14307), .B2(n14750), .A(n14306), .ZN(P1_U2858) );
  NAND2_X1 U17707 ( .A1(n14242), .A2(n14308), .ZN(n14309) );
  NAND2_X1 U17708 ( .A1(n9653), .A2(n14309), .ZN(n15516) );
  NOR2_X1 U17709 ( .A1(n15516), .A2(n15169), .ZN(n14310) );
  AOI21_X1 U17710 ( .B1(P2_EBX_REG_19__SCAN_IN), .B2(n15169), .A(n14310), .ZN(
        n14311) );
  OAI21_X1 U17711 ( .B1(n14312), .B2(n15124), .A(n14311), .ZN(P2_U2868) );
  XOR2_X1 U17712 ( .A(n14677), .B(n14161), .Z(n14315) );
  INV_X1 U17713 ( .A(n14313), .ZN(n14314) );
  AOI21_X1 U17714 ( .B1(n14315), .B2(n14314), .A(n14676), .ZN(n16002) );
  NAND2_X1 U17715 ( .A1(n14317), .A2(n14316), .ZN(n14318) );
  NAND2_X1 U17716 ( .A1(n15908), .A2(n14318), .ZN(n15922) );
  OAI22_X1 U17717 ( .A1(n15922), .A2(n14761), .B1(n15919), .B2(n15945), .ZN(
        n14319) );
  AOI21_X1 U17718 ( .B1(n16002), .B2(n15942), .A(n14319), .ZN(n14320) );
  INV_X1 U17719 ( .A(n14320), .ZN(P1_U2861) );
  INV_X1 U17720 ( .A(n16002), .ZN(n14324) );
  INV_X1 U17721 ( .A(DATAI_11_), .ZN(n14322) );
  MUX2_X1 U17722 ( .A(n14322), .B(n14321), .S(n20099), .Z(n20017) );
  INV_X1 U17723 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14323) );
  OAI222_X1 U17724 ( .A1(n14324), .A2(n14814), .B1(n20017), .B2(n14379), .C1(
        n14323), .C2(n14815), .ZN(P1_U2893) );
  INV_X1 U17725 ( .A(n14358), .ZN(n14325) );
  OAI21_X1 U17726 ( .B1(n14327), .B2(n14326), .A(n14325), .ZN(n14939) );
  INV_X1 U17727 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14352) );
  NAND2_X1 U17728 ( .A1(n14466), .A2(n14352), .ZN(n14331) );
  INV_X1 U17729 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14921) );
  NAND2_X1 U17730 ( .A1(n13781), .A2(n14921), .ZN(n14329) );
  NAND2_X1 U17731 ( .A1(n14467), .A2(n14352), .ZN(n14328) );
  NAND3_X1 U17732 ( .A1(n14329), .A2(n14522), .A3(n14328), .ZN(n14330) );
  AND2_X1 U17733 ( .A1(n14333), .A2(n14332), .ZN(n14334) );
  NOR2_X1 U17734 ( .A1(n14371), .A2(n14334), .ZN(n16076) );
  NOR2_X1 U17735 ( .A1(n15945), .A2(n14352), .ZN(n14335) );
  AOI21_X1 U17736 ( .B1(n16076), .B2(n15941), .A(n14335), .ZN(n14336) );
  OAI21_X1 U17737 ( .B1(n14939), .B2(n14750), .A(n14336), .ZN(P1_U2857) );
  INV_X1 U17738 ( .A(n14337), .ZN(n14339) );
  OAI21_X1 U17739 ( .B1(n14339), .B2(n14338), .A(n9638), .ZN(n15165) );
  INV_X1 U17740 ( .A(n15489), .ZN(n14344) );
  OAI22_X1 U17741 ( .A1(n15206), .A2(n19068), .B1(n14340), .B2(n19069), .ZN(
        n14343) );
  INV_X1 U17742 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n14341) );
  OAI22_X1 U17743 ( .A1(n15210), .A2(n14341), .B1(n15208), .B2(n18185), .ZN(
        n14342) );
  AOI211_X1 U17744 ( .C1(n19099), .C2(n14344), .A(n14343), .B(n14342), .ZN(
        n14345) );
  OAI21_X1 U17745 ( .B1(n15165), .B2(n19103), .A(n14345), .ZN(P2_U2897) );
  NAND2_X1 U17746 ( .A1(n15911), .A2(n15837), .ZN(n19939) );
  INV_X1 U17747 ( .A(n19939), .ZN(n14639) );
  NAND2_X1 U17748 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .ZN(n14350) );
  INV_X1 U17749 ( .A(n14350), .ZN(n14349) );
  INV_X1 U17750 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n16104) );
  INV_X1 U17751 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n19879) );
  INV_X1 U17752 ( .A(n14346), .ZN(n14347) );
  NOR3_X1 U17753 ( .A1(n19879), .A2(n14347), .A3(n19869), .ZN(n15927) );
  NAND2_X1 U17754 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n15927), .ZN(n15928) );
  NOR3_X1 U17755 ( .A1(n16104), .A2(n15064), .A3(n15928), .ZN(n15874) );
  OAI21_X1 U17756 ( .B1(n15874), .B2(n15911), .A(n15837), .ZN(n15914) );
  INV_X1 U17757 ( .A(n15914), .ZN(n14348) );
  OAI21_X1 U17758 ( .B1(n14639), .B2(n14349), .A(n14348), .ZN(n15902) );
  NOR2_X1 U17759 ( .A1(n19940), .A2(n14935), .ZN(n14354) );
  NOR4_X1 U17760 ( .A1(n15911), .A2(n16104), .A3(n15064), .A4(n15928), .ZN(
        n15865) );
  INV_X1 U17761 ( .A(n15865), .ZN(n15900) );
  NOR3_X1 U17762 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n14350), .A3(n15900), 
        .ZN(n14363) );
  AOI211_X1 U17763 ( .C1(n19926), .C2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n19913), .B(n14363), .ZN(n14351) );
  OAI21_X1 U17764 ( .B1(n19895), .B2(n14352), .A(n14351), .ZN(n14353) );
  AOI211_X1 U17765 ( .C1(n15902), .C2(P1_REIP_REG_15__SCAN_IN), .A(n14354), 
        .B(n14353), .ZN(n14356) );
  NAND2_X1 U17766 ( .A1(n16076), .A2(n19945), .ZN(n14355) );
  OAI211_X1 U17767 ( .C1(n14939), .C2(n15891), .A(n14356), .B(n14355), .ZN(
        P1_U2825) );
  OR2_X1 U17768 ( .A1(n14358), .A2(n14357), .ZN(n14359) );
  NAND2_X1 U17769 ( .A1(n14752), .A2(n14359), .ZN(n15980) );
  OAI22_X1 U17770 ( .A1(n14817), .A2(n20112), .B1(n19976), .B2(n14815), .ZN(
        n14360) );
  AOI21_X1 U17771 ( .B1(n15948), .B2(DATAI_16_), .A(n14360), .ZN(n14362) );
  NAND2_X1 U17772 ( .A1(n14819), .A2(BUF1_REG_16__SCAN_IN), .ZN(n14361) );
  OAI211_X1 U17773 ( .C1(n15980), .C2(n14828), .A(n14362), .B(n14361), .ZN(
        P1_U2888) );
  NAND3_X1 U17774 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(P1_REIP_REG_14__SCAN_IN), 
        .A3(P1_REIP_REG_13__SCAN_IN), .ZN(n14482) );
  NOR2_X1 U17775 ( .A1(n14482), .A2(n15900), .ZN(n15896) );
  INV_X1 U17776 ( .A(n15896), .ZN(n14365) );
  NOR2_X1 U17777 ( .A1(n14363), .A2(n15902), .ZN(n14364) );
  MUX2_X1 U17778 ( .A(n14365), .B(n14364), .S(P1_REIP_REG_16__SCAN_IN), .Z(
        n14377) );
  INV_X1 U17779 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n20905) );
  NAND2_X1 U17780 ( .A1(n14366), .A2(n20905), .ZN(n14369) );
  INV_X1 U17781 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n20829) );
  NAND2_X1 U17782 ( .A1(n14467), .A2(n20905), .ZN(n14367) );
  OAI211_X1 U17783 ( .C1(n14475), .C2(n20829), .A(n14367), .B(n13781), .ZN(
        n14368) );
  NOR2_X1 U17784 ( .A1(n14371), .A2(n14370), .ZN(n14372) );
  OR2_X1 U17785 ( .A1(n14756), .A2(n14372), .ZN(n16069) );
  OAI22_X1 U17786 ( .A1(n16069), .A2(n19897), .B1(n19895), .B2(n20905), .ZN(
        n14373) );
  INV_X1 U17787 ( .A(n14373), .ZN(n14374) );
  OAI21_X1 U17788 ( .B1(n15984), .B2(n19940), .A(n14374), .ZN(n14375) );
  AOI211_X1 U17789 ( .C1(n19926), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n19913), .B(n14375), .ZN(n14376) );
  OAI211_X1 U17790 ( .C1(n15980), .C2(n15891), .A(n14377), .B(n14376), .ZN(
        P1_U2824) );
  OAI222_X1 U17791 ( .A1(n14814), .A2(n14939), .B1(n14379), .B2(n14378), .C1(
        n14815), .C2(n13245), .ZN(P1_U2889) );
  NOR2_X1 U17792 ( .A1(n14381), .A2(n14380), .ZN(n14382) );
  MUX2_X1 U17793 ( .A(n18874), .B(n14384), .S(n15169), .Z(n14385) );
  OAI21_X1 U17794 ( .B1(n16220), .B2(n15124), .A(n14385), .ZN(P2_U2867) );
  OAI222_X1 U17795 ( .A1(n16069), .A2(n14761), .B1(n20905), .B2(n15945), .C1(
        n15980), .C2(n14750), .ZN(P1_U2856) );
  INV_X1 U17796 ( .A(n18612), .ZN(n18621) );
  OAI211_X1 U17797 ( .C1(n18621), .C2(n18768), .A(n9591), .B(n18604), .ZN(
        n18146) );
  NOR2_X1 U17798 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18146), .ZN(n14387) );
  NOR2_X1 U17799 ( .A1(n18773), .A2(n14386), .ZN(n18668) );
  NAND2_X1 U17800 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18668), .ZN(n18761) );
  OAI21_X1 U17801 ( .B1(n14387), .B2(n18761), .A(n18262), .ZN(n18153) );
  INV_X1 U17802 ( .A(n18153), .ZN(n14388) );
  INV_X1 U17803 ( .A(n18149), .ZN(n18810) );
  NAND2_X1 U17804 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n17684) );
  AOI22_X1 U17805 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_3__SCAN_IN), .B1(n18810), .B2(n17684), .ZN(n15691) );
  NOR2_X1 U17806 ( .A1(n14388), .A2(n15691), .ZN(n14390) );
  INV_X1 U17807 ( .A(n18239), .ZN(n18504) );
  NOR2_X1 U17808 ( .A1(n18763), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18197) );
  OR2_X1 U17809 ( .A1(n18197), .A2(n14388), .ZN(n15689) );
  OR2_X1 U17810 ( .A1(n18504), .A2(n15689), .ZN(n14389) );
  MUX2_X1 U17811 ( .A(n14390), .B(n14389), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  NAND2_X1 U17812 ( .A1(n15169), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n14391) );
  OAI21_X1 U17813 ( .B1(n14392), .B2(n15169), .A(n14391), .ZN(P2_U2856) );
  NOR2_X1 U17814 ( .A1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n14393) );
  AND2_X1 U17815 ( .A1(n14393), .A2(n14921), .ZN(n14400) );
  NAND2_X1 U17816 ( .A1(n14395), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n14396) );
  INV_X1 U17817 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16119) );
  NOR2_X1 U17818 ( .A1(n9626), .A2(n16119), .ZN(n14398) );
  NAND2_X1 U17819 ( .A1(n15987), .A2(n16119), .ZN(n14399) );
  OR2_X1 U17820 ( .A1(n9625), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14923) );
  NAND2_X1 U17821 ( .A1(n9626), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14401) );
  NAND2_X1 U17822 ( .A1(n14923), .A2(n14401), .ZN(n15975) );
  NAND2_X1 U17823 ( .A1(n9626), .A2(n14921), .ZN(n15973) );
  NAND2_X1 U17824 ( .A1(n14922), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14406) );
  OR2_X2 U17825 ( .A1(n9626), .A2(n16098), .ZN(n15985) );
  NAND2_X1 U17826 ( .A1(n9626), .A2(n16098), .ZN(n14402) );
  NAND2_X1 U17827 ( .A1(n15985), .A2(n14402), .ZN(n14947) );
  INV_X1 U17828 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n16107) );
  NAND2_X1 U17829 ( .A1(n15987), .A2(n16107), .ZN(n14945) );
  NAND2_X1 U17830 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14403) );
  NAND2_X1 U17831 ( .A1(n9626), .A2(n14403), .ZN(n14943) );
  NAND2_X1 U17832 ( .A1(n14945), .A2(n14943), .ZN(n14404) );
  NOR2_X2 U17833 ( .A1(n14947), .A2(n14404), .ZN(n14914) );
  NAND2_X1 U17834 ( .A1(n14914), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n14405) );
  INV_X1 U17835 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n14916) );
  OR2_X1 U17836 ( .A1(n15987), .A2(n14916), .ZN(n14407) );
  NOR2_X1 U17837 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n14941) );
  AND2_X1 U17838 ( .A1(n14941), .A2(n16107), .ZN(n14408) );
  NOR2_X1 U17839 ( .A1(n9626), .A2(n14408), .ZN(n14912) );
  AND3_X1 U17840 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14536) );
  NAND2_X1 U17841 ( .A1(n9619), .A2(n14906), .ZN(n14409) );
  NAND2_X1 U17842 ( .A1(n14409), .A2(n9626), .ZN(n15961) );
  INV_X1 U17843 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14528) );
  INV_X1 U17844 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n16065) );
  INV_X1 U17845 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14891) );
  INV_X1 U17846 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15025) );
  INV_X1 U17847 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14877) );
  INV_X1 U17848 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15009) );
  INV_X1 U17849 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n16045) );
  NAND3_X1 U17850 ( .A1(n14877), .A2(n15009), .A3(n16045), .ZN(n14849) );
  INV_X1 U17851 ( .A(n14849), .ZN(n14410) );
  NAND2_X1 U17852 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15002) );
  NOR2_X1 U17853 ( .A1(n15002), .A2(n15009), .ZN(n14538) );
  INV_X1 U17854 ( .A(n14538), .ZN(n14848) );
  NAND2_X1 U17855 ( .A1(n14847), .A2(n14848), .ZN(n14413) );
  NAND2_X1 U17856 ( .A1(n14412), .A2(n15987), .ZN(n14876) );
  NAND3_X1 U17857 ( .A1(n14413), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14876), .ZN(n14860) );
  AND2_X1 U17858 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14982) );
  AND2_X1 U17859 ( .A1(n9626), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14414) );
  NAND2_X1 U17860 ( .A1(n14982), .A2(n14414), .ZN(n14415) );
  NOR2_X1 U17861 ( .A1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14983) );
  AND2_X1 U17862 ( .A1(n9688), .A2(n14983), .ZN(n14416) );
  AND3_X1 U17863 ( .A1(n14869), .A2(n14416), .A3(n14860), .ZN(n14417) );
  XNOR2_X1 U17864 ( .A(n14420), .B(n14537), .ZN(n14556) );
  NAND2_X1 U17865 ( .A1(n16052), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14550) );
  NAND2_X1 U17866 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14421) );
  OAI211_X1 U17867 ( .C1(n16019), .C2(n14422), .A(n14550), .B(n14421), .ZN(
        n14423) );
  AOI21_X1 U17868 ( .B1(n14599), .B2(n16022), .A(n14423), .ZN(n14424) );
  OAI21_X1 U17869 ( .B1(n14556), .B2(n19850), .A(n14424), .ZN(P1_U2968) );
  XNOR2_X1 U17870 ( .A(n9626), .B(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n14425) );
  XNOR2_X1 U17871 ( .A(n14426), .B(n14425), .ZN(n14436) );
  NAND3_X1 U17872 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n14532) );
  NOR2_X1 U17873 ( .A1(n15060), .A2(n14532), .ZN(n14529) );
  INV_X1 U17874 ( .A(n16131), .ZN(n14545) );
  NOR2_X1 U17875 ( .A1(n14545), .A2(n15059), .ZN(n14543) );
  AOI21_X1 U17876 ( .B1(n14529), .B2(n14427), .A(n14543), .ZN(n16117) );
  OAI22_X1 U17877 ( .A1(n19874), .A2(n16068), .B1(n19879), .B2(n16103), .ZN(
        n14428) );
  AOI21_X1 U17878 ( .B1(n16117), .B2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n14428), .ZN(n14431) );
  NAND2_X1 U17879 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16124) );
  INV_X1 U17880 ( .A(n14429), .ZN(n16083) );
  NAND2_X1 U17881 ( .A1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n16143), .ZN(
        n16140) );
  NOR2_X1 U17882 ( .A1(n16124), .A2(n16140), .ZN(n16118) );
  NAND2_X1 U17883 ( .A1(n16118), .A2(n16119), .ZN(n14430) );
  OAI211_X1 U17884 ( .C1(n14436), .C2(n16111), .A(n14431), .B(n14430), .ZN(
        P1_U3022) );
  OAI22_X1 U17885 ( .A1(n16026), .A2(n11911), .B1(n16103), .B2(n19879), .ZN(
        n14433) );
  NOR2_X1 U17886 ( .A1(n19868), .A2(n20102), .ZN(n14432) );
  AOI211_X1 U17887 ( .C1(n16021), .C2(n14434), .A(n14433), .B(n14432), .ZN(
        n14435) );
  OAI21_X1 U17888 ( .B1(n14436), .B2(n19850), .A(n14435), .ZN(P1_U2990) );
  AOI22_X1 U17889 ( .A1(n14525), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n14524), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14523) );
  NAND2_X1 U17890 ( .A1(n14522), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n14437) );
  NAND2_X1 U17891 ( .A1(n13781), .A2(n14437), .ZN(n14439) );
  NAND2_X1 U17892 ( .A1(n14467), .A2(n14762), .ZN(n14438) );
  NAND2_X1 U17893 ( .A1(n14439), .A2(n14438), .ZN(n14440) );
  OAI21_X1 U17894 ( .B1(n14474), .B2(P1_EBX_REG_17__SCAN_IN), .A(n14440), .ZN(
        n14757) );
  MUX2_X1 U17895 ( .A(n14472), .B(n14522), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n14441) );
  OAI21_X1 U17896 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n14525), .A(
        n14441), .ZN(n14745) );
  INV_X1 U17897 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14742) );
  NAND2_X1 U17898 ( .A1(n14466), .A2(n14742), .ZN(n14445) );
  NAND2_X1 U17899 ( .A1(n13781), .A2(n16065), .ZN(n14443) );
  NAND2_X1 U17900 ( .A1(n14467), .A2(n14742), .ZN(n14442) );
  NAND3_X1 U17901 ( .A1(n14443), .A2(n14522), .A3(n14442), .ZN(n14444) );
  NAND2_X1 U17902 ( .A1(n14445), .A2(n14444), .ZN(n14740) );
  INV_X1 U17903 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15940) );
  NAND2_X1 U17904 ( .A1(n14467), .A2(n15940), .ZN(n14447) );
  NAND2_X1 U17905 ( .A1(n14522), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14446) );
  NAND3_X1 U17906 ( .A1(n14447), .A2(n13781), .A3(n14446), .ZN(n14448) );
  OAI21_X1 U17907 ( .B1(n14472), .B2(P1_EBX_REG_20__SCAN_IN), .A(n14448), .ZN(
        n15800) );
  INV_X1 U17908 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n15846) );
  NAND2_X1 U17909 ( .A1(n14466), .A2(n15846), .ZN(n14452) );
  NAND2_X1 U17910 ( .A1(n13781), .A2(n15025), .ZN(n14450) );
  NAND2_X1 U17911 ( .A1(n14467), .A2(n15846), .ZN(n14449) );
  NAND3_X1 U17912 ( .A1(n14450), .A2(n14522), .A3(n14449), .ZN(n14451) );
  MUX2_X1 U17913 ( .A(n14472), .B(n14522), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n14453) );
  OAI21_X1 U17914 ( .B1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n14525), .A(
        n14453), .ZN(n14728) );
  INV_X1 U17915 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n15824) );
  NAND2_X1 U17916 ( .A1(n14466), .A2(n15824), .ZN(n14457) );
  NAND2_X1 U17917 ( .A1(n13781), .A2(n16045), .ZN(n14455) );
  NAND2_X1 U17918 ( .A1(n14467), .A2(n15824), .ZN(n14454) );
  NAND3_X1 U17919 ( .A1(n14455), .A2(n14522), .A3(n14454), .ZN(n14456) );
  MUX2_X1 U17920 ( .A(n14472), .B(n14522), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n14459) );
  OR2_X1 U17921 ( .A1(n14525), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14458) );
  AND2_X1 U17922 ( .A1(n14459), .A2(n14458), .ZN(n14713) );
  INV_X1 U17923 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n14708) );
  NAND2_X1 U17924 ( .A1(n14466), .A2(n14708), .ZN(n14463) );
  NAND2_X1 U17925 ( .A1(n13781), .A2(n15009), .ZN(n14461) );
  NAND2_X1 U17926 ( .A1(n14467), .A2(n14708), .ZN(n14460) );
  NAND3_X1 U17927 ( .A1(n14461), .A2(n14522), .A3(n14460), .ZN(n14462) );
  NAND2_X1 U17928 ( .A1(n14463), .A2(n14462), .ZN(n14670) );
  MUX2_X1 U17929 ( .A(n14472), .B(n14522), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n14465) );
  OR2_X1 U17930 ( .A1(n14525), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14464) );
  AND2_X1 U17931 ( .A1(n14465), .A2(n14464), .ZN(n14647) );
  INV_X1 U17932 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n20828) );
  NAND2_X1 U17933 ( .A1(n14466), .A2(n20828), .ZN(n14471) );
  INV_X1 U17934 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14992) );
  NAND2_X1 U17935 ( .A1(n13781), .A2(n14992), .ZN(n14469) );
  NAND2_X1 U17936 ( .A1(n14467), .A2(n20828), .ZN(n14468) );
  NAND3_X1 U17937 ( .A1(n14469), .A2(n14522), .A3(n14468), .ZN(n14470) );
  AND2_X1 U17938 ( .A1(n14471), .A2(n14470), .ZN(n14633) );
  MUX2_X1 U17939 ( .A(n14472), .B(n14522), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n14473) );
  OAI21_X1 U17940 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n14525), .A(
        n14473), .ZN(n14619) );
  OAI22_X1 U17941 ( .A1(n14525), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B1(
        n14524), .B2(P1_EBX_REG_29__SCAN_IN), .ZN(n14477) );
  OAI22_X1 U17942 ( .A1(n14477), .A2(n14475), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n14474), .ZN(n14614) );
  NAND2_X1 U17943 ( .A1(n14620), .A2(n14614), .ZN(n14613) );
  NAND2_X1 U17944 ( .A1(n14613), .A2(n14475), .ZN(n14478) );
  INV_X1 U17945 ( .A(n14620), .ZN(n14476) );
  AOI22_X1 U17946 ( .A1(n14478), .A2(n14477), .B1(n14476), .B2(n14522), .ZN(
        n14479) );
  XOR2_X1 U17947 ( .A(n14523), .B(n14479), .Z(n14966) );
  NAND2_X1 U17948 ( .A1(n14835), .A2(n19904), .ZN(n14497) );
  INV_X1 U17949 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n14485) );
  INV_X1 U17950 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14484) );
  INV_X1 U17951 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20707) );
  INV_X1 U17952 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n20830) );
  INV_X1 U17953 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n14483) );
  NOR3_X1 U17954 ( .A1(n20830), .A2(n14483), .A3(n14482), .ZN(n15875) );
  NAND4_X1 U17955 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .A3(n15874), .A4(n15875), .ZN(n15859) );
  NAND2_X1 U17956 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n15825) );
  NOR4_X1 U17957 ( .A1(n14484), .A2(n20707), .A3(n15859), .A4(n15825), .ZN(
        n15813) );
  NAND2_X1 U17958 ( .A1(P1_REIP_REG_24__SCAN_IN), .A2(n15813), .ZN(n14665) );
  NOR2_X1 U17959 ( .A1(n14485), .A2(n14665), .ZN(n14655) );
  NAND2_X1 U17960 ( .A1(n14655), .A2(P1_REIP_REG_26__SCAN_IN), .ZN(n14488) );
  NOR2_X1 U17961 ( .A1(n15911), .A2(n14488), .ZN(n14641) );
  NAND3_X1 U17962 ( .A1(n14641), .A2(P1_REIP_REG_27__SCAN_IN), .A3(
        P1_REIP_REG_28__SCAN_IN), .ZN(n14612) );
  INV_X1 U17963 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n14487) );
  INV_X1 U17964 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14486) );
  OAI21_X1 U17965 ( .B1(n14612), .B2(n14487), .A(n14486), .ZN(n14495) );
  AND2_X1 U17966 ( .A1(P1_REIP_REG_30__SCAN_IN), .A2(P1_REIP_REG_29__SCAN_IN), 
        .ZN(n14491) );
  NOR2_X1 U17967 ( .A1(n14488), .A2(n15918), .ZN(n14638) );
  AND2_X1 U17968 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n14489) );
  NAND2_X1 U17969 ( .A1(n14638), .A2(n14489), .ZN(n14490) );
  NAND2_X1 U17970 ( .A1(n19939), .A2(n14490), .ZN(n14627) );
  OAI21_X1 U17971 ( .B1(n14639), .B2(n14491), .A(n14627), .ZN(n14604) );
  INV_X1 U17972 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14498) );
  NOR2_X1 U17973 ( .A1(n19895), .A2(n14498), .ZN(n14494) );
  INV_X1 U17974 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14492) );
  OAI22_X1 U17975 ( .A1(n14492), .A2(n19941), .B1(n19940), .B2(n14833), .ZN(
        n14493) );
  AOI211_X1 U17976 ( .C1(n14495), .C2(n14604), .A(n14494), .B(n14493), .ZN(
        n14496) );
  OAI211_X1 U17977 ( .C1(n14966), .C2(n19897), .A(n14497), .B(n14496), .ZN(
        P1_U2810) );
  INV_X1 U17978 ( .A(n14835), .ZN(n14769) );
  OAI222_X1 U17979 ( .A1(n14750), .A2(n14769), .B1(n14498), .B2(n15945), .C1(
        n14761), .C2(n14966), .ZN(P1_U2842) );
  AND2_X1 U17980 ( .A1(n14500), .A2(n14499), .ZN(n14501) );
  XOR2_X1 U17981 ( .A(n14505), .B(n14504), .Z(n14519) );
  OAI211_X1 U17982 ( .C1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(n19162), .B(n14506), .ZN(n14512) );
  OAI21_X1 U17983 ( .B1(n9705), .B2(n14508), .A(n14507), .ZN(n19081) );
  INV_X1 U17984 ( .A(n19081), .ZN(n14510) );
  NAND2_X1 U17985 ( .A1(n18902), .A2(P2_REIP_REG_5__SCAN_IN), .ZN(n14516) );
  OAI21_X1 U17986 ( .B1(n18991), .B2(n19179), .A(n14516), .ZN(n14509) );
  AOI21_X1 U17987 ( .B1(n14510), .B2(n16296), .A(n14509), .ZN(n14511) );
  OAI211_X1 U17988 ( .C1(n19164), .C2(n14513), .A(n14512), .B(n14511), .ZN(
        n14514) );
  AOI21_X1 U17989 ( .B1(n14519), .B2(n19188), .A(n14514), .ZN(n14515) );
  OAI21_X1 U17990 ( .B1(n14521), .B2(n19174), .A(n14515), .ZN(P2_U3041) );
  OAI22_X1 U17991 ( .A1(n10754), .A2(n19154), .B1(n15396), .B2(n18990), .ZN(
        n14518) );
  OAI21_X1 U17992 ( .B1(n18991), .B2(n13862), .A(n14516), .ZN(n14517) );
  AOI211_X1 U17993 ( .C1(n14519), .C2(n11114), .A(n14518), .B(n14517), .ZN(
        n14520) );
  OAI21_X1 U17994 ( .B1(n19148), .B2(n14521), .A(n14520), .ZN(P2_U3009) );
  MUX2_X1 U17995 ( .A(n14523), .B(n14522), .S(n14613), .Z(n14527) );
  AOI22_X1 U17996 ( .A1(n14525), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n14524), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14526) );
  INV_X1 U17997 ( .A(n14703), .ZN(n14554) );
  NAND4_X1 U17998 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A4(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15031) );
  NOR2_X1 U17999 ( .A1(n14528), .A2(n15031), .ZN(n14540) );
  NAND3_X1 U18000 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .A3(n14529), .ZN(n15053) );
  NAND2_X1 U18001 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14530) );
  NOR2_X1 U18002 ( .A1(n15053), .A2(n14530), .ZN(n15021) );
  NAND2_X1 U18003 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15021), .ZN(
        n16082) );
  NAND2_X1 U18004 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n14531), .ZN(
        n14534) );
  INV_X1 U18005 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n16120) );
  OR3_X1 U18006 ( .A1(n16120), .A2(n16119), .A3(n14532), .ZN(n15054) );
  NOR3_X1 U18007 ( .A1(n14534), .A2(n14533), .A3(n15054), .ZN(n15056) );
  NAND3_X1 U18008 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A3(n15056), .ZN(n15022) );
  NOR2_X1 U18009 ( .A1(n16098), .A2(n15022), .ZN(n15033) );
  NAND2_X1 U18010 ( .A1(n14535), .A2(n15033), .ZN(n16041) );
  OAI21_X1 U18011 ( .B1(n16082), .B2(n15055), .A(n16041), .ZN(n15042) );
  NAND4_X1 U18012 ( .A1(n14536), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n14540), .A4(n15042), .ZN(n16044) );
  NOR2_X1 U18013 ( .A1(n16044), .A2(n14848), .ZN(n16034) );
  NAND3_X1 U18014 ( .A1(n14993), .A2(n14982), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14961) );
  NAND2_X1 U18015 ( .A1(n14537), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14552) );
  INV_X1 U18016 ( .A(n14982), .ZN(n14549) );
  NOR2_X1 U18017 ( .A1(n14538), .A2(n15794), .ZN(n14546) );
  NAND2_X1 U18018 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n16054) );
  NAND2_X1 U18019 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15024) );
  INV_X1 U18020 ( .A(n15024), .ZN(n14544) );
  NAND2_X1 U18021 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n14540), .ZN(
        n15017) );
  INV_X1 U18022 ( .A(n16082), .ZN(n15032) );
  OAI221_X1 U18023 ( .B1(n15055), .B2(n15032), .C1(n15055), .C2(n14540), .A(
        n14539), .ZN(n14541) );
  AOI221_X1 U18024 ( .B1(n15022), .B2(n14542), .C1(n15017), .C2(n14542), .A(
        n14541), .ZN(n16064) );
  AOI21_X1 U18025 ( .B1(n14544), .B2(n9595), .A(n14543), .ZN(n16051) );
  AOI21_X1 U18026 ( .B1(n14545), .B2(n16054), .A(n16051), .ZN(n15012) );
  OAI21_X1 U18027 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15055), .A(
        n15012), .ZN(n16042) );
  AOI211_X1 U18028 ( .C1(n15002), .C2(n14547), .A(n14546), .B(n16042), .ZN(
        n15010) );
  NAND2_X1 U18029 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n15010), .ZN(
        n16032) );
  INV_X1 U18030 ( .A(n16032), .ZN(n14548) );
  NAND2_X1 U18031 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n14548), .ZN(
        n14980) );
  NAND2_X1 U18032 ( .A1(n15010), .A2(n16131), .ZN(n14981) );
  OAI21_X1 U18033 ( .B1(n14549), .B2(n14980), .A(n14981), .ZN(n14971) );
  OAI211_X1 U18034 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16131), .A(
        n14971), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14962) );
  NAND3_X1 U18035 ( .A1(n14962), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14981), .ZN(n14551) );
  OAI211_X1 U18036 ( .C1(n14961), .C2(n14552), .A(n14551), .B(n14550), .ZN(
        n14553) );
  AOI21_X1 U18037 ( .B1(n16142), .B2(n14554), .A(n14553), .ZN(n14555) );
  OAI21_X1 U18038 ( .B1(n14556), .B2(n16111), .A(n14555), .ZN(P1_U3000) );
  NOR2_X1 U18039 ( .A1(n11634), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n14557) );
  AOI21_X1 U18040 ( .B1(n9621), .B2(n14558), .A(n14557), .ZN(n15734) );
  OAI21_X1 U18041 ( .B1(n15734), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n13902), 
        .ZN(n14559) );
  AOI22_X1 U18042 ( .A1(n14561), .A2(n14562), .B1(n14560), .B2(n14559), .ZN(
        n14565) );
  AOI21_X1 U18043 ( .B1(n15732), .B2(n16151), .A(n14564), .ZN(n14563) );
  OAI22_X1 U18044 ( .A1(n14565), .A2(n14564), .B1(n14563), .B2(n14562), .ZN(
        P1_U3474) );
  NOR2_X1 U18045 ( .A1(n16172), .A2(n15169), .ZN(n14566) );
  AOI21_X1 U18046 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n15169), .A(n14566), .ZN(
        n14567) );
  OAI21_X1 U18047 ( .B1(n14568), .B2(n15124), .A(n14567), .ZN(P2_U2857) );
  NAND2_X1 U18048 ( .A1(n14571), .A2(n14570), .ZN(n15114) );
  INV_X1 U18049 ( .A(n19103), .ZN(n19086) );
  NAND2_X1 U18050 ( .A1(n15114), .A2(n19086), .ZN(n14577) );
  INV_X1 U18051 ( .A(n15406), .ZN(n14574) );
  OAI22_X1 U18052 ( .A1(n15206), .A2(n19051), .B1(n19069), .B2(n14572), .ZN(
        n14573) );
  AOI21_X1 U18053 ( .B1(n14574), .B2(n19099), .A(n14573), .ZN(n14576) );
  AOI22_X1 U18054 ( .A1(n19039), .A2(BUF1_REG_29__SCAN_IN), .B1(n19038), .B2(
        BUF2_REG_29__SCAN_IN), .ZN(n14575) );
  OAI211_X1 U18055 ( .C1(n14569), .C2(n14577), .A(n14576), .B(n14575), .ZN(
        P2_U2890) );
  NAND2_X1 U18056 ( .A1(n14578), .A2(n14579), .ZN(n14586) );
  AOI21_X1 U18057 ( .B1(n14580), .B2(n13095), .A(n14579), .ZN(n14584) );
  NOR2_X1 U18058 ( .A1(n14582), .A2(n14581), .ZN(n14583) );
  NOR2_X1 U18059 ( .A1(n14584), .A2(n14583), .ZN(n14585) );
  NAND2_X1 U18060 ( .A1(n14586), .A2(n14585), .ZN(n15751) );
  OR2_X1 U18061 ( .A1(n14587), .A2(n15762), .ZN(n14591) );
  NAND2_X1 U18062 ( .A1(n14589), .A2(n14588), .ZN(n14590) );
  NAND2_X1 U18063 ( .A1(n14591), .A2(n14590), .ZN(n19844) );
  INV_X1 U18064 ( .A(n19844), .ZN(n14597) );
  OR2_X1 U18065 ( .A1(n14593), .A2(n14592), .ZN(n14594) );
  OAI211_X1 U18066 ( .C1(n14596), .C2(n14595), .A(n14594), .B(n20760), .ZN(
        n20751) );
  NAND2_X1 U18067 ( .A1(n14597), .A2(n20751), .ZN(n15754) );
  AND2_X1 U18068 ( .A1(n15754), .A2(n14598), .ZN(n19852) );
  MUX2_X1 U18069 ( .A(P1_MORE_REG_SCAN_IN), .B(n15751), .S(n19852), .Z(
        P1_U3484) );
  NAND2_X1 U18070 ( .A1(n14599), .A2(n19904), .ZN(n14606) );
  INV_X1 U18071 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n14600) );
  NAND3_X1 U18072 ( .A1(n14600), .A2(P1_REIP_REG_29__SCAN_IN), .A3(
        P1_REIP_REG_30__SCAN_IN), .ZN(n14602) );
  AOI22_X1 U18073 ( .A1(n19938), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19926), .ZN(n14601) );
  OAI21_X1 U18074 ( .B1(n14612), .B2(n14602), .A(n14601), .ZN(n14603) );
  AOI21_X1 U18075 ( .B1(P1_REIP_REG_31__SCAN_IN), .B2(n14604), .A(n14603), 
        .ZN(n14605) );
  OAI211_X1 U18076 ( .C1(n14703), .C2(n19897), .A(n14606), .B(n14605), .ZN(
        P1_U2809) );
  INV_X1 U18077 ( .A(n14627), .ZN(n14617) );
  AOI22_X1 U18078 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19926), .B1(
        n19927), .B2(n14839), .ZN(n14611) );
  NAND2_X1 U18079 ( .A1(n19938), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14610) );
  OAI211_X1 U18080 ( .C1(n14612), .C2(P1_REIP_REG_29__SCAN_IN), .A(n14611), 
        .B(n14610), .ZN(n14616) );
  OAI21_X1 U18081 ( .B1(n14620), .B2(n14614), .A(n14613), .ZN(n14975) );
  NOR2_X1 U18082 ( .A1(n14975), .A2(n19897), .ZN(n14615) );
  AOI211_X1 U18083 ( .C1(n14617), .C2(P1_REIP_REG_29__SCAN_IN), .A(n14616), 
        .B(n14615), .ZN(n14618) );
  OAI21_X1 U18084 ( .B1(n14846), .B2(n15891), .A(n14618), .ZN(P1_U2811) );
  AND2_X1 U18085 ( .A1(n14635), .A2(n14619), .ZN(n14621) );
  OR2_X1 U18086 ( .A1(n14621), .A2(n14620), .ZN(n14988) );
  INV_X1 U18087 ( .A(n14622), .ZN(n14625) );
  INV_X1 U18088 ( .A(n14623), .ZN(n14624) );
  AOI21_X1 U18089 ( .B1(n14625), .B2(n14624), .A(n14607), .ZN(n14857) );
  NAND2_X1 U18090 ( .A1(n14857), .A2(n19904), .ZN(n14632) );
  OAI22_X1 U18091 ( .A1(n14626), .A2(n19941), .B1(n19940), .B2(n14855), .ZN(
        n14630) );
  AOI21_X1 U18092 ( .B1(n14641), .B2(P1_REIP_REG_27__SCAN_IN), .A(
        P1_REIP_REG_28__SCAN_IN), .ZN(n14628) );
  NOR2_X1 U18093 ( .A1(n14628), .A2(n14627), .ZN(n14629) );
  AOI211_X1 U18094 ( .C1(n19938), .C2(P1_EBX_REG_28__SCAN_IN), .A(n14630), .B(
        n14629), .ZN(n14631) );
  OAI211_X1 U18095 ( .C1(n19897), .C2(n14988), .A(n14632), .B(n14631), .ZN(
        P1_U2812) );
  NAND2_X1 U18096 ( .A1(n14649), .A2(n14633), .ZN(n14634) );
  NAND2_X1 U18097 ( .A1(n14635), .A2(n14634), .ZN(n14996) );
  AOI21_X1 U18098 ( .B1(n14637), .B2(n14636), .A(n14623), .ZN(n14866) );
  NAND2_X1 U18099 ( .A1(n14866), .A2(n19904), .ZN(n14646) );
  NOR2_X1 U18100 ( .A1(n14639), .A2(n14638), .ZN(n14654) );
  INV_X1 U18101 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n14640) );
  NAND2_X1 U18102 ( .A1(n14641), .A2(n14640), .ZN(n14643) );
  AOI22_X1 U18103 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19926), .B1(
        n19927), .B2(n14862), .ZN(n14642) );
  OAI211_X1 U18104 ( .C1(n20828), .C2(n19895), .A(n14643), .B(n14642), .ZN(
        n14644) );
  AOI21_X1 U18105 ( .B1(P1_REIP_REG_27__SCAN_IN), .B2(n14654), .A(n14644), 
        .ZN(n14645) );
  OAI211_X1 U18106 ( .C1(n19897), .C2(n14996), .A(n14646), .B(n14645), .ZN(
        P1_U2813) );
  OR2_X1 U18107 ( .A1(n14672), .A2(n14647), .ZN(n14648) );
  NAND2_X1 U18108 ( .A1(n14649), .A2(n14648), .ZN(n16029) );
  INV_X1 U18109 ( .A(n14636), .ZN(n14651) );
  AOI21_X1 U18110 ( .B1(n14652), .B2(n14650), .A(n14651), .ZN(n14874) );
  NAND2_X1 U18111 ( .A1(n14874), .A2(n19904), .ZN(n14661) );
  OAI22_X1 U18112 ( .A1(n14653), .A2(n19941), .B1(n19940), .B2(n14872), .ZN(
        n14659) );
  INV_X1 U18113 ( .A(n14654), .ZN(n14657) );
  AOI21_X1 U18114 ( .B1(n19881), .B2(n14655), .A(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14656) );
  NOR2_X1 U18115 ( .A1(n14657), .A2(n14656), .ZN(n14658) );
  AOI211_X1 U18116 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n19938), .A(n14659), .B(
        n14658), .ZN(n14660) );
  OAI211_X1 U18117 ( .C1(n19897), .C2(n16029), .A(n14661), .B(n14660), .ZN(
        P1_U2814) );
  OAI21_X1 U18118 ( .B1(n14662), .B2(n14663), .A(n14650), .ZN(n14884) );
  NAND2_X1 U18119 ( .A1(n15813), .A2(n15837), .ZN(n14664) );
  AND2_X1 U18120 ( .A1(n19939), .A2(n14664), .ZN(n15826) );
  INV_X1 U18121 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n14667) );
  NAND2_X1 U18122 ( .A1(n14485), .A2(n14665), .ZN(n14666) );
  OAI211_X1 U18123 ( .C1(n14485), .C2(n14667), .A(n19881), .B(n14666), .ZN(
        n14669) );
  AOI22_X1 U18124 ( .A1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n19926), .B1(
        n19927), .B2(n14882), .ZN(n14668) );
  OAI211_X1 U18125 ( .C1(n19895), .C2(n14708), .A(n14669), .B(n14668), .ZN(
        n14674) );
  NOR2_X1 U18126 ( .A1(n14715), .A2(n14670), .ZN(n14671) );
  OR2_X1 U18127 ( .A1(n14672), .A2(n14671), .ZN(n15005) );
  NOR2_X1 U18128 ( .A1(n15005), .A2(n19897), .ZN(n14673) );
  AOI211_X1 U18129 ( .C1(P1_REIP_REG_25__SCAN_IN), .C2(n15826), .A(n14674), 
        .B(n14673), .ZN(n14675) );
  OAI21_X1 U18130 ( .B1(n14884), .B2(n15891), .A(n14675), .ZN(P1_U2815) );
  AOI21_X1 U18131 ( .B1(n14678), .B2(n14677), .A(n14676), .ZN(n14825) );
  INV_X1 U18132 ( .A(n14679), .ZN(n14824) );
  NOR2_X1 U18133 ( .A1(n14825), .A2(n14824), .ZN(n14823) );
  OAI21_X1 U18134 ( .B1(n14823), .B2(n14681), .A(n14680), .ZN(n14952) );
  INV_X1 U18135 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n15901) );
  AOI22_X1 U18136 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n15914), .B1(n15865), 
        .B2(n15901), .ZN(n14690) );
  OAI21_X1 U18137 ( .B1(n15910), .B2(n14683), .A(n14682), .ZN(n14684) );
  INV_X1 U18138 ( .A(n14684), .ZN(n16093) );
  INV_X1 U18139 ( .A(n14948), .ZN(n14685) );
  AOI22_X1 U18140 ( .A1(P1_EBX_REG_13__SCAN_IN), .A2(n19938), .B1(n19927), 
        .B2(n14685), .ZN(n14686) );
  OAI211_X1 U18141 ( .C1(n19941), .C2(n14687), .A(n14686), .B(n15929), .ZN(
        n14688) );
  AOI21_X1 U18142 ( .B1(n16093), .B2(n19945), .A(n14688), .ZN(n14689) );
  OAI211_X1 U18143 ( .C1(n14952), .C2(n15891), .A(n14690), .B(n14689), .ZN(
        P1_U2827) );
  OAI22_X1 U18144 ( .A1(n20800), .A2(n19941), .B1(n14691), .B2(n19940), .ZN(
        n14692) );
  INV_X1 U18145 ( .A(n14692), .ZN(n14693) );
  OAI211_X1 U18146 ( .C1(n14695), .C2(n14694), .A(n14693), .B(n15929), .ZN(
        n14696) );
  AOI221_X1 U18147 ( .B1(P1_REIP_REG_4__SCAN_IN), .B2(n19919), .C1(n14697), 
        .C2(n19919), .A(n14696), .ZN(n14700) );
  AOI22_X1 U18148 ( .A1(n19945), .A2(n14698), .B1(n19938), .B2(
        P1_EBX_REG_4__SCAN_IN), .ZN(n14699) );
  OAI211_X1 U18149 ( .C1(n19949), .C2(n14701), .A(n14700), .B(n14699), .ZN(
        P1_U2836) );
  INV_X1 U18150 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14702) );
  OAI22_X1 U18151 ( .A1(n14703), .A2(n14761), .B1(n15945), .B2(n14702), .ZN(
        P1_U2841) );
  INV_X1 U18152 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14704) );
  OAI222_X1 U18153 ( .A1(n14750), .A2(n14846), .B1(n14704), .B2(n15945), .C1(
        n14975), .C2(n14761), .ZN(P1_U2843) );
  INV_X1 U18154 ( .A(n14857), .ZN(n14782) );
  INV_X1 U18155 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14705) );
  OAI222_X1 U18156 ( .A1(n14750), .A2(n14782), .B1(n14705), .B2(n15945), .C1(
        n14988), .C2(n14761), .ZN(P1_U2844) );
  INV_X1 U18157 ( .A(n14866), .ZN(n14706) );
  OAI222_X1 U18158 ( .A1(n14750), .A2(n14706), .B1(n20828), .B2(n15945), .C1(
        n14996), .C2(n14761), .ZN(P1_U2845) );
  INV_X1 U18159 ( .A(n14874), .ZN(n14789) );
  INV_X1 U18160 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14707) );
  OAI222_X1 U18161 ( .A1(n14750), .A2(n14789), .B1(n14707), .B2(n15945), .C1(
        n16029), .C2(n14761), .ZN(P1_U2846) );
  OAI222_X1 U18162 ( .A1(n15005), .A2(n14761), .B1(n14708), .B2(n15945), .C1(
        n14884), .C2(n14750), .ZN(P1_U2847) );
  OR2_X2 U18163 ( .A1(n15857), .A2(n15858), .ZN(n15855) );
  NOR2_X1 U18164 ( .A1(n15855), .A2(n14710), .ZN(n14718) );
  NOR2_X1 U18165 ( .A1(n14718), .A2(n14711), .ZN(n14712) );
  OR2_X1 U18166 ( .A1(n14662), .A2(n14712), .ZN(n15956) );
  INV_X1 U18167 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14716) );
  NOR2_X1 U18168 ( .A1(n14722), .A2(n14713), .ZN(n14714) );
  OR2_X1 U18169 ( .A1(n14715), .A2(n14714), .ZN(n16038) );
  OAI222_X1 U18170 ( .A1(n14750), .A2(n15956), .B1(n14716), .B2(n15945), .C1(
        n16038), .C2(n14761), .ZN(P1_U2848) );
  INV_X1 U18171 ( .A(n14718), .ZN(n14719) );
  AND2_X1 U18172 ( .A1(n9686), .A2(n14721), .ZN(n14723) );
  OR2_X1 U18173 ( .A1(n14723), .A2(n14722), .ZN(n15834) );
  OAI22_X1 U18174 ( .A1(n15834), .A2(n14761), .B1(n15824), .B2(n15945), .ZN(
        n14724) );
  INV_X1 U18175 ( .A(n14724), .ZN(n14725) );
  OAI21_X1 U18176 ( .B1(n15829), .B2(n14750), .A(n14725), .ZN(P1_U2849) );
  AOI21_X1 U18177 ( .B1(n14727), .B2(n14731), .A(n14726), .ZN(n15964) );
  INV_X1 U18178 ( .A(n15964), .ZN(n14804) );
  NAND2_X1 U18179 ( .A1(n14735), .A2(n14728), .ZN(n14729) );
  AND2_X1 U18180 ( .A1(n9686), .A2(n14729), .ZN(n16053) );
  AOI22_X1 U18181 ( .A1(n16053), .A2(n15941), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n14763), .ZN(n14730) );
  OAI21_X1 U18182 ( .B1(n14804), .B2(n14750), .A(n14730), .ZN(P1_U2850) );
  AOI21_X1 U18183 ( .B1(n14732), .B2(n15855), .A(n9613), .ZN(n14895) );
  INV_X1 U18184 ( .A(n14895), .ZN(n15848) );
  NAND2_X1 U18185 ( .A1(n15797), .A2(n14733), .ZN(n14734) );
  NAND2_X1 U18186 ( .A1(n14735), .A2(n14734), .ZN(n15847) );
  OAI22_X1 U18187 ( .A1(n15847), .A2(n14761), .B1(n15846), .B2(n15945), .ZN(
        n14736) );
  INV_X1 U18188 ( .A(n14736), .ZN(n14737) );
  OAI21_X1 U18189 ( .B1(n15848), .B2(n14750), .A(n14737), .ZN(P1_U2851) );
  OR2_X1 U18190 ( .A1(n14748), .A2(n14738), .ZN(n14739) );
  NAND2_X1 U18191 ( .A1(n15857), .A2(n14739), .ZN(n14904) );
  INV_X1 U18192 ( .A(n14904), .ZN(n15873) );
  OR2_X1 U18193 ( .A1(n9704), .A2(n14740), .ZN(n14741) );
  NAND2_X1 U18194 ( .A1(n15799), .A2(n14741), .ZN(n16060) );
  OAI22_X1 U18195 ( .A1(n16060), .A2(n14761), .B1(n14742), .B2(n15945), .ZN(
        n14743) );
  AOI21_X1 U18196 ( .B1(n15873), .B2(n15942), .A(n14743), .ZN(n14744) );
  INV_X1 U18197 ( .A(n14744), .ZN(P1_U2853) );
  AND2_X1 U18198 ( .A1(n14760), .A2(n14745), .ZN(n14746) );
  OR2_X1 U18199 ( .A1(n9704), .A2(n14746), .ZN(n15880) );
  INV_X1 U18200 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14751) );
  AND2_X1 U18201 ( .A1(n14754), .A2(n14747), .ZN(n14749) );
  OR2_X1 U18202 ( .A1(n14749), .A2(n14748), .ZN(n15881) );
  OAI222_X1 U18203 ( .A1(n15880), .A2(n14761), .B1(n14751), .B2(n15945), .C1(
        n15881), .C2(n14750), .ZN(P1_U2854) );
  INV_X1 U18204 ( .A(n14752), .ZN(n14755) );
  OAI21_X1 U18205 ( .B1(n14755), .B2(n9955), .A(n14754), .ZN(n15892) );
  INV_X1 U18206 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n14762) );
  INV_X1 U18207 ( .A(n14756), .ZN(n14758) );
  NAND2_X1 U18208 ( .A1(n14758), .A2(n9893), .ZN(n14759) );
  NAND2_X1 U18209 ( .A1(n14760), .A2(n14759), .ZN(n15899) );
  OAI222_X1 U18210 ( .A1(n14750), .A2(n15892), .B1(n15945), .B2(n14762), .C1(
        n15899), .C2(n14761), .ZN(P1_U2855) );
  AOI22_X1 U18211 ( .A1(n16093), .A2(n15941), .B1(P1_EBX_REG_13__SCAN_IN), 
        .B2(n14763), .ZN(n14764) );
  OAI21_X1 U18212 ( .B1(n14952), .B2(n14750), .A(n14764), .ZN(P1_U2859) );
  INV_X1 U18213 ( .A(n15948), .ZN(n14792) );
  INV_X1 U18214 ( .A(DATAI_30_), .ZN(n14766) );
  AOI22_X1 U18215 ( .A1(n15947), .A2(n20030), .B1(n15946), .B2(
        P1_EAX_REG_30__SCAN_IN), .ZN(n14765) );
  OAI21_X1 U18216 ( .B1(n14792), .B2(n14766), .A(n14765), .ZN(n14767) );
  AOI21_X1 U18217 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n14819), .A(n14767), .ZN(
        n14768) );
  OAI21_X1 U18218 ( .B1(n14769), .B2(n14828), .A(n14768), .ZN(P1_U2874) );
  INV_X1 U18219 ( .A(DATAI_29_), .ZN(n14773) );
  INV_X1 U18220 ( .A(DATAI_13_), .ZN(n14771) );
  NAND2_X1 U18221 ( .A1(n20099), .A2(BUF1_REG_13__SCAN_IN), .ZN(n14770) );
  OAI21_X1 U18222 ( .B1(n20099), .B2(n14771), .A(n14770), .ZN(n20026) );
  AOI22_X1 U18223 ( .A1(n15947), .A2(n20026), .B1(n15946), .B2(
        P1_EAX_REG_29__SCAN_IN), .ZN(n14772) );
  OAI21_X1 U18224 ( .B1(n14792), .B2(n14773), .A(n14772), .ZN(n14774) );
  AOI21_X1 U18225 ( .B1(BUF1_REG_29__SCAN_IN), .B2(n14819), .A(n14774), .ZN(
        n14775) );
  OAI21_X1 U18226 ( .B1(n14846), .B2(n14828), .A(n14775), .ZN(P1_U2875) );
  INV_X1 U18227 ( .A(DATAI_28_), .ZN(n14779) );
  INV_X1 U18228 ( .A(DATAI_12_), .ZN(n14777) );
  NAND2_X1 U18229 ( .A1(n20099), .A2(BUF1_REG_12__SCAN_IN), .ZN(n14776) );
  OAI21_X1 U18230 ( .B1(n20099), .B2(n14777), .A(n14776), .ZN(n20022) );
  AOI22_X1 U18231 ( .A1(n15947), .A2(n20022), .B1(n15946), .B2(
        P1_EAX_REG_28__SCAN_IN), .ZN(n14778) );
  OAI21_X1 U18232 ( .B1(n14792), .B2(n14779), .A(n14778), .ZN(n14780) );
  AOI21_X1 U18233 ( .B1(BUF1_REG_28__SCAN_IN), .B2(n14819), .A(n14780), .ZN(
        n14781) );
  OAI21_X1 U18234 ( .B1(n14782), .B2(n14828), .A(n14781), .ZN(P1_U2876) );
  INV_X1 U18235 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n15183) );
  NAND2_X1 U18236 ( .A1(n14866), .A2(n15949), .ZN(n14785) );
  OAI22_X1 U18237 ( .A1(n14817), .A2(n20017), .B1(n20021), .B2(n14815), .ZN(
        n14783) );
  AOI21_X1 U18238 ( .B1(n15948), .B2(DATAI_27_), .A(n14783), .ZN(n14784) );
  OAI211_X1 U18239 ( .C1(n15952), .C2(n15183), .A(n14785), .B(n14784), .ZN(
        P1_U2877) );
  OAI22_X1 U18240 ( .A1(n14817), .A2(n20012), .B1(n20016), .B2(n14815), .ZN(
        n14786) );
  AOI21_X1 U18241 ( .B1(n15948), .B2(DATAI_26_), .A(n14786), .ZN(n14788) );
  NAND2_X1 U18242 ( .A1(n14819), .A2(BUF1_REG_26__SCAN_IN), .ZN(n14787) );
  OAI211_X1 U18243 ( .C1(n14789), .C2(n14828), .A(n14788), .B(n14787), .ZN(
        P1_U2878) );
  INV_X1 U18244 ( .A(DATAI_25_), .ZN(n14791) );
  AOI22_X1 U18245 ( .A1(n15947), .A2(n20008), .B1(n15946), .B2(
        P1_EAX_REG_25__SCAN_IN), .ZN(n14790) );
  OAI21_X1 U18246 ( .B1(n14792), .B2(n14791), .A(n14790), .ZN(n14793) );
  AOI21_X1 U18247 ( .B1(n14819), .B2(BUF1_REG_25__SCAN_IN), .A(n14793), .ZN(
        n14794) );
  OAI21_X1 U18248 ( .B1(n14884), .B2(n14828), .A(n14794), .ZN(P1_U2879) );
  OAI22_X1 U18249 ( .A1(n14817), .A2(n20003), .B1(n20007), .B2(n14815), .ZN(
        n14795) );
  AOI21_X1 U18250 ( .B1(n15948), .B2(DATAI_24_), .A(n14795), .ZN(n14797) );
  NAND2_X1 U18251 ( .A1(n14819), .A2(BUF1_REG_24__SCAN_IN), .ZN(n14796) );
  OAI211_X1 U18252 ( .C1(n15956), .C2(n14814), .A(n14797), .B(n14796), .ZN(
        P1_U2880) );
  OAI22_X1 U18253 ( .A1(n14817), .A2(n20144), .B1(n20807), .B2(n14815), .ZN(
        n14798) );
  AOI21_X1 U18254 ( .B1(n15948), .B2(DATAI_23_), .A(n14798), .ZN(n14800) );
  NAND2_X1 U18255 ( .A1(n14819), .A2(BUF1_REG_23__SCAN_IN), .ZN(n14799) );
  OAI211_X1 U18256 ( .C1(n15829), .C2(n14828), .A(n14800), .B(n14799), .ZN(
        P1_U2881) );
  OAI22_X1 U18257 ( .A1(n14817), .A2(n20137), .B1(n19999), .B2(n14815), .ZN(
        n14801) );
  AOI21_X1 U18258 ( .B1(n15948), .B2(DATAI_22_), .A(n14801), .ZN(n14803) );
  NAND2_X1 U18259 ( .A1(n14819), .A2(BUF1_REG_22__SCAN_IN), .ZN(n14802) );
  OAI211_X1 U18260 ( .C1(n14804), .C2(n14814), .A(n14803), .B(n14802), .ZN(
        P1_U2882) );
  OAI22_X1 U18261 ( .A1(n14817), .A2(n20134), .B1(n19995), .B2(n14815), .ZN(
        n14805) );
  AOI21_X1 U18262 ( .B1(n15948), .B2(DATAI_21_), .A(n14805), .ZN(n14807) );
  NAND2_X1 U18263 ( .A1(n14819), .A2(BUF1_REG_21__SCAN_IN), .ZN(n14806) );
  OAI211_X1 U18264 ( .C1(n15848), .C2(n14814), .A(n14807), .B(n14806), .ZN(
        P1_U2883) );
  OAI22_X1 U18265 ( .A1(n14817), .A2(n20128), .B1(n19987), .B2(n14815), .ZN(
        n14808) );
  AOI21_X1 U18266 ( .B1(n15948), .B2(DATAI_19_), .A(n14808), .ZN(n14810) );
  NAND2_X1 U18267 ( .A1(n14819), .A2(BUF1_REG_19__SCAN_IN), .ZN(n14809) );
  OAI211_X1 U18268 ( .C1(n14904), .C2(n14814), .A(n14810), .B(n14809), .ZN(
        P1_U2885) );
  OAI22_X1 U18269 ( .A1(n14817), .A2(n20124), .B1(n19983), .B2(n14815), .ZN(
        n14811) );
  AOI21_X1 U18270 ( .B1(n15948), .B2(DATAI_18_), .A(n14811), .ZN(n14813) );
  NAND2_X1 U18271 ( .A1(n14819), .A2(BUF1_REG_18__SCAN_IN), .ZN(n14812) );
  OAI211_X1 U18272 ( .C1(n15881), .C2(n14814), .A(n14813), .B(n14812), .ZN(
        P1_U2886) );
  OAI22_X1 U18273 ( .A1(n14817), .A2(n20121), .B1(n14816), .B2(n14815), .ZN(
        n14818) );
  AOI21_X1 U18274 ( .B1(n15948), .B2(DATAI_17_), .A(n14818), .ZN(n14821) );
  NAND2_X1 U18275 ( .A1(n14819), .A2(BUF1_REG_17__SCAN_IN), .ZN(n14820) );
  OAI211_X1 U18276 ( .C1(n15892), .C2(n14828), .A(n14821), .B(n14820), .ZN(
        P1_U2887) );
  AOI22_X1 U18277 ( .A1(n14826), .A2(n20026), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n15946), .ZN(n14822) );
  OAI21_X1 U18278 ( .B1(n14952), .B2(n14828), .A(n14822), .ZN(P1_U2891) );
  AOI21_X1 U18279 ( .B1(n14825), .B2(n14824), .A(n14823), .ZN(n15998) );
  INV_X1 U18280 ( .A(n15998), .ZN(n14829) );
  AOI22_X1 U18281 ( .A1(n14826), .A2(n20022), .B1(P1_EAX_REG_12__SCAN_IN), 
        .B2(n15946), .ZN(n14827) );
  OAI21_X1 U18282 ( .B1(n14829), .B2(n14828), .A(n14827), .ZN(P1_U2892) );
  AOI21_X1 U18283 ( .B1(n14831), .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n14830), .ZN(n14969) );
  NAND2_X1 U18284 ( .A1(n16052), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14965) );
  NAND2_X1 U18285 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14832) );
  OAI211_X1 U18286 ( .C1(n16019), .C2(n14833), .A(n14965), .B(n14832), .ZN(
        n14834) );
  AOI21_X1 U18287 ( .B1(n14835), .B2(n16022), .A(n14834), .ZN(n14836) );
  OAI21_X1 U18288 ( .B1(n14969), .B2(n19850), .A(n14836), .ZN(P1_U2969) );
  NAND2_X1 U18289 ( .A1(n16052), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14974) );
  OAI21_X1 U18290 ( .B1(n16026), .B2(n14837), .A(n14974), .ZN(n14838) );
  AOI21_X1 U18291 ( .B1(n14839), .B2(n16021), .A(n14838), .ZN(n14845) );
  NAND2_X1 U18292 ( .A1(n14840), .A2(n14983), .ZN(n14842) );
  NAND2_X1 U18293 ( .A1(n14859), .A2(n14982), .ZN(n14841) );
  XNOR2_X2 U18294 ( .A(n14843), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14970) );
  NAND2_X1 U18295 ( .A1(n14970), .A2(n20093), .ZN(n14844) );
  OAI211_X1 U18296 ( .C1(n14846), .C2(n20102), .A(n14845), .B(n14844), .ZN(
        P1_U2970) );
  NAND2_X1 U18297 ( .A1(n15987), .A2(n14848), .ZN(n14868) );
  NAND2_X1 U18298 ( .A1(n14847), .A2(n14868), .ZN(n14852) );
  OAI21_X1 U18299 ( .B1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n14849), .A(
        n14852), .ZN(n14851) );
  MUX2_X1 U18300 ( .A(n14992), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .S(
        n15987), .Z(n14850) );
  OAI211_X1 U18301 ( .C1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n14852), .A(
        n14851), .B(n14850), .ZN(n14853) );
  XOR2_X1 U18302 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n14853), .Z(
        n14991) );
  NAND2_X1 U18303 ( .A1(n16052), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14984) );
  NAND2_X1 U18304 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14854) );
  OAI211_X1 U18305 ( .C1(n16019), .C2(n14855), .A(n14984), .B(n14854), .ZN(
        n14856) );
  AOI21_X1 U18306 ( .B1(n14857), .B2(n16022), .A(n14856), .ZN(n14858) );
  OAI21_X1 U18307 ( .B1(n19850), .B2(n14991), .A(n14858), .ZN(P1_U2971) );
  MUX2_X1 U18308 ( .A(n14860), .B(n14859), .S(n10059), .Z(n14861) );
  XNOR2_X1 U18309 ( .A(n14861), .B(n14992), .ZN(n15000) );
  NAND2_X1 U18310 ( .A1(n16021), .A2(n14862), .ZN(n14863) );
  NAND2_X1 U18311 ( .A1(n16052), .A2(P1_REIP_REG_27__SCAN_IN), .ZN(n14995) );
  OAI211_X1 U18312 ( .C1(n16026), .C2(n14864), .A(n14863), .B(n14995), .ZN(
        n14865) );
  AOI21_X1 U18313 ( .B1(n14866), .B2(n16022), .A(n14865), .ZN(n14867) );
  OAI21_X1 U18314 ( .B1(n19850), .B2(n15000), .A(n14867), .ZN(P1_U2972) );
  OAI211_X1 U18315 ( .C1(n10059), .C2(n14847), .A(n14869), .B(n14868), .ZN(
        n14870) );
  XOR2_X1 U18316 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n14870), .Z(
        n16028) );
  AOI22_X1 U18317 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n16141), .B2(P1_REIP_REG_26__SCAN_IN), .ZN(n14871) );
  OAI21_X1 U18318 ( .B1(n16019), .B2(n14872), .A(n14871), .ZN(n14873) );
  AOI21_X1 U18319 ( .B1(n14874), .B2(n16022), .A(n14873), .ZN(n14875) );
  OAI21_X1 U18320 ( .B1(n19850), .B2(n16028), .A(n14875), .ZN(P1_U2973) );
  INV_X1 U18321 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14881) );
  NAND2_X1 U18322 ( .A1(n16141), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n15001) );
  NOR2_X1 U18323 ( .A1(n14877), .A2(n15954), .ZN(n14879) );
  NOR3_X1 U18324 ( .A1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n14847), .ZN(n14878) );
  MUX2_X1 U18325 ( .A(n14879), .B(n14878), .S(n10059), .Z(n14880) );
  OAI21_X1 U18326 ( .B1(n14884), .B2(n20102), .A(n14883), .ZN(P1_U2974) );
  XNOR2_X1 U18327 ( .A(n9626), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14885) );
  XNOR2_X1 U18328 ( .A(n14847), .B(n14885), .ZN(n15016) );
  OAI22_X1 U18329 ( .A1(n16026), .A2(n15823), .B1(n16103), .B2(n14484), .ZN(
        n14887) );
  NOR2_X1 U18330 ( .A1(n15829), .A2(n20102), .ZN(n14886) );
  AOI211_X1 U18331 ( .C1(n16021), .C2(n15832), .A(n14887), .B(n14886), .ZN(
        n14888) );
  OAI21_X1 U18332 ( .B1(n15016), .B2(n19850), .A(n14888), .ZN(P1_U2976) );
  NAND2_X1 U18333 ( .A1(n14889), .A2(n10059), .ZN(n15791) );
  NAND3_X1 U18334 ( .A1(n14890), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n9626), .ZN(n15790) );
  OAI22_X1 U18335 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15791), .B1(
        n15790), .B2(n14891), .ZN(n14892) );
  XNOR2_X1 U18336 ( .A(n14892), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15030) );
  NAND2_X1 U18337 ( .A1(n16021), .A2(n15844), .ZN(n14893) );
  NAND2_X1 U18338 ( .A1(n16141), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n15026) );
  OAI211_X1 U18339 ( .C1(n16026), .C2(n15845), .A(n14893), .B(n15026), .ZN(
        n14894) );
  AOI21_X1 U18340 ( .B1(n14895), .B2(n16022), .A(n14894), .ZN(n14896) );
  OAI21_X1 U18341 ( .B1(n15030), .B2(n19850), .A(n14896), .ZN(P1_U2978) );
  NOR2_X1 U18342 ( .A1(n14890), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14897) );
  MUX2_X1 U18343 ( .A(n14897), .B(n14890), .S(n9626), .Z(n14898) );
  XNOR2_X1 U18344 ( .A(n14898), .B(n16065), .ZN(n16062) );
  NAND2_X1 U18345 ( .A1(n16062), .A2(n20093), .ZN(n14903) );
  INV_X1 U18346 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n14899) );
  OAI22_X1 U18347 ( .A1(n16026), .A2(n14900), .B1(n16103), .B2(n14899), .ZN(
        n14901) );
  AOI21_X1 U18348 ( .B1(n16021), .B2(n15867), .A(n14901), .ZN(n14902) );
  OAI211_X1 U18349 ( .C1(n20102), .C2(n14904), .A(n14903), .B(n14902), .ZN(
        P1_U2980) );
  INV_X1 U18350 ( .A(n14890), .ZN(n14905) );
  OAI21_X1 U18351 ( .B1(n14907), .B2(n14906), .A(n14905), .ZN(n15041) );
  NAND2_X1 U18352 ( .A1(n16141), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n15036) );
  OAI21_X1 U18353 ( .B1(n16026), .B2(n14908), .A(n15036), .ZN(n14910) );
  NOR2_X1 U18354 ( .A1(n15881), .A2(n20102), .ZN(n14909) );
  AOI211_X1 U18355 ( .C1(n16021), .C2(n15886), .A(n14910), .B(n14909), .ZN(
        n14911) );
  OAI21_X1 U18356 ( .B1(n19850), .B2(n15041), .A(n14911), .ZN(P1_U2981) );
  INV_X1 U18357 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15043) );
  INV_X1 U18358 ( .A(n14912), .ZN(n14913) );
  NAND2_X1 U18359 ( .A1(n14940), .A2(n14913), .ZN(n14915) );
  NAND2_X1 U18360 ( .A1(n14915), .A2(n14914), .ZN(n15986) );
  AND2_X1 U18361 ( .A1(n15987), .A2(n14916), .ZN(n14917) );
  INV_X1 U18362 ( .A(n14918), .ZN(n14919) );
  OR2_X1 U18363 ( .A1(n15987), .A2(n14921), .ZN(n14932) );
  NAND2_X1 U18364 ( .A1(n14933), .A2(n14932), .ZN(n15974) );
  INV_X1 U18365 ( .A(n15974), .ZN(n14925) );
  NAND2_X1 U18366 ( .A1(n15974), .A2(n14922), .ZN(n15978) );
  INV_X1 U18367 ( .A(n15978), .ZN(n14924) );
  MUX2_X1 U18368 ( .A(n14925), .B(n14924), .S(n14923), .Z(n14926) );
  INV_X1 U18369 ( .A(n15890), .ZN(n14930) );
  NAND2_X1 U18370 ( .A1(n16052), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n15044) );
  OAI21_X1 U18371 ( .B1(n16026), .B2(n14927), .A(n15044), .ZN(n14929) );
  NOR2_X1 U18372 ( .A1(n15892), .A2(n20102), .ZN(n14928) );
  AOI211_X1 U18373 ( .C1(n16021), .C2(n14930), .A(n14929), .B(n14928), .ZN(
        n14931) );
  OAI21_X1 U18374 ( .B1(n10061), .B2(n19850), .A(n14931), .ZN(P1_U2982) );
  NAND2_X1 U18375 ( .A1(n14932), .A2(n15973), .ZN(n14934) );
  XOR2_X1 U18376 ( .A(n14934), .B(n14933), .Z(n16077) );
  NAND2_X1 U18377 ( .A1(n16077), .A2(n20093), .ZN(n14938) );
  AND2_X1 U18378 ( .A1(n16141), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n16075) );
  NOR2_X1 U18379 ( .A1(n16019), .A2(n14935), .ZN(n14936) );
  AOI211_X1 U18380 ( .C1(n20091), .C2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n16075), .B(n14936), .ZN(n14937) );
  OAI211_X1 U18381 ( .C1(n20102), .C2(n14939), .A(n14938), .B(n14937), .ZN(
        P1_U2984) );
  INV_X1 U18382 ( .A(n14940), .ZN(n15049) );
  INV_X1 U18383 ( .A(n14941), .ZN(n14942) );
  AOI22_X1 U18384 ( .A1(n15049), .A2(n14943), .B1(n10059), .B2(n14942), .ZN(
        n15996) );
  INV_X1 U18385 ( .A(n14945), .ZN(n14944) );
  AOI21_X1 U18386 ( .B1(n10059), .B2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n14944), .ZN(n15995) );
  NAND2_X1 U18387 ( .A1(n15996), .A2(n15995), .ZN(n15994) );
  NAND2_X1 U18388 ( .A1(n15994), .A2(n14945), .ZN(n14946) );
  XOR2_X1 U18389 ( .A(n14947), .B(n14946), .Z(n16095) );
  NAND2_X1 U18390 ( .A1(n16095), .A2(n20093), .ZN(n14951) );
  AND2_X1 U18391 ( .A1(n16141), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n16092) );
  NOR2_X1 U18392 ( .A1(n16019), .A2(n14948), .ZN(n14949) );
  AOI211_X1 U18393 ( .C1(n20091), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n16092), .B(n14949), .ZN(n14950) );
  OAI211_X1 U18394 ( .C1(n20102), .C2(n14952), .A(n14951), .B(n14950), .ZN(
        P1_U2986) );
  NAND2_X1 U18395 ( .A1(n16052), .A2(P1_REIP_REG_10__SCAN_IN), .ZN(n16113) );
  INV_X1 U18396 ( .A(n14953), .ZN(n14954) );
  MUX2_X1 U18397 ( .A(n14954), .B(n15049), .S(n9626), .Z(n14955) );
  XOR2_X1 U18398 ( .A(n14955), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .Z(
        n16116) );
  NAND2_X1 U18399 ( .A1(n20093), .A2(n16116), .ZN(n14956) );
  OAI211_X1 U18400 ( .C1(n16026), .C2(n14957), .A(n16113), .B(n14956), .ZN(
        n14958) );
  AOI21_X1 U18401 ( .B1(n15926), .B2(n16021), .A(n14958), .ZN(n14959) );
  OAI21_X1 U18402 ( .B1(n14960), .B2(n20102), .A(n14959), .ZN(P1_U2989) );
  INV_X1 U18403 ( .A(n14961), .ZN(n14963) );
  OAI21_X1 U18404 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14963), .A(
        n14962), .ZN(n14964) );
  OAI211_X1 U18405 ( .C1(n14966), .C2(n16068), .A(n14965), .B(n14964), .ZN(
        n14967) );
  INV_X1 U18406 ( .A(n14967), .ZN(n14968) );
  OAI21_X1 U18407 ( .B1(n14969), .B2(n16111), .A(n14968), .ZN(P1_U3001) );
  INV_X1 U18408 ( .A(n14970), .ZN(n14979) );
  INV_X1 U18409 ( .A(n14971), .ZN(n14977) );
  INV_X1 U18410 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14972) );
  NAND3_X1 U18411 ( .A1(n14993), .A2(n14982), .A3(n14972), .ZN(n14973) );
  OAI211_X1 U18412 ( .C1(n14975), .C2(n16068), .A(n14974), .B(n14973), .ZN(
        n14976) );
  AOI21_X1 U18413 ( .B1(n14977), .B2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n14976), .ZN(n14978) );
  OAI21_X1 U18414 ( .B1(n14979), .B2(n16111), .A(n14978), .ZN(P1_U3002) );
  AND2_X1 U18415 ( .A1(n14981), .A2(n14980), .ZN(n14998) );
  NOR2_X1 U18416 ( .A1(n14983), .A2(n14982), .ZN(n14986) );
  INV_X1 U18417 ( .A(n14984), .ZN(n14985) );
  AOI21_X1 U18418 ( .B1(n14993), .B2(n14986), .A(n14985), .ZN(n14987) );
  OAI21_X1 U18419 ( .B1(n14988), .B2(n16068), .A(n14987), .ZN(n14989) );
  AOI21_X1 U18420 ( .B1(n14998), .B2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        n14989), .ZN(n14990) );
  OAI21_X1 U18421 ( .B1(n14991), .B2(n16111), .A(n14990), .ZN(P1_U3003) );
  NAND2_X1 U18422 ( .A1(n14993), .A2(n14992), .ZN(n14994) );
  OAI211_X1 U18423 ( .C1(n14996), .C2(n16068), .A(n14995), .B(n14994), .ZN(
        n14997) );
  AOI21_X1 U18424 ( .B1(n14998), .B2(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n14997), .ZN(n14999) );
  OAI21_X1 U18425 ( .B1(n15000), .B2(n16111), .A(n14999), .ZN(P1_U3004) );
  INV_X1 U18426 ( .A(n15001), .ZN(n15003) );
  NOR3_X1 U18427 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n15002), .A3(
        n16044), .ZN(n16033) );
  AOI211_X1 U18428 ( .C1(n16144), .C2(n15004), .A(n15003), .B(n16033), .ZN(
        n15008) );
  INV_X1 U18429 ( .A(n15005), .ZN(n15006) );
  NAND2_X1 U18430 ( .A1(n15006), .A2(n16142), .ZN(n15007) );
  OAI211_X1 U18431 ( .C1(n15010), .C2(n15009), .A(n15008), .B(n15007), .ZN(
        P1_U3006) );
  INV_X1 U18432 ( .A(n15834), .ZN(n15014) );
  NAND2_X1 U18433 ( .A1(n16052), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n15011) );
  OAI221_X1 U18434 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n16044), 
        .C1(n16045), .C2(n15012), .A(n15011), .ZN(n15013) );
  AOI21_X1 U18435 ( .B1(n15014), .B2(n16142), .A(n15013), .ZN(n15015) );
  OAI21_X1 U18436 ( .B1(n15016), .B2(n16111), .A(n15015), .ZN(P1_U3008) );
  INV_X1 U18437 ( .A(n15017), .ZN(n15023) );
  NOR3_X1 U18438 ( .A1(n15019), .A2(n15022), .A3(n15018), .ZN(n15020) );
  AOI21_X1 U18439 ( .B1(n15021), .B2(n15061), .A(n15020), .ZN(n15795) );
  OAI21_X1 U18440 ( .B1(n15794), .B2(n15022), .A(n15795), .ZN(n16094) );
  NAND2_X1 U18441 ( .A1(n15023), .A2(n16094), .ZN(n16066) );
  NOR2_X1 U18442 ( .A1(n15024), .A2(n16066), .ZN(n16055) );
  NAND2_X1 U18443 ( .A1(n16055), .A2(n15025), .ZN(n15027) );
  OAI211_X1 U18444 ( .C1(n16068), .C2(n15847), .A(n15027), .B(n15026), .ZN(
        n15028) );
  AOI21_X1 U18445 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n16051), .A(
        n15028), .ZN(n15029) );
  OAI21_X1 U18446 ( .B1(n15030), .B2(n16111), .A(n15029), .ZN(P1_U3010) );
  NOR2_X1 U18447 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n15031), .ZN(
        n15039) );
  INV_X1 U18448 ( .A(n15031), .ZN(n15035) );
  OAI22_X1 U18449 ( .A1(n15057), .A2(n15033), .B1(n15032), .B2(n15055), .ZN(
        n15034) );
  NOR2_X1 U18450 ( .A1(n15059), .A2(n15034), .ZN(n16099) );
  OAI21_X1 U18451 ( .B1(n16131), .B2(n15035), .A(n16099), .ZN(n15046) );
  NAND2_X1 U18452 ( .A1(n15046), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15037) );
  OAI211_X1 U18453 ( .C1(n16068), .C2(n15880), .A(n15037), .B(n15036), .ZN(
        n15038) );
  AOI21_X1 U18454 ( .B1(n15039), .B2(n15042), .A(n15038), .ZN(n15040) );
  OAI21_X1 U18455 ( .B1(n15041), .B2(n16111), .A(n15040), .ZN(P1_U3013) );
  NAND2_X1 U18456 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16067) );
  NAND2_X1 U18457 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n15042), .ZN(
        n16081) );
  OAI21_X1 U18458 ( .B1(n16067), .B2(n16081), .A(n15043), .ZN(n15047) );
  OAI21_X1 U18459 ( .B1(n15899), .B2(n16068), .A(n15044), .ZN(n15045) );
  AOI21_X1 U18460 ( .B1(n15047), .B2(n15046), .A(n15045), .ZN(n15048) );
  OAI21_X1 U18461 ( .B1(n10061), .B2(n16111), .A(n15048), .ZN(P1_U3014) );
  NAND2_X1 U18462 ( .A1(n15987), .A2(n15049), .ZN(n15051) );
  NAND2_X1 U18463 ( .A1(n10059), .A2(n16120), .ZN(n15050) );
  OAI22_X1 U18464 ( .A1(n15051), .A2(n16120), .B1(n14953), .B2(n15050), .ZN(
        n15052) );
  XNOR2_X1 U18465 ( .A(n14290), .B(n15052), .ZN(n16003) );
  NOR2_X1 U18466 ( .A1(n16083), .A2(n15053), .ZN(n15063) );
  NOR2_X1 U18467 ( .A1(n14290), .A2(n15054), .ZN(n16108) );
  OAI22_X1 U18468 ( .A1(n15057), .A2(n15056), .B1(n16108), .B2(n15055), .ZN(
        n15058) );
  AOI211_X1 U18469 ( .C1(n15061), .C2(n15060), .A(n15059), .B(n15058), .ZN(
        n16100) );
  INV_X1 U18470 ( .A(n16100), .ZN(n15062) );
  MUX2_X1 U18471 ( .A(n15063), .B(n15062), .S(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(n15066) );
  INV_X1 U18472 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n15064) );
  OAI22_X1 U18473 ( .A1(n15922), .A2(n16068), .B1(n16103), .B2(n15064), .ZN(
        n15065) );
  AOI211_X1 U18474 ( .C1(n16003), .C2(n16144), .A(n15066), .B(n15065), .ZN(
        n15067) );
  INV_X1 U18475 ( .A(n15067), .ZN(P1_U3020) );
  NAND2_X1 U18476 ( .A1(n9593), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20727) );
  OAI211_X1 U18477 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n9593), .A(n20727), 
        .B(n20602), .ZN(n15069) );
  OAI21_X1 U18478 ( .B1(n15071), .B2(n13348), .A(n15069), .ZN(n15070) );
  MUX2_X1 U18479 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n15070), .S(
        n20736), .Z(P1_U3477) );
  XNOR2_X1 U18480 ( .A(n9620), .B(n20727), .ZN(n15072) );
  OAI22_X1 U18481 ( .A1(n15072), .A2(n20728), .B1(n15071), .B2(n20491), .ZN(
        n15073) );
  MUX2_X1 U18482 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n15073), .S(
        n20736), .Z(P1_U3476) );
  NOR2_X1 U18483 ( .A1(n15075), .A2(n15076), .ZN(n15077) );
  OR2_X1 U18484 ( .A1(n15074), .A2(n15077), .ZN(n15440) );
  OR2_X1 U18485 ( .A1(n15458), .A2(n15079), .ZN(n15080) );
  NAND2_X1 U18486 ( .A1(n15078), .A2(n15080), .ZN(n15446) );
  AOI22_X1 U18487 ( .A1(n15081), .A2(n19022), .B1(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n18997), .ZN(n15083) );
  AOI22_X1 U18488 ( .A1(P2_EBX_REG_25__SCAN_IN), .A2(n19018), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n19017), .ZN(n15082) );
  OAI211_X1 U18489 ( .C1(n15446), .C2(n19001), .A(n15083), .B(n15082), .ZN(
        n15087) );
  AOI211_X1 U18490 ( .C1(n9698), .C2(n15085), .A(n15084), .B(n19677), .ZN(
        n15086) );
  NOR2_X1 U18491 ( .A1(n15087), .A2(n15086), .ZN(n15088) );
  OAI21_X1 U18492 ( .B1(n19004), .B2(n15440), .A(n15088), .ZN(P2_U2830) );
  NAND2_X1 U18493 ( .A1(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n18997), .ZN(
        n15089) );
  OAI211_X1 U18494 ( .C1(n18978), .C2(n15090), .A(n19155), .B(n15089), .ZN(
        n15092) );
  NOR2_X1 U18495 ( .A1(n19001), .A2(n15515), .ZN(n15091) );
  AOI211_X1 U18496 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n19018), .A(n15092), .B(
        n15091), .ZN(n15093) );
  OAI21_X1 U18497 ( .B1(n15516), .B2(n19004), .A(n15093), .ZN(n15097) );
  AOI211_X1 U18498 ( .C1(n15312), .C2(n15095), .A(n15094), .B(n19677), .ZN(
        n15096) );
  AOI211_X1 U18499 ( .C1(n19022), .C2(n15098), .A(n15097), .B(n15096), .ZN(
        n15099) );
  INV_X1 U18500 ( .A(n15099), .ZN(P2_U2836) );
  AOI21_X1 U18501 ( .B1(n15102), .B2(n15101), .A(n15100), .ZN(n16227) );
  NAND2_X1 U18502 ( .A1(n19017), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n15103) );
  OAI211_X1 U18503 ( .C1(n19028), .C2(n15324), .A(n15103), .B(n19155), .ZN(
        n15105) );
  NOR2_X1 U18504 ( .A1(n15325), .A2(n19004), .ZN(n15104) );
  AOI211_X1 U18505 ( .C1(P2_EBX_REG_18__SCAN_IN), .C2(n19018), .A(n15105), .B(
        n15104), .ZN(n15106) );
  OAI21_X1 U18506 ( .B1(n18984), .B2(n15107), .A(n15106), .ZN(n15112) );
  AOI211_X1 U18507 ( .C1(n15110), .C2(n15109), .A(n15108), .B(n19677), .ZN(
        n15111) );
  AOI211_X1 U18508 ( .C1(n19016), .C2(n16227), .A(n15112), .B(n15111), .ZN(
        n15113) );
  INV_X1 U18509 ( .A(n15113), .ZN(P2_U2837) );
  INV_X1 U18510 ( .A(n14569), .ZN(n15115) );
  NAND3_X1 U18511 ( .A1(n15115), .A2(n15150), .A3(n15114), .ZN(n15117) );
  NAND2_X1 U18512 ( .A1(n15169), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n15116) );
  OAI211_X1 U18513 ( .C1(n15410), .C2(n15169), .A(n15117), .B(n15116), .ZN(
        P2_U2858) );
  NAND2_X1 U18514 ( .A1(n15119), .A2(n15118), .ZN(n15121) );
  XNOR2_X1 U18515 ( .A(n15121), .B(n15120), .ZN(n15180) );
  NOR2_X1 U18516 ( .A1(n16181), .A2(n15169), .ZN(n15122) );
  AOI21_X1 U18517 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n15169), .A(n15122), .ZN(
        n15123) );
  OAI21_X1 U18518 ( .B1(n15180), .B2(n15124), .A(n15123), .ZN(P2_U2859) );
  AOI21_X1 U18519 ( .B1(n15127), .B2(n15126), .A(n15125), .ZN(n15128) );
  INV_X1 U18520 ( .A(n15128), .ZN(n15188) );
  NAND2_X1 U18521 ( .A1(n15169), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n15130) );
  NAND2_X1 U18522 ( .A1(n15424), .A2(n15157), .ZN(n15129) );
  OAI211_X1 U18523 ( .C1(n15188), .C2(n15124), .A(n15130), .B(n15129), .ZN(
        P2_U2860) );
  INV_X1 U18524 ( .A(n15131), .ZN(n15132) );
  AOI21_X1 U18525 ( .B1(n15134), .B2(n15133), .A(n15132), .ZN(n15189) );
  NAND2_X1 U18526 ( .A1(n15189), .A2(n15150), .ZN(n15139) );
  OR2_X1 U18527 ( .A1(n15074), .A2(n15135), .ZN(n15136) );
  AND2_X1 U18528 ( .A1(n15137), .A2(n15136), .ZN(n16193) );
  NAND2_X1 U18529 ( .A1(n16193), .A2(n15157), .ZN(n15138) );
  OAI211_X1 U18530 ( .C1(n15157), .C2(n15140), .A(n15139), .B(n15138), .ZN(
        P2_U2861) );
  OAI21_X1 U18531 ( .B1(n15143), .B2(n15142), .A(n15141), .ZN(n15204) );
  MUX2_X1 U18532 ( .A(n15440), .B(n10607), .S(n15169), .Z(n15144) );
  OAI21_X1 U18533 ( .B1(n15204), .B2(n15124), .A(n15144), .ZN(P2_U2862) );
  INV_X1 U18534 ( .A(P2_EBX_REG_24__SCAN_IN), .ZN(n15156) );
  OAI21_X1 U18535 ( .B1(n15147), .B2(n15146), .A(n15145), .ZN(n15149) );
  XNOR2_X1 U18536 ( .A(n15149), .B(n15148), .ZN(n16215) );
  NAND2_X1 U18537 ( .A1(n16215), .A2(n15150), .ZN(n15155) );
  AND2_X1 U18538 ( .A1(n15152), .A2(n15151), .ZN(n15153) );
  OR2_X1 U18539 ( .A1(n15153), .A2(n15075), .ZN(n16203) );
  NAND2_X1 U18540 ( .A1(n15466), .A2(n15157), .ZN(n15154) );
  OAI211_X1 U18541 ( .C1(n15157), .C2(n15156), .A(n15155), .B(n15154), .ZN(
        P2_U2863) );
  OAI21_X1 U18542 ( .B1(n15160), .B2(n15159), .A(n15158), .ZN(n15215) );
  NOR2_X1 U18543 ( .A1(n15470), .A2(n15169), .ZN(n15161) );
  AOI21_X1 U18544 ( .B1(P2_EBX_REG_23__SCAN_IN), .B2(n15169), .A(n15161), .ZN(
        n15162) );
  OAI21_X1 U18545 ( .B1(n15215), .B2(n15124), .A(n15162), .ZN(P2_U2864) );
  INV_X1 U18546 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15163) );
  MUX2_X1 U18547 ( .A(n15485), .B(n15163), .S(n15169), .Z(n15164) );
  OAI21_X1 U18548 ( .B1(n15165), .B2(n15124), .A(n15164), .ZN(P2_U2865) );
  NOR2_X1 U18549 ( .A1(n11119), .A2(n15166), .ZN(n15167) );
  OR2_X1 U18550 ( .A1(n15168), .A2(n15167), .ZN(n18859) );
  MUX2_X1 U18551 ( .A(n18859), .B(n10810), .S(n15169), .Z(n15170) );
  OAI21_X1 U18552 ( .B1(n15171), .B2(n15124), .A(n15170), .ZN(P2_U2866) );
  INV_X1 U18553 ( .A(n15172), .ZN(n15173) );
  AOI22_X1 U18554 ( .A1(n15173), .A2(n19099), .B1(n19039), .B2(
        BUF1_REG_31__SCAN_IN), .ZN(n15175) );
  AOI22_X1 U18555 ( .A1(n19038), .A2(BUF2_REG_31__SCAN_IN), .B1(n19098), .B2(
        P2_EAX_REG_31__SCAN_IN), .ZN(n15174) );
  NAND2_X1 U18556 ( .A1(n15175), .A2(n15174), .ZN(P2_U2888) );
  OAI22_X1 U18557 ( .A1(n15206), .A2(n19053), .B1(n19069), .B2(n15176), .ZN(
        n15177) );
  AOI21_X1 U18558 ( .B1(n19099), .B2(n16179), .A(n15177), .ZN(n15179) );
  AOI22_X1 U18559 ( .A1(n19039), .A2(BUF1_REG_28__SCAN_IN), .B1(n19038), .B2(
        BUF2_REG_28__SCAN_IN), .ZN(n15178) );
  OAI211_X1 U18560 ( .C1(n15180), .C2(n19103), .A(n15179), .B(n15178), .ZN(
        P2_U2891) );
  INV_X1 U18561 ( .A(n15421), .ZN(n15186) );
  OAI22_X1 U18562 ( .A1(n15206), .A2(n19055), .B1(n19069), .B2(n15181), .ZN(
        n15185) );
  INV_X1 U18563 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n15182) );
  OAI22_X1 U18564 ( .A1(n15210), .A2(n15183), .B1(n15208), .B2(n15182), .ZN(
        n15184) );
  AOI211_X1 U18565 ( .C1(n19099), .C2(n15186), .A(n15185), .B(n15184), .ZN(
        n15187) );
  OAI21_X1 U18566 ( .B1(n15188), .B2(n19103), .A(n15187), .ZN(P2_U2892) );
  NAND2_X1 U18567 ( .A1(n15189), .A2(n19086), .ZN(n15196) );
  AOI22_X1 U18568 ( .A1(n19037), .A2(n19057), .B1(n19098), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15195) );
  AOI22_X1 U18569 ( .A1(n19039), .A2(BUF1_REG_26__SCAN_IN), .B1(n19038), .B2(
        BUF2_REG_26__SCAN_IN), .ZN(n15194) );
  NAND2_X1 U18570 ( .A1(n15078), .A2(n15190), .ZN(n15191) );
  AND2_X1 U18571 ( .A1(n15192), .A2(n15191), .ZN(n16192) );
  NAND2_X1 U18572 ( .A1(n19099), .A2(n16192), .ZN(n15193) );
  NAND4_X1 U18573 ( .A1(n15196), .A2(n15195), .A3(n15194), .A4(n15193), .ZN(
        P2_U2893) );
  INV_X1 U18574 ( .A(n15446), .ZN(n15202) );
  OAI22_X1 U18575 ( .A1(n15206), .A2(n19060), .B1(n19069), .B2(n15197), .ZN(
        n15201) );
  INV_X1 U18576 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n15199) );
  INV_X1 U18577 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n15198) );
  OAI22_X1 U18578 ( .A1(n15210), .A2(n15199), .B1(n15208), .B2(n15198), .ZN(
        n15200) );
  AOI211_X1 U18579 ( .C1(n19099), .C2(n15202), .A(n15201), .B(n15200), .ZN(
        n15203) );
  OAI21_X1 U18580 ( .B1(n15204), .B2(n19103), .A(n15203), .ZN(P2_U2894) );
  INV_X1 U18581 ( .A(n15474), .ZN(n15213) );
  OAI22_X1 U18582 ( .A1(n15206), .A2(n19065), .B1(n15205), .B2(n19069), .ZN(
        n15212) );
  INV_X1 U18583 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n15209) );
  INV_X1 U18584 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n15207) );
  OAI22_X1 U18585 ( .A1(n15210), .A2(n15209), .B1(n15208), .B2(n15207), .ZN(
        n15211) );
  AOI211_X1 U18586 ( .C1(n19099), .C2(n15213), .A(n15212), .B(n15211), .ZN(
        n15214) );
  OAI21_X1 U18587 ( .B1(n15215), .B2(n19103), .A(n15214), .ZN(P2_U2896) );
  AOI21_X1 U18588 ( .B1(n15228), .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n15217) );
  NAND2_X1 U18589 ( .A1(n15219), .A2(n15218), .ZN(n15220) );
  XNOR2_X1 U18590 ( .A(n15221), .B(n15220), .ZN(n15412) );
  NOR2_X1 U18591 ( .A1(n19155), .A2(n19748), .ZN(n15401) );
  NOR2_X1 U18592 ( .A1(n15222), .A2(n15396), .ZN(n15223) );
  AOI211_X1 U18593 ( .C1(n15338), .C2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n15401), .B(n15223), .ZN(n15224) );
  OAI21_X1 U18594 ( .B1(n13862), .B2(n15410), .A(n15224), .ZN(n15225) );
  AOI21_X1 U18595 ( .B1(n15412), .B2(n11114), .A(n15225), .ZN(n15226) );
  OAI21_X1 U18596 ( .B1(n15414), .B2(n19148), .A(n15226), .ZN(P2_U2985) );
  XNOR2_X1 U18597 ( .A(n15227), .B(n15417), .ZN(n15427) );
  INV_X1 U18598 ( .A(n15228), .ZN(n15416) );
  NAND2_X1 U18599 ( .A1(n15235), .A2(n15417), .ZN(n15415) );
  NAND3_X1 U18600 ( .A1(n15416), .A2(n16261), .A3(n15415), .ZN(n15234) );
  NAND2_X1 U18601 ( .A1(n15229), .A2(n19141), .ZN(n15230) );
  NAND2_X1 U18602 ( .A1(n18902), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15420) );
  OAI211_X1 U18603 ( .C1(n19154), .C2(n15231), .A(n15230), .B(n15420), .ZN(
        n15232) );
  AOI21_X1 U18604 ( .B1(n19151), .B2(n15424), .A(n15232), .ZN(n15233) );
  OAI211_X1 U18605 ( .C1(n15427), .C2(n19147), .A(n15234), .B(n15233), .ZN(
        P2_U2987) );
  OAI21_X1 U18606 ( .B1(n15250), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15235), .ZN(n15437) );
  NAND2_X1 U18607 ( .A1(n18902), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15430) );
  NAND2_X1 U18608 ( .A1(n15338), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15236) );
  OAI211_X1 U18609 ( .C1(n15237), .C2(n15396), .A(n15430), .B(n15236), .ZN(
        n15244) );
  INV_X1 U18610 ( .A(n15247), .ZN(n15238) );
  AOI21_X1 U18611 ( .B1(n15249), .B2(n15246), .A(n15238), .ZN(n15240) );
  MUX2_X1 U18612 ( .A(n15240), .B(n15246), .S(n15239), .Z(n15242) );
  NOR2_X1 U18613 ( .A1(n15435), .A2(n19147), .ZN(n15243) );
  AOI211_X1 U18614 ( .C1(n19151), .C2(n16193), .A(n15244), .B(n15243), .ZN(
        n15245) );
  OAI21_X1 U18615 ( .B1(n15437), .B2(n19148), .A(n15245), .ZN(P2_U2988) );
  NAND2_X1 U18616 ( .A1(n15247), .A2(n15246), .ZN(n15248) );
  XNOR2_X1 U18617 ( .A(n15249), .B(n15248), .ZN(n15452) );
  INV_X1 U18618 ( .A(n15250), .ZN(n15439) );
  NAND2_X1 U18619 ( .A1(n15454), .A2(n15443), .ZN(n15438) );
  NAND3_X1 U18620 ( .A1(n15439), .A2(n16261), .A3(n15438), .ZN(n15255) );
  NAND2_X1 U18621 ( .A1(n18902), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15445) );
  OAI21_X1 U18622 ( .B1(n19154), .B2(n15251), .A(n15445), .ZN(n15253) );
  NOR2_X1 U18623 ( .A1(n15440), .A2(n13862), .ZN(n15252) );
  AOI211_X1 U18624 ( .C1(n19141), .C2(n9698), .A(n15253), .B(n15252), .ZN(
        n15254) );
  OAI211_X1 U18625 ( .C1(n19147), .C2(n15452), .A(n15255), .B(n15254), .ZN(
        P2_U2989) );
  XNOR2_X1 U18626 ( .A(n15256), .B(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15257) );
  XNOR2_X1 U18627 ( .A(n15258), .B(n15257), .ZN(n15469) );
  NAND2_X1 U18628 ( .A1(n15259), .A2(n15461), .ZN(n15453) );
  NAND3_X1 U18629 ( .A1(n15454), .A2(n16261), .A3(n15453), .ZN(n15264) );
  NOR2_X1 U18630 ( .A1(n19155), .A2(n19739), .ZN(n15460) );
  AOI21_X1 U18631 ( .B1(n15338), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15460), .ZN(n15260) );
  OAI21_X1 U18632 ( .B1(n15261), .B2(n15396), .A(n15260), .ZN(n15262) );
  AOI21_X1 U18633 ( .B1(n15466), .B2(n19151), .A(n15262), .ZN(n15263) );
  OAI211_X1 U18634 ( .C1(n15469), .C2(n19147), .A(n15264), .B(n15263), .ZN(
        P2_U2990) );
  OR2_X1 U18635 ( .A1(n15501), .A2(n15265), .ZN(n15275) );
  NOR2_X1 U18636 ( .A1(n15493), .A2(n15275), .ZN(n15266) );
  OAI21_X1 U18637 ( .B1(n15277), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n15259), .ZN(n15484) );
  XOR2_X1 U18638 ( .A(n15268), .B(n15267), .Z(n15481) );
  NOR2_X1 U18639 ( .A1(n19155), .A2(n19737), .ZN(n15471) );
  NOR2_X1 U18640 ( .A1(n19154), .A2(n15269), .ZN(n15270) );
  AOI211_X1 U18641 ( .C1(n15271), .C2(n19141), .A(n15471), .B(n15270), .ZN(
        n15272) );
  OAI21_X1 U18642 ( .B1(n13862), .B2(n15470), .A(n15272), .ZN(n15273) );
  AOI21_X1 U18643 ( .B1(n15481), .B2(n11114), .A(n15273), .ZN(n15274) );
  OAI21_X1 U18644 ( .B1(n15484), .B2(n19148), .A(n15274), .ZN(P2_U2991) );
  NOR2_X1 U18645 ( .A1(n15276), .A2(n15275), .ZN(n15299) );
  INV_X1 U18646 ( .A(n15277), .ZN(n15278) );
  OAI21_X1 U18647 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15299), .A(
        n15278), .ZN(n15498) );
  NAND2_X1 U18648 ( .A1(n15280), .A2(n15279), .ZN(n15282) );
  NAND2_X1 U18649 ( .A1(n15282), .A2(n15281), .ZN(n15286) );
  NAND2_X1 U18650 ( .A1(n15284), .A2(n15283), .ZN(n15285) );
  XNOR2_X1 U18651 ( .A(n15286), .B(n15285), .ZN(n15496) );
  NOR2_X1 U18652 ( .A1(n19155), .A2(n19735), .ZN(n15486) );
  NOR2_X1 U18653 ( .A1(n15287), .A2(n15396), .ZN(n15288) );
  AOI211_X1 U18654 ( .C1(n15338), .C2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n15486), .B(n15288), .ZN(n15289) );
  OAI21_X1 U18655 ( .B1(n13862), .B2(n15485), .A(n15289), .ZN(n15290) );
  AOI21_X1 U18656 ( .B1(n15496), .B2(n11114), .A(n15290), .ZN(n15291) );
  OAI21_X1 U18657 ( .B1(n15498), .B2(n19148), .A(n15291), .ZN(P2_U2992) );
  AOI21_X1 U18658 ( .B1(n15294), .B2(n15293), .A(n15292), .ZN(n15298) );
  NAND2_X1 U18659 ( .A1(n15296), .A2(n15295), .ZN(n15297) );
  XNOR2_X1 U18660 ( .A(n15298), .B(n15297), .ZN(n15509) );
  AOI21_X1 U18661 ( .B1(n15501), .B2(n15300), .A(n15299), .ZN(n15499) );
  NAND2_X1 U18662 ( .A1(n15499), .A2(n16261), .ZN(n15304) );
  INV_X1 U18663 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19733) );
  OR2_X1 U18664 ( .A1(n19155), .A2(n19733), .ZN(n15503) );
  OAI21_X1 U18665 ( .B1(n19154), .B2(n18858), .A(n15503), .ZN(n15302) );
  NOR2_X1 U18666 ( .A1(n18859), .A2(n13862), .ZN(n15301) );
  AOI211_X1 U18667 ( .C1(n19141), .C2(n18866), .A(n15302), .B(n15301), .ZN(
        n15303) );
  OAI211_X1 U18668 ( .C1(n15509), .C2(n19147), .A(n15304), .B(n15303), .ZN(
        P2_U2993) );
  NOR2_X1 U18669 ( .A1(n15306), .A2(n15305), .ZN(n15308) );
  AOI21_X1 U18670 ( .B1(n15317), .B2(n15320), .A(n15319), .ZN(n15307) );
  XNOR2_X1 U18671 ( .A(n15308), .B(n15307), .ZN(n15521) );
  OAI22_X1 U18672 ( .A1(n15309), .A2(n19154), .B1(n15090), .B2(n19155), .ZN(
        n15311) );
  NOR2_X1 U18673 ( .A1(n15516), .A2(n13862), .ZN(n15310) );
  AOI211_X1 U18674 ( .C1(n15312), .C2(n19141), .A(n15311), .B(n15310), .ZN(
        n15316) );
  INV_X1 U18675 ( .A(n11131), .ZN(n15314) );
  AOI21_X1 U18676 ( .B1(n15513), .B2(n15314), .A(n15313), .ZN(n15519) );
  NAND2_X1 U18677 ( .A1(n15519), .A2(n16261), .ZN(n15315) );
  OAI211_X1 U18678 ( .C1(n15521), .C2(n19147), .A(n15316), .B(n15315), .ZN(
        P2_U2995) );
  INV_X1 U18679 ( .A(n15317), .ZN(n15318) );
  NOR2_X1 U18680 ( .A1(n15319), .A2(n15318), .ZN(n15321) );
  XOR2_X1 U18681 ( .A(n15321), .B(n15320), .Z(n15532) );
  NOR2_X1 U18682 ( .A1(n15322), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15528) );
  NOR3_X1 U18683 ( .A1(n15528), .A2(n11131), .A3(n19148), .ZN(n15328) );
  INV_X1 U18684 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19729) );
  OAI22_X1 U18685 ( .A1(n19729), .A2(n19155), .B1(n15396), .B2(n15323), .ZN(
        n15327) );
  OAI22_X1 U18686 ( .A1(n15325), .A2(n13862), .B1(n15324), .B2(n19154), .ZN(
        n15326) );
  NOR3_X1 U18687 ( .A1(n15328), .A2(n15327), .A3(n15326), .ZN(n15329) );
  OAI21_X1 U18688 ( .B1(n15532), .B2(n19147), .A(n15329), .ZN(P2_U2996) );
  NAND2_X1 U18689 ( .A1(n15331), .A2(n15330), .ZN(n15334) );
  AND2_X1 U18690 ( .A1(n15332), .A2(n9637), .ZN(n15333) );
  XNOR2_X1 U18691 ( .A(n15334), .B(n15333), .ZN(n15541) );
  INV_X1 U18692 ( .A(n15335), .ZN(n15337) );
  INV_X1 U18693 ( .A(n15322), .ZN(n15336) );
  OAI211_X1 U18694 ( .C1(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n15337), .A(
        n15336), .B(n16261), .ZN(n15343) );
  NAND2_X1 U18695 ( .A1(n18893), .A2(n19141), .ZN(n15340) );
  NOR2_X1 U18696 ( .A1(n19155), .A2(n19727), .ZN(n15538) );
  AOI21_X1 U18697 ( .B1(n15338), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n15538), .ZN(n15339) );
  NAND2_X1 U18698 ( .A1(n15340), .A2(n15339), .ZN(n15341) );
  AOI21_X1 U18699 ( .B1(n19151), .B2(n15539), .A(n15341), .ZN(n15342) );
  OAI211_X1 U18700 ( .C1(n15541), .C2(n19147), .A(n15343), .B(n15342), .ZN(
        P2_U2997) );
  NAND2_X1 U18701 ( .A1(n15344), .A2(n15345), .ZN(n15579) );
  INV_X1 U18702 ( .A(n15579), .ZN(n15543) );
  OAI211_X1 U18703 ( .C1(n15543), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n16261), .B(n15335), .ZN(n15354) );
  INV_X1 U18704 ( .A(n15346), .ZN(n15348) );
  AOI221_X1 U18705 ( .B1(n15564), .B2(n15349), .C1(n15348), .C2(n15349), .A(
        n15347), .ZN(n15557) );
  NOR2_X1 U18706 ( .A1(n19155), .A2(n15350), .ZN(n15556) );
  AOI21_X1 U18707 ( .B1(n11114), .B2(n15557), .A(n15556), .ZN(n15351) );
  OAI21_X1 U18708 ( .B1(n9853), .B2(n19154), .A(n15351), .ZN(n15352) );
  AOI21_X1 U18709 ( .B1(n18898), .B2(n19141), .A(n15352), .ZN(n15353) );
  OAI211_X1 U18710 ( .C1(n18903), .C2(n13862), .A(n15354), .B(n15353), .ZN(
        P2_U2998) );
  NAND2_X1 U18711 ( .A1(n15624), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15623) );
  INV_X1 U18712 ( .A(n15623), .ZN(n15366) );
  AND2_X1 U18713 ( .A1(n15344), .A2(n15355), .ZN(n15577) );
  INV_X1 U18714 ( .A(n15577), .ZN(n15356) );
  OAI21_X1 U18715 ( .B1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15594), .A(
        n15356), .ZN(n15593) );
  INV_X1 U18716 ( .A(n15566), .ZN(n15362) );
  INV_X1 U18717 ( .A(n15357), .ZN(n15565) );
  INV_X1 U18718 ( .A(n15358), .ZN(n15361) );
  NAND2_X1 U18719 ( .A1(n15359), .A2(n15565), .ZN(n15360) );
  AOI22_X1 U18720 ( .A1(n15362), .A2(n15565), .B1(n15361), .B2(n15360), .ZN(
        n15591) );
  OAI22_X1 U18721 ( .A1(n10788), .A2(n19155), .B1(n15396), .B2(n18913), .ZN(
        n15364) );
  INV_X1 U18722 ( .A(n18914), .ZN(n15583) );
  OAI22_X1 U18723 ( .A1(n15583), .A2(n13862), .B1(n9855), .B2(n19154), .ZN(
        n15363) );
  AOI211_X1 U18724 ( .C1(n15591), .C2(n11114), .A(n15364), .B(n15363), .ZN(
        n15365) );
  OAI21_X1 U18725 ( .B1(n15593), .B2(n19148), .A(n15365), .ZN(P2_U3000) );
  OR2_X1 U18726 ( .A1(n15623), .A2(n15613), .ZN(n15595) );
  OAI21_X1 U18727 ( .B1(n15366), .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n15595), .ZN(n15622) );
  NAND2_X1 U18728 ( .A1(n15368), .A2(n15367), .ZN(n15370) );
  XOR2_X1 U18729 ( .A(n15370), .B(n15369), .Z(n15620) );
  OAI22_X1 U18730 ( .A1(n11008), .A2(n19155), .B1(n15396), .B2(n15371), .ZN(
        n15374) );
  INV_X1 U18731 ( .A(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n15372) );
  OAI22_X1 U18732 ( .A1(n15617), .A2(n13862), .B1(n15372), .B2(n19154), .ZN(
        n15373) );
  AOI211_X1 U18733 ( .C1(n15620), .C2(n11114), .A(n15374), .B(n15373), .ZN(
        n15375) );
  OAI21_X1 U18734 ( .B1(n15622), .B2(n19148), .A(n15375), .ZN(P2_U3002) );
  INV_X1 U18735 ( .A(n15624), .ZN(n15376) );
  OAI21_X1 U18736 ( .B1(n15344), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n15376), .ZN(n15653) );
  OAI21_X1 U18737 ( .B1(n15390), .B2(n15387), .A(n15388), .ZN(n15381) );
  NAND2_X1 U18738 ( .A1(n10523), .A2(n15379), .ZN(n15380) );
  XNOR2_X1 U18739 ( .A(n15381), .B(n15380), .ZN(n15651) );
  INV_X1 U18740 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19718) );
  OAI22_X1 U18741 ( .A1(n15382), .A2(n19154), .B1(n19718), .B2(n19155), .ZN(
        n15385) );
  INV_X1 U18742 ( .A(n18956), .ZN(n15383) );
  OAI22_X1 U18743 ( .A1(n13862), .A2(n15644), .B1(n15396), .B2(n15383), .ZN(
        n15384) );
  AOI211_X1 U18744 ( .C1(n15651), .C2(n11114), .A(n15385), .B(n15384), .ZN(
        n15386) );
  OAI21_X1 U18745 ( .B1(n15653), .B2(n19148), .A(n15386), .ZN(P2_U3004) );
  NAND2_X1 U18746 ( .A1(n10519), .A2(n15388), .ZN(n15389) );
  XNOR2_X1 U18747 ( .A(n15390), .B(n15389), .ZN(n15655) );
  NAND2_X1 U18748 ( .A1(n15392), .A2(n15391), .ZN(n16252) );
  AOI211_X1 U18749 ( .C1(n16252), .C2(n16253), .A(n15393), .B(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15394) );
  NOR2_X1 U18750 ( .A1(n15394), .A2(n15344), .ZN(n15654) );
  NAND2_X1 U18751 ( .A1(n15654), .A2(n16261), .ZN(n15400) );
  OAI22_X1 U18752 ( .A1(n13806), .A2(n19154), .B1(n15396), .B2(n15395), .ZN(
        n15398) );
  NOR2_X1 U18753 ( .A1(n15659), .A2(n13862), .ZN(n15397) );
  AOI211_X1 U18754 ( .C1(P2_REIP_REG_9__SCAN_IN), .C2(n18902), .A(n15398), .B(
        n15397), .ZN(n15399) );
  OAI211_X1 U18755 ( .C1(n19147), .C2(n15655), .A(n15400), .B(n15399), .ZN(
        P2_U3005) );
  INV_X1 U18756 ( .A(n15401), .ZN(n15405) );
  OAI21_X1 U18757 ( .B1(n15417), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15403) );
  OAI211_X1 U18758 ( .C1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(n15403), .B(n15402), .ZN(
        n15404) );
  OAI211_X1 U18759 ( .C1(n15406), .C2(n19185), .A(n15405), .B(n15404), .ZN(
        n15407) );
  AOI21_X1 U18760 ( .B1(n15408), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n15407), .ZN(n15409) );
  OAI21_X1 U18761 ( .B1(n15410), .B2(n19179), .A(n15409), .ZN(n15411) );
  AOI21_X1 U18762 ( .B1(n15412), .B2(n19188), .A(n15411), .ZN(n15413) );
  OAI21_X1 U18763 ( .B1(n15414), .B2(n19174), .A(n15413), .ZN(P2_U3017) );
  NAND3_X1 U18764 ( .A1(n15416), .A2(n11175), .A3(n15415), .ZN(n15426) );
  NOR2_X1 U18765 ( .A1(n15418), .A2(n15417), .ZN(n15423) );
  OAI211_X1 U18766 ( .C1(n19185), .C2(n15421), .A(n15420), .B(n15419), .ZN(
        n15422) );
  AOI211_X1 U18767 ( .C1(n15424), .C2(n16290), .A(n15423), .B(n15422), .ZN(
        n15425) );
  OAI211_X1 U18768 ( .C1(n15427), .C2(n19157), .A(n15426), .B(n15425), .ZN(
        P2_U3019) );
  INV_X1 U18769 ( .A(n15428), .ZN(n15459) );
  OAI21_X1 U18770 ( .B1(n15461), .B2(n15459), .A(n15534), .ZN(n15441) );
  OAI211_X1 U18771 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n15429), .ZN(n15431) );
  OAI21_X1 U18772 ( .B1(n15442), .B2(n15431), .A(n15430), .ZN(n15432) );
  AOI21_X1 U18773 ( .B1(n16296), .B2(n16192), .A(n15432), .ZN(n15433) );
  OAI21_X1 U18774 ( .B1(n15441), .B2(n15434), .A(n15433), .ZN(n15436) );
  NAND3_X1 U18775 ( .A1(n15439), .A2(n11175), .A3(n15438), .ZN(n15451) );
  INV_X1 U18776 ( .A(n15440), .ZN(n15449) );
  NOR2_X1 U18777 ( .A1(n15441), .A2(n15443), .ZN(n15448) );
  INV_X1 U18778 ( .A(n15442), .ZN(n15462) );
  NAND3_X1 U18779 ( .A1(n15462), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15443), .ZN(n15444) );
  OAI211_X1 U18780 ( .C1(n19185), .C2(n15446), .A(n15445), .B(n15444), .ZN(
        n15447) );
  AOI211_X1 U18781 ( .C1(n15449), .C2(n16290), .A(n15448), .B(n15447), .ZN(
        n15450) );
  OAI211_X1 U18782 ( .C1(n15452), .C2(n19157), .A(n15451), .B(n15450), .ZN(
        P2_U3021) );
  NAND3_X1 U18783 ( .A1(n15454), .A2(n11175), .A3(n15453), .ZN(n15468) );
  NOR2_X1 U18784 ( .A1(n15456), .A2(n15455), .ZN(n15457) );
  OR2_X1 U18785 ( .A1(n15458), .A2(n15457), .ZN(n16213) );
  NAND3_X1 U18786 ( .A1(n15534), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15459), .ZN(n15464) );
  AOI21_X1 U18787 ( .B1(n15462), .B2(n15461), .A(n15460), .ZN(n15463) );
  OAI211_X1 U18788 ( .C1(n19185), .C2(n16213), .A(n15464), .B(n15463), .ZN(
        n15465) );
  AOI21_X1 U18789 ( .B1(n15466), .B2(n16290), .A(n15465), .ZN(n15467) );
  OAI211_X1 U18790 ( .C1(n15469), .C2(n19157), .A(n15468), .B(n15467), .ZN(
        P2_U3022) );
  INV_X1 U18791 ( .A(n15470), .ZN(n15480) );
  INV_X1 U18792 ( .A(n15471), .ZN(n15473) );
  AND2_X1 U18793 ( .A1(n15475), .A2(n15510), .ZN(n15500) );
  AND2_X1 U18794 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15500), .ZN(
        n15476) );
  NAND3_X1 U18795 ( .A1(n15476), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A3(
        n15477), .ZN(n15472) );
  OAI211_X1 U18796 ( .C1(n19185), .C2(n15474), .A(n15473), .B(n15472), .ZN(
        n15479) );
  OAI21_X1 U18797 ( .B1(n15626), .B2(n15475), .A(n15512), .ZN(n15506) );
  AOI21_X1 U18798 ( .B1(n15501), .B2(n15534), .A(n15506), .ZN(n15494) );
  NAND2_X1 U18799 ( .A1(n15476), .A2(n15493), .ZN(n15487) );
  AOI21_X1 U18800 ( .B1(n15494), .B2(n15487), .A(n15477), .ZN(n15478) );
  AOI211_X1 U18801 ( .C1(n15480), .C2(n16290), .A(n15479), .B(n15478), .ZN(
        n15483) );
  NAND2_X1 U18802 ( .A1(n15481), .A2(n19188), .ZN(n15482) );
  OAI211_X1 U18803 ( .C1(n15484), .C2(n19174), .A(n15483), .B(n15482), .ZN(
        P2_U3023) );
  INV_X1 U18804 ( .A(n15485), .ZN(n15491) );
  INV_X1 U18805 ( .A(n15486), .ZN(n15488) );
  OAI211_X1 U18806 ( .C1(n19185), .C2(n15489), .A(n15488), .B(n15487), .ZN(
        n15490) );
  AOI21_X1 U18807 ( .B1(n15491), .B2(n16290), .A(n15490), .ZN(n15492) );
  OAI21_X1 U18808 ( .B1(n15494), .B2(n15493), .A(n15492), .ZN(n15495) );
  AOI21_X1 U18809 ( .B1(n15496), .B2(n19188), .A(n15495), .ZN(n15497) );
  OAI21_X1 U18810 ( .B1(n15498), .B2(n19174), .A(n15497), .ZN(P2_U3024) );
  NAND2_X1 U18811 ( .A1(n15499), .A2(n11175), .ZN(n15508) );
  NAND2_X1 U18812 ( .A1(n15501), .A2(n15500), .ZN(n15502) );
  OAI211_X1 U18813 ( .C1(n19185), .C2(n18870), .A(n15503), .B(n15502), .ZN(
        n15505) );
  NOR2_X1 U18814 ( .A1(n18859), .A2(n19179), .ZN(n15504) );
  AOI211_X1 U18815 ( .C1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15506), .A(
        n15505), .B(n15504), .ZN(n15507) );
  OAI211_X1 U18816 ( .C1(n15509), .C2(n19157), .A(n15508), .B(n15507), .ZN(
        P2_U3025) );
  INV_X1 U18817 ( .A(n15510), .ZN(n15514) );
  NAND2_X1 U18818 ( .A1(P2_REIP_REG_19__SCAN_IN), .A2(n18902), .ZN(n15511) );
  OAI221_X1 U18819 ( .B1(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15514), 
        .C1(n15513), .C2(n15512), .A(n15511), .ZN(n15518) );
  OAI22_X1 U18820 ( .A1(n15516), .A2(n19179), .B1(n15515), .B2(n19185), .ZN(
        n15517) );
  AOI211_X1 U18821 ( .C1(n15519), .C2(n11175), .A(n15518), .B(n15517), .ZN(
        n15520) );
  OAI21_X1 U18822 ( .B1(n15521), .B2(n19157), .A(n15520), .ZN(P2_U3027) );
  NAND2_X1 U18823 ( .A1(n15534), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15526) );
  OAI22_X1 U18824 ( .A1(n19155), .A2(n19729), .B1(
        P2_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n15522), .ZN(n15523) );
  AOI21_X1 U18825 ( .B1(n15524), .B2(n16290), .A(n15523), .ZN(n15525) );
  OAI21_X1 U18826 ( .B1(n15527), .B2(n15526), .A(n15525), .ZN(n15530) );
  NOR3_X1 U18827 ( .A1(n15528), .A2(n11131), .A3(n19174), .ZN(n15529) );
  AOI211_X1 U18828 ( .C1(n16296), .C2(n16227), .A(n15530), .B(n15529), .ZN(
        n15531) );
  OAI21_X1 U18829 ( .B1(n15532), .B2(n19157), .A(n15531), .ZN(P2_U3028) );
  OAI21_X1 U18830 ( .B1(n11175), .B2(n15533), .A(n15335), .ZN(n15536) );
  NAND2_X1 U18831 ( .A1(n15535), .A2(n15534), .ZN(n15574) );
  OAI211_X1 U18832 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15537), .A(
        n15536), .B(n15574), .ZN(n15551) );
  AOI21_X1 U18833 ( .B1(n15544), .B2(n15671), .A(n15551), .ZN(n15550) );
  AOI21_X1 U18834 ( .B1(n15539), .B2(n16290), .A(n15538), .ZN(n15540) );
  OAI21_X1 U18835 ( .B1(n15541), .B2(n19157), .A(n15540), .ZN(n15546) );
  AOI21_X1 U18836 ( .B1(n15543), .B2(n11175), .A(n15542), .ZN(n15562) );
  NOR3_X1 U18837 ( .A1(n15562), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15544), .ZN(n15545) );
  AOI211_X1 U18838 ( .C1(n16296), .C2(n15547), .A(n15546), .B(n15545), .ZN(
        n15548) );
  OAI21_X1 U18839 ( .B1(n15550), .B2(n15549), .A(n15548), .ZN(P2_U3029) );
  NAND2_X1 U18840 ( .A1(n15551), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15561) );
  AND2_X1 U18841 ( .A1(n15553), .A2(n15552), .ZN(n15554) );
  NOR2_X1 U18842 ( .A1(n15555), .A2(n15554), .ZN(n19042) );
  AOI21_X1 U18843 ( .B1(n19188), .B2(n15557), .A(n15556), .ZN(n15558) );
  OAI21_X1 U18844 ( .B1(n19179), .B2(n18903), .A(n15558), .ZN(n15559) );
  AOI21_X1 U18845 ( .B1(n19042), .B2(n16296), .A(n15559), .ZN(n15560) );
  OAI211_X1 U18846 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15562), .A(
        n15561), .B(n15560), .ZN(P2_U3030) );
  NOR2_X1 U18847 ( .A1(n15564), .A2(n15563), .ZN(n15568) );
  NAND2_X1 U18848 ( .A1(n15566), .A2(n15565), .ZN(n15567) );
  XNOR2_X1 U18849 ( .A(n15568), .B(n15567), .ZN(n16232) );
  NAND2_X1 U18850 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n18902), .ZN(n15569) );
  OAI21_X1 U18851 ( .B1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15570), .A(
        n15569), .ZN(n15571) );
  AOI21_X1 U18852 ( .B1(n16290), .B2(n16234), .A(n15571), .ZN(n15572) );
  OAI21_X1 U18853 ( .B1(n15574), .B2(n15573), .A(n15572), .ZN(n15575) );
  AOI21_X1 U18854 ( .B1(n15576), .B2(n16296), .A(n15575), .ZN(n15581) );
  OR2_X1 U18855 ( .A1(n15577), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15578) );
  AND2_X1 U18856 ( .A1(n15579), .A2(n15578), .ZN(n16233) );
  NAND2_X1 U18857 ( .A1(n16233), .A2(n11175), .ZN(n15580) );
  OAI211_X1 U18858 ( .C1(n16232), .C2(n19157), .A(n15581), .B(n15580), .ZN(
        P2_U3031) );
  XNOR2_X1 U18859 ( .A(n15601), .B(n15582), .ZN(n19050) );
  OAI22_X1 U18860 ( .A1(n19179), .A2(n15583), .B1(n10788), .B2(n19155), .ZN(
        n15584) );
  AOI21_X1 U18861 ( .B1(n15586), .B2(n15585), .A(n15584), .ZN(n15589) );
  OAI22_X1 U18862 ( .A1(n15587), .A2(n15614), .B1(n15626), .B2(n15610), .ZN(
        n15604) );
  NAND2_X1 U18863 ( .A1(n15604), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15588) );
  OAI211_X1 U18864 ( .C1(n19050), .C2(n19185), .A(n15589), .B(n15588), .ZN(
        n15590) );
  AOI21_X1 U18865 ( .B1(n15591), .B2(n19188), .A(n15590), .ZN(n15592) );
  OAI21_X1 U18866 ( .B1(n15593), .B2(n19174), .A(n15592), .ZN(P2_U3032) );
  AOI21_X1 U18867 ( .B1(n15596), .B2(n15595), .A(n15594), .ZN(n16242) );
  INV_X1 U18868 ( .A(n16242), .ZN(n15609) );
  AND2_X1 U18869 ( .A1(n15598), .A2(n15597), .ZN(n15599) );
  XNOR2_X1 U18870 ( .A(n15600), .B(n15599), .ZN(n16241) );
  OAI21_X1 U18871 ( .B1(n15615), .B2(n15602), .A(n15601), .ZN(n19052) );
  AOI22_X1 U18872 ( .A1(n16290), .A2(n16240), .B1(P2_REIP_REG_13__SCAN_IN), 
        .B2(n18902), .ZN(n15606) );
  OAI21_X1 U18873 ( .B1(n15613), .B2(n15614), .A(n15596), .ZN(n15603) );
  NAND2_X1 U18874 ( .A1(n15604), .A2(n15603), .ZN(n15605) );
  OAI211_X1 U18875 ( .C1(n19052), .C2(n19185), .A(n15606), .B(n15605), .ZN(
        n15607) );
  AOI21_X1 U18876 ( .B1(n16241), .B2(n19188), .A(n15607), .ZN(n15608) );
  OAI21_X1 U18877 ( .B1(n15609), .B2(n19174), .A(n15608), .ZN(P2_U3033) );
  OR2_X1 U18878 ( .A1(n15626), .A2(n15610), .ZN(n15612) );
  NAND2_X1 U18879 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n18902), .ZN(n15611) );
  OAI221_X1 U18880 ( .B1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n15614), 
        .C1(n15613), .C2(n15612), .A(n15611), .ZN(n15619) );
  AOI21_X1 U18881 ( .B1(n15627), .B2(n15616), .A(n15615), .ZN(n18934) );
  INV_X1 U18882 ( .A(n18934), .ZN(n19054) );
  OAI22_X1 U18883 ( .A1(n19054), .A2(n19185), .B1(n19179), .B2(n15617), .ZN(
        n15618) );
  AOI211_X1 U18884 ( .C1(n15620), .C2(n19188), .A(n15619), .B(n15618), .ZN(
        n15621) );
  OAI21_X1 U18885 ( .B1(n15622), .B2(n19174), .A(n15621), .ZN(P2_U3034) );
  OAI21_X1 U18886 ( .B1(n15624), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15623), .ZN(n16247) );
  INV_X1 U18887 ( .A(n15625), .ZN(n15658) );
  NOR2_X1 U18888 ( .A1(n15626), .A2(n15658), .ZN(n15643) );
  OAI21_X1 U18889 ( .B1(n15629), .B2(n15628), .A(n15627), .ZN(n19056) );
  OAI211_X1 U18890 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n15647), .B(n15630), .ZN(
        n15634) );
  INV_X1 U18891 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n15631) );
  OAI22_X1 U18892 ( .A1(n19179), .A2(n18939), .B1(n15631), .B2(n19155), .ZN(
        n15632) );
  INV_X1 U18893 ( .A(n15632), .ZN(n15633) );
  OAI211_X1 U18894 ( .C1(n19056), .C2(n19185), .A(n15634), .B(n15633), .ZN(
        n15639) );
  NOR2_X1 U18895 ( .A1(n15635), .A2(n9706), .ZN(n15636) );
  XNOR2_X1 U18896 ( .A(n15637), .B(n15636), .ZN(n16248) );
  NOR2_X1 U18897 ( .A1(n16248), .A2(n19157), .ZN(n15638) );
  AOI211_X1 U18898 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15643), .A(
        n15639), .B(n15638), .ZN(n15640) );
  OAI21_X1 U18899 ( .B1(n16247), .B2(n19174), .A(n15640), .ZN(P2_U3035) );
  XNOR2_X1 U18900 ( .A(n15642), .B(n15641), .ZN(n19059) );
  NAND2_X1 U18901 ( .A1(n15643), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15649) );
  OAI22_X1 U18902 ( .A1(n19179), .A2(n15644), .B1(n19718), .B2(n19155), .ZN(
        n15645) );
  AOI21_X1 U18903 ( .B1(n15647), .B2(n15646), .A(n15645), .ZN(n15648) );
  OAI211_X1 U18904 ( .C1(n19185), .C2(n19059), .A(n15649), .B(n15648), .ZN(
        n15650) );
  AOI21_X1 U18905 ( .B1(n15651), .B2(n19188), .A(n15650), .ZN(n15652) );
  OAI21_X1 U18906 ( .B1(n15653), .B2(n19174), .A(n15652), .ZN(P2_U3036) );
  INV_X1 U18907 ( .A(n15654), .ZN(n15664) );
  INV_X1 U18908 ( .A(n15655), .ZN(n15662) );
  NAND2_X1 U18909 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n18902), .ZN(n15656) );
  OAI221_X1 U18910 ( .B1(n15658), .B2(n10526), .C1(n15658), .C2(n15657), .A(
        n15656), .ZN(n15661) );
  OAI22_X1 U18911 ( .A1(n19061), .A2(n19185), .B1(n19179), .B2(n15659), .ZN(
        n15660) );
  AOI211_X1 U18912 ( .C1(n15662), .C2(n19188), .A(n15661), .B(n15660), .ZN(
        n15663) );
  OAI21_X1 U18913 ( .B1(n15664), .B2(n19174), .A(n15663), .ZN(P2_U3037) );
  OAI22_X1 U18914 ( .A1(n15666), .A2(n19179), .B1(n19157), .B2(n15665), .ZN(
        n15667) );
  AOI211_X1 U18915 ( .C1(n15669), .C2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n15668), .B(n15667), .ZN(n15675) );
  NAND2_X1 U18916 ( .A1(n11175), .A2(n15670), .ZN(n15674) );
  OAI211_X1 U18917 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n15671), .B(n19191), .ZN(n15673) );
  NAND2_X1 U18918 ( .A1(n16296), .A2(n19791), .ZN(n15672) );
  NAND4_X1 U18919 ( .A1(n15675), .A2(n15674), .A3(n15673), .A4(n15672), .ZN(
        P2_U3045) );
  INV_X1 U18920 ( .A(n15676), .ZN(n15681) );
  NAND2_X1 U18921 ( .A1(n15681), .A2(n19574), .ZN(n15680) );
  AOI22_X1 U18922 ( .A1(n19575), .A2(n19483), .B1(n19573), .B2(n19463), .ZN(
        n15679) );
  NAND2_X1 U18923 ( .A1(n15684), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n15678) );
  NAND2_X1 U18924 ( .A1(n19576), .A2(n19453), .ZN(n15677) );
  NAND4_X1 U18925 ( .A1(n15680), .A2(n15679), .A3(n15678), .A4(n15677), .ZN(
        P2_U3120) );
  NAND2_X1 U18926 ( .A1(n15681), .A2(n19632), .ZN(n15688) );
  NOR2_X1 U18927 ( .A1(n19216), .A2(n15682), .ZN(n15683) );
  AOI21_X1 U18928 ( .B1(n19630), .B2(n19483), .A(n15683), .ZN(n15687) );
  NAND2_X1 U18929 ( .A1(n15684), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n15686) );
  NAND2_X1 U18930 ( .A1(n19629), .A2(n19453), .ZN(n15685) );
  NAND4_X1 U18931 ( .A1(n15688), .A2(n15687), .A3(n15686), .A4(n15685), .ZN(
        P2_U3127) );
  NAND2_X1 U18932 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18330) );
  INV_X1 U18933 ( .A(n17684), .ZN(n18669) );
  NOR2_X1 U18934 ( .A1(n18149), .A2(n18669), .ZN(n15690) );
  AOI221_X1 U18935 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18330), .C1(n15690), 
        .C2(n18330), .A(n15689), .ZN(n18152) );
  NOR2_X1 U18936 ( .A1(n15691), .A2(n18636), .ZN(n15692) );
  OAI21_X1 U18937 ( .B1(n15692), .B2(n18504), .A(n18153), .ZN(n18150) );
  AOI22_X1 U18938 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18152), .B1(
        n18150), .B2(n18641), .ZN(P3_U2865) );
  AOI211_X1 U18939 ( .C1(n15696), .C2(n15695), .A(n15694), .B(n15693), .ZN(
        n15716) );
  NOR2_X1 U18940 ( .A1(n18164), .A2(n15697), .ZN(n15698) );
  NAND2_X1 U18941 ( .A1(n18598), .A2(n15699), .ZN(n15702) );
  NAND2_X1 U18942 ( .A1(n18164), .A2(n17415), .ZN(n18654) );
  NAND3_X1 U18943 ( .A1(n17356), .A2(n18596), .A3(n18815), .ZN(n15701) );
  NAND4_X1 U18944 ( .A1(n15716), .A2(n15810), .A3(n15702), .A4(n15701), .ZN(
        n18628) );
  NOR2_X1 U18945 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18763), .ZN(n18159) );
  INV_X1 U18946 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18147) );
  NOR2_X1 U18947 ( .A1(n18147), .A2(n18761), .ZN(n15703) );
  INV_X1 U18948 ( .A(n18825), .ZN(n18789) );
  AOI21_X1 U18949 ( .B1(n18612), .B2(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15705) );
  INV_X1 U18950 ( .A(n18622), .ZN(n15704) );
  NOR2_X1 U18951 ( .A1(n15705), .A2(n15704), .ZN(n18650) );
  NAND3_X1 U18952 ( .A1(n18791), .A2(n18789), .A3(n18650), .ZN(n15706) );
  OAI21_X1 U18953 ( .B1(n18791), .B2(n18604), .A(n15706), .ZN(P3_U3284) );
  INV_X1 U18954 ( .A(n18599), .ZN(n15712) );
  NAND2_X1 U18955 ( .A1(n15707), .A2(n18596), .ZN(n15710) );
  OAI21_X1 U18956 ( .B1(n18169), .B2(n9732), .A(n18812), .ZN(n15708) );
  OAI21_X1 U18957 ( .B1(n15709), .B2(n15708), .A(n18815), .ZN(n16519) );
  OAI22_X1 U18958 ( .A1(n15712), .A2(n15711), .B1(n15710), .B2(n16519), .ZN(
        n15713) );
  AOI21_X1 U18959 ( .B1(n18598), .B2(n15714), .A(n15713), .ZN(n15715) );
  INV_X1 U18960 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18080) );
  NOR3_X1 U18961 ( .A1(n18080), .A2(n15717), .A3(n18086), .ZN(n18045) );
  AOI21_X1 U18962 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n17933) );
  INV_X1 U18963 ( .A(n17933), .ZN(n18107) );
  NAND2_X1 U18964 ( .A1(n18045), .A2(n18107), .ZN(n18046) );
  NAND3_X1 U18965 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17934) );
  NOR2_X1 U18966 ( .A1(n18046), .A2(n17934), .ZN(n17955) );
  NAND2_X1 U18967 ( .A1(n17936), .A2(n17955), .ZN(n17886) );
  AOI21_X1 U18968 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n18629), .A(
        n18605), .ZN(n18109) );
  NAND3_X1 U18969 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n18045), .ZN(n18047) );
  NOR2_X1 U18970 ( .A1(n17934), .A2(n18047), .ZN(n17954) );
  NAND2_X1 U18971 ( .A1(n17936), .A2(n17954), .ZN(n15722) );
  OAI22_X1 U18972 ( .A1(n18108), .A2(n17886), .B1(n18109), .B2(n15722), .ZN(
        n16403) );
  NAND2_X1 U18973 ( .A1(n15718), .A2(n16403), .ZN(n17855) );
  NOR3_X1 U18974 ( .A1(n17834), .A2(n18142), .A3(n17855), .ZN(n16397) );
  INV_X1 U18975 ( .A(n18594), .ZN(n17995) );
  NAND2_X1 U18976 ( .A1(n15721), .A2(n17830), .ZN(n16382) );
  INV_X1 U18977 ( .A(n16382), .ZN(n16414) );
  INV_X1 U18978 ( .A(n16410), .ZN(n18600) );
  NAND2_X1 U18979 ( .A1(n17322), .A2(n18140), .ZN(n18062) );
  NOR2_X1 U18980 ( .A1(n15720), .A2(n15719), .ZN(n16415) );
  AOI222_X1 U18981 ( .A1(n15721), .A2(n16397), .B1(n18138), .B2(n16414), .C1(
        n17987), .C2(n16415), .ZN(n15786) );
  INV_X2 U18982 ( .A(n18141), .ZN(n18135) );
  NAND2_X1 U18983 ( .A1(n18125), .A2(n18052), .ZN(n18127) );
  INV_X1 U18984 ( .A(n18108), .ZN(n18627) );
  NOR2_X1 U18985 ( .A1(n18605), .A2(n18627), .ZN(n18027) );
  INV_X1 U18986 ( .A(n18027), .ZN(n17993) );
  NAND2_X1 U18987 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17853) );
  NOR2_X1 U18988 ( .A1(n17854), .A2(n17853), .ZN(n17845) );
  NAND2_X1 U18989 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n17845), .ZN(
        n16365) );
  INV_X1 U18990 ( .A(n17877), .ZN(n15723) );
  INV_X1 U18991 ( .A(n15722), .ZN(n17937) );
  NAND2_X1 U18992 ( .A1(n15723), .A2(n17937), .ZN(n17832) );
  NOR2_X1 U18993 ( .A1(n16365), .A2(n17832), .ZN(n15725) );
  OAI21_X1 U18994 ( .B1(n18790), .B2(n17829), .A(n18629), .ZN(n15724) );
  INV_X1 U18995 ( .A(n17886), .ZN(n17938) );
  NAND2_X1 U18996 ( .A1(n15723), .A2(n17938), .ZN(n17871) );
  OAI21_X1 U18997 ( .B1(n17871), .B2(n16365), .A(n18627), .ZN(n17835) );
  OAI211_X1 U18998 ( .C1(n18110), .C2(n15725), .A(n15724), .B(n17835), .ZN(
        n15781) );
  AOI21_X1 U18999 ( .B1(n17829), .B2(n17993), .A(n15781), .ZN(n16411) );
  NAND2_X1 U19000 ( .A1(n16392), .A2(n17830), .ZN(n16371) );
  AOI22_X1 U19001 ( .A1(n18138), .A2(n16371), .B1(n17987), .B2(n16386), .ZN(
        n15783) );
  OAI221_X1 U19002 ( .B1(n18127), .B2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), 
        .C1(n18127), .C2(n16411), .A(n15783), .ZN(n15726) );
  NOR2_X1 U19003 ( .A1(n18121), .A2(n15726), .ZN(n15731) );
  NAND3_X1 U19004 ( .A1(n16409), .A2(n16410), .A3(n18125), .ZN(n18043) );
  INV_X1 U19005 ( .A(n16413), .ZN(n15727) );
  NOR2_X1 U19006 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17656), .ZN(
        n16406) );
  XOR2_X1 U19007 ( .A(n15729), .B(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .Z(
        n16385) );
  AOI22_X1 U19008 ( .A1(n18100), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n18058), 
        .B2(n16385), .ZN(n15730) );
  OAI221_X1 U19009 ( .B1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15786), 
        .C1(n16383), .C2(n15731), .A(n15730), .ZN(P3_U2833) );
  AOI21_X1 U19010 ( .B1(n15732), .B2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n20519), .ZN(n15733) );
  NAND2_X1 U19011 ( .A1(n15734), .A2(n15733), .ZN(n15736) );
  INV_X1 U19012 ( .A(n15736), .ZN(n15740) );
  INV_X1 U19013 ( .A(n15735), .ZN(n15738) );
  AOI22_X1 U19014 ( .A1(n15738), .A2(n15737), .B1(n20424), .B2(n15736), .ZN(
        n15739) );
  AOI21_X1 U19015 ( .B1(n15740), .B2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n15739), .ZN(n15742) );
  INV_X1 U19016 ( .A(n15742), .ZN(n15744) );
  OAI21_X1 U19017 ( .B1(n15742), .B2(n20488), .A(n15741), .ZN(n15743) );
  OAI21_X1 U19018 ( .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15744), .A(
        n15743), .ZN(n15746) );
  AOI222_X1 U19019 ( .A1(n15746), .A2(n20738), .B1(n15746), .B2(n15745), .C1(
        n20738), .C2(n15745), .ZN(n15747) );
  OR2_X1 U19020 ( .A1(n15747), .A2(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n15760) );
  INV_X1 U19021 ( .A(n15748), .ZN(n15758) );
  INV_X1 U19022 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n15749) );
  AND2_X1 U19023 ( .A1(n19851), .A2(n15749), .ZN(n15755) );
  NOR2_X1 U19024 ( .A1(n15751), .A2(n15750), .ZN(n15752) );
  OAI211_X1 U19025 ( .C1(n15755), .C2(n15754), .A(n15753), .B(n15752), .ZN(
        n15756) );
  AOI21_X1 U19026 ( .B1(n15758), .B2(n15757), .A(n15756), .ZN(n15759) );
  INV_X1 U19027 ( .A(n15775), .ZN(n15766) );
  NAND3_X1 U19028 ( .A1(n15762), .A2(n20120), .A3(n15761), .ZN(n15765) );
  OAI21_X1 U19029 ( .B1(n15763), .B2(n20760), .A(n20660), .ZN(n15764) );
  NAND2_X1 U19030 ( .A1(n15765), .A2(n15764), .ZN(n16158) );
  NOR2_X1 U19031 ( .A1(n20755), .A2(n15767), .ZN(n15768) );
  NOR2_X1 U19032 ( .A1(n16162), .A2(n15768), .ZN(n15773) );
  AOI211_X1 U19033 ( .C1(n20674), .C2(n20752), .A(n15770), .B(n15769), .ZN(
        n15771) );
  NAND2_X1 U19034 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n15771), .ZN(n15772) );
  OAI22_X1 U19035 ( .A1(n15773), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n16162), 
        .B2(n15772), .ZN(n15774) );
  OAI21_X1 U19036 ( .B1(n15775), .B2(n19845), .A(n15774), .ZN(P1_U3161) );
  NAND2_X1 U19037 ( .A1(n16392), .A2(n15782), .ZN(n16377) );
  NAND2_X1 U19038 ( .A1(n15777), .A2(n15776), .ZN(n15778) );
  XOR2_X1 U19039 ( .A(n15778), .B(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .Z(
        n16373) );
  INV_X1 U19040 ( .A(n18052), .ZN(n15779) );
  OAI21_X1 U19041 ( .B1(n15779), .B2(n16392), .A(n18125), .ZN(n15780) );
  OAI21_X1 U19042 ( .B1(n15781), .B2(n15780), .A(n18141), .ZN(n16394) );
  AOI21_X1 U19043 ( .B1(n15783), .B2(n16394), .A(n15782), .ZN(n15784) );
  AOI21_X1 U19044 ( .B1(n18058), .B2(n16373), .A(n15784), .ZN(n15785) );
  NAND2_X1 U19045 ( .A1(n18100), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16367) );
  OAI211_X1 U19046 ( .C1(n15786), .C2(n16377), .A(n15785), .B(n16367), .ZN(
        P3_U2832) );
  INV_X1 U19047 ( .A(HOLD), .ZN(n20670) );
  NAND2_X1 U19048 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(
        P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20664) );
  OAI21_X1 U19049 ( .B1(n20670), .B2(n20663), .A(n20664), .ZN(n15787) );
  OAI21_X1 U19050 ( .B1(n20670), .B2(n11618), .A(n15787), .ZN(n15789) );
  NAND2_X1 U19051 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20674), .ZN(n20669) );
  NAND3_X1 U19052 ( .A1(n15789), .A2(n15788), .A3(n20669), .ZN(P1_U3195) );
  NAND2_X1 U19053 ( .A1(n15791), .A2(n15790), .ZN(n15792) );
  XNOR2_X1 U19054 ( .A(n15792), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15972) );
  NOR3_X1 U19055 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n16065), .A3(
        n16066), .ZN(n15793) );
  AOI21_X1 U19056 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(n16052), .A(n15793), 
        .ZN(n15803) );
  AND2_X1 U19057 ( .A1(n15795), .A2(n15794), .ZN(n15796) );
  OAI21_X1 U19058 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n15796), .A(
        n9595), .ZN(n15801) );
  INV_X1 U19059 ( .A(n15797), .ZN(n15798) );
  AOI21_X1 U19060 ( .B1(n15800), .B2(n15799), .A(n15798), .ZN(n15938) );
  AOI22_X1 U19061 ( .A1(n15801), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        n16142), .B2(n15938), .ZN(n15802) );
  OAI211_X1 U19062 ( .C1(n15972), .C2(n16111), .A(n15803), .B(n15802), .ZN(
        P1_U3011) );
  NOR2_X1 U19063 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n15804) );
  NOR2_X1 U19064 ( .A1(n19822), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19675) );
  INV_X1 U19065 ( .A(n19675), .ZN(n18833) );
  NOR2_X1 U19066 ( .A1(n19825), .A2(n18833), .ZN(n16347) );
  INV_X1 U19067 ( .A(n16363), .ZN(n16348) );
  NOR4_X1 U19068 ( .A1(n15805), .A2(n15804), .A3(n16347), .A4(n16348), .ZN(
        P2_U3178) );
  OAI221_X1 U19069 ( .B1(n15806), .B2(n16363), .C1(n10069), .C2(n16363), .A(
        n19565), .ZN(n19800) );
  NOR2_X1 U19070 ( .A1(n15807), .A2(n19800), .ZN(P2_U3047) );
  NAND2_X1 U19071 ( .A1(n18193), .A2(n17207), .ZN(n17349) );
  INV_X1 U19072 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17413) );
  AOI22_X1 U19073 ( .A1(n17348), .A2(BUF2_REG_0__SCAN_IN), .B1(n17347), .B2(
        n15811), .ZN(n15812) );
  OAI221_X1 U19074 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17349), .C1(n17413), 
        .C2(n17207), .A(n15812), .ZN(P3_U2735) );
  NAND2_X1 U19075 ( .A1(n19881), .A2(n14667), .ZN(n15818) );
  INV_X1 U19076 ( .A(n15813), .ZN(n15817) );
  OAI22_X1 U19077 ( .A1(n15814), .A2(n19941), .B1(n19940), .B2(n15960), .ZN(
        n15815) );
  AOI21_X1 U19078 ( .B1(n19938), .B2(P1_EBX_REG_24__SCAN_IN), .A(n15815), .ZN(
        n15816) );
  OAI21_X1 U19079 ( .B1(n15818), .B2(n15817), .A(n15816), .ZN(n15819) );
  AOI21_X1 U19080 ( .B1(n15826), .B2(P1_REIP_REG_24__SCAN_IN), .A(n15819), 
        .ZN(n15822) );
  OAI22_X1 U19081 ( .A1(n15956), .A2(n15891), .B1(n16038), .B2(n19897), .ZN(
        n15820) );
  INV_X1 U19082 ( .A(n15820), .ZN(n15821) );
  NAND2_X1 U19083 ( .A1(n15822), .A2(n15821), .ZN(P1_U2816) );
  OAI22_X1 U19084 ( .A1(n19895), .A2(n15824), .B1(n19941), .B2(n15823), .ZN(
        n15831) );
  NOR3_X1 U19085 ( .A1(n15911), .A2(n15859), .A3(n15825), .ZN(n15835) );
  AOI21_X1 U19086 ( .B1(P1_REIP_REG_22__SCAN_IN), .B2(n15835), .A(
        P1_REIP_REG_23__SCAN_IN), .ZN(n15828) );
  INV_X1 U19087 ( .A(n15826), .ZN(n15827) );
  OAI22_X1 U19088 ( .A1(n15829), .A2(n15891), .B1(n15828), .B2(n15827), .ZN(
        n15830) );
  OAI21_X1 U19089 ( .B1(n19897), .B2(n15834), .A(n15833), .ZN(P1_U2817) );
  AOI22_X1 U19090 ( .A1(n19938), .A2(P1_EBX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n19926), .ZN(n15841) );
  INV_X1 U19091 ( .A(n15967), .ZN(n15836) );
  AOI22_X1 U19092 ( .A1(n15836), .A2(n19927), .B1(n15835), .B2(n20707), .ZN(
        n15840) );
  AOI22_X1 U19093 ( .A1(n15964), .A2(n19904), .B1(n19945), .B2(n16053), .ZN(
        n15839) );
  NOR2_X1 U19094 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(n15911), .ZN(n15842) );
  INV_X1 U19095 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20704) );
  NOR2_X1 U19096 ( .A1(n15859), .A2(n20704), .ZN(n15843) );
  OAI21_X1 U19097 ( .B1(n15843), .B2(n15911), .A(n15837), .ZN(n15860) );
  OAI21_X1 U19098 ( .B1(n15842), .B2(n15860), .A(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n15838) );
  NAND4_X1 U19099 ( .A1(n15841), .A2(n15840), .A3(n15839), .A4(n15838), .ZN(
        P1_U2818) );
  AOI22_X1 U19100 ( .A1(n15844), .A2(n19927), .B1(n15843), .B2(n15842), .ZN(
        n15852) );
  OAI22_X1 U19101 ( .A1(n19895), .A2(n15846), .B1(n19941), .B2(n15845), .ZN(
        n15850) );
  OAI22_X1 U19102 ( .A1(n15848), .A2(n15891), .B1(n15847), .B2(n19897), .ZN(
        n15849) );
  AOI211_X1 U19103 ( .C1(P1_REIP_REG_21__SCAN_IN), .C2(n15860), .A(n15850), 
        .B(n15849), .ZN(n15851) );
  NAND2_X1 U19104 ( .A1(n15852), .A2(n15851), .ZN(P1_U2819) );
  OAI22_X1 U19105 ( .A1(n19895), .A2(n15940), .B1(n19940), .B2(n15853), .ZN(
        n15854) );
  AOI21_X1 U19106 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19926), .A(
        n15854), .ZN(n15864) );
  INV_X1 U19107 ( .A(n15855), .ZN(n15856) );
  AOI21_X1 U19108 ( .B1(n15858), .B2(n15857), .A(n15856), .ZN(n15969) );
  AOI22_X1 U19109 ( .A1(n15969), .A2(n19904), .B1(n19945), .B2(n15938), .ZN(
        n15863) );
  NOR2_X1 U19110 ( .A1(n15911), .A2(n15859), .ZN(n15861) );
  OAI21_X1 U19111 ( .B1(P1_REIP_REG_20__SCAN_IN), .B2(n15861), .A(n15860), 
        .ZN(n15862) );
  NAND3_X1 U19112 ( .A1(n15864), .A2(n15863), .A3(n15862), .ZN(P1_U2820) );
  INV_X1 U19113 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n15866) );
  NAND2_X1 U19114 ( .A1(n15875), .A2(n15865), .ZN(n15877) );
  NOR3_X1 U19115 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n15866), .A3(n15877), 
        .ZN(n15872) );
  INV_X1 U19116 ( .A(n15867), .ZN(n15870) );
  NAND2_X1 U19117 ( .A1(n19938), .A2(P1_EBX_REG_19__SCAN_IN), .ZN(n15869) );
  AOI21_X1 U19118 ( .B1(n19926), .B2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n19913), .ZN(n15868) );
  OAI211_X1 U19119 ( .C1(n15870), .C2(n19940), .A(n15869), .B(n15868), .ZN(
        n15871) );
  AOI211_X1 U19120 ( .C1(n15873), .C2(n19904), .A(n15872), .B(n15871), .ZN(
        n15879) );
  AOI21_X1 U19121 ( .B1(n15875), .B2(n15874), .A(n15911), .ZN(n15876) );
  OR2_X1 U19122 ( .A1(n15876), .A2(n15918), .ZN(n15895) );
  NOR2_X1 U19123 ( .A1(P1_REIP_REG_18__SCAN_IN), .A2(n15877), .ZN(n15885) );
  OAI21_X1 U19124 ( .B1(n15895), .B2(n15885), .A(P1_REIP_REG_19__SCAN_IN), 
        .ZN(n15878) );
  OAI211_X1 U19125 ( .C1(n16060), .C2(n19897), .A(n15879), .B(n15878), .ZN(
        P1_U2821) );
  OAI22_X1 U19126 ( .A1(n15881), .A2(n15891), .B1(n19897), .B2(n15880), .ZN(
        n15882) );
  INV_X1 U19127 ( .A(n15882), .ZN(n15888) );
  AOI22_X1 U19128 ( .A1(n15895), .A2(P1_REIP_REG_18__SCAN_IN), .B1(n19938), 
        .B2(P1_EBX_REG_18__SCAN_IN), .ZN(n15883) );
  OAI211_X1 U19129 ( .C1(n19941), .C2(n14908), .A(n15883), .B(n15929), .ZN(
        n15884) );
  AOI211_X1 U19130 ( .C1(n19927), .C2(n15886), .A(n15885), .B(n15884), .ZN(
        n15887) );
  NAND2_X1 U19131 ( .A1(n15888), .A2(n15887), .ZN(P1_U2822) );
  AOI21_X1 U19132 ( .B1(n19926), .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .A(
        n19913), .ZN(n15889) );
  OAI21_X1 U19133 ( .B1(n19940), .B2(n15890), .A(n15889), .ZN(n15894) );
  NOR2_X1 U19134 ( .A1(n15892), .A2(n15891), .ZN(n15893) );
  AOI211_X1 U19135 ( .C1(n19938), .C2(P1_EBX_REG_17__SCAN_IN), .A(n15894), .B(
        n15893), .ZN(n15898) );
  OAI221_X1 U19136 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(P1_REIP_REG_16__SCAN_IN), .C1(P1_REIP_REG_17__SCAN_IN), .C2(n15896), .A(n15895), .ZN(n15897) );
  OAI211_X1 U19137 ( .C1(n15899), .C2(n19897), .A(n15898), .B(n15897), .ZN(
        P1_U2823) );
  AOI22_X1 U19138 ( .A1(n15990), .A2(n19927), .B1(n19945), .B2(n16086), .ZN(
        n15906) );
  AOI22_X1 U19139 ( .A1(n19938), .A2(P1_EBX_REG_14__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19926), .ZN(n15905) );
  INV_X1 U19140 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n20696) );
  OAI21_X1 U19141 ( .B1(n15901), .B2(n15900), .A(n20696), .ZN(n15903) );
  AOI22_X1 U19142 ( .A1(n15991), .A2(n19904), .B1(n15903), .B2(n15902), .ZN(
        n15904) );
  NAND4_X1 U19143 ( .A1(n15906), .A2(n15905), .A3(n15904), .A4(n15929), .ZN(
        P1_U2826) );
  AOI22_X1 U19144 ( .A1(n19938), .A2(P1_EBX_REG_12__SCAN_IN), .B1(n19927), 
        .B2(n15999), .ZN(n15917) );
  AND2_X1 U19145 ( .A1(n15908), .A2(n15907), .ZN(n15909) );
  NOR2_X1 U19146 ( .A1(n15910), .A2(n15909), .ZN(n16101) );
  AOI22_X1 U19147 ( .A1(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19926), .B1(
        n19945), .B2(n16101), .ZN(n15916) );
  NOR2_X1 U19148 ( .A1(n15911), .A2(n15928), .ZN(n15920) );
  NAND2_X1 U19149 ( .A1(P1_REIP_REG_11__SCAN_IN), .A2(n15920), .ZN(n15912) );
  NAND2_X1 U19150 ( .A1(n16104), .A2(n15912), .ZN(n15913) );
  AOI22_X1 U19151 ( .A1(n19904), .A2(n15998), .B1(n15914), .B2(n15913), .ZN(
        n15915) );
  NAND4_X1 U19152 ( .A1(n15917), .A2(n15916), .A3(n15915), .A4(n15929), .ZN(
        P1_U2828) );
  AOI21_X1 U19153 ( .B1(n19881), .B2(n15928), .A(n15918), .ZN(n15937) );
  OAI22_X1 U19154 ( .A1(n19895), .A2(n15919), .B1(n19940), .B2(n16006), .ZN(
        n15924) );
  AOI22_X1 U19155 ( .A1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n19926), .B1(
        n15920), .B2(n15064), .ZN(n15921) );
  OAI211_X1 U19156 ( .C1(n15922), .C2(n19897), .A(n15921), .B(n15929), .ZN(
        n15923) );
  AOI211_X1 U19157 ( .C1(n19904), .C2(n16002), .A(n15924), .B(n15923), .ZN(
        n15925) );
  OAI21_X1 U19158 ( .B1(n15937), .B2(n15064), .A(n15925), .ZN(P1_U2829) );
  INV_X1 U19159 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n15936) );
  AOI22_X1 U19160 ( .A1(n15926), .A2(n19927), .B1(n19945), .B2(n16115), .ZN(
        n15935) );
  AND3_X1 U19161 ( .A1(n19881), .A2(n15928), .A3(n15927), .ZN(n15932) );
  NAND2_X1 U19162 ( .A1(n19938), .A2(P1_EBX_REG_10__SCAN_IN), .ZN(n15930) );
  OAI211_X1 U19163 ( .C1(n14957), .C2(n19941), .A(n15930), .B(n15929), .ZN(
        n15931) );
  AOI211_X1 U19164 ( .C1(n15933), .C2(n19904), .A(n15932), .B(n15931), .ZN(
        n15934) );
  OAI211_X1 U19165 ( .C1(n15937), .C2(n15936), .A(n15935), .B(n15934), .ZN(
        P1_U2830) );
  AOI22_X1 U19166 ( .A1(n15969), .A2(n15942), .B1(n15941), .B2(n15938), .ZN(
        n15939) );
  OAI21_X1 U19167 ( .B1(n15945), .B2(n15940), .A(n15939), .ZN(P1_U2852) );
  AOI22_X1 U19168 ( .A1(n15998), .A2(n15942), .B1(n15941), .B2(n16101), .ZN(
        n15943) );
  OAI21_X1 U19169 ( .B1(n15945), .B2(n15944), .A(n15943), .ZN(P1_U2860) );
  INV_X1 U19170 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16442) );
  INV_X1 U19171 ( .A(n20131), .ZN(n19988) );
  AOI22_X1 U19172 ( .A1(n15947), .A2(n19988), .B1(n15946), .B2(
        P1_EAX_REG_20__SCAN_IN), .ZN(n15951) );
  AOI22_X1 U19173 ( .A1(n15969), .A2(n15949), .B1(n15948), .B2(DATAI_20_), 
        .ZN(n15950) );
  OAI211_X1 U19174 ( .C1(n15952), .C2(n16442), .A(n15951), .B(n15950), .ZN(
        P1_U2884) );
  AOI22_X1 U19175 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .B1(
        n16052), .B2(P1_REIP_REG_24__SCAN_IN), .ZN(n15959) );
  NAND2_X1 U19176 ( .A1(n14411), .A2(n15954), .ZN(n15953) );
  MUX2_X1 U19177 ( .A(n15954), .B(n15953), .S(n10059), .Z(n15955) );
  XNOR2_X1 U19178 ( .A(n15955), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n16040) );
  INV_X1 U19179 ( .A(n15956), .ZN(n15957) );
  AOI22_X1 U19180 ( .A1(n16040), .A2(n20093), .B1(n15957), .B2(n16022), .ZN(
        n15958) );
  OAI211_X1 U19181 ( .C1(n16019), .C2(n15960), .A(n15959), .B(n15958), .ZN(
        P1_U2975) );
  AOI22_X1 U19182 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n16052), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15966) );
  NAND2_X1 U19183 ( .A1(n15962), .A2(n15961), .ZN(n15963) );
  XNOR2_X1 U19184 ( .A(n15963), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n16050) );
  AOI22_X1 U19185 ( .A1(n15964), .A2(n16022), .B1(n20093), .B2(n16050), .ZN(
        n15965) );
  OAI211_X1 U19186 ( .C1(n16019), .C2(n15967), .A(n15966), .B(n15965), .ZN(
        P1_U2977) );
  AOI22_X1 U19187 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n16052), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n15971) );
  AOI22_X1 U19188 ( .A1(n15969), .A2(n16022), .B1(n15968), .B2(n16021), .ZN(
        n15970) );
  OAI211_X1 U19189 ( .C1(n15972), .C2(n19850), .A(n15971), .B(n15970), .ZN(
        P1_U2979) );
  AOI22_X1 U19190 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n16052), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15983) );
  NAND2_X1 U19191 ( .A1(n15974), .A2(n15973), .ZN(n15977) );
  INV_X1 U19192 ( .A(n15975), .ZN(n15976) );
  NAND2_X1 U19193 ( .A1(n15977), .A2(n15976), .ZN(n15979) );
  NOR2_X1 U19194 ( .A1(n15980), .A2(n20102), .ZN(n15981) );
  AOI21_X1 U19195 ( .B1(n16071), .B2(n20093), .A(n15981), .ZN(n15982) );
  OAI211_X1 U19196 ( .C1(n16019), .C2(n15984), .A(n15983), .B(n15982), .ZN(
        P1_U2983) );
  NAND2_X1 U19197 ( .A1(n15986), .A2(n15985), .ZN(n15989) );
  XNOR2_X1 U19198 ( .A(n15987), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15988) );
  XNOR2_X1 U19199 ( .A(n15989), .B(n15988), .ZN(n16091) );
  AOI22_X1 U19200 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n16052), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15993) );
  AOI22_X1 U19201 ( .A1(n15991), .A2(n16022), .B1(n15990), .B2(n16021), .ZN(
        n15992) );
  OAI211_X1 U19202 ( .C1(n16091), .C2(n19850), .A(n15993), .B(n15992), .ZN(
        P1_U2985) );
  OAI21_X1 U19203 ( .B1(n15996), .B2(n15995), .A(n15994), .ZN(n15997) );
  INV_X1 U19204 ( .A(n15997), .ZN(n16112) );
  AOI22_X1 U19205 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n16141), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n16001) );
  AOI22_X1 U19206 ( .A1(n16021), .A2(n15999), .B1(n16022), .B2(n15998), .ZN(
        n16000) );
  OAI211_X1 U19207 ( .C1(n16112), .C2(n19850), .A(n16001), .B(n16000), .ZN(
        P1_U2987) );
  AOI22_X1 U19208 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n16052), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n16005) );
  AOI22_X1 U19209 ( .A1(n20093), .A2(n16003), .B1(n16022), .B2(n16002), .ZN(
        n16004) );
  OAI211_X1 U19210 ( .C1(n16019), .C2(n16006), .A(n16005), .B(n16004), .ZN(
        P1_U2988) );
  AOI22_X1 U19211 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n16141), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n16012) );
  NAND2_X1 U19212 ( .A1(n16008), .A2(n16007), .ZN(n16009) );
  NAND2_X1 U19213 ( .A1(n16010), .A2(n16009), .ZN(n16137) );
  AOI22_X1 U19214 ( .A1(n16137), .A2(n20093), .B1(n16022), .B2(n19888), .ZN(
        n16011) );
  OAI211_X1 U19215 ( .C1(n16019), .C2(n19885), .A(n16012), .B(n16011), .ZN(
        P1_U2992) );
  AOI22_X1 U19216 ( .A1(n20091), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n16141), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n16018) );
  NAND2_X1 U19217 ( .A1(n16014), .A2(n16013), .ZN(n16015) );
  XNOR2_X1 U19218 ( .A(n16016), .B(n16015), .ZN(n16145) );
  AOI22_X1 U19219 ( .A1(n16145), .A2(n20093), .B1(n16022), .B2(n19905), .ZN(
        n16017) );
  OAI211_X1 U19220 ( .C1(n16019), .C2(n19910), .A(n16018), .B(n16017), .ZN(
        P1_U2993) );
  INV_X1 U19221 ( .A(n16020), .ZN(n19921) );
  AOI222_X1 U19222 ( .A1(n16023), .A2(n20093), .B1(n16022), .B2(n19921), .C1(
        n19914), .C2(n16021), .ZN(n16025) );
  OAI211_X1 U19223 ( .C1(n16027), .C2(n16026), .A(n16025), .B(n16024), .ZN(
        P1_U2994) );
  INV_X1 U19224 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n16037) );
  INV_X1 U19225 ( .A(n16028), .ZN(n16031) );
  INV_X1 U19226 ( .A(n16029), .ZN(n16030) );
  AOI22_X1 U19227 ( .A1(n16031), .A2(n16144), .B1(n16142), .B2(n16030), .ZN(
        n16036) );
  OAI22_X1 U19228 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n16034), .B1(
        n16033), .B2(n16032), .ZN(n16035) );
  OAI211_X1 U19229 ( .C1(n16037), .C2(n16103), .A(n16036), .B(n16035), .ZN(
        P1_U3005) );
  INV_X1 U19230 ( .A(n16038), .ZN(n16039) );
  AOI22_X1 U19231 ( .A1(n16040), .A2(n16144), .B1(n16142), .B2(n16039), .ZN(
        n16049) );
  NAND2_X1 U19232 ( .A1(n16052), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n16048) );
  NOR2_X1 U19233 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n16041), .ZN(
        n16043) );
  OAI21_X1 U19234 ( .B1(n16043), .B2(n16042), .A(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16047) );
  OR3_X1 U19235 ( .A1(n16045), .A2(n16044), .A3(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n16046) );
  NAND4_X1 U19236 ( .A1(n16049), .A2(n16048), .A3(n16047), .A4(n16046), .ZN(
        P1_U3007) );
  AOI22_X1 U19237 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n16051), .B1(
        n16144), .B2(n16050), .ZN(n16059) );
  NAND2_X1 U19238 ( .A1(n16052), .A2(P1_REIP_REG_22__SCAN_IN), .ZN(n16058) );
  NAND2_X1 U19239 ( .A1(n16053), .A2(n16142), .ZN(n16057) );
  OAI211_X1 U19240 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n16055), .B(n16054), .ZN(
        n16056) );
  NAND4_X1 U19241 ( .A1(n16059), .A2(n16058), .A3(n16057), .A4(n16056), .ZN(
        P1_U3009) );
  OAI22_X1 U19242 ( .A1(n16060), .A2(n16068), .B1(n14899), .B2(n16103), .ZN(
        n16061) );
  AOI21_X1 U19243 ( .B1(n16144), .B2(n16062), .A(n16061), .ZN(n16063) );
  OAI221_X1 U19244 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n16066), 
        .C1(n16065), .C2(n9595), .A(n16063), .ZN(P1_U3012) );
  OAI21_X1 U19245 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n16067), .ZN(n16074) );
  OAI22_X1 U19246 ( .A1(n16069), .A2(n16068), .B1(n16103), .B2(n20830), .ZN(
        n16070) );
  INV_X1 U19247 ( .A(n16070), .ZN(n16073) );
  OAI21_X1 U19248 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16131), .A(
        n16099), .ZN(n16078) );
  AOI22_X1 U19249 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n16078), .B1(
        n16144), .B2(n16071), .ZN(n16072) );
  OAI211_X1 U19250 ( .C1(n16081), .C2(n16074), .A(n16073), .B(n16072), .ZN(
        P1_U3015) );
  AOI21_X1 U19251 ( .B1(n16076), .B2(n16142), .A(n16075), .ZN(n16080) );
  AOI22_X1 U19252 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n16078), .B1(
        n16144), .B2(n16077), .ZN(n16079) );
  OAI211_X1 U19253 ( .C1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n16081), .A(
        n16080), .B(n16079), .ZN(P1_U3016) );
  NOR2_X1 U19254 ( .A1(n16083), .A2(n16082), .ZN(n16085) );
  INV_X1 U19255 ( .A(n16099), .ZN(n16084) );
  MUX2_X1 U19256 ( .A(n16085), .B(n16084), .S(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .Z(n16089) );
  NAND2_X1 U19257 ( .A1(n16086), .A2(n16142), .ZN(n16087) );
  OAI21_X1 U19258 ( .B1(n20696), .B2(n16103), .A(n16087), .ZN(n16088) );
  NOR2_X1 U19259 ( .A1(n16089), .A2(n16088), .ZN(n16090) );
  OAI21_X1 U19260 ( .B1(n16091), .B2(n16111), .A(n16090), .ZN(P1_U3017) );
  AOI21_X1 U19261 ( .B1(n16093), .B2(n16142), .A(n16092), .ZN(n16097) );
  AOI22_X1 U19262 ( .A1(n16095), .A2(n16144), .B1(n16098), .B2(n16094), .ZN(
        n16096) );
  OAI211_X1 U19263 ( .C1(n16099), .C2(n16098), .A(n16097), .B(n16096), .ZN(
        P1_U3018) );
  AOI221_X1 U19264 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n16100), 
        .C1(n16127), .C2(n16100), .A(n16107), .ZN(n16106) );
  NAND2_X1 U19265 ( .A1(n16101), .A2(n16142), .ZN(n16102) );
  OAI21_X1 U19266 ( .B1(n16104), .B2(n16103), .A(n16102), .ZN(n16105) );
  NOR2_X1 U19267 ( .A1(n16106), .A2(n16105), .ZN(n16110) );
  NAND3_X1 U19268 ( .A1(n16108), .A2(n16143), .A3(n16107), .ZN(n16109) );
  OAI211_X1 U19269 ( .C1(n16112), .C2(n16111), .A(n16110), .B(n16109), .ZN(
        P1_U3019) );
  INV_X1 U19270 ( .A(n16113), .ZN(n16114) );
  AOI21_X1 U19271 ( .B1(n16115), .B2(n16142), .A(n16114), .ZN(n16123) );
  AOI22_X1 U19272 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n16117), .B1(
        n16144), .B2(n16116), .ZN(n16122) );
  OAI221_X1 U19273 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n16120), .C2(n16119), .A(
        n16118), .ZN(n16121) );
  NAND3_X1 U19274 ( .A1(n16123), .A2(n16122), .A3(n16121), .ZN(P1_U3021) );
  OAI21_X1 U19275 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16124), .ZN(n16135) );
  AOI21_X1 U19276 ( .B1(n16126), .B2(n16142), .A(n16125), .ZN(n16134) );
  INV_X1 U19277 ( .A(n16128), .ZN(n16130) );
  AOI21_X1 U19278 ( .B1(n14535), .B2(n16130), .A(n16129), .ZN(n16149) );
  OAI21_X1 U19279 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16131), .A(
        n16149), .ZN(n16136) );
  AOI22_X1 U19280 ( .A1(n16132), .A2(n16144), .B1(
        P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n16136), .ZN(n16133) );
  OAI211_X1 U19281 ( .C1(n16140), .C2(n16135), .A(n16134), .B(n16133), .ZN(
        P1_U3023) );
  AOI22_X1 U19282 ( .A1(n19887), .A2(n16142), .B1(n16141), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16139) );
  AOI22_X1 U19283 ( .A1(n16137), .A2(n16144), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16136), .ZN(n16138) );
  OAI211_X1 U19284 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n16140), .A(
        n16139), .B(n16138), .ZN(P1_U3024) );
  INV_X1 U19285 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16148) );
  AOI22_X1 U19286 ( .A1(n19894), .A2(n16142), .B1(n16141), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n16147) );
  AOI22_X1 U19287 ( .A1(n16145), .A2(n16144), .B1(n16143), .B2(n16148), .ZN(
        n16146) );
  OAI211_X1 U19288 ( .C1(n16149), .C2(n16148), .A(n16147), .B(n16146), .ZN(
        P1_U3025) );
  NAND3_X1 U19289 ( .A1(n16152), .A2(n16151), .A3(n16150), .ZN(n16153) );
  OAI21_X1 U19290 ( .B1(n16155), .B2(n16154), .A(n16153), .ZN(P1_U3468) );
  NAND4_X1 U19291 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20752), .A4(n20760), .ZN(n16156) );
  NAND2_X1 U19292 ( .A1(n16157), .A2(n16156), .ZN(n20659) );
  OAI21_X1 U19293 ( .B1(n16159), .B2(n20659), .A(n16158), .ZN(n16160) );
  OAI221_X1 U19294 ( .B1(n20755), .B2(n20493), .C1(n20755), .C2(n20760), .A(
        n16160), .ZN(n16161) );
  AOI221_X1 U19295 ( .B1(n16162), .B2(n13902), .C1(n20756), .C2(n13902), .A(
        n16161), .ZN(P1_U3162) );
  NOR2_X1 U19296 ( .A1(n16162), .A2(n20756), .ZN(n16164) );
  OAI22_X1 U19297 ( .A1(n20493), .A2(n16164), .B1(n16163), .B2(n20756), .ZN(
        P1_U3466) );
  XNOR2_X1 U19298 ( .A(n16168), .B(n16167), .ZN(n16177) );
  AOI22_X1 U19299 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n18997), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19017), .ZN(n16169) );
  OAI21_X1 U19300 ( .B1(n16170), .B2(n18984), .A(n16169), .ZN(n16171) );
  AOI21_X1 U19301 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n19018), .A(n16171), .ZN(
        n16176) );
  INV_X1 U19302 ( .A(n16172), .ZN(n16174) );
  AOI22_X1 U19303 ( .A1(n16174), .A2(n19020), .B1(n19016), .B2(n16173), .ZN(
        n16175) );
  AOI22_X1 U19304 ( .A1(n16178), .A2(n19022), .B1(P2_REIP_REG_28__SCAN_IN), 
        .B2(n19017), .ZN(n16190) );
  AOI22_X1 U19305 ( .A1(P2_EBX_REG_28__SCAN_IN), .A2(n19018), .B1(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n18997), .ZN(n16189) );
  INV_X1 U19306 ( .A(n16179), .ZN(n16180) );
  OAI22_X1 U19307 ( .A1(n16181), .A2(n19004), .B1(n16180), .B2(n19001), .ZN(
        n16182) );
  INV_X1 U19308 ( .A(n16182), .ZN(n16188) );
  AOI21_X1 U19309 ( .B1(n16185), .B2(n16184), .A(n16183), .ZN(n16186) );
  NAND2_X1 U19310 ( .A1(n18993), .A2(n16186), .ZN(n16187) );
  NAND4_X1 U19311 ( .A1(n16190), .A2(n16189), .A3(n16188), .A4(n16187), .ZN(
        P2_U2827) );
  AOI22_X1 U19312 ( .A1(n16191), .A2(n19022), .B1(P2_REIP_REG_26__SCAN_IN), 
        .B2(n19017), .ZN(n16201) );
  AOI22_X1 U19313 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n19018), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n18997), .ZN(n16200) );
  AOI22_X1 U19314 ( .A1(n16193), .A2(n19020), .B1(n16192), .B2(n19016), .ZN(
        n16199) );
  AOI21_X1 U19315 ( .B1(n16196), .B2(n16195), .A(n16194), .ZN(n16197) );
  NAND2_X1 U19316 ( .A1(n18993), .A2(n16197), .ZN(n16198) );
  NAND4_X1 U19317 ( .A1(n16201), .A2(n16200), .A3(n16199), .A4(n16198), .ZN(
        P2_U2829) );
  AOI22_X1 U19318 ( .A1(n16202), .A2(n19022), .B1(P2_REIP_REG_24__SCAN_IN), 
        .B2(n19017), .ZN(n16212) );
  AOI22_X1 U19319 ( .A1(P2_EBX_REG_24__SCAN_IN), .A2(n19018), .B1(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n18997), .ZN(n16211) );
  OAI22_X1 U19320 ( .A1(n16203), .A2(n19004), .B1(n16213), .B2(n19001), .ZN(
        n16204) );
  INV_X1 U19321 ( .A(n16204), .ZN(n16210) );
  AOI21_X1 U19322 ( .B1(n16207), .B2(n16205), .A(n16206), .ZN(n16208) );
  NAND2_X1 U19323 ( .A1(n18993), .A2(n16208), .ZN(n16209) );
  NAND4_X1 U19324 ( .A1(n16212), .A2(n16211), .A3(n16210), .A4(n16209), .ZN(
        P2_U2831) );
  AOI22_X1 U19325 ( .A1(n19037), .A2(n19062), .B1(n19098), .B2(
        P2_EAX_REG_24__SCAN_IN), .ZN(n16218) );
  AOI22_X1 U19326 ( .A1(n19039), .A2(BUF1_REG_24__SCAN_IN), .B1(n19038), .B2(
        BUF2_REG_24__SCAN_IN), .ZN(n16217) );
  INV_X1 U19327 ( .A(n16213), .ZN(n16214) );
  AOI22_X1 U19328 ( .A1(n16215), .A2(n19086), .B1(n19099), .B2(n16214), .ZN(
        n16216) );
  NAND3_X1 U19329 ( .A1(n16218), .A2(n16217), .A3(n16216), .ZN(P2_U2895) );
  AOI22_X1 U19330 ( .A1(n19037), .A2(n16219), .B1(n19098), .B2(
        P2_EAX_REG_20__SCAN_IN), .ZN(n16224) );
  AOI22_X1 U19331 ( .A1(n19039), .A2(BUF1_REG_20__SCAN_IN), .B1(n19038), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16223) );
  OAI22_X1 U19332 ( .A1(n16220), .A2(n19103), .B1(n19046), .B2(n18873), .ZN(
        n16221) );
  INV_X1 U19333 ( .A(n16221), .ZN(n16222) );
  NAND3_X1 U19334 ( .A1(n16224), .A2(n16223), .A3(n16222), .ZN(P2_U2899) );
  AOI22_X1 U19335 ( .A1(n19037), .A2(n16225), .B1(n19098), .B2(
        P2_EAX_REG_18__SCAN_IN), .ZN(n16230) );
  AOI22_X1 U19336 ( .A1(n19039), .A2(BUF1_REG_18__SCAN_IN), .B1(n19038), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n16229) );
  AOI22_X1 U19337 ( .A1(n16227), .A2(n19099), .B1(n19086), .B2(n16226), .ZN(
        n16228) );
  NAND3_X1 U19338 ( .A1(n16230), .A2(n16229), .A3(n16228), .ZN(P2_U2901) );
  AOI22_X1 U19339 ( .A1(P2_REIP_REG_15__SCAN_IN), .A2(n18902), .B1(n19141), 
        .B2(n16231), .ZN(n16237) );
  INV_X1 U19340 ( .A(n16232), .ZN(n16235) );
  AOI222_X1 U19341 ( .A1(n16235), .A2(n11114), .B1(n19151), .B2(n16234), .C1(
        n16261), .C2(n16233), .ZN(n16236) );
  OAI211_X1 U19342 ( .C1(n16238), .C2(n19154), .A(n16237), .B(n16236), .ZN(
        P2_U2999) );
  AOI22_X1 U19343 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n18902), .B1(n19141), 
        .B2(n16239), .ZN(n16244) );
  AOI222_X1 U19344 ( .A1(n16242), .A2(n16261), .B1(n11114), .B2(n16241), .C1(
        n19151), .C2(n16240), .ZN(n16243) );
  OAI211_X1 U19345 ( .C1(n16245), .C2(n19154), .A(n16244), .B(n16243), .ZN(
        P2_U3001) );
  AOI22_X1 U19346 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n18902), .B1(n19141), 
        .B2(n16246), .ZN(n16251) );
  OAI222_X1 U19347 ( .A1(n18939), .A2(n13862), .B1(n19147), .B2(n16248), .C1(
        n19148), .C2(n16247), .ZN(n16249) );
  INV_X1 U19348 ( .A(n16249), .ZN(n16250) );
  OAI211_X1 U19349 ( .C1(n10776), .C2(n19154), .A(n16251), .B(n16250), .ZN(
        P2_U3003) );
  AOI22_X1 U19350 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n18902), .B1(n19141), 
        .B2(n18963), .ZN(n16265) );
  INV_X1 U19351 ( .A(n18968), .ZN(n16280) );
  XOR2_X1 U19352 ( .A(n16253), .B(n16252), .Z(n16281) );
  INV_X1 U19353 ( .A(n16254), .ZN(n16256) );
  OAI21_X1 U19354 ( .B1(n14266), .B2(n16256), .A(n16255), .ZN(n16260) );
  NAND2_X1 U19355 ( .A1(n10518), .A2(n16258), .ZN(n16259) );
  XNOR2_X1 U19356 ( .A(n16260), .B(n16259), .ZN(n16279) );
  AOI22_X1 U19357 ( .A1(n16281), .A2(n16261), .B1(n11114), .B2(n16279), .ZN(
        n16262) );
  INV_X1 U19358 ( .A(n16262), .ZN(n16263) );
  AOI21_X1 U19359 ( .B1(n19151), .B2(n16280), .A(n16263), .ZN(n16264) );
  OAI211_X1 U19360 ( .C1(n16266), .C2(n19154), .A(n16265), .B(n16264), .ZN(
        P2_U3006) );
  AOI22_X1 U19361 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n18902), .B1(n19141), 
        .B2(n16267), .ZN(n16273) );
  OAI22_X1 U19362 ( .A1(n16269), .A2(n19148), .B1(n19147), .B2(n16268), .ZN(
        n16270) );
  AOI21_X1 U19363 ( .B1(n19151), .B2(n16271), .A(n16270), .ZN(n16272) );
  OAI211_X1 U19364 ( .C1(n16274), .C2(n19154), .A(n16273), .B(n16272), .ZN(
        P2_U3008) );
  AOI21_X1 U19365 ( .B1(n16277), .B2(n16276), .A(n16275), .ZN(n18967) );
  AOI22_X1 U19366 ( .A1(n16278), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16296), .B2(n18967), .ZN(n16287) );
  AOI222_X1 U19367 ( .A1(n16281), .A2(n11175), .B1(n16290), .B2(n16280), .C1(
        n16279), .C2(n19188), .ZN(n16286) );
  NAND2_X1 U19368 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n18902), .ZN(n16285) );
  OAI211_X1 U19369 ( .C1(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n16283), .B(n16282), .ZN(n16284) );
  NAND4_X1 U19370 ( .A1(n16287), .A2(n16286), .A3(n16285), .A4(n16284), .ZN(
        P2_U3038) );
  INV_X1 U19371 ( .A(n19075), .ZN(n19768) );
  AOI21_X1 U19372 ( .B1(n16290), .B2(n16289), .A(n16288), .ZN(n16291) );
  OAI21_X1 U19373 ( .B1(n16292), .B2(n19157), .A(n16291), .ZN(n16295) );
  NOR2_X1 U19374 ( .A1(n16293), .A2(n19174), .ZN(n16294) );
  AOI211_X1 U19375 ( .C1(n19768), .C2(n16296), .A(n16295), .B(n16294), .ZN(
        n16297) );
  OAI221_X1 U19376 ( .B1(n16300), .B2(n16299), .C1(n16300), .C2(n16298), .A(
        n16297), .ZN(P2_U3043) );
  INV_X1 U19377 ( .A(n16340), .ZN(n16305) );
  NAND2_X1 U19378 ( .A1(n16305), .A2(n16301), .ZN(n16302) );
  OAI21_X1 U19379 ( .B1(n16305), .B2(n16314), .A(n16302), .ZN(n16322) );
  OR2_X1 U19380 ( .A1(n16305), .A2(n16303), .ZN(n16307) );
  NAND2_X1 U19381 ( .A1(n16305), .A2(n16304), .ZN(n16306) );
  NAND2_X1 U19382 ( .A1(n16307), .A2(n16306), .ZN(n16316) );
  NAND2_X1 U19383 ( .A1(n16311), .A2(n19793), .ZN(n16309) );
  NAND3_X1 U19384 ( .A1(n16309), .A2(n16308), .A3(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n16310) );
  OAI211_X1 U19385 ( .C1(n19793), .C2(n16311), .A(n16340), .B(n16310), .ZN(
        n16312) );
  INV_X1 U19386 ( .A(n16312), .ZN(n16313) );
  OAI21_X1 U19387 ( .B1(n16314), .B2(n19784), .A(n16313), .ZN(n16317) );
  OAI211_X1 U19388 ( .C1(n16322), .C2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n16316), .B(n16317), .ZN(n16315) );
  NAND2_X1 U19389 ( .A1(n16315), .A2(n19775), .ZN(n16320) );
  INV_X1 U19390 ( .A(n16316), .ZN(n16343) );
  INV_X1 U19391 ( .A(n16317), .ZN(n16318) );
  NAND2_X1 U19392 ( .A1(n16343), .A2(n16318), .ZN(n16319) );
  NAND2_X1 U19393 ( .A1(n16320), .A2(n16319), .ZN(n16321) );
  NAND2_X1 U19394 ( .A1(n16321), .A2(n15807), .ZN(n16345) );
  INV_X1 U19395 ( .A(n16322), .ZN(n16342) );
  INV_X1 U19396 ( .A(n16323), .ZN(n16332) );
  INV_X1 U19397 ( .A(n16324), .ZN(n16331) );
  OR2_X1 U19398 ( .A1(n16328), .A2(n16325), .ZN(n16330) );
  INV_X1 U19399 ( .A(n16326), .ZN(n16327) );
  NAND2_X1 U19400 ( .A1(n16328), .A2(n16327), .ZN(n16329) );
  OAI211_X1 U19401 ( .C1(n16332), .C2(n16331), .A(n16330), .B(n16329), .ZN(
        n19813) );
  OAI21_X1 U19402 ( .B1(P2_MORE_REG_SCAN_IN), .B2(P2_FLUSH_REG_SCAN_IN), .A(
        n16333), .ZN(n16336) );
  AOI22_X1 U19403 ( .A1(n16334), .A2(n19829), .B1(n10683), .B2(n19823), .ZN(
        n16335) );
  NAND2_X1 U19404 ( .A1(n16336), .A2(n16335), .ZN(n16337) );
  NOR2_X1 U19405 ( .A1(n19813), .A2(n16337), .ZN(n16338) );
  OAI21_X1 U19406 ( .B1(n16340), .B2(n16339), .A(n16338), .ZN(n16341) );
  AOI21_X1 U19407 ( .B1(n16343), .B2(n16342), .A(n16341), .ZN(n16344) );
  AND2_X1 U19408 ( .A1(n16345), .A2(n16344), .ZN(n16362) );
  AOI211_X1 U19409 ( .C1(n10069), .C2(n16348), .A(n16347), .B(n16346), .ZN(
        n16360) );
  NAND2_X1 U19410 ( .A1(n16362), .A2(n13937), .ZN(n16349) );
  NAND2_X1 U19411 ( .A1(n16349), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n16354) );
  NAND2_X1 U19412 ( .A1(n19818), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16350) );
  AOI21_X1 U19413 ( .B1(n16352), .B2(n16351), .A(n16350), .ZN(n16353) );
  OAI21_X1 U19414 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n16356), .A(n16355), 
        .ZN(n16358) );
  NAND2_X1 U19415 ( .A1(n19679), .A2(n19695), .ZN(n16357) );
  AOI22_X1 U19416 ( .A1(n19679), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n16358), 
        .B2(n16357), .ZN(n16359) );
  OAI211_X1 U19417 ( .C1(n16362), .C2(n16361), .A(n16360), .B(n16359), .ZN(
        P2_U3176) );
  INV_X1 U19418 ( .A(n19679), .ZN(n16364) );
  OAI221_X1 U19419 ( .B1(n19794), .B2(P2_STATE2_REG_0__SCAN_IN), .C1(n19794), 
        .C2(n16364), .A(n16363), .ZN(P2_U3593) );
  INV_X1 U19420 ( .A(n16365), .ZN(n16404) );
  NAND2_X1 U19421 ( .A1(n16404), .A2(n17540), .ZN(n17490) );
  OAI221_X1 U19422 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16369), .C1(
        n16540), .C2(n16368), .A(n16367), .ZN(n16370) );
  AOI21_X1 U19423 ( .B1(n17675), .B2(n16539), .A(n16370), .ZN(n16376) );
  NAND2_X1 U19424 ( .A1(n17815), .A2(n16371), .ZN(n16381) );
  OAI21_X1 U19425 ( .B1(n16372), .B2(n17734), .A(n16381), .ZN(n16374) );
  AOI22_X1 U19426 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16374), .B1(
        n17731), .B2(n16373), .ZN(n16375) );
  OAI211_X1 U19427 ( .C1(n16377), .C2(n17490), .A(n16376), .B(n16375), .ZN(
        P3_U2800) );
  OAI21_X1 U19428 ( .B1(n16378), .B2(n18264), .A(n16550), .ZN(n16379) );
  AOI22_X1 U19429 ( .A1(n18100), .A2(P3_REIP_REG_29__SCAN_IN), .B1(n16380), 
        .B2(n16379), .ZN(n16391) );
  AOI21_X1 U19430 ( .B1(n16383), .B2(n16382), .A(n16381), .ZN(n16384) );
  AOI21_X1 U19431 ( .B1(n16385), .B2(n17731), .A(n16384), .ZN(n16390) );
  OAI211_X1 U19432 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16415), .A(
        n17690), .B(n16386), .ZN(n16389) );
  OAI21_X1 U19433 ( .B1(n16387), .B2(n17675), .A(n16549), .ZN(n16388) );
  NAND4_X1 U19434 ( .A1(n16391), .A2(n16390), .A3(n16389), .A4(n16388), .ZN(
        P3_U2801) );
  INV_X1 U19435 ( .A(n18138), .ZN(n18090) );
  AND3_X1 U19436 ( .A1(n18772), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n16392), .ZN(n16398) );
  OAI22_X1 U19437 ( .A1(n18772), .A2(n16394), .B1(n16393), .B2(n18127), .ZN(
        n16395) );
  AOI211_X1 U19438 ( .C1(n16398), .C2(n16397), .A(n16396), .B(n16395), .ZN(
        n16401) );
  INV_X1 U19439 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18746) );
  NOR2_X1 U19440 ( .A1(n16409), .A2(n18600), .ZN(n18015) );
  INV_X1 U19441 ( .A(n18015), .ZN(n17884) );
  OAI22_X1 U19442 ( .A1(n18016), .A2(n17995), .B1(n18014), .B2(n17884), .ZN(
        n17935) );
  AOI21_X1 U19443 ( .B1(n17936), .B2(n17935), .A(n16403), .ZN(n17878) );
  INV_X1 U19444 ( .A(n17878), .ZN(n17895) );
  NAND2_X1 U19445 ( .A1(n17895), .A2(n18125), .ZN(n17920) );
  NOR2_X1 U19446 ( .A1(n17877), .A2(n17920), .ZN(n17865) );
  NAND2_X1 U19447 ( .A1(n16404), .A2(n17865), .ZN(n17828) );
  NAND2_X1 U19448 ( .A1(n17466), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17479) );
  OAI22_X1 U19449 ( .A1(n18141), .A2(n18746), .B1(n17828), .B2(n17479), .ZN(
        n16405) );
  INV_X1 U19450 ( .A(n16405), .ZN(n16421) );
  AOI21_X1 U19451 ( .B1(n17730), .B2(n17480), .A(n16407), .ZN(n16408) );
  NAND3_X1 U19452 ( .A1(n18140), .A2(n16406), .A3(n16408), .ZN(n16420) );
  INV_X1 U19453 ( .A(n16407), .ZN(n17481) );
  OAI22_X1 U19454 ( .A1(n17656), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B1(
        n17466), .B2(n17730), .ZN(n17475) );
  OR3_X1 U19455 ( .A1(n17481), .A2(n18043), .A3(n17475), .ZN(n16419) );
  INV_X1 U19456 ( .A(n16408), .ZN(n17476) );
  NAND2_X1 U19457 ( .A1(n17476), .A2(n17475), .ZN(n17474) );
  NAND3_X1 U19458 ( .A1(n16410), .A2(n16409), .A3(n17474), .ZN(n16412) );
  OAI211_X1 U19459 ( .C1(n16413), .C2(n16412), .A(n16411), .B(n18126), .ZN(
        n16417) );
  OAI22_X1 U19460 ( .A1(n16415), .A2(n17884), .B1(n16414), .B2(n17995), .ZN(
        n16416) );
  OAI211_X1 U19461 ( .C1(n16417), .C2(n16416), .A(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .B(n18141), .ZN(n16418) );
  NAND4_X1 U19462 ( .A1(n16421), .A2(n16420), .A3(n16419), .A4(n16418), .ZN(
        P3_U2834) );
  NOR3_X1 U19463 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16423) );
  NOR4_X1 U19464 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16422) );
  NAND4_X1 U19465 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16423), .A3(n16422), .A4(
        U215), .ZN(U213) );
  INV_X1 U19466 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n16509) );
  INV_X2 U19467 ( .A(U214), .ZN(n20926) );
  NOR2_X1 U19468 ( .A1(n20926), .A2(n16424), .ZN(n20927) );
  INV_X1 U19469 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16510) );
  OAI222_X1 U19470 ( .A1(U212), .A2(n16509), .B1(n16472), .B2(n16425), .C1(
        U214), .C2(n16510), .ZN(U216) );
  INV_X1 U19471 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n16427) );
  AOI22_X1 U19472 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n20926), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n20925), .ZN(n16426) );
  OAI21_X1 U19473 ( .B1(n16427), .B2(n16472), .A(n16426), .ZN(U217) );
  INV_X1 U19474 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16429) );
  AOI22_X1 U19475 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n20926), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n20925), .ZN(n16428) );
  OAI21_X1 U19476 ( .B1(n16429), .B2(n16472), .A(n16428), .ZN(U218) );
  AOI22_X1 U19477 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n20926), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n20925), .ZN(n16430) );
  OAI21_X1 U19478 ( .B1(n16431), .B2(n16472), .A(n16430), .ZN(U219) );
  AOI22_X1 U19479 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n20926), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n20925), .ZN(n16432) );
  OAI21_X1 U19480 ( .B1(n15183), .B2(n16472), .A(n16432), .ZN(U220) );
  INV_X1 U19481 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16434) );
  AOI22_X1 U19482 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n20926), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n20925), .ZN(n16433) );
  OAI21_X1 U19483 ( .B1(n16434), .B2(n16472), .A(n16433), .ZN(U221) );
  AOI22_X1 U19484 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n20926), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n20925), .ZN(n16435) );
  OAI21_X1 U19485 ( .B1(n15199), .B2(n16472), .A(n16435), .ZN(U222) );
  AOI22_X1 U19486 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n20926), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n20925), .ZN(n16436) );
  OAI21_X1 U19487 ( .B1(n16437), .B2(n16472), .A(n16436), .ZN(U223) );
  AOI22_X1 U19488 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n20926), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n20925), .ZN(n16438) );
  OAI21_X1 U19489 ( .B1(n15209), .B2(n16472), .A(n16438), .ZN(U224) );
  AOI22_X1 U19490 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n20926), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n20925), .ZN(n16439) );
  OAI21_X1 U19491 ( .B1(n14341), .B2(n16472), .A(n16439), .ZN(U225) );
  AOI22_X1 U19492 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n20926), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n20925), .ZN(n16440) );
  OAI21_X1 U19493 ( .B1(n14260), .B2(n16472), .A(n16440), .ZN(U226) );
  AOI22_X1 U19494 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n20926), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n20925), .ZN(n16441) );
  OAI21_X1 U19495 ( .B1(n16442), .B2(n16472), .A(n16441), .ZN(U227) );
  AOI22_X1 U19496 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n20926), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n20925), .ZN(n16443) );
  OAI21_X1 U19497 ( .B1(n14221), .B2(n16472), .A(n16443), .ZN(U228) );
  INV_X1 U19498 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16445) );
  AOI22_X1 U19499 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n20926), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n20925), .ZN(n16444) );
  OAI21_X1 U19500 ( .B1(n16445), .B2(n16472), .A(n16444), .ZN(U229) );
  INV_X1 U19501 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n16447) );
  AOI22_X1 U19502 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n20926), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n20925), .ZN(n16446) );
  OAI21_X1 U19503 ( .B1(n16447), .B2(n16472), .A(n16446), .ZN(U230) );
  INV_X1 U19504 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n16449) );
  AOI22_X1 U19505 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n20926), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n20925), .ZN(n16448) );
  OAI21_X1 U19506 ( .B1(n16449), .B2(n16472), .A(n16448), .ZN(U231) );
  INV_X1 U19507 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n16451) );
  AOI22_X1 U19508 ( .A1(BUF1_REG_15__SCAN_IN), .A2(n20927), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n20926), .ZN(n16450) );
  OAI21_X1 U19509 ( .B1(n16451), .B2(U212), .A(n16450), .ZN(U232) );
  INV_X1 U19510 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n16453) );
  AOI22_X1 U19511 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n20927), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n20926), .ZN(n16452) );
  OAI21_X1 U19512 ( .B1(n16453), .B2(U212), .A(n16452), .ZN(U233) );
  INV_X1 U19513 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16487) );
  AOI22_X1 U19514 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n20927), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n20926), .ZN(n16454) );
  OAI21_X1 U19515 ( .B1(n16487), .B2(U212), .A(n16454), .ZN(U234) );
  INV_X1 U19516 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16456) );
  AOI22_X1 U19517 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n20927), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n20926), .ZN(n16455) );
  OAI21_X1 U19518 ( .B1(n16456), .B2(U212), .A(n16455), .ZN(U236) );
  AOI22_X1 U19519 ( .A1(P1_DATAO_REG_10__SCAN_IN), .A2(n20926), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n20925), .ZN(n16457) );
  OAI21_X1 U19520 ( .B1(n16458), .B2(n16472), .A(n16457), .ZN(U237) );
  INV_X1 U19521 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n16483) );
  AOI22_X1 U19522 ( .A1(BUF1_REG_9__SCAN_IN), .A2(n20927), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n20926), .ZN(n16459) );
  OAI21_X1 U19523 ( .B1(n16483), .B2(U212), .A(n16459), .ZN(U238) );
  AOI22_X1 U19524 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n20926), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n20925), .ZN(n16460) );
  OAI21_X1 U19525 ( .B1(n16461), .B2(n16472), .A(n16460), .ZN(U239) );
  INV_X1 U19526 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16481) );
  AOI22_X1 U19527 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n20927), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n20926), .ZN(n16462) );
  OAI21_X1 U19528 ( .B1(n16481), .B2(U212), .A(n16462), .ZN(U240) );
  INV_X1 U19529 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16480) );
  AOI22_X1 U19530 ( .A1(BUF1_REG_6__SCAN_IN), .A2(n20927), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n20926), .ZN(n16463) );
  OAI21_X1 U19531 ( .B1(n16480), .B2(U212), .A(n16463), .ZN(U241) );
  INV_X1 U19532 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n16479) );
  AOI22_X1 U19533 ( .A1(BUF1_REG_5__SCAN_IN), .A2(n20927), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n20926), .ZN(n16464) );
  OAI21_X1 U19534 ( .B1(n16479), .B2(U212), .A(n16464), .ZN(U242) );
  INV_X1 U19535 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16466) );
  AOI22_X1 U19536 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n20926), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n20925), .ZN(n16465) );
  OAI21_X1 U19537 ( .B1(n16466), .B2(n16472), .A(n16465), .ZN(U243) );
  INV_X1 U19538 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16477) );
  AOI22_X1 U19539 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n20927), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n20926), .ZN(n16467) );
  OAI21_X1 U19540 ( .B1(n16477), .B2(U212), .A(n16467), .ZN(U244) );
  INV_X1 U19541 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16469) );
  AOI22_X1 U19542 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n20926), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n20925), .ZN(n16468) );
  OAI21_X1 U19543 ( .B1(n16469), .B2(n16472), .A(n16468), .ZN(U245) );
  INV_X1 U19544 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n16475) );
  AOI22_X1 U19545 ( .A1(BUF1_REG_1__SCAN_IN), .A2(n20927), .B1(
        P1_DATAO_REG_1__SCAN_IN), .B2(n20926), .ZN(n16470) );
  OAI21_X1 U19546 ( .B1(n16475), .B2(U212), .A(n16470), .ZN(U246) );
  INV_X1 U19547 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16473) );
  AOI22_X1 U19548 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n20926), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n20925), .ZN(n16471) );
  OAI21_X1 U19549 ( .B1(n16473), .B2(n16472), .A(n16471), .ZN(U247) );
  OAI22_X1 U19550 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16507), .ZN(n16474) );
  INV_X1 U19551 ( .A(n16474), .ZN(U251) );
  INV_X1 U19552 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n20810) );
  AOI22_X1 U19553 ( .A1(n16507), .A2(n16475), .B1(n20810), .B2(U215), .ZN(U252) );
  OAI22_X1 U19554 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16497), .ZN(n16476) );
  INV_X1 U19555 ( .A(n16476), .ZN(U253) );
  INV_X1 U19556 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18172) );
  AOI22_X1 U19557 ( .A1(n16507), .A2(n16477), .B1(n18172), .B2(U215), .ZN(U254) );
  OAI22_X1 U19558 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16497), .ZN(n16478) );
  INV_X1 U19559 ( .A(n16478), .ZN(U255) );
  INV_X1 U19560 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18181) );
  AOI22_X1 U19561 ( .A1(n16507), .A2(n16479), .B1(n18181), .B2(U215), .ZN(U256) );
  INV_X1 U19562 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18186) );
  AOI22_X1 U19563 ( .A1(n16507), .A2(n16480), .B1(n18186), .B2(U215), .ZN(U257) );
  INV_X1 U19564 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18190) );
  AOI22_X1 U19565 ( .A1(n16507), .A2(n16481), .B1(n18190), .B2(U215), .ZN(U258) );
  OAI22_X1 U19566 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16497), .ZN(n16482) );
  INV_X1 U19567 ( .A(n16482), .ZN(U259) );
  INV_X1 U19568 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17446) );
  AOI22_X1 U19569 ( .A1(n16507), .A2(n16483), .B1(n17446), .B2(U215), .ZN(U260) );
  OAI22_X1 U19570 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16497), .ZN(n16484) );
  INV_X1 U19571 ( .A(n16484), .ZN(U261) );
  OAI22_X1 U19572 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16497), .ZN(n16485) );
  INV_X1 U19573 ( .A(n16485), .ZN(U262) );
  OAI22_X1 U19574 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16497), .ZN(n16486) );
  INV_X1 U19575 ( .A(n16486), .ZN(U263) );
  INV_X1 U19576 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n20825) );
  AOI22_X1 U19577 ( .A1(n16507), .A2(n16487), .B1(n20825), .B2(U215), .ZN(U264) );
  OAI22_X1 U19578 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16497), .ZN(n16488) );
  INV_X1 U19579 ( .A(n16488), .ZN(U265) );
  OAI22_X1 U19580 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16507), .ZN(n16489) );
  INV_X1 U19581 ( .A(n16489), .ZN(U266) );
  OAI22_X1 U19582 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16497), .ZN(n16490) );
  INV_X1 U19583 ( .A(n16490), .ZN(U267) );
  OAI22_X1 U19584 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16507), .ZN(n16491) );
  INV_X1 U19585 ( .A(n16491), .ZN(U268) );
  OAI22_X1 U19586 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16497), .ZN(n16492) );
  INV_X1 U19587 ( .A(n16492), .ZN(U269) );
  OAI22_X1 U19588 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16507), .ZN(n16493) );
  INV_X1 U19589 ( .A(n16493), .ZN(U270) );
  OAI22_X1 U19590 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16507), .ZN(n16494) );
  INV_X1 U19591 ( .A(n16494), .ZN(U271) );
  OAI22_X1 U19592 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16507), .ZN(n16495) );
  INV_X1 U19593 ( .A(n16495), .ZN(U272) );
  OAI22_X1 U19594 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16507), .ZN(n16496) );
  INV_X1 U19595 ( .A(n16496), .ZN(U273) );
  OAI22_X1 U19596 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16497), .ZN(n16498) );
  INV_X1 U19597 ( .A(n16498), .ZN(U274) );
  OAI22_X1 U19598 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16507), .ZN(n16499) );
  INV_X1 U19599 ( .A(n16499), .ZN(U275) );
  OAI22_X1 U19600 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16507), .ZN(n16500) );
  INV_X1 U19601 ( .A(n16500), .ZN(U276) );
  OAI22_X1 U19602 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16507), .ZN(n16501) );
  INV_X1 U19603 ( .A(n16501), .ZN(U277) );
  OAI22_X1 U19604 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16507), .ZN(n16502) );
  INV_X1 U19605 ( .A(n16502), .ZN(U278) );
  OAI22_X1 U19606 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16507), .ZN(n16503) );
  INV_X1 U19607 ( .A(n16503), .ZN(U279) );
  OAI22_X1 U19608 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16507), .ZN(n16504) );
  INV_X1 U19609 ( .A(n16504), .ZN(U280) );
  OAI22_X1 U19610 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16507), .ZN(n16505) );
  INV_X1 U19611 ( .A(n16505), .ZN(U281) );
  AOI22_X1 U19612 ( .A1(n16507), .A2(n16509), .B1(n16506), .B2(U215), .ZN(U282) );
  INV_X1 U19613 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16508) );
  AOI222_X1 U19614 ( .A1(n16510), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n16509), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16508), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16511) );
  INV_X2 U19615 ( .A(n16513), .ZN(n16512) );
  INV_X1 U19616 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18709) );
  AOI22_X1 U19617 ( .A1(n16512), .A2(n18709), .B1(n19719), .B2(n16513), .ZN(
        U347) );
  INV_X1 U19618 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18707) );
  INV_X1 U19619 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19717) );
  AOI22_X1 U19620 ( .A1(n16512), .A2(n18707), .B1(n19717), .B2(n16513), .ZN(
        U348) );
  INV_X1 U19621 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18704) );
  INV_X1 U19622 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19715) );
  AOI22_X1 U19623 ( .A1(n16512), .A2(n18704), .B1(n19715), .B2(n16513), .ZN(
        U349) );
  INV_X1 U19624 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18703) );
  INV_X1 U19625 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19713) );
  AOI22_X1 U19626 ( .A1(n16512), .A2(n18703), .B1(n19713), .B2(n16513), .ZN(
        U350) );
  INV_X1 U19627 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18701) );
  INV_X1 U19628 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n19711) );
  AOI22_X1 U19629 ( .A1(n16512), .A2(n18701), .B1(n19711), .B2(n16513), .ZN(
        U351) );
  INV_X1 U19630 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18699) );
  INV_X1 U19631 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19709) );
  AOI22_X1 U19632 ( .A1(n16512), .A2(n18699), .B1(n19709), .B2(n16513), .ZN(
        U352) );
  INV_X1 U19633 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18697) );
  INV_X1 U19634 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19707) );
  AOI22_X1 U19635 ( .A1(n16512), .A2(n18697), .B1(n19707), .B2(n16513), .ZN(
        U353) );
  INV_X1 U19636 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18695) );
  INV_X1 U19637 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19705) );
  AOI22_X1 U19638 ( .A1(n16512), .A2(n18695), .B1(n19705), .B2(n16513), .ZN(
        U354) );
  INV_X1 U19639 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18750) );
  INV_X1 U19640 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19753) );
  AOI22_X1 U19641 ( .A1(n16512), .A2(n18750), .B1(n19753), .B2(n16513), .ZN(
        U355) );
  INV_X1 U19642 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18748) );
  INV_X1 U19643 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19749) );
  AOI22_X1 U19644 ( .A1(n16512), .A2(n18748), .B1(n19749), .B2(n16513), .ZN(
        U356) );
  INV_X1 U19645 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18745) );
  INV_X1 U19646 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19747) );
  AOI22_X1 U19647 ( .A1(n16512), .A2(n18745), .B1(n19747), .B2(n16513), .ZN(
        U357) );
  INV_X1 U19648 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18744) );
  INV_X1 U19649 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19745) );
  AOI22_X1 U19650 ( .A1(n16512), .A2(n18744), .B1(n19745), .B2(n16513), .ZN(
        U358) );
  INV_X1 U19651 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18742) );
  INV_X1 U19652 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19744) );
  AOI22_X1 U19653 ( .A1(n16512), .A2(n18742), .B1(n19744), .B2(n16513), .ZN(
        U359) );
  INV_X1 U19654 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18740) );
  INV_X1 U19655 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19742) );
  AOI22_X1 U19656 ( .A1(n16512), .A2(n18740), .B1(n19742), .B2(n16513), .ZN(
        U360) );
  INV_X1 U19657 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18737) );
  INV_X1 U19658 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19740) );
  AOI22_X1 U19659 ( .A1(n16512), .A2(n18737), .B1(n19740), .B2(n16513), .ZN(
        U361) );
  INV_X1 U19660 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18735) );
  INV_X1 U19661 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19738) );
  AOI22_X1 U19662 ( .A1(n16512), .A2(n18735), .B1(n19738), .B2(n16513), .ZN(
        U362) );
  INV_X1 U19663 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18733) );
  INV_X1 U19664 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19736) );
  AOI22_X1 U19665 ( .A1(n16512), .A2(n18733), .B1(n19736), .B2(n16513), .ZN(
        U363) );
  INV_X1 U19666 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18731) );
  INV_X1 U19667 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19734) );
  AOI22_X1 U19668 ( .A1(n16512), .A2(n18731), .B1(n19734), .B2(n16513), .ZN(
        U364) );
  INV_X1 U19669 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18693) );
  INV_X1 U19670 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19703) );
  AOI22_X1 U19671 ( .A1(n16512), .A2(n18693), .B1(n19703), .B2(n16513), .ZN(
        U365) );
  INV_X1 U19672 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18728) );
  INV_X1 U19673 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19732) );
  AOI22_X1 U19674 ( .A1(n16512), .A2(n18728), .B1(n19732), .B2(n16513), .ZN(
        U366) );
  INV_X1 U19675 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18727) );
  INV_X1 U19676 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19731) );
  AOI22_X1 U19677 ( .A1(n16512), .A2(n18727), .B1(n19731), .B2(n16513), .ZN(
        U367) );
  INV_X1 U19678 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18725) );
  INV_X1 U19679 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19730) );
  AOI22_X1 U19680 ( .A1(n16512), .A2(n18725), .B1(n19730), .B2(n16513), .ZN(
        U368) );
  INV_X1 U19681 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18722) );
  INV_X1 U19682 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19728) );
  AOI22_X1 U19683 ( .A1(n16512), .A2(n18722), .B1(n19728), .B2(n16513), .ZN(
        U369) );
  INV_X1 U19684 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18721) );
  INV_X1 U19685 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19726) );
  AOI22_X1 U19686 ( .A1(n16512), .A2(n18721), .B1(n19726), .B2(n16513), .ZN(
        U370) );
  INV_X1 U19687 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18719) );
  INV_X1 U19688 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19725) );
  AOI22_X1 U19689 ( .A1(n16512), .A2(n18719), .B1(n19725), .B2(n16513), .ZN(
        U371) );
  INV_X1 U19690 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18716) );
  INV_X1 U19691 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19723) );
  AOI22_X1 U19692 ( .A1(n16512), .A2(n18716), .B1(n19723), .B2(n16513), .ZN(
        U372) );
  INV_X1 U19693 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18715) );
  INV_X1 U19694 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19722) );
  AOI22_X1 U19695 ( .A1(n16512), .A2(n18715), .B1(n19722), .B2(n16513), .ZN(
        U373) );
  INV_X1 U19696 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18713) );
  INV_X1 U19697 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19721) );
  AOI22_X1 U19698 ( .A1(n16512), .A2(n18713), .B1(n19721), .B2(n16513), .ZN(
        U374) );
  INV_X1 U19699 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18711) );
  INV_X1 U19700 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19720) );
  AOI22_X1 U19701 ( .A1(n16512), .A2(n18711), .B1(n19720), .B2(n16513), .ZN(
        U375) );
  INV_X1 U19702 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18691) );
  INV_X1 U19703 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19701) );
  AOI22_X1 U19704 ( .A1(n16512), .A2(n18691), .B1(n19701), .B2(n16513), .ZN(
        U376) );
  INV_X1 U19705 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18690) );
  NAND2_X1 U19706 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18690), .ZN(n18677) );
  AOI22_X1 U19707 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18677), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18688), .ZN(n18760) );
  AOI21_X1 U19708 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18760), .ZN(n16514) );
  INV_X1 U19709 ( .A(n16514), .ZN(P3_U2633) );
  NAND2_X1 U19710 ( .A1(n18661), .A2(n18763), .ZN(n16517) );
  INV_X1 U19711 ( .A(n16520), .ZN(n16515) );
  OAI21_X1 U19712 ( .B1(n16515), .B2(n17355), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16516) );
  OAI21_X1 U19713 ( .B1(n16517), .B2(n18664), .A(n16516), .ZN(P3_U2634) );
  AOI21_X1 U19714 ( .B1(n18688), .B2(n18690), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16518) );
  AOI22_X1 U19715 ( .A1(n18822), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16518), 
        .B2(n18823), .ZN(P3_U2635) );
  NOR2_X1 U19716 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18673) );
  OAI21_X1 U19717 ( .B1(n18673), .B2(BS16), .A(n18760), .ZN(n18758) );
  OAI21_X1 U19718 ( .B1(n18760), .B2(n18813), .A(n18758), .ZN(P3_U2636) );
  AND3_X1 U19719 ( .A1(n16520), .A2(n18596), .A3(n16519), .ZN(n18601) );
  NOR2_X1 U19720 ( .A1(n18601), .A2(n18811), .ZN(n18804) );
  OAI21_X1 U19721 ( .B1(n18804), .B2(n18147), .A(n16521), .ZN(P3_U2637) );
  NOR4_X1 U19722 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16525) );
  NOR4_X1 U19723 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16524) );
  NOR4_X1 U19724 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16523) );
  NOR4_X1 U19725 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16522) );
  NAND4_X1 U19726 ( .A1(n16525), .A2(n16524), .A3(n16523), .A4(n16522), .ZN(
        n16531) );
  NOR4_X1 U19727 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_3__SCAN_IN), .A3(P3_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_5__SCAN_IN), .ZN(n16529) );
  AOI211_X1 U19728 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_14__SCAN_IN), .B(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16528) );
  NOR4_X1 U19729 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16527) );
  NOR4_X1 U19730 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_7__SCAN_IN), .A3(P3_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_9__SCAN_IN), .ZN(n16526) );
  NAND4_X1 U19731 ( .A1(n16529), .A2(n16528), .A3(n16527), .A4(n16526), .ZN(
        n16530) );
  NOR2_X1 U19732 ( .A1(n16531), .A2(n16530), .ZN(n18802) );
  INV_X1 U19733 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16533) );
  NOR3_X1 U19734 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16534) );
  OAI21_X1 U19735 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16534), .A(n18802), .ZN(
        n16532) );
  OAI21_X1 U19736 ( .B1(n18802), .B2(n16533), .A(n16532), .ZN(P3_U2638) );
  INV_X1 U19737 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18796) );
  INV_X1 U19738 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18759) );
  AOI21_X1 U19739 ( .B1(n18796), .B2(n18759), .A(n16534), .ZN(n16536) );
  INV_X1 U19740 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16535) );
  INV_X1 U19741 ( .A(n18802), .ZN(n18799) );
  AOI22_X1 U19742 ( .A1(n18802), .A2(n16536), .B1(n16535), .B2(n18799), .ZN(
        P3_U2639) );
  NAND2_X1 U19743 ( .A1(n16848), .A2(n16537), .ZN(n16554) );
  XOR2_X1 U19744 ( .A(n16539), .B(n16538), .Z(n16543) );
  INV_X1 U19745 ( .A(n18667), .ZN(n16865) );
  OAI22_X1 U19746 ( .A1(n16558), .A2(n18751), .B1(n16540), .B2(n16875), .ZN(
        n16541) );
  OAI21_X1 U19747 ( .B1(n16883), .B2(n16544), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16545) );
  OAI211_X1 U19748 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16554), .A(n16546), .B(
        n16545), .ZN(P3_U2641) );
  INV_X1 U19749 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18747) );
  AOI211_X1 U19750 ( .C1(n16549), .C2(n16547), .A(n16548), .B(n18667), .ZN(
        n16553) );
  NAND2_X1 U19751 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n16559), .ZN(n16551) );
  OAI22_X1 U19752 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16551), .B1(n16550), 
        .B2(n16875), .ZN(n16552) );
  AOI211_X1 U19753 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16883), .A(n16553), .B(
        n16552), .ZN(n16557) );
  INV_X1 U19754 ( .A(n16554), .ZN(n16555) );
  OAI21_X1 U19755 ( .B1(n16561), .B2(n16934), .A(n16555), .ZN(n16556) );
  OAI211_X1 U19756 ( .C1(n16558), .C2(n18747), .A(n16557), .B(n16556), .ZN(
        P3_U2642) );
  INV_X1 U19757 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16570) );
  AOI22_X1 U19758 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16883), .B1(n16559), 
        .B2(n18746), .ZN(n16569) );
  INV_X1 U19759 ( .A(n16560), .ZN(n16589) );
  OAI21_X1 U19760 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n16573), .A(n16589), 
        .ZN(n16567) );
  AOI211_X1 U19761 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16576), .A(n16561), .B(
        n16887), .ZN(n16566) );
  AOI211_X1 U19762 ( .C1(n16564), .C2(n16563), .A(n16562), .B(n18667), .ZN(
        n16565) );
  AOI211_X1 U19763 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16567), .A(n16566), 
        .B(n16565), .ZN(n16568) );
  OAI211_X1 U19764 ( .C1(n16570), .C2(n16875), .A(n16569), .B(n16568), .ZN(
        P3_U2643) );
  AOI211_X1 U19765 ( .C1(n17483), .C2(n16571), .A(n16572), .B(n18667), .ZN(
        n16575) );
  OAI22_X1 U19766 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16573), .B1(n17487), 
        .B2(n16875), .ZN(n16574) );
  AOI211_X1 U19767 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n16883), .A(n16575), .B(
        n16574), .ZN(n16578) );
  OAI211_X1 U19768 ( .C1(n16580), .C2(n16897), .A(n16848), .B(n16576), .ZN(
        n16577) );
  OAI211_X1 U19769 ( .C1(n16589), .C2(n18743), .A(n16578), .B(n16577), .ZN(
        P3_U2644) );
  NOR2_X1 U19770 ( .A1(n16879), .A2(n16579), .ZN(n16591) );
  AOI21_X1 U19771 ( .B1(P3_REIP_REG_25__SCAN_IN), .B2(n16591), .A(
        P3_REIP_REG_26__SCAN_IN), .ZN(n16590) );
  AOI22_X1 U19772 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16876), .B1(
        n16883), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16588) );
  AOI211_X1 U19773 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16581), .A(n16580), .B(
        n16887), .ZN(n16586) );
  AOI211_X1 U19774 ( .C1(n16584), .C2(n16583), .A(n16582), .B(n18667), .ZN(
        n16585) );
  NOR2_X1 U19775 ( .A1(n16586), .A2(n16585), .ZN(n16587) );
  OAI211_X1 U19776 ( .C1(n16590), .C2(n16589), .A(n16588), .B(n16587), .ZN(
        P3_U2645) );
  INV_X1 U19777 ( .A(n16591), .ZN(n16593) );
  OAI21_X1 U19778 ( .B1(n16605), .B2(n16879), .A(n16891), .ZN(n16620) );
  NOR2_X1 U19779 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16879), .ZN(n16604) );
  NOR2_X1 U19780 ( .A1(n16620), .A2(n16604), .ZN(n16592) );
  MUX2_X1 U19781 ( .A(n16593), .B(n16592), .S(P3_REIP_REG_25__SCAN_IN), .Z(
        n16603) );
  INV_X1 U19782 ( .A(n16594), .ZN(n16595) );
  NAND2_X1 U19783 ( .A1(n16595), .A2(n16848), .ZN(n16606) );
  INV_X1 U19784 ( .A(n16606), .ZN(n16601) );
  OAI21_X1 U19785 ( .B1(n16887), .B2(n16595), .A(n16888), .ZN(n16599) );
  AOI211_X1 U19786 ( .C1(n17509), .C2(n16597), .A(n16596), .B(n18667), .ZN(
        n16598) );
  AOI221_X1 U19787 ( .B1(n16601), .B2(n16600), .C1(n16599), .C2(
        P3_EBX_REG_25__SCAN_IN), .A(n16598), .ZN(n16602) );
  OAI211_X1 U19788 ( .C1(n17507), .C2(n16875), .A(n16603), .B(n16602), .ZN(
        P3_U2646) );
  INV_X1 U19789 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17522) );
  AOI22_X1 U19790 ( .A1(n16883), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16605), 
        .B2(n16604), .ZN(n16613) );
  AOI21_X1 U19791 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n16621), .A(n16606), .ZN(
        n16611) );
  AOI211_X1 U19792 ( .C1(n16609), .C2(n16608), .A(n16607), .B(n18667), .ZN(
        n16610) );
  AOI211_X1 U19793 ( .C1(n16620), .C2(P3_REIP_REG_24__SCAN_IN), .A(n16611), 
        .B(n16610), .ZN(n16612) );
  OAI211_X1 U19794 ( .C1(n17522), .C2(n16875), .A(n16613), .B(n16612), .ZN(
        P3_U2647) );
  NOR2_X1 U19795 ( .A1(n16879), .A2(n16626), .ZN(n16674) );
  INV_X1 U19796 ( .A(n16674), .ZN(n16700) );
  OAI21_X1 U19797 ( .B1(n16614), .B2(n16700), .A(n18734), .ZN(n16619) );
  AOI211_X1 U19798 ( .C1(n17532), .C2(n16616), .A(n16615), .B(n18667), .ZN(
        n16618) );
  OAI22_X1 U19799 ( .A1(n17536), .A2(n16875), .B1(n16888), .B2(n16895), .ZN(
        n16617) );
  AOI211_X1 U19800 ( .C1(n16620), .C2(n16619), .A(n16618), .B(n16617), .ZN(
        n16623) );
  OAI211_X1 U19801 ( .C1(n16624), .C2(n16895), .A(n16848), .B(n16621), .ZN(
        n16622) );
  NAND2_X1 U19802 ( .A1(n16623), .A2(n16622), .ZN(P3_U2648) );
  AOI211_X1 U19803 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16637), .A(n16624), .B(
        n16887), .ZN(n16625) );
  AOI21_X1 U19804 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n16883), .A(n16625), .ZN(
        n16634) );
  NOR2_X1 U19805 ( .A1(n16862), .A2(n16626), .ZN(n16710) );
  AOI21_X1 U19806 ( .B1(n16628), .B2(n16710), .A(n16627), .ZN(n16650) );
  INV_X1 U19807 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18732) );
  INV_X1 U19808 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18730) );
  NAND2_X1 U19809 ( .A1(n16628), .A2(n16674), .ZN(n16643) );
  AOI221_X1 U19810 ( .B1(P3_REIP_REG_22__SCAN_IN), .B2(P3_REIP_REG_21__SCAN_IN), .C1(n18732), .C2(n18730), .A(n16643), .ZN(n16632) );
  AOI211_X1 U19811 ( .C1(n17552), .C2(n16630), .A(n16629), .B(n18667), .ZN(
        n16631) );
  AOI211_X1 U19812 ( .C1(n16650), .C2(P3_REIP_REG_22__SCAN_IN), .A(n16632), 
        .B(n16631), .ZN(n16633) );
  OAI211_X1 U19813 ( .C1(n17549), .C2(n16875), .A(n16634), .B(n16633), .ZN(
        P3_U2649) );
  INV_X1 U19814 ( .A(n16650), .ZN(n16642) );
  AOI211_X1 U19815 ( .C1(n17567), .C2(n16636), .A(n16635), .B(n18667), .ZN(
        n16640) );
  OAI211_X1 U19816 ( .C1(n16644), .C2(n20795), .A(n16848), .B(n16637), .ZN(
        n16638) );
  OAI21_X1 U19817 ( .B1(n20795), .B2(n16888), .A(n16638), .ZN(n16639) );
  AOI211_X1 U19818 ( .C1(n16876), .C2(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(
        n16640), .B(n16639), .ZN(n16641) );
  OAI221_X1 U19819 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n16643), .C1(n18730), 
        .C2(n16642), .A(n16641), .ZN(P3_U2650) );
  AOI211_X1 U19820 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16656), .A(n16644), .B(
        n16887), .ZN(n16645) );
  AOI21_X1 U19821 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16883), .A(n16645), .ZN(
        n16652) );
  NOR3_X1 U19822 ( .A1(n16660), .A2(n16661), .A3(n16700), .ZN(n16649) );
  AOI211_X1 U19823 ( .C1(n17578), .C2(n16647), .A(n16646), .B(n18667), .ZN(
        n16648) );
  AOI221_X1 U19824 ( .B1(n16650), .B2(P3_REIP_REG_20__SCAN_IN), .C1(n16649), 
        .C2(n18729), .A(n16648), .ZN(n16651) );
  OAI211_X1 U19825 ( .C1(n9903), .C2(n16875), .A(n16652), .B(n16651), .ZN(
        P3_U2651) );
  INV_X1 U19826 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18726) );
  INV_X1 U19827 ( .A(n16710), .ZN(n16684) );
  OAI21_X1 U19828 ( .B1(n16660), .B2(n16684), .A(n16889), .ZN(n16677) );
  OAI21_X1 U19829 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16653), .A(
        n17546), .ZN(n17589) );
  INV_X1 U19830 ( .A(n17589), .ZN(n16654) );
  AOI221_X1 U19831 ( .B1(n16655), .B2(n16654), .C1(n16668), .C2(n17589), .A(
        n18667), .ZN(n16659) );
  OAI211_X1 U19832 ( .C1(n16664), .C2(n17011), .A(n16848), .B(n16656), .ZN(
        n16657) );
  OAI211_X1 U19833 ( .C1(n16888), .C2(n17011), .A(n18141), .B(n16657), .ZN(
        n16658) );
  AOI211_X1 U19834 ( .C1(n16876), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16659), .B(n16658), .ZN(n16663) );
  NOR2_X1 U19835 ( .A1(n16660), .A2(n16700), .ZN(n16670) );
  OAI211_X1 U19836 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(P3_REIP_REG_18__SCAN_IN), .A(n16670), .B(n16661), .ZN(n16662) );
  OAI211_X1 U19837 ( .C1(n18726), .C2(n16677), .A(n16663), .B(n16662), .ZN(
        P3_U2652) );
  INV_X1 U19838 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17598) );
  AOI211_X1 U19839 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16680), .A(n16664), .B(
        n16887), .ZN(n16665) );
  AOI211_X1 U19840 ( .C1(n16883), .C2(P3_EBX_REG_18__SCAN_IN), .A(n18135), .B(
        n16665), .ZN(n16673) );
  INV_X1 U19841 ( .A(n16677), .ZN(n16671) );
  INV_X1 U19842 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18724) );
  OAI21_X1 U19843 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17584), .A(
        n16666), .ZN(n17595) );
  AOI211_X1 U19844 ( .C1(n16693), .C2(n17584), .A(n16845), .B(n17595), .ZN(
        n16667) );
  AOI211_X1 U19845 ( .C1(n16668), .C2(n17595), .A(n16667), .B(n18667), .ZN(
        n16669) );
  AOI221_X1 U19846 ( .B1(n16671), .B2(P3_REIP_REG_18__SCAN_IN), .C1(n16670), 
        .C2(n18724), .A(n16669), .ZN(n16672) );
  OAI211_X1 U19847 ( .C1(n17598), .C2(n16875), .A(n16673), .B(n16672), .ZN(
        P3_U2653) );
  INV_X1 U19848 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18720) );
  INV_X1 U19849 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18718) );
  NOR2_X1 U19850 ( .A1(n18720), .A2(n18718), .ZN(n16692) );
  AOI21_X1 U19851 ( .B1(n16692), .B2(n16674), .A(P3_REIP_REG_17__SCAN_IN), 
        .ZN(n16678) );
  AOI21_X1 U19852 ( .B1(n9902), .B2(n16690), .A(n17584), .ZN(n17609) );
  INV_X1 U19853 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16846) );
  NAND2_X1 U19854 ( .A1(n16846), .A2(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n16831) );
  INV_X1 U19855 ( .A(n16831), .ZN(n16866) );
  AOI21_X1 U19856 ( .B1(n17605), .B2(n16866), .A(n16845), .ZN(n16675) );
  XNOR2_X1 U19857 ( .A(n17609), .B(n16675), .ZN(n16676) );
  OAI22_X1 U19858 ( .A1(n16678), .A2(n16677), .B1(n18667), .B2(n16676), .ZN(
        n16679) );
  AOI211_X1 U19859 ( .C1(n16883), .C2(P3_EBX_REG_17__SCAN_IN), .A(n18100), .B(
        n16679), .ZN(n16683) );
  OAI211_X1 U19860 ( .C1(n16685), .C2(n16681), .A(n16848), .B(n16680), .ZN(
        n16682) );
  OAI211_X1 U19861 ( .C1(n16875), .C2(n9902), .A(n16683), .B(n16682), .ZN(
        P3_U2654) );
  NAND2_X1 U19862 ( .A1(n16889), .A2(n16684), .ZN(n16720) );
  AOI211_X1 U19863 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16702), .A(n16685), .B(
        n16887), .ZN(n16688) );
  AOI21_X1 U19864 ( .B1(n16883), .B2(P3_EBX_REG_16__SCAN_IN), .A(n18135), .ZN(
        n16686) );
  INV_X1 U19865 ( .A(n16686), .ZN(n16687) );
  AOI211_X1 U19866 ( .C1(n16876), .C2(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16688), .B(n16687), .ZN(n16698) );
  NOR2_X1 U19867 ( .A1(n16693), .A2(n16689), .ZN(n16701) );
  INV_X1 U19868 ( .A(n16699), .ZN(n16691) );
  OAI21_X1 U19869 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16691), .A(
        n16690), .ZN(n17622) );
  AOI211_X1 U19870 ( .C1(n18720), .C2(n18718), .A(n16692), .B(n16700), .ZN(
        n16696) );
  INV_X1 U19871 ( .A(n16693), .ZN(n16694) );
  AOI211_X1 U19872 ( .C1(n16805), .C2(n16694), .A(n18667), .B(n17622), .ZN(
        n16695) );
  AOI211_X1 U19873 ( .C1(n16701), .C2(n17622), .A(n16696), .B(n16695), .ZN(
        n16697) );
  OAI211_X1 U19874 ( .C1(n18720), .C2(n16720), .A(n16698), .B(n16697), .ZN(
        P3_U2655) );
  OAI21_X1 U19875 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17617), .A(
        n16699), .ZN(n17627) );
  OAI21_X1 U19876 ( .B1(n16845), .B2(n16846), .A(n16865), .ZN(n16886) );
  AOI211_X1 U19877 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n16805), .A(
        n17627), .B(n16886), .ZN(n16708) );
  OAI22_X1 U19878 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16700), .B1(n16888), 
        .B2(n16703), .ZN(n16707) );
  AOI22_X1 U19879 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n16876), .B1(
        n16701), .B2(n17627), .ZN(n16705) );
  OAI211_X1 U19880 ( .C1(n16715), .C2(n16703), .A(n16848), .B(n16702), .ZN(
        n16704) );
  OAI211_X1 U19881 ( .C1(n16720), .C2(n18718), .A(n16705), .B(n16704), .ZN(
        n16706) );
  OR4_X1 U19882 ( .A1(n18135), .A2(n16708), .A3(n16707), .A4(n16706), .ZN(
        P3_U2656) );
  INV_X1 U19883 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18717) );
  INV_X1 U19884 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18714) );
  NAND2_X1 U19885 ( .A1(n16843), .A2(n16709), .ZN(n16733) );
  NOR3_X1 U19886 ( .A1(n16710), .A2(n18714), .A3(n16733), .ZN(n16711) );
  AOI211_X1 U19887 ( .C1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .C2(n16876), .A(
        n18100), .B(n16711), .ZN(n16719) );
  INV_X1 U19888 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17644) );
  NAND2_X1 U19889 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16712), .ZN(
        n16722) );
  AOI21_X1 U19890 ( .B1(n17644), .B2(n16722), .A(n17617), .ZN(n17646) );
  AOI21_X1 U19891 ( .B1(n16712), .B2(n16866), .A(n16845), .ZN(n16730) );
  INV_X1 U19892 ( .A(n17646), .ZN(n16714) );
  INV_X1 U19893 ( .A(n16730), .ZN(n16713) );
  AOI221_X1 U19894 ( .B1(n17646), .B2(n16730), .C1(n16714), .C2(n16713), .A(
        n18667), .ZN(n16717) );
  AOI211_X1 U19895 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16723), .A(n16715), .B(
        n16887), .ZN(n16716) );
  AOI211_X1 U19896 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16883), .A(n16717), .B(
        n16716), .ZN(n16718) );
  OAI211_X1 U19897 ( .C1(n18717), .C2(n16720), .A(n16719), .B(n16718), .ZN(
        P3_U2657) );
  AOI21_X1 U19898 ( .B1(n16843), .B2(n16744), .A(n16862), .ZN(n16749) );
  OAI21_X1 U19899 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n16879), .A(n16749), 
        .ZN(n16729) );
  INV_X1 U19900 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17671) );
  OR2_X1 U19901 ( .A1(n17816), .A2(n17746), .ZN(n16803) );
  NOR2_X1 U19902 ( .A1(n9910), .A2(n16803), .ZN(n16793) );
  NAND2_X1 U19903 ( .A1(n16721), .A2(n16793), .ZN(n17658) );
  NOR2_X1 U19904 ( .A1(n17671), .A2(n17658), .ZN(n16735) );
  OAI21_X1 U19905 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16735), .A(
        n16722), .ZN(n17665) );
  AOI211_X1 U19906 ( .C1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n16805), .A(
        n17665), .B(n16886), .ZN(n16728) );
  AOI22_X1 U19907 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n16876), .B1(
        n16883), .B2(P3_EBX_REG_13__SCAN_IN), .ZN(n16726) );
  OAI211_X1 U19908 ( .C1(n16734), .C2(n16724), .A(n16848), .B(n16723), .ZN(
        n16725) );
  NAND3_X1 U19909 ( .A1(n16726), .A2(n18141), .A3(n16725), .ZN(n16727) );
  AOI211_X1 U19910 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16729), .A(n16728), 
        .B(n16727), .ZN(n16732) );
  NAND3_X1 U19911 ( .A1(n16865), .A2(n16730), .A3(n17665), .ZN(n16731) );
  OAI211_X1 U19912 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16733), .A(n16732), 
        .B(n16731), .ZN(P3_U2658) );
  NAND2_X1 U19913 ( .A1(n16843), .A2(n18712), .ZN(n16743) );
  AOI21_X1 U19914 ( .B1(n16883), .B2(P3_EBX_REG_12__SCAN_IN), .A(n18135), .ZN(
        n16742) );
  AOI211_X1 U19915 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16752), .A(n16734), .B(
        n16887), .ZN(n16740) );
  AOI21_X1 U19916 ( .B1(n17671), .B2(n17658), .A(n16735), .ZN(n17674) );
  INV_X1 U19917 ( .A(n16736), .ZN(n17642) );
  AOI21_X1 U19918 ( .B1(n17642), .B2(n16866), .A(n16845), .ZN(n16737) );
  XNOR2_X1 U19919 ( .A(n17674), .B(n16737), .ZN(n16738) );
  OAI22_X1 U19920 ( .A1(n18667), .A2(n16738), .B1(n18712), .B2(n16749), .ZN(
        n16739) );
  AOI211_X1 U19921 ( .C1(n16876), .C2(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(
        n16740), .B(n16739), .ZN(n16741) );
  OAI211_X1 U19922 ( .C1(n16744), .C2(n16743), .A(n16742), .B(n16741), .ZN(
        P3_U2659) );
  NAND2_X1 U19923 ( .A1(P3_REIP_REG_10__SCAN_IN), .A2(P3_REIP_REG_9__SCAN_IN), 
        .ZN(n16757) );
  INV_X1 U19924 ( .A(n16757), .ZN(n16746) );
  INV_X1 U19925 ( .A(n16745), .ZN(n16785) );
  NOR2_X1 U19926 ( .A1(n16879), .A2(n16785), .ZN(n16773) );
  AOI21_X1 U19927 ( .B1(n16746), .B2(n16773), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16750) );
  INV_X1 U19928 ( .A(n16793), .ZN(n16747) );
  NOR2_X1 U19929 ( .A1(n16764), .A2(n16747), .ZN(n16769) );
  INV_X1 U19930 ( .A(n16769), .ZN(n16762) );
  NOR2_X1 U19931 ( .A1(n16763), .A2(n16762), .ZN(n16761) );
  OAI21_X1 U19932 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16761), .A(
        n17658), .ZN(n17697) );
  AOI21_X1 U19933 ( .B1(n16761), .B2(n16846), .A(n16845), .ZN(n16766) );
  XOR2_X1 U19934 ( .A(n17697), .B(n16766), .Z(n16748) );
  OAI22_X1 U19935 ( .A1(n16750), .A2(n16749), .B1(n18667), .B2(n16748), .ZN(
        n16751) );
  AOI211_X1 U19936 ( .C1(n16883), .C2(P3_EBX_REG_11__SCAN_IN), .A(n18135), .B(
        n16751), .ZN(n16754) );
  OAI211_X1 U19937 ( .C1(n16755), .C2(n17119), .A(n16848), .B(n16752), .ZN(
        n16753) );
  OAI211_X1 U19938 ( .C1(n16875), .C2(n17685), .A(n16754), .B(n16753), .ZN(
        P3_U2660) );
  AOI21_X1 U19939 ( .B1(n16843), .B2(n16785), .A(n16862), .ZN(n16792) );
  INV_X1 U19940 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18708) );
  AOI211_X1 U19941 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16756), .A(n16755), .B(
        n16887), .ZN(n16760) );
  OAI211_X1 U19942 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(P3_REIP_REG_9__SCAN_IN), 
        .A(n16773), .B(n16757), .ZN(n16758) );
  OAI211_X1 U19943 ( .C1(n16763), .C2(n16875), .A(n18141), .B(n16758), .ZN(
        n16759) );
  AOI211_X1 U19944 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16883), .A(n16760), .B(
        n16759), .ZN(n16768) );
  AOI21_X1 U19945 ( .B1(n16763), .B2(n16762), .A(n16761), .ZN(n17706) );
  INV_X1 U19946 ( .A(n17706), .ZN(n16765) );
  AOI21_X1 U19947 ( .B1(n17722), .B2(n16866), .A(n16845), .ZN(n16784) );
  AOI21_X1 U19948 ( .B1(n16805), .B2(n16764), .A(n16784), .ZN(n16771) );
  OAI221_X1 U19949 ( .B1(n17706), .B2(n16766), .C1(n16765), .C2(n16771), .A(
        n16865), .ZN(n16767) );
  OAI211_X1 U19950 ( .C1(n16792), .C2(n18708), .A(n16768), .B(n16767), .ZN(
        P3_U2661) );
  AOI21_X1 U19951 ( .B1(n16848), .B2(n16772), .A(n16883), .ZN(n16779) );
  INV_X1 U19952 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20878) );
  NAND2_X1 U19953 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16793), .ZN(
        n16783) );
  AOI21_X1 U19954 ( .B1(n20878), .B2(n16783), .A(n16769), .ZN(n17716) );
  NAND2_X1 U19955 ( .A1(n20878), .A2(n16846), .ZN(n16770) );
  OAI22_X1 U19956 ( .A1(n17716), .A2(n16771), .B1(n16783), .B2(n16770), .ZN(
        n16777) );
  INV_X1 U19957 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18706) );
  NOR2_X1 U19958 ( .A1(n16772), .A2(n16887), .ZN(n16782) );
  AOI22_X1 U19959 ( .A1(n16773), .A2(n18706), .B1(n16782), .B2(n16780), .ZN(
        n16775) );
  NOR2_X1 U19960 ( .A1(n16805), .A2(n18667), .ZN(n16861) );
  AOI22_X1 U19961 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16876), .B1(
        n17716), .B2(n16861), .ZN(n16774) );
  OAI211_X1 U19962 ( .C1(n16792), .C2(n18706), .A(n16775), .B(n16774), .ZN(
        n16776) );
  AOI211_X1 U19963 ( .C1(n16865), .C2(n16777), .A(n18135), .B(n16776), .ZN(
        n16778) );
  OAI21_X1 U19964 ( .B1(n16780), .B2(n16779), .A(n16778), .ZN(P3_U2662) );
  NAND2_X1 U19965 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16799), .ZN(n16781) );
  AOI22_X1 U19966 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16876), .B1(
        n16782), .B2(n16781), .ZN(n16791) );
  OAI21_X1 U19967 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n16793), .A(
        n16783), .ZN(n17724) );
  XNOR2_X1 U19968 ( .A(n16784), .B(n17724), .ZN(n16789) );
  NAND2_X1 U19969 ( .A1(n16843), .A2(n16785), .ZN(n16786) );
  OAI22_X1 U19970 ( .A1(n16888), .A2(n9828), .B1(n16787), .B2(n16786), .ZN(
        n16788) );
  AOI211_X1 U19971 ( .C1(n16865), .C2(n16789), .A(n18135), .B(n16788), .ZN(
        n16790) );
  OAI211_X1 U19972 ( .C1(n16792), .C2(n18705), .A(n16791), .B(n16790), .ZN(
        P3_U2663) );
  AOI22_X1 U19973 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n16876), .B1(
        n16883), .B2(P3_EBX_REG_7__SCAN_IN), .ZN(n16802) );
  OAI21_X1 U19974 ( .B1(n16794), .B2(n16879), .A(n16891), .ZN(n16812) );
  AOI21_X1 U19975 ( .B1(n9910), .B2(n16803), .A(n16793), .ZN(n17735) );
  OAI21_X1 U19976 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16803), .A(
        n16877), .ZN(n16814) );
  INV_X1 U19977 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18702) );
  NAND3_X1 U19978 ( .A1(n16843), .A2(n16794), .A3(n18702), .ZN(n16797) );
  NOR2_X1 U19979 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16803), .ZN(
        n16795) );
  OAI211_X1 U19980 ( .C1(n16795), .C2(n16845), .A(n16865), .B(n17735), .ZN(
        n16796) );
  OAI211_X1 U19981 ( .C1(n17735), .C2(n16814), .A(n16797), .B(n16796), .ZN(
        n16798) );
  AOI21_X1 U19982 ( .B1(P3_REIP_REG_7__SCAN_IN), .B2(n16812), .A(n16798), .ZN(
        n16801) );
  OAI211_X1 U19983 ( .C1(n16806), .C2(n17121), .A(n16848), .B(n16799), .ZN(
        n16800) );
  NAND4_X1 U19984 ( .A1(n16802), .A2(n16801), .A3(n18141), .A4(n16800), .ZN(
        P3_U2664) );
  NAND2_X1 U19985 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17749), .ZN(
        n16817) );
  INV_X1 U19986 ( .A(n16817), .ZN(n16804) );
  OAI21_X1 U19987 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16804), .A(
        n16803), .ZN(n17753) );
  INV_X1 U19988 ( .A(n17753), .ZN(n16815) );
  OAI21_X1 U19989 ( .B1(n16879), .B2(n16822), .A(n18700), .ZN(n16811) );
  AOI211_X1 U19990 ( .C1(n16805), .C2(n16817), .A(n17753), .B(n16886), .ZN(
        n16810) );
  AOI211_X1 U19991 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16820), .A(n16806), .B(
        n16887), .ZN(n16807) );
  AOI211_X1 U19992 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n16876), .A(
        n18135), .B(n16807), .ZN(n16808) );
  OAI21_X1 U19993 ( .B1(n16888), .B2(n20839), .A(n16808), .ZN(n16809) );
  AOI211_X1 U19994 ( .C1(n16812), .C2(n16811), .A(n16810), .B(n16809), .ZN(
        n16813) );
  OAI21_X1 U19995 ( .B1(n16815), .B2(n16814), .A(n16813), .ZN(P3_U2665) );
  OAI22_X1 U19996 ( .A1(n17765), .A2(n16875), .B1(n16888), .B2(n16821), .ZN(
        n16816) );
  AOI211_X1 U19997 ( .C1(P3_REIP_REG_5__SCAN_IN), .C2(n16862), .A(n18100), .B(
        n16816), .ZN(n16827) );
  NOR2_X1 U19998 ( .A1(n17816), .A2(n17766), .ZN(n16828) );
  OAI21_X1 U19999 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n16828), .A(
        n16817), .ZN(n17771) );
  INV_X1 U20000 ( .A(n17771), .ZN(n16819) );
  AOI21_X1 U20001 ( .B1(n16846), .B2(n16828), .A(n16845), .ZN(n16818) );
  INV_X1 U20002 ( .A(n16818), .ZN(n16832) );
  OAI221_X1 U20003 ( .B1(n16819), .B2(n16818), .C1(n17771), .C2(n16832), .A(
        n16865), .ZN(n16826) );
  OAI211_X1 U20004 ( .C1(n16833), .C2(n16821), .A(n16848), .B(n16820), .ZN(
        n16825) );
  OAI211_X1 U20005 ( .C1(P3_REIP_REG_5__SCAN_IN), .C2(n16823), .A(n16843), .B(
        n16822), .ZN(n16824) );
  NAND4_X1 U20006 ( .A1(n16827), .A2(n16826), .A3(n16825), .A4(n16824), .ZN(
        P3_U2666) );
  AOI21_X1 U20007 ( .B1(n16843), .B2(n16834), .A(n16862), .ZN(n16856) );
  INV_X1 U20008 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n16830) );
  NAND2_X1 U20009 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17782), .ZN(
        n16844) );
  AOI21_X1 U20010 ( .B1(n16830), .B2(n16844), .A(n16828), .ZN(n17783) );
  NAND2_X1 U20011 ( .A1(n18160), .A2(n18806), .ZN(n18829) );
  AOI21_X1 U20012 ( .B1(n9651), .B2(n18604), .A(n18829), .ZN(n16829) );
  AOI211_X1 U20013 ( .C1(n17783), .C2(n16861), .A(n18135), .B(n16829), .ZN(
        n16842) );
  NAND2_X1 U20014 ( .A1(n17782), .A2(n16830), .ZN(n17779) );
  OAI22_X1 U20015 ( .A1(n17783), .A2(n16832), .B1(n16831), .B2(n17779), .ZN(
        n16840) );
  AOI211_X1 U20016 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16847), .A(n16833), .B(
        n16887), .ZN(n16839) );
  AOI22_X1 U20017 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n16876), .B1(
        n16883), .B2(P3_EBX_REG_4__SCAN_IN), .ZN(n16837) );
  INV_X1 U20018 ( .A(n16834), .ZN(n16835) );
  NAND3_X1 U20019 ( .A1(n16843), .A2(n18696), .A3(n16835), .ZN(n16836) );
  NAND2_X1 U20020 ( .A1(n16837), .A2(n16836), .ZN(n16838) );
  AOI211_X1 U20021 ( .C1(n16865), .C2(n16840), .A(n16839), .B(n16838), .ZN(
        n16841) );
  OAI211_X1 U20022 ( .C1(n18696), .C2(n16856), .A(n16842), .B(n16841), .ZN(
        P3_U2667) );
  INV_X1 U20023 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18692) );
  NOR2_X1 U20024 ( .A1(n18796), .A2(n18692), .ZN(n16871) );
  AOI21_X1 U20025 ( .B1(n16843), .B2(n16871), .A(P3_REIP_REG_3__SCAN_IN), .ZN(
        n16857) );
  AOI22_X1 U20026 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n16876), .B1(
        n16883), .B2(P3_EBX_REG_3__SCAN_IN), .ZN(n16855) );
  NOR2_X1 U20027 ( .A1(n17816), .A2(n17811), .ZN(n16860) );
  OAI21_X1 U20028 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n16860), .A(
        n16844), .ZN(n17800) );
  AOI21_X1 U20029 ( .B1(n16860), .B2(n16846), .A(n16845), .ZN(n16864) );
  XNOR2_X1 U20030 ( .A(n17800), .B(n16864), .ZN(n16853) );
  NAND2_X1 U20031 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18612), .ZN(
        n18614) );
  AOI21_X1 U20032 ( .B1(n18768), .B2(n18614), .A(n17125), .ZN(n18764) );
  INV_X1 U20033 ( .A(n18764), .ZN(n16851) );
  OAI211_X1 U20034 ( .C1(n16858), .C2(n16849), .A(n16848), .B(n16847), .ZN(
        n16850) );
  OAI21_X1 U20035 ( .B1(n18829), .B2(n16851), .A(n16850), .ZN(n16852) );
  AOI21_X1 U20036 ( .B1(n16853), .B2(n16865), .A(n16852), .ZN(n16854) );
  OAI211_X1 U20037 ( .C1(n16857), .C2(n16856), .A(n16855), .B(n16854), .ZN(
        P3_U2668) );
  INV_X1 U20038 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17205) );
  INV_X1 U20039 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17199) );
  NAND2_X1 U20040 ( .A1(n17205), .A2(n17199), .ZN(n16859) );
  AOI211_X1 U20041 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16859), .A(n16858), .B(
        n16887), .ZN(n16870) );
  NAND2_X1 U20042 ( .A1(n11361), .A2(n18618), .ZN(n18611) );
  OAI21_X1 U20043 ( .B1(n18621), .B2(n18793), .A(n18611), .ZN(n18774) );
  AOI21_X1 U20044 ( .B1(n17816), .B2(n17811), .A(n16860), .ZN(n16863) );
  AOI22_X1 U20045 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n16862), .B1(n16863), 
        .B2(n16861), .ZN(n16868) );
  INV_X1 U20046 ( .A(n16863), .ZN(n17807) );
  OAI211_X1 U20047 ( .C1(n16866), .C2(n17807), .A(n16865), .B(n16864), .ZN(
        n16867) );
  OAI211_X1 U20048 ( .C1(n18829), .C2(n18774), .A(n16868), .B(n16867), .ZN(
        n16869) );
  AOI211_X1 U20049 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16883), .A(n16870), .B(
        n16869), .ZN(n16874) );
  AOI211_X1 U20050 ( .C1(n18796), .C2(n18692), .A(n16879), .B(n16871), .ZN(
        n16872) );
  INV_X1 U20051 ( .A(n16872), .ZN(n16873) );
  OAI211_X1 U20052 ( .C1(n16875), .C2(n17811), .A(n16874), .B(n16873), .ZN(
        P3_U2669) );
  AOI21_X1 U20053 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16877), .A(
        n16876), .ZN(n16885) );
  NOR2_X1 U20054 ( .A1(n17205), .A2(n17199), .ZN(n17193) );
  AOI21_X1 U20055 ( .B1(n17205), .B2(n17199), .A(n17193), .ZN(n16878) );
  INV_X1 U20056 ( .A(n16878), .ZN(n17200) );
  OAI22_X1 U20057 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16879), .B1(n16887), 
        .B2(n17200), .ZN(n16882) );
  NAND2_X1 U20058 ( .A1(n16880), .A2(n18618), .ZN(n18780) );
  OAI22_X1 U20059 ( .A1(n18796), .A2(n16891), .B1(n18780), .B2(n18829), .ZN(
        n16881) );
  AOI211_X1 U20060 ( .C1(n16883), .C2(P3_EBX_REG_1__SCAN_IN), .A(n16882), .B(
        n16881), .ZN(n16884) );
  OAI221_X1 U20061 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16886), .C1(
        n17816), .C2(n16885), .A(n16884), .ZN(P3_U2670) );
  NAND2_X1 U20062 ( .A1(n16888), .A2(n16887), .ZN(n16890) );
  AOI22_X1 U20063 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n16890), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n16889), .ZN(n16893) );
  NAND3_X1 U20064 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18825), .A3(
        n16891), .ZN(n16892) );
  OAI211_X1 U20065 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18829), .A(
        n16893), .B(n16892), .ZN(P3_U2671) );
  NOR4_X1 U20066 ( .A1(n16896), .A2(n16895), .A3(n16894), .A4(n20795), .ZN(
        n16900) );
  NOR4_X1 U20067 ( .A1(n16934), .A2(n16898), .A3(n16897), .A4(n16981), .ZN(
        n16899) );
  NAND4_X1 U20068 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n16900), .A4(n16899), .ZN(n16903) );
  NAND2_X1 U20069 ( .A1(n17197), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16902) );
  NAND2_X1 U20070 ( .A1(n16930), .A2(n18193), .ZN(n16901) );
  OAI22_X1 U20071 ( .A1(n16930), .A2(n16902), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16901), .ZN(P3_U2672) );
  NAND2_X1 U20072 ( .A1(n16904), .A2(n16903), .ZN(n16905) );
  NAND2_X1 U20073 ( .A1(n16905), .A2(n17197), .ZN(n16929) );
  AOI22_X1 U20074 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17143), .ZN(n16915) );
  AOI22_X1 U20075 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n9607), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16914) );
  AOI22_X1 U20076 ( .A1(n9603), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__7__SCAN_IN), .B2(n17156), .ZN(n16906) );
  OAI21_X1 U20077 ( .B1(n16958), .B2(n17176), .A(n16906), .ZN(n16912) );
  AOI22_X1 U20078 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n9606), .B1(n9605), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16910) );
  AOI22_X1 U20079 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n17160), .B1(
        P3_INSTQUEUE_REG_4__7__SCAN_IN), .B2(n17161), .ZN(n16909) );
  AOI22_X1 U20080 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17125), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n9602), .ZN(n16908) );
  AOI22_X1 U20081 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12941), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16907) );
  NAND4_X1 U20082 ( .A1(n16910), .A2(n16909), .A3(n16908), .A4(n16907), .ZN(
        n16911) );
  AOI211_X1 U20083 ( .C1(n11462), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n16912), .B(n16911), .ZN(n16913) );
  NAND3_X1 U20084 ( .A1(n16915), .A2(n16914), .A3(n16913), .ZN(n16928) );
  BUF_X2 U20085 ( .A(n16916), .Z(n17143) );
  AOI22_X1 U20086 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16920) );
  INV_X2 U20087 ( .A(n16985), .ZN(n17124) );
  AOI22_X1 U20088 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16919) );
  AOI22_X1 U20089 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(n9600), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16918) );
  AOI22_X1 U20090 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12941), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16917) );
  NAND4_X1 U20091 ( .A1(n16920), .A2(n16919), .A3(n16918), .A4(n16917), .ZN(
        n16926) );
  AOI22_X1 U20092 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9623), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16924) );
  AOI22_X1 U20093 ( .A1(n9603), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9602), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16923) );
  AOI22_X1 U20094 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16922) );
  AOI22_X1 U20095 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16921) );
  NAND4_X1 U20096 ( .A1(n16924), .A2(n16923), .A3(n16922), .A4(n16921), .ZN(
        n16925) );
  NOR2_X1 U20097 ( .A1(n16926), .A2(n16925), .ZN(n16933) );
  NOR3_X1 U20098 ( .A1(n16933), .A2(n16931), .A3(n16938), .ZN(n16927) );
  XNOR2_X1 U20099 ( .A(n16928), .B(n16927), .ZN(n17217) );
  OAI22_X1 U20100 ( .A1(n16930), .A2(n16929), .B1(n17217), .B2(n17197), .ZN(
        P3_U2673) );
  NOR2_X1 U20101 ( .A1(n16931), .A2(n16938), .ZN(n16932) );
  XOR2_X1 U20102 ( .A(n16933), .B(n16932), .Z(n17221) );
  AOI22_X1 U20103 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16936), .B1(n16935), 
        .B2(n16934), .ZN(n16937) );
  OAI21_X1 U20104 ( .B1(n17197), .B2(n17221), .A(n16937), .ZN(P3_U2674) );
  OAI21_X1 U20105 ( .B1(n16940), .B2(n16939), .A(n16938), .ZN(n17230) );
  NAND3_X1 U20106 ( .A1(n16942), .A2(P3_EBX_REG_27__SCAN_IN), .A3(n17197), 
        .ZN(n16941) );
  OAI221_X1 U20107 ( .B1(n16942), .B2(P3_EBX_REG_27__SCAN_IN), .C1(n17197), 
        .C2(n17230), .A(n16941), .ZN(P3_U2676) );
  AOI21_X1 U20108 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17197), .A(n9673), .ZN(
        n16946) );
  OAI21_X1 U20109 ( .B1(n16945), .B2(n16944), .A(n16943), .ZN(n17235) );
  OAI22_X1 U20110 ( .A1(n16947), .A2(n16946), .B1(n17197), .B2(n17235), .ZN(
        P3_U2677) );
  AOI21_X1 U20111 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17197), .A(n9674), .ZN(
        n16949) );
  XNOR2_X1 U20112 ( .A(n16948), .B(n16950), .ZN(n17239) );
  OAI22_X1 U20113 ( .A1(n9673), .A2(n16949), .B1(n17197), .B2(n17239), .ZN(
        P3_U2678) );
  AOI21_X1 U20114 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17197), .A(n9675), .ZN(
        n16953) );
  OAI21_X1 U20115 ( .B1(n16952), .B2(n16951), .A(n16950), .ZN(n17244) );
  OAI22_X1 U20116 ( .A1(n9674), .A2(n16953), .B1(n17197), .B2(n17244), .ZN(
        P3_U2679) );
  AOI21_X1 U20117 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17197), .A(n16954), .ZN(
        n16957) );
  XNOR2_X1 U20118 ( .A(n16956), .B(n16955), .ZN(n17249) );
  OAI22_X1 U20119 ( .A1(n9675), .A2(n16957), .B1(n17197), .B2(n17249), .ZN(
        P3_U2680) );
  AOI22_X1 U20120 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9623), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16962) );
  AOI22_X1 U20121 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16961) );
  AOI22_X1 U20122 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16960) );
  AOI22_X1 U20123 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12941), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16959) );
  NAND4_X1 U20124 ( .A1(n16962), .A2(n16961), .A3(n16960), .A4(n16959), .ZN(
        n16968) );
  AOI22_X1 U20125 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17137), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16966) );
  AOI22_X1 U20126 ( .A1(n9603), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16965) );
  AOI22_X1 U20127 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16964) );
  AOI22_X1 U20128 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16963) );
  NAND4_X1 U20129 ( .A1(n16966), .A2(n16965), .A3(n16964), .A4(n16963), .ZN(
        n16967) );
  NOR2_X1 U20130 ( .A1(n16968), .A2(n16967), .ZN(n17251) );
  NAND3_X1 U20131 ( .A1(n16970), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17197), 
        .ZN(n16969) );
  OAI221_X1 U20132 ( .B1(n16970), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17197), 
        .C2(n17251), .A(n16969), .ZN(P3_U2681) );
  AOI22_X1 U20133 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9623), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16974) );
  AOI22_X1 U20134 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16973) );
  AOI22_X1 U20135 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16972) );
  AOI22_X1 U20136 ( .A1(n12941), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n16971) );
  NAND4_X1 U20137 ( .A1(n16974), .A2(n16973), .A3(n16972), .A4(n16971), .ZN(
        n16980) );
  AOI22_X1 U20138 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(n9602), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16978) );
  AOI22_X1 U20139 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n16977) );
  AOI22_X1 U20140 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n16976) );
  AOI22_X1 U20141 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9603), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n16975) );
  NAND4_X1 U20142 ( .A1(n16978), .A2(n16977), .A3(n16976), .A4(n16975), .ZN(
        n16979) );
  NOR2_X1 U20143 ( .A1(n16980), .A2(n16979), .ZN(n17257) );
  AND2_X1 U20144 ( .A1(n17197), .A2(n16981), .ZN(n16995) );
  AOI22_X1 U20145 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16995), .B1(n16982), 
        .B2(n20795), .ZN(n16983) );
  OAI21_X1 U20146 ( .B1(n17257), .B2(n17197), .A(n16983), .ZN(P3_U2682) );
  AOI22_X1 U20147 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16994) );
  AOI22_X1 U20148 ( .A1(n9603), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(n9623), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n16993) );
  AOI22_X1 U20149 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16984) );
  OAI21_X1 U20150 ( .B1(n16985), .B2(n20794), .A(n16984), .ZN(n16991) );
  AOI22_X1 U20151 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n16989) );
  AOI22_X1 U20152 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17137), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16988) );
  AOI22_X1 U20153 ( .A1(n12941), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n16987) );
  AOI22_X1 U20154 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16986) );
  NAND4_X1 U20155 ( .A1(n16989), .A2(n16988), .A3(n16987), .A4(n16986), .ZN(
        n16990) );
  AOI211_X1 U20156 ( .C1(n17020), .C2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A(
        n16991), .B(n16990), .ZN(n16992) );
  NAND3_X1 U20157 ( .A1(n16994), .A2(n16993), .A3(n16992), .ZN(n17261) );
  INV_X1 U20158 ( .A(n17261), .ZN(n16998) );
  OAI21_X1 U20159 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16996), .A(n16995), .ZN(
        n16997) );
  OAI21_X1 U20160 ( .B1(n16998), .B2(n17197), .A(n16997), .ZN(P3_U2683) );
  AOI22_X1 U20161 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17002) );
  AOI22_X1 U20162 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9603), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17001) );
  AOI22_X1 U20163 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17000) );
  AOI22_X1 U20164 ( .A1(n12941), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16999) );
  NAND4_X1 U20165 ( .A1(n17002), .A2(n17001), .A3(n17000), .A4(n16999), .ZN(
        n17008) );
  AOI22_X1 U20166 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n9623), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17006) );
  AOI22_X1 U20167 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17005) );
  AOI22_X1 U20168 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17004) );
  AOI22_X1 U20169 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17003) );
  NAND4_X1 U20170 ( .A1(n17006), .A2(n17005), .A3(n17004), .A4(n17003), .ZN(
        n17007) );
  NOR2_X1 U20171 ( .A1(n17008), .A2(n17007), .ZN(n17269) );
  AND2_X1 U20172 ( .A1(n17197), .A2(n17009), .ZN(n17024) );
  OAI21_X1 U20173 ( .B1(n17292), .B2(n17009), .A(n17011), .ZN(n17010) );
  OAI21_X1 U20174 ( .B1(n17024), .B2(n17011), .A(n17010), .ZN(n17012) );
  OAI21_X1 U20175 ( .B1(n17269), .B2(n17197), .A(n17012), .ZN(P3_U2684) );
  NAND4_X1 U20176 ( .A1(n18193), .A2(P3_EBX_REG_17__SCAN_IN), .A3(
        P3_EBX_REG_16__SCAN_IN), .A4(n17039), .ZN(n17026) );
  AOI22_X1 U20177 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17023) );
  AOI22_X1 U20178 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17022) );
  AOI22_X1 U20179 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(n9606), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17013) );
  OAI21_X1 U20180 ( .B1(n9591), .B2(n17196), .A(n17013), .ZN(n17019) );
  AOI22_X1 U20181 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17017) );
  AOI22_X1 U20182 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9623), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17016) );
  AOI22_X1 U20183 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17015) );
  AOI22_X1 U20184 ( .A1(n9603), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12941), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17014) );
  NAND4_X1 U20185 ( .A1(n17017), .A2(n17016), .A3(n17015), .A4(n17014), .ZN(
        n17018) );
  AOI211_X1 U20186 ( .C1(n17020), .C2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A(
        n17019), .B(n17018), .ZN(n17021) );
  NAND3_X1 U20187 ( .A1(n17023), .A2(n17022), .A3(n17021), .ZN(n17270) );
  AOI22_X1 U20188 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n17024), .B1(n17203), 
        .B2(n17270), .ZN(n17025) );
  OAI21_X1 U20189 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17026), .A(n17025), .ZN(
        P3_U2685) );
  NAND3_X1 U20190 ( .A1(n18193), .A2(P3_EBX_REG_16__SCAN_IN), .A3(n17039), 
        .ZN(n17038) );
  AOI22_X1 U20191 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17030) );
  AOI22_X1 U20192 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n17029) );
  AOI22_X1 U20193 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(n9602), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17028) );
  AOI22_X1 U20194 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12941), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17027) );
  NAND4_X1 U20195 ( .A1(n17030), .A2(n17029), .A3(n17028), .A4(n17027), .ZN(
        n17036) );
  AOI22_X1 U20196 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17034) );
  AOI22_X1 U20197 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9603), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n17033) );
  AOI22_X1 U20198 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17032) );
  AOI22_X1 U20199 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17031) );
  NAND4_X1 U20200 ( .A1(n17034), .A2(n17033), .A3(n17032), .A4(n17031), .ZN(
        n17035) );
  NOR2_X1 U20201 ( .A1(n17036), .A2(n17035), .ZN(n17281) );
  NAND3_X1 U20202 ( .A1(n17038), .A2(P3_EBX_REG_17__SCAN_IN), .A3(n17197), 
        .ZN(n17037) );
  OAI221_X1 U20203 ( .B1(n17038), .B2(P3_EBX_REG_17__SCAN_IN), .C1(n17197), 
        .C2(n17281), .A(n17037), .ZN(P3_U2686) );
  NAND2_X1 U20204 ( .A1(n18193), .A2(n17039), .ZN(n17051) );
  NOR2_X1 U20205 ( .A1(n17203), .A2(n17039), .ZN(n17064) );
  AOI22_X1 U20206 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17049) );
  AOI22_X1 U20207 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17048) );
  AOI22_X1 U20208 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17040) );
  OAI21_X1 U20209 ( .B1(n9591), .B2(n17158), .A(n17040), .ZN(n17046) );
  AOI22_X1 U20210 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9622), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17044) );
  AOI22_X1 U20211 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17137), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17043) );
  AOI22_X1 U20212 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9623), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n17042) );
  AOI22_X1 U20213 ( .A1(n9603), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12941), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17041) );
  NAND4_X1 U20214 ( .A1(n17044), .A2(n17043), .A3(n17042), .A4(n17041), .ZN(
        n17045) );
  AOI211_X1 U20215 ( .C1(n11462), .C2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A(
        n17046), .B(n17045), .ZN(n17047) );
  NAND3_X1 U20216 ( .A1(n17049), .A2(n17048), .A3(n17047), .ZN(n17282) );
  AOI22_X1 U20217 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17064), .B1(n17203), 
        .B2(n17282), .ZN(n17050) );
  OAI21_X1 U20218 ( .B1(P3_EBX_REG_16__SCAN_IN), .B2(n17051), .A(n17050), .ZN(
        P3_U2687) );
  AOI22_X1 U20219 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n17156), .B1(
        n17052), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n17056) );
  AOI22_X1 U20220 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n9603), .B1(n9606), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n17055) );
  AOI22_X1 U20221 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__7__SCAN_IN), .B2(n9602), .ZN(n17054) );
  AOI22_X1 U20222 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n9607), .B1(
        n12941), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17053) );
  NAND4_X1 U20223 ( .A1(n17056), .A2(n17055), .A3(n17054), .A4(n17053), .ZN(
        n17062) );
  AOI22_X1 U20224 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n17125), .ZN(n17060) );
  AOI22_X1 U20225 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n17155), .B1(
        P3_INSTQUEUE_REG_11__7__SCAN_IN), .B2(n17160), .ZN(n17059) );
  AOI22_X1 U20226 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__7__SCAN_IN), .B2(n9605), .ZN(n17058) );
  AOI22_X1 U20227 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n17143), .B1(
        n9623), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n17057) );
  NAND4_X1 U20228 ( .A1(n17060), .A2(n17059), .A3(n17058), .A4(n17057), .ZN(
        n17061) );
  NOR2_X1 U20229 ( .A1(n17062), .A2(n17061), .ZN(n17291) );
  INV_X1 U20230 ( .A(n17063), .ZN(n17065) );
  OAI21_X1 U20231 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17065), .A(n17064), .ZN(
        n17066) );
  OAI21_X1 U20232 ( .B1(n17291), .B2(n17197), .A(n17066), .ZN(P3_U2688) );
  NAND2_X1 U20233 ( .A1(n18193), .A2(n17067), .ZN(n17080) );
  NOR2_X1 U20234 ( .A1(n17203), .A2(n17067), .ZN(n17091) );
  AOI22_X1 U20235 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n17078) );
  AOI22_X1 U20236 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(n9607), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n17077) );
  INV_X1 U20237 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n17069) );
  AOI22_X1 U20238 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17137), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n17068) );
  OAI21_X1 U20239 ( .B1(n11441), .B2(n17069), .A(n17068), .ZN(n17075) );
  AOI22_X1 U20240 ( .A1(n9603), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n9600), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n17073) );
  AOI22_X1 U20241 ( .A1(n17143), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17072) );
  AOI22_X1 U20242 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12941), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17071) );
  AOI22_X1 U20243 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17070) );
  NAND4_X1 U20244 ( .A1(n17073), .A2(n17072), .A3(n17071), .A4(n17070), .ZN(
        n17074) );
  AOI211_X1 U20245 ( .C1(n9596), .C2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n17075), .B(n17074), .ZN(n17076) );
  NAND3_X1 U20246 ( .A1(n17078), .A2(n17077), .A3(n17076), .ZN(n17293) );
  AOI22_X1 U20247 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17091), .B1(n17203), 
        .B2(n17293), .ZN(n17079) );
  OAI21_X1 U20248 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17080), .A(n17079), .ZN(
        P3_U2689) );
  AOI22_X1 U20249 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17084) );
  AOI22_X1 U20250 ( .A1(n9603), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n17083) );
  AOI22_X1 U20251 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9606), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n17082) );
  AOI22_X1 U20252 ( .A1(n12941), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n17081) );
  NAND4_X1 U20253 ( .A1(n17084), .A2(n17083), .A3(n17082), .A4(n17081), .ZN(
        n17090) );
  AOI22_X1 U20254 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17088) );
  AOI22_X1 U20255 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17137), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17087) );
  AOI22_X1 U20256 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n17086) );
  AOI22_X1 U20257 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(n9607), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17085) );
  NAND4_X1 U20258 ( .A1(n17088), .A2(n17087), .A3(n17086), .A4(n17085), .ZN(
        n17089) );
  NOR2_X1 U20259 ( .A1(n17090), .A2(n17089), .ZN(n17298) );
  INV_X1 U20260 ( .A(n17104), .ZN(n17092) );
  OAI21_X1 U20261 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(n17092), .A(n17091), .ZN(
        n17093) );
  OAI21_X1 U20262 ( .B1(n17298), .B2(n17197), .A(n17093), .ZN(P3_U2690) );
  AOI22_X1 U20263 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n17161), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17097) );
  AOI22_X1 U20264 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17096) );
  AOI22_X1 U20265 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17155), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17095) );
  AOI22_X1 U20266 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12941), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17094) );
  NAND4_X1 U20267 ( .A1(n17097), .A2(n17096), .A3(n17095), .A4(n17094), .ZN(
        n17103) );
  AOI22_X1 U20268 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n9602), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17101) );
  AOI22_X1 U20269 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17100) );
  AOI22_X1 U20270 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9603), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n17099) );
  AOI22_X1 U20271 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17098) );
  NAND4_X1 U20272 ( .A1(n17101), .A2(n17100), .A3(n17099), .A4(n17098), .ZN(
        n17102) );
  NOR2_X1 U20273 ( .A1(n17103), .A2(n17102), .ZN(n17302) );
  OAI21_X1 U20274 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n17117), .A(n17104), .ZN(
        n17105) );
  AOI22_X1 U20275 ( .A1(n17203), .A2(n17302), .B1(n17105), .B2(n17197), .ZN(
        P3_U2691) );
  AOI22_X1 U20276 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17116) );
  AOI22_X1 U20277 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17115) );
  AOI22_X1 U20278 ( .A1(n9596), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17106) );
  OAI21_X1 U20279 ( .B1(n17159), .B2(n17190), .A(n17106), .ZN(n17113) );
  AOI22_X1 U20280 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17111) );
  AOI22_X1 U20281 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17161), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17110) );
  AOI22_X1 U20282 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9603), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17109) );
  AOI22_X1 U20283 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17108) );
  NAND4_X1 U20284 ( .A1(n17111), .A2(n17110), .A3(n17109), .A4(n17108), .ZN(
        n17112) );
  AOI211_X1 U20285 ( .C1(n17020), .C2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A(
        n17113), .B(n17112), .ZN(n17114) );
  NAND3_X1 U20286 ( .A1(n17116), .A2(n17115), .A3(n17114), .ZN(n17305) );
  AOI21_X1 U20287 ( .B1(n17119), .B2(n17118), .A(n17117), .ZN(n17120) );
  MUX2_X1 U20288 ( .A(n17305), .B(n17120), .S(n17197), .Z(P3_U2692) );
  NAND2_X1 U20289 ( .A1(n18193), .A2(n17206), .ZN(n17201) );
  INV_X1 U20290 ( .A(n17201), .ZN(n17202) );
  NAND4_X1 U20291 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(P3_EBX_REG_4__SCAN_IN), 
        .A3(n17188), .A4(n17202), .ZN(n17175) );
  NOR3_X1 U20292 ( .A1(n17121), .A2(n20839), .A3(n17175), .ZN(n17172) );
  NAND3_X1 U20293 ( .A1(P3_EBX_REG_9__SCAN_IN), .A2(P3_EBX_REG_8__SCAN_IN), 
        .A3(n17172), .ZN(n17136) );
  NOR2_X1 U20294 ( .A1(n17203), .A2(n17122), .ZN(n17151) );
  AOI22_X1 U20295 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(n9602), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17134) );
  AOI22_X1 U20296 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(n9623), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17133) );
  AOI22_X1 U20297 ( .A1(n9607), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9600), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17123) );
  OAI21_X1 U20298 ( .B1(n17159), .B2(n17196), .A(n17123), .ZN(n17131) );
  AOI22_X1 U20299 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17137), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17129) );
  AOI22_X1 U20300 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9603), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17128) );
  AOI22_X1 U20301 ( .A1(n17160), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17127) );
  AOI22_X1 U20302 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17126) );
  NAND4_X1 U20303 ( .A1(n17129), .A2(n17128), .A3(n17127), .A4(n17126), .ZN(
        n17130) );
  AOI211_X1 U20304 ( .C1(n9596), .C2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A(
        n17131), .B(n17130), .ZN(n17132) );
  NAND3_X1 U20305 ( .A1(n17134), .A2(n17133), .A3(n17132), .ZN(n17308) );
  AOI22_X1 U20306 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17151), .B1(n17203), 
        .B2(n17308), .ZN(n17135) );
  OAI21_X1 U20307 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17136), .A(n17135), .ZN(
        P3_U2693) );
  AOI22_X1 U20308 ( .A1(n17137), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n17142) );
  AOI22_X1 U20309 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n17141) );
  AOI22_X1 U20310 ( .A1(n9606), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(n9607), .B2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n17140) );
  AOI22_X1 U20311 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12941), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17139) );
  NAND4_X1 U20312 ( .A1(n17142), .A2(n17141), .A3(n17140), .A4(n17139), .ZN(
        n17150) );
  AOI22_X1 U20313 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17143), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17148) );
  AOI22_X1 U20314 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9603), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17147) );
  AOI22_X1 U20315 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n17146) );
  AOI22_X1 U20316 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(n9622), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n17145) );
  NAND4_X1 U20317 ( .A1(n17148), .A2(n17147), .A3(n17146), .A4(n17145), .ZN(
        n17149) );
  NOR2_X1 U20318 ( .A1(n17150), .A2(n17149), .ZN(n17313) );
  INV_X1 U20319 ( .A(n17171), .ZN(n17152) );
  OAI21_X1 U20320 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17152), .A(n17151), .ZN(
        n17153) );
  OAI21_X1 U20321 ( .B1(n17313), .B2(n17197), .A(n17153), .ZN(P3_U2694) );
  AOI22_X1 U20322 ( .A1(n17155), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n17154), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17170) );
  AOI22_X1 U20323 ( .A1(n17020), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9603), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17169) );
  AOI22_X1 U20324 ( .A1(n17156), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n9602), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17157) );
  OAI21_X1 U20325 ( .B1(n17159), .B2(n17158), .A(n17157), .ZN(n17167) );
  AOI22_X1 U20326 ( .A1(n9605), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17160), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17165) );
  AOI22_X1 U20327 ( .A1(n17124), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9607), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17164) );
  AOI22_X1 U20328 ( .A1(n17161), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17125), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17163) );
  AOI22_X1 U20329 ( .A1(n9597), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(n9606), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n17162) );
  NAND4_X1 U20330 ( .A1(n17165), .A2(n17164), .A3(n17163), .A4(n17162), .ZN(
        n17166) );
  AOI211_X1 U20331 ( .C1(n11462), .C2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A(
        n17167), .B(n17166), .ZN(n17168) );
  NAND3_X1 U20332 ( .A1(n17170), .A2(n17169), .A3(n17168), .ZN(n17319) );
  INV_X1 U20333 ( .A(n17319), .ZN(n17174) );
  OAI21_X1 U20334 ( .B1(P3_EBX_REG_8__SCAN_IN), .B2(n17172), .A(n17171), .ZN(
        n17173) );
  AOI22_X1 U20335 ( .A1(n17203), .A2(n17174), .B1(n17173), .B2(n17197), .ZN(
        P3_U2695) );
  INV_X1 U20336 ( .A(n17175), .ZN(n17179) );
  AOI22_X1 U20337 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17197), .B1(
        P3_EBX_REG_6__SCAN_IN), .B2(n17179), .ZN(n17177) );
  OAI22_X1 U20338 ( .A1(n9712), .A2(n17177), .B1(n17176), .B2(n17197), .ZN(
        P3_U2696) );
  NAND2_X1 U20339 ( .A1(n17197), .A2(n17178), .ZN(n17182) );
  AOI22_X1 U20340 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n17203), .B1(
        n17179), .B2(n20839), .ZN(n17180) );
  OAI21_X1 U20341 ( .B1(n20839), .B2(n17182), .A(n17180), .ZN(P3_U2697) );
  NOR2_X1 U20342 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17187), .ZN(n17183) );
  OAI22_X1 U20343 ( .A1(n17183), .A2(n17182), .B1(n17181), .B2(n17197), .ZN(
        P3_U2698) );
  OAI21_X1 U20344 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17184), .A(n17197), .ZN(
        n17186) );
  INV_X1 U20345 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17185) );
  OAI22_X1 U20346 ( .A1(n17187), .A2(n17186), .B1(n17185), .B2(n17197), .ZN(
        P3_U2699) );
  AND2_X1 U20347 ( .A1(n17188), .A2(n17202), .ZN(n17192) );
  NOR2_X1 U20348 ( .A1(n17189), .A2(n17201), .ZN(n17194) );
  AOI21_X1 U20349 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17197), .A(n17194), .ZN(
        n17191) );
  OAI22_X1 U20350 ( .A1(n17192), .A2(n17191), .B1(n17190), .B2(n17197), .ZN(
        P3_U2700) );
  AOI221_X1 U20351 ( .B1(n17193), .B2(n17206), .C1(n17292), .C2(n17206), .A(
        P3_EBX_REG_2__SCAN_IN), .ZN(n17195) );
  AOI211_X1 U20352 ( .C1(n17203), .C2(n17196), .A(n17195), .B(n17194), .ZN(
        P3_U2701) );
  OAI222_X1 U20353 ( .A1(n17201), .A2(n17200), .B1(n17199), .B2(n17206), .C1(
        n17198), .C2(n17197), .ZN(P3_U2702) );
  AOI22_X1 U20354 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17203), .B1(
        n17202), .B2(n17205), .ZN(n17204) );
  OAI21_X1 U20355 ( .B1(n17206), .B2(n17205), .A(n17204), .ZN(P3_U2703) );
  INV_X1 U20356 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17362) );
  INV_X1 U20357 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n20862) );
  INV_X1 U20358 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17463) );
  INV_X1 U20359 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17396) );
  NAND4_X1 U20360 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(P3_EAX_REG_5__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17208) );
  INV_X1 U20361 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17389) );
  INV_X1 U20362 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17450) );
  INV_X1 U20363 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17392) );
  INV_X1 U20364 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17394) );
  NOR4_X1 U20365 ( .A1(n17389), .A2(n17450), .A3(n17392), .A4(n17394), .ZN(
        n17209) );
  NOR2_X2 U20366 ( .A1(n17463), .A2(n17294), .ZN(n17288) );
  NAND2_X1 U20367 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .ZN(n17250) );
  NAND4_X1 U20368 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(P3_EAX_REG_19__SCAN_IN), 
        .A3(P3_EAX_REG_18__SCAN_IN), .A4(P3_EAX_REG_17__SCAN_IN), .ZN(n17210)
         );
  NAND2_X1 U20369 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17246), .ZN(n17245) );
  NOR2_X2 U20370 ( .A1(n20862), .A2(n9654), .ZN(n17231) );
  NAND2_X1 U20371 ( .A1(n17214), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17213) );
  NAND2_X1 U20372 ( .A1(n17211), .A2(n17317), .ZN(n17256) );
  OAI21_X1 U20373 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17213), .A(n17212), .ZN(
        P3_U2704) );
  NAND2_X1 U20374 ( .A1(n18182), .A2(n17317), .ZN(n17287) );
  AOI22_X1 U20375 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17276), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17283), .ZN(n17216) );
  OAI211_X1 U20376 ( .C1(n17214), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17340), .B(
        n17213), .ZN(n17215) );
  OAI211_X1 U20377 ( .C1(n17217), .C2(n17342), .A(n17216), .B(n17215), .ZN(
        P3_U2705) );
  AOI22_X1 U20378 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17276), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n17283), .ZN(n17220) );
  OAI211_X1 U20379 ( .C1(n17223), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17340), .B(
        n17218), .ZN(n17219) );
  OAI211_X1 U20380 ( .C1(n17342), .C2(n17221), .A(n17220), .B(n17219), .ZN(
        P3_U2706) );
  AOI22_X1 U20381 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17276), .B1(n17222), .B2(
        n17347), .ZN(n17226) );
  AOI211_X1 U20382 ( .C1(n17362), .C2(n17227), .A(n17223), .B(n17317), .ZN(
        n17224) );
  INV_X1 U20383 ( .A(n17224), .ZN(n17225) );
  OAI211_X1 U20384 ( .C1(n17256), .C2(n18176), .A(n17226), .B(n17225), .ZN(
        P3_U2707) );
  AOI22_X1 U20385 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17276), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n17283), .ZN(n17229) );
  OAI211_X1 U20386 ( .C1(n17231), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17340), .B(
        n17227), .ZN(n17228) );
  OAI211_X1 U20387 ( .C1(n17342), .C2(n17230), .A(n17229), .B(n17228), .ZN(
        P3_U2708) );
  AOI22_X1 U20388 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17276), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17283), .ZN(n17234) );
  AOI211_X1 U20389 ( .C1(n20862), .C2(n9654), .A(n17231), .B(n17317), .ZN(
        n17232) );
  INV_X1 U20390 ( .A(n17232), .ZN(n17233) );
  OAI211_X1 U20391 ( .C1(n17342), .C2(n17235), .A(n17234), .B(n17233), .ZN(
        P3_U2709) );
  AOI22_X1 U20392 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17276), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17283), .ZN(n17238) );
  OAI211_X1 U20393 ( .C1(n17236), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17340), .B(
        n9654), .ZN(n17237) );
  OAI211_X1 U20394 ( .C1(n17239), .C2(n17342), .A(n17238), .B(n17237), .ZN(
        P3_U2710) );
  AOI22_X1 U20395 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17276), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17283), .ZN(n17243) );
  OAI211_X1 U20396 ( .C1(n17241), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17340), .B(
        n17240), .ZN(n17242) );
  OAI211_X1 U20397 ( .C1(n17244), .C2(n17342), .A(n17243), .B(n17242), .ZN(
        P3_U2711) );
  AOI22_X1 U20398 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17276), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17283), .ZN(n17248) );
  OAI211_X1 U20399 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17246), .A(n17340), .B(
        n17245), .ZN(n17247) );
  OAI211_X1 U20400 ( .C1(n17249), .C2(n17342), .A(n17248), .B(n17247), .ZN(
        P3_U2712) );
  INV_X1 U20401 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17379) );
  INV_X1 U20402 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17418) );
  NOR3_X1 U20403 ( .A1(n17292), .A2(n17284), .A3(n17418), .ZN(n17273) );
  INV_X1 U20404 ( .A(n17273), .ZN(n17277) );
  NAND2_X1 U20405 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17271), .ZN(n17266) );
  NAND2_X1 U20406 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17263), .ZN(n17262) );
  NAND2_X1 U20407 ( .A1(n17340), .A2(n17262), .ZN(n17260) );
  OAI21_X1 U20408 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17349), .A(n17260), .ZN(
        n17254) );
  NOR3_X1 U20409 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17250), .A3(n17266), .ZN(
        n17253) );
  INV_X1 U20410 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n18185) );
  OAI22_X1 U20411 ( .A1(n17251), .A2(n17342), .B1(n18185), .B2(n17256), .ZN(
        n17252) );
  AOI211_X1 U20412 ( .C1(P3_EAX_REG_22__SCAN_IN), .C2(n17254), .A(n17253), .B(
        n17252), .ZN(n17255) );
  OAI21_X1 U20413 ( .B1(n18186), .B2(n17287), .A(n17255), .ZN(P3_U2713) );
  INV_X1 U20414 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17373) );
  OAI22_X1 U20415 ( .A1(n17257), .A2(n17342), .B1(n14259), .B2(n17256), .ZN(
        n17258) );
  AOI21_X1 U20416 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17276), .A(n17258), .ZN(
        n17259) );
  OAI221_X1 U20417 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17262), .C1(n17373), 
        .C2(n17260), .A(n17259), .ZN(P3_U2714) );
  INV_X1 U20418 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18177) );
  AOI22_X1 U20419 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17283), .B1(n17347), .B2(
        n17261), .ZN(n17265) );
  OAI211_X1 U20420 ( .C1(n17263), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17340), .B(
        n17262), .ZN(n17264) );
  OAI211_X1 U20421 ( .C1(n17287), .C2(n18177), .A(n17265), .B(n17264), .ZN(
        P3_U2715) );
  AOI22_X1 U20422 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17276), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17283), .ZN(n17268) );
  OAI211_X1 U20423 ( .C1(n17271), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17340), .B(
        n17266), .ZN(n17267) );
  OAI211_X1 U20424 ( .C1(n17269), .C2(n17342), .A(n17268), .B(n17267), .ZN(
        P3_U2716) );
  INV_X1 U20425 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18168) );
  AOI22_X1 U20426 ( .A1(BUF2_REG_18__SCAN_IN), .A2(n17283), .B1(n17347), .B2(
        n17270), .ZN(n17275) );
  INV_X1 U20427 ( .A(n17271), .ZN(n17272) );
  OAI211_X1 U20428 ( .C1(n17273), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17340), .B(
        n17272), .ZN(n17274) );
  OAI211_X1 U20429 ( .C1(n17287), .C2(n18168), .A(n17275), .B(n17274), .ZN(
        P3_U2717) );
  AOI22_X1 U20430 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17276), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17283), .ZN(n17280) );
  INV_X1 U20431 ( .A(n17284), .ZN(n17278) );
  OAI211_X1 U20432 ( .C1(n17278), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17340), .B(
        n17277), .ZN(n17279) );
  OAI211_X1 U20433 ( .C1(n17281), .C2(n17342), .A(n17280), .B(n17279), .ZN(
        P3_U2718) );
  INV_X1 U20434 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18155) );
  AOI22_X1 U20435 ( .A1(BUF2_REG_16__SCAN_IN), .A2(n17283), .B1(n17347), .B2(
        n17282), .ZN(n17286) );
  OAI211_X1 U20436 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17288), .A(n17340), .B(
        n17284), .ZN(n17285) );
  OAI211_X1 U20437 ( .C1(n17287), .C2(n18155), .A(n17286), .B(n17285), .ZN(
        P3_U2719) );
  AOI211_X1 U20438 ( .C1(n17463), .C2(n17294), .A(n17317), .B(n17288), .ZN(
        n17289) );
  AOI21_X1 U20439 ( .B1(n17348), .B2(BUF2_REG_15__SCAN_IN), .A(n17289), .ZN(
        n17290) );
  OAI21_X1 U20440 ( .B1(n17291), .B2(n17342), .A(n17290), .ZN(P3_U2720) );
  NOR3_X1 U20441 ( .A1(n17292), .A2(n17396), .A3(n17321), .ZN(n17312) );
  NAND2_X1 U20442 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17312), .ZN(n17310) );
  INV_X1 U20443 ( .A(n17310), .ZN(n17315) );
  NAND2_X1 U20444 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17315), .ZN(n17307) );
  NOR2_X1 U20445 ( .A1(n17450), .A2(n17307), .ZN(n17301) );
  NAND2_X1 U20446 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17304), .ZN(n17297) );
  AOI22_X1 U20447 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17348), .B1(n17347), .B2(
        n17293), .ZN(n17296) );
  NAND3_X1 U20448 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17340), .A3(n17294), 
        .ZN(n17295) );
  OAI211_X1 U20449 ( .C1(P3_EAX_REG_14__SCAN_IN), .C2(n17297), .A(n17296), .B(
        n17295), .ZN(P3_U2721) );
  INV_X1 U20450 ( .A(n17297), .ZN(n17300) );
  AOI21_X1 U20451 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17340), .A(n17304), .ZN(
        n17299) );
  OAI222_X1 U20452 ( .A1(n17345), .A2(n20825), .B1(n17300), .B2(n17299), .C1(
        n17342), .C2(n17298), .ZN(P3_U2722) );
  INV_X1 U20453 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17452) );
  AOI21_X1 U20454 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17340), .A(n17301), .ZN(
        n17303) );
  OAI222_X1 U20455 ( .A1(n17345), .A2(n17452), .B1(n17304), .B2(n17303), .C1(
        n17342), .C2(n17302), .ZN(P3_U2723) );
  NAND2_X1 U20456 ( .A1(n17340), .A2(n17307), .ZN(n17311) );
  AOI22_X1 U20457 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17348), .B1(n17347), .B2(
        n17305), .ZN(n17306) );
  OAI221_X1 U20458 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17307), .C1(n17450), 
        .C2(n17311), .A(n17306), .ZN(P3_U2724) );
  AOI22_X1 U20459 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17348), .B1(n17347), .B2(
        n17308), .ZN(n17309) );
  OAI221_X1 U20460 ( .B1(n17311), .B2(n17392), .C1(n17311), .C2(n17310), .A(
        n17309), .ZN(P3_U2725) );
  AOI21_X1 U20461 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17340), .A(n17312), .ZN(
        n17314) );
  OAI222_X1 U20462 ( .A1(n17345), .A2(n17446), .B1(n17315), .B2(n17314), .C1(
        n17342), .C2(n17313), .ZN(P3_U2726) );
  AOI211_X1 U20463 ( .C1(n17396), .C2(n17321), .A(n17317), .B(n17316), .ZN(
        n17318) );
  AOI21_X1 U20464 ( .B1(n17347), .B2(n17319), .A(n17318), .ZN(n17320) );
  OAI21_X1 U20465 ( .B1(n17444), .B2(n17345), .A(n17320), .ZN(P3_U2727) );
  INV_X1 U20466 ( .A(n17321), .ZN(n17324) );
  INV_X1 U20467 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17401) );
  INV_X1 U20468 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n20908) );
  INV_X1 U20469 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17436) );
  NOR3_X1 U20470 ( .A1(n17436), .A2(n17413), .A3(n17349), .ZN(n17339) );
  AND2_X1 U20471 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17339), .ZN(n17344) );
  NAND2_X1 U20472 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17344), .ZN(n17332) );
  NOR2_X1 U20473 ( .A1(n20908), .A2(n17332), .ZN(n17335) );
  NAND2_X1 U20474 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17335), .ZN(n17325) );
  NOR2_X1 U20475 ( .A1(n17401), .A2(n17325), .ZN(n17328) );
  AOI21_X1 U20476 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17340), .A(n17328), .ZN(
        n17323) );
  OAI222_X1 U20477 ( .A1(n17345), .A2(n18190), .B1(n17324), .B2(n17323), .C1(
        n17342), .C2(n17322), .ZN(P3_U2728) );
  INV_X1 U20478 ( .A(n17325), .ZN(n17331) );
  AOI21_X1 U20479 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17340), .A(n17331), .ZN(
        n17327) );
  OAI222_X1 U20480 ( .A1(n18186), .A2(n17345), .B1(n17328), .B2(n17327), .C1(
        n17342), .C2(n17326), .ZN(P3_U2729) );
  AOI21_X1 U20481 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17340), .A(n17335), .ZN(
        n17330) );
  OAI222_X1 U20482 ( .A1(n18181), .A2(n17345), .B1(n17331), .B2(n17330), .C1(
        n17342), .C2(n17329), .ZN(P3_U2730) );
  INV_X1 U20483 ( .A(n17332), .ZN(n17338) );
  AOI21_X1 U20484 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17340), .A(n17338), .ZN(
        n17334) );
  OAI222_X1 U20485 ( .A1(n18177), .A2(n17345), .B1(n17335), .B2(n17334), .C1(
        n17342), .C2(n17333), .ZN(P3_U2731) );
  AOI21_X1 U20486 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17340), .A(n17344), .ZN(
        n17337) );
  OAI222_X1 U20487 ( .A1(n18172), .A2(n17345), .B1(n17338), .B2(n17337), .C1(
        n17342), .C2(n17336), .ZN(P3_U2732) );
  AOI21_X1 U20488 ( .B1(P3_EAX_REG_2__SCAN_IN), .B2(n17340), .A(n17339), .ZN(
        n17343) );
  OAI222_X1 U20489 ( .A1(n18168), .A2(n17345), .B1(n17344), .B2(n17343), .C1(
        n17342), .C2(n17341), .ZN(P3_U2733) );
  AOI22_X1 U20490 ( .A1(n17348), .A2(BUF2_REG_1__SCAN_IN), .B1(n17347), .B2(
        n17346), .ZN(n17354) );
  NOR2_X1 U20491 ( .A1(n17413), .A2(n17349), .ZN(n17352) );
  NOR2_X1 U20492 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17349), .ZN(n17351) );
  OAI22_X1 U20493 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17352), .B1(n17351), .B2(
        n17350), .ZN(n17353) );
  NAND2_X1 U20494 ( .A1(n17354), .A2(n17353), .ZN(P3_U2734) );
  NOR2_X2 U20495 ( .A1(n18773), .A2(n17823), .ZN(n18807) );
  NOR2_X4 U20496 ( .A1(n18807), .A2(n17357), .ZN(n17399) );
  AND2_X1 U20497 ( .A1(n17399), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20498 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17433) );
  AOI22_X1 U20499 ( .A1(n18807), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17358) );
  OAI21_X1 U20500 ( .B1(n17433), .B2(n17382), .A(n17358), .ZN(P3_U2737) );
  INV_X1 U20501 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17360) );
  AOI22_X1 U20502 ( .A1(n18807), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17359) );
  OAI21_X1 U20503 ( .B1(n17360), .B2(n17382), .A(n17359), .ZN(P3_U2738) );
  AOI22_X1 U20504 ( .A1(n18807), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17361) );
  OAI21_X1 U20505 ( .B1(n17362), .B2(n17382), .A(n17361), .ZN(P3_U2739) );
  INV_X1 U20506 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17429) );
  AOI22_X1 U20507 ( .A1(n18807), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17363) );
  OAI21_X1 U20508 ( .B1(n17429), .B2(n17382), .A(n17363), .ZN(P3_U2740) );
  AOI22_X1 U20509 ( .A1(n18807), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17364) );
  OAI21_X1 U20510 ( .B1(n20862), .B2(n17382), .A(n17364), .ZN(P3_U2741) );
  INV_X1 U20511 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17366) );
  AOI22_X1 U20512 ( .A1(n18807), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17365) );
  OAI21_X1 U20513 ( .B1(n17366), .B2(n17382), .A(n17365), .ZN(P3_U2742) );
  AOI22_X1 U20514 ( .A1(n18807), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17367) );
  OAI21_X1 U20515 ( .B1(n9728), .B2(n17382), .A(n17367), .ZN(P3_U2743) );
  INV_X1 U20516 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17369) );
  AOI22_X1 U20517 ( .A1(n18807), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17368) );
  OAI21_X1 U20518 ( .B1(n17369), .B2(n17382), .A(n17368), .ZN(P3_U2744) );
  INV_X1 U20519 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17371) );
  AOI22_X1 U20520 ( .A1(n17410), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17370) );
  OAI21_X1 U20521 ( .B1(n17371), .B2(n17382), .A(n17370), .ZN(P3_U2745) );
  AOI22_X1 U20522 ( .A1(n17410), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17372) );
  OAI21_X1 U20523 ( .B1(n17373), .B2(n17382), .A(n17372), .ZN(P3_U2746) );
  INV_X1 U20524 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17375) );
  AOI22_X1 U20525 ( .A1(n17410), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17374) );
  OAI21_X1 U20526 ( .B1(n17375), .B2(n17382), .A(n17374), .ZN(P3_U2747) );
  INV_X1 U20527 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17377) );
  AOI22_X1 U20528 ( .A1(n17410), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17376) );
  OAI21_X1 U20529 ( .B1(n17377), .B2(n17382), .A(n17376), .ZN(P3_U2748) );
  AOI22_X1 U20530 ( .A1(n17410), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17378) );
  OAI21_X1 U20531 ( .B1(n17379), .B2(n17382), .A(n17378), .ZN(P3_U2749) );
  AOI22_X1 U20532 ( .A1(n17410), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17380) );
  OAI21_X1 U20533 ( .B1(n17418), .B2(n17382), .A(n17380), .ZN(P3_U2750) );
  INV_X1 U20534 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17383) );
  AOI22_X1 U20535 ( .A1(n17410), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17381) );
  OAI21_X1 U20536 ( .B1(n17383), .B2(n17382), .A(n17381), .ZN(P3_U2751) );
  AOI22_X1 U20537 ( .A1(n17410), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17384) );
  OAI21_X1 U20538 ( .B1(n17463), .B2(n17412), .A(n17384), .ZN(P3_U2752) );
  INV_X1 U20539 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17458) );
  AOI22_X1 U20540 ( .A1(n17410), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17385) );
  OAI21_X1 U20541 ( .B1(n17458), .B2(n17412), .A(n17385), .ZN(P3_U2753) );
  INV_X1 U20542 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17387) );
  AOI22_X1 U20543 ( .A1(n17410), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17386) );
  OAI21_X1 U20544 ( .B1(n17387), .B2(n17412), .A(n17386), .ZN(P3_U2754) );
  AOI22_X1 U20545 ( .A1(n17410), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17388) );
  OAI21_X1 U20546 ( .B1(n17389), .B2(n17412), .A(n17388), .ZN(P3_U2755) );
  AOI22_X1 U20547 ( .A1(n17410), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17390) );
  OAI21_X1 U20548 ( .B1(n17450), .B2(n17412), .A(n17390), .ZN(P3_U2756) );
  AOI22_X1 U20549 ( .A1(n17410), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17391) );
  OAI21_X1 U20550 ( .B1(n17392), .B2(n17412), .A(n17391), .ZN(P3_U2757) );
  AOI22_X1 U20551 ( .A1(n17410), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17393) );
  OAI21_X1 U20552 ( .B1(n17394), .B2(n17412), .A(n17393), .ZN(P3_U2758) );
  AOI22_X1 U20553 ( .A1(n17410), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17395) );
  OAI21_X1 U20554 ( .B1(n17396), .B2(n17412), .A(n17395), .ZN(P3_U2759) );
  INV_X1 U20555 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17398) );
  AOI22_X1 U20556 ( .A1(n17410), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17397) );
  OAI21_X1 U20557 ( .B1(n17398), .B2(n17412), .A(n17397), .ZN(P3_U2760) );
  AOI22_X1 U20558 ( .A1(n17410), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17400) );
  OAI21_X1 U20559 ( .B1(n17401), .B2(n17412), .A(n17400), .ZN(P3_U2761) );
  INV_X1 U20560 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17403) );
  AOI22_X1 U20561 ( .A1(n17410), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17402) );
  OAI21_X1 U20562 ( .B1(n17403), .B2(n17412), .A(n17402), .ZN(P3_U2762) );
  AOI22_X1 U20563 ( .A1(n17410), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17404) );
  OAI21_X1 U20564 ( .B1(n20908), .B2(n17412), .A(n17404), .ZN(P3_U2763) );
  INV_X1 U20565 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17406) );
  AOI22_X1 U20566 ( .A1(n17410), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17405) );
  OAI21_X1 U20567 ( .B1(n17406), .B2(n17412), .A(n17405), .ZN(P3_U2764) );
  INV_X1 U20568 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17408) );
  AOI22_X1 U20569 ( .A1(n17410), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17407) );
  OAI21_X1 U20570 ( .B1(n17408), .B2(n17412), .A(n17407), .ZN(P3_U2765) );
  AOI22_X1 U20571 ( .A1(n17410), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17409) );
  OAI21_X1 U20572 ( .B1(n17436), .B2(n17412), .A(n17409), .ZN(P3_U2766) );
  AOI22_X1 U20573 ( .A1(n17410), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17399), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17411) );
  OAI21_X1 U20574 ( .B1(n17413), .B2(n17412), .A(n17411), .ZN(P3_U2767) );
  NAND3_X1 U20575 ( .A1(n18164), .A2(n17415), .A3(n17414), .ZN(n17462) );
  AOI22_X1 U20576 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17454), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17453), .ZN(n17416) );
  OAI21_X1 U20577 ( .B1(n18155), .B2(n17456), .A(n17416), .ZN(P3_U2768) );
  AOI22_X1 U20578 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17460), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17453), .ZN(n17417) );
  OAI21_X1 U20579 ( .B1(n17418), .B2(n17462), .A(n17417), .ZN(P3_U2769) );
  AOI22_X1 U20580 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17454), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17453), .ZN(n17419) );
  OAI21_X1 U20581 ( .B1(n18168), .B2(n17456), .A(n17419), .ZN(P3_U2770) );
  AOI22_X1 U20582 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17454), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17453), .ZN(n17420) );
  OAI21_X1 U20583 ( .B1(n18172), .B2(n17456), .A(n17420), .ZN(P3_U2771) );
  AOI22_X1 U20584 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17454), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17453), .ZN(n17421) );
  OAI21_X1 U20585 ( .B1(n18177), .B2(n17456), .A(n17421), .ZN(P3_U2772) );
  AOI22_X1 U20586 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17454), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17453), .ZN(n17422) );
  OAI21_X1 U20587 ( .B1(n18181), .B2(n17456), .A(n17422), .ZN(P3_U2773) );
  AOI22_X1 U20588 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17454), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17453), .ZN(n17423) );
  OAI21_X1 U20589 ( .B1(n18186), .B2(n17456), .A(n17423), .ZN(P3_U2774) );
  AOI22_X1 U20590 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17454), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17453), .ZN(n17424) );
  OAI21_X1 U20591 ( .B1(n18190), .B2(n17456), .A(n17424), .ZN(P3_U2775) );
  AOI22_X1 U20592 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17454), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17453), .ZN(n17425) );
  OAI21_X1 U20593 ( .B1(n17444), .B2(n17456), .A(n17425), .ZN(P3_U2776) );
  AOI22_X1 U20594 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17454), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17453), .ZN(n17426) );
  OAI21_X1 U20595 ( .B1(n17446), .B2(n17456), .A(n17426), .ZN(P3_U2777) );
  INV_X1 U20596 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17448) );
  AOI22_X1 U20597 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17454), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17453), .ZN(n17427) );
  OAI21_X1 U20598 ( .B1(n17448), .B2(n17456), .A(n17427), .ZN(P3_U2778) );
  AOI22_X1 U20599 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17460), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17453), .ZN(n17428) );
  OAI21_X1 U20600 ( .B1(n17429), .B2(n17462), .A(n17428), .ZN(P3_U2779) );
  AOI22_X1 U20601 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17454), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17453), .ZN(n17430) );
  OAI21_X1 U20602 ( .B1(n17452), .B2(n17456), .A(n17430), .ZN(P3_U2780) );
  AOI22_X1 U20603 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17454), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17453), .ZN(n17431) );
  OAI21_X1 U20604 ( .B1(n20825), .B2(n17456), .A(n17431), .ZN(P3_U2781) );
  AOI22_X1 U20605 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17460), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17453), .ZN(n17432) );
  OAI21_X1 U20606 ( .B1(n17433), .B2(n17462), .A(n17432), .ZN(P3_U2782) );
  AOI22_X1 U20607 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17454), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17453), .ZN(n17434) );
  OAI21_X1 U20608 ( .B1(n18155), .B2(n17456), .A(n17434), .ZN(P3_U2783) );
  AOI22_X1 U20609 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17460), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17453), .ZN(n17435) );
  OAI21_X1 U20610 ( .B1(n17436), .B2(n17462), .A(n17435), .ZN(P3_U2784) );
  AOI22_X1 U20611 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17454), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17459), .ZN(n17437) );
  OAI21_X1 U20612 ( .B1(n18168), .B2(n17456), .A(n17437), .ZN(P3_U2785) );
  AOI22_X1 U20613 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17454), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17459), .ZN(n17438) );
  OAI21_X1 U20614 ( .B1(n18172), .B2(n17456), .A(n17438), .ZN(P3_U2786) );
  AOI22_X1 U20615 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17454), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17459), .ZN(n17439) );
  OAI21_X1 U20616 ( .B1(n18177), .B2(n17456), .A(n17439), .ZN(P3_U2787) );
  AOI22_X1 U20617 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17454), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17459), .ZN(n17440) );
  OAI21_X1 U20618 ( .B1(n18181), .B2(n17456), .A(n17440), .ZN(P3_U2788) );
  AOI22_X1 U20619 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17454), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17459), .ZN(n17441) );
  OAI21_X1 U20620 ( .B1(n18186), .B2(n17456), .A(n17441), .ZN(P3_U2789) );
  AOI22_X1 U20621 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(n17454), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17459), .ZN(n17442) );
  OAI21_X1 U20622 ( .B1(n18190), .B2(n17456), .A(n17442), .ZN(P3_U2790) );
  AOI22_X1 U20623 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17454), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17459), .ZN(n17443) );
  OAI21_X1 U20624 ( .B1(n17444), .B2(n17456), .A(n17443), .ZN(P3_U2791) );
  AOI22_X1 U20625 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17454), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17453), .ZN(n17445) );
  OAI21_X1 U20626 ( .B1(n17446), .B2(n17456), .A(n17445), .ZN(P3_U2792) );
  AOI22_X1 U20627 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17454), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17453), .ZN(n17447) );
  OAI21_X1 U20628 ( .B1(n17448), .B2(n17456), .A(n17447), .ZN(P3_U2793) );
  AOI22_X1 U20629 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17460), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17459), .ZN(n17449) );
  OAI21_X1 U20630 ( .B1(n17450), .B2(n17462), .A(n17449), .ZN(P3_U2794) );
  AOI22_X1 U20631 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17454), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17453), .ZN(n17451) );
  OAI21_X1 U20632 ( .B1(n17452), .B2(n17456), .A(n17451), .ZN(P3_U2795) );
  AOI22_X1 U20633 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17454), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17453), .ZN(n17455) );
  OAI21_X1 U20634 ( .B1(n20825), .B2(n17456), .A(n17455), .ZN(P3_U2796) );
  AOI22_X1 U20635 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17460), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17459), .ZN(n17457) );
  OAI21_X1 U20636 ( .B1(n17458), .B2(n17462), .A(n17457), .ZN(P3_U2797) );
  AOI22_X1 U20637 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17460), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17459), .ZN(n17461) );
  OAI21_X1 U20638 ( .B1(n17463), .B2(n17462), .A(n17461), .ZN(P3_U2798) );
  OAI21_X1 U20639 ( .B1(n17464), .B2(n17823), .A(n17822), .ZN(n17465) );
  AOI21_X1 U20640 ( .B1(n18669), .B2(n17467), .A(n17465), .ZN(n17496) );
  OAI21_X1 U20641 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17577), .A(
        n17496), .ZN(n17484) );
  NOR2_X1 U20642 ( .A1(n17690), .A2(n17815), .ZN(n17572) );
  OAI22_X1 U20643 ( .A1(n17837), .A2(n17734), .B1(n17830), .B2(n17827), .ZN(
        n17499) );
  NOR2_X1 U20644 ( .A1(n17829), .A2(n17499), .ZN(n17491) );
  NOR3_X1 U20645 ( .A1(n17572), .A2(n17491), .A3(n17466), .ZN(n17473) );
  NOR2_X1 U20646 ( .A1(n17661), .A2(n17467), .ZN(n17488) );
  OAI211_X1 U20647 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17488), .B(n17468), .ZN(n17470) );
  NAND2_X1 U20648 ( .A1(n18100), .A2(P3_REIP_REG_28__SCAN_IN), .ZN(n17469) );
  OAI211_X1 U20649 ( .C1(n17666), .C2(n17471), .A(n17470), .B(n17469), .ZN(
        n17472) );
  AOI211_X1 U20650 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17484), .A(
        n17473), .B(n17472), .ZN(n17478) );
  OAI211_X1 U20651 ( .C1(n17476), .C2(n17475), .A(n17731), .B(n17474), .ZN(
        n17477) );
  OAI211_X1 U20652 ( .C1(n17479), .C2(n17490), .A(n17478), .B(n17477), .ZN(
        P3_U2802) );
  NAND2_X1 U20653 ( .A1(n17481), .A2(n17480), .ZN(n17482) );
  XOR2_X1 U20654 ( .A(n17482), .B(n17656), .Z(n17844) );
  AOI22_X1 U20655 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17484), .B1(
        n17675), .B2(n17483), .ZN(n17485) );
  NAND2_X1 U20656 ( .A1(n18100), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17842) );
  OAI211_X1 U20657 ( .C1(n17844), .C2(n17721), .A(n17485), .B(n17842), .ZN(
        n17486) );
  AOI21_X1 U20658 ( .B1(n17488), .B2(n17487), .A(n17486), .ZN(n17489) );
  OAI221_X1 U20659 ( .B1(n17491), .B2(n17829), .C1(n17491), .C2(n17490), .A(
        n17489), .ZN(P3_U2803) );
  AOI21_X1 U20660 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17493), .A(
        n17492), .ZN(n17851) );
  NOR2_X1 U20661 ( .A1(n18141), .A2(n18741), .ZN(n17849) );
  NOR2_X2 U20662 ( .A1(n17548), .A2(n17675), .ZN(n17808) );
  AOI21_X1 U20663 ( .B1(n18539), .B2(n17494), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17495) );
  OAI22_X1 U20664 ( .A1(n17808), .A2(n17497), .B1(n17496), .B2(n17495), .ZN(
        n17498) );
  AOI211_X1 U20665 ( .C1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n17499), .A(
        n17849), .B(n17498), .ZN(n17501) );
  INV_X1 U20666 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n20843) );
  NAND3_X1 U20667 ( .A1(n17845), .A2(n17540), .A3(n20843), .ZN(n17500) );
  OAI211_X1 U20668 ( .C1(n17851), .C2(n17721), .A(n17501), .B(n17500), .ZN(
        P3_U2804) );
  XOR2_X1 U20669 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n17502), .Z(
        n17863) );
  NOR2_X1 U20670 ( .A1(n18141), .A2(n18739), .ZN(n17858) );
  INV_X1 U20671 ( .A(n17823), .ZN(n17659) );
  AND2_X1 U20672 ( .A1(n17504), .A2(n18539), .ZN(n17533) );
  AOI211_X1 U20673 ( .C1(n17659), .C2(n17503), .A(n17794), .B(n17533), .ZN(
        n17537) );
  OAI21_X1 U20674 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17577), .A(
        n17537), .ZN(n17521) );
  NOR2_X1 U20675 ( .A1(n17661), .A2(n17504), .ZN(n17523) );
  AOI22_X1 U20676 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n17521), .B1(
        n17523), .B2(n17505), .ZN(n17506) );
  AOI21_X1 U20677 ( .B1(n17522), .B2(n17507), .A(n17506), .ZN(n17508) );
  AOI211_X1 U20678 ( .C1(n17675), .C2(n17509), .A(n17858), .B(n17508), .ZN(
        n17516) );
  AOI21_X1 U20679 ( .B1(n17854), .B2(n17511), .A(n17510), .ZN(n17860) );
  AOI21_X1 U20680 ( .B1(n17513), .B2(n17656), .A(n17512), .ZN(n17514) );
  XOR2_X1 U20681 ( .A(n17514), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17859) );
  AOI22_X1 U20682 ( .A1(n17690), .A2(n17860), .B1(n17731), .B2(n17859), .ZN(
        n17515) );
  OAI211_X1 U20683 ( .C1(n17827), .C2(n17863), .A(n17516), .B(n17515), .ZN(
        P3_U2805) );
  AOI21_X1 U20684 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17518), .A(
        n9609), .ZN(n17876) );
  INV_X1 U20685 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18736) );
  OAI22_X1 U20686 ( .A1(n18141), .A2(n18736), .B1(n17666), .B2(n17519), .ZN(
        n17520) );
  AOI221_X1 U20687 ( .B1(n17523), .B2(n17522), .C1(n17521), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17520), .ZN(n17527) );
  AND2_X1 U20688 ( .A1(n17885), .A2(n17524), .ZN(n17869) );
  NAND2_X1 U20689 ( .A1(n17524), .A2(n17971), .ZN(n17866) );
  INV_X1 U20690 ( .A(n17866), .ZN(n17525) );
  OAI22_X1 U20691 ( .A1(n17869), .A2(n17734), .B1(n17525), .B2(n17827), .ZN(
        n17539) );
  NOR2_X1 U20692 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17870), .ZN(
        n17864) );
  AOI22_X1 U20693 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17539), .B1(
        n17540), .B2(n17864), .ZN(n17526) );
  OAI211_X1 U20694 ( .C1(n17876), .C2(n17721), .A(n17527), .B(n17526), .ZN(
        P3_U2806) );
  AOI22_X1 U20695 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17656), .B1(
        n17528), .B2(n17543), .ZN(n17529) );
  NAND2_X1 U20696 ( .A1(n17573), .A2(n17529), .ZN(n17530) );
  XOR2_X1 U20697 ( .A(n17530), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(
        n17883) );
  AOI22_X1 U20698 ( .A1(n17534), .A2(n17533), .B1(n17532), .B2(n17531), .ZN(
        n17535) );
  NAND2_X1 U20699 ( .A1(n18100), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17882) );
  OAI211_X1 U20700 ( .C1(n17537), .C2(n17536), .A(n17535), .B(n17882), .ZN(
        n17538) );
  AOI221_X1 U20701 ( .B1(n17540), .B2(n17870), .C1(n17539), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n17538), .ZN(n17541) );
  OAI21_X1 U20702 ( .B1(n17721), .B2(n17883), .A(n17541), .ZN(P3_U2807) );
  INV_X1 U20703 ( .A(n17573), .ZN(n17542) );
  AOI221_X1 U20704 ( .B1(n17553), .B2(n17543), .C1(n17559), .C2(n17543), .A(
        n17542), .ZN(n17544) );
  XOR2_X1 U20705 ( .A(n17892), .B(n17544), .Z(n17899) );
  OR2_X1 U20706 ( .A1(n12410), .A2(n17661), .ZN(n17565) );
  AOI211_X1 U20707 ( .C1(n17564), .C2(n17549), .A(n17545), .B(n17565), .ZN(
        n17551) );
  AOI22_X1 U20708 ( .A1(n17659), .A2(n17546), .B1(n18669), .B2(n12410), .ZN(
        n17547) );
  NAND2_X1 U20709 ( .A1(n17547), .A2(n17822), .ZN(n17576) );
  AOI21_X1 U20710 ( .B1(n17548), .B2(n9903), .A(n17576), .ZN(n17563) );
  OAI22_X1 U20711 ( .A1(n17563), .A2(n17549), .B1(n18141), .B2(n18732), .ZN(
        n17550) );
  AOI211_X1 U20712 ( .C1(n17552), .C2(n17675), .A(n17551), .B(n17550), .ZN(
        n17558) );
  INV_X1 U20713 ( .A(n17939), .ZN(n17554) );
  NOR2_X1 U20714 ( .A1(n17554), .A2(n17553), .ZN(n17896) );
  OAI22_X1 U20715 ( .A1(n17734), .A2(n17885), .B1(n17827), .B2(n17971), .ZN(
        n17555) );
  INV_X1 U20716 ( .A(n17555), .ZN(n17625) );
  OAI21_X1 U20717 ( .B1(n17572), .B2(n17896), .A(n17625), .ZN(n17569) );
  NOR2_X1 U20718 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17626), .ZN(
        n17556) );
  AOI22_X1 U20719 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17569), .B1(
        n17896), .B2(n17556), .ZN(n17557) );
  OAI211_X1 U20720 ( .C1(n17721), .C2(n17899), .A(n17558), .B(n17557), .ZN(
        P3_U2808) );
  INV_X1 U20721 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17594) );
  NOR3_X1 U20722 ( .A1(n17656), .A2(n17594), .A3(n17559), .ZN(n17582) );
  INV_X1 U20723 ( .A(n17560), .ZN(n17601) );
  AOI22_X1 U20724 ( .A1(n17568), .A2(n17582), .B1(n17601), .B2(n17561), .ZN(
        n17562) );
  XOR2_X1 U20725 ( .A(n17562), .B(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .Z(
        n17912) );
  NAND2_X1 U20726 ( .A1(n18135), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n17910) );
  OAI221_X1 U20727 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17565), .C1(
        n17564), .C2(n17563), .A(n17910), .ZN(n17566) );
  AOI21_X1 U20728 ( .B1(n17675), .B2(n17567), .A(n17566), .ZN(n17571) );
  INV_X1 U20729 ( .A(n17568), .ZN(n17905) );
  NOR2_X1 U20730 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17905), .ZN(
        n17909) );
  NAND2_X1 U20731 ( .A1(n17939), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17902) );
  NOR2_X1 U20732 ( .A1(n17626), .A2(n17902), .ZN(n17592) );
  AOI22_X1 U20733 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17569), .B1(
        n17909), .B2(n17592), .ZN(n17570) );
  OAI211_X1 U20734 ( .C1(n17912), .C2(n17721), .A(n17571), .B(n17570), .ZN(
        P3_U2809) );
  NOR2_X1 U20735 ( .A1(n17932), .A2(n17902), .ZN(n17915) );
  OAI21_X1 U20736 ( .B1(n17572), .B2(n17915), .A(n17625), .ZN(n17591) );
  OAI221_X1 U20737 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17600), 
        .C1(n17932), .C2(n17582), .A(n17573), .ZN(n17574) );
  XNOR2_X1 U20738 ( .A(n20891), .B(n17574), .ZN(n17925) );
  NAND2_X1 U20739 ( .A1(n17915), .A2(n20891), .ZN(n17919) );
  OAI22_X1 U20740 ( .A1(n17721), .A2(n17925), .B1(n17626), .B2(n17919), .ZN(
        n17575) );
  AOI21_X1 U20741 ( .B1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n17591), .A(
        n17575), .ZN(n17581) );
  NAND2_X1 U20742 ( .A1(n18135), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n17923) );
  OAI221_X1 U20743 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n9677), .C1(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(n18539), .A(n17576), .ZN(
        n17580) );
  OAI21_X1 U20744 ( .B1(n17675), .B2(n17548), .A(n17578), .ZN(n17579) );
  NAND4_X1 U20745 ( .A1(n17581), .A2(n17923), .A3(n17580), .A4(n17579), .ZN(
        P3_U2810) );
  AOI21_X1 U20746 ( .B1(n17601), .B2(n17600), .A(n17582), .ZN(n17583) );
  XOR2_X1 U20747 ( .A(n17583), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Z(
        n17926) );
  AOI21_X1 U20748 ( .B1(n18669), .B2(n17585), .A(n17794), .ZN(n17606) );
  OAI21_X1 U20749 ( .B1(n17584), .B2(n17823), .A(n17606), .ZN(n17597) );
  AOI22_X1 U20750 ( .A1(n18100), .A2(P3_REIP_REG_19__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n17597), .ZN(n17588) );
  NOR2_X1 U20751 ( .A1(n17661), .A2(n17585), .ZN(n17599) );
  OAI211_X1 U20752 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17599), .B(n17586), .ZN(n17587) );
  OAI211_X1 U20753 ( .C1(n17666), .C2(n17589), .A(n17588), .B(n17587), .ZN(
        n17590) );
  AOI221_X1 U20754 ( .B1(n17592), .B2(n17932), .C1(n17591), .C2(
        P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A(n17590), .ZN(n17593) );
  OAI21_X1 U20755 ( .B1(n17926), .B2(n17721), .A(n17593), .ZN(P3_U2811) );
  NAND2_X1 U20756 ( .A1(n17939), .A2(n17594), .ZN(n17946) );
  OAI22_X1 U20757 ( .A1(n18141), .A2(n18724), .B1(n17666), .B2(n17595), .ZN(
        n17596) );
  AOI221_X1 U20758 ( .B1(n17599), .B2(n17598), .C1(n17597), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17596), .ZN(n17604) );
  OAI21_X1 U20759 ( .B1(n17939), .B2(n17626), .A(n17625), .ZN(n17612) );
  AOI21_X1 U20760 ( .B1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n17730), .A(
        n17600), .ZN(n17602) );
  XOR2_X1 U20761 ( .A(n17602), .B(n17601), .Z(n17942) );
  AOI22_X1 U20762 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17612), .B1(
        n17731), .B2(n17942), .ZN(n17603) );
  OAI211_X1 U20763 ( .C1(n17626), .C2(n17946), .A(n17604), .B(n17603), .ZN(
        P3_U2812) );
  NAND2_X1 U20764 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17947), .ZN(
        n17953) );
  AOI21_X1 U20765 ( .B1(n18539), .B2(n17605), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17607) );
  NAND2_X1 U20766 ( .A1(n18135), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n17951) );
  OAI21_X1 U20767 ( .B1(n17607), .B2(n17606), .A(n17951), .ZN(n17608) );
  AOI21_X1 U20768 ( .B1(n17609), .B2(n17531), .A(n17608), .ZN(n17614) );
  OAI21_X1 U20769 ( .B1(n17611), .B2(n17947), .A(n17610), .ZN(n17950) );
  AOI22_X1 U20770 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17612), .B1(
        n17731), .B2(n17950), .ZN(n17613) );
  OAI211_X1 U20771 ( .C1(n17626), .C2(n17953), .A(n17614), .B(n17613), .ZN(
        P3_U2813) );
  NOR2_X1 U20772 ( .A1(n17656), .A2(n17632), .ZN(n17711) );
  INV_X1 U20773 ( .A(n17711), .ZN(n17699) );
  OAI22_X1 U20774 ( .A1(n17730), .A2(n17615), .B1(n17699), .B2(n17831), .ZN(
        n17616) );
  XOR2_X1 U20775 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B(n17616), .Z(
        n17959) );
  AOI21_X1 U20776 ( .B1(n18669), .B2(n17618), .A(n17794), .ZN(n17643) );
  OAI21_X1 U20777 ( .B1(n17617), .B2(n17823), .A(n17643), .ZN(n17629) );
  AOI22_X1 U20778 ( .A1(n18100), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17629), .ZN(n17621) );
  NOR2_X1 U20779 ( .A1(n17661), .A2(n17618), .ZN(n17631) );
  OAI211_X1 U20780 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17631), .B(n17619), .ZN(n17620) );
  OAI211_X1 U20781 ( .C1(n17666), .C2(n17622), .A(n17621), .B(n17620), .ZN(
        n17623) );
  AOI21_X1 U20782 ( .B1(n17731), .B2(n17959), .A(n17623), .ZN(n17624) );
  OAI221_X1 U20783 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17626), 
        .C1(n17962), .C2(n17625), .A(n17624), .ZN(P3_U2814) );
  NOR2_X1 U20784 ( .A1(n17647), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17969) );
  NAND2_X1 U20785 ( .A1(n17690), .A2(n17966), .ZN(n17640) );
  INV_X1 U20786 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17630) );
  NAND2_X1 U20787 ( .A1(n18100), .A2(P3_REIP_REG_15__SCAN_IN), .ZN(n17975) );
  OAI21_X1 U20788 ( .B1(n17666), .B2(n17627), .A(n17975), .ZN(n17628) );
  AOI221_X1 U20789 ( .B1(n17631), .B2(n17630), .C1(n17629), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17628), .ZN(n17639) );
  OAI21_X1 U20790 ( .B1(n17633), .B2(n17632), .A(n9676), .ZN(n17634) );
  OAI221_X1 U20791 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17650), 
        .C1(n18012), .C2(n17730), .A(n17634), .ZN(n17635) );
  XOR2_X1 U20792 ( .A(n12963), .B(n17635), .Z(n17974) );
  NOR2_X1 U20793 ( .A1(n17971), .A2(n17827), .ZN(n17637) );
  NOR2_X1 U20794 ( .A1(n18012), .A2(n18005), .ZN(n17654) );
  INV_X1 U20795 ( .A(n17654), .ZN(n18003) );
  NOR2_X1 U20796 ( .A1(n18016), .A2(n18003), .ZN(n17996) );
  NAND2_X1 U20797 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17996), .ZN(
        n17649) );
  NOR2_X1 U20798 ( .A1(n17650), .A2(n17649), .ZN(n17648) );
  NOR2_X1 U20799 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17648), .ZN(
        n17970) );
  INV_X1 U20800 ( .A(n17970), .ZN(n17636) );
  AOI22_X1 U20801 ( .A1(n17731), .A2(n17974), .B1(n17637), .B2(n17636), .ZN(
        n17638) );
  OAI211_X1 U20802 ( .C1(n17969), .C2(n17640), .A(n17639), .B(n17638), .ZN(
        P3_U2815) );
  NOR3_X1 U20803 ( .A1(n18012), .A2(n18005), .A3(n9935), .ZN(n17980) );
  INV_X1 U20804 ( .A(n17980), .ZN(n17977) );
  OAI22_X1 U20805 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n9676), .B1(
        n17977), .B2(n17699), .ZN(n17641) );
  XOR2_X1 U20806 ( .A(n17650), .B(n17641), .Z(n17991) );
  NAND2_X1 U20807 ( .A1(n18539), .A2(n17642), .ZN(n17687) );
  AOI221_X1 U20808 ( .B1(n17662), .B2(n17644), .C1(n17687), .C2(n17644), .A(
        n17643), .ZN(n17645) );
  NOR2_X1 U20809 ( .A1(n18141), .A2(n18717), .ZN(n17985) );
  AOI211_X1 U20810 ( .C1(n17646), .C2(n17531), .A(n17645), .B(n17985), .ZN(
        n17652) );
  AOI221_X1 U20811 ( .B1(n18014), .B2(n17650), .C1(n17977), .C2(n17650), .A(
        n17647), .ZN(n17986) );
  AOI21_X1 U20812 ( .B1(n17650), .B2(n17649), .A(n17648), .ZN(n17988) );
  AOI22_X1 U20813 ( .A1(n17690), .A2(n17986), .B1(n17815), .B2(n17988), .ZN(
        n17651) );
  OAI211_X1 U20814 ( .C1(n17991), .C2(n17721), .A(n17652), .B(n17651), .ZN(
        P3_U2816) );
  AOI22_X1 U20815 ( .A1(n17654), .A2(n17653), .B1(n17656), .B2(n18012), .ZN(
        n17655) );
  AOI21_X1 U20816 ( .B1(n17656), .B2(n17676), .A(n17655), .ZN(n17657) );
  XOR2_X1 U20817 ( .A(n9935), .B(n17657), .Z(n18001) );
  AOI22_X1 U20818 ( .A1(n17659), .A2(n17658), .B1(n18669), .B2(n16736), .ZN(
        n17660) );
  NAND2_X1 U20819 ( .A1(n17660), .A2(n17822), .ZN(n17673) );
  NOR2_X1 U20820 ( .A1(n17661), .A2(n16736), .ZN(n17672) );
  OAI211_X1 U20821 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17672), .B(n17662), .ZN(n17664) );
  NAND2_X1 U20822 ( .A1(n18135), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17663) );
  OAI211_X1 U20823 ( .C1(n17666), .C2(n17665), .A(n17664), .B(n17663), .ZN(
        n17667) );
  AOI21_X1 U20824 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n17673), .A(
        n17667), .ZN(n17670) );
  NOR2_X1 U20825 ( .A1(n18014), .A2(n18003), .ZN(n17668) );
  OAI22_X1 U20826 ( .A1(n17996), .A2(n17827), .B1(n17668), .B2(n17734), .ZN(
        n17678) );
  NOR2_X1 U20827 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18003), .ZN(
        n17992) );
  AOI22_X1 U20828 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n17678), .B1(
        n17992), .B2(n17717), .ZN(n17669) );
  OAI211_X1 U20829 ( .C1(n17721), .C2(n18001), .A(n17670), .B(n17669), .ZN(
        P3_U2817) );
  AOI22_X1 U20830 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n17673), .B1(
        n17672), .B2(n17671), .ZN(n17683) );
  AOI22_X1 U20831 ( .A1(n18100), .A2(P3_REIP_REG_12__SCAN_IN), .B1(n17675), 
        .B2(n17674), .ZN(n17682) );
  OAI21_X1 U20832 ( .B1(n18005), .B2(n17699), .A(n17676), .ZN(n17677) );
  XOR2_X1 U20833 ( .A(n17677), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n18002) );
  AOI22_X1 U20834 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17678), .B1(
        n17731), .B2(n18002), .ZN(n17681) );
  NAND3_X1 U20835 ( .A1(n17679), .A2(n18012), .A3(n17717), .ZN(n17680) );
  NAND4_X1 U20836 ( .A1(n17683), .A2(n17682), .A3(n17681), .A4(n17680), .ZN(
        P3_U2818) );
  NAND2_X1 U20837 ( .A1(n17822), .A2(n17684), .ZN(n17817) );
  NAND3_X1 U20838 ( .A1(n18539), .A2(n17722), .A3(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17714) );
  NOR2_X1 U20839 ( .A1(n20878), .A2(n17714), .ZN(n17713) );
  NAND2_X1 U20840 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17713), .ZN(
        n17707) );
  OAI21_X1 U20841 ( .B1(n17781), .B2(n17685), .A(n17707), .ZN(n17686) );
  AOI22_X1 U20842 ( .A1(n18100), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n17687), 
        .B2(n17686), .ZN(n17696) );
  NOR2_X1 U20843 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n17692), .ZN(
        n18013) );
  AOI21_X1 U20844 ( .B1(n17711), .B2(n18019), .A(n17688), .ZN(n17689) );
  XOR2_X1 U20845 ( .A(n17689), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(
        n18024) );
  AOI22_X1 U20846 ( .A1(n18014), .A2(n17690), .B1(n17815), .B2(n18016), .ZN(
        n17691) );
  INV_X1 U20847 ( .A(n17691), .ZN(n17718) );
  AOI21_X1 U20848 ( .B1(n17692), .B2(n17717), .A(n17718), .ZN(n17701) );
  OAI22_X1 U20849 ( .A1(n18024), .A2(n17721), .B1(n17701), .B2(n17693), .ZN(
        n17694) );
  AOI21_X1 U20850 ( .B1(n18013), .B2(n17717), .A(n17694), .ZN(n17695) );
  OAI211_X1 U20851 ( .C1(n17808), .C2(n17697), .A(n17696), .B(n17695), .ZN(
        P3_U2819) );
  OAI21_X1 U20852 ( .B1(n18037), .B2(n17699), .A(n17698), .ZN(n17700) );
  XNOR2_X1 U20853 ( .A(n17700), .B(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n18032) );
  INV_X1 U20854 ( .A(n17701), .ZN(n17702) );
  OAI221_X1 U20855 ( .B1(n17717), .B2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), 
        .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(n17702), .ZN(n17703) );
  INV_X1 U20856 ( .A(n17703), .ZN(n17705) );
  NOR2_X1 U20857 ( .A1(n18141), .A2(n18708), .ZN(n17704) );
  AOI211_X1 U20858 ( .C1(n17706), .C2(n17531), .A(n17705), .B(n17704), .ZN(
        n17709) );
  OAI211_X1 U20859 ( .C1(n17713), .C2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n17817), .B(n17707), .ZN(n17708) );
  OAI211_X1 U20860 ( .C1(n18032), .C2(n17721), .A(n17709), .B(n17708), .ZN(
        P3_U2820) );
  NOR2_X1 U20861 ( .A1(n17711), .A2(n17710), .ZN(n17712) );
  XOR2_X1 U20862 ( .A(n17712), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n18044) );
  AOI211_X1 U20863 ( .C1(n17714), .C2(n20878), .A(n17781), .B(n17713), .ZN(
        n17715) );
  NOR2_X1 U20864 ( .A1(n18141), .A2(n18706), .ZN(n18040) );
  AOI211_X1 U20865 ( .C1(n17716), .C2(n17531), .A(n17715), .B(n18040), .ZN(
        n17720) );
  AOI22_X1 U20866 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17718), .B1(
        n17717), .B2(n18037), .ZN(n17719) );
  OAI211_X1 U20867 ( .C1(n18044), .C2(n17721), .A(n17720), .B(n17719), .ZN(
        P3_U2821) );
  AOI21_X1 U20868 ( .B1(n18669), .B2(n17746), .A(n17794), .ZN(n17741) );
  OAI21_X1 U20869 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18264), .A(
        n17741), .ZN(n17726) );
  NOR2_X1 U20870 ( .A1(n18141), .A2(n18705), .ZN(n18053) );
  NAND2_X1 U20871 ( .A1(n18539), .A2(n17722), .ZN(n17723) );
  OAI22_X1 U20872 ( .A1(n17808), .A2(n17724), .B1(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17723), .ZN(n17725) );
  AOI211_X1 U20873 ( .C1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C2(n17726), .A(
        n18053), .B(n17725), .ZN(n17733) );
  AOI21_X1 U20874 ( .B1(n17728), .B2(n18055), .A(n17727), .ZN(n18059) );
  AOI21_X1 U20875 ( .B1(n17730), .B2(n18063), .A(n17729), .ZN(n18057) );
  AOI22_X1 U20876 ( .A1(n17815), .A2(n18059), .B1(n17731), .B2(n18057), .ZN(
        n17732) );
  OAI211_X1 U20877 ( .C1(n17734), .C2(n18063), .A(n17733), .B(n17732), .ZN(
        P3_U2822) );
  NAND2_X1 U20878 ( .A1(n18539), .A2(n9910), .ZN(n17745) );
  AOI22_X1 U20879 ( .A1(n18100), .A2(P3_REIP_REG_7__SCAN_IN), .B1(n17735), 
        .B2(n17531), .ZN(n17744) );
  NAND2_X1 U20880 ( .A1(n17737), .A2(n17736), .ZN(n17738) );
  INV_X1 U20881 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18066) );
  XOR2_X1 U20882 ( .A(n17738), .B(n18066), .Z(n18067) );
  INV_X1 U20883 ( .A(n17797), .ZN(n17826) );
  OAI21_X1 U20884 ( .B1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n17740), .A(
        n17739), .ZN(n18071) );
  OAI22_X1 U20885 ( .A1(n17826), .A2(n18071), .B1(n9910), .B2(n17741), .ZN(
        n17742) );
  AOI21_X1 U20886 ( .B1(n17815), .B2(n18067), .A(n17742), .ZN(n17743) );
  OAI211_X1 U20887 ( .C1(n17746), .C2(n17745), .A(n17744), .B(n17743), .ZN(
        P3_U2823) );
  NAND2_X1 U20888 ( .A1(n18539), .A2(n17749), .ZN(n17757) );
  AOI21_X1 U20889 ( .B1(n18077), .B2(n17748), .A(n17747), .ZN(n18075) );
  AOI22_X1 U20890 ( .A1(n17815), .A2(n18075), .B1(n18135), .B2(
        P3_REIP_REG_6__SCAN_IN), .ZN(n17756) );
  AOI21_X1 U20891 ( .B1(n17749), .B2(n18539), .A(n17781), .ZN(n17768) );
  OAI21_X1 U20892 ( .B1(n17752), .B2(n17751), .A(n17750), .ZN(n18073) );
  OAI22_X1 U20893 ( .A1(n17808), .A2(n17753), .B1(n17826), .B2(n18073), .ZN(
        n17754) );
  AOI21_X1 U20894 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17768), .A(
        n17754), .ZN(n17755) );
  OAI211_X1 U20895 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n17757), .A(
        n17756), .B(n17755), .ZN(P3_U2824) );
  AOI21_X1 U20896 ( .B1(n17760), .B2(n17759), .A(n17758), .ZN(n17761) );
  XOR2_X1 U20897 ( .A(n17761), .B(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(
        n18079) );
  AOI22_X1 U20898 ( .A1(n17797), .A2(n18079), .B1(n18135), .B2(
        P3_REIP_REG_5__SCAN_IN), .ZN(n17770) );
  AOI21_X1 U20899 ( .B1(n17764), .B2(n17763), .A(n17762), .ZN(n18082) );
  OAI21_X1 U20900 ( .B1(n17794), .B2(n17766), .A(n17765), .ZN(n17767) );
  AOI22_X1 U20901 ( .A1(n17815), .A2(n18082), .B1(n17768), .B2(n17767), .ZN(
        n17769) );
  OAI211_X1 U20902 ( .C1(n17808), .C2(n17771), .A(n17770), .B(n17769), .ZN(
        P3_U2825) );
  OAI21_X1 U20903 ( .B1(n17774), .B2(n17773), .A(n17772), .ZN(n18097) );
  OAI21_X1 U20904 ( .B1(n17777), .B2(n17776), .A(n17775), .ZN(n17778) );
  XOR2_X1 U20905 ( .A(n17778), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(
        n18091) );
  OAI22_X1 U20906 ( .A1(n17827), .A2(n18091), .B1(n18264), .B2(n17779), .ZN(
        n17780) );
  AOI21_X1 U20907 ( .B1(n18135), .B2(P3_REIP_REG_4__SCAN_IN), .A(n17780), .ZN(
        n17785) );
  AOI21_X1 U20908 ( .B1(n17782), .B2(n17822), .A(n17781), .ZN(n17796) );
  AOI22_X1 U20909 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17796), .B1(
        n17783), .B2(n17531), .ZN(n17784) );
  OAI211_X1 U20910 ( .C1(n17826), .C2(n18097), .A(n17785), .B(n17784), .ZN(
        P3_U2826) );
  AOI21_X1 U20911 ( .B1(n17788), .B2(n17787), .A(n17786), .ZN(n18101) );
  AOI22_X1 U20912 ( .A1(n17815), .A2(n18101), .B1(n18135), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n17799) );
  AOI21_X1 U20913 ( .B1(n17791), .B2(n17790), .A(n17789), .ZN(n17792) );
  XOR2_X1 U20914 ( .A(n17792), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(
        n18099) );
  OAI21_X1 U20915 ( .B1(n17794), .B2(n17811), .A(n17793), .ZN(n17795) );
  AOI22_X1 U20916 ( .A1(n17797), .A2(n18099), .B1(n17796), .B2(n17795), .ZN(
        n17798) );
  OAI211_X1 U20917 ( .C1(n17808), .C2(n17800), .A(n17799), .B(n17798), .ZN(
        P3_U2827) );
  AOI21_X1 U20918 ( .B1(n17803), .B2(n17802), .A(n17801), .ZN(n18119) );
  NOR2_X1 U20919 ( .A1(n18141), .A2(n18692), .ZN(n18120) );
  OAI21_X1 U20920 ( .B1(n17806), .B2(n17805), .A(n17804), .ZN(n18106) );
  OAI22_X1 U20921 ( .A1(n17808), .A2(n17807), .B1(n17826), .B2(n18106), .ZN(
        n17809) );
  AOI211_X1 U20922 ( .C1(n17815), .C2(n18119), .A(n18120), .B(n17809), .ZN(
        n17810) );
  OAI221_X1 U20923 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18264), .C1(
        n17811), .C2(n17822), .A(n17810), .ZN(P3_U2828) );
  OAI21_X1 U20924 ( .B1(n17820), .B2(n17813), .A(n17812), .ZN(n18134) );
  NAND2_X1 U20925 ( .A1(n18790), .A2(n17821), .ZN(n17814) );
  XNOR2_X1 U20926 ( .A(n17814), .B(n17813), .ZN(n18130) );
  AOI22_X1 U20927 ( .A1(n17815), .A2(n18130), .B1(n18135), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17819) );
  AOI22_X1 U20928 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17817), .B1(
        n17531), .B2(n17816), .ZN(n17818) );
  OAI211_X1 U20929 ( .C1(n17826), .C2(n18134), .A(n17819), .B(n17818), .ZN(
        P3_U2829) );
  AOI21_X1 U20930 ( .B1(n17821), .B2(n18790), .A(n17820), .ZN(n18139) );
  INV_X1 U20931 ( .A(n18139), .ZN(n18137) );
  NAND3_X1 U20932 ( .A1(n18773), .A2(n17823), .A3(n17822), .ZN(n17824) );
  AOI22_X1 U20933 ( .A1(n18135), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17824), .ZN(n17825) );
  OAI221_X1 U20934 ( .B1(n18139), .B2(n17827), .C1(n18137), .C2(n17826), .A(
        n17825), .ZN(P3_U2830) );
  OAI21_X1 U20935 ( .B1(n18142), .B2(n17829), .A(n17828), .ZN(n17841) );
  INV_X1 U20936 ( .A(n17830), .ZN(n17839) );
  INV_X1 U20937 ( .A(n17853), .ZN(n17833) );
  NAND2_X1 U20938 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17954), .ZN(
        n18034) );
  NOR2_X1 U20939 ( .A1(n17831), .A2(n18034), .ZN(n17900) );
  AOI21_X1 U20940 ( .B1(n17900), .B2(n17896), .A(n18616), .ZN(n17891) );
  AOI21_X1 U20941 ( .B1(n18089), .B2(n17832), .A(n17891), .ZN(n17868) );
  OAI21_X1 U20942 ( .B1(n18110), .B2(n17833), .A(n17868), .ZN(n17852) );
  AOI22_X1 U20943 ( .A1(n18605), .A2(n17854), .B1(n18629), .B2(n17834), .ZN(
        n17836) );
  OAI211_X1 U20944 ( .C1(n17837), .C2(n17884), .A(n17836), .B(n17835), .ZN(
        n17838) );
  AOI211_X1 U20945 ( .C1(n18594), .C2(n17839), .A(n17852), .B(n17838), .ZN(
        n17847) );
  OAI211_X1 U20946 ( .C1(n18631), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n17847), .ZN(n17840) );
  AOI22_X1 U20947 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18121), .B1(
        n17841), .B2(n17840), .ZN(n17843) );
  OAI211_X1 U20948 ( .C1(n17844), .C2(n18043), .A(n17843), .B(n17842), .ZN(
        P3_U2835) );
  AOI22_X1 U20949 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18125), .B1(
        n17845), .B2(n17865), .ZN(n17846) );
  AOI21_X1 U20950 ( .B1(n17847), .B2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n17846), .ZN(n17848) );
  AOI211_X1 U20951 ( .C1(n18121), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n17849), .B(n17848), .ZN(n17850) );
  OAI21_X1 U20952 ( .B1(n17851), .B2(n18043), .A(n17850), .ZN(P3_U2836) );
  AOI221_X1 U20953 ( .B1(n17871), .B2(n18627), .C1(n17853), .C2(n18627), .A(
        n17852), .ZN(n17856) );
  AOI221_X1 U20954 ( .B1(n17856), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), 
        .C1(n17855), .C2(n17854), .A(n18142), .ZN(n17857) );
  AOI211_X1 U20955 ( .C1(n18121), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17858), .B(n17857), .ZN(n17862) );
  AOI22_X1 U20956 ( .A1(n17987), .A2(n17860), .B1(n18058), .B2(n17859), .ZN(
        n17861) );
  OAI211_X1 U20957 ( .C1(n18090), .C2(n17863), .A(n17862), .B(n17861), .ZN(
        P3_U2837) );
  AOI22_X1 U20958 ( .A1(n18100), .A2(P3_REIP_REG_24__SCAN_IN), .B1(n17865), 
        .B2(n17864), .ZN(n17875) );
  AOI21_X1 U20959 ( .B1(n18594), .B2(n17866), .A(n18121), .ZN(n17867) );
  OAI211_X1 U20960 ( .C1(n17869), .C2(n17884), .A(n17868), .B(n17867), .ZN(
        n17873) );
  AOI211_X1 U20961 ( .C1(n18627), .C2(n17871), .A(n17870), .B(n17873), .ZN(
        n17872) );
  NOR2_X1 U20962 ( .A1(n18135), .A2(n17872), .ZN(n17879) );
  OAI211_X1 U20963 ( .C1(n18052), .C2(n17873), .A(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n17879), .ZN(n17874) );
  OAI211_X1 U20964 ( .C1(n17876), .C2(n18043), .A(n17875), .B(n17874), .ZN(
        P3_U2838) );
  NOR3_X1 U20965 ( .A1(n18121), .A2(n17878), .A3(n17877), .ZN(n17880) );
  OAI21_X1 U20966 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17880), .A(
        n17879), .ZN(n17881) );
  OAI211_X1 U20967 ( .C1(n17883), .C2(n18043), .A(n17882), .B(n17881), .ZN(
        P3_U2839) );
  NAND2_X1 U20968 ( .A1(n18135), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17898) );
  OAI22_X1 U20969 ( .A1(n17885), .A2(n17884), .B1(n17971), .B2(n17995), .ZN(
        n17901) );
  NOR2_X1 U20970 ( .A1(n18594), .A2(n18015), .ZN(n18018) );
  OAI21_X1 U20971 ( .B1(n17886), .B2(n17902), .A(n18627), .ZN(n17887) );
  OAI221_X1 U20972 ( .B1(n18631), .B2(n17937), .C1(n18631), .C2(n17915), .A(
        n17887), .ZN(n17913) );
  AOI21_X1 U20973 ( .B1(n18605), .B2(n20891), .A(n17913), .ZN(n17888) );
  OAI21_X1 U20974 ( .B1(n17896), .B2(n18018), .A(n17888), .ZN(n17904) );
  AOI22_X1 U20975 ( .A1(n18627), .A2(n17905), .B1(n17906), .B2(n17993), .ZN(
        n17889) );
  NAND2_X1 U20976 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17889), .ZN(
        n17890) );
  NOR4_X1 U20977 ( .A1(n17891), .A2(n17901), .A3(n17904), .A4(n17890), .ZN(
        n17893) );
  OAI22_X1 U20978 ( .A1(n17893), .A2(n18142), .B1(n17892), .B2(n18126), .ZN(
        n17894) );
  OAI221_X1 U20979 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n17896), 
        .C1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .C2(n17895), .A(n17894), .ZN(
        n17897) );
  OAI211_X1 U20980 ( .C1(n17899), .C2(n18043), .A(n17898), .B(n17897), .ZN(
        P3_U2840) );
  NOR2_X1 U20981 ( .A1(n17920), .A2(n17902), .ZN(n17927) );
  NAND2_X1 U20982 ( .A1(n18616), .A2(n18108), .ZN(n18124) );
  INV_X1 U20983 ( .A(n17900), .ZN(n17956) );
  OR2_X1 U20984 ( .A1(n18142), .A2(n17901), .ZN(n17958) );
  AOI221_X1 U20985 ( .B1(n18629), .B2(n17956), .C1(n18629), .C2(n17902), .A(
        n17958), .ZN(n17903) );
  INV_X1 U20986 ( .A(n17903), .ZN(n17917) );
  AOI211_X1 U20987 ( .C1(n17905), .C2(n18124), .A(n17917), .B(n17904), .ZN(
        n17907) );
  NOR3_X1 U20988 ( .A1(n18100), .A2(n17907), .A3(n17906), .ZN(n17908) );
  AOI21_X1 U20989 ( .B1(n17927), .B2(n17909), .A(n17908), .ZN(n17911) );
  OAI211_X1 U20990 ( .C1(n17912), .C2(n18043), .A(n17911), .B(n17910), .ZN(
        P3_U2841) );
  NAND3_X1 U20991 ( .A1(n17932), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(n18124), 
        .ZN(n17918) );
  INV_X1 U20992 ( .A(n17913), .ZN(n17914) );
  OAI21_X1 U20993 ( .B1(n17915), .B2(n18018), .A(n17914), .ZN(n17916) );
  OAI21_X1 U20994 ( .B1(n17917), .B2(n17916), .A(n18141), .ZN(n17931) );
  AND2_X1 U20995 ( .A1(n17918), .A2(n17931), .ZN(n17921) );
  OAI22_X1 U20996 ( .A1(n20891), .A2(n17921), .B1(n17920), .B2(n17919), .ZN(
        n17922) );
  INV_X1 U20997 ( .A(n17922), .ZN(n17924) );
  OAI211_X1 U20998 ( .C1(n17925), .C2(n18043), .A(n17924), .B(n17923), .ZN(
        P3_U2842) );
  INV_X1 U20999 ( .A(n17926), .ZN(n17928) );
  AOI22_X1 U21000 ( .A1(n18058), .A2(n17928), .B1(n17927), .B2(n17932), .ZN(
        n17930) );
  NAND2_X1 U21001 ( .A1(n18135), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17929) );
  OAI211_X1 U21002 ( .C1(n17932), .C2(n17931), .A(n17930), .B(n17929), .ZN(
        P3_U2843) );
  NAND2_X1 U21003 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18088) );
  OAI22_X1 U21004 ( .A1(n17933), .A2(n18108), .B1(n18109), .B2(n18088), .ZN(
        n18098) );
  NAND2_X1 U21005 ( .A1(n18045), .A2(n18098), .ZN(n18065) );
  NOR2_X1 U21006 ( .A1(n17934), .A2(n18065), .ZN(n17981) );
  NOR2_X1 U21007 ( .A1(n17981), .A2(n17935), .ZN(n18006) );
  NAND2_X1 U21008 ( .A1(n17936), .A2(n18038), .ZN(n17963) );
  NOR2_X1 U21009 ( .A1(n18616), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18048) );
  INV_X1 U21010 ( .A(n18048), .ZN(n18111) );
  NAND3_X1 U21011 ( .A1(n17937), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n18111), .ZN(n17941) );
  AOI222_X1 U21012 ( .A1(n17939), .A2(n18108), .B1(n17939), .B2(n17938), .C1(
        n18108), .C2(n18018), .ZN(n17940) );
  AOI211_X1 U21013 ( .C1(n18089), .C2(n17941), .A(n17940), .B(n17958), .ZN(
        n17948) );
  AOI221_X1 U21014 ( .B1(n18110), .B2(n17948), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n17948), .A(n18100), .ZN(
        n17943) );
  AOI22_X1 U21015 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17943), .B1(
        n18058), .B2(n17942), .ZN(n17945) );
  NAND2_X1 U21016 ( .A1(n18135), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17944) );
  OAI211_X1 U21017 ( .C1(n17946), .C2(n17963), .A(n17945), .B(n17944), .ZN(
        P3_U2844) );
  NOR3_X1 U21018 ( .A1(n18135), .A2(n17948), .A3(n17947), .ZN(n17949) );
  AOI21_X1 U21019 ( .B1(n18058), .B2(n17950), .A(n17949), .ZN(n17952) );
  OAI211_X1 U21020 ( .C1(n17963), .C2(n17953), .A(n17952), .B(n17951), .ZN(
        P3_U2845) );
  OAI22_X1 U21021 ( .A1(n18108), .A2(n17955), .B1(n18631), .B2(n17954), .ZN(
        n18033) );
  INV_X1 U21022 ( .A(n18033), .ZN(n18026) );
  OAI21_X1 U21023 ( .B1(n12963), .B2(n18629), .A(n17956), .ZN(n17957) );
  OAI211_X1 U21024 ( .C1(n17965), .C2(n18027), .A(n18026), .B(n17957), .ZN(
        n17964) );
  OAI221_X1 U21025 ( .B1(n17958), .B2(n18052), .C1(n17958), .C2(n17964), .A(
        n18141), .ZN(n17961) );
  AOI22_X1 U21026 ( .A1(n18100), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n18058), 
        .B2(n17959), .ZN(n17960) );
  OAI221_X1 U21027 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17963), 
        .C1(n17962), .C2(n17961), .A(n17960), .ZN(P3_U2846) );
  OAI221_X1 U21028 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n17965), 
        .C1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n17981), .A(n17964), .ZN(
        n17968) );
  NAND2_X1 U21029 ( .A1(n18015), .A2(n17966), .ZN(n17967) );
  AOI221_X1 U21030 ( .B1(n17969), .B2(n17968), .C1(n17967), .C2(n17968), .A(
        n18142), .ZN(n17973) );
  NOR3_X1 U21031 ( .A1(n17971), .A2(n17970), .A3(n18090), .ZN(n17972) );
  AOI211_X1 U21032 ( .C1(n18058), .C2(n17974), .A(n17973), .B(n17972), .ZN(
        n17976) );
  OAI211_X1 U21033 ( .C1(n18126), .C2(n12963), .A(n17976), .B(n17975), .ZN(
        P3_U2847) );
  AOI22_X1 U21034 ( .A1(n18627), .A2(n18003), .B1(n18605), .B2(n17977), .ZN(
        n17978) );
  OAI21_X1 U21035 ( .B1(n18034), .B2(n18003), .A(n18629), .ZN(n17997) );
  NAND4_X1 U21036 ( .A1(n18026), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        n17978), .A4(n17997), .ZN(n17979) );
  AOI21_X1 U21037 ( .B1(n9935), .B2(n18124), .A(n17979), .ZN(n17983) );
  AOI21_X1 U21038 ( .B1(n17981), .B2(n17980), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17982) );
  NOR3_X1 U21039 ( .A1(n17983), .A2(n17982), .A3(n18142), .ZN(n17984) );
  AOI211_X1 U21040 ( .C1(n18121), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17985), .B(n17984), .ZN(n17990) );
  AOI22_X1 U21041 ( .A1(n18138), .A2(n17988), .B1(n17987), .B2(n17986), .ZN(
        n17989) );
  OAI211_X1 U21042 ( .C1(n17991), .C2(n18043), .A(n17990), .B(n17989), .ZN(
        P3_U2848) );
  AOI22_X1 U21043 ( .A1(n18135), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18038), 
        .B2(n17992), .ZN(n18000) );
  OAI21_X1 U21044 ( .B1(n18005), .B2(n18033), .A(n17993), .ZN(n18020) );
  OAI21_X1 U21045 ( .B1(n18014), .B2(n18003), .A(n18015), .ZN(n17994) );
  OAI211_X1 U21046 ( .C1(n17996), .C2(n17995), .A(n18020), .B(n17994), .ZN(
        n18008) );
  OAI211_X1 U21047 ( .C1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n18027), .A(
        n18125), .B(n17997), .ZN(n17998) );
  OAI211_X1 U21048 ( .C1(n18008), .C2(n17998), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n18141), .ZN(n17999) );
  OAI211_X1 U21049 ( .C1(n18001), .C2(n18043), .A(n18000), .B(n17999), .ZN(
        P3_U2849) );
  AOI22_X1 U21050 ( .A1(n18100), .A2(P3_REIP_REG_12__SCAN_IN), .B1(n18058), 
        .B2(n18002), .ZN(n18011) );
  NOR2_X1 U21051 ( .A1(n18034), .A2(n18003), .ZN(n18004) );
  AOI21_X1 U21052 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18616), .A(
        n18004), .ZN(n18009) );
  OAI21_X1 U21053 ( .B1(n18006), .B2(n18005), .A(n18012), .ZN(n18007) );
  OAI211_X1 U21054 ( .C1(n18009), .C2(n18008), .A(n18125), .B(n18007), .ZN(
        n18010) );
  OAI211_X1 U21055 ( .C1(n18126), .C2(n18012), .A(n18011), .B(n18010), .ZN(
        P3_U2850) );
  AOI22_X1 U21056 ( .A1(n18100), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18038), 
        .B2(n18013), .ZN(n18023) );
  AOI22_X1 U21057 ( .A1(n18594), .A2(n18016), .B1(n18015), .B2(n18014), .ZN(
        n18036) );
  OAI21_X1 U21058 ( .B1(n18037), .B2(n18034), .A(n18629), .ZN(n18017) );
  OAI211_X1 U21059 ( .C1(n18019), .C2(n18018), .A(n18036), .B(n18017), .ZN(
        n18029) );
  OAI211_X1 U21060 ( .C1(n18616), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n18125), .B(n18020), .ZN(n18021) );
  OAI211_X1 U21061 ( .C1(n18029), .C2(n18021), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n18141), .ZN(n18022) );
  OAI211_X1 U21062 ( .C1(n18024), .C2(n18043), .A(n18023), .B(n18022), .ZN(
        P3_U2851) );
  NOR2_X1 U21063 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n18037), .ZN(
        n18025) );
  AOI22_X1 U21064 ( .A1(n18100), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n18038), 
        .B2(n18025), .ZN(n18031) );
  OAI211_X1 U21065 ( .C1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n18027), .A(
        n18125), .B(n18026), .ZN(n18028) );
  OAI211_X1 U21066 ( .C1(n18029), .C2(n18028), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B(n18141), .ZN(n18030) );
  OAI211_X1 U21067 ( .C1(n18032), .C2(n18043), .A(n18031), .B(n18030), .ZN(
        P3_U2852) );
  AOI211_X1 U21068 ( .C1(n18629), .C2(n18034), .A(n18142), .B(n18033), .ZN(
        n18035) );
  AOI21_X1 U21069 ( .B1(n18036), .B2(n18035), .A(n18135), .ZN(n18039) );
  AOI22_X1 U21070 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18039), .B1(
        n18038), .B2(n18037), .ZN(n18042) );
  INV_X1 U21071 ( .A(n18040), .ZN(n18041) );
  OAI211_X1 U21072 ( .C1(n18044), .C2(n18043), .A(n18042), .B(n18041), .ZN(
        P3_U2853) );
  NAND2_X1 U21073 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18051) );
  NAND3_X1 U21074 ( .A1(n18045), .A2(n18125), .A3(n18098), .ZN(n18078) );
  NOR2_X1 U21075 ( .A1(n18051), .A2(n18078), .ZN(n18056) );
  INV_X1 U21076 ( .A(n18046), .ZN(n18050) );
  OAI21_X1 U21077 ( .B1(n18048), .B2(n18047), .A(n18089), .ZN(n18049) );
  OAI21_X1 U21078 ( .B1(n18050), .B2(n18108), .A(n18049), .ZN(n18072) );
  AOI21_X1 U21079 ( .B1(n18052), .B2(n18051), .A(n18072), .ZN(n18064) );
  OAI21_X1 U21080 ( .B1(n18064), .B2(n18127), .A(n18126), .ZN(n18054) );
  AOI221_X1 U21081 ( .B1(n18056), .B2(n18055), .C1(n18054), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18053), .ZN(n18061) );
  AOI22_X1 U21082 ( .A1(n18138), .A2(n18059), .B1(n18058), .B2(n18057), .ZN(
        n18060) );
  OAI211_X1 U21083 ( .C1(n18063), .C2(n18062), .A(n18061), .B(n18060), .ZN(
        P3_U2854) );
  INV_X1 U21084 ( .A(n18140), .ZN(n18133) );
  AOI22_X1 U21085 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n18121), .B1(
        n18135), .B2(P3_REIP_REG_7__SCAN_IN), .ZN(n18070) );
  AOI221_X1 U21086 ( .B1(n18077), .B2(n18066), .C1(n18065), .C2(n18066), .A(
        n18064), .ZN(n18068) );
  AOI22_X1 U21087 ( .A1(n18125), .A2(n18068), .B1(n18138), .B2(n18067), .ZN(
        n18069) );
  OAI211_X1 U21088 ( .C1(n18133), .C2(n18071), .A(n18070), .B(n18069), .ZN(
        P3_U2855) );
  OAI21_X1 U21089 ( .B1(n18142), .B2(n18072), .A(n18141), .ZN(n18085) );
  OAI22_X1 U21090 ( .A1(n18141), .A2(n18700), .B1(n18133), .B2(n18073), .ZN(
        n18074) );
  AOI21_X1 U21091 ( .B1(n18138), .B2(n18075), .A(n18074), .ZN(n18076) );
  OAI221_X1 U21092 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18078), .C1(
        n18077), .C2(n18085), .A(n18076), .ZN(P3_U2856) );
  AOI22_X1 U21093 ( .A1(n18100), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18140), 
        .B2(n18079), .ZN(n18084) );
  NAND3_X1 U21094 ( .A1(n18125), .A2(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n18098), .ZN(n18092) );
  NOR3_X1 U21095 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18080), .A3(
        n18092), .ZN(n18081) );
  AOI21_X1 U21096 ( .B1(n18082), .B2(n18138), .A(n18081), .ZN(n18083) );
  OAI211_X1 U21097 ( .C1(n18086), .C2(n18085), .A(n18084), .B(n18083), .ZN(
        P3_U2857) );
  OAI211_X1 U21098 ( .C1(n18108), .C2(n18107), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n18111), .ZN(n18087) );
  AOI21_X1 U21099 ( .B1(n18089), .B2(n18088), .A(n18087), .ZN(n18105) );
  OAI21_X1 U21100 ( .B1(n18105), .B2(n18127), .A(n18126), .ZN(n18094) );
  OAI22_X1 U21101 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18092), .B1(
        n18091), .B2(n18090), .ZN(n18093) );
  AOI21_X1 U21102 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n18094), .A(
        n18093), .ZN(n18096) );
  NAND2_X1 U21103 ( .A1(n18135), .A2(P3_REIP_REG_4__SCAN_IN), .ZN(n18095) );
  OAI211_X1 U21104 ( .C1(n18097), .C2(n18133), .A(n18096), .B(n18095), .ZN(
        P3_U2858) );
  OAI21_X1 U21105 ( .B1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n18098), .A(
        n18125), .ZN(n18104) );
  AOI22_X1 U21106 ( .A1(n18100), .A2(P3_REIP_REG_3__SCAN_IN), .B1(n18140), 
        .B2(n18099), .ZN(n18103) );
  AOI22_X1 U21107 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18121), .B1(
        n18138), .B2(n18101), .ZN(n18102) );
  OAI211_X1 U21108 ( .C1(n18105), .C2(n18104), .A(n18103), .B(n18102), .ZN(
        P3_U2859) );
  OAI22_X1 U21109 ( .A1(n18108), .A2(n18107), .B1(n18600), .B2(n18106), .ZN(
        n18118) );
  INV_X1 U21110 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18771) );
  NOR2_X1 U21111 ( .A1(n18771), .A2(n18109), .ZN(n18116) );
  NOR2_X1 U21112 ( .A1(n18771), .A2(n18790), .ZN(n18113) );
  AOI21_X1 U21113 ( .B1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n18111), .A(
        n18110), .ZN(n18112) );
  AOI21_X1 U21114 ( .B1(n18113), .B2(n18627), .A(n18112), .ZN(n18114) );
  INV_X1 U21115 ( .A(n18114), .ZN(n18115) );
  MUX2_X1 U21116 ( .A(n18116), .B(n18115), .S(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n18117) );
  AOI211_X1 U21117 ( .C1(n18594), .C2(n18119), .A(n18118), .B(n18117), .ZN(
        n18123) );
  AOI21_X1 U21118 ( .B1(n18121), .B2(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A(
        n18120), .ZN(n18122) );
  OAI21_X1 U21119 ( .B1(n18123), .B2(n18142), .A(n18122), .ZN(P3_U2860) );
  NAND3_X1 U21120 ( .A1(n18125), .A2(n18790), .A3(n18124), .ZN(n18144) );
  AOI21_X1 U21121 ( .B1(n18126), .B2(n18144), .A(n18771), .ZN(n18129) );
  AOI211_X1 U21122 ( .C1(n18631), .C2(n18790), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B(n18127), .ZN(n18128) );
  AOI211_X1 U21123 ( .C1(n18138), .C2(n18130), .A(n18129), .B(n18128), .ZN(
        n18132) );
  NAND2_X1 U21124 ( .A1(n18135), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18131) );
  OAI211_X1 U21125 ( .C1(n18134), .C2(n18133), .A(n18132), .B(n18131), .ZN(
        P3_U2861) );
  AND2_X1 U21126 ( .A1(n18135), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18136) );
  AOI221_X1 U21127 ( .B1(n18140), .B2(n18139), .C1(n18138), .C2(n18137), .A(
        n18136), .ZN(n18145) );
  OAI211_X1 U21128 ( .C1(n18605), .C2(n18142), .A(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B(n18141), .ZN(n18143) );
  NAND3_X1 U21129 ( .A1(n18145), .A2(n18144), .A3(n18143), .ZN(P3_U2862) );
  AOI211_X1 U21130 ( .C1(n18147), .C2(n18146), .A(n18661), .B(n18773), .ZN(
        n18655) );
  OAI21_X1 U21131 ( .B1(n18655), .B2(n18197), .A(n18153), .ZN(n18148) );
  OAI221_X1 U21132 ( .B1(n18634), .B2(n18149), .C1(n18634), .C2(n18153), .A(
        n18148), .ZN(P3_U2863) );
  NAND2_X1 U21133 ( .A1(n20792), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18287) );
  NAND2_X1 U21134 ( .A1(n18641), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18421) );
  INV_X1 U21135 ( .A(n18421), .ZN(n18397) );
  NAND2_X1 U21136 ( .A1(n18504), .A2(n18397), .ZN(n18448) );
  AND2_X1 U21137 ( .A1(n18287), .A2(n18448), .ZN(n18151) );
  OAI22_X1 U21138 ( .A1(n18152), .A2(n20792), .B1(n18151), .B2(n18150), .ZN(
        P3_U2866) );
  INV_X1 U21139 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18644) );
  NOR2_X1 U21140 ( .A1(n18644), .A2(n18153), .ZN(P3_U2867) );
  NAND2_X1 U21141 ( .A1(n18539), .A2(BUF2_REG_16__SCAN_IN), .ZN(n18509) );
  NAND2_X1 U21142 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18156) );
  INV_X1 U21143 ( .A(n18156), .ZN(n18476) );
  NOR2_X1 U21144 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18636), .ZN(
        n18398) );
  NAND2_X1 U21145 ( .A1(n18476), .A2(n18398), .ZN(n18208) );
  NOR2_X1 U21146 ( .A1(n18156), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18538) );
  NAND2_X1 U21147 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18538), .ZN(
        n18576) );
  INV_X1 U21148 ( .A(n18576), .ZN(n18586) );
  NOR2_X2 U21149 ( .A1(n18154), .A2(n18264), .ZN(n18540) );
  NOR2_X2 U21150 ( .A1(n18262), .A2(n18155), .ZN(n18534) );
  INV_X1 U21151 ( .A(n18533), .ZN(n18662) );
  NOR2_X1 U21152 ( .A1(n20792), .A2(n18330), .ZN(n18537) );
  NAND2_X1 U21153 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18537), .ZN(
        n18544) );
  NOR2_X1 U21154 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18261) );
  NOR2_X1 U21155 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18240) );
  NAND2_X1 U21156 ( .A1(n18261), .A2(n18240), .ZN(n18260) );
  NAND2_X1 U21157 ( .A1(n18544), .A2(n18260), .ZN(n18157) );
  INV_X1 U21158 ( .A(n18157), .ZN(n18217) );
  NOR2_X1 U21159 ( .A1(n18662), .A2(n18217), .ZN(n18191) );
  AOI22_X1 U21160 ( .A1(n18586), .A2(n18540), .B1(n18534), .B2(n18191), .ZN(
        n18162) );
  NOR2_X1 U21161 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18634), .ZN(
        n18374) );
  NOR2_X1 U21162 ( .A1(n18398), .A2(n18374), .ZN(n18449) );
  NOR2_X1 U21163 ( .A1(n18449), .A2(n18156), .ZN(n18505) );
  AOI21_X1 U21164 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18262), .ZN(n18502) );
  AOI22_X1 U21165 ( .A1(n18539), .A2(n18505), .B1(n18502), .B2(n18157), .ZN(
        n18194) );
  INV_X1 U21166 ( .A(n18260), .ZN(n18253) );
  NAND2_X1 U21167 ( .A1(n18159), .A2(n18158), .ZN(n18192) );
  NOR2_X1 U21168 ( .A1(n18160), .A2(n18192), .ZN(n18506) );
  AOI22_X1 U21169 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18194), .B1(
        n18253), .B2(n18506), .ZN(n18161) );
  OAI211_X1 U21170 ( .C1(n18509), .C2(n18208), .A(n18162), .B(n18161), .ZN(
        P3_U2868) );
  INV_X1 U21171 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n18163) );
  NOR2_X1 U21172 ( .A1(n18264), .A2(n18163), .ZN(n18546) );
  INV_X1 U21173 ( .A(n18546), .ZN(n18483) );
  NAND2_X1 U21174 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n18539), .ZN(n18550) );
  INV_X1 U21175 ( .A(n18550), .ZN(n18480) );
  NOR2_X2 U21176 ( .A1(n18262), .A2(n20810), .ZN(n18545) );
  AOI22_X1 U21177 ( .A1(n18586), .A2(n18480), .B1(n18191), .B2(n18545), .ZN(
        n18166) );
  NOR2_X2 U21178 ( .A1(n18164), .A2(n18192), .ZN(n18547) );
  AOI22_X1 U21179 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18194), .B1(
        n18253), .B2(n18547), .ZN(n18165) );
  OAI211_X1 U21180 ( .C1(n18208), .C2(n18483), .A(n18166), .B(n18165), .ZN(
        P3_U2869) );
  INV_X1 U21181 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n18167) );
  NOR2_X1 U21182 ( .A1(n18264), .A2(n18167), .ZN(n18552) );
  INV_X1 U21183 ( .A(n18552), .ZN(n18430) );
  NAND2_X1 U21184 ( .A1(BUF2_REG_26__SCAN_IN), .A2(n18539), .ZN(n18556) );
  INV_X1 U21185 ( .A(n18556), .ZN(n18427) );
  NOR2_X2 U21186 ( .A1(n18262), .A2(n18168), .ZN(n18551) );
  AOI22_X1 U21187 ( .A1(n18586), .A2(n18427), .B1(n18191), .B2(n18551), .ZN(
        n18171) );
  NOR2_X2 U21188 ( .A1(n18169), .A2(n18192), .ZN(n18553) );
  AOI22_X1 U21189 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18194), .B1(
        n18253), .B2(n18553), .ZN(n18170) );
  OAI211_X1 U21190 ( .C1(n18208), .C2(n18430), .A(n18171), .B(n18170), .ZN(
        P3_U2870) );
  NAND2_X1 U21191 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18539), .ZN(n18434) );
  INV_X1 U21192 ( .A(n18208), .ZN(n18528) );
  NAND2_X1 U21193 ( .A1(n18539), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18562) );
  INV_X1 U21194 ( .A(n18562), .ZN(n18431) );
  NOR2_X2 U21195 ( .A1(n18262), .A2(n18172), .ZN(n18557) );
  AOI22_X1 U21196 ( .A1(n18528), .A2(n18431), .B1(n18191), .B2(n18557), .ZN(
        n18175) );
  NOR2_X2 U21197 ( .A1(n18173), .A2(n18192), .ZN(n18559) );
  AOI22_X1 U21198 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18194), .B1(
        n18253), .B2(n18559), .ZN(n18174) );
  OAI211_X1 U21199 ( .C1(n18576), .C2(n18434), .A(n18175), .B(n18174), .ZN(
        P3_U2871) );
  NOR2_X1 U21200 ( .A1(n18176), .A2(n18264), .ZN(n18564) );
  INV_X1 U21201 ( .A(n18564), .ZN(n18519) );
  NAND2_X1 U21202 ( .A1(n18539), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18568) );
  INV_X1 U21203 ( .A(n18568), .ZN(n18516) );
  NOR2_X2 U21204 ( .A1(n18262), .A2(n18177), .ZN(n18563) );
  AOI22_X1 U21205 ( .A1(n18528), .A2(n18516), .B1(n18191), .B2(n18563), .ZN(
        n18180) );
  NOR2_X2 U21206 ( .A1(n18178), .A2(n18192), .ZN(n18565) );
  AOI22_X1 U21207 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18194), .B1(
        n18253), .B2(n18565), .ZN(n18179) );
  OAI211_X1 U21208 ( .C1(n18576), .C2(n18519), .A(n18180), .B(n18179), .ZN(
        P3_U2872) );
  NOR2_X1 U21209 ( .A1(n18264), .A2(n14259), .ZN(n18462) );
  INV_X1 U21210 ( .A(n18462), .ZN(n18575) );
  NAND2_X1 U21211 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n18539), .ZN(n18465) );
  INV_X1 U21212 ( .A(n18465), .ZN(n18570) );
  NOR2_X2 U21213 ( .A1(n18262), .A2(n18181), .ZN(n18571) );
  AOI22_X1 U21214 ( .A1(n18586), .A2(n18570), .B1(n18191), .B2(n18571), .ZN(
        n18184) );
  NOR2_X2 U21215 ( .A1(n18182), .A2(n18192), .ZN(n18572) );
  AOI22_X1 U21216 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18194), .B1(
        n18253), .B2(n18572), .ZN(n18183) );
  OAI211_X1 U21217 ( .C1(n18208), .C2(n18575), .A(n18184), .B(n18183), .ZN(
        P3_U2873) );
  NOR2_X1 U21218 ( .A1(n18264), .A2(n18185), .ZN(n18578) );
  NAND2_X1 U21219 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18539), .ZN(n18582) );
  NOR2_X2 U21220 ( .A1(n18262), .A2(n18186), .ZN(n18577) );
  AOI22_X1 U21221 ( .A1(n18586), .A2(n18493), .B1(n18191), .B2(n18577), .ZN(
        n18189) );
  NOR2_X2 U21222 ( .A1(n18187), .A2(n18192), .ZN(n18579) );
  AOI22_X1 U21223 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18194), .B1(
        n18253), .B2(n18579), .ZN(n18188) );
  OAI211_X1 U21224 ( .C1(n18208), .C2(n18496), .A(n18189), .B(n18188), .ZN(
        P3_U2874) );
  NOR2_X1 U21225 ( .A1(n15207), .A2(n18264), .ZN(n18585) );
  INV_X1 U21226 ( .A(n18585), .ZN(n18532) );
  NAND2_X1 U21227 ( .A1(n18539), .A2(BUF2_REG_31__SCAN_IN), .ZN(n18593) );
  INV_X1 U21228 ( .A(n18593), .ZN(n18527) );
  NOR2_X2 U21229 ( .A1(n18190), .A2(n18262), .ZN(n18584) );
  AOI22_X1 U21230 ( .A1(n18586), .A2(n18527), .B1(n18191), .B2(n18584), .ZN(
        n18196) );
  NOR2_X2 U21231 ( .A1(n18193), .A2(n18192), .ZN(n18587) );
  AOI22_X1 U21232 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18194), .B1(
        n18253), .B2(n18587), .ZN(n18195) );
  OAI211_X1 U21233 ( .C1(n18208), .C2(n18532), .A(n18196), .B(n18195), .ZN(
        P3_U2875) );
  NAND2_X1 U21234 ( .A1(n18240), .A2(n18374), .ZN(n18286) );
  INV_X1 U21235 ( .A(n18509), .ZN(n18535) );
  INV_X1 U21236 ( .A(n18544), .ZN(n18588) );
  INV_X1 U21237 ( .A(n18240), .ZN(n18237) );
  NAND2_X1 U21238 ( .A1(n18636), .A2(n18533), .ZN(n18375) );
  NOR2_X1 U21239 ( .A1(n18237), .A2(n18375), .ZN(n18213) );
  AOI22_X1 U21240 ( .A1(n18535), .A2(n18588), .B1(n18534), .B2(n18213), .ZN(
        n18199) );
  NOR2_X1 U21241 ( .A1(n18262), .A2(n18197), .ZN(n18536) );
  INV_X1 U21242 ( .A(n18536), .ZN(n18238) );
  NOR2_X1 U21243 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18238), .ZN(
        n18475) );
  AOI22_X1 U21244 ( .A1(n18539), .A2(n18537), .B1(n18240), .B2(n18475), .ZN(
        n18214) );
  AOI22_X1 U21245 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18214), .B1(
        n18528), .B2(n18540), .ZN(n18198) );
  OAI211_X1 U21246 ( .C1(n18543), .C2(n18286), .A(n18199), .B(n18198), .ZN(
        P3_U2876) );
  AOI22_X1 U21247 ( .A1(n18528), .A2(n18480), .B1(n18545), .B2(n18213), .ZN(
        n18201) );
  AOI22_X1 U21248 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18214), .B1(
        n18547), .B2(n18279), .ZN(n18200) );
  OAI211_X1 U21249 ( .C1(n18544), .C2(n18483), .A(n18201), .B(n18200), .ZN(
        P3_U2877) );
  AOI22_X1 U21250 ( .A1(n18528), .A2(n18427), .B1(n18551), .B2(n18213), .ZN(
        n18203) );
  AOI22_X1 U21251 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18214), .B1(
        n18553), .B2(n18279), .ZN(n18202) );
  OAI211_X1 U21252 ( .C1(n18544), .C2(n18430), .A(n18203), .B(n18202), .ZN(
        P3_U2878) );
  AOI22_X1 U21253 ( .A1(n18588), .A2(n18431), .B1(n18557), .B2(n18213), .ZN(
        n18205) );
  AOI22_X1 U21254 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18214), .B1(
        n18559), .B2(n18279), .ZN(n18204) );
  OAI211_X1 U21255 ( .C1(n18208), .C2(n18434), .A(n18205), .B(n18204), .ZN(
        P3_U2879) );
  AOI22_X1 U21256 ( .A1(n18588), .A2(n18516), .B1(n18563), .B2(n18213), .ZN(
        n18207) );
  AOI22_X1 U21257 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18214), .B1(
        n18565), .B2(n18279), .ZN(n18206) );
  OAI211_X1 U21258 ( .C1(n18208), .C2(n18519), .A(n18207), .B(n18206), .ZN(
        P3_U2880) );
  AOI22_X1 U21259 ( .A1(n18528), .A2(n18570), .B1(n18571), .B2(n18213), .ZN(
        n18210) );
  AOI22_X1 U21260 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18214), .B1(
        n18572), .B2(n18279), .ZN(n18209) );
  OAI211_X1 U21261 ( .C1(n18544), .C2(n18575), .A(n18210), .B(n18209), .ZN(
        P3_U2881) );
  AOI22_X1 U21262 ( .A1(n18528), .A2(n18493), .B1(n18577), .B2(n18213), .ZN(
        n18212) );
  AOI22_X1 U21263 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18214), .B1(
        n18579), .B2(n18279), .ZN(n18211) );
  OAI211_X1 U21264 ( .C1(n18544), .C2(n18496), .A(n18212), .B(n18211), .ZN(
        P3_U2882) );
  AOI22_X1 U21265 ( .A1(n18528), .A2(n18527), .B1(n18584), .B2(n18213), .ZN(
        n18216) );
  AOI22_X1 U21266 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18214), .B1(
        n18587), .B2(n18279), .ZN(n18215) );
  OAI211_X1 U21267 ( .C1(n18544), .C2(n18532), .A(n18216), .B(n18215), .ZN(
        P3_U2883) );
  NAND2_X1 U21268 ( .A1(n18398), .A2(n18240), .ZN(n18308) );
  NOR2_X1 U21269 ( .A1(n18279), .A2(n18301), .ZN(n18265) );
  NOR2_X1 U21270 ( .A1(n18662), .A2(n18265), .ZN(n18233) );
  AOI22_X1 U21271 ( .A1(n18535), .A2(n18253), .B1(n18534), .B2(n18233), .ZN(
        n18220) );
  INV_X1 U21272 ( .A(n18262), .ZN(n18451) );
  OAI21_X1 U21273 ( .B1(n18217), .B2(n18239), .A(n18265), .ZN(n18218) );
  OAI211_X1 U21274 ( .C1(n18301), .C2(n18763), .A(n18451), .B(n18218), .ZN(
        n18234) );
  AOI22_X1 U21275 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18234), .B1(
        n18588), .B2(n18540), .ZN(n18219) );
  OAI211_X1 U21276 ( .C1(n18543), .C2(n18308), .A(n18220), .B(n18219), .ZN(
        P3_U2884) );
  AOI22_X1 U21277 ( .A1(n18588), .A2(n18480), .B1(n18545), .B2(n18233), .ZN(
        n18222) );
  AOI22_X1 U21278 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18234), .B1(
        n18547), .B2(n18301), .ZN(n18221) );
  OAI211_X1 U21279 ( .C1(n18260), .C2(n18483), .A(n18222), .B(n18221), .ZN(
        P3_U2885) );
  AOI22_X1 U21280 ( .A1(n18253), .A2(n18552), .B1(n18551), .B2(n18233), .ZN(
        n18224) );
  AOI22_X1 U21281 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18234), .B1(
        n18553), .B2(n18301), .ZN(n18223) );
  OAI211_X1 U21282 ( .C1(n18544), .C2(n18556), .A(n18224), .B(n18223), .ZN(
        P3_U2886) );
  AOI22_X1 U21283 ( .A1(n18253), .A2(n18431), .B1(n18557), .B2(n18233), .ZN(
        n18226) );
  AOI22_X1 U21284 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18234), .B1(
        n18559), .B2(n18301), .ZN(n18225) );
  OAI211_X1 U21285 ( .C1(n18544), .C2(n18434), .A(n18226), .B(n18225), .ZN(
        P3_U2887) );
  AOI22_X1 U21286 ( .A1(n18588), .A2(n18564), .B1(n18563), .B2(n18233), .ZN(
        n18228) );
  AOI22_X1 U21287 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18234), .B1(
        n18565), .B2(n18301), .ZN(n18227) );
  OAI211_X1 U21288 ( .C1(n18260), .C2(n18568), .A(n18228), .B(n18227), .ZN(
        P3_U2888) );
  AOI22_X1 U21289 ( .A1(n18253), .A2(n18462), .B1(n18571), .B2(n18233), .ZN(
        n18230) );
  AOI22_X1 U21290 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18234), .B1(
        n18572), .B2(n18301), .ZN(n18229) );
  OAI211_X1 U21291 ( .C1(n18544), .C2(n18465), .A(n18230), .B(n18229), .ZN(
        P3_U2889) );
  AOI22_X1 U21292 ( .A1(n18588), .A2(n18493), .B1(n18577), .B2(n18233), .ZN(
        n18232) );
  AOI22_X1 U21293 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18234), .B1(
        n18579), .B2(n18301), .ZN(n18231) );
  OAI211_X1 U21294 ( .C1(n18260), .C2(n18496), .A(n18232), .B(n18231), .ZN(
        P3_U2890) );
  AOI22_X1 U21295 ( .A1(n18588), .A2(n18527), .B1(n18584), .B2(n18233), .ZN(
        n18236) );
  AOI22_X1 U21296 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18234), .B1(
        n18587), .B2(n18301), .ZN(n18235) );
  OAI211_X1 U21297 ( .C1(n18260), .C2(n18532), .A(n18236), .B(n18235), .ZN(
        P3_U2891) );
  NOR2_X1 U21298 ( .A1(n18636), .A2(n18237), .ZN(n18288) );
  AND2_X1 U21299 ( .A1(n18533), .A2(n18288), .ZN(n18256) );
  AOI22_X1 U21300 ( .A1(n18253), .A2(n18540), .B1(n18534), .B2(n18256), .ZN(
        n18242) );
  AOI21_X1 U21301 ( .B1(n18636), .B2(n18239), .A(n18238), .ZN(n18332) );
  NAND2_X1 U21302 ( .A1(n18240), .A2(n18332), .ZN(n18257) );
  NAND2_X1 U21303 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18288), .ZN(
        n18329) );
  AOI22_X1 U21304 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18257), .B1(
        n18506), .B2(n18322), .ZN(n18241) );
  OAI211_X1 U21305 ( .C1(n18509), .C2(n18286), .A(n18242), .B(n18241), .ZN(
        P3_U2892) );
  AOI22_X1 U21306 ( .A1(n18546), .A2(n18279), .B1(n18545), .B2(n18256), .ZN(
        n18244) );
  AOI22_X1 U21307 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18257), .B1(
        n18547), .B2(n18322), .ZN(n18243) );
  OAI211_X1 U21308 ( .C1(n18260), .C2(n18550), .A(n18244), .B(n18243), .ZN(
        P3_U2893) );
  AOI22_X1 U21309 ( .A1(n18253), .A2(n18427), .B1(n18551), .B2(n18256), .ZN(
        n18246) );
  AOI22_X1 U21310 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18257), .B1(
        n18553), .B2(n18322), .ZN(n18245) );
  OAI211_X1 U21311 ( .C1(n18430), .C2(n18286), .A(n18246), .B(n18245), .ZN(
        P3_U2894) );
  INV_X1 U21312 ( .A(n18434), .ZN(n18558) );
  AOI22_X1 U21313 ( .A1(n18253), .A2(n18558), .B1(n18557), .B2(n18256), .ZN(
        n18248) );
  AOI22_X1 U21314 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18257), .B1(
        n18559), .B2(n18322), .ZN(n18247) );
  OAI211_X1 U21315 ( .C1(n18562), .C2(n18286), .A(n18248), .B(n18247), .ZN(
        P3_U2895) );
  AOI22_X1 U21316 ( .A1(n18253), .A2(n18564), .B1(n18563), .B2(n18256), .ZN(
        n18250) );
  AOI22_X1 U21317 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18257), .B1(
        n18565), .B2(n18322), .ZN(n18249) );
  OAI211_X1 U21318 ( .C1(n18568), .C2(n18286), .A(n18250), .B(n18249), .ZN(
        P3_U2896) );
  AOI22_X1 U21319 ( .A1(n18462), .A2(n18279), .B1(n18571), .B2(n18256), .ZN(
        n18252) );
  AOI22_X1 U21320 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18257), .B1(
        n18572), .B2(n18322), .ZN(n18251) );
  OAI211_X1 U21321 ( .C1(n18260), .C2(n18465), .A(n18252), .B(n18251), .ZN(
        P3_U2897) );
  AOI22_X1 U21322 ( .A1(n18253), .A2(n18493), .B1(n18577), .B2(n18256), .ZN(
        n18255) );
  AOI22_X1 U21323 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18257), .B1(
        n18579), .B2(n18322), .ZN(n18254) );
  OAI211_X1 U21324 ( .C1(n18496), .C2(n18286), .A(n18255), .B(n18254), .ZN(
        P3_U2898) );
  AOI22_X1 U21325 ( .A1(n18585), .A2(n18279), .B1(n18584), .B2(n18256), .ZN(
        n18259) );
  AOI22_X1 U21326 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18257), .B1(
        n18587), .B2(n18322), .ZN(n18258) );
  OAI211_X1 U21327 ( .C1(n18260), .C2(n18593), .A(n18259), .B(n18258), .ZN(
        P3_U2899) );
  INV_X1 U21328 ( .A(n18261), .ZN(n18637) );
  NOR2_X2 U21329 ( .A1(n18637), .A2(n18287), .ZN(n18345) );
  INV_X1 U21330 ( .A(n18345), .ZN(n18352) );
  NAND2_X1 U21331 ( .A1(n18329), .A2(n18352), .ZN(n18309) );
  INV_X1 U21332 ( .A(n18309), .ZN(n18263) );
  NOR2_X1 U21333 ( .A1(n18662), .A2(n18263), .ZN(n18282) );
  AOI22_X1 U21334 ( .A1(n18535), .A2(n18301), .B1(n18534), .B2(n18282), .ZN(
        n18268) );
  OAI22_X1 U21335 ( .A1(n18265), .A2(n18264), .B1(n18263), .B2(n18262), .ZN(
        n18266) );
  OAI21_X1 U21336 ( .B1(n18345), .B2(n18763), .A(n18266), .ZN(n18283) );
  AOI22_X1 U21337 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18283), .B1(
        n18540), .B2(n18279), .ZN(n18267) );
  OAI211_X1 U21338 ( .C1(n18543), .C2(n18352), .A(n18268), .B(n18267), .ZN(
        P3_U2900) );
  AOI22_X1 U21339 ( .A1(n18546), .A2(n18301), .B1(n18545), .B2(n18282), .ZN(
        n18270) );
  AOI22_X1 U21340 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18283), .B1(
        n18547), .B2(n18345), .ZN(n18269) );
  OAI211_X1 U21341 ( .C1(n18550), .C2(n18286), .A(n18270), .B(n18269), .ZN(
        P3_U2901) );
  AOI22_X1 U21342 ( .A1(n18427), .A2(n18279), .B1(n18551), .B2(n18282), .ZN(
        n18272) );
  AOI22_X1 U21343 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18283), .B1(
        n18553), .B2(n18345), .ZN(n18271) );
  OAI211_X1 U21344 ( .C1(n18430), .C2(n18308), .A(n18272), .B(n18271), .ZN(
        P3_U2902) );
  AOI22_X1 U21345 ( .A1(n18431), .A2(n18301), .B1(n18557), .B2(n18282), .ZN(
        n18274) );
  AOI22_X1 U21346 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18283), .B1(
        n18559), .B2(n18345), .ZN(n18273) );
  OAI211_X1 U21347 ( .C1(n18434), .C2(n18286), .A(n18274), .B(n18273), .ZN(
        P3_U2903) );
  AOI22_X1 U21348 ( .A1(n18564), .A2(n18279), .B1(n18563), .B2(n18282), .ZN(
        n18276) );
  AOI22_X1 U21349 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18283), .B1(
        n18565), .B2(n18345), .ZN(n18275) );
  OAI211_X1 U21350 ( .C1(n18568), .C2(n18308), .A(n18276), .B(n18275), .ZN(
        P3_U2904) );
  AOI22_X1 U21351 ( .A1(n18462), .A2(n18301), .B1(n18571), .B2(n18282), .ZN(
        n18278) );
  AOI22_X1 U21352 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18283), .B1(
        n18572), .B2(n18345), .ZN(n18277) );
  OAI211_X1 U21353 ( .C1(n18465), .C2(n18286), .A(n18278), .B(n18277), .ZN(
        P3_U2905) );
  AOI22_X1 U21354 ( .A1(n18577), .A2(n18282), .B1(n18493), .B2(n18279), .ZN(
        n18281) );
  AOI22_X1 U21355 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18283), .B1(
        n18579), .B2(n18345), .ZN(n18280) );
  OAI211_X1 U21356 ( .C1(n18496), .C2(n18308), .A(n18281), .B(n18280), .ZN(
        P3_U2906) );
  AOI22_X1 U21357 ( .A1(n18585), .A2(n18301), .B1(n18584), .B2(n18282), .ZN(
        n18285) );
  AOI22_X1 U21358 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18283), .B1(
        n18587), .B2(n18345), .ZN(n18284) );
  OAI211_X1 U21359 ( .C1(n18593), .C2(n18286), .A(n18285), .B(n18284), .ZN(
        P3_U2907) );
  INV_X1 U21360 ( .A(n18287), .ZN(n18331) );
  NAND2_X1 U21361 ( .A1(n18374), .A2(n18331), .ZN(n18362) );
  NOR2_X1 U21362 ( .A1(n18375), .A2(n18287), .ZN(n18304) );
  AOI22_X1 U21363 ( .A1(n18540), .A2(n18301), .B1(n18534), .B2(n18304), .ZN(
        n18290) );
  AOI22_X1 U21364 ( .A1(n18539), .A2(n18288), .B1(n18475), .B2(n18331), .ZN(
        n18305) );
  AOI22_X1 U21365 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18305), .B1(
        n18535), .B2(n18322), .ZN(n18289) );
  OAI211_X1 U21366 ( .C1(n18543), .C2(n18362), .A(n18290), .B(n18289), .ZN(
        P3_U2908) );
  AOI22_X1 U21367 ( .A1(n18546), .A2(n18322), .B1(n18545), .B2(n18304), .ZN(
        n18292) );
  INV_X1 U21368 ( .A(n18362), .ZN(n18370) );
  AOI22_X1 U21369 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18305), .B1(
        n18547), .B2(n18370), .ZN(n18291) );
  OAI211_X1 U21370 ( .C1(n18550), .C2(n18308), .A(n18292), .B(n18291), .ZN(
        P3_U2909) );
  AOI22_X1 U21371 ( .A1(n18552), .A2(n18322), .B1(n18551), .B2(n18304), .ZN(
        n18294) );
  AOI22_X1 U21372 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18305), .B1(
        n18553), .B2(n18370), .ZN(n18293) );
  OAI211_X1 U21373 ( .C1(n18556), .C2(n18308), .A(n18294), .B(n18293), .ZN(
        P3_U2910) );
  AOI22_X1 U21374 ( .A1(n18558), .A2(n18301), .B1(n18557), .B2(n18304), .ZN(
        n18296) );
  AOI22_X1 U21375 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18305), .B1(
        n18559), .B2(n18370), .ZN(n18295) );
  OAI211_X1 U21376 ( .C1(n18562), .C2(n18329), .A(n18296), .B(n18295), .ZN(
        P3_U2911) );
  AOI22_X1 U21377 ( .A1(n18564), .A2(n18301), .B1(n18563), .B2(n18304), .ZN(
        n18298) );
  AOI22_X1 U21378 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18305), .B1(
        n18565), .B2(n18370), .ZN(n18297) );
  OAI211_X1 U21379 ( .C1(n18568), .C2(n18329), .A(n18298), .B(n18297), .ZN(
        P3_U2912) );
  AOI22_X1 U21380 ( .A1(n18462), .A2(n18322), .B1(n18571), .B2(n18304), .ZN(
        n18300) );
  AOI22_X1 U21381 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18305), .B1(
        n18572), .B2(n18370), .ZN(n18299) );
  OAI211_X1 U21382 ( .C1(n18465), .C2(n18308), .A(n18300), .B(n18299), .ZN(
        P3_U2913) );
  AOI22_X1 U21383 ( .A1(n18577), .A2(n18304), .B1(n18493), .B2(n18301), .ZN(
        n18303) );
  AOI22_X1 U21384 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18305), .B1(
        n18579), .B2(n18370), .ZN(n18302) );
  OAI211_X1 U21385 ( .C1(n18496), .C2(n18329), .A(n18303), .B(n18302), .ZN(
        P3_U2914) );
  AOI22_X1 U21386 ( .A1(n18585), .A2(n18322), .B1(n18584), .B2(n18304), .ZN(
        n18307) );
  AOI22_X1 U21387 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18305), .B1(
        n18587), .B2(n18370), .ZN(n18306) );
  OAI211_X1 U21388 ( .C1(n18593), .C2(n18308), .A(n18307), .B(n18306), .ZN(
        P3_U2915) );
  NAND2_X1 U21389 ( .A1(n18398), .A2(n18331), .ZN(n18396) );
  NAND2_X1 U21390 ( .A1(n18362), .A2(n18396), .ZN(n18353) );
  AND2_X1 U21391 ( .A1(n18533), .A2(n18353), .ZN(n18325) );
  AOI22_X1 U21392 ( .A1(n18535), .A2(n18345), .B1(n18534), .B2(n18325), .ZN(
        n18311) );
  OAI221_X1 U21393 ( .B1(n18353), .B2(n18504), .C1(n18353), .C2(n18309), .A(
        n18502), .ZN(n18326) );
  AOI22_X1 U21394 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18326), .B1(
        n18540), .B2(n18322), .ZN(n18310) );
  OAI211_X1 U21395 ( .C1(n18543), .C2(n18396), .A(n18311), .B(n18310), .ZN(
        P3_U2916) );
  AOI22_X1 U21396 ( .A1(n18480), .A2(n18322), .B1(n18545), .B2(n18325), .ZN(
        n18313) );
  INV_X1 U21397 ( .A(n18396), .ZN(n18387) );
  AOI22_X1 U21398 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18326), .B1(
        n18547), .B2(n18387), .ZN(n18312) );
  OAI211_X1 U21399 ( .C1(n18483), .C2(n18352), .A(n18313), .B(n18312), .ZN(
        P3_U2917) );
  AOI22_X1 U21400 ( .A1(n18552), .A2(n18345), .B1(n18551), .B2(n18325), .ZN(
        n18315) );
  AOI22_X1 U21401 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18326), .B1(
        n18553), .B2(n18387), .ZN(n18314) );
  OAI211_X1 U21402 ( .C1(n18556), .C2(n18329), .A(n18315), .B(n18314), .ZN(
        P3_U2918) );
  AOI22_X1 U21403 ( .A1(n18431), .A2(n18345), .B1(n18557), .B2(n18325), .ZN(
        n18317) );
  AOI22_X1 U21404 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18326), .B1(
        n18559), .B2(n18387), .ZN(n18316) );
  OAI211_X1 U21405 ( .C1(n18434), .C2(n18329), .A(n18317), .B(n18316), .ZN(
        P3_U2919) );
  AOI22_X1 U21406 ( .A1(n18516), .A2(n18345), .B1(n18563), .B2(n18325), .ZN(
        n18319) );
  AOI22_X1 U21407 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18326), .B1(
        n18565), .B2(n18387), .ZN(n18318) );
  OAI211_X1 U21408 ( .C1(n18519), .C2(n18329), .A(n18319), .B(n18318), .ZN(
        P3_U2920) );
  AOI22_X1 U21409 ( .A1(n18462), .A2(n18345), .B1(n18571), .B2(n18325), .ZN(
        n18321) );
  AOI22_X1 U21410 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18326), .B1(
        n18572), .B2(n18387), .ZN(n18320) );
  OAI211_X1 U21411 ( .C1(n18465), .C2(n18329), .A(n18321), .B(n18320), .ZN(
        P3_U2921) );
  AOI22_X1 U21412 ( .A1(n18577), .A2(n18325), .B1(n18493), .B2(n18322), .ZN(
        n18324) );
  AOI22_X1 U21413 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18326), .B1(
        n18579), .B2(n18387), .ZN(n18323) );
  OAI211_X1 U21414 ( .C1(n18496), .C2(n18352), .A(n18324), .B(n18323), .ZN(
        P3_U2922) );
  AOI22_X1 U21415 ( .A1(n18585), .A2(n18345), .B1(n18584), .B2(n18325), .ZN(
        n18328) );
  AOI22_X1 U21416 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18326), .B1(
        n18587), .B2(n18387), .ZN(n18327) );
  OAI211_X1 U21417 ( .C1(n18593), .C2(n18329), .A(n18328), .B(n18327), .ZN(
        P3_U2923) );
  INV_X1 U21418 ( .A(n9716), .ZN(n18420) );
  NOR2_X1 U21419 ( .A1(n18330), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18376) );
  AND2_X1 U21420 ( .A1(n18533), .A2(n18376), .ZN(n18348) );
  AOI22_X1 U21421 ( .A1(n18535), .A2(n18370), .B1(n18534), .B2(n18348), .ZN(
        n18334) );
  NAND2_X1 U21422 ( .A1(n18332), .A2(n18331), .ZN(n18349) );
  AOI22_X1 U21423 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18349), .B1(
        n18540), .B2(n18345), .ZN(n18333) );
  OAI211_X1 U21424 ( .C1(n18543), .C2(n18420), .A(n18334), .B(n18333), .ZN(
        P3_U2924) );
  AOI22_X1 U21425 ( .A1(n18546), .A2(n18370), .B1(n18545), .B2(n18348), .ZN(
        n18336) );
  AOI22_X1 U21426 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18349), .B1(
        n18547), .B2(n9716), .ZN(n18335) );
  OAI211_X1 U21427 ( .C1(n18550), .C2(n18352), .A(n18336), .B(n18335), .ZN(
        P3_U2925) );
  AOI22_X1 U21428 ( .A1(n18427), .A2(n18345), .B1(n18551), .B2(n18348), .ZN(
        n18338) );
  AOI22_X1 U21429 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18349), .B1(
        n18553), .B2(n9716), .ZN(n18337) );
  OAI211_X1 U21430 ( .C1(n18430), .C2(n18362), .A(n18338), .B(n18337), .ZN(
        P3_U2926) );
  AOI22_X1 U21431 ( .A1(n18558), .A2(n18345), .B1(n18557), .B2(n18348), .ZN(
        n18340) );
  AOI22_X1 U21432 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18349), .B1(
        n18559), .B2(n9716), .ZN(n18339) );
  OAI211_X1 U21433 ( .C1(n18562), .C2(n18362), .A(n18340), .B(n18339), .ZN(
        P3_U2927) );
  AOI22_X1 U21434 ( .A1(n18516), .A2(n18370), .B1(n18563), .B2(n18348), .ZN(
        n18342) );
  AOI22_X1 U21435 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18349), .B1(
        n18565), .B2(n9716), .ZN(n18341) );
  OAI211_X1 U21436 ( .C1(n18519), .C2(n18352), .A(n18342), .B(n18341), .ZN(
        P3_U2928) );
  AOI22_X1 U21437 ( .A1(n18571), .A2(n18348), .B1(n18570), .B2(n18345), .ZN(
        n18344) );
  AOI22_X1 U21438 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18349), .B1(
        n18572), .B2(n9716), .ZN(n18343) );
  OAI211_X1 U21439 ( .C1(n18575), .C2(n18362), .A(n18344), .B(n18343), .ZN(
        P3_U2929) );
  AOI22_X1 U21440 ( .A1(n18577), .A2(n18348), .B1(n18493), .B2(n18345), .ZN(
        n18347) );
  AOI22_X1 U21441 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18349), .B1(
        n18579), .B2(n9716), .ZN(n18346) );
  OAI211_X1 U21442 ( .C1(n18496), .C2(n18362), .A(n18347), .B(n18346), .ZN(
        P3_U2930) );
  AOI22_X1 U21443 ( .A1(n18585), .A2(n18370), .B1(n18584), .B2(n18348), .ZN(
        n18351) );
  AOI22_X1 U21444 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18349), .B1(
        n18587), .B2(n9716), .ZN(n18350) );
  OAI211_X1 U21445 ( .C1(n18593), .C2(n18352), .A(n18351), .B(n18350), .ZN(
        P3_U2931) );
  NOR2_X2 U21446 ( .A1(n18637), .A2(n18421), .ZN(n18437) );
  INV_X1 U21447 ( .A(n18437), .ZN(n18446) );
  NAND2_X1 U21448 ( .A1(n18420), .A2(n18446), .ZN(n18399) );
  AND2_X1 U21449 ( .A1(n18533), .A2(n18399), .ZN(n18369) );
  AOI22_X1 U21450 ( .A1(n18535), .A2(n18387), .B1(n18534), .B2(n18369), .ZN(
        n18355) );
  OAI221_X1 U21451 ( .B1(n18399), .B2(n18504), .C1(n18399), .C2(n18353), .A(
        n18502), .ZN(n18371) );
  AOI22_X1 U21452 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18371), .B1(
        n18540), .B2(n18370), .ZN(n18354) );
  OAI211_X1 U21453 ( .C1(n18543), .C2(n18446), .A(n18355), .B(n18354), .ZN(
        P3_U2932) );
  AOI22_X1 U21454 ( .A1(n18546), .A2(n18387), .B1(n18545), .B2(n18369), .ZN(
        n18357) );
  AOI22_X1 U21455 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18371), .B1(
        n18547), .B2(n18437), .ZN(n18356) );
  OAI211_X1 U21456 ( .C1(n18550), .C2(n18362), .A(n18357), .B(n18356), .ZN(
        P3_U2933) );
  AOI22_X1 U21457 ( .A1(n18427), .A2(n18370), .B1(n18551), .B2(n18369), .ZN(
        n18359) );
  AOI22_X1 U21458 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18371), .B1(
        n18553), .B2(n18437), .ZN(n18358) );
  OAI211_X1 U21459 ( .C1(n18430), .C2(n18396), .A(n18359), .B(n18358), .ZN(
        P3_U2934) );
  AOI22_X1 U21460 ( .A1(n18431), .A2(n18387), .B1(n18557), .B2(n18369), .ZN(
        n18361) );
  AOI22_X1 U21461 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18371), .B1(
        n18559), .B2(n18437), .ZN(n18360) );
  OAI211_X1 U21462 ( .C1(n18434), .C2(n18362), .A(n18361), .B(n18360), .ZN(
        P3_U2935) );
  AOI22_X1 U21463 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18371), .B1(
        n18563), .B2(n18369), .ZN(n18364) );
  AOI22_X1 U21464 ( .A1(n18564), .A2(n18370), .B1(n18565), .B2(n18437), .ZN(
        n18363) );
  OAI211_X1 U21465 ( .C1(n18568), .C2(n18396), .A(n18364), .B(n18363), .ZN(
        P3_U2936) );
  AOI22_X1 U21466 ( .A1(n18571), .A2(n18369), .B1(n18570), .B2(n18370), .ZN(
        n18366) );
  AOI22_X1 U21467 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18371), .B1(
        n18572), .B2(n18437), .ZN(n18365) );
  OAI211_X1 U21468 ( .C1(n18575), .C2(n18396), .A(n18366), .B(n18365), .ZN(
        P3_U2937) );
  AOI22_X1 U21469 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18371), .B1(
        n18577), .B2(n18369), .ZN(n18368) );
  AOI22_X1 U21470 ( .A1(n18579), .A2(n18437), .B1(n18493), .B2(n18370), .ZN(
        n18367) );
  OAI211_X1 U21471 ( .C1(n18496), .C2(n18396), .A(n18368), .B(n18367), .ZN(
        P3_U2938) );
  AOI22_X1 U21472 ( .A1(n18527), .A2(n18370), .B1(n18584), .B2(n18369), .ZN(
        n18373) );
  AOI22_X1 U21473 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18371), .B1(
        n18587), .B2(n18437), .ZN(n18372) );
  OAI211_X1 U21474 ( .C1(n18532), .C2(n18396), .A(n18373), .B(n18372), .ZN(
        P3_U2939) );
  NAND2_X1 U21475 ( .A1(n18374), .A2(n18397), .ZN(n18468) );
  NOR2_X1 U21476 ( .A1(n18375), .A2(n18421), .ZN(n18392) );
  AOI22_X1 U21477 ( .A1(n18540), .A2(n18387), .B1(n18534), .B2(n18392), .ZN(
        n18378) );
  NOR2_X1 U21478 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18421), .ZN(
        n18422) );
  AOI22_X1 U21479 ( .A1(n18539), .A2(n18376), .B1(n18536), .B2(n18422), .ZN(
        n18393) );
  AOI22_X1 U21480 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18393), .B1(
        n18535), .B2(n9716), .ZN(n18377) );
  OAI211_X1 U21481 ( .C1(n18543), .C2(n18468), .A(n18378), .B(n18377), .ZN(
        P3_U2940) );
  AOI22_X1 U21482 ( .A1(n18480), .A2(n18387), .B1(n18545), .B2(n18392), .ZN(
        n18380) );
  INV_X1 U21483 ( .A(n18468), .ZN(n18470) );
  AOI22_X1 U21484 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18393), .B1(
        n18547), .B2(n18470), .ZN(n18379) );
  OAI211_X1 U21485 ( .C1(n18483), .C2(n18420), .A(n18380), .B(n18379), .ZN(
        P3_U2941) );
  AOI22_X1 U21486 ( .A1(n18427), .A2(n18387), .B1(n18551), .B2(n18392), .ZN(
        n18382) );
  AOI22_X1 U21487 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18393), .B1(
        n18553), .B2(n18470), .ZN(n18381) );
  OAI211_X1 U21488 ( .C1(n18430), .C2(n18420), .A(n18382), .B(n18381), .ZN(
        P3_U2942) );
  AOI22_X1 U21489 ( .A1(n18558), .A2(n18387), .B1(n18557), .B2(n18392), .ZN(
        n18384) );
  AOI22_X1 U21490 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18393), .B1(
        n18559), .B2(n18470), .ZN(n18383) );
  OAI211_X1 U21491 ( .C1(n18562), .C2(n18420), .A(n18384), .B(n18383), .ZN(
        P3_U2943) );
  AOI22_X1 U21492 ( .A1(n18564), .A2(n18387), .B1(n18563), .B2(n18392), .ZN(
        n18386) );
  AOI22_X1 U21493 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18393), .B1(
        n18565), .B2(n18470), .ZN(n18385) );
  OAI211_X1 U21494 ( .C1(n18568), .C2(n18420), .A(n18386), .B(n18385), .ZN(
        P3_U2944) );
  AOI22_X1 U21495 ( .A1(n18571), .A2(n18392), .B1(n18570), .B2(n18387), .ZN(
        n18389) );
  AOI22_X1 U21496 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18393), .B1(
        n18572), .B2(n18470), .ZN(n18388) );
  OAI211_X1 U21497 ( .C1(n18575), .C2(n18420), .A(n18389), .B(n18388), .ZN(
        P3_U2945) );
  AOI22_X1 U21498 ( .A1(n18578), .A2(n9716), .B1(n18577), .B2(n18392), .ZN(
        n18391) );
  AOI22_X1 U21499 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18393), .B1(
        n18579), .B2(n18470), .ZN(n18390) );
  OAI211_X1 U21500 ( .C1(n18582), .C2(n18396), .A(n18391), .B(n18390), .ZN(
        P3_U2946) );
  AOI22_X1 U21501 ( .A1(n18585), .A2(n9716), .B1(n18584), .B2(n18392), .ZN(
        n18395) );
  AOI22_X1 U21502 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18393), .B1(
        n18587), .B2(n18470), .ZN(n18394) );
  OAI211_X1 U21503 ( .C1(n18593), .C2(n18396), .A(n18395), .B(n18394), .ZN(
        P3_U2947) );
  NAND2_X1 U21504 ( .A1(n18398), .A2(n18397), .ZN(n18501) );
  AOI21_X1 U21505 ( .B1(n18468), .B2(n18501), .A(n18662), .ZN(n18416) );
  AOI22_X1 U21506 ( .A1(n18540), .A2(n9716), .B1(n18534), .B2(n18416), .ZN(
        n18402) );
  NAND2_X1 U21507 ( .A1(n18468), .A2(n18501), .ZN(n18400) );
  OAI221_X1 U21508 ( .B1(n18400), .B2(n18504), .C1(n18400), .C2(n18399), .A(
        n18502), .ZN(n18417) );
  AOI22_X1 U21509 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18417), .B1(
        n18535), .B2(n18437), .ZN(n18401) );
  OAI211_X1 U21510 ( .C1(n18543), .C2(n18501), .A(n18402), .B(n18401), .ZN(
        P3_U2948) );
  AOI22_X1 U21511 ( .A1(n18546), .A2(n18437), .B1(n18545), .B2(n18416), .ZN(
        n18404) );
  INV_X1 U21512 ( .A(n18501), .ZN(n18492) );
  AOI22_X1 U21513 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18417), .B1(
        n18547), .B2(n18492), .ZN(n18403) );
  OAI211_X1 U21514 ( .C1(n18550), .C2(n18420), .A(n18404), .B(n18403), .ZN(
        P3_U2949) );
  AOI22_X1 U21515 ( .A1(n18552), .A2(n18437), .B1(n18551), .B2(n18416), .ZN(
        n18406) );
  AOI22_X1 U21516 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18417), .B1(
        n18553), .B2(n18492), .ZN(n18405) );
  OAI211_X1 U21517 ( .C1(n18556), .C2(n18420), .A(n18406), .B(n18405), .ZN(
        P3_U2950) );
  AOI22_X1 U21518 ( .A1(n18431), .A2(n18437), .B1(n18557), .B2(n18416), .ZN(
        n18408) );
  AOI22_X1 U21519 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18417), .B1(
        n18559), .B2(n18492), .ZN(n18407) );
  OAI211_X1 U21520 ( .C1(n18434), .C2(n18420), .A(n18408), .B(n18407), .ZN(
        P3_U2951) );
  AOI22_X1 U21521 ( .A1(n18564), .A2(n9716), .B1(n18563), .B2(n18416), .ZN(
        n18410) );
  AOI22_X1 U21522 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18417), .B1(
        n18565), .B2(n18492), .ZN(n18409) );
  OAI211_X1 U21523 ( .C1(n18568), .C2(n18446), .A(n18410), .B(n18409), .ZN(
        P3_U2952) );
  AOI22_X1 U21524 ( .A1(n18462), .A2(n18437), .B1(n18571), .B2(n18416), .ZN(
        n18412) );
  AOI22_X1 U21525 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18417), .B1(
        n18572), .B2(n18492), .ZN(n18411) );
  OAI211_X1 U21526 ( .C1(n18465), .C2(n18420), .A(n18412), .B(n18411), .ZN(
        P3_U2953) );
  AOI22_X1 U21527 ( .A1(n18577), .A2(n18416), .B1(n18493), .B2(n9716), .ZN(
        n18415) );
  AOI22_X1 U21528 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18417), .B1(
        n18579), .B2(n18492), .ZN(n18414) );
  OAI211_X1 U21529 ( .C1(n18496), .C2(n18446), .A(n18415), .B(n18414), .ZN(
        P3_U2954) );
  AOI22_X1 U21530 ( .A1(n18585), .A2(n18437), .B1(n18584), .B2(n18416), .ZN(
        n18419) );
  AOI22_X1 U21531 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18417), .B1(
        n18587), .B2(n18492), .ZN(n18418) );
  OAI211_X1 U21532 ( .C1(n18593), .C2(n18420), .A(n18419), .B(n18418), .ZN(
        P3_U2955) );
  NOR2_X1 U21533 ( .A1(n18636), .A2(n18421), .ZN(n18477) );
  NAND2_X1 U21534 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18477), .ZN(
        n18524) );
  AND2_X1 U21535 ( .A1(n18533), .A2(n18477), .ZN(n18442) );
  AOI22_X1 U21536 ( .A1(n18535), .A2(n18470), .B1(n18534), .B2(n18442), .ZN(
        n18424) );
  AOI22_X1 U21537 ( .A1(n18539), .A2(n18422), .B1(n18536), .B2(n18477), .ZN(
        n18443) );
  AOI22_X1 U21538 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18443), .B1(
        n18540), .B2(n18437), .ZN(n18423) );
  OAI211_X1 U21539 ( .C1(n18543), .C2(n18524), .A(n18424), .B(n18423), .ZN(
        P3_U2956) );
  AOI22_X1 U21540 ( .A1(n18546), .A2(n18470), .B1(n18545), .B2(n18442), .ZN(
        n18426) );
  INV_X1 U21541 ( .A(n18524), .ZN(n18526) );
  AOI22_X1 U21542 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18443), .B1(
        n18547), .B2(n18526), .ZN(n18425) );
  OAI211_X1 U21543 ( .C1(n18550), .C2(n18446), .A(n18426), .B(n18425), .ZN(
        P3_U2957) );
  AOI22_X1 U21544 ( .A1(n18427), .A2(n18437), .B1(n18551), .B2(n18442), .ZN(
        n18429) );
  AOI22_X1 U21545 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18443), .B1(
        n18553), .B2(n18526), .ZN(n18428) );
  OAI211_X1 U21546 ( .C1(n18430), .C2(n18468), .A(n18429), .B(n18428), .ZN(
        P3_U2958) );
  AOI22_X1 U21547 ( .A1(n18431), .A2(n18470), .B1(n18557), .B2(n18442), .ZN(
        n18433) );
  AOI22_X1 U21548 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18443), .B1(
        n18559), .B2(n18526), .ZN(n18432) );
  OAI211_X1 U21549 ( .C1(n18434), .C2(n18446), .A(n18433), .B(n18432), .ZN(
        P3_U2959) );
  AOI22_X1 U21550 ( .A1(n18564), .A2(n18437), .B1(n18563), .B2(n18442), .ZN(
        n18436) );
  AOI22_X1 U21551 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18443), .B1(
        n18565), .B2(n18526), .ZN(n18435) );
  OAI211_X1 U21552 ( .C1(n18568), .C2(n18468), .A(n18436), .B(n18435), .ZN(
        P3_U2960) );
  AOI22_X1 U21553 ( .A1(n18571), .A2(n18442), .B1(n18570), .B2(n18437), .ZN(
        n18439) );
  AOI22_X1 U21554 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18443), .B1(
        n18572), .B2(n18526), .ZN(n18438) );
  OAI211_X1 U21555 ( .C1(n18575), .C2(n18468), .A(n18439), .B(n18438), .ZN(
        P3_U2961) );
  AOI22_X1 U21556 ( .A1(n18578), .A2(n18470), .B1(n18577), .B2(n18442), .ZN(
        n18441) );
  AOI22_X1 U21557 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18443), .B1(
        n18579), .B2(n18526), .ZN(n18440) );
  OAI211_X1 U21558 ( .C1(n18582), .C2(n18446), .A(n18441), .B(n18440), .ZN(
        P3_U2962) );
  AOI22_X1 U21559 ( .A1(n18585), .A2(n18470), .B1(n18584), .B2(n18442), .ZN(
        n18445) );
  AOI22_X1 U21560 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18443), .B1(
        n18587), .B2(n18526), .ZN(n18444) );
  OAI211_X1 U21561 ( .C1(n18593), .C2(n18446), .A(n18445), .B(n18444), .ZN(
        P3_U2963) );
  INV_X1 U21562 ( .A(n18538), .ZN(n18474) );
  NOR2_X2 U21563 ( .A1(n18474), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18569) );
  INV_X1 U21564 ( .A(n18569), .ZN(n18592) );
  NAND2_X1 U21565 ( .A1(n18524), .A2(n18592), .ZN(n18503) );
  INV_X1 U21566 ( .A(n18503), .ZN(n18447) );
  NOR2_X1 U21567 ( .A1(n18662), .A2(n18447), .ZN(n18469) );
  AOI22_X1 U21568 ( .A1(n18535), .A2(n18492), .B1(n18534), .B2(n18469), .ZN(
        n18453) );
  OAI21_X1 U21569 ( .B1(n18449), .B2(n18448), .A(n18447), .ZN(n18450) );
  OAI211_X1 U21570 ( .C1(n18569), .C2(n18763), .A(n18451), .B(n18450), .ZN(
        n18471) );
  AOI22_X1 U21571 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18471), .B1(
        n18540), .B2(n18470), .ZN(n18452) );
  OAI211_X1 U21572 ( .C1(n18543), .C2(n18592), .A(n18453), .B(n18452), .ZN(
        P3_U2964) );
  AOI22_X1 U21573 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18471), .B1(
        n18545), .B2(n18469), .ZN(n18455) );
  AOI22_X1 U21574 ( .A1(n18547), .A2(n18569), .B1(n18480), .B2(n18470), .ZN(
        n18454) );
  OAI211_X1 U21575 ( .C1(n18483), .C2(n18501), .A(n18455), .B(n18454), .ZN(
        P3_U2965) );
  AOI22_X1 U21576 ( .A1(n18552), .A2(n18492), .B1(n18551), .B2(n18469), .ZN(
        n18457) );
  AOI22_X1 U21577 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18471), .B1(
        n18553), .B2(n18569), .ZN(n18456) );
  OAI211_X1 U21578 ( .C1(n18556), .C2(n18468), .A(n18457), .B(n18456), .ZN(
        P3_U2966) );
  AOI22_X1 U21579 ( .A1(n18558), .A2(n18470), .B1(n18557), .B2(n18469), .ZN(
        n18459) );
  AOI22_X1 U21580 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18471), .B1(
        n18559), .B2(n18569), .ZN(n18458) );
  OAI211_X1 U21581 ( .C1(n18562), .C2(n18501), .A(n18459), .B(n18458), .ZN(
        P3_U2967) );
  AOI22_X1 U21582 ( .A1(n18516), .A2(n18492), .B1(n18563), .B2(n18469), .ZN(
        n18461) );
  AOI22_X1 U21583 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18471), .B1(
        n18565), .B2(n18569), .ZN(n18460) );
  OAI211_X1 U21584 ( .C1(n18519), .C2(n18468), .A(n18461), .B(n18460), .ZN(
        P3_U2968) );
  AOI22_X1 U21585 ( .A1(n18462), .A2(n18492), .B1(n18571), .B2(n18469), .ZN(
        n18464) );
  AOI22_X1 U21586 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18471), .B1(
        n18572), .B2(n18569), .ZN(n18463) );
  OAI211_X1 U21587 ( .C1(n18465), .C2(n18468), .A(n18464), .B(n18463), .ZN(
        P3_U2969) );
  AOI22_X1 U21588 ( .A1(n18578), .A2(n18492), .B1(n18577), .B2(n18469), .ZN(
        n18467) );
  AOI22_X1 U21589 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18471), .B1(
        n18579), .B2(n18569), .ZN(n18466) );
  OAI211_X1 U21590 ( .C1(n18582), .C2(n18468), .A(n18467), .B(n18466), .ZN(
        P3_U2970) );
  AOI22_X1 U21591 ( .A1(n18527), .A2(n18470), .B1(n18584), .B2(n18469), .ZN(
        n18473) );
  AOI22_X1 U21592 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18471), .B1(
        n18587), .B2(n18569), .ZN(n18472) );
  OAI211_X1 U21593 ( .C1(n18532), .C2(n18501), .A(n18473), .B(n18472), .ZN(
        P3_U2971) );
  NOR2_X1 U21594 ( .A1(n18662), .A2(n18474), .ZN(n18497) );
  AOI22_X1 U21595 ( .A1(n18540), .A2(n18492), .B1(n18534), .B2(n18497), .ZN(
        n18479) );
  AOI22_X1 U21596 ( .A1(n18539), .A2(n18477), .B1(n18476), .B2(n18475), .ZN(
        n18498) );
  AOI22_X1 U21597 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18498), .B1(
        n18506), .B2(n18586), .ZN(n18478) );
  OAI211_X1 U21598 ( .C1(n18509), .C2(n18524), .A(n18479), .B(n18478), .ZN(
        P3_U2972) );
  AOI22_X1 U21599 ( .A1(n18480), .A2(n18492), .B1(n18545), .B2(n18497), .ZN(
        n18482) );
  AOI22_X1 U21600 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18498), .B1(
        n18586), .B2(n18547), .ZN(n18481) );
  OAI211_X1 U21601 ( .C1(n18483), .C2(n18524), .A(n18482), .B(n18481), .ZN(
        P3_U2973) );
  AOI22_X1 U21602 ( .A1(n18552), .A2(n18526), .B1(n18551), .B2(n18497), .ZN(
        n18485) );
  AOI22_X1 U21603 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18498), .B1(
        n18586), .B2(n18553), .ZN(n18484) );
  OAI211_X1 U21604 ( .C1(n18556), .C2(n18501), .A(n18485), .B(n18484), .ZN(
        P3_U2974) );
  AOI22_X1 U21605 ( .A1(n18558), .A2(n18492), .B1(n18557), .B2(n18497), .ZN(
        n18487) );
  AOI22_X1 U21606 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18498), .B1(
        n18586), .B2(n18559), .ZN(n18486) );
  OAI211_X1 U21607 ( .C1(n18562), .C2(n18524), .A(n18487), .B(n18486), .ZN(
        P3_U2975) );
  AOI22_X1 U21608 ( .A1(n18516), .A2(n18526), .B1(n18563), .B2(n18497), .ZN(
        n18489) );
  AOI22_X1 U21609 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18498), .B1(
        n18586), .B2(n18565), .ZN(n18488) );
  OAI211_X1 U21610 ( .C1(n18519), .C2(n18501), .A(n18489), .B(n18488), .ZN(
        P3_U2976) );
  AOI22_X1 U21611 ( .A1(n18571), .A2(n18497), .B1(n18570), .B2(n18492), .ZN(
        n18491) );
  AOI22_X1 U21612 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18498), .B1(
        n18586), .B2(n18572), .ZN(n18490) );
  OAI211_X1 U21613 ( .C1(n18575), .C2(n18524), .A(n18491), .B(n18490), .ZN(
        P3_U2977) );
  AOI22_X1 U21614 ( .A1(n18577), .A2(n18497), .B1(n18493), .B2(n18492), .ZN(
        n18495) );
  AOI22_X1 U21615 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18498), .B1(
        n18586), .B2(n18579), .ZN(n18494) );
  OAI211_X1 U21616 ( .C1(n18496), .C2(n18524), .A(n18495), .B(n18494), .ZN(
        P3_U2978) );
  AOI22_X1 U21617 ( .A1(n18585), .A2(n18526), .B1(n18584), .B2(n18497), .ZN(
        n18500) );
  AOI22_X1 U21618 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18498), .B1(
        n18586), .B2(n18587), .ZN(n18499) );
  OAI211_X1 U21619 ( .C1(n18593), .C2(n18501), .A(n18500), .B(n18499), .ZN(
        P3_U2979) );
  AND2_X1 U21620 ( .A1(n18533), .A2(n18505), .ZN(n18525) );
  AOI22_X1 U21621 ( .A1(n18540), .A2(n18526), .B1(n18534), .B2(n18525), .ZN(
        n18508) );
  OAI221_X1 U21622 ( .B1(n18505), .B2(n18504), .C1(n18505), .C2(n18503), .A(
        n18502), .ZN(n18529) );
  AOI22_X1 U21623 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18529), .B1(
        n18528), .B2(n18506), .ZN(n18507) );
  OAI211_X1 U21624 ( .C1(n18509), .C2(n18592), .A(n18508), .B(n18507), .ZN(
        P3_U2980) );
  AOI22_X1 U21625 ( .A1(n18546), .A2(n18569), .B1(n18545), .B2(n18525), .ZN(
        n18511) );
  AOI22_X1 U21626 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18529), .B1(
        n18528), .B2(n18547), .ZN(n18510) );
  OAI211_X1 U21627 ( .C1(n18550), .C2(n18524), .A(n18511), .B(n18510), .ZN(
        P3_U2981) );
  AOI22_X1 U21628 ( .A1(n18552), .A2(n18569), .B1(n18551), .B2(n18525), .ZN(
        n18513) );
  AOI22_X1 U21629 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18529), .B1(
        n18528), .B2(n18553), .ZN(n18512) );
  OAI211_X1 U21630 ( .C1(n18556), .C2(n18524), .A(n18513), .B(n18512), .ZN(
        P3_U2982) );
  AOI22_X1 U21631 ( .A1(n18558), .A2(n18526), .B1(n18557), .B2(n18525), .ZN(
        n18515) );
  AOI22_X1 U21632 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18529), .B1(
        n18528), .B2(n18559), .ZN(n18514) );
  OAI211_X1 U21633 ( .C1(n18562), .C2(n18592), .A(n18515), .B(n18514), .ZN(
        P3_U2983) );
  AOI22_X1 U21634 ( .A1(n18516), .A2(n18569), .B1(n18563), .B2(n18525), .ZN(
        n18518) );
  AOI22_X1 U21635 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18529), .B1(
        n18528), .B2(n18565), .ZN(n18517) );
  OAI211_X1 U21636 ( .C1(n18519), .C2(n18524), .A(n18518), .B(n18517), .ZN(
        P3_U2984) );
  AOI22_X1 U21637 ( .A1(n18571), .A2(n18525), .B1(n18570), .B2(n18526), .ZN(
        n18521) );
  AOI22_X1 U21638 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18529), .B1(
        n18528), .B2(n18572), .ZN(n18520) );
  OAI211_X1 U21639 ( .C1(n18575), .C2(n18592), .A(n18521), .B(n18520), .ZN(
        P3_U2985) );
  AOI22_X1 U21640 ( .A1(n18578), .A2(n18569), .B1(n18577), .B2(n18525), .ZN(
        n18523) );
  AOI22_X1 U21641 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18529), .B1(
        n18528), .B2(n18579), .ZN(n18522) );
  OAI211_X1 U21642 ( .C1(n18582), .C2(n18524), .A(n18523), .B(n18522), .ZN(
        P3_U2986) );
  AOI22_X1 U21643 ( .A1(n18527), .A2(n18526), .B1(n18584), .B2(n18525), .ZN(
        n18531) );
  AOI22_X1 U21644 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18529), .B1(
        n18528), .B2(n18587), .ZN(n18530) );
  OAI211_X1 U21645 ( .C1(n18532), .C2(n18592), .A(n18531), .B(n18530), .ZN(
        P3_U2987) );
  AND2_X1 U21646 ( .A1(n18533), .A2(n18537), .ZN(n18583) );
  AOI22_X1 U21647 ( .A1(n18535), .A2(n18586), .B1(n18534), .B2(n18583), .ZN(
        n18542) );
  AOI22_X1 U21648 ( .A1(n18539), .A2(n18538), .B1(n18537), .B2(n18536), .ZN(
        n18589) );
  AOI22_X1 U21649 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18589), .B1(
        n18540), .B2(n18569), .ZN(n18541) );
  OAI211_X1 U21650 ( .C1(n18544), .C2(n18543), .A(n18542), .B(n18541), .ZN(
        P3_U2988) );
  AOI22_X1 U21651 ( .A1(n18586), .A2(n18546), .B1(n18545), .B2(n18583), .ZN(
        n18549) );
  AOI22_X1 U21652 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18589), .B1(
        n18588), .B2(n18547), .ZN(n18548) );
  OAI211_X1 U21653 ( .C1(n18550), .C2(n18592), .A(n18549), .B(n18548), .ZN(
        P3_U2989) );
  AOI22_X1 U21654 ( .A1(n18586), .A2(n18552), .B1(n18551), .B2(n18583), .ZN(
        n18555) );
  AOI22_X1 U21655 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18589), .B1(
        n18588), .B2(n18553), .ZN(n18554) );
  OAI211_X1 U21656 ( .C1(n18556), .C2(n18592), .A(n18555), .B(n18554), .ZN(
        P3_U2990) );
  AOI22_X1 U21657 ( .A1(n18558), .A2(n18569), .B1(n18557), .B2(n18583), .ZN(
        n18561) );
  AOI22_X1 U21658 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18589), .B1(
        n18588), .B2(n18559), .ZN(n18560) );
  OAI211_X1 U21659 ( .C1(n18576), .C2(n18562), .A(n18561), .B(n18560), .ZN(
        P3_U2991) );
  AOI22_X1 U21660 ( .A1(n18564), .A2(n18569), .B1(n18563), .B2(n18583), .ZN(
        n18567) );
  AOI22_X1 U21661 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18589), .B1(
        n18588), .B2(n18565), .ZN(n18566) );
  OAI211_X1 U21662 ( .C1(n18576), .C2(n18568), .A(n18567), .B(n18566), .ZN(
        P3_U2992) );
  AOI22_X1 U21663 ( .A1(n18571), .A2(n18583), .B1(n18570), .B2(n18569), .ZN(
        n18574) );
  AOI22_X1 U21664 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18589), .B1(
        n18588), .B2(n18572), .ZN(n18573) );
  OAI211_X1 U21665 ( .C1(n18576), .C2(n18575), .A(n18574), .B(n18573), .ZN(
        P3_U2993) );
  AOI22_X1 U21666 ( .A1(n18586), .A2(n18578), .B1(n18577), .B2(n18583), .ZN(
        n18581) );
  AOI22_X1 U21667 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18589), .B1(
        n18588), .B2(n18579), .ZN(n18580) );
  OAI211_X1 U21668 ( .C1(n18582), .C2(n18592), .A(n18581), .B(n18580), .ZN(
        P3_U2994) );
  AOI22_X1 U21669 ( .A1(n18586), .A2(n18585), .B1(n18584), .B2(n18583), .ZN(
        n18591) );
  AOI22_X1 U21670 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18589), .B1(
        n18588), .B2(n18587), .ZN(n18590) );
  OAI211_X1 U21671 ( .C1(n18593), .C2(n18592), .A(n18591), .B(n18590), .ZN(
        P3_U2995) );
  NOR2_X1 U21672 ( .A1(n18627), .A2(n18594), .ZN(n18597) );
  OAI222_X1 U21673 ( .A1(n18600), .A2(n18599), .B1(n18598), .B2(n18597), .C1(
        n18596), .C2(n18595), .ZN(n18805) );
  OAI21_X1 U21674 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18601), .ZN(n18602) );
  OAI211_X1 U21675 ( .C1(n18604), .C2(n18628), .A(n18603), .B(n18602), .ZN(
        n18649) );
  NOR2_X1 U21676 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18605), .ZN(
        n18632) );
  INV_X1 U21677 ( .A(n18632), .ZN(n18606) );
  AOI22_X1 U21678 ( .A1(n18612), .A2(n18606), .B1(n18627), .B2(n18611), .ZN(
        n18607) );
  NOR2_X1 U21679 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18607), .ZN(
        n18765) );
  OAI21_X1 U21680 ( .B1(n18610), .B2(n18609), .A(n18608), .ZN(n18620) );
  OAI21_X1 U21681 ( .B1(n18612), .B2(n18631), .A(n18611), .ZN(n18613) );
  AOI21_X1 U21682 ( .B1(n18620), .B2(n18614), .A(n18613), .ZN(n18766) );
  NAND2_X1 U21683 ( .A1(n18628), .A2(n18766), .ZN(n18615) );
  AOI22_X1 U21684 ( .A1(n18628), .A2(n18765), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18615), .ZN(n18647) );
  INV_X1 U21685 ( .A(n18628), .ZN(n18639) );
  NOR2_X1 U21686 ( .A1(n18616), .A2(n18793), .ZN(n18617) );
  OAI21_X1 U21687 ( .B1(n18617), .B2(n18619), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18625) );
  OAI221_X1 U21688 ( .B1(n18620), .B2(n18786), .C1(n18620), .C2(n18619), .A(
        n18618), .ZN(n18624) );
  OAI211_X1 U21689 ( .C1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n18622), .B(n18621), .ZN(
        n18623) );
  OAI221_X1 U21690 ( .B1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B2(n18625), 
        .C1(n11361), .C2(n18624), .A(n18623), .ZN(n18626) );
  AOI21_X1 U21691 ( .B1(n18627), .B2(n18774), .A(n18626), .ZN(n18776) );
  AOI22_X1 U21692 ( .A1(n18639), .A2(n11361), .B1(n18776), .B2(n18628), .ZN(
        n18643) );
  NOR2_X1 U21693 ( .A1(n18630), .A2(n18629), .ZN(n18633) );
  AOI22_X1 U21694 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18631), .B1(
        n18633), .B2(n18793), .ZN(n18788) );
  OAI22_X1 U21695 ( .A1(n18633), .A2(n18780), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18632), .ZN(n18784) );
  OR3_X1 U21696 ( .A1(n18788), .A2(n18636), .A3(n18634), .ZN(n18635) );
  AOI22_X1 U21697 ( .A1(n18788), .A2(n18636), .B1(n18784), .B2(n18635), .ZN(
        n18638) );
  OAI21_X1 U21698 ( .B1(n18639), .B2(n18638), .A(n18637), .ZN(n18642) );
  AND2_X1 U21699 ( .A1(n18643), .A2(n18642), .ZN(n18640) );
  OAI221_X1 U21700 ( .B1(n18643), .B2(n18642), .C1(n18641), .C2(n18640), .A(
        n18644), .ZN(n18646) );
  AOI21_X1 U21701 ( .B1(n18644), .B2(n20792), .A(n18643), .ZN(n18645) );
  AOI222_X1 U21702 ( .A1(n18647), .A2(n18646), .B1(n18647), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18646), .C2(n18645), .ZN(
        n18648) );
  NOR4_X1 U21703 ( .A1(n18650), .A2(n18805), .A3(n18649), .A4(n18648), .ZN(
        n18660) );
  INV_X1 U21704 ( .A(n18775), .ZN(n18787) );
  NOR2_X1 U21705 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18817) );
  AOI22_X1 U21706 ( .A1(n18787), .A2(n18817), .B1(n18681), .B2(n18807), .ZN(
        n18651) );
  INV_X1 U21707 ( .A(n18651), .ZN(n18657) );
  OAI211_X1 U21708 ( .C1(n18654), .C2(n18653), .A(n18652), .B(n18660), .ZN(
        n18762) );
  OAI21_X1 U21709 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18815), .A(n18762), 
        .ZN(n18663) );
  NOR2_X1 U21710 ( .A1(n18655), .A2(n18663), .ZN(n18656) );
  MUX2_X1 U21711 ( .A(n18657), .B(n18656), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18659) );
  OAI211_X1 U21712 ( .C1(n18660), .C2(n18811), .A(n18659), .B(n18658), .ZN(
        P3_U2996) );
  NAND2_X1 U21713 ( .A1(n18681), .A2(n18807), .ZN(n18666) );
  NAND3_X1 U21714 ( .A1(n18681), .A2(n18668), .A3(n18661), .ZN(n18671) );
  OR3_X1 U21715 ( .A1(n18664), .A2(n18663), .A3(n18662), .ZN(n18665) );
  NAND4_X1 U21716 ( .A1(n18667), .A2(n18666), .A3(n18671), .A4(n18665), .ZN(
        P3_U2997) );
  OR3_X1 U21717 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18669), .A3(n18668), 
        .ZN(n18670) );
  AND3_X1 U21718 ( .A1(n18671), .A2(n18761), .A3(n18670), .ZN(P3_U2998) );
  AND2_X1 U21719 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18672), .ZN(
        P3_U2999) );
  AND2_X1 U21720 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18672), .ZN(
        P3_U3000) );
  AND2_X1 U21721 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18672), .ZN(
        P3_U3001) );
  AND2_X1 U21722 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18672), .ZN(
        P3_U3002) );
  AND2_X1 U21723 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18672), .ZN(
        P3_U3003) );
  AND2_X1 U21724 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18672), .ZN(
        P3_U3004) );
  AND2_X1 U21725 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18672), .ZN(
        P3_U3005) );
  AND2_X1 U21726 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18672), .ZN(
        P3_U3006) );
  AND2_X1 U21727 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18672), .ZN(
        P3_U3007) );
  AND2_X1 U21728 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18672), .ZN(
        P3_U3008) );
  AND2_X1 U21729 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18672), .ZN(
        P3_U3009) );
  AND2_X1 U21730 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18672), .ZN(
        P3_U3010) );
  AND2_X1 U21731 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18672), .ZN(
        P3_U3011) );
  AND2_X1 U21732 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18672), .ZN(
        P3_U3012) );
  AND2_X1 U21733 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18672), .ZN(
        P3_U3013) );
  AND2_X1 U21734 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18672), .ZN(
        P3_U3014) );
  AND2_X1 U21735 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18672), .ZN(
        P3_U3015) );
  AND2_X1 U21736 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18672), .ZN(
        P3_U3016) );
  AND2_X1 U21737 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18672), .ZN(
        P3_U3017) );
  AND2_X1 U21738 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18672), .ZN(
        P3_U3018) );
  AND2_X1 U21739 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18672), .ZN(
        P3_U3019) );
  AND2_X1 U21740 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18672), .ZN(
        P3_U3020) );
  AND2_X1 U21741 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18672), .ZN(P3_U3021) );
  AND2_X1 U21742 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18672), .ZN(P3_U3022) );
  AND2_X1 U21743 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18672), .ZN(P3_U3023) );
  AND2_X1 U21744 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18672), .ZN(P3_U3024) );
  AND2_X1 U21745 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18672), .ZN(P3_U3025) );
  AND2_X1 U21746 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18672), .ZN(P3_U3026) );
  AND2_X1 U21747 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18672), .ZN(P3_U3027) );
  AND2_X1 U21748 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18672), .ZN(P3_U3028) );
  OAI21_X1 U21749 ( .B1(n18673), .B2(n20670), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18674) );
  AOI22_X1 U21750 ( .A1(n18688), .A2(n18690), .B1(n18823), .B2(n18674), .ZN(
        n18676) );
  INV_X1 U21751 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18675) );
  NAND3_X1 U21752 ( .A1(NA), .A2(n18688), .A3(n18675), .ZN(n18683) );
  OAI211_X1 U21753 ( .C1(n18677), .C2(n18815), .A(n18676), .B(n18683), .ZN(
        P3_U3029) );
  AOI21_X1 U21754 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(HOLD), .A(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18678) );
  AOI21_X1 U21755 ( .B1(HOLD), .B2(P3_STATE_REG_2__SCAN_IN), .A(n18678), .ZN(
        n18679) );
  AOI22_X1 U21756 ( .A1(n18681), .A2(P3_STATE_REG_1__SCAN_IN), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n18679), .ZN(n18680) );
  NAND2_X1 U21757 ( .A1(n18680), .A2(n18812), .ZN(P3_U3030) );
  NAND2_X1 U21758 ( .A1(n18681), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18684) );
  INV_X1 U21759 ( .A(n18684), .ZN(n18682) );
  AOI21_X1 U21760 ( .B1(n18688), .B2(n18683), .A(n18682), .ZN(n18689) );
  NOR2_X1 U21761 ( .A1(n18690), .A2(n20670), .ZN(n18686) );
  OAI22_X1 U21762 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18684), .ZN(n18685) );
  OAI22_X1 U21763 ( .A1(n18686), .A2(n18685), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18687) );
  OAI22_X1 U21764 ( .A1(n18689), .A2(n18690), .B1(n18688), .B2(n18687), .ZN(
        P3_U3031) );
  OAI222_X1 U21765 ( .A1(n18796), .A2(n18752), .B1(n18691), .B2(n18822), .C1(
        n18692), .C2(n18738), .ZN(P3_U3032) );
  INV_X1 U21766 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18694) );
  OAI222_X1 U21767 ( .A1(n18738), .A2(n18694), .B1(n18693), .B2(n18822), .C1(
        n18692), .C2(n18752), .ZN(P3_U3033) );
  OAI222_X1 U21768 ( .A1(n18738), .A2(n18696), .B1(n18695), .B2(n18822), .C1(
        n18694), .C2(n18752), .ZN(P3_U3034) );
  INV_X1 U21769 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18698) );
  OAI222_X1 U21770 ( .A1(n18738), .A2(n18698), .B1(n18697), .B2(n18822), .C1(
        n18696), .C2(n18752), .ZN(P3_U3035) );
  OAI222_X1 U21771 ( .A1(n18738), .A2(n18700), .B1(n18699), .B2(n18822), .C1(
        n18698), .C2(n18752), .ZN(P3_U3036) );
  OAI222_X1 U21772 ( .A1(n18738), .A2(n18702), .B1(n18701), .B2(n18822), .C1(
        n18700), .C2(n18752), .ZN(P3_U3037) );
  OAI222_X1 U21773 ( .A1(n18738), .A2(n18705), .B1(n18703), .B2(n18822), .C1(
        n18702), .C2(n18752), .ZN(P3_U3038) );
  OAI222_X1 U21774 ( .A1(n18705), .A2(n18752), .B1(n18704), .B2(n18822), .C1(
        n18706), .C2(n18738), .ZN(P3_U3039) );
  OAI222_X1 U21775 ( .A1(n18738), .A2(n18708), .B1(n18707), .B2(n18822), .C1(
        n18706), .C2(n18752), .ZN(P3_U3040) );
  INV_X1 U21776 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18710) );
  OAI222_X1 U21777 ( .A1(n18738), .A2(n18710), .B1(n18709), .B2(n18822), .C1(
        n18708), .C2(n18752), .ZN(P3_U3041) );
  OAI222_X1 U21778 ( .A1(n18738), .A2(n18712), .B1(n18711), .B2(n18822), .C1(
        n18710), .C2(n18752), .ZN(P3_U3042) );
  OAI222_X1 U21779 ( .A1(n18738), .A2(n18714), .B1(n18713), .B2(n18822), .C1(
        n18712), .C2(n18752), .ZN(P3_U3043) );
  OAI222_X1 U21780 ( .A1(n18738), .A2(n18717), .B1(n18715), .B2(n18822), .C1(
        n18714), .C2(n18752), .ZN(P3_U3044) );
  OAI222_X1 U21781 ( .A1(n18717), .A2(n18752), .B1(n18716), .B2(n18822), .C1(
        n18718), .C2(n18738), .ZN(P3_U3045) );
  OAI222_X1 U21782 ( .A1(n18738), .A2(n18720), .B1(n18719), .B2(n18822), .C1(
        n18718), .C2(n18752), .ZN(P3_U3046) );
  INV_X1 U21783 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18723) );
  OAI222_X1 U21784 ( .A1(n18738), .A2(n18723), .B1(n18721), .B2(n18822), .C1(
        n18720), .C2(n18752), .ZN(P3_U3047) );
  OAI222_X1 U21785 ( .A1(n18723), .A2(n18752), .B1(n18722), .B2(n18822), .C1(
        n18724), .C2(n18738), .ZN(P3_U3048) );
  OAI222_X1 U21786 ( .A1(n18738), .A2(n18726), .B1(n18725), .B2(n18822), .C1(
        n18724), .C2(n18752), .ZN(P3_U3049) );
  OAI222_X1 U21787 ( .A1(n18738), .A2(n18729), .B1(n18727), .B2(n18822), .C1(
        n18726), .C2(n18752), .ZN(P3_U3050) );
  OAI222_X1 U21788 ( .A1(n18729), .A2(n18752), .B1(n18728), .B2(n18822), .C1(
        n18730), .C2(n18738), .ZN(P3_U3051) );
  OAI222_X1 U21789 ( .A1(n18738), .A2(n18732), .B1(n18731), .B2(n18822), .C1(
        n18730), .C2(n18752), .ZN(P3_U3052) );
  OAI222_X1 U21790 ( .A1(n18738), .A2(n18734), .B1(n18733), .B2(n18822), .C1(
        n18732), .C2(n18752), .ZN(P3_U3053) );
  OAI222_X1 U21791 ( .A1(n18738), .A2(n18736), .B1(n18735), .B2(n18822), .C1(
        n18734), .C2(n18752), .ZN(P3_U3054) );
  OAI222_X1 U21792 ( .A1(n18738), .A2(n18739), .B1(n18737), .B2(n18822), .C1(
        n18736), .C2(n18752), .ZN(P3_U3055) );
  OAI222_X1 U21793 ( .A1(n18738), .A2(n18741), .B1(n18740), .B2(n18822), .C1(
        n18739), .C2(n18752), .ZN(P3_U3056) );
  OAI222_X1 U21794 ( .A1(n18738), .A2(n18743), .B1(n18742), .B2(n18822), .C1(
        n18741), .C2(n18752), .ZN(P3_U3057) );
  OAI222_X1 U21795 ( .A1(n18738), .A2(n18746), .B1(n18744), .B2(n18822), .C1(
        n18743), .C2(n18752), .ZN(P3_U3058) );
  OAI222_X1 U21796 ( .A1(n18746), .A2(n18752), .B1(n18745), .B2(n18822), .C1(
        n18747), .C2(n18738), .ZN(P3_U3059) );
  OAI222_X1 U21797 ( .A1(n18738), .A2(n18751), .B1(n18748), .B2(n18822), .C1(
        n18747), .C2(n18752), .ZN(P3_U3060) );
  OAI222_X1 U21798 ( .A1(n18752), .A2(n18751), .B1(n18750), .B2(n18822), .C1(
        n18749), .C2(n18738), .ZN(P3_U3061) );
  OAI22_X1 U21799 ( .A1(n18823), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18822), .ZN(n18753) );
  INV_X1 U21800 ( .A(n18753), .ZN(P3_U3274) );
  OAI22_X1 U21801 ( .A1(n18823), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18822), .ZN(n18754) );
  INV_X1 U21802 ( .A(n18754), .ZN(P3_U3275) );
  OAI22_X1 U21803 ( .A1(n18823), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18822), .ZN(n18755) );
  INV_X1 U21804 ( .A(n18755), .ZN(P3_U3276) );
  OAI22_X1 U21805 ( .A1(n18823), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18822), .ZN(n18756) );
  INV_X1 U21806 ( .A(n18756), .ZN(P3_U3277) );
  OAI21_X1 U21807 ( .B1(n18760), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18758), 
        .ZN(n18757) );
  INV_X1 U21808 ( .A(n18757), .ZN(P3_U3280) );
  OAI21_X1 U21809 ( .B1(n18760), .B2(n18759), .A(n18758), .ZN(P3_U3281) );
  OAI221_X1 U21810 ( .B1(n18763), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18763), 
        .C2(n18762), .A(n18761), .ZN(P3_U3282) );
  AOI22_X1 U21811 ( .A1(n18789), .A2(n18765), .B1(n18787), .B2(n18764), .ZN(
        n18770) );
  OAI21_X1 U21812 ( .B1(n18825), .B2(n18766), .A(n18791), .ZN(n18767) );
  INV_X1 U21813 ( .A(n18767), .ZN(n18769) );
  OAI22_X1 U21814 ( .A1(n18794), .A2(n18770), .B1(n18769), .B2(n18768), .ZN(
        P3_U3285) );
  OAI22_X1 U21815 ( .A1(n18772), .A2(n18771), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18782) );
  INV_X1 U21816 ( .A(n18782), .ZN(n18778) );
  NOR2_X1 U21817 ( .A1(n18773), .A2(n18790), .ZN(n18781) );
  OAI22_X1 U21818 ( .A1(n18776), .A2(n18825), .B1(n18775), .B2(n18774), .ZN(
        n18777) );
  AOI21_X1 U21819 ( .B1(n18778), .B2(n18781), .A(n18777), .ZN(n18779) );
  AOI22_X1 U21820 ( .A1(n18794), .A2(n11361), .B1(n18779), .B2(n18791), .ZN(
        P3_U3288) );
  INV_X1 U21821 ( .A(n18780), .ZN(n18783) );
  AOI222_X1 U21822 ( .A1(n18784), .A2(n18789), .B1(n18787), .B2(n18783), .C1(
        n18782), .C2(n18781), .ZN(n18785) );
  AOI22_X1 U21823 ( .A1(n18794), .A2(n18786), .B1(n18785), .B2(n18791), .ZN(
        P3_U3289) );
  AOI222_X1 U21824 ( .A1(n18790), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18789), 
        .B2(n18788), .C1(n18793), .C2(n18787), .ZN(n18792) );
  AOI22_X1 U21825 ( .A1(n18794), .A2(n18793), .B1(n18792), .B2(n18791), .ZN(
        P3_U3290) );
  AOI21_X1 U21826 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18795) );
  OAI22_X1 U21827 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n18796), .B1(
        P3_REIP_REG_1__SCAN_IN), .B2(n18795), .ZN(n18798) );
  INV_X1 U21828 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18797) );
  AOI22_X1 U21829 ( .A1(n18802), .A2(n18798), .B1(n18797), .B2(n18799), .ZN(
        P3_U3292) );
  NOR2_X1 U21830 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n18801) );
  INV_X1 U21831 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18800) );
  AOI22_X1 U21832 ( .A1(n18802), .A2(n18801), .B1(n18800), .B2(n18799), .ZN(
        P3_U3293) );
  INV_X1 U21833 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18803) );
  AOI22_X1 U21834 ( .A1(n18822), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18803), 
        .B2(n18823), .ZN(P3_U3294) );
  MUX2_X1 U21835 ( .A(P3_MORE_REG_SCAN_IN), .B(n18805), .S(n18804), .Z(
        P3_U3295) );
  AOI21_X1 U21836 ( .B1(n18815), .B2(n18807), .A(n18806), .ZN(n18808) );
  INV_X1 U21837 ( .A(n18808), .ZN(n18809) );
  AOI21_X1 U21838 ( .B1(n18811), .B2(n18810), .A(n18809), .ZN(n18821) );
  AOI21_X1 U21839 ( .B1(n18814), .B2(n18813), .A(n18812), .ZN(n18816) );
  OAI211_X1 U21840 ( .C1(n18826), .C2(n18816), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18815), .ZN(n18818) );
  AOI21_X1 U21841 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18818), .A(n18817), 
        .ZN(n18820) );
  NAND2_X1 U21842 ( .A1(n18821), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18819) );
  OAI21_X1 U21843 ( .B1(n18821), .B2(n18820), .A(n18819), .ZN(P3_U3296) );
  OAI22_X1 U21844 ( .A1(n18823), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18822), .ZN(n18824) );
  INV_X1 U21845 ( .A(n18824), .ZN(P3_U3297) );
  OAI21_X1 U21846 ( .B1(n18825), .B2(P3_STATE2_REG_2__SCAN_IN), .A(n18827), 
        .ZN(n18830) );
  OAI22_X1 U21847 ( .A1(n18830), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18827), 
        .B2(n18826), .ZN(n18828) );
  INV_X1 U21848 ( .A(n18828), .ZN(P3_U3298) );
  OAI21_X1 U21849 ( .B1(n18830), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n18829), 
        .ZN(n18831) );
  INV_X1 U21850 ( .A(n18831), .ZN(P3_U3299) );
  INV_X1 U21851 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19681) );
  INV_X1 U21852 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19700) );
  NAND2_X1 U21853 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19700), .ZN(n19689) );
  INV_X1 U21854 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19692) );
  NAND2_X1 U21855 ( .A1(n19681), .A2(n19692), .ZN(n19685) );
  OAI21_X1 U21856 ( .B1(n19681), .B2(n19689), .A(n19685), .ZN(n19761) );
  AOI21_X1 U21857 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19761), .ZN(n18832) );
  INV_X1 U21858 ( .A(n18832), .ZN(P2_U2815) );
  INV_X1 U21859 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18835) );
  OAI22_X1 U21860 ( .A1(n19819), .A2(n18835), .B1(n18834), .B2(n18833), .ZN(
        P2_U2816) );
  INV_X2 U21861 ( .A(n19838), .ZN(n19837) );
  AOI22_X1 U21862 ( .A1(n19837), .A2(n18835), .B1(P2_D_C_N_REG_SCAN_IN), .B2(
        n19838), .ZN(n18836) );
  OAI21_X1 U21863 ( .B1(P2_STATE_REG_2__SCAN_IN), .B2(n19685), .A(n18836), 
        .ZN(P2_U2817) );
  OAI21_X1 U21864 ( .B1(n19691), .B2(BS16), .A(n19761), .ZN(n19759) );
  OAI21_X1 U21865 ( .B1(n19761), .B2(n19382), .A(n19759), .ZN(P2_U2818) );
  NOR4_X1 U21866 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18840) );
  NOR4_X1 U21867 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18839) );
  NOR4_X1 U21868 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18838) );
  NOR4_X1 U21869 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18837) );
  NAND4_X1 U21870 ( .A1(n18840), .A2(n18839), .A3(n18838), .A4(n18837), .ZN(
        n18846) );
  NOR4_X1 U21871 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_4__SCAN_IN), .A3(P2_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_6__SCAN_IN), .ZN(n18844) );
  AOI211_X1 U21872 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_11__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18843) );
  NOR4_X1 U21873 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n18842) );
  NOR4_X1 U21874 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_8__SCAN_IN), .A3(P2_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_10__SCAN_IN), .ZN(n18841) );
  NAND4_X1 U21875 ( .A1(n18844), .A2(n18843), .A3(n18842), .A4(n18841), .ZN(
        n18845) );
  NOR2_X1 U21876 ( .A1(n18846), .A2(n18845), .ZN(n18857) );
  INV_X1 U21877 ( .A(n18857), .ZN(n18855) );
  NOR2_X1 U21878 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18855), .ZN(n18849) );
  INV_X1 U21879 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18847) );
  AOI22_X1 U21880 ( .A1(n18849), .A2(n18850), .B1(n18855), .B2(n18847), .ZN(
        P2_U2820) );
  OR3_X1 U21881 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18854) );
  INV_X1 U21882 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18848) );
  AOI22_X1 U21883 ( .A1(n18849), .A2(n18854), .B1(n18855), .B2(n18848), .ZN(
        P2_U2821) );
  INV_X1 U21884 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19760) );
  NAND2_X1 U21885 ( .A1(n18849), .A2(n19760), .ZN(n18853) );
  OAI21_X1 U21886 ( .B1(n18850), .B2(n19702), .A(n18857), .ZN(n18851) );
  OAI21_X1 U21887 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18857), .A(n18851), 
        .ZN(n18852) );
  OAI221_X1 U21888 ( .B1(n18853), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18853), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18852), .ZN(P2_U2822) );
  INV_X1 U21889 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18856) );
  OAI221_X1 U21890 ( .B1(n18857), .B2(n18856), .C1(n18855), .C2(n18854), .A(
        n18853), .ZN(P2_U2823) );
  OAI22_X1 U21891 ( .A1(n18978), .A2(n19733), .B1(n19028), .B2(n18858), .ZN(
        n18861) );
  NOR2_X1 U21892 ( .A1(n18859), .A2(n19004), .ZN(n18860) );
  AOI211_X1 U21893 ( .C1(P2_EBX_REG_21__SCAN_IN), .C2(n19018), .A(n18861), .B(
        n18860), .ZN(n18862) );
  OAI21_X1 U21894 ( .B1(n18863), .B2(n18984), .A(n18862), .ZN(n18868) );
  AOI211_X1 U21895 ( .C1(n18866), .C2(n18865), .A(n18864), .B(n19677), .ZN(
        n18867) );
  NOR2_X1 U21896 ( .A1(n18868), .A2(n18867), .ZN(n18869) );
  OAI21_X1 U21897 ( .B1(n18870), .B2(n19001), .A(n18869), .ZN(P2_U2834) );
  AOI22_X1 U21898 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18997), .B1(
        P2_REIP_REG_20__SCAN_IN), .B2(n19017), .ZN(n18883) );
  INV_X1 U21899 ( .A(n18871), .ZN(n18872) );
  AOI22_X1 U21900 ( .A1(n18872), .A2(n19022), .B1(P2_EBX_REG_20__SCAN_IN), 
        .B2(n19018), .ZN(n18882) );
  OAI22_X1 U21901 ( .A1(n18874), .A2(n19004), .B1(n18873), .B2(n19001), .ZN(
        n18875) );
  INV_X1 U21902 ( .A(n18875), .ZN(n18881) );
  AOI21_X1 U21903 ( .B1(n18878), .B2(n18877), .A(n18876), .ZN(n18879) );
  NAND2_X1 U21904 ( .A1(n18993), .A2(n18879), .ZN(n18880) );
  NAND4_X1 U21905 ( .A1(n18883), .A2(n18882), .A3(n18881), .A4(n18880), .ZN(
        P2_U2835) );
  AOI22_X1 U21906 ( .A1(n18884), .A2(n19022), .B1(P2_EBX_REG_17__SCAN_IN), 
        .B2(n19018), .ZN(n18885) );
  OAI211_X1 U21907 ( .C1(n19727), .C2(n18978), .A(n18885), .B(n19155), .ZN(
        n18889) );
  OAI22_X1 U21908 ( .A1(n18887), .A2(n19001), .B1(n19004), .B2(n18886), .ZN(
        n18888) );
  AOI211_X1 U21909 ( .C1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(n18997), .A(
        n18889), .B(n18888), .ZN(n18895) );
  INV_X1 U21910 ( .A(n18890), .ZN(n18892) );
  OAI221_X1 U21911 ( .B1(n18893), .B2(n18892), .C1(n18891), .C2(n18890), .A(
        n18993), .ZN(n18894) );
  NAND2_X1 U21912 ( .A1(n18895), .A2(n18894), .ZN(P2_U2838) );
  NAND2_X1 U21913 ( .A1(n9838), .A2(n18896), .ZN(n18897) );
  XOR2_X1 U21914 ( .A(n18898), .B(n18897), .Z(n18907) );
  AOI22_X1 U21915 ( .A1(n19018), .A2(P2_EBX_REG_16__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n18997), .ZN(n18899) );
  OAI21_X1 U21916 ( .B1(n18900), .B2(n18984), .A(n18899), .ZN(n18901) );
  AOI211_X1 U21917 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n19017), .A(n18902), 
        .B(n18901), .ZN(n18906) );
  NOR2_X1 U21918 ( .A1(n18903), .A2(n19004), .ZN(n18904) );
  AOI21_X1 U21919 ( .B1(n19042), .B2(n19016), .A(n18904), .ZN(n18905) );
  OAI211_X1 U21920 ( .C1(n19677), .C2(n18907), .A(n18906), .B(n18905), .ZN(
        P2_U2839) );
  AOI22_X1 U21921 ( .A1(n18908), .A2(n19022), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n19018), .ZN(n18909) );
  OAI211_X1 U21922 ( .C1(n10788), .C2(n18978), .A(n18909), .B(n19155), .ZN(
        n18910) );
  AOI21_X1 U21923 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n18997), .A(
        n18910), .ZN(n18917) );
  NAND2_X1 U21924 ( .A1(n9838), .A2(n18911), .ZN(n18912) );
  XOR2_X1 U21925 ( .A(n18913), .B(n18912), .Z(n18915) );
  AOI22_X1 U21926 ( .A1(n18915), .A2(n18993), .B1(n19020), .B2(n18914), .ZN(
        n18916) );
  OAI211_X1 U21927 ( .C1(n19050), .C2(n19001), .A(n18917), .B(n18916), .ZN(
        P2_U2841) );
  NOR2_X1 U21928 ( .A1(n11247), .A2(n18918), .ZN(n18920) );
  XOR2_X1 U21929 ( .A(n18920), .B(n18919), .Z(n18927) );
  AOI22_X1 U21930 ( .A1(n18921), .A2(n19022), .B1(P2_EBX_REG_13__SCAN_IN), 
        .B2(n19018), .ZN(n18922) );
  OAI211_X1 U21931 ( .C1(n11011), .C2(n18978), .A(n18922), .B(n19155), .ZN(
        n18925) );
  OAI22_X1 U21932 ( .A1(n19052), .A2(n19001), .B1(n19004), .B2(n18923), .ZN(
        n18924) );
  AOI211_X1 U21933 ( .C1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .C2(n18997), .A(
        n18925), .B(n18924), .ZN(n18926) );
  OAI21_X1 U21934 ( .B1(n19677), .B2(n18927), .A(n18926), .ZN(P2_U2842) );
  NAND2_X1 U21935 ( .A1(n9838), .A2(n18928), .ZN(n18945) );
  XOR2_X1 U21936 ( .A(n18929), .B(n18945), .Z(n18937) );
  AOI22_X1 U21937 ( .A1(n18930), .A2(n19022), .B1(P2_EBX_REG_12__SCAN_IN), 
        .B2(n19018), .ZN(n18931) );
  OAI211_X1 U21938 ( .C1(n11008), .C2(n18978), .A(n18931), .B(n19155), .ZN(
        n18932) );
  AOI21_X1 U21939 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18997), .A(
        n18932), .ZN(n18936) );
  AOI22_X1 U21940 ( .A1(n18934), .A2(n19016), .B1(n19020), .B2(n18933), .ZN(
        n18935) );
  OAI211_X1 U21941 ( .C1(n19677), .C2(n18937), .A(n18936), .B(n18935), .ZN(
        P2_U2843) );
  AOI22_X1 U21942 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n18997), .B1(
        P2_REIP_REG_11__SCAN_IN), .B2(n19017), .ZN(n18938) );
  OAI211_X1 U21943 ( .C1(n19004), .C2(n18939), .A(n18938), .B(n19155), .ZN(
        n18940) );
  AOI21_X1 U21944 ( .B1(n19018), .B2(P2_EBX_REG_11__SCAN_IN), .A(n18940), .ZN(
        n18943) );
  NAND2_X1 U21945 ( .A1(n18941), .A2(n19022), .ZN(n18942) );
  OAI211_X1 U21946 ( .C1(n19056), .C2(n19001), .A(n18943), .B(n18942), .ZN(
        n18944) );
  INV_X1 U21947 ( .A(n18944), .ZN(n18949) );
  INV_X1 U21948 ( .A(n18945), .ZN(n18946) );
  OAI211_X1 U21949 ( .C1(n18947), .C2(n18950), .A(n18993), .B(n18946), .ZN(
        n18948) );
  OAI211_X1 U21950 ( .C1(n19027), .C2(n18950), .A(n18949), .B(n18948), .ZN(
        P2_U2844) );
  AOI22_X1 U21951 ( .A1(n18951), .A2(n19022), .B1(P2_EBX_REG_10__SCAN_IN), 
        .B2(n19018), .ZN(n18952) );
  OAI211_X1 U21952 ( .C1(n19718), .C2(n18978), .A(n18952), .B(n19155), .ZN(
        n18953) );
  AOI21_X1 U21953 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18997), .A(
        n18953), .ZN(n18960) );
  NAND2_X1 U21954 ( .A1(n9838), .A2(n18954), .ZN(n18955) );
  XNOR2_X1 U21955 ( .A(n18956), .B(n18955), .ZN(n18958) );
  AOI22_X1 U21956 ( .A1(n18958), .A2(n18993), .B1(n19020), .B2(n18957), .ZN(
        n18959) );
  OAI211_X1 U21957 ( .C1(n19001), .C2(n19059), .A(n18960), .B(n18959), .ZN(
        P2_U2845) );
  NAND2_X1 U21958 ( .A1(n9838), .A2(n18961), .ZN(n18962) );
  XOR2_X1 U21959 ( .A(n18963), .B(n18962), .Z(n18972) );
  AOI22_X1 U21960 ( .A1(n19018), .A2(P2_EBX_REG_8__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18997), .ZN(n18964) );
  OAI21_X1 U21961 ( .B1(n18965), .B2(n18984), .A(n18964), .ZN(n18966) );
  AOI211_X1 U21962 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n19017), .A(n18902), .B(
        n18966), .ZN(n18971) );
  INV_X1 U21963 ( .A(n18967), .ZN(n19064) );
  OAI22_X1 U21964 ( .A1(n18968), .A2(n19004), .B1(n19001), .B2(n19064), .ZN(
        n18969) );
  INV_X1 U21965 ( .A(n18969), .ZN(n18970) );
  OAI211_X1 U21966 ( .C1(n19677), .C2(n18972), .A(n18971), .B(n18970), .ZN(
        P2_U2847) );
  NOR2_X1 U21967 ( .A1(n11247), .A2(n18973), .ZN(n18974) );
  XOR2_X1 U21968 ( .A(n18975), .B(n18974), .Z(n18983) );
  AOI22_X1 U21969 ( .A1(n19022), .A2(n18976), .B1(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18997), .ZN(n18977) );
  OAI211_X1 U21970 ( .C1(n19712), .C2(n18978), .A(n18977), .B(n19155), .ZN(
        n18981) );
  OAI22_X1 U21971 ( .A1(n19066), .A2(n19001), .B1(n19004), .B2(n18979), .ZN(
        n18980) );
  AOI211_X1 U21972 ( .C1(P2_EBX_REG_7__SCAN_IN), .C2(n19018), .A(n18981), .B(
        n18980), .ZN(n18982) );
  OAI21_X1 U21973 ( .B1(n19677), .B2(n18983), .A(n18982), .ZN(P2_U2848) );
  OAI22_X1 U21974 ( .A1(n19002), .A2(n10755), .B1(n18985), .B2(n18984), .ZN(
        n18986) );
  AOI211_X1 U21975 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19017), .A(n18902), .B(
        n18986), .ZN(n18996) );
  NOR2_X1 U21976 ( .A1(n11247), .A2(n18987), .ZN(n18989) );
  XNOR2_X1 U21977 ( .A(n18990), .B(n18989), .ZN(n18994) );
  OAI22_X1 U21978 ( .A1(n19081), .A2(n19001), .B1(n19004), .B2(n18991), .ZN(
        n18992) );
  AOI21_X1 U21979 ( .B1(n18994), .B2(n18993), .A(n18992), .ZN(n18995) );
  OAI211_X1 U21980 ( .C1(n10754), .C2(n19028), .A(n18996), .B(n18995), .ZN(
        P2_U2850) );
  AOI22_X1 U21981 ( .A1(n19022), .A2(n18998), .B1(
        P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n18997), .ZN(n19013) );
  XNOR2_X1 U21982 ( .A(n19000), .B(n18999), .ZN(n19156) );
  OAI22_X1 U21983 ( .A1(n19002), .A2(n10750), .B1(n19001), .B2(n19156), .ZN(
        n19003) );
  AOI211_X1 U21984 ( .C1(P2_REIP_REG_4__SCAN_IN), .C2(n19017), .A(n18902), .B(
        n19003), .ZN(n19012) );
  OAI22_X1 U21985 ( .A1(n19084), .A2(n19005), .B1(n19004), .B2(n19163), .ZN(
        n19006) );
  INV_X1 U21986 ( .A(n19006), .ZN(n19011) );
  AND2_X1 U21987 ( .A1(n9838), .A2(n19007), .ZN(n19009) );
  AOI21_X1 U21988 ( .B1(n19140), .B2(n19009), .A(n19677), .ZN(n19008) );
  OAI21_X1 U21989 ( .B1(n19140), .B2(n19009), .A(n19008), .ZN(n19010) );
  NAND4_X1 U21990 ( .A1(n19013), .A2(n19012), .A3(n19011), .A4(n19010), .ZN(
        P2_U2851) );
  INV_X1 U21991 ( .A(n19014), .ZN(n19015) );
  AOI22_X1 U21992 ( .A1(n19017), .A2(P2_REIP_REG_0__SCAN_IN), .B1(n19016), 
        .B2(n19015), .ZN(n19026) );
  NAND2_X1 U21993 ( .A1(n19018), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n19025) );
  NAND2_X1 U21994 ( .A1(n19020), .A2(n19019), .ZN(n19024) );
  NAND2_X1 U21995 ( .A1(n19022), .A2(n19021), .ZN(n19023) );
  AND4_X1 U21996 ( .A1(n19026), .A2(n19025), .A3(n19024), .A4(n19023), .ZN(
        n19033) );
  NAND2_X1 U21997 ( .A1(n19028), .A2(n19027), .ZN(n19031) );
  AOI22_X1 U21998 ( .A1(n19031), .A2(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19030), .B2(n19029), .ZN(n19032) );
  OAI211_X1 U21999 ( .C1(n19035), .C2(n19034), .A(n19033), .B(n19032), .ZN(
        P2_U2855) );
  AOI22_X1 U22000 ( .A1(n19037), .A2(n19036), .B1(n19098), .B2(
        P2_EAX_REG_16__SCAN_IN), .ZN(n19045) );
  AOI22_X1 U22001 ( .A1(n19039), .A2(BUF1_REG_16__SCAN_IN), .B1(n19038), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n19044) );
  NOR2_X1 U22002 ( .A1(n19040), .A2(n19103), .ZN(n19041) );
  AOI21_X1 U22003 ( .B1(n19042), .B2(n19099), .A(n19041), .ZN(n19043) );
  NAND3_X1 U22004 ( .A1(n19045), .A2(n19044), .A3(n19043), .ZN(P2_U2903) );
  OAI222_X1 U22005 ( .A1(n19048), .A2(n19082), .B1(n19111), .B2(n19069), .C1(
        n19047), .C2(n19107), .ZN(P2_U2904) );
  INV_X1 U22006 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19113) );
  OAI222_X1 U22007 ( .A1(n19050), .A2(n19082), .B1(n19113), .B2(n19069), .C1(
        n19107), .C2(n19049), .ZN(P2_U2905) );
  INV_X1 U22008 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19115) );
  OAI222_X1 U22009 ( .A1(n19052), .A2(n19082), .B1(n19115), .B2(n19069), .C1(
        n19107), .C2(n19051), .ZN(P2_U2906) );
  OAI222_X1 U22010 ( .A1(n19054), .A2(n19082), .B1(n13132), .B2(n19069), .C1(
        n19107), .C2(n19053), .ZN(P2_U2907) );
  INV_X1 U22011 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19118) );
  OAI222_X1 U22012 ( .A1(n19056), .A2(n19082), .B1(n19118), .B2(n19069), .C1(
        n19107), .C2(n19055), .ZN(P2_U2908) );
  AOI22_X1 U22013 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19098), .B1(n19057), 
        .B2(n19071), .ZN(n19058) );
  OAI21_X1 U22014 ( .B1(n19082), .B2(n19059), .A(n19058), .ZN(P2_U2909) );
  INV_X1 U22015 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19121) );
  OAI222_X1 U22016 ( .A1(n19061), .A2(n19082), .B1(n19121), .B2(n19069), .C1(
        n19107), .C2(n19060), .ZN(P2_U2910) );
  AOI22_X1 U22017 ( .A1(P2_EAX_REG_8__SCAN_IN), .A2(n19098), .B1(n19062), .B2(
        n19071), .ZN(n19063) );
  OAI21_X1 U22018 ( .B1(n19082), .B2(n19064), .A(n19063), .ZN(P2_U2911) );
  OAI222_X1 U22019 ( .A1(n19066), .A2(n19082), .B1(n19125), .B2(n19069), .C1(
        n19107), .C2(n19065), .ZN(P2_U2912) );
  INV_X1 U22020 ( .A(n19067), .ZN(n19070) );
  OAI222_X1 U22021 ( .A1(n19070), .A2(n19082), .B1(n19128), .B2(n19069), .C1(
        n19107), .C2(n19068), .ZN(P2_U2913) );
  AOI22_X1 U22022 ( .A1(P2_EAX_REG_5__SCAN_IN), .A2(n19098), .B1(n19072), .B2(
        n19071), .ZN(n19080) );
  AOI21_X1 U22023 ( .B1(n19777), .B2(n19074), .A(n19073), .ZN(n19092) );
  XNOR2_X1 U22024 ( .A(n19076), .B(n19075), .ZN(n19093) );
  NOR2_X1 U22025 ( .A1(n19092), .A2(n19093), .ZN(n19091) );
  NOR2_X1 U22026 ( .A1(n19766), .A2(n19768), .ZN(n19077) );
  OAI21_X1 U22027 ( .B1(n19091), .B2(n19077), .A(n19156), .ZN(n19085) );
  INV_X1 U22028 ( .A(n19084), .ZN(n19078) );
  NAND3_X1 U22029 ( .A1(n19085), .A2(n19078), .A3(n19086), .ZN(n19079) );
  OAI211_X1 U22030 ( .C1(n19082), .C2(n19081), .A(n19080), .B(n19079), .ZN(
        P2_U2914) );
  INV_X1 U22031 ( .A(n19156), .ZN(n19083) );
  AOI22_X1 U22032 ( .A1(n19099), .A2(n19083), .B1(n19098), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n19089) );
  XNOR2_X1 U22033 ( .A(n19085), .B(n19084), .ZN(n19087) );
  NAND2_X1 U22034 ( .A1(n19087), .A2(n19086), .ZN(n19088) );
  OAI211_X1 U22035 ( .C1(n19090), .C2(n19107), .A(n19089), .B(n19088), .ZN(
        P2_U2915) );
  AOI22_X1 U22036 ( .A1(n19768), .A2(n19099), .B1(n19098), .B2(
        P2_EAX_REG_3__SCAN_IN), .ZN(n19096) );
  AOI21_X1 U22037 ( .B1(n19093), .B2(n19092), .A(n19091), .ZN(n19094) );
  OR2_X1 U22038 ( .A1(n19094), .A2(n19103), .ZN(n19095) );
  OAI211_X1 U22039 ( .C1(n19097), .C2(n19107), .A(n19096), .B(n19095), .ZN(
        P2_U2916) );
  AOI22_X1 U22040 ( .A1(n19099), .A2(n19791), .B1(n19098), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19106) );
  AOI21_X1 U22041 ( .B1(n19102), .B2(n19101), .A(n19100), .ZN(n19104) );
  OR2_X1 U22042 ( .A1(n19104), .A2(n19103), .ZN(n19105) );
  OAI211_X1 U22043 ( .C1(n19108), .C2(n19107), .A(n19106), .B(n19105), .ZN(
        P2_U2918) );
  AND2_X1 U22044 ( .A1(n19126), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(P2_U2920)
         );
  AOI22_X1 U22045 ( .A1(n19821), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19110) );
  OAI21_X1 U22046 ( .B1(n19111), .B2(n19139), .A(n19110), .ZN(P2_U2936) );
  AOI22_X1 U22047 ( .A1(n19821), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19112) );
  OAI21_X1 U22048 ( .B1(n19113), .B2(n19139), .A(n19112), .ZN(P2_U2937) );
  AOI22_X1 U22049 ( .A1(n19821), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19114) );
  OAI21_X1 U22050 ( .B1(n19115), .B2(n19139), .A(n19114), .ZN(P2_U2938) );
  AOI22_X1 U22051 ( .A1(n19821), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19116) );
  OAI21_X1 U22052 ( .B1(n13132), .B2(n19139), .A(n19116), .ZN(P2_U2939) );
  AOI22_X1 U22053 ( .A1(n19821), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19117) );
  OAI21_X1 U22054 ( .B1(n19118), .B2(n19139), .A(n19117), .ZN(P2_U2940) );
  AOI22_X1 U22055 ( .A1(n19821), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19119) );
  OAI21_X1 U22056 ( .B1(n10980), .B2(n19139), .A(n19119), .ZN(P2_U2941) );
  AOI22_X1 U22057 ( .A1(n19821), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19120) );
  OAI21_X1 U22058 ( .B1(n19121), .B2(n19139), .A(n19120), .ZN(P2_U2942) );
  AOI22_X1 U22059 ( .A1(n19821), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19122) );
  OAI21_X1 U22060 ( .B1(n19123), .B2(n19139), .A(n19122), .ZN(P2_U2943) );
  AOI22_X1 U22061 ( .A1(n19821), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19124) );
  OAI21_X1 U22062 ( .B1(n19125), .B2(n19139), .A(n19124), .ZN(P2_U2944) );
  AOI22_X1 U22063 ( .A1(n19821), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19127) );
  OAI21_X1 U22064 ( .B1(n19128), .B2(n19139), .A(n19127), .ZN(P2_U2945) );
  INV_X1 U22065 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19130) );
  AOI22_X1 U22066 ( .A1(n19821), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19129) );
  OAI21_X1 U22067 ( .B1(n19130), .B2(n19139), .A(n19129), .ZN(P2_U2946) );
  INV_X1 U22068 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19132) );
  AOI22_X1 U22069 ( .A1(n19821), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19131) );
  OAI21_X1 U22070 ( .B1(n19132), .B2(n19139), .A(n19131), .ZN(P2_U2947) );
  AOI22_X1 U22071 ( .A1(n19821), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19133) );
  OAI21_X1 U22072 ( .B1(n10910), .B2(n19139), .A(n19133), .ZN(P2_U2948) );
  AOI22_X1 U22073 ( .A1(n19821), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19134) );
  OAI21_X1 U22074 ( .B1(n19135), .B2(n19139), .A(n19134), .ZN(P2_U2949) );
  AOI22_X1 U22075 ( .A1(n19821), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19136) );
  OAI21_X1 U22076 ( .B1(n19137), .B2(n19139), .A(n19136), .ZN(P2_U2950) );
  AOI22_X1 U22077 ( .A1(n19821), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19126), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19138) );
  OAI21_X1 U22078 ( .B1(n13122), .B2(n19139), .A(n19138), .ZN(P2_U2951) );
  AOI22_X1 U22079 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n18902), .B1(n19141), 
        .B2(n19140), .ZN(n19153) );
  INV_X1 U22080 ( .A(n19163), .ZN(n19150) );
  XNOR2_X1 U22081 ( .A(n19142), .B(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n19143) );
  XNOR2_X1 U22082 ( .A(n19144), .B(n19143), .ZN(n19168) );
  XNOR2_X1 U22083 ( .A(n19146), .B(n19145), .ZN(n19158) );
  OAI22_X1 U22084 ( .A1(n19168), .A2(n19148), .B1(n19147), .B2(n19158), .ZN(
        n19149) );
  AOI21_X1 U22085 ( .B1(n19151), .B2(n19150), .A(n19149), .ZN(n19152) );
  OAI211_X1 U22086 ( .C1(n10749), .C2(n19154), .A(n19153), .B(n19152), .ZN(
        P2_U3010) );
  INV_X1 U22087 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19706) );
  NOR2_X1 U22088 ( .A1(n19706), .A2(n19155), .ZN(n19160) );
  OAI22_X1 U22089 ( .A1(n19158), .A2(n19157), .B1(n19185), .B2(n19156), .ZN(
        n19159) );
  AOI211_X1 U22090 ( .C1(n19162), .C2(n19161), .A(n19160), .B(n19159), .ZN(
        n19167) );
  OAI22_X1 U22091 ( .A1(n19164), .A2(n19161), .B1(n19179), .B2(n19163), .ZN(
        n19165) );
  INV_X1 U22092 ( .A(n19165), .ZN(n19166) );
  OAI211_X1 U22093 ( .C1(n19174), .C2(n19168), .A(n19167), .B(n19166), .ZN(
        P2_U3042) );
  INV_X1 U22094 ( .A(n19169), .ZN(n19171) );
  NOR2_X1 U22095 ( .A1(n19171), .A2(n19170), .ZN(n19176) );
  INV_X1 U22096 ( .A(n19172), .ZN(n19173) );
  OAI22_X1 U22097 ( .A1(n19176), .A2(n19175), .B1(n19174), .B2(n19173), .ZN(
        n19181) );
  OAI21_X1 U22098 ( .B1(n19179), .B2(n19178), .A(n19177), .ZN(n19180) );
  NOR2_X1 U22099 ( .A1(n19181), .A2(n19180), .ZN(n19184) );
  NAND2_X1 U22100 ( .A1(n19182), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n19183) );
  OAI211_X1 U22101 ( .C1(n19777), .C2(n19185), .A(n19184), .B(n19183), .ZN(
        n19186) );
  INV_X1 U22102 ( .A(n19186), .ZN(n19190) );
  NAND2_X1 U22103 ( .A1(n19188), .A2(n19187), .ZN(n19189) );
  OAI211_X1 U22104 ( .C1(n19192), .C2(n19191), .A(n19190), .B(n19189), .ZN(
        P2_U3044) );
  INV_X1 U22105 ( .A(n19271), .ZN(n19272) );
  NAND2_X1 U22106 ( .A1(n19272), .A2(n19793), .ZN(n19230) );
  NOR2_X1 U22107 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19230), .ZN(
        n19217) );
  AOI22_X1 U22108 ( .A1(n19576), .A2(n19669), .B1(n19573), .B2(n19217), .ZN(
        n19202) );
  NOR3_X1 U22109 ( .A1(n19197), .A2(n19217), .A3(n19528), .ZN(n19196) );
  OAI21_X1 U22110 ( .B1(n19669), .B2(n19241), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19194) );
  NAND2_X1 U22111 ( .A1(n19194), .A2(n19764), .ZN(n19200) );
  AOI221_X1 U22112 ( .B1(n19794), .B2(n19200), .C1(n19794), .C2(n19662), .A(
        n19217), .ZN(n19195) );
  NOR2_X1 U22113 ( .A1(n19662), .A2(n19217), .ZN(n19199) );
  OAI21_X1 U22114 ( .B1(n19197), .B2(n19217), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19198) );
  AOI22_X1 U22115 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19219), .B1(
        n19574), .B2(n19218), .ZN(n19201) );
  OAI211_X1 U22116 ( .C1(n19537), .C2(n19254), .A(n19202), .B(n19201), .ZN(
        P2_U3048) );
  AOI22_X1 U22117 ( .A1(n19638), .A2(n19669), .B1(n14064), .B2(n19217), .ZN(
        n19204) );
  AOI22_X1 U22118 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19219), .B1(
        n19637), .B2(n19218), .ZN(n19203) );
  OAI211_X1 U22119 ( .C1(n19540), .C2(n19254), .A(n19204), .B(n19203), .ZN(
        P2_U3049) );
  AOI22_X1 U22120 ( .A1(n19645), .A2(n19669), .B1(n19643), .B2(n19217), .ZN(
        n19206) );
  AOI22_X1 U22121 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19219), .B1(
        n19644), .B2(n19218), .ZN(n19205) );
  OAI211_X1 U22122 ( .C1(n19543), .C2(n19254), .A(n19206), .B(n19205), .ZN(
        P2_U3050) );
  AOI22_X1 U22123 ( .A1(n19651), .A2(n19669), .B1(n19649), .B2(n19217), .ZN(
        n19209) );
  AOI22_X1 U22124 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19219), .B1(
        n19650), .B2(n19218), .ZN(n19208) );
  OAI211_X1 U22125 ( .C1(n19546), .C2(n19254), .A(n19209), .B(n19208), .ZN(
        P2_U3051) );
  AOI22_X1 U22126 ( .A1(n19658), .A2(n19669), .B1(n19655), .B2(n19217), .ZN(
        n19211) );
  AOI22_X1 U22127 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19219), .B1(
        n19656), .B2(n19218), .ZN(n19210) );
  OAI211_X1 U22128 ( .C1(n19592), .C2(n19254), .A(n19211), .B(n19210), .ZN(
        P2_U3052) );
  AOI22_X1 U22129 ( .A1(n19549), .A2(n19669), .B1(n19593), .B2(n19217), .ZN(
        n19213) );
  AOI22_X1 U22130 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19219), .B1(
        n19594), .B2(n19218), .ZN(n19212) );
  OAI211_X1 U22131 ( .C1(n19552), .C2(n19254), .A(n19213), .B(n19212), .ZN(
        P2_U3053) );
  AOI22_X1 U22132 ( .A1(n19666), .A2(n19669), .B1(n19663), .B2(n19217), .ZN(
        n19215) );
  AOI22_X1 U22133 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19219), .B1(
        n19664), .B2(n19218), .ZN(n19214) );
  OAI211_X1 U22134 ( .C1(n19603), .C2(n19254), .A(n19215), .B(n19214), .ZN(
        P2_U3054) );
  AOI22_X1 U22135 ( .A1(n19629), .A2(n19669), .B1(n19627), .B2(n19217), .ZN(
        n19221) );
  AOI22_X1 U22136 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19219), .B1(
        n19632), .B2(n19218), .ZN(n19220) );
  OAI211_X1 U22137 ( .C1(n19561), .C2(n19254), .A(n19221), .B(n19220), .ZN(
        P2_U3055) );
  INV_X1 U22138 ( .A(n19222), .ZN(n19224) );
  NOR2_X1 U22139 ( .A1(n19223), .A2(n19271), .ZN(n19249) );
  NOR3_X1 U22140 ( .A1(n19224), .A2(n19249), .A3(n19528), .ZN(n19229) );
  INV_X1 U22141 ( .A(n19230), .ZN(n19225) );
  AOI21_X1 U22142 ( .B1(n19794), .B2(n19225), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19226) );
  NOR2_X1 U22143 ( .A1(n19229), .A2(n19226), .ZN(n19250) );
  AOI22_X1 U22144 ( .A1(n19250), .A2(n19574), .B1(n19249), .B2(n19573), .ZN(
        n19234) );
  INV_X1 U22145 ( .A(n19227), .ZN(n19350) );
  NAND2_X1 U22146 ( .A1(n19350), .A2(n19228), .ZN(n19231) );
  AOI21_X1 U22147 ( .B1(n19231), .B2(n19230), .A(n19229), .ZN(n19232) );
  OAI211_X1 U22148 ( .C1(n19249), .C2(n19794), .A(n19232), .B(n19533), .ZN(
        n19251) );
  AOI22_X1 U22149 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19251), .B1(
        n19241), .B2(n19576), .ZN(n19233) );
  OAI211_X1 U22150 ( .C1(n19537), .C2(n19244), .A(n19234), .B(n19233), .ZN(
        P2_U3056) );
  AOI22_X1 U22151 ( .A1(n19250), .A2(n19637), .B1(n14064), .B2(n19249), .ZN(
        n19236) );
  AOI22_X1 U22152 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19251), .B1(
        n19241), .B2(n19638), .ZN(n19235) );
  OAI211_X1 U22153 ( .C1(n19540), .C2(n19244), .A(n19236), .B(n19235), .ZN(
        P2_U3057) );
  AOI22_X1 U22154 ( .A1(n19250), .A2(n19644), .B1(n19249), .B2(n19643), .ZN(
        n19238) );
  AOI22_X1 U22155 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19251), .B1(
        n19241), .B2(n19645), .ZN(n19237) );
  OAI211_X1 U22156 ( .C1(n19543), .C2(n19244), .A(n19238), .B(n19237), .ZN(
        P2_U3058) );
  AOI22_X1 U22157 ( .A1(n19250), .A2(n19650), .B1(n19649), .B2(n19249), .ZN(
        n19240) );
  AOI22_X1 U22158 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19251), .B1(
        n19241), .B2(n19651), .ZN(n19239) );
  OAI211_X1 U22159 ( .C1(n19546), .C2(n19244), .A(n19240), .B(n19239), .ZN(
        P2_U3059) );
  AOI22_X1 U22160 ( .A1(n19250), .A2(n19656), .B1(n19249), .B2(n19655), .ZN(
        n19243) );
  AOI22_X1 U22161 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19251), .B1(
        n19241), .B2(n19658), .ZN(n19242) );
  OAI211_X1 U22162 ( .C1(n19592), .C2(n19244), .A(n19243), .B(n19242), .ZN(
        P2_U3060) );
  AOI22_X1 U22163 ( .A1(n19250), .A2(n19594), .B1(n19249), .B2(n19593), .ZN(
        n19246) );
  AOI22_X1 U22164 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19251), .B1(
        n19267), .B2(n19595), .ZN(n19245) );
  OAI211_X1 U22165 ( .C1(n19598), .C2(n19254), .A(n19246), .B(n19245), .ZN(
        P2_U3061) );
  AOI22_X1 U22166 ( .A1(n19250), .A2(n19664), .B1(n19663), .B2(n19249), .ZN(
        n19248) );
  AOI22_X1 U22167 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19251), .B1(
        n19267), .B2(n19668), .ZN(n19247) );
  OAI211_X1 U22168 ( .C1(n19516), .C2(n19254), .A(n19248), .B(n19247), .ZN(
        P2_U3062) );
  INV_X1 U22169 ( .A(n19629), .ZN(n19610) );
  AOI22_X1 U22170 ( .A1(n19250), .A2(n19632), .B1(n19627), .B2(n19249), .ZN(
        n19253) );
  AOI22_X1 U22171 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19251), .B1(
        n19267), .B2(n19630), .ZN(n19252) );
  OAI211_X1 U22172 ( .C1(n19610), .C2(n19254), .A(n19253), .B(n19252), .ZN(
        P2_U3063) );
  AOI22_X1 U22173 ( .A1(n19266), .A2(n19637), .B1(n14064), .B2(n19265), .ZN(
        n19256) );
  AOI22_X1 U22174 ( .A1(n19303), .A2(n19639), .B1(n19267), .B2(n19638), .ZN(
        n19255) );
  OAI211_X1 U22175 ( .C1(n19270), .C2(n12612), .A(n19256), .B(n19255), .ZN(
        P2_U3065) );
  AOI22_X1 U22176 ( .A1(n19266), .A2(n19644), .B1(n19643), .B2(n19265), .ZN(
        n19258) );
  AOI22_X1 U22177 ( .A1(n19303), .A2(n19646), .B1(n19267), .B2(n19645), .ZN(
        n19257) );
  OAI211_X1 U22178 ( .C1(n19270), .C2(n12598), .A(n19258), .B(n19257), .ZN(
        P2_U3066) );
  AOI22_X1 U22179 ( .A1(n19266), .A2(n19650), .B1(n19649), .B2(n19265), .ZN(
        n19260) );
  AOI22_X1 U22180 ( .A1(n19303), .A2(n19652), .B1(n19267), .B2(n19651), .ZN(
        n19259) );
  OAI211_X1 U22181 ( .C1(n19270), .C2(n12585), .A(n19260), .B(n19259), .ZN(
        P2_U3067) );
  AOI22_X1 U22182 ( .A1(n19266), .A2(n19656), .B1(n19655), .B2(n19265), .ZN(
        n19262) );
  AOI22_X1 U22183 ( .A1(n19267), .A2(n19658), .B1(n19303), .B2(n19657), .ZN(
        n19261) );
  OAI211_X1 U22184 ( .C1(n19270), .C2(n12572), .A(n19262), .B(n19261), .ZN(
        P2_U3068) );
  AOI22_X1 U22185 ( .A1(n19266), .A2(n19594), .B1(n19593), .B2(n19265), .ZN(
        n19264) );
  AOI22_X1 U22186 ( .A1(n19303), .A2(n19595), .B1(n19267), .B2(n19549), .ZN(
        n19263) );
  OAI211_X1 U22187 ( .C1(n19270), .C2(n12559), .A(n19264), .B(n19263), .ZN(
        P2_U3069) );
  AOI22_X1 U22188 ( .A1(n19266), .A2(n19632), .B1(n19627), .B2(n19265), .ZN(
        n19269) );
  AOI22_X1 U22189 ( .A1(n19303), .A2(n19630), .B1(n19267), .B2(n19629), .ZN(
        n19268) );
  OAI211_X1 U22190 ( .C1(n19270), .C2(n12667), .A(n19269), .B(n19268), .ZN(
        P2_U3071) );
  INV_X1 U22191 ( .A(n19487), .ZN(n19762) );
  AOI21_X1 U22192 ( .B1(n19350), .B2(n19762), .A(n19771), .ZN(n19275) );
  NOR2_X1 U22193 ( .A1(n19793), .A2(n19271), .ZN(n19279) );
  AND2_X1 U22194 ( .A1(n19490), .A2(n19272), .ZN(n19302) );
  INV_X1 U22195 ( .A(n19302), .ZN(n19276) );
  AOI21_X1 U22196 ( .B1(n19277), .B2(n19276), .A(n19528), .ZN(n19273) );
  AOI22_X1 U22197 ( .A1(n19575), .A2(n19343), .B1(n19573), .B2(n19302), .ZN(
        n19282) );
  INV_X1 U22198 ( .A(n19275), .ZN(n19280) );
  OAI211_X1 U22199 ( .C1(n19277), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19276), 
        .B(n19771), .ZN(n19278) );
  OAI211_X1 U22200 ( .C1(n19280), .C2(n19279), .A(n19533), .B(n19278), .ZN(
        n19304) );
  AOI22_X1 U22201 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19304), .B1(
        n19303), .B2(n19576), .ZN(n19281) );
  OAI211_X1 U22202 ( .C1(n19308), .C2(n19283), .A(n19282), .B(n19281), .ZN(
        P2_U3072) );
  AOI22_X1 U22203 ( .A1(n19639), .A2(n19343), .B1(n14064), .B2(n19302), .ZN(
        n19285) );
  AOI22_X1 U22204 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19304), .B1(
        n19303), .B2(n19638), .ZN(n19284) );
  OAI211_X1 U22205 ( .C1(n19308), .C2(n19286), .A(n19285), .B(n19284), .ZN(
        P2_U3073) );
  AOI22_X1 U22206 ( .A1(n19645), .A2(n19303), .B1(n19643), .B2(n19302), .ZN(
        n19288) );
  AOI22_X1 U22207 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19304), .B1(
        n19343), .B2(n19646), .ZN(n19287) );
  OAI211_X1 U22208 ( .C1(n19308), .C2(n19289), .A(n19288), .B(n19287), .ZN(
        P2_U3074) );
  AOI22_X1 U22209 ( .A1(n19652), .A2(n19343), .B1(n19649), .B2(n19302), .ZN(
        n19291) );
  AOI22_X1 U22210 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19304), .B1(
        n19303), .B2(n19651), .ZN(n19290) );
  OAI211_X1 U22211 ( .C1(n19308), .C2(n19292), .A(n19291), .B(n19290), .ZN(
        P2_U3075) );
  AOI22_X1 U22212 ( .A1(n19657), .A2(n19343), .B1(n19655), .B2(n19302), .ZN(
        n19294) );
  AOI22_X1 U22213 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19304), .B1(
        n19303), .B2(n19658), .ZN(n19293) );
  OAI211_X1 U22214 ( .C1(n19308), .C2(n19295), .A(n19294), .B(n19293), .ZN(
        P2_U3076) );
  AOI22_X1 U22215 ( .A1(n19595), .A2(n19343), .B1(n19593), .B2(n19302), .ZN(
        n19297) );
  AOI22_X1 U22216 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19304), .B1(
        n19303), .B2(n19549), .ZN(n19296) );
  OAI211_X1 U22217 ( .C1(n19308), .C2(n19298), .A(n19297), .B(n19296), .ZN(
        P2_U3077) );
  AOI22_X1 U22218 ( .A1(n19666), .A2(n19303), .B1(n19663), .B2(n19302), .ZN(
        n19300) );
  AOI22_X1 U22219 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19304), .B1(
        n19343), .B2(n19668), .ZN(n19299) );
  OAI211_X1 U22220 ( .C1(n19308), .C2(n19301), .A(n19300), .B(n19299), .ZN(
        P2_U3078) );
  INV_X1 U22221 ( .A(n19632), .ZN(n19307) );
  AOI22_X1 U22222 ( .A1(n19629), .A2(n19303), .B1(n19627), .B2(n19302), .ZN(
        n19306) );
  AOI22_X1 U22223 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19304), .B1(
        n19343), .B2(n19630), .ZN(n19305) );
  OAI211_X1 U22224 ( .C1(n19308), .C2(n19307), .A(n19306), .B(n19305), .ZN(
        P2_U3079) );
  NAND3_X1 U22225 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n19775), .A3(
        n19793), .ZN(n19356) );
  NOR2_X1 U22226 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19356), .ZN(
        n19341) );
  NOR3_X1 U22227 ( .A1(n19309), .A2(n19341), .A3(n19528), .ZN(n19320) );
  INV_X1 U22228 ( .A(n19320), .ZN(n19316) );
  INV_X1 U22229 ( .A(n19341), .ZN(n19314) );
  NOR2_X1 U22230 ( .A1(n19311), .A2(n19310), .ZN(n19529) );
  NAND2_X1 U22231 ( .A1(n19529), .A2(n19775), .ZN(n19317) );
  OAI21_X1 U22232 ( .B1(n19343), .B2(n19373), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19313) );
  AOI22_X1 U22233 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19314), .B1(n19317), 
        .B2(n19313), .ZN(n19315) );
  INV_X1 U22234 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n19323) );
  INV_X1 U22235 ( .A(n19317), .ZN(n19318) );
  AOI21_X1 U22236 ( .B1(n19794), .B2(n19318), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19319) );
  NOR2_X1 U22237 ( .A1(n19320), .A2(n19319), .ZN(n19342) );
  AOI22_X1 U22238 ( .A1(n19342), .A2(n19574), .B1(n19341), .B2(n19573), .ZN(
        n19322) );
  AOI22_X1 U22239 ( .A1(n19343), .A2(n19576), .B1(n19373), .B2(n19575), .ZN(
        n19321) );
  OAI211_X1 U22240 ( .C1(n19347), .C2(n19323), .A(n19322), .B(n19321), .ZN(
        P2_U3080) );
  INV_X1 U22241 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n19326) );
  AOI22_X1 U22242 ( .A1(n19342), .A2(n19637), .B1(n14064), .B2(n19341), .ZN(
        n19325) );
  AOI22_X1 U22243 ( .A1(n19373), .A2(n19639), .B1(n19343), .B2(n19638), .ZN(
        n19324) );
  OAI211_X1 U22244 ( .C1(n19347), .C2(n19326), .A(n19325), .B(n19324), .ZN(
        P2_U3081) );
  INV_X1 U22245 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n19329) );
  AOI22_X1 U22246 ( .A1(n19342), .A2(n19644), .B1(n19341), .B2(n19643), .ZN(
        n19328) );
  AOI22_X1 U22247 ( .A1(n19373), .A2(n19646), .B1(n19343), .B2(n19645), .ZN(
        n19327) );
  OAI211_X1 U22248 ( .C1(n19347), .C2(n19329), .A(n19328), .B(n19327), .ZN(
        P2_U3082) );
  INV_X1 U22249 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n19332) );
  AOI22_X1 U22250 ( .A1(n19342), .A2(n19650), .B1(n19649), .B2(n19341), .ZN(
        n19331) );
  AOI22_X1 U22251 ( .A1(n19373), .A2(n19652), .B1(n19343), .B2(n19651), .ZN(
        n19330) );
  OAI211_X1 U22252 ( .C1(n19347), .C2(n19332), .A(n19331), .B(n19330), .ZN(
        P2_U3083) );
  INV_X1 U22253 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n19335) );
  AOI22_X1 U22254 ( .A1(n19342), .A2(n19656), .B1(n19341), .B2(n19655), .ZN(
        n19334) );
  AOI22_X1 U22255 ( .A1(n19343), .A2(n19658), .B1(n19373), .B2(n19657), .ZN(
        n19333) );
  OAI211_X1 U22256 ( .C1(n19347), .C2(n19335), .A(n19334), .B(n19333), .ZN(
        P2_U3084) );
  INV_X1 U22257 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n19338) );
  AOI22_X1 U22258 ( .A1(n19342), .A2(n19594), .B1(n19341), .B2(n19593), .ZN(
        n19337) );
  AOI22_X1 U22259 ( .A1(n19373), .A2(n19595), .B1(n19343), .B2(n19549), .ZN(
        n19336) );
  OAI211_X1 U22260 ( .C1(n19347), .C2(n19338), .A(n19337), .B(n19336), .ZN(
        P2_U3085) );
  AOI22_X1 U22261 ( .A1(n19342), .A2(n19664), .B1(n19663), .B2(n19341), .ZN(
        n19340) );
  AOI22_X1 U22262 ( .A1(n19373), .A2(n19668), .B1(n19343), .B2(n19666), .ZN(
        n19339) );
  OAI211_X1 U22263 ( .C1(n19347), .C2(n12632), .A(n19340), .B(n19339), .ZN(
        P2_U3086) );
  INV_X1 U22264 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n19346) );
  AOI22_X1 U22265 ( .A1(n19342), .A2(n19632), .B1(n19627), .B2(n19341), .ZN(
        n19345) );
  AOI22_X1 U22266 ( .A1(n19373), .A2(n19630), .B1(n19343), .B2(n19629), .ZN(
        n19344) );
  OAI211_X1 U22267 ( .C1(n19347), .C2(n19346), .A(n19345), .B(n19344), .ZN(
        P2_U3087) );
  NOR2_X1 U22268 ( .A1(n19802), .A2(n19356), .ZN(n19384) );
  AOI22_X1 U22269 ( .A1(n19576), .A2(n19373), .B1(n19573), .B2(n19384), .ZN(
        n19359) );
  INV_X1 U22270 ( .A(n19562), .ZN(n19349) );
  AOI21_X1 U22271 ( .B1(n19350), .B2(n19349), .A(n19771), .ZN(n19354) );
  INV_X1 U22272 ( .A(n19351), .ZN(n19352) );
  NOR2_X1 U22273 ( .A1(n19352), .A2(n19384), .ZN(n19355) );
  AOI22_X1 U22274 ( .A1(n19354), .A2(n19356), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n19355), .ZN(n19353) );
  OAI211_X1 U22275 ( .C1(n19384), .C2(n19794), .A(n19353), .B(n19533), .ZN(
        n19375) );
  INV_X1 U22276 ( .A(n19354), .ZN(n19357) );
  OAI22_X1 U22277 ( .A1(n19357), .A2(n19356), .B1(n19355), .B2(n19528), .ZN(
        n19374) );
  AOI22_X1 U22278 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19375), .B1(
        n19574), .B2(n19374), .ZN(n19358) );
  OAI211_X1 U22279 ( .C1(n19537), .C2(n19407), .A(n19359), .B(n19358), .ZN(
        P2_U3088) );
  AOI22_X1 U22280 ( .A1(n19639), .A2(n19399), .B1(n14064), .B2(n19384), .ZN(
        n19361) );
  AOI22_X1 U22281 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19375), .B1(
        n19637), .B2(n19374), .ZN(n19360) );
  OAI211_X1 U22282 ( .C1(n19583), .C2(n19366), .A(n19361), .B(n19360), .ZN(
        P2_U3089) );
  AOI22_X1 U22283 ( .A1(n19646), .A2(n19399), .B1(n19643), .B2(n19384), .ZN(
        n19363) );
  AOI22_X1 U22284 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19375), .B1(
        n19644), .B2(n19374), .ZN(n19362) );
  OAI211_X1 U22285 ( .C1(n19586), .C2(n19366), .A(n19363), .B(n19362), .ZN(
        P2_U3090) );
  AOI22_X1 U22286 ( .A1(n19652), .A2(n19399), .B1(n19649), .B2(n19384), .ZN(
        n19365) );
  AOI22_X1 U22287 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19375), .B1(
        n19650), .B2(n19374), .ZN(n19364) );
  OAI211_X1 U22288 ( .C1(n19589), .C2(n19366), .A(n19365), .B(n19364), .ZN(
        P2_U3091) );
  AOI22_X1 U22289 ( .A1(n19658), .A2(n19373), .B1(n19655), .B2(n19384), .ZN(
        n19368) );
  AOI22_X1 U22290 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19375), .B1(
        n19656), .B2(n19374), .ZN(n19367) );
  OAI211_X1 U22291 ( .C1(n19592), .C2(n19407), .A(n19368), .B(n19367), .ZN(
        P2_U3092) );
  AOI22_X1 U22292 ( .A1(n19549), .A2(n19373), .B1(n19593), .B2(n19384), .ZN(
        n19370) );
  AOI22_X1 U22293 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19375), .B1(
        n19594), .B2(n19374), .ZN(n19369) );
  OAI211_X1 U22294 ( .C1(n19552), .C2(n19407), .A(n19370), .B(n19369), .ZN(
        P2_U3093) );
  AOI22_X1 U22295 ( .A1(n19666), .A2(n19373), .B1(n19663), .B2(n19384), .ZN(
        n19372) );
  AOI22_X1 U22296 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19375), .B1(
        n19664), .B2(n19374), .ZN(n19371) );
  OAI211_X1 U22297 ( .C1(n19603), .C2(n19407), .A(n19372), .B(n19371), .ZN(
        P2_U3094) );
  AOI22_X1 U22298 ( .A1(n19629), .A2(n19373), .B1(n19627), .B2(n19384), .ZN(
        n19377) );
  AOI22_X1 U22299 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19375), .B1(
        n19632), .B2(n19374), .ZN(n19376) );
  OAI211_X1 U22300 ( .C1(n19561), .C2(n19407), .A(n19377), .B(n19376), .ZN(
        P2_U3095) );
  NOR2_X1 U22301 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19378), .ZN(
        n19402) );
  NOR2_X1 U22302 ( .A1(n19384), .A2(n19402), .ZN(n19379) );
  OR2_X1 U22303 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19379), .ZN(n19381) );
  NOR3_X1 U22304 ( .A1(n10271), .A2(n19402), .A3(n19528), .ZN(n19385) );
  AOI21_X1 U22305 ( .B1(n19528), .B2(n19381), .A(n19385), .ZN(n19403) );
  AOI22_X1 U22306 ( .A1(n19403), .A2(n19574), .B1(n19402), .B2(n19573), .ZN(
        n19388) );
  AOI21_X1 U22307 ( .B1(n19407), .B2(n19419), .A(n19382), .ZN(n19383) );
  AOI221_X1 U22308 ( .B1(n19794), .B2(n19384), .C1(n19794), .C2(n19383), .A(
        n19402), .ZN(n19386) );
  AOI22_X1 U22309 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19404), .B1(
        n19399), .B2(n19576), .ZN(n19387) );
  OAI211_X1 U22310 ( .C1(n19537), .C2(n19419), .A(n19388), .B(n19387), .ZN(
        P2_U3096) );
  AOI22_X1 U22311 ( .A1(n19403), .A2(n19637), .B1(n14064), .B2(n19402), .ZN(
        n19390) );
  AOI22_X1 U22312 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19404), .B1(
        n19421), .B2(n19639), .ZN(n19389) );
  OAI211_X1 U22313 ( .C1(n19583), .C2(n19407), .A(n19390), .B(n19389), .ZN(
        P2_U3097) );
  AOI22_X1 U22314 ( .A1(n19403), .A2(n19644), .B1(n19402), .B2(n19643), .ZN(
        n19392) );
  AOI22_X1 U22315 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19404), .B1(
        n19399), .B2(n19645), .ZN(n19391) );
  OAI211_X1 U22316 ( .C1(n19543), .C2(n19419), .A(n19392), .B(n19391), .ZN(
        P2_U3098) );
  AOI22_X1 U22317 ( .A1(n19403), .A2(n19650), .B1(n19649), .B2(n19402), .ZN(
        n19394) );
  AOI22_X1 U22318 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19404), .B1(
        n19421), .B2(n19652), .ZN(n19393) );
  OAI211_X1 U22319 ( .C1(n19589), .C2(n19407), .A(n19394), .B(n19393), .ZN(
        P2_U3099) );
  AOI22_X1 U22320 ( .A1(n19403), .A2(n19656), .B1(n19402), .B2(n19655), .ZN(
        n19396) );
  AOI22_X1 U22321 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19404), .B1(
        n19399), .B2(n19658), .ZN(n19395) );
  OAI211_X1 U22322 ( .C1(n19592), .C2(n19419), .A(n19396), .B(n19395), .ZN(
        P2_U3100) );
  AOI22_X1 U22323 ( .A1(n19403), .A2(n19594), .B1(n19402), .B2(n19593), .ZN(
        n19398) );
  AOI22_X1 U22324 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19404), .B1(
        n19421), .B2(n19595), .ZN(n19397) );
  OAI211_X1 U22325 ( .C1(n19598), .C2(n19407), .A(n19398), .B(n19397), .ZN(
        P2_U3101) );
  AOI22_X1 U22326 ( .A1(n19403), .A2(n19664), .B1(n19663), .B2(n19402), .ZN(
        n19401) );
  AOI22_X1 U22327 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19404), .B1(
        n19399), .B2(n19666), .ZN(n19400) );
  OAI211_X1 U22328 ( .C1(n19603), .C2(n19419), .A(n19401), .B(n19400), .ZN(
        P2_U3102) );
  AOI22_X1 U22329 ( .A1(n19403), .A2(n19632), .B1(n19627), .B2(n19402), .ZN(
        n19406) );
  AOI22_X1 U22330 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19404), .B1(
        n19421), .B2(n19630), .ZN(n19405) );
  OAI211_X1 U22331 ( .C1(n19610), .C2(n19407), .A(n19406), .B(n19405), .ZN(
        P2_U3103) );
  AOI22_X1 U22332 ( .A1(n19420), .A2(n19637), .B1(n19432), .B2(n14064), .ZN(
        n19409) );
  AOI22_X1 U22333 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19416), .B1(
        n19421), .B2(n19638), .ZN(n19408) );
  OAI211_X1 U22334 ( .C1(n19540), .C2(n19458), .A(n19409), .B(n19408), .ZN(
        P2_U3105) );
  INV_X1 U22335 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n20816) );
  AOI22_X1 U22336 ( .A1(n19420), .A2(n19644), .B1(n19432), .B2(n19643), .ZN(
        n19411) );
  AOI22_X1 U22337 ( .A1(n19444), .A2(n19646), .B1(n19421), .B2(n19645), .ZN(
        n19410) );
  OAI211_X1 U22338 ( .C1(n19425), .C2(n20816), .A(n19411), .B(n19410), .ZN(
        P2_U3106) );
  AOI22_X1 U22339 ( .A1(n19420), .A2(n19650), .B1(n19432), .B2(n19649), .ZN(
        n19413) );
  AOI22_X1 U22340 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19416), .B1(
        n19421), .B2(n19651), .ZN(n19412) );
  OAI211_X1 U22341 ( .C1(n19546), .C2(n19458), .A(n19413), .B(n19412), .ZN(
        P2_U3107) );
  AOI22_X1 U22342 ( .A1(n19420), .A2(n19656), .B1(n19432), .B2(n19655), .ZN(
        n19415) );
  AOI22_X1 U22343 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19416), .B1(
        n19421), .B2(n19658), .ZN(n19414) );
  OAI211_X1 U22344 ( .C1(n19592), .C2(n19458), .A(n19415), .B(n19414), .ZN(
        P2_U3108) );
  AOI22_X1 U22345 ( .A1(n19420), .A2(n19664), .B1(n19432), .B2(n19663), .ZN(
        n19418) );
  AOI22_X1 U22346 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19416), .B1(
        n19444), .B2(n19668), .ZN(n19417) );
  OAI211_X1 U22347 ( .C1(n19516), .C2(n19419), .A(n19418), .B(n19417), .ZN(
        P2_U3110) );
  INV_X1 U22348 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n19424) );
  AOI22_X1 U22349 ( .A1(n19420), .A2(n19632), .B1(n19432), .B2(n19627), .ZN(
        n19423) );
  AOI22_X1 U22350 ( .A1(n19444), .A2(n19630), .B1(n19421), .B2(n19629), .ZN(
        n19422) );
  OAI211_X1 U22351 ( .C1(n19425), .C2(n19424), .A(n19423), .B(n19422), .ZN(
        P2_U3111) );
  NOR2_X1 U22352 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19426), .ZN(
        n19452) );
  AOI22_X1 U22353 ( .A1(n19576), .A2(n19444), .B1(n19573), .B2(n19452), .ZN(
        n19437) );
  NAND2_X1 U22354 ( .A1(n19458), .A2(n19447), .ZN(n19427) );
  AOI21_X1 U22355 ( .B1(n19427), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19771), 
        .ZN(n19431) );
  AOI21_X1 U22356 ( .B1(n19433), .B2(n19794), .A(n19764), .ZN(n19428) );
  AOI21_X1 U22357 ( .B1(n19431), .B2(n19429), .A(n19428), .ZN(n19430) );
  OAI21_X1 U22358 ( .B1(n19452), .B2(n19430), .A(n19533), .ZN(n19455) );
  OAI21_X1 U22359 ( .B1(n19432), .B2(n19452), .A(n19431), .ZN(n19435) );
  OAI21_X1 U22360 ( .B1(n19433), .B2(n19452), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19434) );
  NAND2_X1 U22361 ( .A1(n19435), .A2(n19434), .ZN(n19454) );
  AOI22_X1 U22362 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19455), .B1(
        n19574), .B2(n19454), .ZN(n19436) );
  OAI211_X1 U22363 ( .C1(n19537), .C2(n19447), .A(n19437), .B(n19436), .ZN(
        P2_U3112) );
  AOI22_X1 U22364 ( .A1(n19639), .A2(n19453), .B1(n14064), .B2(n19452), .ZN(
        n19439) );
  AOI22_X1 U22365 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19455), .B1(
        n19454), .B2(n19637), .ZN(n19438) );
  OAI211_X1 U22366 ( .C1(n19583), .C2(n19458), .A(n19439), .B(n19438), .ZN(
        P2_U3113) );
  AOI22_X1 U22367 ( .A1(n19646), .A2(n19453), .B1(n19643), .B2(n19452), .ZN(
        n19441) );
  AOI22_X1 U22368 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19455), .B1(
        n19454), .B2(n19644), .ZN(n19440) );
  OAI211_X1 U22369 ( .C1(n19586), .C2(n19458), .A(n19441), .B(n19440), .ZN(
        P2_U3114) );
  AOI22_X1 U22370 ( .A1(n19652), .A2(n19453), .B1(n19649), .B2(n19452), .ZN(
        n19443) );
  AOI22_X1 U22371 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19455), .B1(
        n19454), .B2(n19650), .ZN(n19442) );
  OAI211_X1 U22372 ( .C1(n19589), .C2(n19458), .A(n19443), .B(n19442), .ZN(
        P2_U3115) );
  AOI22_X1 U22373 ( .A1(n19658), .A2(n19444), .B1(n19655), .B2(n19452), .ZN(
        n19446) );
  AOI22_X1 U22374 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19455), .B1(
        n19454), .B2(n19656), .ZN(n19445) );
  OAI211_X1 U22375 ( .C1(n19592), .C2(n19447), .A(n19446), .B(n19445), .ZN(
        P2_U3116) );
  AOI22_X1 U22376 ( .A1(n19595), .A2(n19453), .B1(n19593), .B2(n19452), .ZN(
        n19449) );
  AOI22_X1 U22377 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19455), .B1(
        n19454), .B2(n19594), .ZN(n19448) );
  OAI211_X1 U22378 ( .C1(n19598), .C2(n19458), .A(n19449), .B(n19448), .ZN(
        P2_U3117) );
  AOI22_X1 U22379 ( .A1(n19668), .A2(n19453), .B1(n19663), .B2(n19452), .ZN(
        n19451) );
  AOI22_X1 U22380 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19455), .B1(
        n19454), .B2(n19664), .ZN(n19450) );
  OAI211_X1 U22381 ( .C1(n19516), .C2(n19458), .A(n19451), .B(n19450), .ZN(
        P2_U3118) );
  AOI22_X1 U22382 ( .A1(n19630), .A2(n19453), .B1(n19627), .B2(n19452), .ZN(
        n19457) );
  AOI22_X1 U22383 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19455), .B1(
        n19454), .B2(n19632), .ZN(n19456) );
  OAI211_X1 U22384 ( .C1(n19610), .C2(n19458), .A(n19457), .B(n19456), .ZN(
        P2_U3119) );
  NOR2_X1 U22385 ( .A1(n19459), .A2(n19489), .ZN(n19481) );
  OAI21_X1 U22386 ( .B1(n19460), .B2(n19481), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19461) );
  OAI21_X1 U22387 ( .B1(n19489), .B2(n19462), .A(n19461), .ZN(n19482) );
  AOI22_X1 U22388 ( .A1(n19482), .A2(n19574), .B1(n19481), .B2(n19573), .ZN(
        n19468) );
  AOI221_X1 U22389 ( .B1(n19508), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19483), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19463), .ZN(n19464) );
  AOI211_X1 U22390 ( .C1(P2_STATE2_REG_2__SCAN_IN), .C2(n19465), .A(
        P2_STATE2_REG_3__SCAN_IN), .B(n19464), .ZN(n19466) );
  OAI21_X1 U22391 ( .B1(n19466), .B2(n19481), .A(n19533), .ZN(n19484) );
  AOI22_X1 U22392 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19484), .B1(
        n19483), .B2(n19576), .ZN(n19467) );
  OAI211_X1 U22393 ( .C1(n19537), .C2(n19522), .A(n19468), .B(n19467), .ZN(
        P2_U3128) );
  AOI22_X1 U22394 ( .A1(n19482), .A2(n19637), .B1(n14064), .B2(n19481), .ZN(
        n19470) );
  AOI22_X1 U22395 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19484), .B1(
        n19483), .B2(n19638), .ZN(n19469) );
  OAI211_X1 U22396 ( .C1(n19540), .C2(n19522), .A(n19470), .B(n19469), .ZN(
        P2_U3129) );
  AOI22_X1 U22397 ( .A1(n19482), .A2(n19644), .B1(n19481), .B2(n19643), .ZN(
        n19472) );
  AOI22_X1 U22398 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19484), .B1(
        n19483), .B2(n19645), .ZN(n19471) );
  OAI211_X1 U22399 ( .C1(n19543), .C2(n19522), .A(n19472), .B(n19471), .ZN(
        P2_U3130) );
  AOI22_X1 U22400 ( .A1(n19482), .A2(n19650), .B1(n19649), .B2(n19481), .ZN(
        n19474) );
  AOI22_X1 U22401 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19484), .B1(
        n19483), .B2(n19651), .ZN(n19473) );
  OAI211_X1 U22402 ( .C1(n19546), .C2(n19522), .A(n19474), .B(n19473), .ZN(
        P2_U3131) );
  AOI22_X1 U22403 ( .A1(n19482), .A2(n19656), .B1(n19481), .B2(n19655), .ZN(
        n19476) );
  AOI22_X1 U22404 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19484), .B1(
        n19483), .B2(n19658), .ZN(n19475) );
  OAI211_X1 U22405 ( .C1(n19592), .C2(n19522), .A(n19476), .B(n19475), .ZN(
        P2_U3132) );
  AOI22_X1 U22406 ( .A1(n19482), .A2(n19594), .B1(n19481), .B2(n19593), .ZN(
        n19478) );
  AOI22_X1 U22407 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19484), .B1(
        n19483), .B2(n19549), .ZN(n19477) );
  OAI211_X1 U22408 ( .C1(n19552), .C2(n19522), .A(n19478), .B(n19477), .ZN(
        P2_U3133) );
  AOI22_X1 U22409 ( .A1(n19482), .A2(n19664), .B1(n19663), .B2(n19481), .ZN(
        n19480) );
  AOI22_X1 U22410 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19484), .B1(
        n19483), .B2(n19666), .ZN(n19479) );
  OAI211_X1 U22411 ( .C1(n19603), .C2(n19522), .A(n19480), .B(n19479), .ZN(
        P2_U3134) );
  AOI22_X1 U22412 ( .A1(n19482), .A2(n19632), .B1(n19627), .B2(n19481), .ZN(
        n19486) );
  AOI22_X1 U22413 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19484), .B1(
        n19483), .B2(n19629), .ZN(n19485) );
  OAI211_X1 U22414 ( .C1(n19561), .C2(n19522), .A(n19486), .B(n19485), .ZN(
        P2_U3135) );
  NOR2_X2 U22415 ( .A1(n19488), .A2(n19487), .ZN(n19557) );
  INV_X1 U22416 ( .A(n19557), .ZN(n19511) );
  INV_X1 U22417 ( .A(n19489), .ZN(n19492) );
  AND2_X1 U22418 ( .A1(n19490), .A2(n19492), .ZN(n19517) );
  NOR3_X1 U22419 ( .A1(n19491), .A2(n19517), .A3(n19528), .ZN(n19496) );
  NAND2_X1 U22420 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19492), .ZN(
        n19497) );
  INV_X1 U22421 ( .A(n19497), .ZN(n19493) );
  AOI21_X1 U22422 ( .B1(n19794), .B2(n19493), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19494) );
  NOR2_X1 U22423 ( .A1(n19496), .A2(n19494), .ZN(n19518) );
  AOI22_X1 U22424 ( .A1(n19518), .A2(n19574), .B1(n19517), .B2(n19573), .ZN(
        n19501) );
  NAND2_X1 U22425 ( .A1(n19495), .A2(n19762), .ZN(n19498) );
  AOI21_X1 U22426 ( .B1(n19498), .B2(n19497), .A(n19496), .ZN(n19499) );
  OAI211_X1 U22427 ( .C1(n19517), .C2(n19794), .A(n19499), .B(n19533), .ZN(
        n19519) );
  AOI22_X1 U22428 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19519), .B1(
        n19508), .B2(n19576), .ZN(n19500) );
  OAI211_X1 U22429 ( .C1(n19537), .C2(n19511), .A(n19501), .B(n19500), .ZN(
        P2_U3136) );
  AOI22_X1 U22430 ( .A1(n19518), .A2(n19637), .B1(n14064), .B2(n19517), .ZN(
        n19503) );
  AOI22_X1 U22431 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19519), .B1(
        n19508), .B2(n19638), .ZN(n19502) );
  OAI211_X1 U22432 ( .C1(n19540), .C2(n19511), .A(n19503), .B(n19502), .ZN(
        P2_U3137) );
  AOI22_X1 U22433 ( .A1(n19518), .A2(n19644), .B1(n19517), .B2(n19643), .ZN(
        n19505) );
  AOI22_X1 U22434 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19519), .B1(
        n19557), .B2(n19646), .ZN(n19504) );
  OAI211_X1 U22435 ( .C1(n19586), .C2(n19522), .A(n19505), .B(n19504), .ZN(
        P2_U3138) );
  AOI22_X1 U22436 ( .A1(n19518), .A2(n19650), .B1(n19649), .B2(n19517), .ZN(
        n19507) );
  AOI22_X1 U22437 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19519), .B1(
        n19557), .B2(n19652), .ZN(n19506) );
  OAI211_X1 U22438 ( .C1(n19589), .C2(n19522), .A(n19507), .B(n19506), .ZN(
        P2_U3139) );
  AOI22_X1 U22439 ( .A1(n19518), .A2(n19656), .B1(n19517), .B2(n19655), .ZN(
        n19510) );
  AOI22_X1 U22440 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19519), .B1(
        n19508), .B2(n19658), .ZN(n19509) );
  OAI211_X1 U22441 ( .C1(n19592), .C2(n19511), .A(n19510), .B(n19509), .ZN(
        P2_U3140) );
  AOI22_X1 U22442 ( .A1(n19518), .A2(n19594), .B1(n19517), .B2(n19593), .ZN(
        n19513) );
  AOI22_X1 U22443 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19519), .B1(
        n19557), .B2(n19595), .ZN(n19512) );
  OAI211_X1 U22444 ( .C1(n19598), .C2(n19522), .A(n19513), .B(n19512), .ZN(
        P2_U3141) );
  AOI22_X1 U22445 ( .A1(n19518), .A2(n19664), .B1(n19663), .B2(n19517), .ZN(
        n19515) );
  AOI22_X1 U22446 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19519), .B1(
        n19557), .B2(n19668), .ZN(n19514) );
  OAI211_X1 U22447 ( .C1(n19516), .C2(n19522), .A(n19515), .B(n19514), .ZN(
        P2_U3142) );
  AOI22_X1 U22448 ( .A1(n19518), .A2(n19632), .B1(n19627), .B2(n19517), .ZN(
        n19521) );
  AOI22_X1 U22449 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19519), .B1(
        n19557), .B2(n19630), .ZN(n19520) );
  OAI211_X1 U22450 ( .C1(n19610), .C2(n19522), .A(n19521), .B(n19520), .ZN(
        P2_U3143) );
  NOR2_X1 U22451 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19572), .ZN(
        n19555) );
  NOR2_X1 U22452 ( .A1(n19524), .A2(n19555), .ZN(n19530) );
  INV_X1 U22453 ( .A(n19525), .ZN(n19527) );
  INV_X1 U22454 ( .A(n19529), .ZN(n19526) );
  OAI22_X1 U22455 ( .A1(n19530), .A2(n19528), .B1(n19527), .B2(n19526), .ZN(
        n19556) );
  AOI22_X1 U22456 ( .A1(n19556), .A2(n19574), .B1(n19555), .B2(n19573), .ZN(
        n19536) );
  OAI21_X1 U22457 ( .B1(n19599), .B2(n19557), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19532) );
  NAND2_X1 U22458 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19529), .ZN(
        n19531) );
  AOI22_X1 U22459 ( .A1(n19532), .A2(n19531), .B1(P2_STATE2_REG_2__SCAN_IN), 
        .B2(n19530), .ZN(n19534) );
  OAI211_X1 U22460 ( .C1(n19555), .C2(n19794), .A(n19534), .B(n19533), .ZN(
        n19558) );
  AOI22_X1 U22461 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19558), .B1(
        n19557), .B2(n19576), .ZN(n19535) );
  OAI211_X1 U22462 ( .C1(n19537), .C2(n19609), .A(n19536), .B(n19535), .ZN(
        P2_U3144) );
  AOI22_X1 U22463 ( .A1(n19556), .A2(n19637), .B1(n14064), .B2(n19555), .ZN(
        n19539) );
  AOI22_X1 U22464 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19558), .B1(
        n19557), .B2(n19638), .ZN(n19538) );
  OAI211_X1 U22465 ( .C1(n19540), .C2(n19609), .A(n19539), .B(n19538), .ZN(
        P2_U3145) );
  AOI22_X1 U22466 ( .A1(n19556), .A2(n19644), .B1(n19555), .B2(n19643), .ZN(
        n19542) );
  AOI22_X1 U22467 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19558), .B1(
        n19557), .B2(n19645), .ZN(n19541) );
  OAI211_X1 U22468 ( .C1(n19543), .C2(n19609), .A(n19542), .B(n19541), .ZN(
        P2_U3146) );
  AOI22_X1 U22469 ( .A1(n19556), .A2(n19650), .B1(n19649), .B2(n19555), .ZN(
        n19545) );
  AOI22_X1 U22470 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19558), .B1(
        n19557), .B2(n19651), .ZN(n19544) );
  OAI211_X1 U22471 ( .C1(n19546), .C2(n19609), .A(n19545), .B(n19544), .ZN(
        P2_U3147) );
  AOI22_X1 U22472 ( .A1(n19556), .A2(n19656), .B1(n19555), .B2(n19655), .ZN(
        n19548) );
  AOI22_X1 U22473 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19558), .B1(
        n19557), .B2(n19658), .ZN(n19547) );
  OAI211_X1 U22474 ( .C1(n19592), .C2(n19609), .A(n19548), .B(n19547), .ZN(
        P2_U3148) );
  AOI22_X1 U22475 ( .A1(n19556), .A2(n19594), .B1(n19555), .B2(n19593), .ZN(
        n19551) );
  AOI22_X1 U22476 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19558), .B1(
        n19557), .B2(n19549), .ZN(n19550) );
  OAI211_X1 U22477 ( .C1(n19552), .C2(n19609), .A(n19551), .B(n19550), .ZN(
        P2_U3149) );
  AOI22_X1 U22478 ( .A1(n19556), .A2(n19664), .B1(n19663), .B2(n19555), .ZN(
        n19554) );
  AOI22_X1 U22479 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19558), .B1(
        n19557), .B2(n19666), .ZN(n19553) );
  OAI211_X1 U22480 ( .C1(n19603), .C2(n19609), .A(n19554), .B(n19553), .ZN(
        P2_U3150) );
  AOI22_X1 U22481 ( .A1(n19556), .A2(n19632), .B1(n19627), .B2(n19555), .ZN(
        n19560) );
  AOI22_X1 U22482 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19558), .B1(
        n19557), .B2(n19629), .ZN(n19559) );
  OAI211_X1 U22483 ( .C1(n19561), .C2(n19609), .A(n19560), .B(n19559), .ZN(
        P2_U3151) );
  OAI21_X1 U22484 ( .B1(n19563), .B2(n19562), .A(n19572), .ZN(n19569) );
  OR2_X1 U22485 ( .A1(n19564), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19567) );
  NOR2_X1 U22486 ( .A1(n19764), .A2(n19604), .ZN(n19566) );
  AOI21_X1 U22487 ( .B1(n19567), .B2(n19566), .A(n19565), .ZN(n19568) );
  INV_X1 U22488 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n19579) );
  OAI21_X1 U22489 ( .B1(n19570), .B2(n19604), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19571) );
  OAI21_X1 U22490 ( .B1(n19572), .B2(n19771), .A(n19571), .ZN(n19605) );
  AOI22_X1 U22491 ( .A1(n19605), .A2(n19574), .B1(n19604), .B2(n19573), .ZN(
        n19578) );
  AOI22_X1 U22492 ( .A1(n19599), .A2(n19576), .B1(n19628), .B2(n19575), .ZN(
        n19577) );
  OAI211_X1 U22493 ( .C1(n19580), .C2(n19579), .A(n19578), .B(n19577), .ZN(
        P2_U3152) );
  AOI22_X1 U22494 ( .A1(n19605), .A2(n19637), .B1(n14064), .B2(n19604), .ZN(
        n19582) );
  AOI22_X1 U22495 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19606), .B1(
        n19628), .B2(n19639), .ZN(n19581) );
  OAI211_X1 U22496 ( .C1(n19583), .C2(n19609), .A(n19582), .B(n19581), .ZN(
        P2_U3153) );
  AOI22_X1 U22497 ( .A1(n19605), .A2(n19644), .B1(n19604), .B2(n19643), .ZN(
        n19585) );
  AOI22_X1 U22498 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19606), .B1(
        n19628), .B2(n19646), .ZN(n19584) );
  OAI211_X1 U22499 ( .C1(n19586), .C2(n19609), .A(n19585), .B(n19584), .ZN(
        P2_U3154) );
  AOI22_X1 U22500 ( .A1(n19605), .A2(n19650), .B1(n19649), .B2(n19604), .ZN(
        n19588) );
  AOI22_X1 U22501 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19606), .B1(
        n19628), .B2(n19652), .ZN(n19587) );
  OAI211_X1 U22502 ( .C1(n19589), .C2(n19609), .A(n19588), .B(n19587), .ZN(
        P2_U3155) );
  AOI22_X1 U22503 ( .A1(n19605), .A2(n19656), .B1(n19604), .B2(n19655), .ZN(
        n19591) );
  AOI22_X1 U22504 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19606), .B1(
        n19599), .B2(n19658), .ZN(n19590) );
  OAI211_X1 U22505 ( .C1(n19592), .C2(n19602), .A(n19591), .B(n19590), .ZN(
        P2_U3156) );
  AOI22_X1 U22506 ( .A1(n19605), .A2(n19594), .B1(n19604), .B2(n19593), .ZN(
        n19597) );
  AOI22_X1 U22507 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19606), .B1(
        n19628), .B2(n19595), .ZN(n19596) );
  OAI211_X1 U22508 ( .C1(n19598), .C2(n19609), .A(n19597), .B(n19596), .ZN(
        P2_U3157) );
  AOI22_X1 U22509 ( .A1(n19605), .A2(n19664), .B1(n19663), .B2(n19604), .ZN(
        n19601) );
  AOI22_X1 U22510 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19606), .B1(
        n19599), .B2(n19666), .ZN(n19600) );
  OAI211_X1 U22511 ( .C1(n19603), .C2(n19602), .A(n19601), .B(n19600), .ZN(
        P2_U3158) );
  AOI22_X1 U22512 ( .A1(n19605), .A2(n19632), .B1(n19627), .B2(n19604), .ZN(
        n19608) );
  AOI22_X1 U22513 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19606), .B1(
        n19628), .B2(n19630), .ZN(n19607) );
  OAI211_X1 U22514 ( .C1(n19610), .C2(n19609), .A(n19608), .B(n19607), .ZN(
        P2_U3159) );
  INV_X1 U22515 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n19613) );
  AOI22_X1 U22516 ( .A1(n19638), .A2(n19628), .B1(n14064), .B2(n19626), .ZN(
        n19612) );
  AOI22_X1 U22517 ( .A1(n19637), .A2(n19631), .B1(n19667), .B2(n19639), .ZN(
        n19611) );
  OAI211_X1 U22518 ( .C1(n19636), .C2(n19613), .A(n19612), .B(n19611), .ZN(
        P2_U3161) );
  INV_X1 U22519 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n19616) );
  AOI22_X1 U22520 ( .A1(n19646), .A2(n19667), .B1(n19643), .B2(n19626), .ZN(
        n19615) );
  AOI22_X1 U22521 ( .A1(n19644), .A2(n19631), .B1(n19628), .B2(n19645), .ZN(
        n19614) );
  OAI211_X1 U22522 ( .C1(n19636), .C2(n19616), .A(n19615), .B(n19614), .ZN(
        P2_U3162) );
  INV_X1 U22523 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n19619) );
  AOI22_X1 U22524 ( .A1(n19652), .A2(n19667), .B1(n19649), .B2(n19626), .ZN(
        n19618) );
  AOI22_X1 U22525 ( .A1(n19650), .A2(n19631), .B1(n19628), .B2(n19651), .ZN(
        n19617) );
  OAI211_X1 U22526 ( .C1(n19636), .C2(n19619), .A(n19618), .B(n19617), .ZN(
        P2_U3163) );
  INV_X1 U22527 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n19622) );
  AOI22_X1 U22528 ( .A1(n19658), .A2(n19628), .B1(n19655), .B2(n19626), .ZN(
        n19621) );
  AOI22_X1 U22529 ( .A1(n19656), .A2(n19631), .B1(n19667), .B2(n19657), .ZN(
        n19620) );
  OAI211_X1 U22530 ( .C1(n19636), .C2(n19622), .A(n19621), .B(n19620), .ZN(
        P2_U3164) );
  INV_X1 U22531 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n19625) );
  AOI22_X1 U22532 ( .A1(n19668), .A2(n19667), .B1(n19663), .B2(n19626), .ZN(
        n19624) );
  AOI22_X1 U22533 ( .A1(n19664), .A2(n19631), .B1(n19628), .B2(n19666), .ZN(
        n19623) );
  OAI211_X1 U22534 ( .C1(n19636), .C2(n19625), .A(n19624), .B(n19623), .ZN(
        P2_U3166) );
  INV_X1 U22535 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n19635) );
  AOI22_X1 U22536 ( .A1(n19629), .A2(n19628), .B1(n19627), .B2(n19626), .ZN(
        n19634) );
  AOI22_X1 U22537 ( .A1(n19632), .A2(n19631), .B1(n19667), .B2(n19630), .ZN(
        n19633) );
  OAI211_X1 U22538 ( .C1(n19636), .C2(n19635), .A(n19634), .B(n19633), .ZN(
        P2_U3167) );
  INV_X1 U22539 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n19642) );
  AOI22_X1 U22540 ( .A1(n19665), .A2(n19637), .B1(n14064), .B2(n19662), .ZN(
        n19641) );
  AOI22_X1 U22541 ( .A1(n19669), .A2(n19639), .B1(n19667), .B2(n19638), .ZN(
        n19640) );
  OAI211_X1 U22542 ( .C1(n19672), .C2(n19642), .A(n19641), .B(n19640), .ZN(
        P2_U3169) );
  AOI22_X1 U22543 ( .A1(n19665), .A2(n19644), .B1(n19662), .B2(n19643), .ZN(
        n19648) );
  AOI22_X1 U22544 ( .A1(n19669), .A2(n19646), .B1(n19667), .B2(n19645), .ZN(
        n19647) );
  OAI211_X1 U22545 ( .C1(n19672), .C2(n10321), .A(n19648), .B(n19647), .ZN(
        P2_U3170) );
  AOI22_X1 U22546 ( .A1(n19665), .A2(n19650), .B1(n19649), .B2(n19662), .ZN(
        n19654) );
  AOI22_X1 U22547 ( .A1(n19669), .A2(n19652), .B1(n19667), .B2(n19651), .ZN(
        n19653) );
  OAI211_X1 U22548 ( .C1(n19672), .C2(n10353), .A(n19654), .B(n19653), .ZN(
        P2_U3171) );
  INV_X1 U22549 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n19661) );
  AOI22_X1 U22550 ( .A1(n19665), .A2(n19656), .B1(n19662), .B2(n19655), .ZN(
        n19660) );
  AOI22_X1 U22551 ( .A1(n19667), .A2(n19658), .B1(n19669), .B2(n19657), .ZN(
        n19659) );
  OAI211_X1 U22552 ( .C1(n19672), .C2(n19661), .A(n19660), .B(n19659), .ZN(
        P2_U3172) );
  AOI22_X1 U22553 ( .A1(n19665), .A2(n19664), .B1(n19663), .B2(n19662), .ZN(
        n19671) );
  AOI22_X1 U22554 ( .A1(n19669), .A2(n19668), .B1(n19667), .B2(n19666), .ZN(
        n19670) );
  OAI211_X1 U22555 ( .C1(n19672), .C2(n10412), .A(n19671), .B(n19670), .ZN(
        P2_U3174) );
  NOR2_X1 U22556 ( .A1(n19695), .A2(n19822), .ZN(n19674) );
  AOI21_X1 U22557 ( .B1(n19763), .B2(n19674), .A(n19673), .ZN(n19678) );
  OAI211_X1 U22558 ( .C1(n19679), .C2(n19675), .A(n19695), .B(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19676) );
  OAI211_X1 U22559 ( .C1(n19679), .C2(n19678), .A(n19677), .B(n19676), .ZN(
        P2_U3177) );
  AND2_X1 U22560 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19680), .ZN(
        P2_U3179) );
  AND2_X1 U22561 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19680), .ZN(
        P2_U3180) );
  AND2_X1 U22562 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19680), .ZN(
        P2_U3181) );
  AND2_X1 U22563 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19680), .ZN(
        P2_U3182) );
  AND2_X1 U22564 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19680), .ZN(
        P2_U3183) );
  AND2_X1 U22565 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19680), .ZN(
        P2_U3184) );
  AND2_X1 U22566 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19680), .ZN(
        P2_U3185) );
  AND2_X1 U22567 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19680), .ZN(
        P2_U3186) );
  AND2_X1 U22568 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19680), .ZN(
        P2_U3187) );
  AND2_X1 U22569 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19680), .ZN(
        P2_U3188) );
  AND2_X1 U22570 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19680), .ZN(
        P2_U3189) );
  AND2_X1 U22571 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19680), .ZN(
        P2_U3190) );
  AND2_X1 U22572 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19680), .ZN(
        P2_U3191) );
  AND2_X1 U22573 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19680), .ZN(
        P2_U3192) );
  AND2_X1 U22574 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19680), .ZN(
        P2_U3193) );
  AND2_X1 U22575 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19680), .ZN(
        P2_U3194) );
  AND2_X1 U22576 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19680), .ZN(
        P2_U3195) );
  AND2_X1 U22577 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19680), .ZN(
        P2_U3196) );
  AND2_X1 U22578 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19680), .ZN(
        P2_U3197) );
  AND2_X1 U22579 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19680), .ZN(
        P2_U3198) );
  AND2_X1 U22580 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19680), .ZN(
        P2_U3199) );
  AND2_X1 U22581 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19680), .ZN(
        P2_U3200) );
  AND2_X1 U22582 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19680), .ZN(P2_U3201) );
  AND2_X1 U22583 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19680), .ZN(P2_U3202) );
  AND2_X1 U22584 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19680), .ZN(P2_U3203) );
  AND2_X1 U22585 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19680), .ZN(P2_U3204) );
  AND2_X1 U22586 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19680), .ZN(P2_U3205) );
  AND2_X1 U22587 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19680), .ZN(P2_U3206) );
  AND2_X1 U22588 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19680), .ZN(P2_U3207) );
  AND2_X1 U22589 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19680), .ZN(P2_U3208) );
  NOR2_X1 U22590 ( .A1(n19692), .A2(n19825), .ZN(n19690) );
  INV_X1 U22591 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19836) );
  OR3_X1 U22592 ( .A1(n19690), .A2(n19836), .A3(n19681), .ZN(n19683) );
  AOI211_X1 U22593 ( .C1(n20670), .C2(P2_REQUESTPENDING_REG_SCAN_IN), .A(
        n19691), .B(n19837), .ZN(n19682) );
  INV_X1 U22594 ( .A(NA), .ZN(n20676) );
  NOR2_X1 U22595 ( .A1(n20676), .A2(n19685), .ZN(n19697) );
  AOI211_X1 U22596 ( .C1(n19700), .C2(n19683), .A(n19682), .B(n19697), .ZN(
        n19684) );
  INV_X1 U22597 ( .A(n19684), .ZN(P2_U3209) );
  AOI21_X1 U22598 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20670), .A(n19700), 
        .ZN(n19693) );
  NOR2_X1 U22599 ( .A1(n19836), .A2(n19693), .ZN(n19686) );
  AOI21_X1 U22600 ( .B1(n19686), .B2(n19685), .A(n19690), .ZN(n19688) );
  OAI211_X1 U22601 ( .C1(n20670), .C2(n19689), .A(n19688), .B(n19687), .ZN(
        P2_U3210) );
  AOI22_X1 U22602 ( .A1(n19691), .A2(n19836), .B1(n19690), .B2(n20676), .ZN(
        n19699) );
  OAI21_X1 U22603 ( .B1(P2_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .ZN(n19698) );
  NOR2_X1 U22604 ( .A1(n19692), .A2(n19700), .ZN(n19694) );
  AOI21_X1 U22605 ( .B1(n19695), .B2(n19694), .A(n19693), .ZN(n19696) );
  OAI22_X1 U22606 ( .A1(n19699), .A2(n19698), .B1(n19697), .B2(n19696), .ZN(
        P2_U3211) );
  OAI222_X1 U22607 ( .A1(n19751), .A2(n19702), .B1(n19701), .B2(n19837), .C1(
        n19704), .C2(n19750), .ZN(P2_U3212) );
  OAI222_X1 U22608 ( .A1(n19751), .A2(n19704), .B1(n19703), .B2(n19837), .C1(
        n13701), .C2(n19750), .ZN(P2_U3213) );
  OAI222_X1 U22609 ( .A1(n19751), .A2(n13701), .B1(n19705), .B2(n19837), .C1(
        n19706), .C2(n19750), .ZN(P2_U3214) );
  INV_X1 U22610 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n19708) );
  OAI222_X1 U22611 ( .A1(n19750), .A2(n19708), .B1(n19707), .B2(n19837), .C1(
        n19706), .C2(n19751), .ZN(P2_U3215) );
  OAI222_X1 U22612 ( .A1(n19750), .A2(n19710), .B1(n19709), .B2(n19837), .C1(
        n19708), .C2(n19751), .ZN(P2_U3216) );
  OAI222_X1 U22613 ( .A1(n19750), .A2(n19712), .B1(n19711), .B2(n19837), .C1(
        n19710), .C2(n19751), .ZN(P2_U3217) );
  INV_X1 U22614 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19714) );
  OAI222_X1 U22615 ( .A1(n19750), .A2(n19714), .B1(n19713), .B2(n19837), .C1(
        n19712), .C2(n19751), .ZN(P2_U3218) );
  INV_X1 U22616 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19716) );
  OAI222_X1 U22617 ( .A1(n19750), .A2(n19716), .B1(n19715), .B2(n19837), .C1(
        n19714), .C2(n19751), .ZN(P2_U3219) );
  OAI222_X1 U22618 ( .A1(n19750), .A2(n19718), .B1(n19717), .B2(n19837), .C1(
        n19716), .C2(n19751), .ZN(P2_U3220) );
  OAI222_X1 U22619 ( .A1(n19750), .A2(n15631), .B1(n19719), .B2(n19837), .C1(
        n19718), .C2(n19751), .ZN(P2_U3221) );
  OAI222_X1 U22620 ( .A1(n19750), .A2(n11008), .B1(n19720), .B2(n19837), .C1(
        n15631), .C2(n19751), .ZN(P2_U3222) );
  OAI222_X1 U22621 ( .A1(n19750), .A2(n11011), .B1(n19721), .B2(n19837), .C1(
        n11008), .C2(n19751), .ZN(P2_U3223) );
  OAI222_X1 U22622 ( .A1(n19750), .A2(n10788), .B1(n19722), .B2(n19837), .C1(
        n11011), .C2(n19751), .ZN(P2_U3224) );
  INV_X1 U22623 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19724) );
  OAI222_X1 U22624 ( .A1(n19750), .A2(n19724), .B1(n19723), .B2(n19837), .C1(
        n10788), .C2(n19751), .ZN(P2_U3225) );
  OAI222_X1 U22625 ( .A1(n19750), .A2(n15350), .B1(n19725), .B2(n19837), .C1(
        n19724), .C2(n19751), .ZN(P2_U3226) );
  OAI222_X1 U22626 ( .A1(n19750), .A2(n19727), .B1(n19726), .B2(n19837), .C1(
        n15350), .C2(n19751), .ZN(P2_U3227) );
  OAI222_X1 U22627 ( .A1(n19750), .A2(n19729), .B1(n19728), .B2(n19837), .C1(
        n19727), .C2(n19751), .ZN(P2_U3228) );
  OAI222_X1 U22628 ( .A1(n19750), .A2(n15090), .B1(n19730), .B2(n19837), .C1(
        n19729), .C2(n19751), .ZN(P2_U3229) );
  OAI222_X1 U22629 ( .A1(n19750), .A2(n11122), .B1(n19731), .B2(n19837), .C1(
        n15090), .C2(n19751), .ZN(P2_U3230) );
  OAI222_X1 U22630 ( .A1(n19750), .A2(n19733), .B1(n19732), .B2(n19837), .C1(
        n11122), .C2(n19751), .ZN(P2_U3231) );
  OAI222_X1 U22631 ( .A1(n19750), .A2(n19735), .B1(n19734), .B2(n19837), .C1(
        n19733), .C2(n19751), .ZN(P2_U3232) );
  OAI222_X1 U22632 ( .A1(n19750), .A2(n19737), .B1(n19736), .B2(n19837), .C1(
        n19735), .C2(n19751), .ZN(P2_U3233) );
  OAI222_X1 U22633 ( .A1(n19750), .A2(n19739), .B1(n19738), .B2(n19837), .C1(
        n19737), .C2(n19751), .ZN(P2_U3234) );
  INV_X1 U22634 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19741) );
  OAI222_X1 U22635 ( .A1(n19750), .A2(n19741), .B1(n19740), .B2(n19837), .C1(
        n19739), .C2(n19751), .ZN(P2_U3235) );
  INV_X1 U22636 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19743) );
  OAI222_X1 U22637 ( .A1(n19750), .A2(n19743), .B1(n19742), .B2(n19837), .C1(
        n19741), .C2(n19751), .ZN(P2_U3236) );
  OAI222_X1 U22638 ( .A1(n19750), .A2(n19746), .B1(n19744), .B2(n19837), .C1(
        n19743), .C2(n19751), .ZN(P2_U3237) );
  OAI222_X1 U22639 ( .A1(n19751), .A2(n19746), .B1(n19745), .B2(n19837), .C1(
        n12467), .C2(n19750), .ZN(P2_U3238) );
  OAI222_X1 U22640 ( .A1(n19750), .A2(n19748), .B1(n19747), .B2(n19837), .C1(
        n12467), .C2(n19751), .ZN(P2_U3239) );
  OAI222_X1 U22641 ( .A1(n19750), .A2(n19752), .B1(n19749), .B2(n19837), .C1(
        n19748), .C2(n19751), .ZN(P2_U3240) );
  OAI222_X1 U22642 ( .A1(n19750), .A2(n19754), .B1(n19753), .B2(n19837), .C1(
        n19752), .C2(n19751), .ZN(P2_U3241) );
  OAI22_X1 U22643 ( .A1(n19838), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19837), .ZN(n19755) );
  INV_X1 U22644 ( .A(n19755), .ZN(P2_U3585) );
  MUX2_X1 U22645 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .B(P2_BE_N_REG_2__SCAN_IN), .S(n19838), .Z(P2_U3586) );
  OAI22_X1 U22646 ( .A1(n19838), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19837), .ZN(n19756) );
  INV_X1 U22647 ( .A(n19756), .ZN(P2_U3587) );
  OAI22_X1 U22648 ( .A1(n19838), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19837), .ZN(n19757) );
  INV_X1 U22649 ( .A(n19757), .ZN(P2_U3588) );
  OAI21_X1 U22650 ( .B1(n19761), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19759), 
        .ZN(n19758) );
  INV_X1 U22651 ( .A(n19758), .ZN(P2_U3591) );
  OAI21_X1 U22652 ( .B1(n19761), .B2(n19760), .A(n19759), .ZN(P2_U3592) );
  INV_X1 U22653 ( .A(n19800), .ZN(n19803) );
  AND2_X1 U22654 ( .A1(n19764), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19789) );
  NAND2_X1 U22655 ( .A1(n19762), .A2(n19789), .ZN(n19778) );
  NAND2_X1 U22656 ( .A1(n19787), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19765) );
  AOI21_X1 U22657 ( .B1(n19765), .B2(n19764), .A(n19763), .ZN(n19776) );
  NAND2_X1 U22658 ( .A1(n19778), .A2(n19776), .ZN(n19767) );
  NAND2_X1 U22659 ( .A1(n19767), .A2(n19766), .ZN(n19770) );
  NAND2_X1 U22660 ( .A1(n19768), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19769) );
  OAI211_X1 U22661 ( .C1(n19772), .C2(n19771), .A(n19770), .B(n19769), .ZN(
        n19773) );
  INV_X1 U22662 ( .A(n19773), .ZN(n19774) );
  AOI22_X1 U22663 ( .A1(n19803), .A2(n19775), .B1(n19774), .B2(n19800), .ZN(
        P2_U3602) );
  INV_X1 U22664 ( .A(n19776), .ZN(n19781) );
  NOR2_X1 U22665 ( .A1(n19777), .A2(n19794), .ZN(n19780) );
  INV_X1 U22666 ( .A(n19778), .ZN(n19779) );
  AOI211_X1 U22667 ( .C1(n19782), .C2(n19781), .A(n19780), .B(n19779), .ZN(
        n19783) );
  AOI22_X1 U22668 ( .A1(n19803), .A2(n19784), .B1(n19783), .B2(n19800), .ZN(
        P2_U3603) );
  INV_X1 U22669 ( .A(n19785), .ZN(n19795) );
  AND2_X1 U22670 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19786) );
  NOR2_X1 U22671 ( .A1(n19795), .A2(n19786), .ZN(n19788) );
  MUX2_X1 U22672 ( .A(n19789), .B(n19788), .S(n19787), .Z(n19790) );
  AOI21_X1 U22673 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19791), .A(n19790), 
        .ZN(n19792) );
  AOI22_X1 U22674 ( .A1(n19803), .A2(n19793), .B1(n19792), .B2(n19800), .ZN(
        P2_U3604) );
  OAI22_X1 U22675 ( .A1(n19796), .A2(n19795), .B1(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n19794), .ZN(n19797) );
  AOI21_X1 U22676 ( .B1(n19799), .B2(n19798), .A(n19797), .ZN(n19801) );
  AOI22_X1 U22677 ( .A1(n19803), .A2(n19802), .B1(n19801), .B2(n19800), .ZN(
        P2_U3605) );
  INV_X1 U22678 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19804) );
  AOI22_X1 U22679 ( .A1(n19837), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19804), 
        .B2(n19838), .ZN(P2_U3608) );
  INV_X1 U22680 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n19817) );
  INV_X1 U22681 ( .A(n19805), .ZN(n19816) );
  AOI21_X1 U22682 ( .B1(n19808), .B2(n19807), .A(n19806), .ZN(n19812) );
  NOR3_X1 U22683 ( .A1(n19810), .A2(n10069), .A3(n19809), .ZN(n19811) );
  NOR2_X1 U22684 ( .A1(n19812), .A2(n19811), .ZN(n19815) );
  NOR2_X1 U22685 ( .A1(n19816), .A2(n19813), .ZN(n19814) );
  AOI22_X1 U22686 ( .A1(n19817), .A2(n19816), .B1(n19815), .B2(n19814), .ZN(
        P2_U3609) );
  AOI21_X1 U22687 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19818), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19820) );
  AOI211_X1 U22688 ( .C1(n19821), .C2(n19825), .A(n19820), .B(n19819), .ZN(
        n19835) );
  NOR4_X1 U22689 ( .A1(n19828), .A2(n19829), .A3(n19823), .A4(n19822), .ZN(
        n19827) );
  AOI21_X1 U22690 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19825), .A(n19824), 
        .ZN(n19826) );
  NOR2_X1 U22691 ( .A1(n19827), .A2(n19826), .ZN(n19834) );
  NAND2_X1 U22692 ( .A1(n19828), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19831) );
  AND3_X1 U22693 ( .A1(n19831), .A2(n19830), .A3(n19829), .ZN(n19832) );
  NOR2_X1 U22694 ( .A1(n19835), .A2(n19832), .ZN(n19833) );
  AOI22_X1 U22695 ( .A1(n19836), .A2(n19835), .B1(n19834), .B2(n19833), .ZN(
        P2_U3610) );
  OAI22_X1 U22696 ( .A1(n19838), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19837), .ZN(n19839) );
  INV_X1 U22697 ( .A(n19839), .ZN(P2_U3611) );
  NAND2_X1 U22698 ( .A1(n19840), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .ZN(n19842)
         );
  NAND3_X1 U22699 ( .A1(n19842), .A2(n19847), .A3(n19841), .ZN(P1_U2801) );
  OAI21_X1 U22700 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(n20663), .A(
        P1_STATE_REG_0__SCAN_IN), .ZN(n20679) );
  INV_X2 U22701 ( .A(n20750), .ZN(n20748) );
  OAI21_X1 U22702 ( .B1(n20679), .B2(P1_ADS_N_REG_SCAN_IN), .A(n20748), .ZN(
        n19843) );
  INV_X1 U22703 ( .A(n19843), .ZN(P1_U2802) );
  OAI21_X1 U22704 ( .B1(n19845), .B2(n19844), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19846) );
  OAI21_X1 U22705 ( .B1(n19847), .B2(n20756), .A(n19846), .ZN(P1_U2803) );
  NOR2_X1 U22706 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19849) );
  OAI21_X1 U22707 ( .B1(n19849), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20748), .ZN(
        n19848) );
  OAI21_X1 U22708 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20748), .A(n19848), 
        .ZN(P1_U2804) );
  NAND2_X1 U22709 ( .A1(n20679), .A2(n20748), .ZN(n20662) );
  INV_X1 U22710 ( .A(n20662), .ZN(n20726) );
  OAI21_X1 U22711 ( .B1(BS16), .B2(n19849), .A(n20726), .ZN(n20724) );
  OAI21_X1 U22712 ( .B1(n20726), .B2(n20753), .A(n20724), .ZN(P1_U2805) );
  OAI21_X1 U22713 ( .B1(n19852), .B2(n19851), .A(n19850), .ZN(P1_U2806) );
  NOR4_X1 U22714 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_21__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19856) );
  NOR4_X1 U22715 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19855) );
  NOR4_X1 U22716 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19854) );
  NOR4_X1 U22717 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19853) );
  NAND4_X1 U22718 ( .A1(n19856), .A2(n19855), .A3(n19854), .A4(n19853), .ZN(
        n19862) );
  NOR4_X1 U22719 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_3__SCAN_IN), .A3(P1_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_6__SCAN_IN), .ZN(n19860) );
  AOI211_X1 U22720 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_19__SCAN_IN), .B(
        P1_DATAWIDTH_REG_4__SCAN_IN), .ZN(n19859) );
  NOR4_X1 U22721 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19858) );
  NOR4_X1 U22722 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_8__SCAN_IN), .A3(P1_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19857) );
  NAND4_X1 U22723 ( .A1(n19860), .A2(n19859), .A3(n19858), .A4(n19857), .ZN(
        n19861) );
  NOR2_X1 U22724 ( .A1(n19862), .A2(n19861), .ZN(n20747) );
  INV_X1 U22725 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19864) );
  NOR3_X1 U22726 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19865) );
  OAI21_X1 U22727 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19865), .A(n20747), .ZN(
        n19863) );
  OAI21_X1 U22728 ( .B1(n20747), .B2(n19864), .A(n19863), .ZN(P1_U2807) );
  INV_X1 U22729 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20725) );
  AOI21_X1 U22730 ( .B1(n20740), .B2(n20725), .A(n19865), .ZN(n19867) );
  INV_X1 U22731 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19866) );
  INV_X1 U22732 ( .A(n20747), .ZN(n20742) );
  AOI22_X1 U22733 ( .A1(n20747), .A2(n19867), .B1(n19866), .B2(n20742), .ZN(
        P1_U2808) );
  INV_X1 U22734 ( .A(n19868), .ZN(n19877) );
  NOR3_X1 U22735 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n19869), .A3(n19924), .ZN(
        n19876) );
  AOI21_X1 U22736 ( .B1(n19926), .B2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n19913), .ZN(n19870) );
  OAI21_X1 U22737 ( .B1(n19940), .B2(n19871), .A(n19870), .ZN(n19872) );
  AOI21_X1 U22738 ( .B1(n19938), .B2(P1_EBX_REG_9__SCAN_IN), .A(n19872), .ZN(
        n19873) );
  OAI21_X1 U22739 ( .B1(n19874), .B2(n19897), .A(n19873), .ZN(n19875) );
  AOI211_X1 U22740 ( .C1(n19877), .C2(n19904), .A(n19876), .B(n19875), .ZN(
        n19878) );
  OAI21_X1 U22741 ( .B1(n19880), .B2(n19879), .A(n19878), .ZN(P1_U2831) );
  NAND2_X1 U22742 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .ZN(n19882) );
  AOI21_X1 U22743 ( .B1(n19881), .B2(n19882), .A(n19919), .ZN(n19901) );
  INV_X1 U22744 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n19893) );
  OR3_X1 U22745 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19882), .A3(n19924), .ZN(
        n19891) );
  NAND2_X1 U22746 ( .A1(n19938), .A2(P1_EBX_REG_7__SCAN_IN), .ZN(n19884) );
  AOI21_X1 U22747 ( .B1(n19926), .B2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n19913), .ZN(n19883) );
  OAI211_X1 U22748 ( .C1(n19940), .C2(n19885), .A(n19884), .B(n19883), .ZN(
        n19886) );
  AOI21_X1 U22749 ( .B1(n19945), .B2(n19887), .A(n19886), .ZN(n19890) );
  NAND2_X1 U22750 ( .A1(n19888), .A2(n19904), .ZN(n19889) );
  AND3_X1 U22751 ( .A1(n19891), .A2(n19890), .A3(n19889), .ZN(n19892) );
  OAI21_X1 U22752 ( .B1(n19901), .B2(n19893), .A(n19892), .ZN(P1_U2833) );
  INV_X1 U22753 ( .A(n19894), .ZN(n19898) );
  OAI22_X1 U22754 ( .A1(n19898), .A2(n19897), .B1(n19896), .B2(n19895), .ZN(
        n19899) );
  AOI211_X1 U22755 ( .C1(n19926), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n19913), .B(n19899), .ZN(n19909) );
  INV_X1 U22756 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n19900) );
  NOR2_X1 U22757 ( .A1(n19900), .A2(n19924), .ZN(n19903) );
  INV_X1 U22758 ( .A(n19901), .ZN(n19902) );
  MUX2_X1 U22759 ( .A(n19903), .B(n19902), .S(P1_REIP_REG_6__SCAN_IN), .Z(
        n19907) );
  AND2_X1 U22760 ( .A1(n19905), .A2(n19904), .ZN(n19906) );
  NOR2_X1 U22761 ( .A1(n19907), .A2(n19906), .ZN(n19908) );
  OAI211_X1 U22762 ( .C1(n19910), .C2(n19940), .A(n19909), .B(n19908), .ZN(
        P1_U2834) );
  INV_X1 U22763 ( .A(n19911), .ZN(n19912) );
  NAND2_X1 U22764 ( .A1(n19945), .A2(n19912), .ZN(n19918) );
  NAND2_X1 U22765 ( .A1(n19938), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n19917) );
  AOI21_X1 U22766 ( .B1(n19927), .B2(n19914), .A(n19913), .ZN(n19916) );
  NAND2_X1 U22767 ( .A1(n19926), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n19915) );
  AND4_X1 U22768 ( .A1(n19918), .A2(n19917), .A3(n19916), .A4(n19915), .ZN(
        n19923) );
  INV_X1 U22769 ( .A(n19949), .ZN(n19920) );
  AOI22_X1 U22770 ( .A1(n19921), .A2(n19920), .B1(P1_REIP_REG_5__SCAN_IN), 
        .B2(n19919), .ZN(n19922) );
  OAI211_X1 U22771 ( .C1(P1_REIP_REG_5__SCAN_IN), .C2(n19924), .A(n19923), .B(
        n19922), .ZN(P1_U2835) );
  INV_X1 U22772 ( .A(n19925), .ZN(n19928) );
  AOI222_X1 U22773 ( .A1(n20735), .A2(n19943), .B1(n19928), .B2(n19927), .C1(
        n19926), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n19936) );
  AOI221_X1 U22774 ( .B1(P1_REIP_REG_3__SCAN_IN), .B2(P1_REIP_REG_2__SCAN_IN), 
        .C1(n20684), .C2(n20682), .A(n19929), .ZN(n19934) );
  AOI22_X1 U22775 ( .A1(n19930), .A2(n19945), .B1(n19938), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n19931) );
  OAI21_X1 U22776 ( .B1(n19932), .B2(n19949), .A(n19931), .ZN(n19933) );
  NOR2_X1 U22777 ( .A1(n19934), .A2(n19933), .ZN(n19935) );
  OAI211_X1 U22778 ( .C1(n19937), .C2(n20684), .A(n19936), .B(n19935), .ZN(
        P1_U2837) );
  AOI22_X1 U22779 ( .A1(n19939), .A2(P1_REIP_REG_0__SCAN_IN), .B1(n19938), 
        .B2(P1_EBX_REG_0__SCAN_IN), .ZN(n19948) );
  NAND2_X1 U22780 ( .A1(n19941), .A2(n19940), .ZN(n19946) );
  INV_X1 U22781 ( .A(n19942), .ZN(n19944) );
  AOI222_X1 U22782 ( .A1(n19946), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19945), .B2(n19944), .C1(n9621), .C2(n19943), .ZN(n19947) );
  OAI211_X1 U22783 ( .C1(n19949), .C2(n20097), .A(n19948), .B(n19947), .ZN(
        P1_U2840) );
  AOI22_X1 U22784 ( .A1(n20761), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n19962), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19951) );
  OAI21_X1 U22785 ( .B1(n13245), .B2(n19970), .A(n19951), .ZN(P1_U2921) );
  INV_X1 U22786 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20089) );
  AOI22_X1 U22787 ( .A1(n20761), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n19962), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19952) );
  OAI21_X1 U22788 ( .B1(n20089), .B2(n19970), .A(n19952), .ZN(P1_U2922) );
  INV_X1 U22789 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20083) );
  AOI22_X1 U22790 ( .A1(n20761), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n19962), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19953) );
  OAI21_X1 U22791 ( .B1(n20083), .B2(n19970), .A(n19953), .ZN(P1_U2923) );
  INV_X1 U22792 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n20079) );
  AOI22_X1 U22793 ( .A1(n20761), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n19962), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19954) );
  OAI21_X1 U22794 ( .B1(n20079), .B2(n19970), .A(n19954), .ZN(P1_U2924) );
  AOI22_X1 U22795 ( .A1(n20761), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n19962), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19955) );
  OAI21_X1 U22796 ( .B1(n14323), .B2(n19970), .A(n19955), .ZN(P1_U2925) );
  AOI22_X1 U22797 ( .A1(n20761), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n19962), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19956) );
  OAI21_X1 U22798 ( .B1(n14213), .B2(n19970), .A(n19956), .ZN(P1_U2926) );
  INV_X1 U22799 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n20069) );
  AOI22_X1 U22800 ( .A1(n20761), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n19962), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19957) );
  OAI21_X1 U22801 ( .B1(n20069), .B2(n19970), .A(n19957), .ZN(P1_U2927) );
  AOI22_X1 U22802 ( .A1(n20761), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n19962), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19958) );
  OAI21_X1 U22803 ( .B1(n14028), .B2(n19970), .A(n19958), .ZN(P1_U2928) );
  AOI22_X1 U22804 ( .A1(n19968), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n19962), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19959) );
  OAI21_X1 U22805 ( .B1(n11878), .B2(n19970), .A(n19959), .ZN(P1_U2929) );
  AOI22_X1 U22806 ( .A1(n19968), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n19962), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19960) );
  OAI21_X1 U22807 ( .B1(n11870), .B2(n19970), .A(n19960), .ZN(P1_U2930) );
  AOI22_X1 U22808 ( .A1(n19968), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n19962), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19961) );
  OAI21_X1 U22809 ( .B1(n13728), .B2(n19970), .A(n19961), .ZN(P1_U2931) );
  AOI22_X1 U22810 ( .A1(n19968), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n19962), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19963) );
  OAI21_X1 U22811 ( .B1(n20053), .B2(n19970), .A(n19963), .ZN(P1_U2932) );
  AOI22_X1 U22812 ( .A1(n19968), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n19967), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19964) );
  OAI21_X1 U22813 ( .B1(n20049), .B2(n19970), .A(n19964), .ZN(P1_U2933) );
  AOI22_X1 U22814 ( .A1(n19968), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n19967), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19965) );
  OAI21_X1 U22815 ( .B1(n20866), .B2(n19970), .A(n19965), .ZN(P1_U2934) );
  AOI22_X1 U22816 ( .A1(n19968), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n19967), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19966) );
  OAI21_X1 U22817 ( .B1(n20042), .B2(n19970), .A(n19966), .ZN(P1_U2935) );
  AOI22_X1 U22818 ( .A1(n19968), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n19967), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19969) );
  OAI21_X1 U22819 ( .B1(n20038), .B2(n19970), .A(n19969), .ZN(P1_U2936) );
  INV_X1 U22820 ( .A(n20112), .ZN(n19972) );
  NAND2_X1 U22821 ( .A1(n20031), .A2(n19972), .ZN(n20036) );
  INV_X2 U22822 ( .A(n19973), .ZN(n20084) );
  NAND2_X1 U22823 ( .A1(n20084), .A2(P1_UWORD_REG_0__SCAN_IN), .ZN(n19974) );
  AND2_X1 U22824 ( .A1(n20036), .A2(n19974), .ZN(n19975) );
  OAI21_X1 U22825 ( .B1(n19976), .B2(n20088), .A(n19975), .ZN(P1_U2937) );
  INV_X1 U22826 ( .A(n20121), .ZN(n19977) );
  NAND2_X1 U22827 ( .A1(n20031), .A2(n19977), .ZN(n20040) );
  NAND2_X1 U22828 ( .A1(n20084), .A2(P1_UWORD_REG_1__SCAN_IN), .ZN(n19978) );
  AND2_X1 U22829 ( .A1(n20040), .A2(n19978), .ZN(n19979) );
  OAI21_X1 U22830 ( .B1(n14816), .B2(n20088), .A(n19979), .ZN(P1_U2938) );
  INV_X1 U22831 ( .A(n20124), .ZN(n19980) );
  NAND2_X1 U22832 ( .A1(n20031), .A2(n19980), .ZN(n20044) );
  NAND2_X1 U22833 ( .A1(n20084), .A2(P1_UWORD_REG_2__SCAN_IN), .ZN(n19981) );
  AND2_X1 U22834 ( .A1(n20044), .A2(n19981), .ZN(n19982) );
  OAI21_X1 U22835 ( .B1(n19983), .B2(n20088), .A(n19982), .ZN(P1_U2939) );
  INV_X1 U22836 ( .A(n20128), .ZN(n19984) );
  NAND2_X1 U22837 ( .A1(n20031), .A2(n19984), .ZN(n20047) );
  NAND2_X1 U22838 ( .A1(n20084), .A2(P1_UWORD_REG_3__SCAN_IN), .ZN(n19985) );
  AND2_X1 U22839 ( .A1(n20047), .A2(n19985), .ZN(n19986) );
  OAI21_X1 U22840 ( .B1(n19987), .B2(n20088), .A(n19986), .ZN(P1_U2940) );
  NAND2_X1 U22841 ( .A1(n20031), .A2(n19988), .ZN(n20051) );
  NAND2_X1 U22842 ( .A1(n20084), .A2(P1_UWORD_REG_4__SCAN_IN), .ZN(n19989) );
  AND2_X1 U22843 ( .A1(n20051), .A2(n19989), .ZN(n19990) );
  OAI21_X1 U22844 ( .B1(n19991), .B2(n20088), .A(n19990), .ZN(P1_U2941) );
  INV_X1 U22845 ( .A(n20134), .ZN(n19992) );
  NAND2_X1 U22846 ( .A1(n20031), .A2(n19992), .ZN(n20055) );
  NAND2_X1 U22847 ( .A1(n20084), .A2(P1_UWORD_REG_5__SCAN_IN), .ZN(n19993) );
  AND2_X1 U22848 ( .A1(n20055), .A2(n19993), .ZN(n19994) );
  OAI21_X1 U22849 ( .B1(n19995), .B2(n20088), .A(n19994), .ZN(P1_U2942) );
  INV_X1 U22850 ( .A(n20137), .ZN(n19996) );
  NAND2_X1 U22851 ( .A1(n20031), .A2(n19996), .ZN(n20058) );
  NAND2_X1 U22852 ( .A1(n20084), .A2(P1_UWORD_REG_6__SCAN_IN), .ZN(n19997) );
  AND2_X1 U22853 ( .A1(n20058), .A2(n19997), .ZN(n19998) );
  OAI21_X1 U22854 ( .B1(n19999), .B2(n20088), .A(n19998), .ZN(P1_U2943) );
  INV_X1 U22855 ( .A(n20144), .ZN(n20000) );
  NAND2_X1 U22856 ( .A1(n20031), .A2(n20000), .ZN(n20061) );
  NAND2_X1 U22857 ( .A1(n20084), .A2(P1_UWORD_REG_7__SCAN_IN), .ZN(n20001) );
  AND2_X1 U22858 ( .A1(n20061), .A2(n20001), .ZN(n20002) );
  OAI21_X1 U22859 ( .B1(n20807), .B2(n20088), .A(n20002), .ZN(P1_U2944) );
  INV_X1 U22860 ( .A(n20003), .ZN(n20004) );
  NAND2_X1 U22861 ( .A1(n20031), .A2(n20004), .ZN(n20064) );
  NAND2_X1 U22862 ( .A1(n20084), .A2(P1_UWORD_REG_8__SCAN_IN), .ZN(n20005) );
  AND2_X1 U22863 ( .A1(n20064), .A2(n20005), .ZN(n20006) );
  OAI21_X1 U22864 ( .B1(n20007), .B2(n20088), .A(n20006), .ZN(P1_U2945) );
  NAND2_X1 U22865 ( .A1(n20031), .A2(n20008), .ZN(n20067) );
  NAND2_X1 U22866 ( .A1(n20084), .A2(P1_UWORD_REG_9__SCAN_IN), .ZN(n20009) );
  AND2_X1 U22867 ( .A1(n20067), .A2(n20009), .ZN(n20010) );
  OAI21_X1 U22868 ( .B1(n20011), .B2(n20088), .A(n20010), .ZN(P1_U2946) );
  INV_X1 U22869 ( .A(n20012), .ZN(n20013) );
  NAND2_X1 U22870 ( .A1(n20031), .A2(n20013), .ZN(n20071) );
  NAND2_X1 U22871 ( .A1(n20084), .A2(P1_UWORD_REG_10__SCAN_IN), .ZN(n20014) );
  AND2_X1 U22872 ( .A1(n20071), .A2(n20014), .ZN(n20015) );
  OAI21_X1 U22873 ( .B1(n20016), .B2(n20088), .A(n20015), .ZN(P1_U2947) );
  INV_X1 U22874 ( .A(n20017), .ZN(n20018) );
  NAND2_X1 U22875 ( .A1(n20031), .A2(n20018), .ZN(n20074) );
  NAND2_X1 U22876 ( .A1(n20084), .A2(P1_UWORD_REG_11__SCAN_IN), .ZN(n20019) );
  AND2_X1 U22877 ( .A1(n20074), .A2(n20019), .ZN(n20020) );
  OAI21_X1 U22878 ( .B1(n20021), .B2(n20088), .A(n20020), .ZN(P1_U2948) );
  NAND2_X1 U22879 ( .A1(n20031), .A2(n20022), .ZN(n20077) );
  NAND2_X1 U22880 ( .A1(n20084), .A2(P1_UWORD_REG_12__SCAN_IN), .ZN(n20023) );
  AND2_X1 U22881 ( .A1(n20077), .A2(n20023), .ZN(n20024) );
  OAI21_X1 U22882 ( .B1(n20025), .B2(n20088), .A(n20024), .ZN(P1_U2949) );
  NAND2_X1 U22883 ( .A1(n20031), .A2(n20026), .ZN(n20081) );
  NAND2_X1 U22884 ( .A1(n20084), .A2(P1_UWORD_REG_13__SCAN_IN), .ZN(n20027) );
  AND2_X1 U22885 ( .A1(n20081), .A2(n20027), .ZN(n20028) );
  OAI21_X1 U22886 ( .B1(n20029), .B2(n20088), .A(n20028), .ZN(P1_U2950) );
  NAND2_X1 U22887 ( .A1(n20031), .A2(n20030), .ZN(n20086) );
  NAND2_X1 U22888 ( .A1(n20084), .A2(P1_UWORD_REG_14__SCAN_IN), .ZN(n20032) );
  AND2_X1 U22889 ( .A1(n20086), .A2(n20032), .ZN(n20033) );
  OAI21_X1 U22890 ( .B1(n20034), .B2(n20088), .A(n20033), .ZN(P1_U2951) );
  NAND2_X1 U22891 ( .A1(n20084), .A2(P1_LWORD_REG_0__SCAN_IN), .ZN(n20035) );
  AND2_X1 U22892 ( .A1(n20036), .A2(n20035), .ZN(n20037) );
  OAI21_X1 U22893 ( .B1(n20038), .B2(n20088), .A(n20037), .ZN(P1_U2952) );
  NAND2_X1 U22894 ( .A1(n20084), .A2(P1_LWORD_REG_1__SCAN_IN), .ZN(n20039) );
  AND2_X1 U22895 ( .A1(n20040), .A2(n20039), .ZN(n20041) );
  OAI21_X1 U22896 ( .B1(n20042), .B2(n20088), .A(n20041), .ZN(P1_U2953) );
  NAND2_X1 U22897 ( .A1(n20084), .A2(P1_LWORD_REG_2__SCAN_IN), .ZN(n20043) );
  AND2_X1 U22898 ( .A1(n20044), .A2(n20043), .ZN(n20045) );
  OAI21_X1 U22899 ( .B1(n20866), .B2(n20088), .A(n20045), .ZN(P1_U2954) );
  NAND2_X1 U22900 ( .A1(n20084), .A2(P1_LWORD_REG_3__SCAN_IN), .ZN(n20046) );
  AND2_X1 U22901 ( .A1(n20047), .A2(n20046), .ZN(n20048) );
  OAI21_X1 U22902 ( .B1(n20049), .B2(n20088), .A(n20048), .ZN(P1_U2955) );
  NAND2_X1 U22903 ( .A1(n20084), .A2(P1_LWORD_REG_4__SCAN_IN), .ZN(n20050) );
  AND2_X1 U22904 ( .A1(n20051), .A2(n20050), .ZN(n20052) );
  OAI21_X1 U22905 ( .B1(n20053), .B2(n20088), .A(n20052), .ZN(P1_U2956) );
  NAND2_X1 U22906 ( .A1(n20084), .A2(P1_LWORD_REG_5__SCAN_IN), .ZN(n20054) );
  AND2_X1 U22907 ( .A1(n20055), .A2(n20054), .ZN(n20056) );
  OAI21_X1 U22908 ( .B1(n13728), .B2(n20088), .A(n20056), .ZN(P1_U2957) );
  NAND2_X1 U22909 ( .A1(n20084), .A2(P1_LWORD_REG_6__SCAN_IN), .ZN(n20057) );
  AND2_X1 U22910 ( .A1(n20058), .A2(n20057), .ZN(n20059) );
  OAI21_X1 U22911 ( .B1(n11870), .B2(n20088), .A(n20059), .ZN(P1_U2958) );
  NAND2_X1 U22912 ( .A1(n20084), .A2(P1_LWORD_REG_7__SCAN_IN), .ZN(n20060) );
  AND2_X1 U22913 ( .A1(n20061), .A2(n20060), .ZN(n20062) );
  OAI21_X1 U22914 ( .B1(n11878), .B2(n20088), .A(n20062), .ZN(P1_U2959) );
  NAND2_X1 U22915 ( .A1(n20084), .A2(P1_LWORD_REG_8__SCAN_IN), .ZN(n20063) );
  AND2_X1 U22916 ( .A1(n20064), .A2(n20063), .ZN(n20065) );
  OAI21_X1 U22917 ( .B1(n14028), .B2(n20088), .A(n20065), .ZN(P1_U2960) );
  NAND2_X1 U22918 ( .A1(n20084), .A2(P1_LWORD_REG_9__SCAN_IN), .ZN(n20066) );
  AND2_X1 U22919 ( .A1(n20067), .A2(n20066), .ZN(n20068) );
  OAI21_X1 U22920 ( .B1(n20069), .B2(n20088), .A(n20068), .ZN(P1_U2961) );
  NAND2_X1 U22921 ( .A1(n20084), .A2(P1_LWORD_REG_10__SCAN_IN), .ZN(n20070) );
  AND2_X1 U22922 ( .A1(n20071), .A2(n20070), .ZN(n20072) );
  OAI21_X1 U22923 ( .B1(n14213), .B2(n20088), .A(n20072), .ZN(P1_U2962) );
  NAND2_X1 U22924 ( .A1(n20084), .A2(P1_LWORD_REG_11__SCAN_IN), .ZN(n20073) );
  AND2_X1 U22925 ( .A1(n20074), .A2(n20073), .ZN(n20075) );
  OAI21_X1 U22926 ( .B1(n14323), .B2(n20088), .A(n20075), .ZN(P1_U2963) );
  NAND2_X1 U22927 ( .A1(n20084), .A2(P1_LWORD_REG_12__SCAN_IN), .ZN(n20076) );
  AND2_X1 U22928 ( .A1(n20077), .A2(n20076), .ZN(n20078) );
  OAI21_X1 U22929 ( .B1(n20079), .B2(n20088), .A(n20078), .ZN(P1_U2964) );
  NAND2_X1 U22930 ( .A1(n20084), .A2(P1_LWORD_REG_13__SCAN_IN), .ZN(n20080) );
  AND2_X1 U22931 ( .A1(n20081), .A2(n20080), .ZN(n20082) );
  OAI21_X1 U22932 ( .B1(n20083), .B2(n20088), .A(n20082), .ZN(P1_U2965) );
  NAND2_X1 U22933 ( .A1(n20084), .A2(P1_LWORD_REG_14__SCAN_IN), .ZN(n20085) );
  AND2_X1 U22934 ( .A1(n20086), .A2(n20085), .ZN(n20087) );
  OAI21_X1 U22935 ( .B1(n20089), .B2(n20088), .A(n20087), .ZN(P1_U2966) );
  OR2_X1 U22936 ( .A1(n20091), .A2(n20090), .ZN(n20092) );
  AOI22_X1 U22937 ( .A1(n20094), .A2(n20093), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20092), .ZN(n20096) );
  OAI211_X1 U22938 ( .C1(n20097), .C2(n20102), .A(n20096), .B(n20095), .ZN(
        P1_U2999) );
  NOR2_X1 U22939 ( .A1(n20098), .A2(n20736), .ZN(P1_U3032) );
  AOI22_X1 U22940 ( .A1(DATAI_16_), .A2(n20100), .B1(BUF1_REG_16__SCAN_IN), 
        .B2(n20140), .ZN(n20561) );
  AOI22_X1 U22941 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20140), .B1(DATAI_24_), 
        .B2(n20100), .ZN(n20611) );
  INV_X1 U22942 ( .A(n20611), .ZN(n20558) );
  NOR2_X2 U22943 ( .A1(n20142), .A2(n20105), .ZN(n20600) );
  NOR3_X1 U22944 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20153) );
  NAND2_X1 U22945 ( .A1(n20519), .A2(n20153), .ZN(n20110) );
  INV_X1 U22946 ( .A(n20110), .ZN(n20143) );
  AOI22_X1 U22947 ( .A1(n20653), .A2(n20558), .B1(n20600), .B2(n20143), .ZN(
        n20119) );
  NOR2_X1 U22948 ( .A1(n20428), .A2(n20373), .ZN(n20115) );
  NAND2_X1 U22949 ( .A1(n20114), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20549) );
  INV_X1 U22950 ( .A(n20549), .ZN(n20106) );
  AOI21_X1 U22951 ( .B1(n20175), .B2(n20107), .A(n20753), .ZN(n20108) );
  NOR2_X1 U22952 ( .A1(n20108), .A2(n20728), .ZN(n20113) );
  INV_X1 U22953 ( .A(n20491), .ZN(n20109) );
  OR2_X1 U22954 ( .A1(n20735), .A2(n20109), .ZN(n20179) );
  OR2_X1 U22955 ( .A1(n20179), .A2(n20553), .ZN(n20116) );
  AOI22_X1 U22956 ( .A1(n20113), .A2(n20116), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20110), .ZN(n20111) );
  OAI211_X1 U22957 ( .C1(n20115), .C2(n20752), .A(n20430), .B(n20111), .ZN(
        n20146) );
  NOR2_X2 U22958 ( .A1(n20112), .A2(n20265), .ZN(n20601) );
  INV_X1 U22959 ( .A(n20113), .ZN(n20117) );
  NOR2_X1 U22960 ( .A1(n20114), .A2(n20752), .ZN(n20266) );
  INV_X1 U22961 ( .A(n20266), .ZN(n20432) );
  INV_X1 U22962 ( .A(n20115), .ZN(n20260) );
  AOI22_X1 U22963 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20146), .B1(
        n20601), .B2(n20145), .ZN(n20118) );
  OAI211_X1 U22964 ( .C1(n20561), .C2(n20175), .A(n20119), .B(n20118), .ZN(
        P1_U3033) );
  AOI22_X1 U22965 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n20140), .B1(DATAI_17_), 
        .B2(n20100), .ZN(n20565) );
  AOI22_X1 U22966 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n20140), .B1(DATAI_25_), 
        .B2(n20100), .ZN(n20617) );
  INV_X1 U22967 ( .A(n20617), .ZN(n20562) );
  NOR2_X2 U22968 ( .A1(n20142), .A2(n20120), .ZN(n20612) );
  AOI22_X1 U22969 ( .A1(n20653), .A2(n20562), .B1(n20612), .B2(n20143), .ZN(
        n20123) );
  NOR2_X2 U22970 ( .A1(n20121), .A2(n20265), .ZN(n20613) );
  AOI22_X1 U22971 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20146), .B1(
        n20613), .B2(n20145), .ZN(n20122) );
  OAI211_X1 U22972 ( .C1(n20565), .C2(n20175), .A(n20123), .B(n20122), .ZN(
        P1_U3034) );
  AOI22_X1 U22973 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20140), .B1(DATAI_18_), 
        .B2(n20100), .ZN(n20569) );
  INV_X1 U22974 ( .A(n20623), .ZN(n20566) );
  AOI22_X1 U22975 ( .A1(n20653), .A2(n20566), .B1(n20618), .B2(n20143), .ZN(
        n20126) );
  NOR2_X2 U22976 ( .A1(n20124), .A2(n20265), .ZN(n20619) );
  AOI22_X1 U22977 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20146), .B1(
        n20619), .B2(n20145), .ZN(n20125) );
  OAI211_X1 U22978 ( .C1(n20569), .C2(n20175), .A(n20126), .B(n20125), .ZN(
        P1_U3035) );
  AOI22_X1 U22979 ( .A1(DATAI_19_), .A2(n20100), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n20140), .ZN(n20573) );
  AOI22_X1 U22980 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20140), .B1(DATAI_27_), 
        .B2(n20100), .ZN(n20629) );
  INV_X1 U22981 ( .A(n20629), .ZN(n20570) );
  NOR2_X2 U22982 ( .A1(n20142), .A2(n20127), .ZN(n20624) );
  AOI22_X1 U22983 ( .A1(n20653), .A2(n20570), .B1(n20624), .B2(n20143), .ZN(
        n20130) );
  NOR2_X2 U22984 ( .A1(n20128), .A2(n20265), .ZN(n20625) );
  AOI22_X1 U22985 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20146), .B1(
        n20625), .B2(n20145), .ZN(n20129) );
  OAI211_X1 U22986 ( .C1(n20573), .C2(n20175), .A(n20130), .B(n20129), .ZN(
        P1_U3036) );
  AOI22_X1 U22987 ( .A1(DATAI_20_), .A2(n20100), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n20140), .ZN(n20577) );
  AOI22_X1 U22988 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20140), .B1(DATAI_28_), 
        .B2(n20100), .ZN(n20635) );
  INV_X1 U22989 ( .A(n20635), .ZN(n20574) );
  NOR2_X2 U22990 ( .A1(n20142), .A2(n11626), .ZN(n20630) );
  AOI22_X1 U22991 ( .A1(n20653), .A2(n20574), .B1(n20630), .B2(n20143), .ZN(
        n20133) );
  NOR2_X2 U22992 ( .A1(n20131), .A2(n20265), .ZN(n20631) );
  AOI22_X1 U22993 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20146), .B1(
        n20631), .B2(n20145), .ZN(n20132) );
  OAI211_X1 U22994 ( .C1(n20577), .C2(n20175), .A(n20133), .B(n20132), .ZN(
        P1_U3037) );
  AOI22_X1 U22995 ( .A1(DATAI_21_), .A2(n20100), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n20140), .ZN(n20581) );
  AOI22_X1 U22996 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20140), .B1(DATAI_29_), 
        .B2(n20100), .ZN(n20641) );
  INV_X1 U22997 ( .A(n20641), .ZN(n20578) );
  AOI22_X1 U22998 ( .A1(n20653), .A2(n20578), .B1(n20636), .B2(n20143), .ZN(
        n20136) );
  NOR2_X2 U22999 ( .A1(n20134), .A2(n20265), .ZN(n20637) );
  AOI22_X1 U23000 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20146), .B1(
        n20637), .B2(n20145), .ZN(n20135) );
  OAI211_X1 U23001 ( .C1(n20581), .C2(n20175), .A(n20136), .B(n20135), .ZN(
        P1_U3038) );
  AOI22_X1 U23002 ( .A1(DATAI_22_), .A2(n20100), .B1(BUF1_REG_22__SCAN_IN), 
        .B2(n20140), .ZN(n20585) );
  AOI22_X1 U23003 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20140), .B1(DATAI_30_), 
        .B2(n20100), .ZN(n20647) );
  INV_X1 U23004 ( .A(n20647), .ZN(n20582) );
  NOR2_X2 U23005 ( .A1(n20142), .A2(n9938), .ZN(n20642) );
  AOI22_X1 U23006 ( .A1(n20653), .A2(n20582), .B1(n20642), .B2(n20143), .ZN(
        n20139) );
  NOR2_X2 U23007 ( .A1(n20137), .A2(n20265), .ZN(n20643) );
  AOI22_X1 U23008 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20146), .B1(
        n20643), .B2(n20145), .ZN(n20138) );
  OAI211_X1 U23009 ( .C1(n20585), .C2(n20175), .A(n20139), .B(n20138), .ZN(
        P1_U3039) );
  AOI22_X1 U23010 ( .A1(DATAI_23_), .A2(n20100), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n20140), .ZN(n20593) );
  AOI22_X1 U23011 ( .A1(DATAI_31_), .A2(n20100), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20140), .ZN(n20658) );
  INV_X1 U23012 ( .A(n20658), .ZN(n20588) );
  NOR2_X2 U23013 ( .A1(n20142), .A2(n20141), .ZN(n20649) );
  AOI22_X1 U23014 ( .A1(n20653), .A2(n20588), .B1(n20649), .B2(n20143), .ZN(
        n20148) );
  NOR2_X2 U23015 ( .A1(n20144), .A2(n20265), .ZN(n20650) );
  AOI22_X1 U23016 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20146), .B1(
        n20650), .B2(n20145), .ZN(n20147) );
  OAI211_X1 U23017 ( .C1(n20593), .C2(n20175), .A(n20148), .B(n20147), .ZN(
        P1_U3040) );
  INV_X1 U23018 ( .A(n20179), .ZN(n20216) );
  INV_X1 U23019 ( .A(n20149), .ZN(n20520) );
  INV_X1 U23020 ( .A(n20153), .ZN(n20150) );
  NOR2_X1 U23021 ( .A1(n20519), .A2(n20150), .ZN(n20169) );
  AOI21_X1 U23022 ( .B1(n20216), .B2(n20520), .A(n20169), .ZN(n20151) );
  OAI22_X1 U23023 ( .A1(n20151), .A2(n20728), .B1(n20150), .B2(n20752), .ZN(
        n20170) );
  AOI22_X1 U23024 ( .A1(n20601), .A2(n20170), .B1(n20600), .B2(n20169), .ZN(
        n20155) );
  OAI211_X1 U23025 ( .C1(n20217), .C2(n20753), .A(n20602), .B(n20151), .ZN(
        n20152) );
  OAI211_X1 U23026 ( .C1(n20602), .C2(n20153), .A(n20606), .B(n20152), .ZN(
        n20172) );
  OR2_X1 U23027 ( .A1(n9593), .A2(n13249), .ZN(n20525) );
  INV_X1 U23028 ( .A(n20210), .ZN(n20171) );
  INV_X1 U23029 ( .A(n20561), .ZN(n20608) );
  AOI22_X1 U23030 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20172), .B1(
        n20171), .B2(n20608), .ZN(n20154) );
  OAI211_X1 U23031 ( .C1(n20611), .C2(n20175), .A(n20155), .B(n20154), .ZN(
        P1_U3041) );
  AOI22_X1 U23032 ( .A1(n20613), .A2(n20170), .B1(n20612), .B2(n20169), .ZN(
        n20157) );
  INV_X1 U23033 ( .A(n20175), .ZN(n20166) );
  AOI22_X1 U23034 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20172), .B1(
        n20166), .B2(n20562), .ZN(n20156) );
  OAI211_X1 U23035 ( .C1(n20565), .C2(n20210), .A(n20157), .B(n20156), .ZN(
        P1_U3042) );
  AOI22_X1 U23036 ( .A1(n20619), .A2(n20170), .B1(n20618), .B2(n20169), .ZN(
        n20159) );
  AOI22_X1 U23037 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20172), .B1(
        n20166), .B2(n20566), .ZN(n20158) );
  OAI211_X1 U23038 ( .C1(n20569), .C2(n20210), .A(n20159), .B(n20158), .ZN(
        P1_U3043) );
  AOI22_X1 U23039 ( .A1(n20625), .A2(n20170), .B1(n20624), .B2(n20169), .ZN(
        n20161) );
  AOI22_X1 U23040 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20172), .B1(
        n20166), .B2(n20570), .ZN(n20160) );
  OAI211_X1 U23041 ( .C1(n20573), .C2(n20210), .A(n20161), .B(n20160), .ZN(
        P1_U3044) );
  AOI22_X1 U23042 ( .A1(n20631), .A2(n20170), .B1(n20630), .B2(n20169), .ZN(
        n20163) );
  INV_X1 U23043 ( .A(n20577), .ZN(n20632) );
  AOI22_X1 U23044 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20172), .B1(
        n20171), .B2(n20632), .ZN(n20162) );
  OAI211_X1 U23045 ( .C1(n20635), .C2(n20175), .A(n20163), .B(n20162), .ZN(
        P1_U3045) );
  AOI22_X1 U23046 ( .A1(n20637), .A2(n20170), .B1(n20636), .B2(n20169), .ZN(
        n20165) );
  AOI22_X1 U23047 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20172), .B1(
        n20166), .B2(n20578), .ZN(n20164) );
  OAI211_X1 U23048 ( .C1(n20581), .C2(n20210), .A(n20165), .B(n20164), .ZN(
        P1_U3046) );
  AOI22_X1 U23049 ( .A1(n20643), .A2(n20170), .B1(n20642), .B2(n20169), .ZN(
        n20168) );
  AOI22_X1 U23050 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20172), .B1(
        n20166), .B2(n20582), .ZN(n20167) );
  OAI211_X1 U23051 ( .C1(n20585), .C2(n20210), .A(n20168), .B(n20167), .ZN(
        P1_U3047) );
  AOI22_X1 U23052 ( .A1(n20650), .A2(n20170), .B1(n20649), .B2(n20169), .ZN(
        n20174) );
  INV_X1 U23053 ( .A(n20593), .ZN(n20652) );
  AOI22_X1 U23054 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20172), .B1(
        n20171), .B2(n20652), .ZN(n20173) );
  OAI211_X1 U23055 ( .C1(n20658), .C2(n20175), .A(n20174), .B(n20173), .ZN(
        P1_U3048) );
  AND2_X1 U23056 ( .A1(n9593), .A2(n13249), .ZN(n20546) );
  INV_X1 U23057 ( .A(n20546), .ZN(n20312) );
  INV_X1 U23058 ( .A(n20600), .ZN(n20212) );
  NAND3_X1 U23059 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20738), .A3(
        n20488), .ZN(n20221) );
  OR2_X1 U23060 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20221), .ZN(
        n20204) );
  OAI22_X1 U23061 ( .A1(n20210), .A2(n20611), .B1(n20212), .B2(n20204), .ZN(
        n20176) );
  INV_X1 U23062 ( .A(n20176), .ZN(n20185) );
  INV_X1 U23063 ( .A(n20217), .ZN(n20178) );
  NAND3_X1 U23064 ( .A1(n20343), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(n20487), 
        .ZN(n20177) );
  NAND2_X1 U23065 ( .A1(n20177), .A2(n20602), .ZN(n20425) );
  OAI21_X1 U23066 ( .B1(n20178), .B2(n20728), .A(n20425), .ZN(n20181) );
  OR2_X1 U23067 ( .A1(n20179), .A2(n13348), .ZN(n20182) );
  AOI22_X1 U23068 ( .A1(n20181), .A2(n20182), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20204), .ZN(n20180) );
  NAND2_X1 U23069 ( .A1(n20428), .A2(n20738), .ZN(n20319) );
  NAND2_X1 U23070 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20319), .ZN(n20316) );
  NAND3_X1 U23071 ( .A1(n20430), .A2(n20180), .A3(n20316), .ZN(n20207) );
  INV_X1 U23072 ( .A(n20181), .ZN(n20183) );
  OAI22_X1 U23073 ( .A1(n20183), .A2(n20182), .B1(n20432), .B2(n20319), .ZN(
        n20206) );
  AOI22_X1 U23074 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20207), .B1(
        n20601), .B2(n20206), .ZN(n20184) );
  OAI211_X1 U23075 ( .C1(n20561), .C2(n20257), .A(n20185), .B(n20184), .ZN(
        P1_U3049) );
  INV_X1 U23076 ( .A(n20612), .ZN(n20226) );
  OAI22_X1 U23077 ( .A1(n20210), .A2(n20617), .B1(n20226), .B2(n20204), .ZN(
        n20186) );
  INV_X1 U23078 ( .A(n20186), .ZN(n20188) );
  AOI22_X1 U23079 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20207), .B1(
        n20613), .B2(n20206), .ZN(n20187) );
  OAI211_X1 U23080 ( .C1(n20565), .C2(n20257), .A(n20188), .B(n20187), .ZN(
        P1_U3050) );
  INV_X1 U23081 ( .A(n20618), .ZN(n20230) );
  OAI22_X1 U23082 ( .A1(n20257), .A2(n20569), .B1(n20230), .B2(n20204), .ZN(
        n20189) );
  INV_X1 U23083 ( .A(n20189), .ZN(n20191) );
  AOI22_X1 U23084 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20207), .B1(
        n20619), .B2(n20206), .ZN(n20190) );
  OAI211_X1 U23085 ( .C1(n20623), .C2(n20210), .A(n20191), .B(n20190), .ZN(
        P1_U3051) );
  INV_X1 U23086 ( .A(n20624), .ZN(n20234) );
  OAI22_X1 U23087 ( .A1(n20257), .A2(n20573), .B1(n20234), .B2(n20204), .ZN(
        n20192) );
  INV_X1 U23088 ( .A(n20192), .ZN(n20194) );
  AOI22_X1 U23089 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20207), .B1(
        n20625), .B2(n20206), .ZN(n20193) );
  OAI211_X1 U23090 ( .C1(n20629), .C2(n20210), .A(n20194), .B(n20193), .ZN(
        P1_U3052) );
  INV_X1 U23091 ( .A(n20630), .ZN(n20238) );
  OAI22_X1 U23092 ( .A1(n20210), .A2(n20635), .B1(n20238), .B2(n20204), .ZN(
        n20195) );
  INV_X1 U23093 ( .A(n20195), .ZN(n20197) );
  AOI22_X1 U23094 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20207), .B1(
        n20631), .B2(n20206), .ZN(n20196) );
  OAI211_X1 U23095 ( .C1(n20577), .C2(n20257), .A(n20197), .B(n20196), .ZN(
        P1_U3053) );
  INV_X1 U23096 ( .A(n20636), .ZN(n20242) );
  OAI22_X1 U23097 ( .A1(n20210), .A2(n20641), .B1(n20242), .B2(n20204), .ZN(
        n20198) );
  INV_X1 U23098 ( .A(n20198), .ZN(n20200) );
  AOI22_X1 U23099 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20207), .B1(
        n20637), .B2(n20206), .ZN(n20199) );
  OAI211_X1 U23100 ( .C1(n20581), .C2(n20257), .A(n20200), .B(n20199), .ZN(
        P1_U3054) );
  INV_X1 U23101 ( .A(n20642), .ZN(n20246) );
  OAI22_X1 U23102 ( .A1(n20257), .A2(n20585), .B1(n20246), .B2(n20204), .ZN(
        n20201) );
  INV_X1 U23103 ( .A(n20201), .ZN(n20203) );
  AOI22_X1 U23104 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20207), .B1(
        n20643), .B2(n20206), .ZN(n20202) );
  OAI211_X1 U23105 ( .C1(n20647), .C2(n20210), .A(n20203), .B(n20202), .ZN(
        P1_U3055) );
  INV_X1 U23106 ( .A(n20649), .ZN(n20251) );
  OAI22_X1 U23107 ( .A1(n20257), .A2(n20593), .B1(n20251), .B2(n20204), .ZN(
        n20205) );
  INV_X1 U23108 ( .A(n20205), .ZN(n20209) );
  AOI22_X1 U23109 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20207), .B1(
        n20650), .B2(n20206), .ZN(n20208) );
  OAI211_X1 U23110 ( .C1(n20658), .C2(n20210), .A(n20209), .B(n20208), .ZN(
        P1_U3056) );
  INV_X1 U23111 ( .A(n20458), .ZN(n20211) );
  NAND2_X1 U23112 ( .A1(n20211), .A2(n20738), .ZN(n20250) );
  OAI22_X1 U23113 ( .A1(n20262), .A2(n20561), .B1(n20212), .B2(n20250), .ZN(
        n20213) );
  INV_X1 U23114 ( .A(n20213), .ZN(n20225) );
  AND2_X1 U23115 ( .A1(n20214), .A2(n9621), .ZN(n20595) );
  INV_X1 U23116 ( .A(n20250), .ZN(n20215) );
  AOI21_X1 U23117 ( .B1(n20216), .B2(n20595), .A(n20215), .ZN(n20223) );
  OR2_X1 U23118 ( .A1(n20217), .A2(n20727), .ZN(n20218) );
  AOI22_X1 U23119 ( .A1(n20223), .A2(n20220), .B1(n20728), .B2(n20221), .ZN(
        n20219) );
  NAND2_X1 U23120 ( .A1(n20606), .A2(n20219), .ZN(n20254) );
  INV_X1 U23121 ( .A(n20220), .ZN(n20222) );
  OAI22_X1 U23122 ( .A1(n20223), .A2(n20222), .B1(n20752), .B2(n20221), .ZN(
        n20253) );
  AOI22_X1 U23123 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20254), .B1(
        n20601), .B2(n20253), .ZN(n20224) );
  OAI211_X1 U23124 ( .C1(n20611), .C2(n20257), .A(n20225), .B(n20224), .ZN(
        P1_U3057) );
  OAI22_X1 U23125 ( .A1(n20262), .A2(n20565), .B1(n20226), .B2(n20250), .ZN(
        n20227) );
  INV_X1 U23126 ( .A(n20227), .ZN(n20229) );
  AOI22_X1 U23127 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20254), .B1(
        n20613), .B2(n20253), .ZN(n20228) );
  OAI211_X1 U23128 ( .C1(n20617), .C2(n20257), .A(n20229), .B(n20228), .ZN(
        P1_U3058) );
  OAI22_X1 U23129 ( .A1(n20262), .A2(n20569), .B1(n20230), .B2(n20250), .ZN(
        n20231) );
  INV_X1 U23130 ( .A(n20231), .ZN(n20233) );
  AOI22_X1 U23131 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20254), .B1(
        n20619), .B2(n20253), .ZN(n20232) );
  OAI211_X1 U23132 ( .C1(n20623), .C2(n20257), .A(n20233), .B(n20232), .ZN(
        P1_U3059) );
  OAI22_X1 U23133 ( .A1(n20262), .A2(n20573), .B1(n20234), .B2(n20250), .ZN(
        n20235) );
  INV_X1 U23134 ( .A(n20235), .ZN(n20237) );
  AOI22_X1 U23135 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20254), .B1(
        n20625), .B2(n20253), .ZN(n20236) );
  OAI211_X1 U23136 ( .C1(n20629), .C2(n20257), .A(n20237), .B(n20236), .ZN(
        P1_U3060) );
  OAI22_X1 U23137 ( .A1(n20262), .A2(n20577), .B1(n20238), .B2(n20250), .ZN(
        n20239) );
  INV_X1 U23138 ( .A(n20239), .ZN(n20241) );
  AOI22_X1 U23139 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20254), .B1(
        n20631), .B2(n20253), .ZN(n20240) );
  OAI211_X1 U23140 ( .C1(n20635), .C2(n20257), .A(n20241), .B(n20240), .ZN(
        P1_U3061) );
  OAI22_X1 U23141 ( .A1(n20262), .A2(n20581), .B1(n20242), .B2(n20250), .ZN(
        n20243) );
  INV_X1 U23142 ( .A(n20243), .ZN(n20245) );
  AOI22_X1 U23143 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20254), .B1(
        n20637), .B2(n20253), .ZN(n20244) );
  OAI211_X1 U23144 ( .C1(n20641), .C2(n20257), .A(n20245), .B(n20244), .ZN(
        P1_U3062) );
  OAI22_X1 U23145 ( .A1(n20262), .A2(n20585), .B1(n20246), .B2(n20250), .ZN(
        n20247) );
  INV_X1 U23146 ( .A(n20247), .ZN(n20249) );
  AOI22_X1 U23147 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20254), .B1(
        n20643), .B2(n20253), .ZN(n20248) );
  OAI211_X1 U23148 ( .C1(n20647), .C2(n20257), .A(n20249), .B(n20248), .ZN(
        P1_U3063) );
  OAI22_X1 U23149 ( .A1(n20262), .A2(n20593), .B1(n20251), .B2(n20250), .ZN(
        n20252) );
  INV_X1 U23150 ( .A(n20252), .ZN(n20256) );
  AOI22_X1 U23151 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20254), .B1(
        n20650), .B2(n20253), .ZN(n20255) );
  OAI211_X1 U23152 ( .C1(n20658), .C2(n20257), .A(n20256), .B(n20255), .ZN(
        P1_U3064) );
  NOR3_X1 U23153 ( .A1(n20488), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20291) );
  INV_X1 U23154 ( .A(n20291), .ZN(n20288) );
  NOR2_X1 U23155 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20288), .ZN(
        n20283) );
  OR2_X1 U23156 ( .A1(n20491), .A2(n20259), .ZN(n20314) );
  NAND2_X1 U23157 ( .A1(n13348), .A2(n20602), .ZN(n20261) );
  OAI22_X1 U23158 ( .A1(n20314), .A2(n20261), .B1(n20260), .B2(n20549), .ZN(
        n20282) );
  AOI22_X1 U23159 ( .A1(n20600), .A2(n20283), .B1(n20601), .B2(n20282), .ZN(
        n20269) );
  INV_X1 U23160 ( .A(n20311), .ZN(n20263) );
  OAI21_X1 U23161 ( .B1(n20284), .B2(n20263), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20264) );
  OAI21_X1 U23162 ( .B1(n20553), .B2(n20314), .A(n20264), .ZN(n20267) );
  AOI22_X1 U23163 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20285), .B1(
        n20284), .B2(n20558), .ZN(n20268) );
  OAI211_X1 U23164 ( .C1(n20561), .C2(n20311), .A(n20269), .B(n20268), .ZN(
        P1_U3065) );
  AOI22_X1 U23165 ( .A1(n20612), .A2(n20283), .B1(n20613), .B2(n20282), .ZN(
        n20271) );
  AOI22_X1 U23166 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20285), .B1(
        n20284), .B2(n20562), .ZN(n20270) );
  OAI211_X1 U23167 ( .C1(n20565), .C2(n20311), .A(n20271), .B(n20270), .ZN(
        P1_U3066) );
  AOI22_X1 U23168 ( .A1(n20618), .A2(n20283), .B1(n20619), .B2(n20282), .ZN(
        n20273) );
  AOI22_X1 U23169 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20285), .B1(
        n20284), .B2(n20566), .ZN(n20272) );
  OAI211_X1 U23170 ( .C1(n20569), .C2(n20311), .A(n20273), .B(n20272), .ZN(
        P1_U3067) );
  AOI22_X1 U23171 ( .A1(n20624), .A2(n20283), .B1(n20625), .B2(n20282), .ZN(
        n20275) );
  AOI22_X1 U23172 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20285), .B1(
        n20284), .B2(n20570), .ZN(n20274) );
  OAI211_X1 U23173 ( .C1(n20573), .C2(n20311), .A(n20275), .B(n20274), .ZN(
        P1_U3068) );
  AOI22_X1 U23174 ( .A1(n20630), .A2(n20283), .B1(n20631), .B2(n20282), .ZN(
        n20277) );
  AOI22_X1 U23175 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20285), .B1(
        n20284), .B2(n20574), .ZN(n20276) );
  OAI211_X1 U23176 ( .C1(n20577), .C2(n20311), .A(n20277), .B(n20276), .ZN(
        P1_U3069) );
  AOI22_X1 U23177 ( .A1(n20636), .A2(n20283), .B1(n20637), .B2(n20282), .ZN(
        n20279) );
  AOI22_X1 U23178 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20285), .B1(
        n20284), .B2(n20578), .ZN(n20278) );
  OAI211_X1 U23179 ( .C1(n20581), .C2(n20311), .A(n20279), .B(n20278), .ZN(
        P1_U3070) );
  AOI22_X1 U23180 ( .A1(n20642), .A2(n20283), .B1(n20643), .B2(n20282), .ZN(
        n20281) );
  AOI22_X1 U23181 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20285), .B1(
        n20284), .B2(n20582), .ZN(n20280) );
  OAI211_X1 U23182 ( .C1(n20585), .C2(n20311), .A(n20281), .B(n20280), .ZN(
        P1_U3071) );
  AOI22_X1 U23183 ( .A1(n20649), .A2(n20283), .B1(n20650), .B2(n20282), .ZN(
        n20287) );
  AOI22_X1 U23184 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20285), .B1(
        n20284), .B2(n20588), .ZN(n20286) );
  OAI211_X1 U23185 ( .C1(n20593), .C2(n20311), .A(n20287), .B(n20286), .ZN(
        P1_U3072) );
  NOR2_X1 U23186 ( .A1(n20519), .A2(n20288), .ZN(n20307) );
  INV_X1 U23187 ( .A(n20314), .ZN(n20344) );
  AOI21_X1 U23188 ( .B1(n20344), .B2(n20520), .A(n20307), .ZN(n20289) );
  OAI22_X1 U23189 ( .A1(n20289), .A2(n20728), .B1(n20288), .B2(n20752), .ZN(
        n20306) );
  AOI22_X1 U23190 ( .A1(n20600), .A2(n20307), .B1(n20601), .B2(n20306), .ZN(
        n20293) );
  OAI211_X1 U23191 ( .C1(n20729), .C2(n20753), .A(n20602), .B(n20289), .ZN(
        n20290) );
  OAI211_X1 U23192 ( .C1(n20602), .C2(n20291), .A(n20606), .B(n20290), .ZN(
        n20308) );
  AOI22_X1 U23193 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20308), .B1(
        n20338), .B2(n20608), .ZN(n20292) );
  OAI211_X1 U23194 ( .C1(n20611), .C2(n20311), .A(n20293), .B(n20292), .ZN(
        P1_U3073) );
  AOI22_X1 U23195 ( .A1(n20612), .A2(n20307), .B1(n20613), .B2(n20306), .ZN(
        n20295) );
  INV_X1 U23196 ( .A(n20565), .ZN(n20614) );
  AOI22_X1 U23197 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20308), .B1(
        n20338), .B2(n20614), .ZN(n20294) );
  OAI211_X1 U23198 ( .C1(n20617), .C2(n20311), .A(n20295), .B(n20294), .ZN(
        P1_U3074) );
  AOI22_X1 U23199 ( .A1(n20618), .A2(n20307), .B1(n20619), .B2(n20306), .ZN(
        n20297) );
  INV_X1 U23200 ( .A(n20569), .ZN(n20620) );
  AOI22_X1 U23201 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20308), .B1(
        n20338), .B2(n20620), .ZN(n20296) );
  OAI211_X1 U23202 ( .C1(n20623), .C2(n20311), .A(n20297), .B(n20296), .ZN(
        P1_U3075) );
  AOI22_X1 U23203 ( .A1(n20624), .A2(n20307), .B1(n20625), .B2(n20306), .ZN(
        n20299) );
  INV_X1 U23204 ( .A(n20573), .ZN(n20626) );
  AOI22_X1 U23205 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20308), .B1(
        n20338), .B2(n20626), .ZN(n20298) );
  OAI211_X1 U23206 ( .C1(n20629), .C2(n20311), .A(n20299), .B(n20298), .ZN(
        P1_U3076) );
  AOI22_X1 U23207 ( .A1(n20630), .A2(n20307), .B1(n20631), .B2(n20306), .ZN(
        n20301) );
  AOI22_X1 U23208 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20308), .B1(
        n20338), .B2(n20632), .ZN(n20300) );
  OAI211_X1 U23209 ( .C1(n20635), .C2(n20311), .A(n20301), .B(n20300), .ZN(
        P1_U3077) );
  AOI22_X1 U23210 ( .A1(n20636), .A2(n20307), .B1(n20637), .B2(n20306), .ZN(
        n20303) );
  INV_X1 U23211 ( .A(n20581), .ZN(n20638) );
  AOI22_X1 U23212 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20308), .B1(
        n20338), .B2(n20638), .ZN(n20302) );
  OAI211_X1 U23213 ( .C1(n20641), .C2(n20311), .A(n20303), .B(n20302), .ZN(
        P1_U3078) );
  AOI22_X1 U23214 ( .A1(n20642), .A2(n20307), .B1(n20643), .B2(n20306), .ZN(
        n20305) );
  INV_X1 U23215 ( .A(n20585), .ZN(n20644) );
  AOI22_X1 U23216 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20308), .B1(
        n20338), .B2(n20644), .ZN(n20304) );
  OAI211_X1 U23217 ( .C1(n20647), .C2(n20311), .A(n20305), .B(n20304), .ZN(
        P1_U3079) );
  AOI22_X1 U23218 ( .A1(n20649), .A2(n20307), .B1(n20650), .B2(n20306), .ZN(
        n20310) );
  AOI22_X1 U23219 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20308), .B1(
        n20338), .B2(n20652), .ZN(n20309) );
  OAI211_X1 U23220 ( .C1(n20658), .C2(n20311), .A(n20310), .B(n20309), .ZN(
        P1_U3080) );
  INV_X1 U23221 ( .A(n20345), .ZN(n20348) );
  NAND2_X1 U23222 ( .A1(n20519), .A2(n20348), .ZN(n20315) );
  INV_X1 U23223 ( .A(n20315), .ZN(n20337) );
  AOI22_X1 U23224 ( .A1(n20338), .A2(n20558), .B1(n20600), .B2(n20337), .ZN(
        n20323) );
  OAI21_X1 U23225 ( .B1(n20313), .B2(n20728), .A(n20425), .ZN(n20318) );
  OR2_X1 U23226 ( .A1(n20314), .A2(n13348), .ZN(n20320) );
  AOI22_X1 U23227 ( .A1(n20318), .A2(n20320), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20315), .ZN(n20317) );
  NAND3_X1 U23228 ( .A1(n20556), .A2(n20317), .A3(n20316), .ZN(n20340) );
  INV_X1 U23229 ( .A(n20318), .ZN(n20321) );
  OAI22_X1 U23230 ( .A1(n20321), .A2(n20320), .B1(n20549), .B2(n20319), .ZN(
        n20339) );
  AOI22_X1 U23231 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20340), .B1(
        n20601), .B2(n20339), .ZN(n20322) );
  OAI211_X1 U23232 ( .C1(n20561), .C2(n20361), .A(n20323), .B(n20322), .ZN(
        P1_U3081) );
  AOI22_X1 U23233 ( .A1(n20338), .A2(n20562), .B1(n20612), .B2(n20337), .ZN(
        n20325) );
  AOI22_X1 U23234 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20340), .B1(
        n20613), .B2(n20339), .ZN(n20324) );
  OAI211_X1 U23235 ( .C1(n20565), .C2(n20361), .A(n20325), .B(n20324), .ZN(
        P1_U3082) );
  AOI22_X1 U23236 ( .A1(n20366), .A2(n20620), .B1(n20618), .B2(n20337), .ZN(
        n20327) );
  AOI22_X1 U23237 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20340), .B1(
        n20619), .B2(n20339), .ZN(n20326) );
  OAI211_X1 U23238 ( .C1(n20623), .C2(n20336), .A(n20327), .B(n20326), .ZN(
        P1_U3083) );
  AOI22_X1 U23239 ( .A1(n20338), .A2(n20570), .B1(n20624), .B2(n20337), .ZN(
        n20329) );
  AOI22_X1 U23240 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20340), .B1(
        n20625), .B2(n20339), .ZN(n20328) );
  OAI211_X1 U23241 ( .C1(n20573), .C2(n20361), .A(n20329), .B(n20328), .ZN(
        P1_U3084) );
  AOI22_X1 U23242 ( .A1(n20338), .A2(n20574), .B1(n20630), .B2(n20337), .ZN(
        n20331) );
  AOI22_X1 U23243 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20340), .B1(
        n20631), .B2(n20339), .ZN(n20330) );
  OAI211_X1 U23244 ( .C1(n20577), .C2(n20361), .A(n20331), .B(n20330), .ZN(
        P1_U3085) );
  AOI22_X1 U23245 ( .A1(n20366), .A2(n20638), .B1(n20636), .B2(n20337), .ZN(
        n20333) );
  AOI22_X1 U23246 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20340), .B1(
        n20637), .B2(n20339), .ZN(n20332) );
  OAI211_X1 U23247 ( .C1(n20641), .C2(n20336), .A(n20333), .B(n20332), .ZN(
        P1_U3086) );
  AOI22_X1 U23248 ( .A1(n20366), .A2(n20644), .B1(n20642), .B2(n20337), .ZN(
        n20335) );
  AOI22_X1 U23249 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20340), .B1(
        n20643), .B2(n20339), .ZN(n20334) );
  OAI211_X1 U23250 ( .C1(n20647), .C2(n20336), .A(n20335), .B(n20334), .ZN(
        P1_U3087) );
  AOI22_X1 U23251 ( .A1(n20338), .A2(n20588), .B1(n20649), .B2(n20337), .ZN(
        n20342) );
  AOI22_X1 U23252 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20340), .B1(
        n20650), .B2(n20339), .ZN(n20341) );
  OAI211_X1 U23253 ( .C1(n20593), .C2(n20361), .A(n20342), .B(n20341), .ZN(
        P1_U3088) );
  AOI21_X1 U23254 ( .B1(n20344), .B2(n20595), .A(n20365), .ZN(n20346) );
  OAI22_X1 U23255 ( .A1(n20346), .A2(n20728), .B1(n20345), .B2(n20752), .ZN(
        n20364) );
  AOI22_X1 U23256 ( .A1(n20600), .A2(n20365), .B1(n20601), .B2(n20364), .ZN(
        n20350) );
  OAI211_X1 U23257 ( .C1(n20729), .C2(n20727), .A(n20602), .B(n20346), .ZN(
        n20347) );
  OAI211_X1 U23258 ( .C1(n20348), .C2(n20602), .A(n20606), .B(n20347), .ZN(
        n20367) );
  AOI22_X1 U23259 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20367), .B1(
        n20366), .B2(n20558), .ZN(n20349) );
  OAI211_X1 U23260 ( .C1(n20561), .C2(n20370), .A(n20350), .B(n20349), .ZN(
        P1_U3089) );
  AOI22_X1 U23261 ( .A1(n20612), .A2(n20365), .B1(n20613), .B2(n20364), .ZN(
        n20352) );
  AOI22_X1 U23262 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20367), .B1(
        n20366), .B2(n20562), .ZN(n20351) );
  OAI211_X1 U23263 ( .C1(n20565), .C2(n20370), .A(n20352), .B(n20351), .ZN(
        P1_U3090) );
  AOI22_X1 U23264 ( .A1(n20618), .A2(n20365), .B1(n20619), .B2(n20364), .ZN(
        n20354) );
  AOI22_X1 U23265 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20367), .B1(
        n20395), .B2(n20620), .ZN(n20353) );
  OAI211_X1 U23266 ( .C1(n20623), .C2(n20361), .A(n20354), .B(n20353), .ZN(
        P1_U3091) );
  AOI22_X1 U23267 ( .A1(n20624), .A2(n20365), .B1(n20625), .B2(n20364), .ZN(
        n20356) );
  AOI22_X1 U23268 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20367), .B1(
        n20366), .B2(n20570), .ZN(n20355) );
  OAI211_X1 U23269 ( .C1(n20573), .C2(n20370), .A(n20356), .B(n20355), .ZN(
        P1_U3092) );
  AOI22_X1 U23270 ( .A1(n20630), .A2(n20365), .B1(n20631), .B2(n20364), .ZN(
        n20358) );
  AOI22_X1 U23271 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20367), .B1(
        n20366), .B2(n20574), .ZN(n20357) );
  OAI211_X1 U23272 ( .C1(n20577), .C2(n20370), .A(n20358), .B(n20357), .ZN(
        P1_U3093) );
  AOI22_X1 U23273 ( .A1(n20636), .A2(n20365), .B1(n20637), .B2(n20364), .ZN(
        n20360) );
  AOI22_X1 U23274 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20367), .B1(
        n20395), .B2(n20638), .ZN(n20359) );
  OAI211_X1 U23275 ( .C1(n20641), .C2(n20361), .A(n20360), .B(n20359), .ZN(
        P1_U3094) );
  AOI22_X1 U23276 ( .A1(n20642), .A2(n20365), .B1(n20643), .B2(n20364), .ZN(
        n20363) );
  AOI22_X1 U23277 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20367), .B1(
        n20366), .B2(n20582), .ZN(n20362) );
  OAI211_X1 U23278 ( .C1(n20585), .C2(n20370), .A(n20363), .B(n20362), .ZN(
        P1_U3095) );
  AOI22_X1 U23279 ( .A1(n20649), .A2(n20365), .B1(n20650), .B2(n20364), .ZN(
        n20369) );
  AOI22_X1 U23280 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20367), .B1(
        n20366), .B2(n20588), .ZN(n20368) );
  OAI211_X1 U23281 ( .C1(n20593), .C2(n20370), .A(n20369), .B(n20368), .ZN(
        P1_U3096) );
  NOR3_X1 U23282 ( .A1(n20738), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20402) );
  INV_X1 U23283 ( .A(n20402), .ZN(n20399) );
  NOR2_X1 U23284 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20399), .ZN(
        n20394) );
  NAND2_X1 U23285 ( .A1(n20735), .A2(n20491), .ZN(n20426) );
  INV_X1 U23286 ( .A(n20426), .ZN(n20459) );
  AOI21_X1 U23287 ( .B1(n20459), .B2(n13348), .A(n20394), .ZN(n20376) );
  INV_X1 U23288 ( .A(n20428), .ZN(n20374) );
  NAND2_X1 U23289 ( .A1(n20374), .A2(n20373), .ZN(n20495) );
  OAI22_X1 U23290 ( .A1(n20376), .A2(n20728), .B1(n20432), .B2(n20495), .ZN(
        n20393) );
  AOI22_X1 U23291 ( .A1(n20600), .A2(n20394), .B1(n20393), .B2(n20601), .ZN(
        n20380) );
  INV_X1 U23292 ( .A(n20423), .ZN(n20375) );
  OAI21_X1 U23293 ( .B1(n20375), .B2(n20395), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20377) );
  NAND2_X1 U23294 ( .A1(n20377), .A2(n20376), .ZN(n20378) );
  AOI22_X1 U23295 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20396), .B1(
        n20395), .B2(n20558), .ZN(n20379) );
  OAI211_X1 U23296 ( .C1(n20561), .C2(n20423), .A(n20380), .B(n20379), .ZN(
        P1_U3097) );
  AOI22_X1 U23297 ( .A1(n20612), .A2(n20394), .B1(n20393), .B2(n20613), .ZN(
        n20382) );
  AOI22_X1 U23298 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20396), .B1(
        n20395), .B2(n20562), .ZN(n20381) );
  OAI211_X1 U23299 ( .C1(n20565), .C2(n20423), .A(n20382), .B(n20381), .ZN(
        P1_U3098) );
  AOI22_X1 U23300 ( .A1(n20618), .A2(n20394), .B1(n20393), .B2(n20619), .ZN(
        n20384) );
  AOI22_X1 U23301 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20396), .B1(
        n20395), .B2(n20566), .ZN(n20383) );
  OAI211_X1 U23302 ( .C1(n20569), .C2(n20423), .A(n20384), .B(n20383), .ZN(
        P1_U3099) );
  AOI22_X1 U23303 ( .A1(n20624), .A2(n20394), .B1(n20393), .B2(n20625), .ZN(
        n20386) );
  AOI22_X1 U23304 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20396), .B1(
        n20395), .B2(n20570), .ZN(n20385) );
  OAI211_X1 U23305 ( .C1(n20573), .C2(n20423), .A(n20386), .B(n20385), .ZN(
        P1_U3100) );
  AOI22_X1 U23306 ( .A1(n20630), .A2(n20394), .B1(n20393), .B2(n20631), .ZN(
        n20388) );
  AOI22_X1 U23307 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20396), .B1(
        n20395), .B2(n20574), .ZN(n20387) );
  OAI211_X1 U23308 ( .C1(n20577), .C2(n20423), .A(n20388), .B(n20387), .ZN(
        P1_U3101) );
  AOI22_X1 U23309 ( .A1(n20636), .A2(n20394), .B1(n20393), .B2(n20637), .ZN(
        n20390) );
  AOI22_X1 U23310 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20396), .B1(
        n20395), .B2(n20578), .ZN(n20389) );
  OAI211_X1 U23311 ( .C1(n20581), .C2(n20423), .A(n20390), .B(n20389), .ZN(
        P1_U3102) );
  AOI22_X1 U23312 ( .A1(n20642), .A2(n20394), .B1(n20393), .B2(n20643), .ZN(
        n20392) );
  AOI22_X1 U23313 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20396), .B1(
        n20395), .B2(n20582), .ZN(n20391) );
  OAI211_X1 U23314 ( .C1(n20585), .C2(n20423), .A(n20392), .B(n20391), .ZN(
        P1_U3103) );
  AOI22_X1 U23315 ( .A1(n20649), .A2(n20394), .B1(n20393), .B2(n20650), .ZN(
        n20398) );
  AOI22_X1 U23316 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20396), .B1(
        n20395), .B2(n20588), .ZN(n20397) );
  OAI211_X1 U23317 ( .C1(n20593), .C2(n20423), .A(n20398), .B(n20397), .ZN(
        P1_U3104) );
  NOR2_X1 U23318 ( .A1(n20519), .A2(n20399), .ZN(n20419) );
  AOI21_X1 U23319 ( .B1(n20459), .B2(n20520), .A(n20419), .ZN(n20400) );
  OAI22_X1 U23320 ( .A1(n20400), .A2(n20728), .B1(n20399), .B2(n20752), .ZN(
        n20418) );
  AOI22_X1 U23321 ( .A1(n20600), .A2(n20419), .B1(n20418), .B2(n20601), .ZN(
        n20405) );
  INV_X1 U23322 ( .A(n20457), .ZN(n20462) );
  OAI211_X1 U23323 ( .C1(n20462), .C2(n20753), .A(n20602), .B(n20400), .ZN(
        n20401) );
  OAI211_X1 U23324 ( .C1(n20602), .C2(n20402), .A(n20606), .B(n20401), .ZN(
        n20420) );
  INV_X1 U23325 ( .A(n20525), .ZN(n20403) );
  AOI22_X1 U23326 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20420), .B1(
        n20447), .B2(n20608), .ZN(n20404) );
  OAI211_X1 U23327 ( .C1(n20611), .C2(n20423), .A(n20405), .B(n20404), .ZN(
        P1_U3105) );
  AOI22_X1 U23328 ( .A1(n20612), .A2(n20419), .B1(n20418), .B2(n20613), .ZN(
        n20407) );
  AOI22_X1 U23329 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20420), .B1(
        n20447), .B2(n20614), .ZN(n20406) );
  OAI211_X1 U23330 ( .C1(n20617), .C2(n20423), .A(n20407), .B(n20406), .ZN(
        P1_U3106) );
  AOI22_X1 U23331 ( .A1(n20618), .A2(n20419), .B1(n20418), .B2(n20619), .ZN(
        n20409) );
  AOI22_X1 U23332 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20420), .B1(
        n20447), .B2(n20620), .ZN(n20408) );
  OAI211_X1 U23333 ( .C1(n20623), .C2(n20423), .A(n20409), .B(n20408), .ZN(
        P1_U3107) );
  AOI22_X1 U23334 ( .A1(n20624), .A2(n20419), .B1(n20418), .B2(n20625), .ZN(
        n20411) );
  AOI22_X1 U23335 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20420), .B1(
        n20447), .B2(n20626), .ZN(n20410) );
  OAI211_X1 U23336 ( .C1(n20629), .C2(n20423), .A(n20411), .B(n20410), .ZN(
        P1_U3108) );
  AOI22_X1 U23337 ( .A1(n20630), .A2(n20419), .B1(n20418), .B2(n20631), .ZN(
        n20413) );
  AOI22_X1 U23338 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20420), .B1(
        n20447), .B2(n20632), .ZN(n20412) );
  OAI211_X1 U23339 ( .C1(n20635), .C2(n20423), .A(n20413), .B(n20412), .ZN(
        P1_U3109) );
  AOI22_X1 U23340 ( .A1(n20636), .A2(n20419), .B1(n20418), .B2(n20637), .ZN(
        n20415) );
  AOI22_X1 U23341 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20420), .B1(
        n20447), .B2(n20638), .ZN(n20414) );
  OAI211_X1 U23342 ( .C1(n20641), .C2(n20423), .A(n20415), .B(n20414), .ZN(
        P1_U3110) );
  AOI22_X1 U23343 ( .A1(n20642), .A2(n20419), .B1(n20418), .B2(n20643), .ZN(
        n20417) );
  AOI22_X1 U23344 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20420), .B1(
        n20447), .B2(n20644), .ZN(n20416) );
  OAI211_X1 U23345 ( .C1(n20647), .C2(n20423), .A(n20417), .B(n20416), .ZN(
        P1_U3111) );
  AOI22_X1 U23346 ( .A1(n20649), .A2(n20419), .B1(n20418), .B2(n20650), .ZN(
        n20422) );
  AOI22_X1 U23347 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20420), .B1(
        n20447), .B2(n20652), .ZN(n20421) );
  OAI211_X1 U23348 ( .C1(n20658), .C2(n20423), .A(n20422), .B(n20421), .ZN(
        P1_U3112) );
  NOR3_X1 U23349 ( .A1(n20738), .A2(n20424), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20464) );
  NAND2_X1 U23350 ( .A1(n20519), .A2(n20464), .ZN(n20427) );
  INV_X1 U23351 ( .A(n20427), .ZN(n20450) );
  AOI22_X1 U23352 ( .A1(n20483), .A2(n20608), .B1(n20600), .B2(n20450), .ZN(
        n20436) );
  OAI21_X1 U23353 ( .B1(n20457), .B2(n20728), .A(n20425), .ZN(n20431) );
  OR2_X1 U23354 ( .A1(n20426), .A2(n13348), .ZN(n20433) );
  AOI22_X1 U23355 ( .A1(n20431), .A2(n20433), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20427), .ZN(n20429) );
  NAND2_X1 U23356 ( .A1(n20428), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20550) );
  NAND2_X1 U23357 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20550), .ZN(n20555) );
  NAND3_X1 U23358 ( .A1(n20430), .A2(n20429), .A3(n20555), .ZN(n20452) );
  INV_X1 U23359 ( .A(n20431), .ZN(n20434) );
  OAI22_X1 U23360 ( .A1(n20434), .A2(n20433), .B1(n20432), .B2(n20550), .ZN(
        n20451) );
  AOI22_X1 U23361 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20452), .B1(
        n20601), .B2(n20451), .ZN(n20435) );
  OAI211_X1 U23362 ( .C1(n20611), .C2(n20455), .A(n20436), .B(n20435), .ZN(
        P1_U3113) );
  AOI22_X1 U23363 ( .A1(n20483), .A2(n20614), .B1(n20612), .B2(n20450), .ZN(
        n20438) );
  AOI22_X1 U23364 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20452), .B1(
        n20613), .B2(n20451), .ZN(n20437) );
  OAI211_X1 U23365 ( .C1(n20617), .C2(n20455), .A(n20438), .B(n20437), .ZN(
        P1_U3114) );
  AOI22_X1 U23366 ( .A1(n20483), .A2(n20620), .B1(n20618), .B2(n20450), .ZN(
        n20440) );
  AOI22_X1 U23367 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20452), .B1(
        n20619), .B2(n20451), .ZN(n20439) );
  OAI211_X1 U23368 ( .C1(n20623), .C2(n20455), .A(n20440), .B(n20439), .ZN(
        P1_U3115) );
  AOI22_X1 U23369 ( .A1(n20447), .A2(n20570), .B1(n20624), .B2(n20450), .ZN(
        n20442) );
  AOI22_X1 U23370 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20452), .B1(
        n20625), .B2(n20451), .ZN(n20441) );
  OAI211_X1 U23371 ( .C1(n20573), .C2(n20478), .A(n20442), .B(n20441), .ZN(
        P1_U3116) );
  AOI22_X1 U23372 ( .A1(n20447), .A2(n20574), .B1(n20630), .B2(n20450), .ZN(
        n20444) );
  AOI22_X1 U23373 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20452), .B1(
        n20631), .B2(n20451), .ZN(n20443) );
  OAI211_X1 U23374 ( .C1(n20577), .C2(n20478), .A(n20444), .B(n20443), .ZN(
        P1_U3117) );
  AOI22_X1 U23375 ( .A1(n20447), .A2(n20578), .B1(n20636), .B2(n20450), .ZN(
        n20446) );
  AOI22_X1 U23376 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20452), .B1(
        n20637), .B2(n20451), .ZN(n20445) );
  OAI211_X1 U23377 ( .C1(n20581), .C2(n20478), .A(n20446), .B(n20445), .ZN(
        P1_U3118) );
  AOI22_X1 U23378 ( .A1(n20447), .A2(n20582), .B1(n20642), .B2(n20450), .ZN(
        n20449) );
  AOI22_X1 U23379 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20452), .B1(
        n20643), .B2(n20451), .ZN(n20448) );
  OAI211_X1 U23380 ( .C1(n20585), .C2(n20478), .A(n20449), .B(n20448), .ZN(
        P1_U3119) );
  AOI22_X1 U23381 ( .A1(n20483), .A2(n20652), .B1(n20649), .B2(n20450), .ZN(
        n20454) );
  AOI22_X1 U23382 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20452), .B1(
        n20650), .B2(n20451), .ZN(n20453) );
  OAI211_X1 U23383 ( .C1(n20658), .C2(n20455), .A(n20454), .B(n20453), .ZN(
        P1_U3120) );
  NOR2_X1 U23384 ( .A1(n20458), .A2(n20738), .ZN(n20482) );
  AOI21_X1 U23385 ( .B1(n20459), .B2(n20595), .A(n20482), .ZN(n20461) );
  INV_X1 U23386 ( .A(n20464), .ZN(n20460) );
  OAI22_X1 U23387 ( .A1(n20461), .A2(n20728), .B1(n20460), .B2(n20752), .ZN(
        n20481) );
  AOI22_X1 U23388 ( .A1(n20600), .A2(n20482), .B1(n20481), .B2(n20601), .ZN(
        n20466) );
  OAI211_X1 U23389 ( .C1(n20462), .C2(n20727), .A(n20602), .B(n20461), .ZN(
        n20463) );
  OAI211_X1 U23390 ( .C1(n20602), .C2(n20464), .A(n20606), .B(n20463), .ZN(
        n20484) );
  AOI22_X1 U23391 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20484), .B1(
        n20483), .B2(n20558), .ZN(n20465) );
  OAI211_X1 U23392 ( .C1(n20561), .C2(n20518), .A(n20466), .B(n20465), .ZN(
        P1_U3121) );
  AOI22_X1 U23393 ( .A1(n20612), .A2(n20482), .B1(n20481), .B2(n20613), .ZN(
        n20468) );
  INV_X1 U23394 ( .A(n20518), .ZN(n20475) );
  AOI22_X1 U23395 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20484), .B1(
        n20475), .B2(n20614), .ZN(n20467) );
  OAI211_X1 U23396 ( .C1(n20617), .C2(n20478), .A(n20468), .B(n20467), .ZN(
        P1_U3122) );
  AOI22_X1 U23397 ( .A1(n20618), .A2(n20482), .B1(n20481), .B2(n20619), .ZN(
        n20470) );
  AOI22_X1 U23398 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20484), .B1(
        n20475), .B2(n20620), .ZN(n20469) );
  OAI211_X1 U23399 ( .C1(n20623), .C2(n20478), .A(n20470), .B(n20469), .ZN(
        P1_U3123) );
  AOI22_X1 U23400 ( .A1(n20624), .A2(n20482), .B1(n20481), .B2(n20625), .ZN(
        n20472) );
  AOI22_X1 U23401 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20484), .B1(
        n20475), .B2(n20626), .ZN(n20471) );
  OAI211_X1 U23402 ( .C1(n20629), .C2(n20478), .A(n20472), .B(n20471), .ZN(
        P1_U3124) );
  AOI22_X1 U23403 ( .A1(n20630), .A2(n20482), .B1(n20481), .B2(n20631), .ZN(
        n20474) );
  AOI22_X1 U23404 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20484), .B1(
        n20475), .B2(n20632), .ZN(n20473) );
  OAI211_X1 U23405 ( .C1(n20635), .C2(n20478), .A(n20474), .B(n20473), .ZN(
        P1_U3125) );
  AOI22_X1 U23406 ( .A1(n20636), .A2(n20482), .B1(n20481), .B2(n20637), .ZN(
        n20477) );
  AOI22_X1 U23407 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20484), .B1(
        n20475), .B2(n20638), .ZN(n20476) );
  OAI211_X1 U23408 ( .C1(n20641), .C2(n20478), .A(n20477), .B(n20476), .ZN(
        P1_U3126) );
  AOI22_X1 U23409 ( .A1(n20642), .A2(n20482), .B1(n20481), .B2(n20643), .ZN(
        n20480) );
  AOI22_X1 U23410 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20484), .B1(
        n20483), .B2(n20582), .ZN(n20479) );
  OAI211_X1 U23411 ( .C1(n20585), .C2(n20518), .A(n20480), .B(n20479), .ZN(
        P1_U3127) );
  AOI22_X1 U23412 ( .A1(n20649), .A2(n20482), .B1(n20481), .B2(n20650), .ZN(
        n20486) );
  AOI22_X1 U23413 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20484), .B1(
        n20483), .B2(n20588), .ZN(n20485) );
  OAI211_X1 U23414 ( .C1(n20593), .C2(n20518), .A(n20486), .B(n20485), .ZN(
        P1_U3128) );
  NOR3_X1 U23415 ( .A1(n20488), .A2(n20738), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20524) );
  INV_X1 U23416 ( .A(n20524), .ZN(n20521) );
  NOR2_X1 U23417 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20521), .ZN(
        n20512) );
  AOI22_X1 U23418 ( .A1(n20513), .A2(n20608), .B1(n20600), .B2(n20512), .ZN(
        n20499) );
  NAND2_X1 U23419 ( .A1(n20518), .A2(n20545), .ZN(n20489) );
  AOI21_X1 U23420 ( .B1(n20489), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20728), 
        .ZN(n20494) );
  NAND2_X1 U23421 ( .A1(n20594), .A2(n13348), .ZN(n20496) );
  AOI22_X1 U23422 ( .A1(n20494), .A2(n20496), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20495), .ZN(n20492) );
  OAI211_X1 U23423 ( .C1(n20512), .C2(n20493), .A(n20556), .B(n20492), .ZN(
        n20515) );
  INV_X1 U23424 ( .A(n20494), .ZN(n20497) );
  AOI22_X1 U23425 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20515), .B1(
        n20601), .B2(n20514), .ZN(n20498) );
  OAI211_X1 U23426 ( .C1(n20611), .C2(n20518), .A(n20499), .B(n20498), .ZN(
        P1_U3129) );
  AOI22_X1 U23427 ( .A1(n20513), .A2(n20614), .B1(n20612), .B2(n20512), .ZN(
        n20501) );
  AOI22_X1 U23428 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20515), .B1(
        n20613), .B2(n20514), .ZN(n20500) );
  OAI211_X1 U23429 ( .C1(n20617), .C2(n20518), .A(n20501), .B(n20500), .ZN(
        P1_U3130) );
  AOI22_X1 U23430 ( .A1(n20513), .A2(n20620), .B1(n20618), .B2(n20512), .ZN(
        n20503) );
  AOI22_X1 U23431 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20515), .B1(
        n20619), .B2(n20514), .ZN(n20502) );
  OAI211_X1 U23432 ( .C1(n20623), .C2(n20518), .A(n20503), .B(n20502), .ZN(
        P1_U3131) );
  AOI22_X1 U23433 ( .A1(n20513), .A2(n20626), .B1(n20624), .B2(n20512), .ZN(
        n20505) );
  AOI22_X1 U23434 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20515), .B1(
        n20625), .B2(n20514), .ZN(n20504) );
  OAI211_X1 U23435 ( .C1(n20629), .C2(n20518), .A(n20505), .B(n20504), .ZN(
        P1_U3132) );
  AOI22_X1 U23436 ( .A1(n20513), .A2(n20632), .B1(n20630), .B2(n20512), .ZN(
        n20507) );
  AOI22_X1 U23437 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20515), .B1(
        n20631), .B2(n20514), .ZN(n20506) );
  OAI211_X1 U23438 ( .C1(n20635), .C2(n20518), .A(n20507), .B(n20506), .ZN(
        P1_U3133) );
  AOI22_X1 U23439 ( .A1(n20513), .A2(n20638), .B1(n20636), .B2(n20512), .ZN(
        n20509) );
  AOI22_X1 U23440 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20515), .B1(
        n20637), .B2(n20514), .ZN(n20508) );
  OAI211_X1 U23441 ( .C1(n20641), .C2(n20518), .A(n20509), .B(n20508), .ZN(
        P1_U3134) );
  AOI22_X1 U23442 ( .A1(n20513), .A2(n20644), .B1(n20642), .B2(n20512), .ZN(
        n20511) );
  AOI22_X1 U23443 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20515), .B1(
        n20643), .B2(n20514), .ZN(n20510) );
  OAI211_X1 U23444 ( .C1(n20647), .C2(n20518), .A(n20511), .B(n20510), .ZN(
        P1_U3135) );
  AOI22_X1 U23445 ( .A1(n20513), .A2(n20652), .B1(n20649), .B2(n20512), .ZN(
        n20517) );
  AOI22_X1 U23446 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20515), .B1(
        n20650), .B2(n20514), .ZN(n20516) );
  OAI211_X1 U23447 ( .C1(n20658), .C2(n20518), .A(n20517), .B(n20516), .ZN(
        P1_U3136) );
  NOR2_X1 U23448 ( .A1(n20519), .A2(n20521), .ZN(n20541) );
  AOI21_X1 U23449 ( .B1(n20594), .B2(n20520), .A(n20541), .ZN(n20522) );
  OAI22_X1 U23450 ( .A1(n20522), .A2(n20728), .B1(n20521), .B2(n20752), .ZN(
        n20540) );
  AOI22_X1 U23451 ( .A1(n20600), .A2(n20541), .B1(n20601), .B2(n20540), .ZN(
        n20527) );
  NOR3_X1 U23452 ( .A1(n20603), .A2(n20728), .A3(n20753), .ZN(n20523) );
  OAI21_X1 U23453 ( .B1(n20524), .B2(n20523), .A(n20606), .ZN(n20542) );
  NOR2_X2 U23454 ( .A1(n20603), .A2(n20525), .ZN(n20589) );
  AOI22_X1 U23455 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20542), .B1(
        n20589), .B2(n20608), .ZN(n20526) );
  OAI211_X1 U23456 ( .C1(n20611), .C2(n20545), .A(n20527), .B(n20526), .ZN(
        P1_U3137) );
  AOI22_X1 U23457 ( .A1(n20612), .A2(n20541), .B1(n20613), .B2(n20540), .ZN(
        n20529) );
  AOI22_X1 U23458 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20542), .B1(
        n20589), .B2(n20614), .ZN(n20528) );
  OAI211_X1 U23459 ( .C1(n20617), .C2(n20545), .A(n20529), .B(n20528), .ZN(
        P1_U3138) );
  AOI22_X1 U23460 ( .A1(n20618), .A2(n20541), .B1(n20619), .B2(n20540), .ZN(
        n20531) );
  AOI22_X1 U23461 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20542), .B1(
        n20589), .B2(n20620), .ZN(n20530) );
  OAI211_X1 U23462 ( .C1(n20623), .C2(n20545), .A(n20531), .B(n20530), .ZN(
        P1_U3139) );
  AOI22_X1 U23463 ( .A1(n20624), .A2(n20541), .B1(n20625), .B2(n20540), .ZN(
        n20533) );
  AOI22_X1 U23464 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20542), .B1(
        n20589), .B2(n20626), .ZN(n20532) );
  OAI211_X1 U23465 ( .C1(n20629), .C2(n20545), .A(n20533), .B(n20532), .ZN(
        P1_U3140) );
  AOI22_X1 U23466 ( .A1(n20630), .A2(n20541), .B1(n20631), .B2(n20540), .ZN(
        n20535) );
  AOI22_X1 U23467 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20542), .B1(
        n20589), .B2(n20632), .ZN(n20534) );
  OAI211_X1 U23468 ( .C1(n20635), .C2(n20545), .A(n20535), .B(n20534), .ZN(
        P1_U3141) );
  AOI22_X1 U23469 ( .A1(n20636), .A2(n20541), .B1(n20637), .B2(n20540), .ZN(
        n20537) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20542), .B1(
        n20589), .B2(n20638), .ZN(n20536) );
  OAI211_X1 U23471 ( .C1(n20641), .C2(n20545), .A(n20537), .B(n20536), .ZN(
        P1_U3142) );
  AOI22_X1 U23472 ( .A1(n20642), .A2(n20541), .B1(n20643), .B2(n20540), .ZN(
        n20539) );
  AOI22_X1 U23473 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20542), .B1(
        n20589), .B2(n20644), .ZN(n20538) );
  OAI211_X1 U23474 ( .C1(n20647), .C2(n20545), .A(n20539), .B(n20538), .ZN(
        P1_U3143) );
  AOI22_X1 U23475 ( .A1(n20649), .A2(n20541), .B1(n20650), .B2(n20540), .ZN(
        n20544) );
  AOI22_X1 U23476 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20542), .B1(
        n20589), .B2(n20652), .ZN(n20543) );
  OAI211_X1 U23477 ( .C1(n20658), .C2(n20545), .A(n20544), .B(n20543), .ZN(
        P1_U3144) );
  INV_X1 U23478 ( .A(n20603), .ZN(n20547) );
  NOR2_X1 U23479 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20604), .ZN(
        n20587) );
  NAND3_X1 U23480 ( .A1(n20594), .A2(n20553), .A3(n20602), .ZN(n20548) );
  OAI21_X1 U23481 ( .B1(n20550), .B2(n20549), .A(n20548), .ZN(n20586) );
  AOI22_X1 U23482 ( .A1(n20600), .A2(n20587), .B1(n20601), .B2(n20586), .ZN(
        n20560) );
  NOR3_X1 U23483 ( .A1(n20753), .A2(n20603), .A3(n20551), .ZN(n20552) );
  AOI21_X1 U23484 ( .B1(n20594), .B2(n20553), .A(n20552), .ZN(n20554) );
  NOR2_X1 U23485 ( .A1(n20554), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20557) );
  AOI22_X1 U23486 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20558), .ZN(n20559) );
  OAI211_X1 U23487 ( .C1(n20561), .C2(n20657), .A(n20560), .B(n20559), .ZN(
        P1_U3145) );
  AOI22_X1 U23488 ( .A1(n20612), .A2(n20587), .B1(n20613), .B2(n20586), .ZN(
        n20564) );
  AOI22_X1 U23489 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20562), .ZN(n20563) );
  OAI211_X1 U23490 ( .C1(n20565), .C2(n20657), .A(n20564), .B(n20563), .ZN(
        P1_U3146) );
  AOI22_X1 U23491 ( .A1(n20618), .A2(n20587), .B1(n20619), .B2(n20586), .ZN(
        n20568) );
  AOI22_X1 U23492 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20566), .ZN(n20567) );
  OAI211_X1 U23493 ( .C1(n20569), .C2(n20657), .A(n20568), .B(n20567), .ZN(
        P1_U3147) );
  AOI22_X1 U23494 ( .A1(n20624), .A2(n20587), .B1(n20625), .B2(n20586), .ZN(
        n20572) );
  AOI22_X1 U23495 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20570), .ZN(n20571) );
  OAI211_X1 U23496 ( .C1(n20573), .C2(n20657), .A(n20572), .B(n20571), .ZN(
        P1_U3148) );
  AOI22_X1 U23497 ( .A1(n20630), .A2(n20587), .B1(n20631), .B2(n20586), .ZN(
        n20576) );
  AOI22_X1 U23498 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20574), .ZN(n20575) );
  OAI211_X1 U23499 ( .C1(n20577), .C2(n20657), .A(n20576), .B(n20575), .ZN(
        P1_U3149) );
  AOI22_X1 U23500 ( .A1(n20636), .A2(n20587), .B1(n20637), .B2(n20586), .ZN(
        n20580) );
  AOI22_X1 U23501 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20578), .ZN(n20579) );
  OAI211_X1 U23502 ( .C1(n20581), .C2(n20657), .A(n20580), .B(n20579), .ZN(
        P1_U3150) );
  AOI22_X1 U23503 ( .A1(n20642), .A2(n20587), .B1(n20643), .B2(n20586), .ZN(
        n20584) );
  AOI22_X1 U23504 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20582), .ZN(n20583) );
  OAI211_X1 U23505 ( .C1(n20585), .C2(n20657), .A(n20584), .B(n20583), .ZN(
        P1_U3151) );
  AOI22_X1 U23506 ( .A1(n20649), .A2(n20587), .B1(n20650), .B2(n20586), .ZN(
        n20592) );
  AOI22_X1 U23507 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20590), .B1(
        n20589), .B2(n20588), .ZN(n20591) );
  OAI211_X1 U23508 ( .C1(n20593), .C2(n20657), .A(n20592), .B(n20591), .ZN(
        P1_U3152) );
  INV_X1 U23509 ( .A(n20594), .ZN(n20598) );
  INV_X1 U23510 ( .A(n20595), .ZN(n20597) );
  INV_X1 U23511 ( .A(n20648), .ZN(n20596) );
  OAI21_X1 U23512 ( .B1(n20598), .B2(n20597), .A(n20596), .ZN(n20607) );
  INV_X1 U23513 ( .A(n20607), .ZN(n20599) );
  OAI22_X1 U23514 ( .A1(n20599), .A2(n20728), .B1(n20604), .B2(n20752), .ZN(
        n20651) );
  AOI22_X1 U23515 ( .A1(n20651), .A2(n20601), .B1(n20600), .B2(n20648), .ZN(
        n20610) );
  OAI21_X1 U23516 ( .B1(n20603), .B2(n20727), .A(n20602), .ZN(n20731) );
  NAND2_X1 U23517 ( .A1(n20604), .A2(n20728), .ZN(n20605) );
  OAI211_X1 U23518 ( .C1(n20731), .C2(n20607), .A(n20606), .B(n20605), .ZN(
        n20654) );
  AOI22_X1 U23519 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20608), .ZN(n20609) );
  OAI211_X1 U23520 ( .C1(n20611), .C2(n20657), .A(n20610), .B(n20609), .ZN(
        P1_U3153) );
  AOI22_X1 U23521 ( .A1(n20651), .A2(n20613), .B1(n20612), .B2(n20648), .ZN(
        n20616) );
  AOI22_X1 U23522 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20614), .ZN(n20615) );
  OAI211_X1 U23523 ( .C1(n20617), .C2(n20657), .A(n20616), .B(n20615), .ZN(
        P1_U3154) );
  AOI22_X1 U23524 ( .A1(n20651), .A2(n20619), .B1(n20618), .B2(n20648), .ZN(
        n20622) );
  AOI22_X1 U23525 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20620), .ZN(n20621) );
  OAI211_X1 U23526 ( .C1(n20623), .C2(n20657), .A(n20622), .B(n20621), .ZN(
        P1_U3155) );
  AOI22_X1 U23527 ( .A1(n20651), .A2(n20625), .B1(n20624), .B2(n20648), .ZN(
        n20628) );
  AOI22_X1 U23528 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20626), .ZN(n20627) );
  OAI211_X1 U23529 ( .C1(n20629), .C2(n20657), .A(n20628), .B(n20627), .ZN(
        P1_U3156) );
  AOI22_X1 U23530 ( .A1(n20651), .A2(n20631), .B1(n20630), .B2(n20648), .ZN(
        n20634) );
  AOI22_X1 U23531 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20632), .ZN(n20633) );
  OAI211_X1 U23532 ( .C1(n20635), .C2(n20657), .A(n20634), .B(n20633), .ZN(
        P1_U3157) );
  AOI22_X1 U23533 ( .A1(n20651), .A2(n20637), .B1(n20636), .B2(n20648), .ZN(
        n20640) );
  AOI22_X1 U23534 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20638), .ZN(n20639) );
  OAI211_X1 U23535 ( .C1(n20641), .C2(n20657), .A(n20640), .B(n20639), .ZN(
        P1_U3158) );
  AOI22_X1 U23536 ( .A1(n20651), .A2(n20643), .B1(n20642), .B2(n20648), .ZN(
        n20646) );
  AOI22_X1 U23537 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20644), .ZN(n20645) );
  OAI211_X1 U23538 ( .C1(n20647), .C2(n20657), .A(n20646), .B(n20645), .ZN(
        P1_U3159) );
  AOI22_X1 U23539 ( .A1(n20651), .A2(n20650), .B1(n20649), .B2(n20648), .ZN(
        n20656) );
  AOI22_X1 U23540 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20654), .B1(
        n20653), .B2(n20652), .ZN(n20655) );
  OAI211_X1 U23541 ( .C1(n20658), .C2(n20657), .A(n20656), .B(n20655), .ZN(
        P1_U3160) );
  AOI21_X1 U23542 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20756), .A(n20659), 
        .ZN(n20661) );
  NAND2_X1 U23543 ( .A1(n20661), .A2(n20660), .ZN(P1_U3163) );
  AND2_X1 U23544 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20662), .ZN(
        P1_U3164) );
  AND2_X1 U23545 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20662), .ZN(
        P1_U3165) );
  AND2_X1 U23546 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20662), .ZN(
        P1_U3166) );
  AND2_X1 U23547 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20662), .ZN(
        P1_U3167) );
  AND2_X1 U23548 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20662), .ZN(
        P1_U3168) );
  AND2_X1 U23549 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20662), .ZN(
        P1_U3169) );
  AND2_X1 U23550 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20662), .ZN(
        P1_U3170) );
  AND2_X1 U23551 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20662), .ZN(
        P1_U3171) );
  AND2_X1 U23552 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20662), .ZN(
        P1_U3172) );
  AND2_X1 U23553 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20662), .ZN(
        P1_U3173) );
  AND2_X1 U23554 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20662), .ZN(
        P1_U3174) );
  AND2_X1 U23555 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20662), .ZN(
        P1_U3175) );
  AND2_X1 U23556 ( .A1(n20662), .A2(P1_DATAWIDTH_REG_19__SCAN_IN), .ZN(
        P1_U3176) );
  AND2_X1 U23557 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20662), .ZN(
        P1_U3177) );
  AND2_X1 U23558 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20662), .ZN(
        P1_U3178) );
  AND2_X1 U23559 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20662), .ZN(
        P1_U3179) );
  AND2_X1 U23560 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20662), .ZN(
        P1_U3180) );
  AND2_X1 U23561 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20662), .ZN(
        P1_U3181) );
  AND2_X1 U23562 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20662), .ZN(
        P1_U3182) );
  AND2_X1 U23563 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20662), .ZN(
        P1_U3183) );
  AND2_X1 U23564 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20662), .ZN(
        P1_U3184) );
  AND2_X1 U23565 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20662), .ZN(
        P1_U3185) );
  AND2_X1 U23566 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(n20662), .ZN(P1_U3186) );
  AND2_X1 U23567 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20662), .ZN(P1_U3187) );
  AND2_X1 U23568 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20662), .ZN(P1_U3188) );
  AND2_X1 U23569 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20662), .ZN(P1_U3189) );
  AND2_X1 U23570 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20662), .ZN(P1_U3190) );
  AND2_X1 U23571 ( .A1(n20662), .A2(P1_DATAWIDTH_REG_4__SCAN_IN), .ZN(P1_U3191) );
  AND2_X1 U23572 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20662), .ZN(P1_U3192) );
  AND2_X1 U23573 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20662), .ZN(P1_U3193) );
  NAND2_X1 U23574 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20669), .ZN(n20675) );
  INV_X1 U23575 ( .A(n20675), .ZN(n20667) );
  NAND2_X1 U23576 ( .A1(n20663), .A2(n11618), .ZN(n20665) );
  NAND2_X1 U23577 ( .A1(n20676), .A2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n20668) );
  AOI22_X1 U23578 ( .A1(HOLD), .A2(n20665), .B1(n20668), .B2(n20664), .ZN(
        n20666) );
  OAI22_X1 U23579 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20667), .B1(n20750), 
        .B2(n20666), .ZN(P1_U3194) );
  INV_X1 U23580 ( .A(n20668), .ZN(n20673) );
  INV_X1 U23581 ( .A(n20669), .ZN(n20672) );
  AOI21_X1 U23582 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n11618), .A(n20670), .ZN(n20671) );
  AOI21_X1 U23583 ( .B1(n20673), .B2(n20672), .A(n20671), .ZN(n20680) );
  NAND3_X1 U23584 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20674), .A3(n20676), 
        .ZN(n20678) );
  OAI211_X1 U23585 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n20676), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20675), .ZN(n20677) );
  OAI221_X1 U23586 ( .B1(n20680), .B2(n20679), .C1(n20680), .C2(n20678), .A(
        n20677), .ZN(P1_U3196) );
  OR2_X1 U23587 ( .A1(n20748), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20706) );
  INV_X1 U23588 ( .A(P1_ADDRESS_REG_0__SCAN_IN), .ZN(n20801) );
  OR2_X1 U23589 ( .A1(n11618), .A2(n20748), .ZN(n20703) );
  OAI222_X1 U23590 ( .A1(n20706), .A2(n20682), .B1(n20801), .B2(n20750), .C1(
        n20740), .C2(n20703), .ZN(P1_U3197) );
  OAI222_X1 U23591 ( .A1(n20703), .A2(n20682), .B1(n20681), .B2(n20750), .C1(
        n20684), .C2(n20706), .ZN(P1_U3198) );
  INV_X1 U23592 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20826) );
  OAI222_X1 U23593 ( .A1(n20703), .A2(n20684), .B1(n20826), .B2(n20750), .C1(
        n20683), .C2(n20706), .ZN(P1_U3199) );
  INV_X1 U23594 ( .A(n20703), .ZN(n20717) );
  AOI222_X1 U23595 ( .A1(n20716), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20748), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20717), .ZN(n20685) );
  INV_X1 U23596 ( .A(n20685), .ZN(P1_U3200) );
  AOI222_X1 U23597 ( .A1(n20717), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20748), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20716), .ZN(n20686) );
  INV_X1 U23598 ( .A(n20686), .ZN(P1_U3201) );
  AOI222_X1 U23599 ( .A1(n20717), .A2(P1_REIP_REG_6__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20748), .C1(P1_REIP_REG_7__SCAN_IN), 
        .C2(n20716), .ZN(n20687) );
  INV_X1 U23600 ( .A(n20687), .ZN(P1_U3202) );
  AOI222_X1 U23601 ( .A1(n20717), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_6__SCAN_IN), .B2(n20748), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20716), .ZN(n20688) );
  INV_X1 U23602 ( .A(n20688), .ZN(P1_U3203) );
  AOI222_X1 U23603 ( .A1(n20717), .A2(P1_REIP_REG_8__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20748), .C1(P1_REIP_REG_9__SCAN_IN), 
        .C2(n20716), .ZN(n20689) );
  INV_X1 U23604 ( .A(n20689), .ZN(P1_U3204) );
  AOI222_X1 U23605 ( .A1(n20717), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20748), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20716), .ZN(n20690) );
  INV_X1 U23606 ( .A(n20690), .ZN(P1_U3205) );
  AOI222_X1 U23607 ( .A1(n20717), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20748), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n20716), .ZN(n20691) );
  INV_X1 U23608 ( .A(n20691), .ZN(P1_U3206) );
  AOI222_X1 U23609 ( .A1(n20717), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20748), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20716), .ZN(n20692) );
  INV_X1 U23610 ( .A(n20692), .ZN(P1_U3207) );
  AOI222_X1 U23611 ( .A1(n20716), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20748), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20717), .ZN(n20693) );
  INV_X1 U23612 ( .A(n20693), .ZN(P1_U3208) );
  AOI222_X1 U23613 ( .A1(n20717), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20748), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20716), .ZN(n20694) );
  INV_X1 U23614 ( .A(n20694), .ZN(P1_U3209) );
  AOI22_X1 U23615 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20748), .B1(
        P1_REIP_REG_15__SCAN_IN), .B2(n20716), .ZN(n20695) );
  OAI21_X1 U23616 ( .B1(n20696), .B2(n20703), .A(n20695), .ZN(P1_U3210) );
  AOI22_X1 U23617 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(n20748), .B1(
        P1_REIP_REG_15__SCAN_IN), .B2(n20717), .ZN(n20697) );
  OAI21_X1 U23618 ( .B1(n20830), .B2(n20706), .A(n20697), .ZN(P1_U3211) );
  AOI222_X1 U23619 ( .A1(n20716), .A2(P1_REIP_REG_17__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n20748), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20717), .ZN(n20698) );
  INV_X1 U23620 ( .A(n20698), .ZN(P1_U3212) );
  AOI222_X1 U23621 ( .A1(n20717), .A2(P1_REIP_REG_17__SCAN_IN), .B1(
        P1_ADDRESS_REG_16__SCAN_IN), .B2(n20748), .C1(P1_REIP_REG_18__SCAN_IN), 
        .C2(n20716), .ZN(n20699) );
  INV_X1 U23622 ( .A(n20699), .ZN(P1_U3213) );
  AOI222_X1 U23623 ( .A1(n20717), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20748), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20716), .ZN(n20700) );
  INV_X1 U23624 ( .A(n20700), .ZN(P1_U3214) );
  AOI222_X1 U23625 ( .A1(n20716), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20748), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20717), .ZN(n20701) );
  INV_X1 U23626 ( .A(n20701), .ZN(P1_U3215) );
  AOI22_X1 U23627 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(n20748), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(n20716), .ZN(n20702) );
  OAI21_X1 U23628 ( .B1(n20704), .B2(n20703), .A(n20702), .ZN(P1_U3216) );
  AOI22_X1 U23629 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(n20748), .B1(
        P1_REIP_REG_21__SCAN_IN), .B2(n20717), .ZN(n20705) );
  OAI21_X1 U23630 ( .B1(n20707), .B2(n20706), .A(n20705), .ZN(P1_U3217) );
  AOI222_X1 U23631 ( .A1(n20717), .A2(P1_REIP_REG_22__SCAN_IN), .B1(
        P1_ADDRESS_REG_21__SCAN_IN), .B2(n20748), .C1(P1_REIP_REG_23__SCAN_IN), 
        .C2(n20716), .ZN(n20708) );
  INV_X1 U23632 ( .A(n20708), .ZN(P1_U3218) );
  AOI222_X1 U23633 ( .A1(n20717), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20748), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n20716), .ZN(n20709) );
  INV_X1 U23634 ( .A(n20709), .ZN(P1_U3219) );
  AOI222_X1 U23635 ( .A1(n20717), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20748), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20716), .ZN(n20710) );
  INV_X1 U23636 ( .A(n20710), .ZN(P1_U3220) );
  AOI222_X1 U23637 ( .A1(n20717), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20748), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20716), .ZN(n20711) );
  INV_X1 U23638 ( .A(n20711), .ZN(P1_U3221) );
  AOI222_X1 U23639 ( .A1(n20717), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20748), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20716), .ZN(n20712) );
  INV_X1 U23640 ( .A(n20712), .ZN(P1_U3222) );
  AOI222_X1 U23641 ( .A1(n20717), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20748), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20716), .ZN(n20713) );
  INV_X1 U23642 ( .A(n20713), .ZN(P1_U3223) );
  AOI222_X1 U23643 ( .A1(n20717), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20748), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20716), .ZN(n20714) );
  INV_X1 U23644 ( .A(n20714), .ZN(P1_U3224) );
  AOI222_X1 U23645 ( .A1(n20717), .A2(P1_REIP_REG_29__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20748), .C1(P1_REIP_REG_30__SCAN_IN), 
        .C2(n20716), .ZN(n20715) );
  INV_X1 U23646 ( .A(n20715), .ZN(P1_U3225) );
  AOI222_X1 U23647 ( .A1(n20717), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20748), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20716), .ZN(n20718) );
  INV_X1 U23648 ( .A(n20718), .ZN(P1_U3226) );
  OAI22_X1 U23649 ( .A1(n20748), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20750), .ZN(n20719) );
  INV_X1 U23650 ( .A(n20719), .ZN(P1_U3458) );
  OAI22_X1 U23651 ( .A1(n20748), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20750), .ZN(n20720) );
  INV_X1 U23652 ( .A(n20720), .ZN(P1_U3459) );
  OAI22_X1 U23653 ( .A1(n20748), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20750), .ZN(n20721) );
  INV_X1 U23654 ( .A(n20721), .ZN(P1_U3460) );
  OAI22_X1 U23655 ( .A1(n20748), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20750), .ZN(n20722) );
  INV_X1 U23656 ( .A(n20722), .ZN(P1_U3461) );
  OAI21_X1 U23657 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20726), .A(n20724), 
        .ZN(n20723) );
  INV_X1 U23658 ( .A(n20723), .ZN(P1_U3464) );
  OAI21_X1 U23659 ( .B1(n20726), .B2(n20725), .A(n20724), .ZN(P1_U3465) );
  INV_X1 U23660 ( .A(n20736), .ZN(n20739) );
  NOR3_X1 U23661 ( .A1(n20729), .A2(n20728), .A3(n20727), .ZN(n20733) );
  NOR2_X1 U23662 ( .A1(n20731), .A2(n20730), .ZN(n20732) );
  AOI211_X1 U23663 ( .C1(n20735), .C2(n20734), .A(n20733), .B(n20732), .ZN(
        n20737) );
  AOI22_X1 U23664 ( .A1(n20739), .A2(n20738), .B1(n20737), .B2(n20736), .ZN(
        P1_U3475) );
  AOI21_X1 U23665 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20741) );
  AOI22_X1 U23666 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20741), .B2(n20740), .ZN(n20744) );
  INV_X1 U23667 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20743) );
  AOI22_X1 U23668 ( .A1(n20747), .A2(n20744), .B1(n20743), .B2(n20742), .ZN(
        P1_U3481) );
  INV_X1 U23669 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20746) );
  OAI21_X1 U23670 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20747), .ZN(n20745) );
  OAI21_X1 U23671 ( .B1(n20747), .B2(n20746), .A(n20745), .ZN(P1_U3482) );
  INV_X1 U23672 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20749) );
  AOI22_X1 U23673 ( .A1(n20750), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20749), 
        .B2(n20748), .ZN(P1_U3483) );
  AOI211_X1 U23674 ( .C1(n20754), .C2(n20753), .A(n20752), .B(n20751), .ZN(
        n20757) );
  OAI21_X1 U23675 ( .B1(n20757), .B2(n20756), .A(n20755), .ZN(n20763) );
  AOI211_X1 U23676 ( .C1(n20761), .C2(n20760), .A(n20759), .B(n20758), .ZN(
        n20762) );
  MUX2_X1 U23677 ( .A(n20763), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n20762), 
        .Z(P1_U3485) );
  MUX2_X1 U23678 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n20748), .Z(P1_U3486) );
  NAND2_X1 U23679 ( .A1(keyinput34), .A2(keyinput0), .ZN(n20770) );
  NOR2_X1 U23680 ( .A1(keyinput49), .A2(keyinput40), .ZN(n20768) );
  NAND3_X1 U23681 ( .A1(keyinput32), .A2(keyinput57), .A3(keyinput25), .ZN(
        n20766) );
  INV_X1 U23682 ( .A(keyinput21), .ZN(n20764) );
  NAND3_X1 U23683 ( .A1(keyinput55), .A2(keyinput18), .A3(n20764), .ZN(n20765)
         );
  NOR4_X1 U23684 ( .A1(keyinput58), .A2(keyinput23), .A3(n20766), .A4(n20765), 
        .ZN(n20767) );
  NAND4_X1 U23685 ( .A1(keyinput8), .A2(keyinput28), .A3(n20768), .A4(n20767), 
        .ZN(n20769) );
  NOR4_X1 U23686 ( .A1(keyinput11), .A2(keyinput60), .A3(n20770), .A4(n20769), 
        .ZN(n20924) );
  NAND4_X1 U23687 ( .A1(keyinput12), .A2(keyinput16), .A3(keyinput13), .A4(
        keyinput61), .ZN(n20789) );
  NOR3_X1 U23688 ( .A1(keyinput14), .A2(keyinput2), .A3(keyinput41), .ZN(
        n20774) );
  NAND3_X1 U23689 ( .A1(keyinput47), .A2(keyinput51), .A3(keyinput36), .ZN(
        n20772) );
  NAND3_X1 U23690 ( .A1(keyinput44), .A2(keyinput35), .A3(keyinput20), .ZN(
        n20771) );
  NOR4_X1 U23691 ( .A1(keyinput24), .A2(keyinput43), .A3(n20772), .A4(n20771), 
        .ZN(n20773) );
  NAND3_X1 U23692 ( .A1(keyinput29), .A2(n20774), .A3(n20773), .ZN(n20788) );
  NOR2_X1 U23693 ( .A1(keyinput22), .A2(keyinput4), .ZN(n20779) );
  NAND4_X1 U23694 ( .A1(keyinput42), .A2(keyinput7), .A3(keyinput59), .A4(
        keyinput33), .ZN(n20777) );
  NAND3_X1 U23695 ( .A1(keyinput26), .A2(keyinput52), .A3(keyinput1), .ZN(
        n20776) );
  NAND4_X1 U23696 ( .A1(keyinput30), .A2(keyinput31), .A3(keyinput5), .A4(
        keyinput6), .ZN(n20775) );
  NOR4_X1 U23697 ( .A1(keyinput38), .A2(n20777), .A3(n20776), .A4(n20775), 
        .ZN(n20778) );
  NAND4_X1 U23698 ( .A1(keyinput9), .A2(keyinput27), .A3(n20779), .A4(n20778), 
        .ZN(n20787) );
  NOR2_X1 U23699 ( .A1(keyinput15), .A2(keyinput54), .ZN(n20785) );
  NAND3_X1 U23700 ( .A1(keyinput45), .A2(keyinput19), .A3(keyinput37), .ZN(
        n20783) );
  NOR2_X1 U23701 ( .A1(keyinput50), .A2(keyinput63), .ZN(n20781) );
  NOR4_X1 U23702 ( .A1(keyinput62), .A2(keyinput17), .A3(keyinput46), .A4(
        keyinput39), .ZN(n20780) );
  NAND4_X1 U23703 ( .A1(keyinput56), .A2(keyinput10), .A3(n20781), .A4(n20780), 
        .ZN(n20782) );
  NOR3_X1 U23704 ( .A1(keyinput48), .A2(n20783), .A3(n20782), .ZN(n20784) );
  NAND4_X1 U23705 ( .A1(keyinput53), .A2(keyinput3), .A3(n20785), .A4(n20784), 
        .ZN(n20786) );
  NOR4_X1 U23706 ( .A1(n20789), .A2(n20788), .A3(n20787), .A4(n20786), .ZN(
        n20923) );
  INV_X1 U23707 ( .A(keyinput14), .ZN(n20791) );
  AOI22_X1 U23708 ( .A1(n20792), .A2(keyinput29), .B1(
        P2_DATAWIDTH_REG_11__SCAN_IN), .B2(n20791), .ZN(n20790) );
  OAI221_X1 U23709 ( .B1(n20792), .B2(keyinput29), .C1(n20791), .C2(
        P2_DATAWIDTH_REG_11__SCAN_IN), .A(n20790), .ZN(n20805) );
  AOI22_X1 U23710 ( .A1(n20795), .A2(keyinput2), .B1(n20794), .B2(keyinput41), 
        .ZN(n20793) );
  OAI221_X1 U23711 ( .B1(n20795), .B2(keyinput2), .C1(n20794), .C2(keyinput41), 
        .A(n20793), .ZN(n20804) );
  INV_X1 U23712 ( .A(P2_UWORD_REG_14__SCAN_IN), .ZN(n20798) );
  INV_X1 U23713 ( .A(P1_LWORD_REG_6__SCAN_IN), .ZN(n20797) );
  AOI22_X1 U23714 ( .A1(n20798), .A2(keyinput47), .B1(n20797), .B2(keyinput51), 
        .ZN(n20796) );
  OAI221_X1 U23715 ( .B1(n20798), .B2(keyinput47), .C1(n20797), .C2(keyinput51), .A(n20796), .ZN(n20803) );
  AOI22_X1 U23716 ( .A1(n20801), .A2(keyinput36), .B1(n20800), .B2(keyinput24), 
        .ZN(n20799) );
  OAI221_X1 U23717 ( .B1(n20801), .B2(keyinput36), .C1(n20800), .C2(keyinput24), .A(n20799), .ZN(n20802) );
  NOR4_X1 U23718 ( .A1(n20805), .A2(n20804), .A3(n20803), .A4(n20802), .ZN(
        n20854) );
  AOI22_X1 U23719 ( .A1(n20808), .A2(keyinput12), .B1(n20807), .B2(keyinput16), 
        .ZN(n20806) );
  OAI221_X1 U23720 ( .B1(n20808), .B2(keyinput12), .C1(n20807), .C2(keyinput16), .A(n20806), .ZN(n20820) );
  AOI22_X1 U23721 ( .A1(n20811), .A2(keyinput13), .B1(keyinput61), .B2(n20810), 
        .ZN(n20809) );
  OAI221_X1 U23722 ( .B1(n20811), .B2(keyinput13), .C1(n20810), .C2(keyinput61), .A(n20809), .ZN(n20819) );
  INV_X1 U23723 ( .A(keyinput44), .ZN(n20813) );
  AOI22_X1 U23724 ( .A1(n10980), .A2(keyinput35), .B1(
        P3_ADDRESS_REG_16__SCAN_IN), .B2(n20813), .ZN(n20812) );
  OAI221_X1 U23725 ( .B1(n10980), .B2(keyinput35), .C1(n20813), .C2(
        P3_ADDRESS_REG_16__SCAN_IN), .A(n20812), .ZN(n20818) );
  INV_X1 U23726 ( .A(keyinput20), .ZN(n20815) );
  AOI22_X1 U23727 ( .A1(n20816), .A2(keyinput43), .B1(
        P3_DATAWIDTH_REG_11__SCAN_IN), .B2(n20815), .ZN(n20814) );
  OAI221_X1 U23728 ( .B1(n20816), .B2(keyinput43), .C1(n20815), .C2(
        P3_DATAWIDTH_REG_11__SCAN_IN), .A(n20814), .ZN(n20817) );
  NOR4_X1 U23729 ( .A1(n20820), .A2(n20819), .A3(n20818), .A4(n20817), .ZN(
        n20853) );
  INV_X1 U23730 ( .A(P3_DATAO_REG_16__SCAN_IN), .ZN(n20823) );
  INV_X1 U23731 ( .A(keyinput9), .ZN(n20822) );
  AOI22_X1 U23732 ( .A1(n20823), .A2(keyinput22), .B1(
        P1_DATAWIDTH_REG_4__SCAN_IN), .B2(n20822), .ZN(n20821) );
  OAI221_X1 U23733 ( .B1(n20823), .B2(keyinput22), .C1(n20822), .C2(
        P1_DATAWIDTH_REG_4__SCAN_IN), .A(n20821), .ZN(n20836) );
  AOI22_X1 U23734 ( .A1(n20826), .A2(keyinput59), .B1(n20825), .B2(keyinput33), 
        .ZN(n20824) );
  OAI221_X1 U23735 ( .B1(n20826), .B2(keyinput59), .C1(n20825), .C2(keyinput33), .A(n20824), .ZN(n20835) );
  AOI22_X1 U23736 ( .A1(n20829), .A2(keyinput27), .B1(keyinput4), .B2(n20828), 
        .ZN(n20827) );
  OAI221_X1 U23737 ( .B1(n20829), .B2(keyinput27), .C1(n20828), .C2(keyinput4), 
        .A(n20827), .ZN(n20834) );
  XOR2_X1 U23738 ( .A(n20830), .B(keyinput42), .Z(n20832) );
  XNOR2_X1 U23739 ( .A(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B(keyinput7), .ZN(
        n20831) );
  NAND2_X1 U23740 ( .A1(n20832), .A2(n20831), .ZN(n20833) );
  NOR4_X1 U23741 ( .A1(n20836), .A2(n20835), .A3(n20834), .A4(n20833), .ZN(
        n20852) );
  INV_X1 U23742 ( .A(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n20838) );
  AOI22_X1 U23743 ( .A1(n20839), .A2(keyinput26), .B1(n20838), .B2(keyinput52), 
        .ZN(n20837) );
  OAI221_X1 U23744 ( .B1(n20839), .B2(keyinput26), .C1(n20838), .C2(keyinput52), .A(n20837), .ZN(n20850) );
  INV_X1 U23745 ( .A(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n20841) );
  AOI22_X1 U23746 ( .A1(n10268), .A2(keyinput1), .B1(keyinput38), .B2(n20841), 
        .ZN(n20840) );
  OAI221_X1 U23747 ( .B1(n10268), .B2(keyinput1), .C1(n20841), .C2(keyinput38), 
        .A(n20840), .ZN(n20849) );
  AOI22_X1 U23748 ( .A1(n20843), .A2(keyinput30), .B1(n13245), .B2(keyinput31), 
        .ZN(n20842) );
  OAI221_X1 U23749 ( .B1(n20843), .B2(keyinput30), .C1(n13245), .C2(keyinput31), .A(n20842), .ZN(n20848) );
  INV_X1 U23750 ( .A(DATAI_0_), .ZN(n20846) );
  INV_X1 U23751 ( .A(keyinput5), .ZN(n20845) );
  AOI22_X1 U23752 ( .A1(n20846), .A2(keyinput6), .B1(P3_DATAO_REG_15__SCAN_IN), 
        .B2(n20845), .ZN(n20844) );
  OAI221_X1 U23753 ( .B1(n20846), .B2(keyinput6), .C1(n20845), .C2(
        P3_DATAO_REG_15__SCAN_IN), .A(n20844), .ZN(n20847) );
  NOR4_X1 U23754 ( .A1(n20850), .A2(n20849), .A3(n20848), .A4(n20847), .ZN(
        n20851) );
  NAND4_X1 U23755 ( .A1(n20854), .A2(n20853), .A3(n20852), .A4(n20851), .ZN(
        n20922) );
  INV_X1 U23756 ( .A(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n20857) );
  INV_X1 U23757 ( .A(P3_EBX_REG_14__SCAN_IN), .ZN(n20856) );
  AOI22_X1 U23758 ( .A1(n20857), .A2(keyinput10), .B1(keyinput63), .B2(n20856), 
        .ZN(n20855) );
  OAI221_X1 U23759 ( .B1(n20857), .B2(keyinput10), .C1(n20856), .C2(keyinput63), .A(n20855), .ZN(n20870) );
  INV_X1 U23760 ( .A(P3_UWORD_REG_6__SCAN_IN), .ZN(n20860) );
  INV_X1 U23761 ( .A(keyinput56), .ZN(n20859) );
  AOI22_X1 U23762 ( .A1(n20860), .A2(keyinput50), .B1(
        P3_ADDRESS_REG_18__SCAN_IN), .B2(n20859), .ZN(n20858) );
  OAI221_X1 U23763 ( .B1(n20860), .B2(keyinput50), .C1(n20859), .C2(
        P3_ADDRESS_REG_18__SCAN_IN), .A(n20858), .ZN(n20869) );
  INV_X1 U23764 ( .A(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n20863) );
  AOI22_X1 U23765 ( .A1(n20863), .A2(keyinput46), .B1(keyinput39), .B2(n20862), 
        .ZN(n20861) );
  OAI221_X1 U23766 ( .B1(n20863), .B2(keyinput46), .C1(n20862), .C2(keyinput39), .A(n20861), .ZN(n20868) );
  INV_X1 U23767 ( .A(keyinput62), .ZN(n20865) );
  AOI22_X1 U23768 ( .A1(n20866), .A2(keyinput17), .B1(
        P1_DATAWIDTH_REG_19__SCAN_IN), .B2(n20865), .ZN(n20864) );
  OAI221_X1 U23769 ( .B1(n20866), .B2(keyinput17), .C1(n20865), .C2(
        P1_DATAWIDTH_REG_19__SCAN_IN), .A(n20864), .ZN(n20867) );
  NOR4_X1 U23770 ( .A1(n20870), .A2(n20869), .A3(n20868), .A4(n20867), .ZN(
        n20920) );
  INV_X1 U23771 ( .A(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n20873) );
  INV_X1 U23772 ( .A(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n20872) );
  AOI22_X1 U23773 ( .A1(n20873), .A2(keyinput53), .B1(keyinput3), .B2(n20872), 
        .ZN(n20871) );
  OAI221_X1 U23774 ( .B1(n20873), .B2(keyinput53), .C1(n20872), .C2(keyinput3), 
        .A(n20871), .ZN(n20885) );
  INV_X1 U23775 ( .A(keyinput15), .ZN(n20875) );
  AOI22_X1 U23776 ( .A1(n15140), .A2(keyinput54), .B1(
        P3_ADDRESS_REG_29__SCAN_IN), .B2(n20875), .ZN(n20874) );
  OAI221_X1 U23777 ( .B1(n15140), .B2(keyinput54), .C1(n20875), .C2(
        P3_ADDRESS_REG_29__SCAN_IN), .A(n20874), .ZN(n20884) );
  AOI22_X1 U23778 ( .A1(n20878), .A2(keyinput48), .B1(n20877), .B2(keyinput37), 
        .ZN(n20876) );
  OAI221_X1 U23779 ( .B1(n20878), .B2(keyinput48), .C1(n20877), .C2(keyinput37), .A(n20876), .ZN(n20883) );
  INV_X1 U23780 ( .A(P1_UWORD_REG_6__SCAN_IN), .ZN(n20880) );
  AOI22_X1 U23781 ( .A1(n20881), .A2(keyinput45), .B1(n20880), .B2(keyinput19), 
        .ZN(n20879) );
  OAI221_X1 U23782 ( .B1(n20881), .B2(keyinput45), .C1(n20880), .C2(keyinput19), .A(n20879), .ZN(n20882) );
  NOR4_X1 U23783 ( .A1(n20885), .A2(n20884), .A3(n20883), .A4(n20882), .ZN(
        n20919) );
  INV_X1 U23784 ( .A(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n20888) );
  INV_X1 U23785 ( .A(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n20887) );
  AOI22_X1 U23786 ( .A1(n20888), .A2(keyinput32), .B1(n20887), .B2(keyinput57), 
        .ZN(n20886) );
  OAI221_X1 U23787 ( .B1(n20888), .B2(keyinput32), .C1(n20887), .C2(keyinput57), .A(n20886), .ZN(n20900) );
  INV_X1 U23788 ( .A(P1_UWORD_REG_11__SCAN_IN), .ZN(n20890) );
  AOI22_X1 U23789 ( .A1(n20891), .A2(keyinput23), .B1(keyinput21), .B2(n20890), 
        .ZN(n20889) );
  OAI221_X1 U23790 ( .B1(n20891), .B2(keyinput23), .C1(n20890), .C2(keyinput21), .A(n20889), .ZN(n20899) );
  INV_X1 U23791 ( .A(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n20893) );
  AOI22_X1 U23792 ( .A1(n13121), .A2(keyinput25), .B1(n20893), .B2(keyinput58), 
        .ZN(n20892) );
  OAI221_X1 U23793 ( .B1(n13121), .B2(keyinput25), .C1(n20893), .C2(keyinput58), .A(n20892), .ZN(n20898) );
  INV_X1 U23794 ( .A(keyinput18), .ZN(n20894) );
  XOR2_X1 U23795 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .B(n20894), .Z(n20896) );
  XNOR2_X1 U23796 ( .A(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B(keyinput55), .ZN(
        n20895) );
  NAND2_X1 U23797 ( .A1(n20896), .A2(n20895), .ZN(n20897) );
  NOR4_X1 U23798 ( .A1(n20900), .A2(n20899), .A3(n20898), .A4(n20897), .ZN(
        n20918) );
  INV_X1 U23799 ( .A(P1_UWORD_REG_13__SCAN_IN), .ZN(n20903) );
  INV_X1 U23800 ( .A(keyinput60), .ZN(n20902) );
  AOI22_X1 U23801 ( .A1(n20903), .A2(keyinput0), .B1(
        P3_DATAWIDTH_REG_14__SCAN_IN), .B2(n20902), .ZN(n20901) );
  OAI221_X1 U23802 ( .B1(n20903), .B2(keyinput0), .C1(n20902), .C2(
        P3_DATAWIDTH_REG_14__SCAN_IN), .A(n20901), .ZN(n20916) );
  AOI22_X1 U23803 ( .A1(n20906), .A2(keyinput34), .B1(n20905), .B2(keyinput11), 
        .ZN(n20904) );
  OAI221_X1 U23804 ( .B1(n20906), .B2(keyinput34), .C1(n20905), .C2(keyinput11), .A(n20904), .ZN(n20915) );
  INV_X1 U23805 ( .A(P2_UWORD_REG_9__SCAN_IN), .ZN(n20909) );
  AOI22_X1 U23806 ( .A1(n20909), .A2(keyinput49), .B1(n20908), .B2(keyinput40), 
        .ZN(n20907) );
  OAI221_X1 U23807 ( .B1(n20909), .B2(keyinput49), .C1(n20908), .C2(keyinput40), .A(n20907), .ZN(n20914) );
  INV_X1 U23808 ( .A(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n20912) );
  INV_X1 U23809 ( .A(P1_UWORD_REG_7__SCAN_IN), .ZN(n20911) );
  AOI22_X1 U23810 ( .A1(n20912), .A2(keyinput8), .B1(keyinput28), .B2(n20911), 
        .ZN(n20910) );
  OAI221_X1 U23811 ( .B1(n20912), .B2(keyinput8), .C1(n20911), .C2(keyinput28), 
        .A(n20910), .ZN(n20913) );
  NOR4_X1 U23812 ( .A1(n20916), .A2(n20915), .A3(n20914), .A4(n20913), .ZN(
        n20917) );
  NAND4_X1 U23813 ( .A1(n20920), .A2(n20919), .A3(n20918), .A4(n20917), .ZN(
        n20921) );
  AOI211_X1 U23814 ( .C1(n20924), .C2(n20923), .A(n20922), .B(n20921), .ZN(
        n20929) );
  AOI222_X1 U23815 ( .A1(BUF1_REG_12__SCAN_IN), .A2(n20927), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n20926), .C1(P2_DATAO_REG_12__SCAN_IN), 
        .C2(n20925), .ZN(n20928) );
  XNOR2_X1 U23816 ( .A(n20929), .B(n20928), .ZN(U235) );
  AND2_X1 U12300 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n11235) );
  AND2_X2 U12363 ( .A1(n11125), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n11190) );
  NOR2_X2 U12347 ( .A1(n11223), .A2(n11224), .ZN(n11222) );
  NOR2_X2 U11219 ( .A1(n16184), .A2(n16185), .ZN(n16183) );
  NOR2_X2 U11557 ( .A1(n18877), .A2(n18878), .ZN(n18876) );
  NOR2_X2 U14336 ( .A1(n16207), .A2(n16205), .ZN(n16206) );
  NOR2_X2 U14337 ( .A1(n9698), .A2(n15085), .ZN(n15084) );
  CLKBUF_X2 U11174 ( .A(n11492), .Z(n9608) );
  NAND2_X1 U11153 ( .A1(n10174), .A2(n10175), .ZN(n14014) );
  OAI211_X1 U13118 ( .C1(n10224), .C2(n19822), .A(n10223), .B(n10222), .ZN(
        n10245) );
  OR3_X1 U12304 ( .A1(n11207), .A2(n9850), .A3(n11202), .ZN(n9656) );
  INV_X1 U11146 ( .A(n18605), .ZN(n18631) );
  CLKBUF_X1 U11036 ( .A(n11738), .Z(n11653) );
  CLKBUF_X1 U11063 ( .A(n13394), .Z(n11762) );
  NOR2_X2 U11083 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13948) );
  CLKBUF_X1 U11108 ( .A(n11547), .Z(n12341) );
  OR2_X2 U11112 ( .A1(n13497), .A2(n19822), .ZN(n10748) );
  NAND2_X1 U11114 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18786), .ZN(
        n11289) );
  NOR2_X2 U11140 ( .A1(n19809), .A2(n10848), .ZN(n10199) );
  CLKBUF_X1 U11150 ( .A(n11398), .Z(n9600) );
  NOR2_X1 U11209 ( .A1(n16195), .A2(n16196), .ZN(n16194) );
  AND4_X1 U11345 ( .A1(n11123), .A2(n9642), .A3(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A4(n11234), .ZN(n11227) );
  CLKBUF_X1 U11556 ( .A(n11773), .Z(n9621) );
  AND2_X1 U11640 ( .A1(n9837), .A2(n15222), .ZN(n16165) );
  NOR2_X1 U11641 ( .A1(n13066), .A2(n15229), .ZN(n13065) );
  NOR2_X1 U12051 ( .A1(n15271), .A2(n13052), .ZN(n13051) );
  INV_X1 U12205 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n19822) );
  INV_X1 U12241 ( .A(n17808), .ZN(n17531) );
  CLKBUF_X1 U12340 ( .A(n16064), .Z(n9595) );
  CLKBUF_X1 U12349 ( .A(n16497), .Z(n16507) );
  CLKBUF_X1 U12429 ( .A(n18807), .Z(n17410) );
endmodule

