

module b14_C_gen_AntiSAT_k_128_8 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, 
        U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, 
        U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, 
        U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, 
        U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, 
        U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, 
        U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, 
        U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, 
        U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, 
        U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, 
        U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, 
        U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, 
        U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, 
        U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, 
        U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, 
        U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, 
        U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, 
        U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, 
        U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, 
        U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, 
        U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, 
        U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, 
        U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, 
        U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, 
        U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722;

  CLKBUF_X2 U2285 ( .A(n2964), .Z(n3680) );
  XNOR2_X1 U2286 ( .A(n2318), .B(IR_REG_2__SCAN_IN), .ZN(n4366) );
  NAND2_X1 U2287 ( .A1(n2654), .A2(n2244), .ZN(n2759) );
  INV_X1 U2288 ( .A(IR_REG_5__SCAN_IN), .ZN(n2353) );
  INV_X1 U2289 ( .A(IR_REG_6__SCAN_IN), .ZN(n2366) );
  NOR2_X1 U2290 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2272)
         );
  INV_X1 U2292 ( .A(n2068), .ZN(n3675) );
  INV_X2 U2293 ( .A(n2312), .ZN(n3409) );
  NOR2_X1 U2294 ( .A1(n2811), .A2(n3103), .ZN(n2816) );
  NOR2_X1 U2295 ( .A1(n2816), .A2(n2101), .ZN(n2877) );
  AND2_X1 U2296 ( .A1(n3225), .A2(n3275), .ZN(n3169) );
  AND2_X1 U2297 ( .A1(n2510), .A2(n2076), .ZN(n2275) );
  INV_X1 U2298 ( .A(IR_REG_7__SCAN_IN), .ZN(n2405) );
  INV_X1 U2299 ( .A(IR_REG_31__SCAN_IN), .ZN(n2378) );
  AND2_X1 U2300 ( .A1(n2668), .A2(n2053), .ZN(n2752) );
  XNOR2_X2 U2301 ( .A(n2617), .B(n2616), .ZN(n2623) );
  NAND2_X2 U2302 ( .A1(n2615), .A2(IR_REG_31__SCAN_IN), .ZN(n2617) );
  NOR2_X1 U2303 ( .A1(n4449), .A2(REG1_REG_16__SCAN_IN), .ZN(n4450) );
  NAND2_X1 U2304 ( .A1(n3744), .A2(n3743), .ZN(n3742) );
  AND2_X1 U2305 ( .A1(n3753), .A2(n3755), .ZN(n3630) );
  OR2_X1 U2306 ( .A1(n3632), .A2(n3631), .ZN(n3633) );
  NOR2_X1 U2307 ( .A1(n2102), .A2(n2139), .ZN(n2101) );
  AND2_X2 U2308 ( .A1(n2741), .A2(n4476), .ZN(n4367) );
  INV_X1 U2309 ( .A(n2103), .ZN(n2102) );
  OR2_X1 U2310 ( .A1(n2782), .A2(n2781), .ZN(n2142) );
  INV_X2 U2311 ( .A(n2887), .ZN(n2958) );
  NAND2_X1 U2312 ( .A1(n2807), .A2(n2104), .ZN(n2103) );
  INV_X4 U2313 ( .A(n3682), .ZN(n2960) );
  INV_X2 U2314 ( .A(n2068), .ZN(n2043) );
  OR2_X1 U2315 ( .A1(n3459), .A2(n2651), .ZN(n2843) );
  NAND2_X2 U2316 ( .A1(n2288), .A2(n2756), .ZN(n2311) );
  INV_X1 U2317 ( .A(n2752), .ZN(n2764) );
  NAND2_X1 U2318 ( .A1(n4358), .A2(n2284), .ZN(n2312) );
  INV_X2 U2319 ( .A(n2319), .ZN(n2333) );
  XNOR2_X1 U2320 ( .A(n2282), .B(IR_REG_30__SCAN_IN), .ZN(n4358) );
  XNOR2_X1 U2321 ( .A(n2612), .B(n2611), .ZN(n3459) );
  NAND2_X1 U2322 ( .A1(n2759), .A2(IR_REG_31__SCAN_IN), .ZN(n2282) );
  NOR2_X1 U2323 ( .A1(n2518), .A2(IR_REG_18__SCAN_IN), .ZN(n2610) );
  NOR2_X1 U2324 ( .A1(IR_REG_4__SCAN_IN), .A2(IR_REG_3__SCAN_IN), .ZN(n2106)
         );
  INV_X1 U2325 ( .A(IR_REG_8__SCAN_IN), .ZN(n2388) );
  NOR2_X1 U2326 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2270)
         );
  NOR2_X1 U2327 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2273)
         );
  NOR2_X2 U2328 ( .A1(n4009), .A2(n3689), .ZN(n2719) );
  OR2_X2 U2329 ( .A1(n4031), .A2(n3713), .ZN(n4009) );
  MUX2_X1 U2330 ( .A(n2711), .B(n2710), .S(IR_REG_28__SCAN_IN), .Z(n2044) );
  MUX2_X1 U2331 ( .A(n2711), .B(n2710), .S(IR_REG_28__SCAN_IN), .Z(n2045) );
  INV_X4 U2332 ( .A(n2333), .ZN(n2512) );
  NAND2_X1 U2333 ( .A1(n2829), .A2(n2841), .ZN(n2887) );
  NAND2_X1 U2334 ( .A1(n2654), .A2(n2280), .ZN(n2283) );
  OR2_X1 U2335 ( .A1(n2311), .A2(n2295), .ZN(n2299) );
  NOR2_X1 U2336 ( .A1(n3874), .A2(n2229), .ZN(n2228) );
  OR2_X1 U2337 ( .A1(n3515), .A2(n2411), .ZN(n2413) );
  NAND2_X1 U2338 ( .A1(n2902), .A2(n3034), .ZN(n3501) );
  NAND2_X1 U2339 ( .A1(n2321), .A2(n2320), .ZN(n3007) );
  INV_X1 U2340 ( .A(n2759), .ZN(n2192) );
  NAND4_X1 U2341 ( .A1(n2388), .A2(n2366), .A3(n2353), .A4(n2405), .ZN(n2258)
         );
  OR2_X1 U2342 ( .A1(n2580), .A2(n2579), .ZN(n2598) );
  NAND2_X1 U2343 ( .A1(n3610), .A2(n2213), .ZN(n2215) );
  AND2_X1 U2344 ( .A1(n3886), .A2(n3800), .ZN(n2213) );
  OR2_X1 U2345 ( .A1(n2964), .A2(n2902), .ZN(n2108) );
  NAND2_X1 U2346 ( .A1(n2933), .A2(n2136), .ZN(n2135) );
  NAND2_X1 U2347 ( .A1(n4366), .A2(REG2_REG_2__SCAN_IN), .ZN(n2136) );
  INV_X1 U2348 ( .A(n4510), .ZN(n3958) );
  NAND2_X1 U2349 ( .A1(n4372), .A2(n4373), .ZN(n4371) );
  NAND2_X1 U2350 ( .A1(n4392), .A2(n4393), .ZN(n4391) );
  NAND2_X1 U2351 ( .A1(n3907), .A2(n3782), .ZN(n2450) );
  AOI21_X1 U2352 ( .B1(n2715), .B2(n4203), .A(n2252), .ZN(n3996) );
  INV_X1 U2353 ( .A(n4203), .ZN(n4159) );
  INV_X1 U2354 ( .A(IR_REG_28__SCAN_IN), .ZN(n2280) );
  AND2_X1 U2355 ( .A1(n2132), .A2(n2276), .ZN(n2131) );
  INV_X1 U2356 ( .A(IR_REG_20__SCAN_IN), .ZN(n2616) );
  NOR2_X1 U2357 ( .A1(n4460), .A2(n3977), .ZN(n4471) );
  NAND2_X1 U2358 ( .A1(n4471), .A2(n4472), .ZN(n4469) );
  AND2_X1 U2359 ( .A1(n2391), .A2(n3162), .ZN(n2409) );
  INV_X1 U2360 ( .A(n2650), .ZN(n3538) );
  OR2_X1 U2361 ( .A1(n3538), .A2(n3447), .ZN(n2129) );
  INV_X1 U2362 ( .A(n2187), .ZN(n2182) );
  INV_X1 U2363 ( .A(n2577), .ZN(n2185) );
  INV_X1 U2364 ( .A(n2488), .ZN(n2196) );
  NAND2_X1 U2365 ( .A1(n2487), .A2(n2486), .ZN(n2488) );
  INV_X1 U2366 ( .A(n3490), .ZN(n2115) );
  NAND2_X1 U2367 ( .A1(n3490), .A2(n2114), .ZN(n2113) );
  INV_X1 U2368 ( .A(n3517), .ZN(n2118) );
  INV_X1 U2369 ( .A(IR_REG_26__SCAN_IN), .ZN(n2200) );
  INV_X1 U2370 ( .A(IR_REG_17__SCAN_IN), .ZN(n2509) );
  INV_X1 U2371 ( .A(n2254), .ZN(n2208) );
  NOR2_X1 U2372 ( .A1(n3187), .A2(n3186), .ZN(n2212) );
  NAND2_X1 U2373 ( .A1(n3187), .A2(n3186), .ZN(n2211) );
  INV_X1 U2374 ( .A(n2212), .ZN(n2210) );
  NOR2_X1 U2375 ( .A1(n2225), .A2(n2224), .ZN(n2223) );
  INV_X1 U2376 ( .A(n3822), .ZN(n2224) );
  NAND2_X1 U2377 ( .A1(n3875), .A2(n2230), .ZN(n2226) );
  AND2_X1 U2378 ( .A1(n3599), .A2(n3598), .ZN(n3720) );
  AOI21_X1 U2379 ( .B1(n2243), .B2(n3575), .A(n2240), .ZN(n2239) );
  NOR2_X1 U2380 ( .A1(n3370), .A2(n2241), .ZN(n2240) );
  AND2_X1 U2381 ( .A1(n3586), .A2(n3585), .ZN(n3777) );
  NOR2_X1 U2382 ( .A1(n3656), .A2(n3658), .ZN(n3654) );
  NAND2_X1 U2383 ( .A1(n2548), .A2(REG3_REG_23__SCAN_IN), .ZN(n2558) );
  INV_X1 U2384 ( .A(n2550), .ZN(n2548) );
  OR2_X1 U2385 ( .A1(n2558), .A2(n4698), .ZN(n2570) );
  NAND2_X1 U2386 ( .A1(n2959), .A2(n3660), .ZN(n2962) );
  NOR2_X1 U2387 ( .A1(n3575), .A2(n3576), .ZN(n2242) );
  NAND2_X1 U2388 ( .A1(n2239), .A2(n3776), .ZN(n2235) );
  INV_X1 U2389 ( .A(n3777), .ZN(n2238) );
  NAND2_X1 U2390 ( .A1(n3828), .A2(n2204), .ZN(n2203) );
  OAI22_X1 U2391 ( .A1(n2902), .A2(n2887), .B1(n2842), .B2(n3682), .ZN(n2845)
         );
  AND2_X1 U2392 ( .A1(n2592), .A2(n2591), .ZN(n3674) );
  AND2_X1 U2393 ( .A1(n2081), .A2(n2080), .ZN(n2782) );
  NAND2_X1 U2394 ( .A1(n2054), .A2(n4364), .ZN(n2081) );
  XNOR2_X1 U2395 ( .A(n2103), .B(n4363), .ZN(n2811) );
  OR2_X1 U2396 ( .A1(n2879), .A2(n2093), .ZN(n2092) );
  AND2_X1 U2397 ( .A1(n4362), .A2(REG2_REG_7__SCAN_IN), .ZN(n2093) );
  NAND2_X1 U2398 ( .A1(n4371), .A2(n3962), .ZN(n3964) );
  NAND2_X1 U2399 ( .A1(n4383), .A2(REG2_REG_10__SCAN_IN), .ZN(n4382) );
  NAND2_X1 U2400 ( .A1(n4391), .A2(n3966), .ZN(n3968) );
  NAND2_X1 U2401 ( .A1(n4394), .A2(n3945), .ZN(n3946) );
  NAND2_X1 U2402 ( .A1(n4403), .A2(REG2_REG_12__SCAN_IN), .ZN(n4402) );
  OAI21_X1 U2403 ( .B1(n4415), .B2(n4411), .A(n2137), .ZN(n3948) );
  OR2_X1 U2404 ( .A1(n3956), .A2(REG2_REG_13__SCAN_IN), .ZN(n2137) );
  NAND2_X1 U2405 ( .A1(n4438), .A2(n3973), .ZN(n3975) );
  NOR2_X1 U2406 ( .A1(n4433), .A2(n2094), .ZN(n3951) );
  AND2_X1 U2407 ( .A1(n3955), .A2(REG2_REG_15__SCAN_IN), .ZN(n2094) );
  NAND2_X1 U2408 ( .A1(n4454), .A2(n2148), .ZN(n2147) );
  NAND2_X1 U2409 ( .A1(n4463), .A2(n2491), .ZN(n2148) );
  NAND2_X1 U2410 ( .A1(n2719), .A2(n3994), .ZN(n4215) );
  NOR2_X1 U2411 ( .A1(n2127), .A2(n4005), .ZN(n2126) );
  INV_X1 U2412 ( .A(n3544), .ZN(n2127) );
  AOI21_X1 U2413 ( .B1(n4110), .B2(n2536), .A(n2535), .ZN(n4101) );
  AND2_X1 U2414 ( .A1(n4133), .A2(n4115), .ZN(n2535) );
  NAND2_X1 U2415 ( .A1(n2160), .A2(n2047), .ZN(n2158) );
  NAND2_X1 U2416 ( .A1(n2047), .A2(n2256), .ZN(n2159) );
  AND2_X1 U2417 ( .A1(n4294), .A2(n3616), .ZN(n2498) );
  NAND2_X1 U2418 ( .A1(n4206), .A2(n4205), .ZN(n4204) );
  INV_X1 U2419 ( .A(n4205), .ZN(n2197) );
  NAND2_X1 U2420 ( .A1(n3261), .A2(n2488), .ZN(n2198) );
  AND2_X1 U2421 ( .A1(n3429), .A2(n3493), .ZN(n4205) );
  AND2_X1 U2422 ( .A1(n2245), .A2(n2066), .ZN(n2165) );
  NAND2_X1 U2423 ( .A1(n2164), .A2(n2162), .ZN(n3200) );
  NOR2_X1 U2424 ( .A1(n2163), .A2(n2462), .ZN(n2162) );
  OR2_X1 U2425 ( .A1(n2416), .A2(n2172), .ZN(n2170) );
  AND2_X1 U2426 ( .A1(n2167), .A2(n2174), .ZN(n2171) );
  NAND2_X1 U2427 ( .A1(n2176), .A2(n2175), .ZN(n2180) );
  INV_X1 U2428 ( .A(n2427), .ZN(n2175) );
  INV_X1 U2429 ( .A(n3168), .ZN(n2176) );
  AND2_X1 U2430 ( .A1(n3295), .A2(n3297), .ZN(n3455) );
  OAI21_X1 U2431 ( .B1(n3058), .B2(n3054), .A(n3487), .ZN(n3083) );
  AOI21_X1 U2432 ( .B1(n3007), .B2(n2335), .A(n2255), .ZN(n2992) );
  OR2_X1 U2433 ( .A1(n2992), .A2(n2994), .ZN(n3056) );
  NAND2_X1 U2434 ( .A1(n2301), .A2(REG1_REG_0__SCAN_IN), .ZN(n2307) );
  OR2_X1 U2435 ( .A1(n2303), .A2(n2309), .ZN(n2316) );
  AND2_X1 U2436 ( .A1(n2586), .A2(n2585), .ZN(n4237) );
  INV_X1 U2437 ( .A(n3909), .ZN(n3308) );
  AND4_X1 U2438 ( .A1(n2435), .A2(n2434), .A3(n2433), .A4(n2432), .ZN(n3745)
         );
  INV_X1 U2439 ( .A(n3747), .ZN(n3365) );
  INV_X1 U2440 ( .A(n3911), .ZN(n3238) );
  NAND2_X1 U2441 ( .A1(n2652), .A2(n3443), .ZN(n4203) );
  NAND2_X1 U2442 ( .A1(n2752), .A2(n2676), .ZN(n2763) );
  NAND2_X1 U2443 ( .A1(n2841), .A2(n4497), .ZN(n2860) );
  NAND2_X1 U2444 ( .A1(n2190), .A2(n2189), .ZN(n2284) );
  NAND2_X1 U2445 ( .A1(n2283), .A2(n2057), .ZN(n2189) );
  AOI21_X1 U2446 ( .B1(IR_REG_22__SCAN_IN), .B2(IR_REG_31__SCAN_IN), .A(
        IR_REG_23__SCAN_IN), .ZN(n2219) );
  NOR2_X2 U2447 ( .A1(n2618), .A2(IR_REG_21__SCAN_IN), .ZN(n2673) );
  INV_X1 U2448 ( .A(IR_REG_9__SCAN_IN), .ZN(n2259) );
  NAND2_X1 U2449 ( .A1(n3840), .A2(n3842), .ZN(n3590) );
  OAI21_X1 U2450 ( .B1(n3840), .B2(n3842), .A(n3841), .ZN(n3589) );
  NAND2_X1 U2451 ( .A1(n2851), .A2(n2068), .ZN(n2854) );
  CLKBUF_X1 U2452 ( .A(n2892), .Z(n2857) );
  AND2_X1 U2453 ( .A1(n2538), .A2(n2529), .ZN(n4117) );
  INV_X1 U2454 ( .A(n3884), .ZN(n3897) );
  NAND2_X1 U2455 ( .A1(n2576), .A2(n2575), .ZN(n4063) );
  OR2_X1 U2456 ( .A1(n3793), .A2(n2658), .ZN(n2576) );
  INV_X1 U2457 ( .A(n4050), .ZN(n4234) );
  INV_X1 U2458 ( .A(n4156), .ZN(n4284) );
  INV_X1 U2459 ( .A(n4287), .ZN(n3904) );
  INV_X1 U2460 ( .A(n3593), .ZN(n3905) );
  OR2_X1 U2461 ( .A1(n2149), .A2(n2775), .ZN(n2088) );
  NAND2_X1 U2462 ( .A1(n4395), .A2(n4396), .ZN(n4394) );
  XNOR2_X1 U2463 ( .A(n3968), .B(n4506), .ZN(n4408) );
  XNOR2_X1 U2464 ( .A(n3975), .B(n3974), .ZN(n4449) );
  NAND2_X1 U2465 ( .A1(n2146), .A2(n4413), .ZN(n2145) );
  NAND2_X1 U2466 ( .A1(n2147), .A2(n4466), .ZN(n2146) );
  AOI21_X1 U2467 ( .B1(n4468), .B2(ADDR_REG_18__SCAN_IN), .A(n4467), .ZN(n2144) );
  NOR2_X1 U2468 ( .A1(n2147), .A2(n4466), .ZN(n4465) );
  XNOR2_X1 U2469 ( .A(n2098), .B(n3979), .ZN(n3984) );
  NAND2_X1 U2470 ( .A1(n4469), .A2(n2070), .ZN(n2098) );
  AND2_X1 U2471 ( .A1(n3923), .A2(n3918), .ZN(n4470) );
  NOR2_X1 U2472 ( .A1(n4465), .A2(n2097), .ZN(n2096) );
  AND2_X1 U2473 ( .A1(n3954), .A2(REG2_REG_18__SCAN_IN), .ZN(n2097) );
  INV_X1 U2474 ( .A(DATAI_1_), .ZN(n2153) );
  AND2_X1 U2475 ( .A1(n3996), .A2(n2130), .ZN(n2724) );
  AOI21_X1 U2476 ( .B1(n3992), .B2(n4521), .A(n2717), .ZN(n2130) );
  INV_X2 U2477 ( .A(n4527), .ZN(n4529) );
  XNOR2_X1 U2478 ( .A(n2614), .B(IR_REG_19__SCAN_IN), .ZN(n4360) );
  XNOR2_X1 U2479 ( .A(n2089), .B(IR_REG_1__SCAN_IN), .ZN(n2149) );
  NAND2_X1 U2480 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2089)
         );
  INV_X1 U2481 ( .A(n3680), .ZN(n3669) );
  AND2_X1 U2482 ( .A1(n2251), .A2(n3493), .ZN(n2116) );
  NOR2_X1 U2483 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2271)
         );
  NOR2_X1 U2484 ( .A1(n2528), .A2(n3766), .ZN(n2537) );
  NAND2_X1 U2485 ( .A1(n2960), .A2(n3069), .ZN(n2964) );
  AND2_X1 U2486 ( .A1(n2463), .A2(REG3_REG_15__SCAN_IN), .ZN(n2285) );
  NOR2_X1 U2487 ( .A1(n2501), .A2(n2500), .ZN(n2513) );
  INV_X1 U2488 ( .A(n2417), .ZN(n2168) );
  AOI21_X1 U2489 ( .B1(n2177), .B2(n2427), .A(n2063), .ZN(n2174) );
  NOR2_X1 U2490 ( .A1(n2430), .A2(n2429), .ZN(n2428) );
  NAND2_X1 U2491 ( .A1(n3169), .A2(n3365), .ZN(n3170) );
  NAND2_X1 U2492 ( .A1(n2977), .A2(n2979), .ZN(n2978) );
  INV_X1 U2493 ( .A(IR_REG_27__SCAN_IN), .ZN(n2276) );
  NOR2_X1 U2494 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2266)
         );
  NOR2_X1 U2495 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2264)
         );
  NOR2_X1 U2496 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2265)
         );
  INV_X1 U2497 ( .A(n2258), .ZN(n2232) );
  OR3_X1 U2498 ( .A1(n2436), .A2(IR_REG_12__SCAN_IN), .A3(n2260), .ZN(n2459)
         );
  INV_X1 U2499 ( .A(IR_REG_2__SCAN_IN), .ZN(n2107) );
  NAND2_X1 U2500 ( .A1(n2537), .A2(REG3_REG_22__SCAN_IN), .ZN(n2550) );
  NAND2_X1 U2501 ( .A1(n2073), .A2(n2072), .ZN(n3011) );
  OR2_X1 U2502 ( .A1(n2333), .A2(n2797), .ZN(n2073) );
  NAND2_X1 U2503 ( .A1(n2333), .A2(DATAI_3_), .ZN(n2072) );
  AND2_X1 U2504 ( .A1(n2253), .A2(n3615), .ZN(n2214) );
  INV_X2 U2505 ( .A(n2958), .ZN(n3683) );
  INV_X1 U2506 ( .A(n4140), .ZN(n4131) );
  NAND2_X1 U2507 ( .A1(n2428), .A2(REG3_REG_12__SCAN_IN), .ZN(n2453) );
  OR2_X1 U2508 ( .A1(n2453), .A2(n2452), .ZN(n2464) );
  NOR2_X1 U2509 ( .A1(n3853), .A2(n2202), .ZN(n2201) );
  INV_X1 U2510 ( .A(n3641), .ZN(n2202) );
  OAI21_X1 U2511 ( .B1(n3605), .B2(n3720), .A(n3607), .ZN(n3886) );
  AND4_X1 U2512 ( .A1(n2495), .A2(n2494), .A3(n2493), .A4(n2492), .ZN(n4294)
         );
  NAND2_X1 U2513 ( .A1(n2133), .A2(n4364), .ZN(n2085) );
  NAND2_X1 U2514 ( .A1(n2142), .A2(n2141), .ZN(n2140) );
  NAND2_X1 U2515 ( .A1(n2105), .A2(REG2_REG_5__SCAN_IN), .ZN(n2141) );
  NAND2_X1 U2516 ( .A1(n2105), .A2(REG1_REG_5__SCAN_IN), .ZN(n2104) );
  AOI21_X1 U2517 ( .B1(n2819), .B2(REG2_REG_6__SCAN_IN), .A(n2138), .ZN(n2821)
         );
  AND2_X1 U2518 ( .A1(n2140), .A2(n4363), .ZN(n2138) );
  NOR2_X1 U2519 ( .A1(n2821), .A2(n2820), .ZN(n2879) );
  XNOR2_X1 U2520 ( .A(n2092), .B(n2091), .ZN(n3941) );
  NAND2_X1 U2521 ( .A1(n2100), .A2(n2099), .ZN(n4372) );
  OR2_X1 U2522 ( .A1(n3961), .A2(n4361), .ZN(n2099) );
  NAND2_X1 U2523 ( .A1(n3959), .A2(REG1_REG_8__SCAN_IN), .ZN(n2100) );
  NAND2_X1 U2524 ( .A1(n4387), .A2(n3965), .ZN(n4392) );
  NAND2_X1 U2525 ( .A1(n4419), .A2(n3970), .ZN(n3971) );
  XNOR2_X1 U2526 ( .A(n3951), .B(n3974), .ZN(n4446) );
  NAND2_X1 U2527 ( .A1(n4446), .A2(n4444), .ZN(n4445) );
  AND2_X1 U2528 ( .A1(n2607), .A2(n2606), .ZN(n3684) );
  OR2_X1 U2529 ( .A1(n3699), .A2(n2658), .ZN(n2607) );
  NAND2_X1 U2530 ( .A1(n2125), .A2(n2123), .ZN(n2708) );
  AOI21_X1 U2531 ( .B1(n2126), .B2(n2129), .A(n2124), .ZN(n2123) );
  INV_X1 U2532 ( .A(n3416), .ZN(n2124) );
  NOR2_X1 U2533 ( .A1(n2058), .A2(n2185), .ZN(n2184) );
  OR2_X1 U2534 ( .A1(n2056), .A2(n2182), .ZN(n2181) );
  AND2_X1 U2535 ( .A1(n2598), .A2(n2581), .ZN(n4033) );
  OR2_X1 U2536 ( .A1(n4055), .A2(n3447), .ZN(n4021) );
  AOI21_X1 U2537 ( .B1(n2048), .B2(n2159), .A(n2155), .ZN(n2154) );
  INV_X1 U2538 ( .A(n3463), .ZN(n2155) );
  NAND2_X1 U2539 ( .A1(n2513), .A2(REG3_REG_19__SCAN_IN), .ZN(n2521) );
  AND3_X1 U2540 ( .A1(n2508), .A2(n2507), .A3(n2506), .ZN(n4156) );
  INV_X1 U2541 ( .A(n4175), .ZN(n4181) );
  OR2_X1 U2542 ( .A1(n2489), .A2(n4686), .ZN(n2501) );
  AOI21_X1 U2543 ( .B1(n2194), .B2(n2046), .A(n2193), .ZN(n3400) );
  INV_X1 U2544 ( .A(n2195), .ZN(n2193) );
  AOI21_X1 U2545 ( .B1(n2046), .B2(n2196), .A(n2199), .ZN(n2195) );
  NAND2_X1 U2546 ( .A1(n2111), .A2(n2109), .ZN(n3428) );
  AND2_X1 U2547 ( .A1(n2110), .A2(n3528), .ZN(n2109) );
  NAND2_X1 U2548 ( .A1(n2055), .A2(n2115), .ZN(n2110) );
  OR2_X1 U2549 ( .A1(n2419), .A2(n4701), .ZN(n2430) );
  INV_X1 U2550 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2429) );
  NAND2_X1 U2551 ( .A1(n2112), .A2(n3490), .ZN(n3294) );
  NAND2_X1 U2552 ( .A1(n3167), .A2(n3486), .ZN(n2112) );
  OR2_X1 U2553 ( .A1(n3082), .A2(n2417), .ZN(n2173) );
  INV_X1 U2554 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2369) );
  INV_X1 U2555 ( .A(n2121), .ZN(n2120) );
  AOI21_X1 U2556 ( .B1(n2121), .B2(n2119), .A(n2118), .ZN(n2117) );
  AND2_X1 U2557 ( .A1(n2122), .A2(n3520), .ZN(n2121) );
  INV_X1 U2558 ( .A(n3280), .ZN(n3275) );
  NAND2_X1 U2559 ( .A1(n2398), .A2(REG3_REG_8__SCAN_IN), .ZN(n2382) );
  AND2_X1 U2560 ( .A1(n2627), .A2(n3518), .ZN(n3515) );
  AND4_X1 U2561 ( .A1(n2404), .A2(n2403), .A3(n2402), .A4(n2401), .ZN(n3190)
         );
  INV_X1 U2562 ( .A(n3913), .ZN(n3144) );
  AND2_X1 U2563 ( .A1(n2736), .A2(n2768), .ZN(n2827) );
  OR2_X1 U2564 ( .A1(n2763), .A2(D_REG_1__SCAN_IN), .ZN(n2826) );
  NAND2_X1 U2565 ( .A1(n2625), .A2(n3512), .ZN(n3058) );
  OR2_X1 U2566 ( .A1(n2995), .A2(n2624), .ZN(n2625) );
  NAND2_X1 U2567 ( .A1(n2982), .A2(n3501), .ZN(n2732) );
  NAND2_X1 U2568 ( .A1(n2732), .A2(n3471), .ZN(n2731) );
  INV_X1 U2569 ( .A(n4302), .ZN(n3069) );
  OR2_X1 U2570 ( .A1(n2977), .A2(n3496), .ZN(n2982) );
  NAND2_X1 U2571 ( .A1(n4043), .A2(n4032), .ZN(n4031) );
  AND2_X1 U2572 ( .A1(n4061), .A2(n4045), .ZN(n4043) );
  NOR2_X1 U2573 ( .A1(n4082), .A2(n4242), .ZN(n4061) );
  OR2_X1 U2574 ( .A1(n4097), .A2(n3644), .ZN(n4082) );
  NAND2_X1 U2575 ( .A1(n4113), .A2(n4095), .ZN(n4097) );
  AND2_X1 U2576 ( .A1(n4138), .A2(n4115), .ZN(n4113) );
  INV_X1 U2577 ( .A(n4260), .ZN(n4115) );
  NOR2_X1 U2578 ( .A1(n2045), .A2(n4540), .ZN(n4260) );
  NOR2_X2 U2579 ( .A1(n4161), .A2(n4131), .ZN(n4138) );
  NAND2_X1 U2580 ( .A1(n4182), .A2(n4181), .ZN(n4180) );
  NAND2_X1 U2581 ( .A1(n3327), .A2(n3591), .ZN(n3262) );
  INV_X1 U2582 ( .A(n3726), .ZN(n3591) );
  AND2_X1 U2583 ( .A1(n3325), .A2(n3588), .ZN(n3327) );
  NOR2_X2 U2584 ( .A1(n3302), .A2(n3782), .ZN(n3325) );
  INV_X1 U2585 ( .A(n3374), .ZN(n3372) );
  NAND2_X1 U2586 ( .A1(n2075), .A2(n2074), .ZN(n3226) );
  INV_X1 U2587 ( .A(n3086), .ZN(n2075) );
  INV_X1 U2588 ( .A(n3236), .ZN(n3252) );
  INV_X1 U2589 ( .A(n3147), .ZN(n3143) );
  NAND2_X1 U2590 ( .A1(n3084), .A2(n3143), .ZN(n3086) );
  AND4_X1 U2591 ( .A1(n2350), .A2(n2349), .A3(n2348), .A4(n2347), .ZN(n3125)
         );
  INV_X1 U2592 ( .A(n3133), .ZN(n3126) );
  NAND2_X1 U2593 ( .A1(n3017), .A2(n3016), .ZN(n3018) );
  INV_X1 U2594 ( .A(n3011), .ZN(n3016) );
  AND2_X1 U2595 ( .A1(n2909), .A2(n2623), .ZN(n4302) );
  INV_X1 U2596 ( .A(n4293), .ZN(n4283) );
  INV_X1 U2597 ( .A(n4220), .ZN(n4295) );
  INV_X1 U2598 ( .A(n4261), .ZN(n4299) );
  INV_X1 U2599 ( .A(n2283), .ZN(n2656) );
  AND2_X1 U2600 ( .A1(n2053), .A2(n2279), .ZN(n2710) );
  NAND2_X1 U2601 ( .A1(n2218), .A2(IR_REG_31__SCAN_IN), .ZN(n2680) );
  NAND2_X1 U2602 ( .A1(n2673), .A2(n2620), .ZN(n2218) );
  XNOR2_X1 U2603 ( .A(n2621), .B(n2620), .ZN(n2830) );
  INV_X1 U2604 ( .A(IR_REG_21__SCAN_IN), .ZN(n2611) );
  AND2_X1 U2605 ( .A1(n2485), .A2(n2484), .ZN(n3955) );
  INV_X1 U2606 ( .A(IR_REG_3__SCAN_IN), .ZN(n2330) );
  NOR2_X2 U2607 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2317)
         );
  INV_X1 U2608 ( .A(n2207), .ZN(n2206) );
  OAI21_X1 U2609 ( .B1(n2212), .B2(n2208), .A(n2211), .ZN(n2207) );
  NAND3_X1 U2610 ( .A1(n2222), .A2(n2221), .A3(n2050), .ZN(n3712) );
  NAND2_X1 U2611 ( .A1(n3659), .A2(n2062), .ZN(n2222) );
  OAI21_X1 U2612 ( .B1(n3742), .B2(n2242), .A(n2239), .ZN(n2233) );
  XOR2_X1 U2613 ( .A(n3612), .B(n3611), .Z(n3800) );
  AND4_X1 U2614 ( .A1(n2341), .A2(n2340), .A3(n2339), .A4(n2338), .ZN(n3132)
         );
  NAND2_X1 U2615 ( .A1(n2296), .A2(REG3_REG_1__SCAN_IN), .ZN(n2298) );
  OR2_X1 U2616 ( .A1(n2303), .A2(n2294), .ZN(n2300) );
  NAND2_X1 U2617 ( .A1(n2238), .A2(n2237), .ZN(n2236) );
  NAND2_X1 U2618 ( .A1(n2235), .A2(n2238), .ZN(n2234) );
  INV_X1 U2619 ( .A(n2242), .ZN(n2237) );
  AND2_X1 U2620 ( .A1(n2534), .A2(n2533), .ZN(n4133) );
  NAND2_X1 U2621 ( .A1(n2203), .A2(n3641), .ZN(n3852) );
  NAND2_X1 U2622 ( .A1(n3742), .A2(n3370), .ZN(n3577) );
  NAND2_X1 U2623 ( .A1(n2889), .A2(n2890), .ZN(n2891) );
  AOI21_X1 U2624 ( .B1(n3789), .B2(n3790), .A(n3791), .ZN(n3877) );
  INV_X1 U2625 ( .A(n4237), .ZN(n4046) );
  NAND2_X1 U2626 ( .A1(n2556), .A2(n2555), .ZN(n4243) );
  OR2_X1 U2627 ( .A1(n2728), .A2(n2841), .ZN(n3903) );
  INV_X1 U2628 ( .A(n4294), .ZN(n4195) );
  INV_X1 U2629 ( .A(n3745), .ZN(n3908) );
  NAND4_X1 U2630 ( .A1(n2376), .A2(n2375), .A3(n2374), .A4(n2373), .ZN(n3910)
         );
  NAND2_X1 U2631 ( .A1(n2248), .A2(n2386), .ZN(n3911) );
  AND3_X1 U2632 ( .A1(n2385), .A2(n2384), .A3(n2383), .ZN(n2248) );
  INV_X1 U2633 ( .A(n3190), .ZN(n3912) );
  AND3_X1 U2634 ( .A1(n2326), .A2(n2325), .A3(n2324), .ZN(n2328) );
  OR2_X1 U2635 ( .A1(n2303), .A2(n2322), .ZN(n2326) );
  INV_X1 U2636 ( .A(n2902), .ZN(n3917) );
  NAND2_X1 U2637 ( .A1(n2777), .A2(n2778), .ZN(n2933) );
  XNOR2_X1 U2638 ( .A(n2135), .B(n2797), .ZN(n2796) );
  INV_X1 U2639 ( .A(n2142), .ZN(n2804) );
  XNOR2_X1 U2640 ( .A(n2140), .B(n2139), .ZN(n2819) );
  OAI22_X1 U2641 ( .A1(n3941), .A2(n4478), .B1(n4361), .B2(n2090), .ZN(n4375)
         );
  INV_X1 U2642 ( .A(n2092), .ZN(n2090) );
  NAND2_X1 U2643 ( .A1(n4382), .A2(n3944), .ZN(n4395) );
  NAND2_X1 U2644 ( .A1(n4407), .A2(n3969), .ZN(n4420) );
  NAND2_X1 U2645 ( .A1(n4420), .A2(n4421), .ZN(n4419) );
  NAND2_X1 U2646 ( .A1(n4402), .A2(n3947), .ZN(n4415) );
  XNOR2_X1 U2647 ( .A(n3971), .B(n4432), .ZN(n4429) );
  XNOR2_X1 U2648 ( .A(n3948), .B(n4432), .ZN(n4425) );
  NOR2_X1 U2649 ( .A1(n4435), .A2(n4434), .ZN(n4433) );
  NOR2_X1 U2650 ( .A1(n4450), .A2(n3976), .ZN(n4459) );
  INV_X1 U2651 ( .A(n3684), .ZN(n4224) );
  NAND2_X1 U2652 ( .A1(n2128), .A2(n2126), .ZN(n4008) );
  NAND2_X1 U2653 ( .A1(n2128), .A2(n3544), .ZN(n4006) );
  NAND2_X1 U2654 ( .A1(n2186), .A2(n2577), .ZN(n4020) );
  NAND2_X1 U2655 ( .A1(n2568), .A2(n2187), .ZN(n2186) );
  AND2_X1 U2656 ( .A1(n2564), .A2(n2563), .ZN(n4050) );
  AND2_X1 U2657 ( .A1(n2527), .A2(n2526), .ZN(n4120) );
  NAND2_X1 U2658 ( .A1(n2157), .A2(n2158), .ZN(n4125) );
  OR2_X1 U2659 ( .A1(n4171), .A2(n2159), .ZN(n2157) );
  NAND2_X1 U2660 ( .A1(n4170), .A2(n2256), .ZN(n4148) );
  NAND2_X1 U2661 ( .A1(n4204), .A2(n3493), .ZN(n3398) );
  AND4_X1 U2662 ( .A1(n2293), .A2(n2292), .A3(n2291), .A4(n2290), .ZN(n4287)
         );
  NAND2_X1 U2663 ( .A1(n2198), .A2(n2247), .ZN(n4191) );
  AND2_X1 U2664 ( .A1(n2198), .A2(n2046), .ZN(n4190) );
  AND4_X1 U2665 ( .A1(n2470), .A2(n2469), .A3(n2468), .A4(n2467), .ZN(n3593)
         );
  AND2_X1 U2666 ( .A1(n2164), .A2(n2166), .ZN(n3201) );
  NAND2_X1 U2667 ( .A1(n2451), .A2(n2245), .ZN(n3324) );
  NAND2_X1 U2668 ( .A1(n2180), .A2(n2178), .ZN(n3304) );
  INV_X1 U2669 ( .A(n2179), .ZN(n2178) );
  NAND4_X1 U2670 ( .A1(n2425), .A2(n2424), .A3(n2423), .A4(n2422), .ZN(n3909)
         );
  OR2_X1 U2671 ( .A1(n2311), .A2(n2418), .ZN(n2424) );
  INV_X1 U2672 ( .A(n3910), .ZN(n3276) );
  OR2_X1 U2673 ( .A1(n2860), .A2(n2740), .ZN(n4476) );
  INV_X1 U2674 ( .A(n4210), .ZN(n4112) );
  AND2_X1 U2675 ( .A1(n3056), .A2(n2993), .ZN(n4520) );
  INV_X1 U2676 ( .A(n2959), .ZN(n2965) );
  NAND4_X1 U2677 ( .A1(n2307), .A2(n2306), .A3(n2305), .A4(n2304), .ZN(n2852)
         );
  OR2_X1 U2678 ( .A1(n2303), .A2(n2302), .ZN(n2306) );
  INV_X1 U2679 ( .A(n3701), .ZN(n4196) );
  INV_X1 U2680 ( .A(n2885), .ZN(n3916) );
  AND2_X1 U2681 ( .A1(n3697), .A2(n2665), .ZN(n2666) );
  AND3_X1 U2682 ( .A1(n3350), .A2(n3349), .A3(n3348), .ZN(n3353) );
  NAND2_X1 U2683 ( .A1(n2763), .A2(n2762), .ZN(n4496) );
  AND2_X1 U2684 ( .A1(n2280), .A2(n2281), .ZN(n2244) );
  INV_X1 U2685 ( .A(IR_REG_29__SCAN_IN), .ZN(n2281) );
  NAND2_X1 U2686 ( .A1(n2217), .A2(n2216), .ZN(n2674) );
  AOI21_X1 U2687 ( .B1(n2219), .B2(n2378), .A(n2378), .ZN(n2216) );
  INV_X1 U2688 ( .A(n3955), .ZN(n4502) );
  INV_X1 U2689 ( .A(n3967), .ZN(n4506) );
  OR2_X1 U2690 ( .A1(n2380), .A2(n2379), .ZN(n4510) );
  AND2_X1 U2691 ( .A1(n2408), .A2(n2407), .ZN(n4362) );
  CLKBUF_X1 U2692 ( .A(n2856), .Z(n2847) );
  INV_X1 U2693 ( .A(n2143), .ZN(n4474) );
  OAI21_X1 U2694 ( .B1(n4465), .B2(n2145), .A(n2144), .ZN(n2143) );
  XNOR2_X1 U2695 ( .A(n2096), .B(n2095), .ZN(n3986) );
  INV_X1 U2696 ( .A(n3953), .ZN(n2095) );
  OR2_X1 U2697 ( .A1(n4367), .A2(n4370), .ZN(n2078) );
  OAI211_X1 U2698 ( .C1(n2724), .C2(n4533), .A(n2723), .B(n2069), .ZN(U3547)
         );
  NAND2_X1 U2699 ( .A1(n2722), .A2(n3227), .ZN(n2723) );
  NAND2_X1 U2700 ( .A1(n2722), .A2(n3232), .ZN(n2726) );
  NAND2_X1 U2701 ( .A1(n2151), .A2(n2150), .ZN(U3351) );
  NAND2_X1 U2702 ( .A1(U3149), .A2(DATAI_1_), .ZN(n2150) );
  AND2_X1 U2703 ( .A1(n2197), .A2(n2247), .ZN(n2046) );
  NAND2_X1 U2704 ( .A1(n3835), .A2(n4162), .ZN(n2047) );
  NAND2_X1 U2705 ( .A1(n2135), .A2(n4365), .ZN(n2134) );
  INV_X1 U2706 ( .A(n3193), .ZN(n2074) );
  AND2_X1 U2707 ( .A1(n2158), .A2(n2064), .ZN(n2048) );
  INV_X1 U2708 ( .A(n4364), .ZN(n2948) );
  AND2_X1 U2709 ( .A1(n3246), .A2(n3245), .ZN(n2049) );
  NOR2_X1 U2710 ( .A1(n3780), .A2(n3588), .ZN(n2462) );
  INV_X1 U2711 ( .A(n2809), .ZN(n2105) );
  INV_X1 U2712 ( .A(n3578), .ZN(n3782) );
  NAND2_X1 U2713 ( .A1(n2227), .A2(n2226), .ZN(n2050) );
  NAND2_X1 U2714 ( .A1(n3497), .A2(n3501), .ZN(n2977) );
  INV_X2 U2715 ( .A(n4533), .ZN(n4535) );
  INV_X1 U2716 ( .A(n2296), .ZN(n2658) );
  OR2_X1 U2717 ( .A1(n3262), .A2(n2486), .ZN(n2051) );
  NAND2_X1 U2718 ( .A1(n2519), .A2(IR_REG_31__SCAN_IN), .ZN(n2614) );
  AND2_X1 U2719 ( .A1(n2108), .A2(n2846), .ZN(n2052) );
  NAND2_X1 U2720 ( .A1(n2215), .A2(n3615), .ZN(n3808) );
  NAND2_X1 U2721 ( .A1(n2510), .A2(n2132), .ZN(n2053) );
  NAND2_X1 U2722 ( .A1(n2328), .A2(n2327), .ZN(n2959) );
  AND4_X1 U2723 ( .A1(n2316), .A2(n2315), .A3(n2314), .A4(n2313), .ZN(n2885)
         );
  NAND2_X1 U2724 ( .A1(n2086), .A2(n2134), .ZN(n2054) );
  NAND2_X1 U2725 ( .A1(n2678), .A2(n2677), .ZN(n2841) );
  NAND2_X1 U2726 ( .A1(n3819), .A2(n2220), .ZN(n3789) );
  AND2_X1 U2727 ( .A1(n2632), .A2(n2113), .ZN(n2055) );
  AND2_X1 U2728 ( .A1(n4237), .A2(n4032), .ZN(n2056) );
  NAND2_X1 U2729 ( .A1(n3659), .A2(n3658), .ZN(n3819) );
  OAI21_X1 U2730 ( .B1(n2319), .B2(n2153), .A(n2152), .ZN(n3034) );
  NAND2_X1 U2731 ( .A1(n2317), .A2(n2107), .ZN(n2329) );
  INV_X1 U2732 ( .A(n2275), .ZN(n2669) );
  AND2_X1 U2733 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_29__SCAN_IN), .ZN(n2057)
         );
  NOR2_X1 U2734 ( .A1(n4237), .A2(n4032), .ZN(n2058) );
  INV_X1 U2735 ( .A(n2231), .ZN(n2351) );
  NAND2_X1 U2736 ( .A1(n2274), .A2(n2200), .ZN(n2059) );
  AND2_X1 U2737 ( .A1(n2134), .A2(n2948), .ZN(n2060) );
  NOR2_X1 U2738 ( .A1(n2351), .A2(n2258), .ZN(n2269) );
  OAI21_X1 U2739 ( .B1(n4174), .B2(n2161), .A(n2520), .ZN(n2160) );
  XNOR2_X1 U2740 ( .A(n2845), .B(n2043), .ZN(n2889) );
  INV_X1 U2741 ( .A(n2134), .ZN(n2133) );
  AND2_X1 U2742 ( .A1(n2849), .A2(n2848), .ZN(n2851) );
  AND2_X1 U2743 ( .A1(n2342), .A2(n2332), .ZN(n4365) );
  INV_X1 U2744 ( .A(n2177), .ZN(n2172) );
  NOR2_X1 U2745 ( .A1(n3455), .A2(n2179), .ZN(n2177) );
  NAND2_X1 U2746 ( .A1(n2275), .A2(n2274), .ZN(n2671) );
  NAND2_X1 U2747 ( .A1(n3910), .A2(n3275), .ZN(n2061) );
  INV_X1 U2748 ( .A(n3576), .ZN(n2241) );
  INV_X1 U2749 ( .A(n4363), .ZN(n2139) );
  NAND2_X1 U2750 ( .A1(n2156), .A2(n2154), .ZN(n4110) );
  OAI21_X1 U2751 ( .B1(n3742), .B2(n2236), .A(n2234), .ZN(n3840) );
  INV_X1 U2752 ( .A(n3518), .ZN(n2119) );
  INV_X1 U2753 ( .A(n2233), .ZN(n3775) );
  INV_X1 U2754 ( .A(n3472), .ZN(n2163) );
  INV_X1 U2755 ( .A(n3790), .ZN(n2229) );
  AND2_X1 U2756 ( .A1(n2228), .A2(n3658), .ZN(n2062) );
  OR2_X1 U2757 ( .A1(n2902), .A2(n3034), .ZN(n3497) );
  NOR2_X1 U2758 ( .A1(n4180), .A2(n3758), .ZN(n2079) );
  NAND2_X1 U2759 ( .A1(n3370), .A2(n2241), .ZN(n2243) );
  AND2_X1 U2760 ( .A1(n3745), .A2(n3372), .ZN(n2063) );
  INV_X1 U2761 ( .A(n3791), .ZN(n2230) );
  NAND2_X1 U2762 ( .A1(n4262), .A2(n4131), .ZN(n2064) );
  INV_X1 U2763 ( .A(n3874), .ZN(n2227) );
  AND4_X1 U2764 ( .A1(n2447), .A2(n2446), .A3(n2445), .A4(n2444), .ZN(n3580)
         );
  OAI21_X1 U2765 ( .B1(n3994), .B2(n4220), .A(n2716), .ZN(n2717) );
  OR2_X1 U2766 ( .A1(n4265), .A2(n4095), .ZN(n2065) );
  NAND2_X1 U2767 ( .A1(n3780), .A2(n3588), .ZN(n2066) );
  NAND2_X1 U2768 ( .A1(n2171), .A2(n2170), .ZN(n3287) );
  XNOR2_X1 U2769 ( .A(n2674), .B(IR_REG_24__SCAN_IN), .ZN(n2678) );
  INV_X1 U2770 ( .A(n3486), .ZN(n2114) );
  AND2_X1 U2771 ( .A1(n3502), .A2(n3505), .ZN(n3471) );
  INV_X1 U2772 ( .A(n3471), .ZN(n2320) );
  AND2_X1 U2773 ( .A1(n2180), .A2(n2177), .ZN(n2067) );
  INV_X1 U2774 ( .A(n2462), .ZN(n2166) );
  AND2_X1 U2775 ( .A1(n2844), .A2(n2843), .ZN(n2068) );
  OR2_X1 U2776 ( .A1(n4535), .A2(n2718), .ZN(n2069) );
  INV_X1 U2777 ( .A(n4361), .ZN(n2091) );
  OR2_X1 U2778 ( .A1(n4498), .A2(n3978), .ZN(n2070) );
  AND2_X1 U2779 ( .A1(n2085), .A2(n2083), .ZN(n2071) );
  NOR2_X2 U2780 ( .A1(n3226), .A2(n3252), .ZN(n3225) );
  NOR2_X2 U2781 ( .A1(n3062), .A2(n3126), .ZN(n3084) );
  NOR2_X2 U2782 ( .A1(n2077), .A2(n2059), .ZN(n2132) );
  NAND4_X1 U2783 ( .A1(n2270), .A2(n2273), .A3(n2272), .A4(n2271), .ZN(n2077)
         );
  INV_X1 U2784 ( .A(n2077), .ZN(n2076) );
  NAND2_X1 U2785 ( .A1(n4369), .A2(n2078), .ZN(U3261) );
  INV_X1 U2786 ( .A(n2079), .ZN(n4161) );
  NOR2_X4 U2787 ( .A1(n4194), .A2(n4282), .ZN(n4182) );
  AND2_X2 U2788 ( .A1(n2131), .A2(n2510), .ZN(n2654) );
  NAND3_X1 U2789 ( .A1(n2071), .A2(REG2_REG_4__SCAN_IN), .A3(n2082), .ZN(n2080) );
  NAND2_X1 U2790 ( .A1(n2071), .A2(n2082), .ZN(n2942) );
  NAND2_X1 U2791 ( .A1(n2060), .A2(n2086), .ZN(n2082) );
  NAND2_X1 U2792 ( .A1(n2796), .A2(REG2_REG_3__SCAN_IN), .ZN(n2086) );
  NAND2_X1 U2793 ( .A1(n2796), .A2(n2084), .ZN(n2083) );
  NOR2_X1 U2794 ( .A1(n2948), .A2(n2323), .ZN(n2084) );
  NAND2_X1 U2795 ( .A1(n2088), .A2(n2087), .ZN(n3933) );
  NAND2_X1 U2796 ( .A1(n2149), .A2(n2775), .ZN(n2087) );
  AND3_X2 U2797 ( .A1(n2317), .A2(n2107), .A3(n2106), .ZN(n2231) );
  AND4_X2 U2798 ( .A1(n2300), .A2(n2299), .A3(n2297), .A4(n2298), .ZN(n2902)
         );
  NAND2_X1 U2799 ( .A1(n3167), .A2(n2055), .ZN(n2111) );
  NAND2_X1 U2800 ( .A1(n4204), .A2(n2116), .ZN(n4150) );
  OAI21_X1 U2801 ( .B1(n3065), .B2(n2120), .A(n2117), .ZN(n3154) );
  OAI21_X1 U2802 ( .B1(n3065), .B2(n2628), .A(n3518), .ZN(n3220) );
  NAND2_X1 U2803 ( .A1(n3518), .A2(n2628), .ZN(n2122) );
  NAND2_X1 U2804 ( .A1(n4055), .A2(n2126), .ZN(n2125) );
  OR2_X1 U2805 ( .A1(n4055), .A2(n2129), .ZN(n2128) );
  NOR2_X1 U2806 ( .A1(n2192), .A2(n2191), .ZN(n2190) );
  NAND2_X1 U2807 ( .A1(n2149), .A2(REG2_REG_1__SCAN_IN), .ZN(n2930) );
  NAND2_X1 U2808 ( .A1(n2149), .A2(REG1_REG_1__SCAN_IN), .ZN(n2786) );
  NAND2_X1 U2809 ( .A1(n2149), .A2(STATE_REG_SCAN_IN), .ZN(n2151) );
  XNOR2_X1 U2810 ( .A(n2149), .B(n2295), .ZN(n3930) );
  NAND2_X1 U2811 ( .A1(n2045), .A2(n2149), .ZN(n2152) );
  NAND2_X1 U2812 ( .A1(n3927), .A2(n2149), .ZN(n3937) );
  NAND2_X1 U2813 ( .A1(n4171), .A2(n2048), .ZN(n2156) );
  INV_X1 U2814 ( .A(n2256), .ZN(n2161) );
  NAND2_X1 U2815 ( .A1(n4171), .A2(n4174), .ZN(n4170) );
  NAND2_X1 U2816 ( .A1(n2451), .A2(n2165), .ZN(n2164) );
  INV_X1 U2817 ( .A(n3082), .ZN(n2169) );
  NAND3_X1 U2818 ( .A1(n2168), .A2(n2177), .A3(n2169), .ZN(n2167) );
  NAND2_X1 U2819 ( .A1(n2416), .A2(n2173), .ZN(n3168) );
  NOR2_X1 U2820 ( .A1(n3308), .A2(n3365), .ZN(n2179) );
  INV_X1 U2821 ( .A(n2568), .ZN(n2183) );
  OAI22_X1 U2822 ( .A1(n2183), .A2(n2181), .B1(n2056), .B2(n2184), .ZN(n4004)
         );
  NAND2_X1 U2823 ( .A1(n2568), .A2(n2567), .ZN(n4041) );
  NOR2_X1 U2824 ( .A1(n2578), .A2(n2188), .ZN(n2187) );
  INV_X1 U2825 ( .A(n2567), .ZN(n2188) );
  NOR2_X1 U2826 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_29__SCAN_IN), .ZN(n2191)
         );
  INV_X1 U2827 ( .A(n3261), .ZN(n2194) );
  AND2_X1 U2828 ( .A1(n3904), .A2(n4296), .ZN(n2199) );
  AND3_X2 U2829 ( .A1(n2231), .A2(n2268), .A3(n2232), .ZN(n2510) );
  NAND2_X1 U2830 ( .A1(n2203), .A2(n2201), .ZN(n3734) );
  NAND2_X1 U2831 ( .A1(n3828), .A2(n3831), .ZN(n3767) );
  NOR2_X1 U2832 ( .A1(n3642), .A2(n2205), .ZN(n2204) );
  INV_X1 U2833 ( .A(n3831), .ZN(n2205) );
  NOR2_X1 U2834 ( .A1(n3141), .A2(n2254), .ZN(n3189) );
  NAND2_X1 U2835 ( .A1(n2209), .A2(n2206), .ZN(n3248) );
  NAND2_X1 U2836 ( .A1(n3141), .A2(n2210), .ZN(n2209) );
  NAND2_X1 U2837 ( .A1(n2215), .A2(n2214), .ZN(n3754) );
  NAND2_X1 U2838 ( .A1(n2673), .A2(n2219), .ZN(n2217) );
  NAND2_X1 U2839 ( .A1(n3820), .A2(n3822), .ZN(n2220) );
  NAND2_X1 U2840 ( .A1(n3820), .A2(n2223), .ZN(n2221) );
  INV_X1 U2841 ( .A(n2228), .ZN(n2225) );
  NAND4_X1 U2842 ( .A1(n2231), .A2(n2509), .A3(n2232), .A4(n2268), .ZN(n2518)
         );
  OR2_X1 U2843 ( .A1(n2310), .A2(n2874), .ZN(n2304) );
  NAND2_X1 U2844 ( .A1(n4358), .A2(n2756), .ZN(n2310) );
  NAND2_X1 U2845 ( .A1(n2869), .A2(n2871), .ZN(n2870) );
  INV_X1 U2846 ( .A(n4367), .ZN(n4187) );
  OR2_X1 U2847 ( .A1(n3907), .A2(n3782), .ZN(n2245) );
  AND2_X1 U2848 ( .A1(n4195), .A2(n4282), .ZN(n2246) );
  AND4_X1 U2849 ( .A1(n2481), .A2(n2480), .A3(n2479), .A4(n2478), .ZN(n4300)
         );
  INV_X1 U2850 ( .A(n4300), .ZN(n2487) );
  OR2_X1 U2851 ( .A1(n2487), .A2(n2486), .ZN(n2247) );
  NAND2_X1 U2852 ( .A1(n4535), .A2(n4302), .ZN(n4292) );
  NAND2_X1 U2853 ( .A1(n4529), .A2(n4302), .ZN(n4355) );
  INV_X1 U2854 ( .A(n2623), .ZN(n2651) );
  OR2_X1 U2855 ( .A1(n3706), .A2(n4292), .ZN(n2249) );
  OR2_X1 U2856 ( .A1(n3706), .A2(n4355), .ZN(n2250) );
  NAND2_X1 U2857 ( .A1(n4195), .A2(n3616), .ZN(n2251) );
  AND2_X1 U2858 ( .A1(n3987), .A2(n3900), .ZN(n2252) );
  NOR2_X1 U2859 ( .A1(n3862), .A2(n3626), .ZN(n2253) );
  AND2_X1 U2860 ( .A1(n3140), .A2(n3139), .ZN(n2254) );
  AND2_X1 U2861 ( .A1(n2959), .A2(n3011), .ZN(n2255) );
  OR2_X1 U2862 ( .A1(n4284), .A2(n4175), .ZN(n2256) );
  OR2_X1 U2863 ( .A1(n3905), .A2(n3726), .ZN(n2257) );
  INV_X1 U2864 ( .A(n3780), .ZN(n3906) );
  AND4_X1 U2865 ( .A1(n2458), .A2(n2457), .A3(n2456), .A4(n2455), .ZN(n3780)
         );
  NAND2_X1 U2866 ( .A1(n3910), .A2(n3280), .ZN(n2391) );
  OR2_X1 U2867 ( .A1(n2830), .A2(n4360), .ZN(n2844) );
  AND2_X1 U2868 ( .A1(n2649), .A2(n4022), .ZN(n2650) );
  INV_X1 U2869 ( .A(n3596), .ZN(n2486) );
  NOR2_X1 U2870 ( .A1(n2464), .A2(n4660), .ZN(n2463) );
  NAND2_X1 U2871 ( .A1(n3614), .A2(n3613), .ZN(n3615) );
  INV_X1 U2872 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2452) );
  INV_X1 U2873 ( .A(n2570), .ZN(n2569) );
  NOR2_X1 U2874 ( .A1(n2764), .A2(n2751), .ZN(n2677) );
  INV_X1 U2875 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2396) );
  INV_X1 U2876 ( .A(IR_REG_25__SCAN_IN), .ZN(n2274) );
  AND4_X1 U2877 ( .A1(n2267), .A2(n2266), .A3(n2265), .A4(n2264), .ZN(n2268)
         );
  OR2_X1 U2878 ( .A1(n3599), .A2(n3598), .ZN(n3721) );
  INV_X1 U2879 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4701) );
  NAND2_X1 U2880 ( .A1(n2285), .A2(REG3_REG_16__SCAN_IN), .ZN(n2489) );
  INV_X1 U2881 ( .A(n2052), .ZN(n2890) );
  NAND2_X1 U2882 ( .A1(n2569), .A2(REG3_REG_25__SCAN_IN), .ZN(n2580) );
  NAND2_X1 U2883 ( .A1(n2359), .A2(REG3_REG_6__SCAN_IN), .ZN(n2397) );
  OR2_X1 U2884 ( .A1(n2382), .A2(n2369), .ZN(n2419) );
  NOR2_X1 U2885 ( .A1(n2397), .A2(n2396), .ZN(n2398) );
  INV_X1 U2886 ( .A(n3616), .ZN(n4282) );
  AND2_X1 U2887 ( .A1(n3508), .A2(n3512), .ZN(n2994) );
  AND3_X1 U2888 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2359) );
  NAND2_X1 U2889 ( .A1(n3829), .A2(n3830), .ZN(n3828) );
  OR2_X1 U2890 ( .A1(n2865), .A2(n2863), .ZN(n3856) );
  OR2_X1 U2891 ( .A1(n2865), .A2(n2864), .ZN(n3857) );
  NAND2_X1 U2892 ( .A1(n3604), .A2(n3603), .ZN(n3887) );
  INV_X1 U2893 ( .A(n4365), .ZN(n2797) );
  INV_X1 U2894 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4660) );
  AOI21_X1 U2895 ( .B1(n2705), .B2(n3482), .A(n2704), .ZN(n2706) );
  INV_X1 U2896 ( .A(n3454), .ZN(n2637) );
  AND2_X1 U2897 ( .A1(n3507), .A2(n3504), .ZN(n3452) );
  OR2_X1 U2898 ( .A1(n2763), .A2(D_REG_0__SCAN_IN), .ZN(n2696) );
  NOR2_X1 U2899 ( .A1(n2319), .A2(n4658), .ZN(n4233) );
  INV_X1 U2900 ( .A(n2546), .ZN(n4095) );
  OR2_X1 U2901 ( .A1(n2763), .A2(n2692), .ZN(n2736) );
  INV_X1 U2902 ( .A(n3856), .ZN(n3891) );
  NOR2_X1 U2903 ( .A1(n3044), .A2(n3045), .ZN(n3121) );
  OR2_X1 U2904 ( .A1(n2521), .A2(n4669), .ZN(n2528) );
  INV_X1 U2905 ( .A(n3857), .ZN(n3889) );
  AND2_X1 U2906 ( .A1(n2544), .A2(n2543), .ZN(n4265) );
  AND2_X1 U2907 ( .A1(n2780), .A2(n2779), .ZN(n3923) );
  AND2_X1 U2908 ( .A1(n3923), .A2(n3559), .ZN(n4413) );
  OR2_X1 U2909 ( .A1(n3077), .A2(n3515), .ZN(n4523) );
  AND2_X1 U2910 ( .A1(n2358), .A2(n2357), .ZN(n3082) );
  INV_X1 U2911 ( .A(n4164), .ZN(n4490) );
  AND2_X1 U2912 ( .A1(n4106), .A2(n4261), .ZN(n4012) );
  NAND2_X1 U2913 ( .A1(n2696), .A2(n2695), .ZN(n2738) );
  INV_X1 U2914 ( .A(n3758), .ZN(n4162) );
  NAND2_X1 U2915 ( .A1(n4137), .A2(n3309), .ZN(n4521) );
  AND2_X1 U2916 ( .A1(n2912), .A2(n2830), .ZN(n4519) );
  INV_X1 U2917 ( .A(n2284), .ZN(n2756) );
  INV_X1 U2918 ( .A(n2830), .ZN(n3562) );
  AND2_X1 U2919 ( .A1(n2440), .A2(n2448), .ZN(n3957) );
  AND2_X1 U2920 ( .A1(n2780), .A2(n2773), .ZN(n4468) );
  AND2_X1 U2921 ( .A1(n2970), .A2(n2969), .ZN(n3895) );
  OR2_X1 U2922 ( .A1(n2865), .A2(n2859), .ZN(n3884) );
  INV_X1 U2923 ( .A(n3674), .ZN(n4028) );
  INV_X1 U2924 ( .A(n4120), .ZN(n4262) );
  INV_X1 U2925 ( .A(n3580), .ZN(n3907) );
  INV_X1 U2926 ( .A(n3132), .ZN(n3915) );
  INV_X1 U2927 ( .A(n4413), .ZN(n4464) );
  OR2_X1 U2928 ( .A1(n4183), .A2(n3069), .ZN(n4164) );
  OR2_X1 U2929 ( .A1(n2700), .A2(n2738), .ZN(n4533) );
  AND3_X1 U2930 ( .A1(n4526), .A2(n4525), .A3(n4524), .ZN(n4534) );
  OR2_X1 U2931 ( .A1(n2700), .A2(n2828), .ZN(n4527) );
  INV_X1 U2932 ( .A(n2678), .ZN(n2765) );
  AND2_X1 U2933 ( .A1(n2771), .A2(STATE_REG_SCAN_IN), .ZN(n4497) );
  INV_X1 U2934 ( .A(n3956), .ZN(n4505) );
  AND2_X1 U2935 ( .A1(n2368), .A2(n2387), .ZN(n4363) );
  NAND2_X1 U2936 ( .A1(n2269), .A2(n2259), .ZN(n2436) );
  NOR2_X2 U2937 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2267)
         );
  INV_X1 U2938 ( .A(n2267), .ZN(n2260) );
  NOR2_X1 U2939 ( .A1(n2459), .A2(IR_REG_13__SCAN_IN), .ZN(n2471) );
  INV_X1 U2940 ( .A(IR_REG_14__SCAN_IN), .ZN(n2261) );
  NAND2_X1 U2941 ( .A1(n2471), .A2(n2261), .ZN(n2262) );
  NAND2_X1 U2942 ( .A1(n2262), .A2(IR_REG_31__SCAN_IN), .ZN(n2483) );
  INV_X1 U2943 ( .A(IR_REG_15__SCAN_IN), .ZN(n2482) );
  NAND2_X1 U2944 ( .A1(n2483), .A2(n2482), .ZN(n2485) );
  NAND2_X1 U2945 ( .A1(n2485), .A2(IR_REG_31__SCAN_IN), .ZN(n2263) );
  XNOR2_X1 U2946 ( .A(n2263), .B(IR_REG_16__SCAN_IN), .ZN(n3974) );
  INV_X1 U2947 ( .A(n2654), .ZN(n2278) );
  NAND2_X1 U2948 ( .A1(n2276), .A2(n2378), .ZN(n2277) );
  NAND2_X1 U2949 ( .A1(n2278), .A2(n2277), .ZN(n2711) );
  AND2_X1 U2950 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2279)
         );
  MUX2_X2 U2951 ( .A(n2711), .B(n2710), .S(IR_REG_28__SCAN_IN), .Z(n2319) );
  MUX2_X1 U2952 ( .A(DATAI_16_), .B(n3974), .S(n2512), .Z(n4296) );
  INV_X1 U2953 ( .A(n4358), .ZN(n2288) );
  NAND2_X1 U2954 ( .A1(n2288), .A2(n2284), .ZN(n2303) );
  INV_X1 U2955 ( .A(n2303), .ZN(n3410) );
  NAND2_X1 U2956 ( .A1(n3410), .A2(REG0_REG_16__SCAN_IN), .ZN(n2293) );
  OR2_X1 U2957 ( .A1(n2312), .A2(n4444), .ZN(n2292) );
  INV_X1 U2958 ( .A(n2285), .ZN(n2477) );
  INV_X1 U2959 ( .A(REG3_REG_16__SCAN_IN), .ZN(n2286) );
  NAND2_X1 U2960 ( .A1(n2477), .A2(n2286), .ZN(n2287) );
  NAND2_X1 U2961 ( .A1(n2489), .A2(n2287), .ZN(n4198) );
  OR2_X1 U2962 ( .A1(n2658), .A2(n4198), .ZN(n2291) );
  INV_X1 U2963 ( .A(n2311), .ZN(n2301) );
  INV_X1 U2964 ( .A(REG1_REG_16__SCAN_IN), .ZN(n2289) );
  OR2_X1 U2965 ( .A1(n2311), .A2(n2289), .ZN(n2290) );
  INV_X1 U2966 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2294) );
  INV_X1 U2967 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2295) );
  INV_X1 U2968 ( .A(n2310), .ZN(n2296) );
  NAND2_X1 U2969 ( .A1(n3409), .A2(REG2_REG_1__SCAN_IN), .ZN(n2297) );
  INV_X1 U2970 ( .A(n3034), .ZN(n2842) );
  INV_X1 U2971 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2302) );
  INV_X1 U2972 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2916) );
  OR2_X1 U2973 ( .A1(n2312), .A2(n2916), .ZN(n2305) );
  INV_X1 U2974 ( .A(REG3_REG_0__SCAN_IN), .ZN(n2874) );
  MUX2_X1 U2975 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(n2044), .Z(n2987) );
  AND2_X1 U2976 ( .A1(n2852), .A2(n2987), .ZN(n2979) );
  NAND2_X1 U2977 ( .A1(n3917), .A2(n3034), .ZN(n2308) );
  NAND2_X1 U2978 ( .A1(n2978), .A2(n2308), .ZN(n2729) );
  INV_X1 U2979 ( .A(n2729), .ZN(n2321) );
  INV_X1 U2980 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2309) );
  INV_X1 U2981 ( .A(REG3_REG_2__SCAN_IN), .ZN(n2923) );
  OR2_X1 U2982 ( .A1(n2310), .A2(n2923), .ZN(n2315) );
  INV_X1 U2983 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2906) );
  OR2_X1 U2984 ( .A1(n2311), .A2(n2906), .ZN(n2314) );
  INV_X1 U2985 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2774) );
  OR2_X1 U2986 ( .A1(n2312), .A2(n2774), .ZN(n2313) );
  OR2_X1 U2987 ( .A1(n2317), .A2(n2378), .ZN(n2318) );
  MUX2_X1 U2988 ( .A(DATAI_2_), .B(n4366), .S(n2045), .Z(n2900) );
  NAND2_X1 U2989 ( .A1(n2885), .A2(n2900), .ZN(n3502) );
  INV_X1 U2990 ( .A(n2900), .ZN(n2888) );
  NAND2_X1 U2991 ( .A1(n3916), .A2(n2888), .ZN(n3505) );
  NAND2_X1 U2992 ( .A1(n2885), .A2(n2888), .ZN(n3006) );
  INV_X1 U2993 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2322) );
  OR2_X1 U2994 ( .A1(n2658), .A2(REG3_REG_3__SCAN_IN), .ZN(n2325) );
  INV_X1 U2995 ( .A(REG2_REG_3__SCAN_IN), .ZN(n2323) );
  OR2_X1 U2996 ( .A1(n2312), .A2(n2323), .ZN(n2324) );
  INV_X1 U2997 ( .A(REG1_REG_3__SCAN_IN), .ZN(n3020) );
  OR2_X1 U2998 ( .A1(n2311), .A2(n3020), .ZN(n2327) );
  NAND2_X1 U2999 ( .A1(n2329), .A2(IR_REG_31__SCAN_IN), .ZN(n2331) );
  NAND2_X1 U3000 ( .A1(n2331), .A2(n2330), .ZN(n2342) );
  OR2_X1 U3001 ( .A1(n2331), .A2(n2330), .ZN(n2332) );
  NAND2_X1 U3002 ( .A1(n2965), .A2(n3016), .ZN(n2334) );
  AND2_X1 U3003 ( .A1(n3006), .A2(n2334), .ZN(n2335) );
  NAND2_X1 U3004 ( .A1(n3409), .A2(REG2_REG_4__SCAN_IN), .ZN(n2341) );
  INV_X1 U3005 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2336) );
  OR2_X1 U3006 ( .A1(n2303), .A2(n2336), .ZN(n2340) );
  XNOR2_X1 U3007 ( .A(REG3_REG_4__SCAN_IN), .B(REG3_REG_3__SCAN_IN), .ZN(n3051) );
  OR2_X1 U3008 ( .A1(n2658), .A2(n3051), .ZN(n2339) );
  INV_X1 U3009 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2337) );
  OR2_X1 U3010 ( .A1(n2311), .A2(n2337), .ZN(n2338) );
  NAND2_X1 U3011 ( .A1(n2342), .A2(IR_REG_31__SCAN_IN), .ZN(n2343) );
  XNOR2_X1 U3012 ( .A(n2343), .B(IR_REG_4__SCAN_IN), .ZN(n4364) );
  MUX2_X1 U3013 ( .A(DATAI_4_), .B(n4364), .S(n2512), .Z(n3048) );
  NAND2_X1 U3014 ( .A1(n3132), .A2(n3048), .ZN(n3508) );
  INV_X1 U3015 ( .A(n3048), .ZN(n3039) );
  NAND2_X1 U3016 ( .A1(n3915), .A2(n3039), .ZN(n3512) );
  NAND2_X1 U3017 ( .A1(n3915), .A2(n3048), .ZN(n3055) );
  AOI21_X1 U3018 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        REG3_REG_5__SCAN_IN), .ZN(n2344) );
  NOR2_X1 U3019 ( .A1(n2344), .A2(n2359), .ZN(n3112) );
  NAND2_X1 U3020 ( .A1(n2296), .A2(n3112), .ZN(n2350) );
  INV_X1 U3021 ( .A(REG0_REG_5__SCAN_IN), .ZN(n2345) );
  OR2_X1 U3022 ( .A1(n2303), .A2(n2345), .ZN(n2349) );
  INV_X1 U3023 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2808) );
  OR2_X1 U3024 ( .A1(n2311), .A2(n2808), .ZN(n2348) );
  INV_X1 U3025 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2346) );
  OR2_X1 U3026 ( .A1(n2312), .A2(n2346), .ZN(n2347) );
  INV_X1 U3027 ( .A(n3125), .ZN(n3914) );
  INV_X1 U3028 ( .A(DATAI_5_), .ZN(n4569) );
  NAND2_X1 U3029 ( .A1(n2351), .A2(IR_REG_31__SCAN_IN), .ZN(n2352) );
  MUX2_X1 U3030 ( .A(n2352), .B(IR_REG_31__SCAN_IN), .S(n2353), .Z(n2354) );
  NAND2_X1 U3031 ( .A1(n2231), .A2(n2353), .ZN(n2365) );
  NAND2_X1 U3032 ( .A1(n2354), .A2(n2365), .ZN(n2809) );
  MUX2_X1 U3033 ( .A(n4569), .B(n2809), .S(n2512), .Z(n3133) );
  NAND2_X1 U3034 ( .A1(n3914), .A2(n3126), .ZN(n2355) );
  AND2_X1 U3035 ( .A1(n3055), .A2(n2355), .ZN(n2356) );
  NAND2_X1 U3036 ( .A1(n3056), .A2(n2356), .ZN(n2358) );
  NAND2_X1 U3037 ( .A1(n3125), .A2(n3133), .ZN(n2357) );
  NAND2_X1 U3038 ( .A1(n3410), .A2(REG0_REG_6__SCAN_IN), .ZN(n2363) );
  INV_X1 U3039 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3087) );
  OR2_X1 U3040 ( .A1(n2312), .A2(n3087), .ZN(n2362) );
  OAI21_X1 U3041 ( .B1(n2359), .B2(REG3_REG_6__SCAN_IN), .A(n2397), .ZN(n3150)
         );
  OR2_X1 U3042 ( .A1(n2658), .A2(n3150), .ZN(n2361) );
  OR2_X1 U3043 ( .A1(n2311), .A2(n3103), .ZN(n2360) );
  NAND4_X1 U3044 ( .A1(n2363), .A2(n2362), .A3(n2361), .A4(n2360), .ZN(n3913)
         );
  NAND2_X1 U3045 ( .A1(n2365), .A2(IR_REG_31__SCAN_IN), .ZN(n2364) );
  MUX2_X1 U3046 ( .A(n2364), .B(IR_REG_31__SCAN_IN), .S(n2366), .Z(n2368) );
  INV_X1 U3047 ( .A(n2365), .ZN(n2367) );
  NAND2_X1 U3048 ( .A1(n2367), .A2(n2366), .ZN(n2387) );
  MUX2_X1 U3049 ( .A(DATAI_6_), .B(n4363), .S(n2512), .Z(n3147) );
  AND2_X1 U3050 ( .A1(n3913), .A2(n3147), .ZN(n3074) );
  NAND2_X1 U3051 ( .A1(n3410), .A2(REG0_REG_9__SCAN_IN), .ZN(n2376) );
  NAND2_X1 U3052 ( .A1(n2382), .A2(n2369), .ZN(n2370) );
  NAND2_X1 U3053 ( .A1(n2419), .A2(n2370), .ZN(n3283) );
  OR2_X1 U3054 ( .A1(n2658), .A2(n3283), .ZN(n2375) );
  INV_X1 U3055 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2371) );
  OR2_X1 U3056 ( .A1(n2311), .A2(n2371), .ZN(n2374) );
  INV_X1 U3057 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2372) );
  OR2_X1 U3058 ( .A1(n2312), .A2(n2372), .ZN(n2373) );
  NOR2_X1 U3059 ( .A1(n2269), .A2(n2378), .ZN(n2377) );
  MUX2_X1 U3060 ( .A(n2378), .B(n2377), .S(IR_REG_9__SCAN_IN), .Z(n2380) );
  INV_X1 U3061 ( .A(n2436), .ZN(n2379) );
  MUX2_X1 U3062 ( .A(DATAI_9_), .B(n3958), .S(n2512), .Z(n3280) );
  NAND2_X1 U3063 ( .A1(n3410), .A2(REG0_REG_8__SCAN_IN), .ZN(n2385) );
  INV_X1 U3064 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4478) );
  OR2_X1 U3065 ( .A1(n2312), .A2(n4478), .ZN(n2384) );
  OR2_X1 U3066 ( .A1(n2398), .A2(REG3_REG_8__SCAN_IN), .ZN(n2381) );
  NAND2_X1 U3067 ( .A1(n2382), .A2(n2381), .ZN(n4477) );
  OR2_X1 U3068 ( .A1(n2658), .A2(n4477), .ZN(n2383) );
  OR2_X1 U3069 ( .A1(n2311), .A2(n3230), .ZN(n2386) );
  INV_X1 U3070 ( .A(DATAI_8_), .ZN(n2390) );
  NAND2_X1 U3071 ( .A1(n2387), .A2(IR_REG_31__SCAN_IN), .ZN(n2406) );
  NAND2_X1 U3072 ( .A1(n2406), .A2(n2405), .ZN(n2408) );
  NAND2_X1 U3073 ( .A1(n2408), .A2(IR_REG_31__SCAN_IN), .ZN(n2389) );
  XNOR2_X1 U3074 ( .A(n2389), .B(n2388), .ZN(n4361) );
  MUX2_X1 U3075 ( .A(n2390), .B(n4361), .S(n2512), .Z(n3236) );
  NAND2_X1 U3076 ( .A1(n3911), .A2(n3252), .ZN(n3162) );
  NAND2_X1 U3077 ( .A1(n3238), .A2(n3236), .ZN(n3161) );
  INV_X1 U3078 ( .A(n3161), .ZN(n2392) );
  NAND2_X1 U3079 ( .A1(n2409), .A2(n2392), .ZN(n2394) );
  NAND2_X1 U3080 ( .A1(n3276), .A2(n3275), .ZN(n2393) );
  NAND2_X1 U3081 ( .A1(n2394), .A2(n2393), .ZN(n2411) );
  NAND2_X1 U3082 ( .A1(n3410), .A2(REG0_REG_7__SCAN_IN), .ZN(n2404) );
  INV_X1 U3083 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2395) );
  OR2_X1 U3084 ( .A1(n2312), .A2(n2395), .ZN(n2403) );
  AND2_X1 U3085 ( .A1(n2397), .A2(n2396), .ZN(n2399) );
  OR2_X1 U3086 ( .A1(n2399), .A2(n2398), .ZN(n3196) );
  OR2_X1 U3087 ( .A1(n2658), .A2(n3196), .ZN(n2402) );
  INV_X1 U3088 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2400) );
  OR2_X1 U3089 ( .A1(n2311), .A2(n2400), .ZN(n2401) );
  OR2_X1 U3090 ( .A1(n2406), .A2(n2405), .ZN(n2407) );
  MUX2_X1 U3091 ( .A(DATAI_7_), .B(n4362), .S(n2512), .Z(n3193) );
  NAND2_X1 U3092 ( .A1(n3912), .A2(n3193), .ZN(n3160) );
  AND2_X1 U3093 ( .A1(n3160), .A2(n2409), .ZN(n2410) );
  NOR2_X1 U3094 ( .A1(n2411), .A2(n2410), .ZN(n2415) );
  OR2_X1 U3095 ( .A1(n3074), .A2(n2415), .ZN(n2417) );
  NAND2_X1 U3096 ( .A1(n3190), .A2(n3193), .ZN(n2627) );
  NAND2_X1 U3097 ( .A1(n3912), .A2(n2074), .ZN(n3518) );
  OR2_X1 U3098 ( .A1(n3147), .A2(n3913), .ZN(n3075) );
  INV_X1 U3099 ( .A(n3075), .ZN(n2412) );
  NOR2_X1 U3100 ( .A1(n2413), .A2(n2412), .ZN(n2414) );
  OR2_X1 U3101 ( .A1(n2415), .A2(n2414), .ZN(n2416) );
  NAND2_X1 U3102 ( .A1(n3410), .A2(REG0_REG_10__SCAN_IN), .ZN(n2425) );
  INV_X1 U3103 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2418) );
  NAND2_X1 U3104 ( .A1(n2419), .A2(n4701), .ZN(n2420) );
  NAND2_X1 U3105 ( .A1(n2430), .A2(n2420), .ZN(n3748) );
  OR2_X1 U3106 ( .A1(n2658), .A2(n3748), .ZN(n2423) );
  INV_X1 U3107 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2421) );
  OR2_X1 U3108 ( .A1(n2312), .A2(n2421), .ZN(n2422) );
  NAND2_X1 U3109 ( .A1(n2436), .A2(IR_REG_31__SCAN_IN), .ZN(n2426) );
  XNOR2_X1 U3110 ( .A(n2426), .B(IR_REG_10__SCAN_IN), .ZN(n3963) );
  MUX2_X1 U3111 ( .A(DATAI_10_), .B(n3963), .S(n2512), .Z(n3747) );
  NOR2_X1 U3112 ( .A1(n3909), .A2(n3747), .ZN(n2427) );
  NAND2_X1 U3113 ( .A1(n3410), .A2(REG0_REG_11__SCAN_IN), .ZN(n2435) );
  INV_X1 U3114 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3314) );
  OR2_X1 U3115 ( .A1(n2311), .A2(n3314), .ZN(n2434) );
  INV_X1 U3116 ( .A(n2428), .ZN(n2442) );
  NAND2_X1 U3117 ( .A1(n2430), .A2(n2429), .ZN(n2431) );
  NAND2_X1 U3118 ( .A1(n2442), .A2(n2431), .ZN(n3567) );
  OR2_X1 U3119 ( .A1(n2658), .A2(n3567), .ZN(n2433) );
  INV_X1 U3120 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3568) );
  OR2_X1 U3121 ( .A1(n2312), .A2(n3568), .ZN(n2432) );
  OR2_X1 U3122 ( .A1(n2436), .A2(IR_REG_10__SCAN_IN), .ZN(n2437) );
  NAND2_X1 U3123 ( .A1(n2437), .A2(IR_REG_31__SCAN_IN), .ZN(n2439) );
  INV_X1 U3124 ( .A(IR_REG_11__SCAN_IN), .ZN(n2438) );
  OR2_X1 U3125 ( .A1(n2439), .A2(n2438), .ZN(n2440) );
  NAND2_X1 U3126 ( .A1(n2439), .A2(n2438), .ZN(n2448) );
  MUX2_X1 U3127 ( .A(DATAI_11_), .B(n3957), .S(n2512), .Z(n3374) );
  NAND2_X1 U3128 ( .A1(n3745), .A2(n3374), .ZN(n3295) );
  NAND2_X1 U3129 ( .A1(n3908), .A2(n3372), .ZN(n3297) );
  NAND2_X1 U3130 ( .A1(n3410), .A2(REG0_REG_12__SCAN_IN), .ZN(n2447) );
  INV_X1 U3131 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3289) );
  OR2_X1 U3132 ( .A1(n2312), .A2(n3289), .ZN(n2446) );
  INV_X1 U3133 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2441) );
  NAND2_X1 U3134 ( .A1(n2442), .A2(n2441), .ZN(n2443) );
  NAND2_X1 U3135 ( .A1(n2453), .A2(n2443), .ZN(n3785) );
  OR2_X1 U3136 ( .A1(n2658), .A2(n3785), .ZN(n2445) );
  INV_X1 U3137 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3351) );
  OR2_X1 U3138 ( .A1(n2311), .A2(n3351), .ZN(n2444) );
  NAND2_X1 U3139 ( .A1(n2448), .A2(IR_REG_31__SCAN_IN), .ZN(n2449) );
  XNOR2_X1 U3140 ( .A(n2449), .B(IR_REG_12__SCAN_IN), .ZN(n3967) );
  MUX2_X1 U3141 ( .A(n4657), .B(n4506), .S(n2512), .Z(n3578) );
  NAND2_X1 U3142 ( .A1(n3287), .A2(n2450), .ZN(n2451) );
  NAND2_X1 U3143 ( .A1(n3410), .A2(REG0_REG_13__SCAN_IN), .ZN(n2458) );
  INV_X1 U3144 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4412) );
  OR2_X1 U3145 ( .A1(n2312), .A2(n4412), .ZN(n2457) );
  NAND2_X1 U3146 ( .A1(n2453), .A2(n2452), .ZN(n2454) );
  NAND2_X1 U3147 ( .A1(n2464), .A2(n2454), .ZN(n3847) );
  OR2_X1 U31480 ( .A1(n2658), .A2(n3847), .ZN(n2456) );
  INV_X1 U31490 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3382) );
  OR2_X1 U3150 ( .A1(n2311), .A2(n3382), .ZN(n2455) );
  INV_X1 U3151 ( .A(DATAI_13_), .ZN(n2461) );
  NAND2_X1 U3152 ( .A1(n2459), .A2(IR_REG_31__SCAN_IN), .ZN(n2460) );
  XNOR2_X1 U3153 ( .A(n2460), .B(IR_REG_13__SCAN_IN), .ZN(n3956) );
  MUX2_X1 U3154 ( .A(n2461), .B(n4505), .S(n2512), .Z(n3588) );
  INV_X1 U3155 ( .A(n3588), .ZN(n3844) );
  NAND2_X1 U3156 ( .A1(n3410), .A2(REG0_REG_14__SCAN_IN), .ZN(n2470) );
  INV_X1 U3157 ( .A(REG1_REG_14__SCAN_IN), .ZN(n3338) );
  OR2_X1 U3158 ( .A1(n2311), .A2(n3338), .ZN(n2469) );
  INV_X1 U3159 ( .A(n2463), .ZN(n2475) );
  NAND2_X1 U3160 ( .A1(n2464), .A2(n4660), .ZN(n2465) );
  NAND2_X1 U3161 ( .A1(n2475), .A2(n2465), .ZN(n3729) );
  OR2_X1 U3162 ( .A1(n2658), .A2(n3729), .ZN(n2468) );
  INV_X1 U3163 ( .A(REG2_REG_14__SCAN_IN), .ZN(n2466) );
  OR2_X1 U3164 ( .A1(n2312), .A2(n2466), .ZN(n2467) );
  OR2_X1 U3165 ( .A1(n2471), .A2(n2378), .ZN(n2472) );
  XNOR2_X1 U3166 ( .A(n2472), .B(IR_REG_14__SCAN_IN), .ZN(n4503) );
  MUX2_X1 U3167 ( .A(DATAI_14_), .B(n4503), .S(n2512), .Z(n3726) );
  NAND2_X1 U3168 ( .A1(n3593), .A2(n3726), .ZN(n3421) );
  NAND2_X1 U3169 ( .A1(n3905), .A2(n3591), .ZN(n3492) );
  NAND2_X1 U3170 ( .A1(n3421), .A2(n3492), .ZN(n3472) );
  NAND2_X1 U3171 ( .A1(n3200), .A2(n2257), .ZN(n3261) );
  NAND2_X1 U3172 ( .A1(n3410), .A2(REG0_REG_15__SCAN_IN), .ZN(n2481) );
  INV_X1 U3173 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2473) );
  OR2_X1 U3174 ( .A1(n2312), .A2(n2473), .ZN(n2480) );
  INV_X1 U3175 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2474) );
  NAND2_X1 U3176 ( .A1(n2475), .A2(n2474), .ZN(n2476) );
  NAND2_X1 U3177 ( .A1(n2477), .A2(n2476), .ZN(n3894) );
  OR2_X1 U3178 ( .A1(n2658), .A2(n3894), .ZN(n2479) );
  INV_X1 U3179 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3392) );
  OR2_X1 U3180 ( .A1(n2311), .A2(n3392), .ZN(n2478) );
  INV_X1 U3181 ( .A(DATAI_15_), .ZN(n4681) );
  OR2_X1 U3182 ( .A1(n2483), .A2(n2482), .ZN(n2484) );
  MUX2_X1 U3183 ( .A(n4681), .B(n4502), .S(n2512), .Z(n3596) );
  NAND2_X1 U3184 ( .A1(n4287), .A2(n4296), .ZN(n3429) );
  INV_X1 U3185 ( .A(n4296), .ZN(n3608) );
  NAND2_X1 U3186 ( .A1(n3904), .A2(n3608), .ZN(n3493) );
  INV_X1 U3187 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4686) );
  NAND2_X1 U3188 ( .A1(n2489), .A2(n4686), .ZN(n2490) );
  AND2_X1 U3189 ( .A1(n2501), .A2(n2490), .ZN(n3812) );
  NAND2_X1 U3190 ( .A1(n2296), .A2(n3812), .ZN(n2495) );
  INV_X1 U3191 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4353) );
  OR2_X1 U3192 ( .A1(n2303), .A2(n4353), .ZN(n2494) );
  INV_X1 U3193 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4290) );
  OR2_X1 U3194 ( .A1(n2311), .A2(n4290), .ZN(n2493) );
  INV_X1 U3195 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2491) );
  OR2_X1 U3196 ( .A1(n2312), .A2(n2491), .ZN(n2492) );
  INV_X1 U3197 ( .A(DATAI_17_), .ZN(n2497) );
  OR2_X1 U3198 ( .A1(n2510), .A2(n2378), .ZN(n2496) );
  XNOR2_X1 U3199 ( .A(n2496), .B(IR_REG_17__SCAN_IN), .ZN(n4499) );
  INV_X1 U3200 ( .A(n4499), .ZN(n4463) );
  MUX2_X1 U3201 ( .A(n2497), .B(n4463), .S(n2045), .Z(n3616) );
  NOR2_X1 U3202 ( .A1(n3400), .A2(n2498), .ZN(n2499) );
  NOR2_X1 U3203 ( .A1(n2499), .A2(n2246), .ZN(n4171) );
  INV_X1 U3204 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2500) );
  INV_X1 U3205 ( .A(n2513), .ZN(n2514) );
  NAND2_X1 U3206 ( .A1(n2501), .A2(n2500), .ZN(n2502) );
  NAND2_X1 U3207 ( .A1(n2514), .A2(n2502), .ZN(n4184) );
  OR2_X1 U3208 ( .A1(n4184), .A2(n2658), .ZN(n2508) );
  INV_X1 U3209 ( .A(REG0_REG_18__SCAN_IN), .ZN(n2503) );
  OR2_X1 U32100 ( .A1(n2303), .A2(n2503), .ZN(n2505) );
  INV_X1 U32110 ( .A(REG1_REG_18__SCAN_IN), .ZN(n3978) );
  OR2_X1 U32120 ( .A1(n2311), .A2(n3978), .ZN(n2504) );
  AND2_X1 U32130 ( .A1(n2505), .A2(n2504), .ZN(n2507) );
  NAND2_X1 U32140 ( .A1(n3409), .A2(REG2_REG_18__SCAN_IN), .ZN(n2506) );
  NAND2_X1 U32150 ( .A1(n2518), .A2(IR_REG_31__SCAN_IN), .ZN(n2511) );
  XNOR2_X1 U32160 ( .A(n2511), .B(IR_REG_18__SCAN_IN), .ZN(n3954) );
  MUX2_X1 U32170 ( .A(DATAI_18_), .B(n3954), .S(n2319), .Z(n4175) );
  NAND2_X1 U32180 ( .A1(n4156), .A2(n4175), .ZN(n4151) );
  NAND2_X1 U32190 ( .A1(n4284), .A2(n4181), .ZN(n4152) );
  NAND2_X1 U32200 ( .A1(n4151), .A2(n4152), .ZN(n4174) );
  INV_X1 U32210 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4277) );
  INV_X1 U32220 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4685) );
  NAND2_X1 U32230 ( .A1(n2514), .A2(n4685), .ZN(n2515) );
  NAND2_X1 U32240 ( .A1(n2521), .A2(n2515), .ZN(n4165) );
  OR2_X1 U32250 ( .A1(n4165), .A2(n2658), .ZN(n2517) );
  AOI22_X1 U32260 ( .A1(n3409), .A2(REG2_REG_19__SCAN_IN), .B1(n3410), .B2(
        REG0_REG_19__SCAN_IN), .ZN(n2516) );
  OAI211_X1 U32270 ( .C1(n2311), .C2(n4277), .A(n2517), .B(n2516), .ZN(n4176)
         );
  INV_X1 U32280 ( .A(n2610), .ZN(n2519) );
  MUX2_X1 U32290 ( .A(DATAI_19_), .B(n4360), .S(n2319), .Z(n3758) );
  NAND2_X1 U32300 ( .A1(n4176), .A2(n3758), .ZN(n2520) );
  INV_X1 U32310 ( .A(n4176), .ZN(n3835) );
  INV_X1 U32320 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4669) );
  NAND2_X1 U32330 ( .A1(n2521), .A2(n4669), .ZN(n2522) );
  NAND2_X1 U32340 ( .A1(n2528), .A2(n2522), .ZN(n4141) );
  OR2_X1 U32350 ( .A1(n4141), .A2(n2658), .ZN(n2527) );
  INV_X1 U32360 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4273) );
  NAND2_X1 U32370 ( .A1(n3409), .A2(REG2_REG_20__SCAN_IN), .ZN(n2524) );
  NAND2_X1 U32380 ( .A1(n3410), .A2(REG0_REG_20__SCAN_IN), .ZN(n2523) );
  OAI211_X1 U32390 ( .C1(n4273), .C2(n2311), .A(n2524), .B(n2523), .ZN(n2525)
         );
  INV_X1 U32400 ( .A(n2525), .ZN(n2526) );
  NAND2_X1 U32410 ( .A1(n2333), .A2(DATAI_20_), .ZN(n4140) );
  NAND2_X1 U32420 ( .A1(n4120), .A2(n4140), .ZN(n3463) );
  INV_X1 U32430 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3766) );
  INV_X1 U32440 ( .A(n2537), .ZN(n2538) );
  NAND2_X1 U32450 ( .A1(n2528), .A2(n3766), .ZN(n2529) );
  NAND2_X1 U32460 ( .A1(n4117), .A2(n2296), .ZN(n2534) );
  INV_X1 U32470 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4268) );
  NAND2_X1 U32480 ( .A1(n3410), .A2(REG0_REG_21__SCAN_IN), .ZN(n2531) );
  NAND2_X1 U32490 ( .A1(n3409), .A2(REG2_REG_21__SCAN_IN), .ZN(n2530) );
  OAI211_X1 U32500 ( .C1(n2311), .C2(n4268), .A(n2531), .B(n2530), .ZN(n2532)
         );
  INV_X1 U32510 ( .A(n2532), .ZN(n2533) );
  INV_X1 U32520 ( .A(n4133), .ZN(n3902) );
  INV_X1 U32530 ( .A(DATAI_21_), .ZN(n4540) );
  NAND2_X1 U32540 ( .A1(n3902), .A2(n4260), .ZN(n2536) );
  INV_X1 U32550 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3855) );
  NAND2_X1 U32560 ( .A1(n2538), .A2(n3855), .ZN(n2539) );
  NAND2_X1 U32570 ( .A1(n2550), .A2(n2539), .ZN(n3854) );
  OR2_X1 U32580 ( .A1(n3854), .A2(n2658), .ZN(n2544) );
  INV_X1 U32590 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4258) );
  NAND2_X1 U32600 ( .A1(n3410), .A2(REG0_REG_22__SCAN_IN), .ZN(n2541) );
  NAND2_X1 U32610 ( .A1(n3409), .A2(REG2_REG_22__SCAN_IN), .ZN(n2540) );
  OAI211_X1 U32620 ( .C1(n2311), .C2(n4258), .A(n2541), .B(n2540), .ZN(n2542)
         );
  INV_X1 U32630 ( .A(n2542), .ZN(n2543) );
  INV_X1 U32640 ( .A(DATAI_22_), .ZN(n2545) );
  NOR2_X1 U32650 ( .A1(n2045), .A2(n2545), .ZN(n2546) );
  NAND2_X1 U32660 ( .A1(n4265), .A2(n2546), .ZN(n4076) );
  INV_X1 U32670 ( .A(n4265), .ZN(n4116) );
  NAND2_X1 U32680 ( .A1(n4116), .A2(n4095), .ZN(n2644) );
  NAND2_X1 U32690 ( .A1(n4076), .A2(n2644), .ZN(n4100) );
  NAND2_X1 U32700 ( .A1(n4101), .A2(n4100), .ZN(n4102) );
  NAND2_X1 U32710 ( .A1(n4102), .A2(n2065), .ZN(n4072) );
  INV_X1 U32720 ( .A(DATAI_23_), .ZN(n2547) );
  NOR2_X1 U32730 ( .A1(n2045), .A2(n2547), .ZN(n3644) );
  INV_X1 U32740 ( .A(REG3_REG_23__SCAN_IN), .ZN(n2549) );
  NAND2_X1 U32750 ( .A1(n2550), .A2(n2549), .ZN(n2551) );
  NAND2_X1 U32760 ( .A1(n2558), .A2(n2551), .ZN(n4085) );
  OR2_X1 U32770 ( .A1(n4085), .A2(n2658), .ZN(n2556) );
  INV_X1 U32780 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4253) );
  NAND2_X1 U32790 ( .A1(n3409), .A2(REG2_REG_23__SCAN_IN), .ZN(n2553) );
  NAND2_X1 U32800 ( .A1(n3410), .A2(REG0_REG_23__SCAN_IN), .ZN(n2552) );
  OAI211_X1 U32810 ( .C1(n4253), .C2(n2311), .A(n2553), .B(n2552), .ZN(n2554)
         );
  INV_X1 U32820 ( .A(n2554), .ZN(n2555) );
  OR2_X1 U32830 ( .A1(n3644), .A2(n4243), .ZN(n2557) );
  NAND2_X1 U32840 ( .A1(n4072), .A2(n2557), .ZN(n4058) );
  NAND2_X1 U32850 ( .A1(n4243), .A2(n3644), .ZN(n4057) );
  INV_X1 U32860 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4698) );
  NAND2_X1 U32870 ( .A1(n2558), .A2(n4698), .ZN(n2559) );
  AND2_X1 U32880 ( .A1(n2570), .A2(n2559), .ZN(n4064) );
  NAND2_X1 U32890 ( .A1(n4064), .A2(n2296), .ZN(n2564) );
  INV_X1 U32900 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4249) );
  NAND2_X1 U32910 ( .A1(n3409), .A2(REG2_REG_24__SCAN_IN), .ZN(n2561) );
  NAND2_X1 U32920 ( .A1(n3410), .A2(REG0_REG_24__SCAN_IN), .ZN(n2560) );
  OAI211_X1 U32930 ( .C1(n4249), .C2(n2311), .A(n2561), .B(n2560), .ZN(n2562)
         );
  INV_X1 U32940 ( .A(n2562), .ZN(n2563) );
  NAND2_X1 U32950 ( .A1(n2333), .A2(DATAI_24_), .ZN(n3823) );
  OR2_X1 U32960 ( .A1(n4050), .A2(n3823), .ZN(n2565) );
  AND2_X1 U32970 ( .A1(n4057), .A2(n2565), .ZN(n2566) );
  NAND2_X1 U32980 ( .A1(n4058), .A2(n2566), .ZN(n2568) );
  NAND2_X1 U32990 ( .A1(n4050), .A2(n3823), .ZN(n2567) );
  INV_X1 U33000 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4542) );
  NAND2_X1 U33010 ( .A1(n2570), .A2(n4542), .ZN(n2571) );
  NAND2_X1 U33020 ( .A1(n2580), .A2(n2571), .ZN(n3793) );
  INV_X1 U33030 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4240) );
  NAND2_X1 U33040 ( .A1(n3409), .A2(REG2_REG_25__SCAN_IN), .ZN(n2573) );
  NAND2_X1 U33050 ( .A1(n3410), .A2(REG0_REG_25__SCAN_IN), .ZN(n2572) );
  OAI211_X1 U33060 ( .C1(n4240), .C2(n2311), .A(n2573), .B(n2572), .ZN(n2574)
         );
  INV_X1 U33070 ( .A(n2574), .ZN(n2575) );
  INV_X1 U33080 ( .A(DATAI_25_), .ZN(n4658) );
  NOR2_X1 U33090 ( .A1(n4063), .A2(n4233), .ZN(n2578) );
  NAND2_X1 U33100 ( .A1(n4063), .A2(n4233), .ZN(n2577) );
  INV_X1 U33110 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2579) );
  NAND2_X1 U33120 ( .A1(n2580), .A2(n2579), .ZN(n2581) );
  NAND2_X1 U33130 ( .A1(n4033), .A2(n2296), .ZN(n2586) );
  INV_X1 U33140 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4231) );
  NAND2_X1 U33150 ( .A1(n3409), .A2(REG2_REG_26__SCAN_IN), .ZN(n2583) );
  NAND2_X1 U33160 ( .A1(n3410), .A2(REG0_REG_26__SCAN_IN), .ZN(n2582) );
  OAI211_X1 U33170 ( .C1(n4231), .C2(n2311), .A(n2583), .B(n2582), .ZN(n2584)
         );
  INV_X1 U33180 ( .A(n2584), .ZN(n2585) );
  NAND2_X1 U33190 ( .A1(n2333), .A2(DATAI_26_), .ZN(n4032) );
  XNOR2_X1 U33200 ( .A(n2598), .B(REG3_REG_27__SCAN_IN), .ZN(n4011) );
  NAND2_X1 U33210 ( .A1(n4011), .A2(n2296), .ZN(n2592) );
  INV_X1 U33220 ( .A(REG1_REG_27__SCAN_IN), .ZN(n2589) );
  NAND2_X1 U33230 ( .A1(n3409), .A2(REG2_REG_27__SCAN_IN), .ZN(n2588) );
  NAND2_X1 U33240 ( .A1(n3410), .A2(REG0_REG_27__SCAN_IN), .ZN(n2587) );
  OAI211_X1 U33250 ( .C1(n2589), .C2(n2311), .A(n2588), .B(n2587), .ZN(n2590)
         );
  INV_X1 U33260 ( .A(n2590), .ZN(n2591) );
  NAND2_X1 U33270 ( .A1(n2333), .A2(DATAI_27_), .ZN(n4221) );
  NAND2_X1 U33280 ( .A1(n3674), .A2(n4221), .ZN(n2593) );
  NAND2_X1 U33290 ( .A1(n4004), .A2(n2593), .ZN(n2595) );
  INV_X1 U33300 ( .A(n4221), .ZN(n3713) );
  NAND2_X1 U33310 ( .A1(n4028), .A2(n3713), .ZN(n2594) );
  NAND2_X1 U33320 ( .A1(n2595), .A2(n2594), .ZN(n2705) );
  INV_X1 U33330 ( .A(REG3_REG_27__SCAN_IN), .ZN(n2597) );
  INV_X1 U33340 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2596) );
  OAI21_X1 U33350 ( .B1(n2598), .B2(n2597), .A(n2596), .ZN(n2601) );
  INV_X1 U33360 ( .A(n2598), .ZN(n2600) );
  AND2_X1 U33370 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG3_REG_28__SCAN_IN), .ZN(
        n2599) );
  NAND2_X1 U33380 ( .A1(n2600), .A2(n2599), .ZN(n3997) );
  NAND2_X1 U33390 ( .A1(n2601), .A2(n3997), .ZN(n3699) );
  INV_X1 U33400 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2604) );
  NAND2_X1 U33410 ( .A1(n3409), .A2(REG2_REG_28__SCAN_IN), .ZN(n2603) );
  NAND2_X1 U33420 ( .A1(n3410), .A2(REG0_REG_28__SCAN_IN), .ZN(n2602) );
  OAI211_X1 U33430 ( .C1(n2604), .C2(n2311), .A(n2603), .B(n2602), .ZN(n2605)
         );
  INV_X1 U33440 ( .A(n2605), .ZN(n2606) );
  INV_X1 U33450 ( .A(DATAI_28_), .ZN(n2608) );
  NOR2_X1 U33460 ( .A1(n2045), .A2(n2608), .ZN(n3689) );
  NAND2_X1 U33470 ( .A1(n3684), .A2(n3689), .ZN(n3417) );
  INV_X1 U33480 ( .A(n3689), .ZN(n3700) );
  NAND2_X1 U33490 ( .A1(n4224), .A2(n3700), .ZN(n3413) );
  NAND2_X1 U33500 ( .A1(n3417), .A2(n3413), .ZN(n3482) );
  XNOR2_X1 U33510 ( .A(n2705), .B(n3482), .ZN(n3710) );
  NOR2_X1 U33520 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2609) );
  NAND2_X1 U3353 ( .A1(n2610), .A2(n2609), .ZN(n2618) );
  NAND2_X1 U33540 ( .A1(n2618), .A2(IR_REG_31__SCAN_IN), .ZN(n2612) );
  INV_X1 U3355 ( .A(IR_REG_19__SCAN_IN), .ZN(n2613) );
  NAND2_X1 U3356 ( .A1(n2614), .A2(n2613), .ZN(n2615) );
  INV_X1 U3357 ( .A(n2673), .ZN(n2619) );
  NAND2_X1 U3358 ( .A1(n2619), .A2(IR_REG_31__SCAN_IN), .ZN(n2621) );
  INV_X1 U3359 ( .A(IR_REG_22__SCAN_IN), .ZN(n2620) );
  XNOR2_X1 U3360 ( .A(n2843), .B(n3562), .ZN(n2622) );
  INV_X1 U3361 ( .A(n4360), .ZN(n3982) );
  NAND2_X1 U3362 ( .A1(n2622), .A2(n3982), .ZN(n4137) );
  AND2_X1 U3363 ( .A1(n2623), .A2(n4360), .ZN(n2912) );
  INV_X1 U3364 ( .A(n4519), .ZN(n3309) );
  INV_X1 U3365 ( .A(n4521), .ZN(n4306) );
  INV_X1 U3366 ( .A(n2852), .ZN(n2981) );
  NAND2_X1 U3367 ( .A1(n2981), .A2(n2987), .ZN(n3496) );
  NAND2_X1 U3368 ( .A1(n2731), .A2(n3502), .ZN(n3010) );
  NAND2_X1 U3369 ( .A1(n2965), .A2(n3011), .ZN(n3507) );
  NAND2_X1 U3370 ( .A1(n2959), .A2(n3016), .ZN(n3504) );
  NAND2_X1 U3371 ( .A1(n3010), .A2(n3452), .ZN(n3009) );
  NAND2_X1 U3372 ( .A1(n3009), .A2(n3507), .ZN(n2995) );
  INV_X1 U3373 ( .A(n3508), .ZN(n2624) );
  AND2_X1 U3374 ( .A1(n3914), .A2(n3133), .ZN(n3054) );
  NAND2_X1 U3375 ( .A1(n3125), .A2(n3126), .ZN(n3487) );
  NAND2_X1 U3376 ( .A1(n3913), .A2(n3143), .ZN(n3510) );
  NAND2_X1 U3377 ( .A1(n3083), .A2(n3510), .ZN(n2626) );
  NAND2_X1 U3378 ( .A1(n3144), .A2(n3147), .ZN(n3514) );
  NAND2_X1 U3379 ( .A1(n2626), .A2(n3514), .ZN(n3065) );
  INV_X1 U3380 ( .A(n2627), .ZN(n2628) );
  NAND2_X1 U3381 ( .A1(n3238), .A2(n3252), .ZN(n3520) );
  NAND2_X1 U3382 ( .A1(n3911), .A2(n3236), .ZN(n3517) );
  INV_X1 U3383 ( .A(n3154), .ZN(n2629) );
  NAND2_X1 U3384 ( .A1(n2629), .A2(n2061), .ZN(n2630) );
  NAND2_X1 U3385 ( .A1(n3276), .A2(n3280), .ZN(n3521) );
  NAND2_X1 U3386 ( .A1(n2630), .A2(n3521), .ZN(n3167) );
  NAND2_X1 U3387 ( .A1(n3909), .A2(n3365), .ZN(n3486) );
  NAND2_X1 U3388 ( .A1(n3308), .A2(n3747), .ZN(n3490) );
  NAND2_X1 U3389 ( .A1(n3907), .A2(n3578), .ZN(n3316) );
  NAND2_X1 U3390 ( .A1(n3906), .A2(n3588), .ZN(n2631) );
  NAND2_X1 U3391 ( .A1(n3316), .A2(n2631), .ZN(n3525) );
  INV_X1 U3392 ( .A(n3297), .ZN(n3527) );
  NOR2_X1 U3393 ( .A1(n3525), .A2(n3527), .ZN(n2632) );
  NAND2_X1 U3394 ( .A1(n3580), .A2(n3782), .ZN(n3318) );
  NAND2_X1 U3395 ( .A1(n3295), .A2(n3318), .ZN(n2635) );
  INV_X1 U3396 ( .A(n3525), .ZN(n2634) );
  NOR2_X1 U3397 ( .A1(n3906), .A2(n3588), .ZN(n2633) );
  AOI21_X1 U3398 ( .B1(n2635), .B2(n2634), .A(n2633), .ZN(n3528) );
  NAND2_X1 U3399 ( .A1(n3428), .A2(n2163), .ZN(n2636) );
  NAND2_X1 U3400 ( .A1(n2636), .A2(n3421), .ZN(n3258) );
  INV_X1 U3401 ( .A(n3258), .ZN(n2638) );
  NAND2_X1 U3402 ( .A1(n4300), .A2(n2486), .ZN(n3427) );
  NAND2_X1 U3403 ( .A1(n2487), .A2(n3596), .ZN(n3491) );
  NAND2_X1 U3404 ( .A1(n3427), .A2(n3491), .ZN(n3454) );
  NAND2_X1 U3405 ( .A1(n2638), .A2(n2637), .ZN(n3259) );
  NAND2_X1 U3406 ( .A1(n3259), .A2(n3491), .ZN(n4206) );
  INV_X1 U3407 ( .A(n4150), .ZN(n2639) );
  NAND2_X1 U3408 ( .A1(n4176), .A2(n4162), .ZN(n3464) );
  NAND2_X1 U3409 ( .A1(n3464), .A2(n4152), .ZN(n3422) );
  NAND2_X1 U3410 ( .A1(n2639), .A2(n3424), .ZN(n4128) );
  NAND2_X1 U3411 ( .A1(n4262), .A2(n4140), .ZN(n3423) );
  INV_X1 U3412 ( .A(n3423), .ZN(n2643) );
  NAND2_X1 U3413 ( .A1(n4294), .A2(n4282), .ZN(n4149) );
  AND2_X1 U3414 ( .A1(n4151), .A2(n4149), .ZN(n2640) );
  OR2_X1 U3415 ( .A1(n4176), .A2(n4162), .ZN(n3465) );
  OAI21_X1 U3416 ( .B1(n3422), .B2(n2640), .A(n3465), .ZN(n4126) );
  NOR2_X1 U3417 ( .A1(n4262), .A2(n4140), .ZN(n2641) );
  OR2_X1 U3418 ( .A1(n4126), .A2(n2641), .ZN(n2642) );
  NAND2_X1 U3419 ( .A1(n2642), .A2(n3423), .ZN(n3535) );
  OAI21_X1 U3420 ( .B1(n4128), .B2(n2643), .A(n3535), .ZN(n4108) );
  NAND2_X1 U3421 ( .A1(n4133), .A2(n4260), .ZN(n3462) );
  AND2_X1 U3422 ( .A1(n4076), .A2(n3462), .ZN(n3536) );
  INV_X1 U3423 ( .A(n3536), .ZN(n2646) );
  INV_X1 U3424 ( .A(n3644), .ZN(n4083) );
  NAND2_X1 U3425 ( .A1(n4243), .A2(n4083), .ZN(n3448) );
  NAND2_X1 U3426 ( .A1(n3448), .A2(n2644), .ZN(n3485) );
  NOR2_X1 U3427 ( .A1(n4133), .A2(n4260), .ZN(n4073) );
  AND2_X1 U3428 ( .A1(n4076), .A2(n4073), .ZN(n2645) );
  NOR2_X1 U3429 ( .A1(n3485), .A2(n2645), .ZN(n3434) );
  OAI21_X1 U3430 ( .B1(n4108), .B2(n2646), .A(n3434), .ZN(n2647) );
  INV_X1 U3431 ( .A(n4243), .ZN(n4067) );
  NAND2_X1 U3432 ( .A1(n4067), .A2(n3644), .ZN(n3449) );
  NAND2_X1 U3433 ( .A1(n2647), .A2(n3449), .ZN(n4055) );
  NOR2_X1 U3434 ( .A1(n4234), .A2(n3823), .ZN(n3447) );
  INV_X1 U3435 ( .A(n4032), .ZN(n2648) );
  NAND2_X1 U3436 ( .A1(n4237), .A2(n2648), .ZN(n2649) );
  INV_X1 U3437 ( .A(n4063), .ZN(n4246) );
  NAND2_X1 U3438 ( .A1(n4246), .A2(n4233), .ZN(n4022) );
  INV_X1 U3439 ( .A(n4233), .ZN(n4045) );
  NAND2_X1 U3440 ( .A1(n4063), .A2(n4045), .ZN(n3445) );
  NAND2_X1 U3441 ( .A1(n4234), .A2(n3823), .ZN(n4038) );
  NAND2_X1 U3442 ( .A1(n3445), .A2(n4038), .ZN(n4023) );
  AND2_X1 U3443 ( .A1(n4046), .A2(n4032), .ZN(n3415) );
  AOI21_X1 U3444 ( .B1(n2650), .B2(n4023), .A(n3415), .ZN(n3544) );
  XNOR2_X1 U3445 ( .A(n4028), .B(n4221), .ZN(n4005) );
  OR2_X1 U3446 ( .A1(n4028), .A2(n4221), .ZN(n3416) );
  XOR2_X1 U3447 ( .A(n3482), .B(n2708), .Z(n2653) );
  NAND2_X1 U3448 ( .A1(n3562), .A2(n4360), .ZN(n2652) );
  INV_X1 U3449 ( .A(n3459), .ZN(n4359) );
  NAND2_X1 U3450 ( .A1(n4359), .A2(n2651), .ZN(n3443) );
  NAND2_X1 U3451 ( .A1(n2653), .A2(n4203), .ZN(n3697) );
  NOR2_X1 U3452 ( .A1(n2654), .A2(n2378), .ZN(n2655) );
  MUX2_X1 U3453 ( .A(n2378), .B(n2655), .S(IR_REG_28__SCAN_IN), .Z(n2657) );
  OR2_X1 U3454 ( .A1(n2657), .A2(n2656), .ZN(n2920) );
  NAND2_X1 U3455 ( .A1(n3562), .A2(n4359), .ZN(n2835) );
  NOR2_X2 U3456 ( .A1(n2920), .A2(n2835), .ZN(n4261) );
  OR2_X1 U3457 ( .A1(n3997), .A2(n2658), .ZN(n2663) );
  INV_X1 U34580 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2718) );
  NAND2_X1 U34590 ( .A1(n3409), .A2(REG2_REG_29__SCAN_IN), .ZN(n2660) );
  NAND2_X1 U3460 ( .A1(n3410), .A2(REG0_REG_29__SCAN_IN), .ZN(n2659) );
  OAI211_X1 U3461 ( .C1(n2718), .C2(n2311), .A(n2660), .B(n2659), .ZN(n2661)
         );
  INV_X1 U3462 ( .A(n2661), .ZN(n2662) );
  NAND2_X1 U3463 ( .A1(n2663), .A2(n2662), .ZN(n3901) );
  INV_X1 U3464 ( .A(n3901), .ZN(n3702) );
  INV_X1 U3465 ( .A(n2835), .ZN(n2772) );
  NAND2_X1 U3466 ( .A1(n2920), .A2(n2772), .ZN(n4293) );
  NAND2_X1 U34670 ( .A1(n2830), .A2(n3459), .ZN(n2834) );
  OR2_X1 U3468 ( .A1(n2834), .A2(n2623), .ZN(n4220) );
  OAI22_X1 U34690 ( .A1(n3702), .A2(n4293), .B1(n3700), .B2(n4220), .ZN(n2664)
         );
  AOI21_X1 U3470 ( .B1(n4261), .B2(n4028), .A(n2664), .ZN(n2665) );
  OAI21_X1 U34710 ( .B1(n3710), .B2(n4306), .A(n2666), .ZN(n2701) );
  NAND2_X1 U3472 ( .A1(n2671), .A2(IR_REG_31__SCAN_IN), .ZN(n2667) );
  MUX2_X1 U34730 ( .A(IR_REG_31__SCAN_IN), .B(n2667), .S(IR_REG_26__SCAN_IN), 
        .Z(n2668) );
  NAND2_X1 U3474 ( .A1(n2669), .A2(IR_REG_31__SCAN_IN), .ZN(n2670) );
  MUX2_X1 U34750 ( .A(IR_REG_31__SCAN_IN), .B(n2670), .S(IR_REG_25__SCAN_IN), 
        .Z(n2672) );
  NAND2_X1 U3476 ( .A1(n2672), .A2(n2671), .ZN(n2751) );
  NAND2_X1 U34770 ( .A1(n2751), .A2(B_REG_SCAN_IN), .ZN(n2675) );
  INV_X1 U3478 ( .A(IR_REG_23__SCAN_IN), .ZN(n2679) );
  MUX2_X1 U34790 ( .A(n2675), .B(B_REG_SCAN_IN), .S(n2678), .Z(n2676) );
  NAND2_X1 U3480 ( .A1(n2764), .A2(n2751), .ZN(n2768) );
  NAND2_X1 U34810 ( .A1(n2826), .A2(n2768), .ZN(n2694) );
  XNOR2_X1 U3482 ( .A(n2680), .B(n2679), .ZN(n2771) );
  NAND2_X1 U34830 ( .A1(n4519), .A2(n3459), .ZN(n2740) );
  AND2_X1 U3484 ( .A1(n2623), .A2(n3982), .ZN(n2833) );
  OR2_X1 U34850 ( .A1(n2835), .A2(n2833), .ZN(n2838) );
  NAND2_X1 U3486 ( .A1(n2740), .A2(n2838), .ZN(n2681) );
  NOR2_X1 U34870 ( .A1(n2860), .A2(n2681), .ZN(n2693) );
  NOR4_X1 U3488 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2685) );
  NOR4_X1 U34890 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2684) );
  NOR4_X1 U3490 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2683) );
  NOR4_X1 U34910 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2682) );
  NAND4_X1 U3492 ( .A1(n2685), .A2(n2684), .A3(n2683), .A4(n2682), .ZN(n2691)
         );
  NOR2_X1 U34930 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_3__SCAN_IN), .ZN(n2689) );
  NOR4_X1 U3494 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2688) );
  NOR4_X1 U34950 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2687) );
  NOR4_X1 U3496 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2686) );
  NAND4_X1 U34970 ( .A1(n2689), .A2(n2688), .A3(n2687), .A4(n2686), .ZN(n2690)
         );
  NOR2_X1 U3498 ( .A1(n2691), .A2(n2690), .ZN(n2692) );
  NAND3_X1 U34990 ( .A1(n2694), .A2(n2693), .A3(n2736), .ZN(n2700) );
  NAND2_X1 U3500 ( .A1(n2765), .A2(n2764), .ZN(n2695) );
  INV_X1 U35010 ( .A(n2738), .ZN(n2828) );
  MUX2_X1 U3502 ( .A(REG0_REG_28__SCAN_IN), .B(n2701), .S(n4529), .Z(n2697) );
  INV_X1 U35030 ( .A(n2697), .ZN(n2699) );
  INV_X1 U3504 ( .A(n2987), .ZN(n2910) );
  NAND2_X1 U35050 ( .A1(n2842), .A2(n2910), .ZN(n2989) );
  NOR2_X1 U35060 ( .A1(n2989), .A2(n2900), .ZN(n3017) );
  OR2_X2 U35070 ( .A1(n3018), .A2(n3048), .ZN(n3062) );
  OR2_X2 U35080 ( .A1(n3170), .A2(n3374), .ZN(n3302) );
  OR2_X2 U35090 ( .A1(n2051), .A2(n4296), .ZN(n4194) );
  INV_X1 U35100 ( .A(n3823), .ZN(n4242) );
  AND2_X1 U35110 ( .A1(n4009), .A2(n3689), .ZN(n2698) );
  OR2_X1 U35120 ( .A1(n2698), .A2(n2719), .ZN(n3706) );
  INV_X1 U35130 ( .A(n2834), .ZN(n2909) );
  NAND2_X1 U35140 ( .A1(n2699), .A2(n2250), .ZN(U3514) );
  MUX2_X1 U35150 ( .A(REG1_REG_28__SCAN_IN), .B(n2701), .S(n4535), .Z(n2702)
         );
  INV_X1 U35160 ( .A(n2702), .ZN(n2703) );
  NAND2_X1 U35170 ( .A1(n2703), .A2(n2249), .ZN(U3546) );
  NOR2_X1 U35180 ( .A1(n3684), .A2(n3700), .ZN(n2704) );
  NAND2_X1 U35190 ( .A1(n2333), .A2(DATAI_29_), .ZN(n3994) );
  XNOR2_X1 U35200 ( .A(n3901), .B(n3994), .ZN(n3483) );
  XNOR2_X1 U35210 ( .A(n2706), .B(n3483), .ZN(n3992) );
  INV_X1 U35220 ( .A(n3417), .ZN(n2707) );
  AOI21_X1 U35230 ( .B1(n2708), .B2(n3413), .A(n2707), .ZN(n2709) );
  XNOR2_X1 U35240 ( .A(n2709), .B(n3483), .ZN(n2715) );
  NOR2_X1 U35250 ( .A1(n2711), .A2(n2710), .ZN(n2921) );
  AOI21_X1 U35260 ( .B1(B_REG_SCAN_IN), .B2(n2921), .A(n4293), .ZN(n3987) );
  INV_X1 U35270 ( .A(REG1_REG_30__SCAN_IN), .ZN(n2714) );
  NAND2_X1 U35280 ( .A1(n3409), .A2(REG2_REG_30__SCAN_IN), .ZN(n2713) );
  NAND2_X1 U35290 ( .A1(n3410), .A2(REG0_REG_30__SCAN_IN), .ZN(n2712) );
  OAI211_X1 U35300 ( .C1(n2311), .C2(n2714), .A(n2713), .B(n2712), .ZN(n3900)
         );
  NAND2_X1 U35310 ( .A1(n4224), .A2(n4261), .ZN(n2716) );
  INV_X1 U35320 ( .A(n2719), .ZN(n2720) );
  INV_X1 U35330 ( .A(n3994), .ZN(n3414) );
  NAND2_X1 U35340 ( .A1(n2720), .A2(n3414), .ZN(n2721) );
  NAND2_X1 U35350 ( .A1(n4215), .A2(n2721), .ZN(n3998) );
  INV_X1 U35360 ( .A(n3998), .ZN(n2722) );
  INV_X1 U35370 ( .A(REG0_REG_29__SCAN_IN), .ZN(n2725) );
  MUX2_X1 U35380 ( .A(n2725), .B(n2724), .S(n4529), .Z(n2727) );
  NAND2_X1 U35390 ( .A1(n2727), .A2(n2726), .ZN(U3515) );
  INV_X2 U35400 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U35410 ( .A(n4497), .ZN(n2728) );
  INV_X2 U35420 ( .A(n3903), .ZN(U4043) );
  NAND2_X1 U35430 ( .A1(n2729), .A2(n3471), .ZN(n2730) );
  NAND2_X1 U35440 ( .A1(n3007), .A2(n2730), .ZN(n2905) );
  INV_X1 U35450 ( .A(n4137), .ZN(n2998) );
  NAND2_X1 U35460 ( .A1(n2905), .A2(n2998), .ZN(n2735) );
  OAI21_X1 U35470 ( .B1(n3471), .B2(n2732), .A(n2731), .ZN(n2733) );
  NAND2_X1 U35480 ( .A1(n2733), .A2(n4203), .ZN(n2734) );
  NAND2_X1 U35490 ( .A1(n2735), .A2(n2734), .ZN(n2903) );
  INV_X1 U35500 ( .A(n2838), .ZN(n2737) );
  NOR2_X1 U35510 ( .A1(n2860), .A2(n2737), .ZN(n2739) );
  NAND4_X1 U35520 ( .A1(n2827), .A2(n2739), .A3(n2738), .A4(n2826), .ZN(n2741)
         );
  INV_X1 U35530 ( .A(n4367), .ZN(n4106) );
  MUX2_X1 U35540 ( .A(REG2_REG_2__SCAN_IN), .B(n2903), .S(n4106), .Z(n2749) );
  NAND2_X1 U35550 ( .A1(n4187), .A2(n3982), .ZN(n4183) );
  XNOR2_X1 U35560 ( .A(n2989), .B(n2900), .ZN(n2941) );
  NOR2_X1 U35570 ( .A1(n4164), .A2(n2941), .ZN(n2748) );
  NAND2_X1 U35580 ( .A1(n4106), .A2(n4295), .ZN(n4015) );
  INV_X1 U35590 ( .A(n2843), .ZN(n2829) );
  NAND2_X1 U35600 ( .A1(n2829), .A2(n4360), .ZN(n3078) );
  INV_X1 U35610 ( .A(n3078), .ZN(n2742) );
  NAND2_X1 U35620 ( .A1(n4106), .A2(n2742), .ZN(n4147) );
  INV_X1 U35630 ( .A(n4147), .ZN(n4491) );
  NAND2_X1 U35640 ( .A1(n2905), .A2(n4491), .ZN(n2744) );
  INV_X1 U35650 ( .A(n4476), .ZN(n4486) );
  NAND2_X1 U35660 ( .A1(n4486), .A2(REG3_REG_2__SCAN_IN), .ZN(n2743) );
  OAI211_X1 U35670 ( .C1(n4015), .C2(n2888), .A(n2744), .B(n2743), .ZN(n2747)
         );
  NAND2_X1 U35680 ( .A1(n4106), .A2(n4283), .ZN(n3701) );
  NAND2_X1 U35690 ( .A1(n4012), .A2(n3917), .ZN(n2745) );
  OAI21_X1 U35700 ( .B1(n2965), .B2(n3701), .A(n2745), .ZN(n2746) );
  OR4_X1 U35710 ( .A1(n2749), .A2(n2748), .A3(n2747), .A4(n2746), .ZN(U3288)
         );
  NAND2_X1 U35720 ( .A1(U3149), .A2(DATAI_25_), .ZN(n2750) );
  OAI21_X1 U35730 ( .B1(n2751), .B2(U3149), .A(n2750), .ZN(U3327) );
  INV_X1 U35740 ( .A(DATAI_26_), .ZN(n4695) );
  NAND2_X1 U35750 ( .A1(n2752), .A2(STATE_REG_SCAN_IN), .ZN(n2753) );
  OAI21_X1 U35760 ( .B1(STATE_REG_SCAN_IN), .B2(n4695), .A(n2753), .ZN(U3326)
         );
  INV_X1 U35770 ( .A(DATAI_27_), .ZN(n4683) );
  NAND2_X1 U35780 ( .A1(n2921), .A2(STATE_REG_SCAN_IN), .ZN(n2754) );
  OAI21_X1 U35790 ( .B1(STATE_REG_SCAN_IN), .B2(n4683), .A(n2754), .ZN(U3325)
         );
  NAND2_X1 U35800 ( .A1(n3562), .A2(STATE_REG_SCAN_IN), .ZN(n2755) );
  OAI21_X1 U35810 ( .B1(STATE_REG_SCAN_IN), .B2(n2545), .A(n2755), .ZN(U3330)
         );
  INV_X1 U3582 ( .A(DATAI_29_), .ZN(n4661) );
  NAND2_X1 U3583 ( .A1(n2756), .A2(STATE_REG_SCAN_IN), .ZN(n2757) );
  OAI21_X1 U3584 ( .B1(STATE_REG_SCAN_IN), .B2(n4661), .A(n2757), .ZN(U3323)
         );
  INV_X1 U3585 ( .A(DATAI_24_), .ZN(n4636) );
  NAND2_X1 U3586 ( .A1(n2678), .A2(STATE_REG_SCAN_IN), .ZN(n2758) );
  OAI21_X1 U3587 ( .B1(STATE_REG_SCAN_IN), .B2(n4636), .A(n2758), .ZN(U3328)
         );
  INV_X1 U3588 ( .A(DATAI_31_), .ZN(n4537) );
  OR4_X1 U3589 ( .A1(n2759), .A2(IR_REG_30__SCAN_IN), .A3(n2378), .A4(U3149), 
        .ZN(n2760) );
  OAI21_X1 U3590 ( .B1(STATE_REG_SCAN_IN), .B2(n4537), .A(n2760), .ZN(U3321)
         );
  INV_X1 U3591 ( .A(n2920), .ZN(n2917) );
  NAND2_X1 U3592 ( .A1(n2917), .A2(STATE_REG_SCAN_IN), .ZN(n2761) );
  OAI21_X1 U3593 ( .B1(STATE_REG_SCAN_IN), .B2(n2608), .A(n2761), .ZN(U3324)
         );
  INV_X1 U3594 ( .A(n2860), .ZN(n2762) );
  INV_X1 U3595 ( .A(D_REG_0__SCAN_IN), .ZN(n2767) );
  AND2_X1 U3596 ( .A1(n4497), .A2(n2764), .ZN(n2766) );
  AOI22_X1 U3597 ( .A1(n4496), .A2(n2767), .B1(n2766), .B2(n2765), .ZN(U3458)
         );
  INV_X1 U3598 ( .A(D_REG_1__SCAN_IN), .ZN(n2770) );
  INV_X1 U3599 ( .A(n2768), .ZN(n2769) );
  AOI22_X1 U3600 ( .A1(n4496), .A2(n2770), .B1(n2769), .B2(n4497), .ZN(U3459)
         );
  OR2_X1 U3601 ( .A1(n2771), .A2(U3149), .ZN(n3564) );
  NAND2_X1 U3602 ( .A1(n2860), .A2(n3564), .ZN(n2780) );
  AOI21_X1 U3603 ( .B1(n2772), .B2(n2771), .A(n2319), .ZN(n2779) );
  INV_X1 U3604 ( .A(n2779), .ZN(n2773) );
  NOR2_X1 U3605 ( .A1(n4468), .A2(U4043), .ZN(U3148) );
  INV_X1 U3606 ( .A(n4366), .ZN(n2926) );
  MUX2_X1 U3607 ( .A(REG2_REG_2__SCAN_IN), .B(n2774), .S(n4366), .Z(n2778) );
  INV_X1 U3608 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2775) );
  AND2_X1 U3609 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n2776)
         );
  NAND2_X1 U3610 ( .A1(n3933), .A2(n2776), .ZN(n3932) );
  NAND2_X1 U3611 ( .A1(n3932), .A2(n2930), .ZN(n2777) );
  MUX2_X1 U3612 ( .A(REG2_REG_5__SCAN_IN), .B(n2346), .S(n2809), .Z(n2781) );
  INV_X1 U3613 ( .A(n2921), .ZN(n3918) );
  NOR2_X1 U3614 ( .A1(n2920), .A2(n3918), .ZN(n3559) );
  AOI211_X1 U3615 ( .C1(n2782), .C2(n2781), .A(n2804), .B(n4464), .ZN(n2785)
         );
  NAND2_X1 U3616 ( .A1(n3923), .A2(n2920), .ZN(n4475) );
  INV_X1 U3617 ( .A(REG3_REG_5__SCAN_IN), .ZN(n4655) );
  NOR2_X1 U3618 ( .A1(STATE_REG_SCAN_IN), .A2(n4655), .ZN(n3135) );
  AOI21_X1 U3619 ( .B1(n4468), .B2(ADDR_REG_5__SCAN_IN), .A(n3135), .ZN(n2783)
         );
  OAI21_X1 U3620 ( .B1(n4475), .B2(n2809), .A(n2783), .ZN(n2784) );
  NOR2_X1 U3621 ( .A1(n2785), .A2(n2784), .ZN(n2795) );
  XNOR2_X1 U3622 ( .A(n2809), .B(REG1_REG_5__SCAN_IN), .ZN(n2793) );
  XNOR2_X1 U3623 ( .A(n4366), .B(n2906), .ZN(n2929) );
  AND2_X1 U3624 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3929)
         );
  NAND2_X1 U3625 ( .A1(n3930), .A2(n3929), .ZN(n3928) );
  NAND2_X1 U3626 ( .A1(n3928), .A2(n2786), .ZN(n2928) );
  NAND2_X1 U3627 ( .A1(n2929), .A2(n2928), .ZN(n2927) );
  NAND2_X1 U3628 ( .A1(n4366), .A2(REG1_REG_2__SCAN_IN), .ZN(n2787) );
  NAND2_X1 U3629 ( .A1(n2927), .A2(n2787), .ZN(n2788) );
  XNOR2_X1 U3630 ( .A(n2788), .B(n2797), .ZN(n2800) );
  NAND2_X1 U3631 ( .A1(n2800), .A2(REG1_REG_3__SCAN_IN), .ZN(n2799) );
  NAND2_X1 U3632 ( .A1(n2788), .A2(n4365), .ZN(n2789) );
  NAND2_X1 U3633 ( .A1(n2799), .A2(n2789), .ZN(n2790) );
  INV_X1 U3634 ( .A(n2790), .ZN(n2791) );
  XNOR2_X1 U3635 ( .A(n2790), .B(n2948), .ZN(n2944) );
  NAND2_X1 U3636 ( .A1(n2944), .A2(REG1_REG_4__SCAN_IN), .ZN(n2943) );
  OAI21_X1 U3637 ( .B1(n2791), .B2(n2948), .A(n2943), .ZN(n2792) );
  NAND2_X1 U3638 ( .A1(n2792), .A2(n2793), .ZN(n2807) );
  OAI211_X1 U3639 ( .C1(n2793), .C2(n2792), .A(n4470), .B(n2807), .ZN(n2794)
         );
  NAND2_X1 U3640 ( .A1(n2795), .A2(n2794), .ZN(U3245) );
  XNOR2_X1 U3641 ( .A(n2796), .B(REG2_REG_3__SCAN_IN), .ZN(n2803) );
  INV_X1 U3642 ( .A(REG3_REG_3__SCAN_IN), .ZN(n4680) );
  NOR2_X1 U3643 ( .A1(STATE_REG_SCAN_IN), .A2(n4680), .ZN(n2971) );
  NOR2_X1 U3644 ( .A1(n4475), .A2(n2797), .ZN(n2798) );
  AOI211_X1 U3645 ( .C1(n4468), .C2(ADDR_REG_3__SCAN_IN), .A(n2971), .B(n2798), 
        .ZN(n2802) );
  OAI211_X1 U3646 ( .C1(REG1_REG_3__SCAN_IN), .C2(n2800), .A(n4470), .B(n2799), 
        .ZN(n2801) );
  OAI211_X1 U3647 ( .C1(n2803), .C2(n4464), .A(n2802), .B(n2801), .ZN(U3243)
         );
  XNOR2_X1 U3648 ( .A(n2819), .B(REG2_REG_6__SCAN_IN), .ZN(n2815) );
  INV_X1 U3649 ( .A(n4475), .ZN(n3927) );
  INV_X1 U3650 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2805) );
  NOR2_X1 U3651 ( .A1(STATE_REG_SCAN_IN), .A2(n2805), .ZN(n3146) );
  AOI21_X1 U3652 ( .B1(n4468), .B2(ADDR_REG_6__SCAN_IN), .A(n3146), .ZN(n2806)
         );
  INV_X1 U3653 ( .A(n2806), .ZN(n2813) );
  INV_X1 U3654 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3103) );
  INV_X1 U3655 ( .A(n4470), .ZN(n2810) );
  AOI211_X1 U3656 ( .C1(n2811), .C2(n3103), .A(n2816), .B(n2810), .ZN(n2812)
         );
  AOI211_X1 U3657 ( .C1(n3927), .C2(n4363), .A(n2813), .B(n2812), .ZN(n2814)
         );
  OAI21_X1 U3658 ( .B1(n2815), .B2(n4464), .A(n2814), .ZN(U3246) );
  MUX2_X1 U3659 ( .A(REG1_REG_7__SCAN_IN), .B(n2400), .S(n4362), .Z(n2817) );
  XNOR2_X1 U3660 ( .A(n2877), .B(n2817), .ZN(n2824) );
  INV_X1 U3661 ( .A(n4362), .ZN(n2875) );
  NOR2_X1 U3662 ( .A1(STATE_REG_SCAN_IN), .A2(n2396), .ZN(n3192) );
  AOI21_X1 U3663 ( .B1(n4468), .B2(ADDR_REG_7__SCAN_IN), .A(n3192), .ZN(n2818)
         );
  OAI21_X1 U3664 ( .B1(n4475), .B2(n2875), .A(n2818), .ZN(n2823) );
  MUX2_X1 U3665 ( .A(n2395), .B(REG2_REG_7__SCAN_IN), .S(n4362), .Z(n2820) );
  AOI211_X1 U3666 ( .C1(n2821), .C2(n2820), .A(n4464), .B(n2879), .ZN(n2822)
         );
  AOI211_X1 U3667 ( .C1(n4470), .C2(n2824), .A(n2823), .B(n2822), .ZN(n2825)
         );
  INV_X1 U3668 ( .A(n2825), .ZN(U3247) );
  NAND3_X1 U3669 ( .A1(n2828), .A2(n2827), .A3(n2826), .ZN(n2865) );
  INV_X1 U3670 ( .A(n2844), .ZN(n2831) );
  NAND2_X1 U3671 ( .A1(n4497), .A2(n2831), .ZN(n2832) );
  NOR2_X1 U3672 ( .A1(n3679), .A2(n2832), .ZN(n3560) );
  NAND2_X1 U3673 ( .A1(n2865), .A2(n3560), .ZN(n2968) );
  INV_X1 U3674 ( .A(n2968), .ZN(n2840) );
  OR2_X1 U3675 ( .A1(n2834), .A2(n2833), .ZN(n2836) );
  NAND2_X1 U3676 ( .A1(n2836), .A2(n2835), .ZN(n2858) );
  NAND2_X1 U3677 ( .A1(n2858), .A2(n4220), .ZN(n2837) );
  NAND2_X1 U3678 ( .A1(n2865), .A2(n2837), .ZN(n2839) );
  NAND2_X1 U3679 ( .A1(n2839), .A2(n2838), .ZN(n2967) );
  NOR3_X1 U3680 ( .A1(n2840), .A2(n2967), .A3(n2860), .ZN(n2895) );
  INV_X1 U3681 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3029) );
  NAND2_X4 U3682 ( .A1(n2841), .A2(n2843), .ZN(n3682) );
  NAND2_X1 U3683 ( .A1(n2958), .A2(n3034), .ZN(n2846) );
  XNOR2_X1 U3684 ( .A(n2889), .B(n2052), .ZN(n2856) );
  NAND2_X1 U3685 ( .A1(n2852), .A2(n2958), .ZN(n2849) );
  NAND2_X1 U3686 ( .A1(n2960), .A2(n2987), .ZN(n2848) );
  INV_X1 U3687 ( .A(n2841), .ZN(n2966) );
  NAND2_X1 U3688 ( .A1(n2966), .A2(REG1_REG_0__SCAN_IN), .ZN(n2850) );
  NAND2_X1 U3689 ( .A1(n2851), .A2(n2850), .ZN(n2869) );
  AOI22_X1 U3690 ( .A1(n2958), .A2(n2987), .B1(n2966), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2853) );
  OAI21_X1 U3691 ( .B1(n2981), .B2(n2964), .A(n2853), .ZN(n2871) );
  NAND2_X1 U3692 ( .A1(n2854), .A2(n2870), .ZN(n2855) );
  NAND2_X1 U3693 ( .A1(n2856), .A2(n2855), .ZN(n2892) );
  OR2_X1 U3694 ( .A1(n2860), .A2(n2858), .ZN(n2859) );
  OAI211_X1 U3695 ( .C1(n2847), .C2(n2855), .A(n2857), .B(n3897), .ZN(n2868)
         );
  OR2_X1 U3696 ( .A1(n2860), .A2(n4220), .ZN(n2861) );
  OR2_X1 U3697 ( .A1(n2865), .A2(n2861), .ZN(n2862) );
  NAND2_X1 U3698 ( .A1(n2862), .A2(n4476), .ZN(n3890) );
  NAND2_X1 U3699 ( .A1(n3560), .A2(n2917), .ZN(n2863) );
  NAND2_X1 U3700 ( .A1(n3560), .A2(n2920), .ZN(n2864) );
  OAI22_X1 U3701 ( .A1(n2981), .A2(n3856), .B1(n3857), .B2(n2885), .ZN(n2866)
         );
  AOI21_X1 U3702 ( .B1(n3034), .B2(n3890), .A(n2866), .ZN(n2867) );
  OAI211_X1 U3703 ( .C1(n2895), .C2(n3029), .A(n2868), .B(n2867), .ZN(U3219)
         );
  OAI21_X1 U3704 ( .B1(n2869), .B2(n2871), .A(n2870), .ZN(n2918) );
  OAI22_X1 U3705 ( .A1(n2918), .A2(n3884), .B1(n3857), .B2(n2902), .ZN(n2872)
         );
  AOI21_X1 U3706 ( .B1(n2987), .B2(n3890), .A(n2872), .ZN(n2873) );
  OAI21_X1 U3707 ( .B1(n2895), .B2(n2874), .A(n2873), .ZN(U3229) );
  NOR2_X1 U3708 ( .A1(n4362), .A2(REG1_REG_7__SCAN_IN), .ZN(n2876) );
  OAI22_X1 U3709 ( .A1(n2877), .A2(n2876), .B1(n2400), .B2(n2875), .ZN(n3960)
         );
  XNOR2_X1 U3710 ( .A(n3960), .B(n4361), .ZN(n3959) );
  XOR2_X1 U3711 ( .A(REG1_REG_8__SCAN_IN), .B(n3959), .Z(n2878) );
  NAND2_X1 U3712 ( .A1(n2878), .A2(n4470), .ZN(n2884) );
  XNOR2_X1 U3713 ( .A(REG2_REG_8__SCAN_IN), .B(n3941), .ZN(n2880) );
  NAND2_X1 U3714 ( .A1(n4413), .A2(n2880), .ZN(n2881) );
  NAND2_X1 U3715 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3250) );
  NAND2_X1 U3716 ( .A1(n2881), .A2(n3250), .ZN(n2882) );
  AOI21_X1 U3717 ( .B1(n4468), .B2(ADDR_REG_8__SCAN_IN), .A(n2882), .ZN(n2883)
         );
  OAI211_X1 U3718 ( .C1(n4475), .C2(n4361), .A(n2884), .B(n2883), .ZN(U3248)
         );
  OAI22_X1 U3719 ( .A1(n2885), .A2(n3683), .B1(n3682), .B2(n2888), .ZN(n2886)
         );
  XNOR2_X1 U3720 ( .A(n2886), .B(n2043), .ZN(n2954) );
  INV_X2 U3721 ( .A(n2958), .ZN(n3679) );
  OAI22_X1 U3722 ( .A1(n2885), .A2(n2964), .B1(n3679), .B2(n2888), .ZN(n2953)
         );
  XNOR2_X1 U3723 ( .A(n2954), .B(n2953), .ZN(n2894) );
  NAND2_X1 U3724 ( .A1(n2892), .A2(n2891), .ZN(n2893) );
  NOR2_X1 U3725 ( .A1(n2893), .A2(n2894), .ZN(n2955) );
  AOI21_X1 U3726 ( .B1(n2894), .B2(n2893), .A(n2955), .ZN(n2899) );
  OAI22_X1 U3727 ( .A1(n2965), .A2(n3857), .B1(n3856), .B2(n2902), .ZN(n2897)
         );
  NOR2_X1 U3728 ( .A1(n2895), .A2(n2923), .ZN(n2896) );
  AOI211_X1 U3729 ( .C1(n2900), .C2(n3890), .A(n2897), .B(n2896), .ZN(n2898)
         );
  OAI21_X1 U3730 ( .B1(n2899), .B2(n3884), .A(n2898), .ZN(U3234) );
  AOI22_X1 U3731 ( .A1(n2959), .A2(n4283), .B1(n2900), .B2(n4295), .ZN(n2901)
         );
  OAI21_X1 U3732 ( .B1(n2902), .B2(n4299), .A(n2901), .ZN(n2904) );
  AOI211_X1 U3733 ( .C1(n4519), .C2(n2905), .A(n2904), .B(n2903), .ZN(n2938)
         );
  OAI22_X1 U3734 ( .A1(n4292), .A2(n2941), .B1(n4535), .B2(n2906), .ZN(n2907)
         );
  INV_X1 U3735 ( .A(n2907), .ZN(n2908) );
  OAI21_X1 U3736 ( .B1(n2938), .B2(n4533), .A(n2908), .ZN(U3520) );
  NAND2_X1 U3737 ( .A1(n2987), .A2(n2909), .ZN(n4511) );
  NAND2_X1 U3738 ( .A1(n2852), .A2(n2910), .ZN(n3498) );
  NAND2_X1 U3739 ( .A1(n3496), .A2(n3498), .ZN(n4515) );
  NAND2_X1 U3740 ( .A1(n4137), .A2(n4159), .ZN(n2911) );
  AOI22_X1 U3741 ( .A1(n4515), .A2(n2911), .B1(n4283), .B2(n3917), .ZN(n4512)
         );
  OAI21_X1 U3742 ( .B1(n2912), .B2(n4511), .A(n4512), .ZN(n2913) );
  AOI22_X1 U3743 ( .A1(n2913), .A2(n4187), .B1(REG3_REG_0__SCAN_IN), .B2(n4486), .ZN(n2915) );
  NAND2_X1 U3744 ( .A1(n4491), .A2(n4515), .ZN(n2914) );
  OAI211_X1 U3745 ( .C1(n4106), .C2(n2916), .A(n2915), .B(n2914), .ZN(U3290)
         );
  INV_X1 U3746 ( .A(IR_REG_0__SCAN_IN), .ZN(n3919) );
  OAI21_X1 U3747 ( .B1(REG2_REG_0__SCAN_IN), .B2(n3918), .A(n2917), .ZN(n3921)
         );
  NAND2_X1 U3748 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3931) );
  NOR2_X1 U3749 ( .A1(n2918), .A2(n2921), .ZN(n2919) );
  AOI211_X1 U3750 ( .C1(n2921), .C2(n3931), .A(n2920), .B(n2919), .ZN(n2922)
         );
  AOI211_X1 U3751 ( .C1(n3919), .C2(n3921), .A(n3903), .B(n2922), .ZN(n2949)
         );
  NOR2_X1 U3752 ( .A1(n2923), .A2(STATE_REG_SCAN_IN), .ZN(n2924) );
  AOI21_X1 U3753 ( .B1(n4468), .B2(ADDR_REG_2__SCAN_IN), .A(n2924), .ZN(n2925)
         );
  OAI21_X1 U3754 ( .B1(n4475), .B2(n2926), .A(n2925), .ZN(n2937) );
  OAI211_X1 U3755 ( .C1(n2929), .C2(n2928), .A(n4470), .B(n2927), .ZN(n2935)
         );
  MUX2_X1 U3756 ( .A(n2774), .B(REG2_REG_2__SCAN_IN), .S(n4366), .Z(n2931) );
  NAND3_X1 U3757 ( .A1(n2931), .A2(n3932), .A3(n2930), .ZN(n2932) );
  NAND3_X1 U3758 ( .A1(n4413), .A2(n2933), .A3(n2932), .ZN(n2934) );
  NAND2_X1 U3759 ( .A1(n2935), .A2(n2934), .ZN(n2936) );
  OR3_X1 U3760 ( .A1(n2949), .A2(n2937), .A3(n2936), .ZN(U3242) );
  OR2_X1 U3761 ( .A1(n2938), .A2(n4527), .ZN(n2940) );
  NAND2_X1 U3762 ( .A1(n4527), .A2(REG0_REG_2__SCAN_IN), .ZN(n2939) );
  OAI211_X1 U3763 ( .C1(n2941), .C2(n4355), .A(n2940), .B(n2939), .ZN(U3471)
         );
  XNOR2_X1 U3764 ( .A(n2942), .B(REG2_REG_4__SCAN_IN), .ZN(n2951) );
  OAI211_X1 U3765 ( .C1(REG1_REG_4__SCAN_IN), .C2(n2944), .A(n4470), .B(n2943), 
        .ZN(n2947) );
  NAND2_X1 U3766 ( .A1(REG3_REG_4__SCAN_IN), .A2(U3149), .ZN(n3046) );
  INV_X1 U3767 ( .A(n3046), .ZN(n2945) );
  AOI21_X1 U3768 ( .B1(n4468), .B2(ADDR_REG_4__SCAN_IN), .A(n2945), .ZN(n2946)
         );
  OAI211_X1 U3769 ( .C1(n4475), .C2(n2948), .A(n2947), .B(n2946), .ZN(n2950)
         );
  AOI211_X1 U3770 ( .C1(n4413), .C2(n2951), .A(n2950), .B(n2949), .ZN(n2952)
         );
  INV_X1 U3771 ( .A(n2952), .ZN(U3244) );
  INV_X1 U3772 ( .A(n2953), .ZN(n2957) );
  INV_X1 U3773 ( .A(n2954), .ZN(n2956) );
  AOI21_X1 U3774 ( .B1(n2957), .B2(n2956), .A(n2955), .ZN(n3043) );
  NAND2_X1 U3775 ( .A1(n2960), .A2(n3011), .ZN(n2961) );
  NAND2_X1 U3776 ( .A1(n2962), .A2(n2961), .ZN(n2963) );
  XNOR2_X1 U3777 ( .A(n2963), .B(n3675), .ZN(n3041) );
  OAI22_X1 U3778 ( .A1(n2965), .A2(n3680), .B1(n3679), .B2(n3016), .ZN(n3040)
         );
  XNOR2_X1 U3779 ( .A(n3041), .B(n3040), .ZN(n3042) );
  XNOR2_X1 U3780 ( .A(n3043), .B(n3042), .ZN(n2975) );
  OAI21_X1 U3781 ( .B1(n2967), .B2(n2966), .A(STATE_REG_SCAN_IN), .ZN(n2970)
         );
  AND2_X1 U3782 ( .A1(n2968), .A2(n3564), .ZN(n2969) );
  AOI21_X1 U3783 ( .B1(n3889), .B2(n3915), .A(n2971), .ZN(n2973) );
  AOI22_X1 U3784 ( .A1(n3891), .A2(n3916), .B1(n3890), .B2(n3011), .ZN(n2972)
         );
  OAI211_X1 U3785 ( .C1(n3895), .C2(REG3_REG_3__SCAN_IN), .A(n2973), .B(n2972), 
        .ZN(n2974) );
  AOI21_X1 U3786 ( .B1(n2975), .B2(n3897), .A(n2974), .ZN(n2976) );
  INV_X1 U3787 ( .A(n2976), .ZN(U3215) );
  OAI21_X1 U3788 ( .B1(n2977), .B2(n2979), .A(n2978), .ZN(n3030) );
  INV_X1 U3789 ( .A(n3030), .ZN(n2986) );
  AOI22_X1 U3790 ( .A1(n3916), .A2(n4283), .B1(n4295), .B2(n3034), .ZN(n2980)
         );
  OAI21_X1 U3791 ( .B1(n2981), .B2(n4299), .A(n2980), .ZN(n2985) );
  INV_X1 U3792 ( .A(n2982), .ZN(n2983) );
  AOI21_X1 U3793 ( .B1(n2977), .B2(n3496), .A(n2983), .ZN(n2984) );
  OAI22_X1 U3794 ( .A1(n2984), .A2(n4159), .B1(n4137), .B2(n3030), .ZN(n3031)
         );
  AOI211_X1 U3795 ( .C1(n4519), .C2(n2986), .A(n2985), .B(n3031), .ZN(n3028)
         );
  NAND2_X1 U3796 ( .A1(n3034), .A2(n2987), .ZN(n2988) );
  NAND2_X1 U3797 ( .A1(n2989), .A2(n2988), .ZN(n3037) );
  OAI22_X1 U3798 ( .A1(n4292), .A2(n3037), .B1(n4535), .B2(n2295), .ZN(n2990)
         );
  INV_X1 U3799 ( .A(n2990), .ZN(n2991) );
  OAI21_X1 U3800 ( .B1(n3028), .B2(n4533), .A(n2991), .ZN(U3519) );
  NAND2_X1 U3801 ( .A1(n2992), .A2(n2994), .ZN(n2993) );
  INV_X1 U3802 ( .A(n4520), .ZN(n3005) );
  INV_X1 U3803 ( .A(n2994), .ZN(n3473) );
  XNOR2_X1 U3804 ( .A(n2995), .B(n3473), .ZN(n3000) );
  AOI22_X1 U3805 ( .A1(n2959), .A2(n4261), .B1(n3048), .B2(n4295), .ZN(n2996)
         );
  OAI21_X1 U3806 ( .B1(n3125), .B2(n4293), .A(n2996), .ZN(n2997) );
  AOI21_X1 U3807 ( .B1(n4520), .B2(n2998), .A(n2997), .ZN(n2999) );
  OAI21_X1 U3808 ( .B1(n4159), .B2(n3000), .A(n2999), .ZN(n4517) );
  INV_X1 U3809 ( .A(n3018), .ZN(n3001) );
  OAI211_X1 U3810 ( .C1(n3001), .C2(n3039), .A(n4302), .B(n3062), .ZN(n4516)
         );
  OAI22_X1 U3811 ( .A1(n4516), .A2(n4360), .B1(n4476), .B2(n3051), .ZN(n3002)
         );
  OAI21_X1 U3812 ( .B1(n4517), .B2(n3002), .A(n4187), .ZN(n3004) );
  NAND2_X1 U3813 ( .A1(n4367), .A2(REG2_REG_4__SCAN_IN), .ZN(n3003) );
  OAI211_X1 U3814 ( .C1(n3005), .C2(n4147), .A(n3004), .B(n3003), .ZN(U3286)
         );
  NAND2_X1 U3815 ( .A1(n3007), .A2(n3006), .ZN(n3008) );
  XNOR2_X1 U3816 ( .A(n3008), .B(n3452), .ZN(n4487) );
  OAI21_X1 U3817 ( .B1(n3452), .B2(n3010), .A(n3009), .ZN(n3015) );
  AOI22_X1 U3818 ( .A1(n3916), .A2(n4261), .B1(n4295), .B2(n3011), .ZN(n3012)
         );
  OAI21_X1 U3819 ( .B1(n3132), .B2(n4293), .A(n3012), .ZN(n3014) );
  NOR2_X1 U3820 ( .A1(n4487), .A2(n4137), .ZN(n3013) );
  AOI211_X1 U3821 ( .C1(n4203), .C2(n3015), .A(n3014), .B(n3013), .ZN(n4495)
         );
  OAI21_X1 U3822 ( .B1(n4487), .B2(n3309), .A(n4495), .ZN(n3023) );
  OR2_X1 U3823 ( .A1(n3017), .A2(n3016), .ZN(n3019) );
  NAND2_X1 U3824 ( .A1(n3019), .A2(n3018), .ZN(n4488) );
  OAI22_X1 U3825 ( .A1(n4292), .A2(n4488), .B1(n4535), .B2(n3020), .ZN(n3021)
         );
  AOI21_X1 U3826 ( .B1(n3023), .B2(n4535), .A(n3021), .ZN(n3022) );
  INV_X1 U3827 ( .A(n3022), .ZN(U3521) );
  NAND2_X1 U3828 ( .A1(n3023), .A2(n4529), .ZN(n3025) );
  NAND2_X1 U3829 ( .A1(n4527), .A2(REG0_REG_3__SCAN_IN), .ZN(n3024) );
  OAI211_X1 U3830 ( .C1(n4488), .C2(n4355), .A(n3025), .B(n3024), .ZN(U3473)
         );
  OAI22_X1 U3831 ( .A1(n4355), .A2(n3037), .B1(n4529), .B2(n2294), .ZN(n3026)
         );
  INV_X1 U3832 ( .A(n3026), .ZN(n3027) );
  OAI21_X1 U3833 ( .B1(n3028), .B2(n4527), .A(n3027), .ZN(U3469) );
  INV_X1 U3834 ( .A(n4015), .ZN(n4197) );
  OAI22_X1 U3835 ( .A1(n4147), .A2(n3030), .B1(n3029), .B2(n4476), .ZN(n3033)
         );
  MUX2_X1 U3836 ( .A(REG2_REG_1__SCAN_IN), .B(n3031), .S(n4106), .Z(n3032) );
  AOI211_X1 U3837 ( .C1(n4197), .C2(n3034), .A(n3033), .B(n3032), .ZN(n3036)
         );
  AOI22_X1 U3838 ( .A1(n4196), .A2(n3916), .B1(n4012), .B2(n2852), .ZN(n3035)
         );
  OAI211_X1 U3839 ( .C1(n4164), .C2(n3037), .A(n3036), .B(n3035), .ZN(U3289)
         );
  OAI22_X1 U3840 ( .A1(n3132), .A2(n3679), .B1(n3682), .B2(n3039), .ZN(n3038)
         );
  XNOR2_X1 U3841 ( .A(n3038), .B(n2043), .ZN(n3122) );
  OAI22_X1 U3842 ( .A1(n3132), .A2(n3680), .B1(n3679), .B2(n3039), .ZN(n3123)
         );
  XNOR2_X1 U3843 ( .A(n3122), .B(n3123), .ZN(n3045) );
  OAI22_X1 U3844 ( .A1(n3043), .A2(n3042), .B1(n3041), .B2(n3040), .ZN(n3044)
         );
  AOI211_X1 U3845 ( .C1(n3045), .C2(n3044), .A(n3884), .B(n3121), .ZN(n3053)
         );
  OAI21_X1 U3846 ( .B1(n3857), .B2(n3125), .A(n3046), .ZN(n3047) );
  INV_X1 U3847 ( .A(n3047), .ZN(n3050) );
  AOI22_X1 U3848 ( .A1(n3891), .A2(n2959), .B1(n3890), .B2(n3048), .ZN(n3049)
         );
  OAI211_X1 U3849 ( .C1(n3895), .C2(n3051), .A(n3050), .B(n3049), .ZN(n3052)
         );
  OR2_X1 U3850 ( .A1(n3053), .A2(n3052), .ZN(U3227) );
  INV_X1 U3851 ( .A(n3054), .ZN(n3511) );
  NAND2_X1 U3852 ( .A1(n3511), .A2(n3487), .ZN(n3470) );
  NAND2_X1 U3853 ( .A1(n3056), .A2(n3055), .ZN(n3057) );
  XOR2_X1 U3854 ( .A(n3470), .B(n3057), .Z(n3118) );
  XNOR2_X1 U3855 ( .A(n3058), .B(n3470), .ZN(n3059) );
  NAND2_X1 U3856 ( .A1(n3059), .A2(n4203), .ZN(n3120) );
  AOI22_X1 U3857 ( .A1(n3913), .A2(n4283), .B1(n4295), .B2(n3126), .ZN(n3060)
         );
  OAI211_X1 U3858 ( .C1(n3132), .C2(n4299), .A(n3120), .B(n3060), .ZN(n3061)
         );
  AOI21_X1 U3859 ( .B1(n3118), .B2(n4521), .A(n3061), .ZN(n3097) );
  INV_X1 U3860 ( .A(n4355), .ZN(n3232) );
  AND2_X1 U3861 ( .A1(n3062), .A2(n3126), .ZN(n3063) );
  NOR2_X1 U3862 ( .A1(n3084), .A2(n3063), .ZN(n3111) );
  AOI22_X1 U3863 ( .A1(n3232), .A2(n3111), .B1(REG0_REG_5__SCAN_IN), .B2(n4527), .ZN(n3064) );
  OAI21_X1 U3864 ( .B1(n3097), .B2(n4527), .A(n3064), .ZN(U3477) );
  XNOR2_X1 U3865 ( .A(n3065), .B(n3515), .ZN(n3068) );
  AOI22_X1 U3866 ( .A1(n3911), .A2(n4283), .B1(n4295), .B2(n3193), .ZN(n3066)
         );
  OAI21_X1 U3867 ( .B1(n3144), .B2(n4299), .A(n3066), .ZN(n3067) );
  AOI21_X1 U3868 ( .B1(n3068), .B2(n4203), .A(n3067), .ZN(n4526) );
  AOI21_X1 U3869 ( .B1(n3086), .B2(n3193), .A(n3069), .ZN(n3070) );
  NAND2_X1 U3870 ( .A1(n3070), .A2(n3226), .ZN(n4525) );
  INV_X1 U3871 ( .A(n4525), .ZN(n3073) );
  INV_X1 U3872 ( .A(n4183), .ZN(n3072) );
  OAI22_X1 U3873 ( .A1(n4187), .A2(n2395), .B1(n3196), .B2(n4476), .ZN(n3071)
         );
  AOI21_X1 U3874 ( .B1(n3073), .B2(n3072), .A(n3071), .ZN(n3081) );
  OR2_X1 U3875 ( .A1(n3082), .A2(n3074), .ZN(n3076) );
  NAND2_X1 U3876 ( .A1(n3076), .A2(n3075), .ZN(n3077) );
  NAND2_X1 U3877 ( .A1(n3077), .A2(n3515), .ZN(n4522) );
  NAND2_X1 U3878 ( .A1(n4137), .A2(n3078), .ZN(n3079) );
  NAND2_X1 U3879 ( .A1(n4187), .A2(n3079), .ZN(n4210) );
  NAND3_X1 U3880 ( .A1(n4523), .A2(n4522), .A3(n4112), .ZN(n3080) );
  OAI211_X1 U3881 ( .C1(n4526), .C2(n4367), .A(n3081), .B(n3080), .ZN(U3283)
         );
  AND2_X1 U3882 ( .A1(n3514), .A2(n3510), .ZN(n3450) );
  XOR2_X1 U3883 ( .A(n3082), .B(n3450), .Z(n3102) );
  XNOR2_X1 U3884 ( .A(n3083), .B(n3450), .ZN(n3100) );
  NAND2_X1 U3885 ( .A1(n4187), .A2(n4203), .ZN(n3209) );
  INV_X1 U3886 ( .A(n3209), .ZN(n3093) );
  OR2_X1 U3887 ( .A1(n3084), .A2(n3143), .ZN(n3085) );
  NAND2_X1 U3888 ( .A1(n3086), .A2(n3085), .ZN(n3107) );
  OAI22_X1 U3889 ( .A1(n4106), .A2(n3087), .B1(n3150), .B2(n4476), .ZN(n3088)
         );
  AOI21_X1 U3890 ( .B1(n4012), .B2(n3914), .A(n3088), .ZN(n3091) );
  OAI22_X1 U3891 ( .A1(n3190), .A2(n3701), .B1(n4015), .B2(n3143), .ZN(n3089)
         );
  INV_X1 U3892 ( .A(n3089), .ZN(n3090) );
  OAI211_X1 U3893 ( .C1(n4164), .C2(n3107), .A(n3091), .B(n3090), .ZN(n3092)
         );
  AOI21_X1 U3894 ( .B1(n3100), .B2(n3093), .A(n3092), .ZN(n3094) );
  OAI21_X1 U3895 ( .B1(n3102), .B2(n4210), .A(n3094), .ZN(U3284) );
  NAND2_X1 U3896 ( .A1(n4533), .A2(REG1_REG_5__SCAN_IN), .ZN(n3096) );
  INV_X1 U3897 ( .A(n4292), .ZN(n3227) );
  NAND2_X1 U3898 ( .A1(n3227), .A2(n3111), .ZN(n3095) );
  OAI211_X1 U3899 ( .C1(n3097), .C2(n4533), .A(n3096), .B(n3095), .ZN(U3523)
         );
  AOI22_X1 U3900 ( .A1(n3912), .A2(n4283), .B1(n3147), .B2(n4295), .ZN(n3098)
         );
  OAI21_X1 U3901 ( .B1(n3125), .B2(n4299), .A(n3098), .ZN(n3099) );
  AOI21_X1 U3902 ( .B1(n3100), .B2(n4203), .A(n3099), .ZN(n3101) );
  OAI21_X1 U3903 ( .B1(n3102), .B2(n4306), .A(n3101), .ZN(n3109) );
  OAI22_X1 U3904 ( .A1(n4292), .A2(n3107), .B1(n4535), .B2(n3103), .ZN(n3104)
         );
  AOI21_X1 U3905 ( .B1(n3109), .B2(n4535), .A(n3104), .ZN(n3105) );
  INV_X1 U3906 ( .A(n3105), .ZN(U3524) );
  INV_X1 U3907 ( .A(REG0_REG_6__SCAN_IN), .ZN(n3106) );
  OAI22_X1 U3908 ( .A1(n4355), .A2(n3107), .B1(n4529), .B2(n3106), .ZN(n3108)
         );
  AOI21_X1 U3909 ( .B1(n3109), .B2(n4529), .A(n3108), .ZN(n3110) );
  INV_X1 U3910 ( .A(n3110), .ZN(U3479) );
  INV_X1 U3911 ( .A(n3111), .ZN(n3116) );
  INV_X1 U3912 ( .A(n3112), .ZN(n3138) );
  OAI22_X1 U3913 ( .A1(n4106), .A2(n2346), .B1(n3138), .B2(n4476), .ZN(n3114)
         );
  OAI22_X1 U3914 ( .A1(n3144), .A2(n3701), .B1(n4015), .B2(n3133), .ZN(n3113)
         );
  AOI211_X1 U3915 ( .C1(n4012), .C2(n3915), .A(n3114), .B(n3113), .ZN(n3115)
         );
  OAI21_X1 U3916 ( .B1(n4164), .B2(n3116), .A(n3115), .ZN(n3117) );
  AOI21_X1 U3917 ( .B1(n3118), .B2(n4112), .A(n3117), .ZN(n3119) );
  OAI21_X1 U3918 ( .B1(n4367), .B2(n3120), .A(n3119), .ZN(U3285) );
  AOI21_X1 U3919 ( .B1(n3123), .B2(n3122), .A(n3121), .ZN(n3130) );
  OAI22_X1 U3920 ( .A1(n3125), .A2(n3679), .B1(n3682), .B2(n3133), .ZN(n3124)
         );
  XNOR2_X1 U3921 ( .A(n3124), .B(n3675), .ZN(n3140) );
  OR2_X1 U3922 ( .A1(n3125), .A2(n3680), .ZN(n3128) );
  NAND2_X1 U3923 ( .A1(n3660), .A2(n3126), .ZN(n3127) );
  NAND2_X1 U3924 ( .A1(n3128), .A2(n3127), .ZN(n3139) );
  XNOR2_X1 U3925 ( .A(n3140), .B(n3139), .ZN(n3129) );
  NOR2_X1 U3926 ( .A1(n3130), .A2(n3129), .ZN(n3141) );
  AOI211_X1 U3927 ( .C1(n3130), .C2(n3129), .A(n3884), .B(n3141), .ZN(n3131)
         );
  INV_X1 U3928 ( .A(n3131), .ZN(n3137) );
  INV_X1 U3929 ( .A(n3890), .ZN(n3881) );
  OAI22_X1 U3930 ( .A1(n3881), .A2(n3133), .B1(n3132), .B2(n3856), .ZN(n3134)
         );
  AOI211_X1 U3931 ( .C1(n3889), .C2(n3913), .A(n3135), .B(n3134), .ZN(n3136)
         );
  OAI211_X1 U3932 ( .C1(n3895), .C2(n3138), .A(n3137), .B(n3136), .ZN(U3224)
         );
  OAI22_X1 U3933 ( .A1(n3144), .A2(n3679), .B1(n3682), .B2(n3143), .ZN(n3142)
         );
  XNOR2_X1 U3934 ( .A(n3142), .B(n3675), .ZN(n3187) );
  OAI22_X1 U3935 ( .A1(n3144), .A2(n3680), .B1(n3679), .B2(n3143), .ZN(n3186)
         );
  XNOR2_X1 U3936 ( .A(n3187), .B(n3188), .ZN(n3145) );
  XNOR2_X1 U3937 ( .A(n3189), .B(n3145), .ZN(n3152) );
  AOI21_X1 U3938 ( .B1(n3889), .B2(n3912), .A(n3146), .ZN(n3149) );
  AOI22_X1 U3939 ( .A1(n3891), .A2(n3914), .B1(n3890), .B2(n3147), .ZN(n3148)
         );
  OAI211_X1 U3940 ( .C1(n3895), .C2(n3150), .A(n3149), .B(n3148), .ZN(n3151)
         );
  AOI21_X1 U3941 ( .B1(n3152), .B2(n3897), .A(n3151), .ZN(n3153) );
  INV_X1 U3942 ( .A(n3153), .ZN(U3236) );
  AND2_X1 U3943 ( .A1(n2061), .A2(n3521), .ZN(n3453) );
  XOR2_X1 U3944 ( .A(n3154), .B(n3453), .Z(n3155) );
  NAND2_X1 U3945 ( .A1(n3155), .A2(n4203), .ZN(n3179) );
  INV_X1 U3946 ( .A(n3225), .ZN(n3156) );
  AOI21_X1 U3947 ( .B1(n3280), .B2(n3156), .A(n3169), .ZN(n3183) );
  AOI22_X1 U3948 ( .A1(n4196), .A2(n3909), .B1(n4012), .B2(n3911), .ZN(n3157)
         );
  OAI21_X1 U3949 ( .B1(n3275), .B2(n4015), .A(n3157), .ZN(n3159) );
  OAI22_X1 U3950 ( .A1(n3283), .A2(n4476), .B1(n2372), .B2(n4106), .ZN(n3158)
         );
  AOI211_X1 U3951 ( .C1(n3183), .C2(n4490), .A(n3159), .B(n3158), .ZN(n3166)
         );
  NAND2_X1 U3952 ( .A1(n4523), .A2(n3160), .ZN(n3219) );
  NAND2_X1 U3953 ( .A1(n3219), .A2(n3161), .ZN(n3163) );
  NAND2_X1 U3954 ( .A1(n3163), .A2(n3162), .ZN(n3164) );
  XNOR2_X1 U3955 ( .A(n3164), .B(n3453), .ZN(n3181) );
  NAND2_X1 U3956 ( .A1(n3181), .A2(n4112), .ZN(n3165) );
  OAI211_X1 U3957 ( .C1(n3179), .C2(n4367), .A(n3166), .B(n3165), .ZN(U3281)
         );
  NAND2_X1 U3958 ( .A1(n3490), .A2(n3486), .ZN(n3468) );
  XNOR2_X1 U3959 ( .A(n3167), .B(n3468), .ZN(n3212) );
  XNOR2_X1 U3960 ( .A(n3168), .B(n3468), .ZN(n3214) );
  NAND2_X1 U3961 ( .A1(n3214), .A2(n4112), .ZN(n3177) );
  INV_X1 U3962 ( .A(n3169), .ZN(n3171) );
  INV_X1 U3963 ( .A(n3170), .ZN(n3303) );
  AOI21_X1 U3964 ( .B1(n3747), .B2(n3171), .A(n3303), .ZN(n3216) );
  INV_X1 U3965 ( .A(n4012), .ZN(n4202) );
  AOI22_X1 U3966 ( .A1(n4197), .A2(n3747), .B1(n4196), .B2(n3908), .ZN(n3174)
         );
  INV_X1 U3967 ( .A(n3748), .ZN(n3172) );
  AOI22_X1 U3968 ( .A1(n4367), .A2(REG2_REG_10__SCAN_IN), .B1(n3172), .B2(
        n4486), .ZN(n3173) );
  OAI211_X1 U3969 ( .C1(n3276), .C2(n4202), .A(n3174), .B(n3173), .ZN(n3175)
         );
  AOI21_X1 U3970 ( .B1(n3216), .B2(n4490), .A(n3175), .ZN(n3176) );
  OAI211_X1 U3971 ( .C1(n3212), .C2(n3209), .A(n3177), .B(n3176), .ZN(U3280)
         );
  AOI22_X1 U3972 ( .A1(n3909), .A2(n4283), .B1(n4295), .B2(n3280), .ZN(n3178)
         );
  OAI211_X1 U3973 ( .C1(n3238), .C2(n4299), .A(n3179), .B(n3178), .ZN(n3180)
         );
  AOI21_X1 U3974 ( .B1(n3181), .B2(n4521), .A(n3180), .ZN(n3185) );
  AOI22_X1 U3975 ( .A1(n3183), .A2(n3227), .B1(REG1_REG_9__SCAN_IN), .B2(n4533), .ZN(n3182) );
  OAI21_X1 U3976 ( .B1(n3185), .B2(n4533), .A(n3182), .ZN(U3527) );
  AOI22_X1 U3977 ( .A1(n3183), .A2(n3232), .B1(REG0_REG_9__SCAN_IN), .B2(n4527), .ZN(n3184) );
  OAI21_X1 U3978 ( .B1(n3185), .B2(n4527), .A(n3184), .ZN(U3485) );
  INV_X1 U3979 ( .A(n3186), .ZN(n3188) );
  OAI22_X1 U3980 ( .A1(n3190), .A2(n3680), .B1(n3679), .B2(n2074), .ZN(n3246)
         );
  OAI22_X1 U3981 ( .A1(n3190), .A2(n3683), .B1(n3682), .B2(n2074), .ZN(n3191)
         );
  XNOR2_X1 U3982 ( .A(n3191), .B(n3675), .ZN(n3245) );
  XOR2_X1 U3983 ( .A(n3246), .B(n3245), .Z(n3247) );
  XOR2_X1 U3984 ( .A(n3248), .B(n3247), .Z(n3198) );
  AOI21_X1 U3985 ( .B1(n3889), .B2(n3911), .A(n3192), .ZN(n3195) );
  AOI22_X1 U3986 ( .A1(n3891), .A2(n3913), .B1(n3890), .B2(n3193), .ZN(n3194)
         );
  OAI211_X1 U3987 ( .C1(n3895), .C2(n3196), .A(n3195), .B(n3194), .ZN(n3197)
         );
  AOI21_X1 U3988 ( .B1(n3198), .B2(n3897), .A(n3197), .ZN(n3199) );
  INV_X1 U3989 ( .A(n3199), .ZN(U3210) );
  XNOR2_X1 U3990 ( .A(n3428), .B(n3472), .ZN(n3335) );
  OAI21_X1 U3991 ( .B1(n3201), .B2(n3472), .A(n3200), .ZN(n3337) );
  NAND2_X1 U3992 ( .A1(n3337), .A2(n4112), .ZN(n3208) );
  OAI21_X1 U3993 ( .B1(n3327), .B2(n3591), .A(n3262), .ZN(n3343) );
  INV_X1 U3994 ( .A(n3343), .ZN(n3206) );
  AOI22_X1 U3995 ( .A1(n4197), .A2(n3726), .B1(n4196), .B2(n2487), .ZN(n3204)
         );
  INV_X1 U3996 ( .A(n3729), .ZN(n3202) );
  AOI22_X1 U3997 ( .A1(n4367), .A2(REG2_REG_14__SCAN_IN), .B1(n3202), .B2(
        n4486), .ZN(n3203) );
  OAI211_X1 U3998 ( .C1(n3780), .C2(n4202), .A(n3204), .B(n3203), .ZN(n3205)
         );
  AOI21_X1 U3999 ( .B1(n3206), .B2(n4490), .A(n3205), .ZN(n3207) );
  OAI211_X1 U4000 ( .C1(n3335), .C2(n3209), .A(n3208), .B(n3207), .ZN(U3276)
         );
  OAI22_X1 U4001 ( .A1(n3745), .A2(n4293), .B1(n4220), .B2(n3365), .ZN(n3210)
         );
  AOI21_X1 U4002 ( .B1(n4261), .B2(n3910), .A(n3210), .ZN(n3211) );
  OAI21_X1 U4003 ( .B1(n3212), .B2(n4159), .A(n3211), .ZN(n3213) );
  AOI21_X1 U4004 ( .B1(n4521), .B2(n3214), .A(n3213), .ZN(n3218) );
  AOI22_X1 U4005 ( .A1(n3216), .A2(n3232), .B1(REG0_REG_10__SCAN_IN), .B2(
        n4527), .ZN(n3215) );
  OAI21_X1 U4006 ( .B1(n3218), .B2(n4527), .A(n3215), .ZN(U3487) );
  AOI22_X1 U4007 ( .A1(n3216), .A2(n3227), .B1(REG1_REG_10__SCAN_IN), .B2(
        n4533), .ZN(n3217) );
  OAI21_X1 U4008 ( .B1(n3218), .B2(n4533), .A(n3217), .ZN(U3528) );
  INV_X1 U4009 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3230) );
  AND2_X1 U4010 ( .A1(n3520), .A2(n3517), .ZN(n3451) );
  XOR2_X1 U4011 ( .A(n3451), .B(n3219), .Z(n4480) );
  XOR2_X1 U4012 ( .A(n3451), .B(n3220), .Z(n3224) );
  AOI22_X1 U4013 ( .A1(n3912), .A2(n4261), .B1(n3252), .B2(n4295), .ZN(n3221)
         );
  OAI21_X1 U4014 ( .B1(n3276), .B2(n4293), .A(n3221), .ZN(n3223) );
  NOR2_X1 U4015 ( .A1(n4480), .A2(n4137), .ZN(n3222) );
  AOI211_X1 U4016 ( .C1(n4203), .C2(n3224), .A(n3223), .B(n3222), .ZN(n4485)
         );
  OAI21_X1 U4017 ( .B1(n3309), .B2(n4480), .A(n4485), .ZN(n3231) );
  NAND2_X1 U4018 ( .A1(n3231), .A2(n4535), .ZN(n3229) );
  AOI21_X1 U4019 ( .B1(n3252), .B2(n3226), .A(n3225), .ZN(n4481) );
  NAND2_X1 U4020 ( .A1(n4481), .A2(n3227), .ZN(n3228) );
  OAI211_X1 U4021 ( .C1(n4535), .C2(n3230), .A(n3229), .B(n3228), .ZN(U3526)
         );
  INV_X1 U4022 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3235) );
  NAND2_X1 U4023 ( .A1(n3231), .A2(n4529), .ZN(n3234) );
  NAND2_X1 U4024 ( .A1(n4481), .A2(n3232), .ZN(n3233) );
  OAI211_X1 U4025 ( .C1(n4529), .C2(n3235), .A(n3234), .B(n3233), .ZN(U3483)
         );
  OAI22_X1 U4026 ( .A1(n3238), .A2(n3683), .B1(n3682), .B2(n3236), .ZN(n3237)
         );
  XNOR2_X1 U4027 ( .A(n3237), .B(n2043), .ZN(n3241) );
  OR2_X1 U4028 ( .A1(n3238), .A2(n3680), .ZN(n3240) );
  NAND2_X1 U4029 ( .A1(n3660), .A2(n3252), .ZN(n3239) );
  NAND2_X1 U4030 ( .A1(n3240), .A2(n3239), .ZN(n3242) );
  NAND2_X1 U4031 ( .A1(n3241), .A2(n3242), .ZN(n3271) );
  INV_X1 U4032 ( .A(n3241), .ZN(n3244) );
  INV_X1 U4033 ( .A(n3242), .ZN(n3243) );
  NAND2_X1 U4034 ( .A1(n3244), .A2(n3243), .ZN(n3273) );
  NAND2_X1 U4035 ( .A1(n3271), .A2(n3273), .ZN(n3249) );
  AOI21_X1 U4036 ( .B1(n3248), .B2(n3247), .A(n2049), .ZN(n3272) );
  XOR2_X1 U4037 ( .A(n3249), .B(n3272), .Z(n3256) );
  OAI21_X1 U4038 ( .B1(n3857), .B2(n3276), .A(n3250), .ZN(n3251) );
  INV_X1 U4039 ( .A(n3251), .ZN(n3254) );
  AOI22_X1 U4040 ( .A1(n3891), .A2(n3912), .B1(n3890), .B2(n3252), .ZN(n3253)
         );
  OAI211_X1 U4041 ( .C1(n3895), .C2(n4477), .A(n3254), .B(n3253), .ZN(n3255)
         );
  AOI21_X1 U4042 ( .B1(n3256), .B2(n3897), .A(n3255), .ZN(n3257) );
  INV_X1 U40430 ( .A(n3257), .ZN(U3218) );
  AOI21_X1 U4044 ( .B1(n3258), .B2(n3454), .A(n4159), .ZN(n3260) );
  NAND2_X1 U4045 ( .A1(n3260), .A2(n3259), .ZN(n3389) );
  XNOR2_X1 U4046 ( .A(n3261), .B(n3454), .ZN(n3391) );
  NAND2_X1 U4047 ( .A1(n3391), .A2(n4112), .ZN(n3270) );
  INV_X1 U4048 ( .A(n3262), .ZN(n3263) );
  OAI21_X1 U4049 ( .B1(n3263), .B2(n3596), .A(n2051), .ZN(n3397) );
  INV_X1 U4050 ( .A(n3397), .ZN(n3268) );
  AOI22_X1 U4051 ( .A1(n2486), .A2(n4197), .B1(n4196), .B2(n3904), .ZN(n3266)
         );
  INV_X1 U4052 ( .A(n3894), .ZN(n3264) );
  AOI22_X1 U4053 ( .A1(n4367), .A2(REG2_REG_15__SCAN_IN), .B1(n3264), .B2(
        n4486), .ZN(n3265) );
  OAI211_X1 U4054 ( .C1(n3593), .C2(n4202), .A(n3266), .B(n3265), .ZN(n3267)
         );
  AOI21_X1 U4055 ( .B1(n3268), .B2(n4490), .A(n3267), .ZN(n3269) );
  OAI211_X1 U4056 ( .C1(n4367), .C2(n3389), .A(n3270), .B(n3269), .ZN(U3275)
         );
  NAND2_X1 U4057 ( .A1(n3272), .A2(n3271), .ZN(n3274) );
  NAND2_X1 U4058 ( .A1(n3274), .A2(n3273), .ZN(n3361) );
  OAI22_X1 U4059 ( .A1(n3276), .A2(n3680), .B1(n3679), .B2(n3275), .ZN(n3357)
         );
  NAND2_X1 U4060 ( .A1(n3910), .A2(n3660), .ZN(n3278) );
  NAND2_X1 U4061 ( .A1(n2960), .A2(n3280), .ZN(n3277) );
  NAND2_X1 U4062 ( .A1(n3278), .A2(n3277), .ZN(n3279) );
  XNOR2_X1 U4063 ( .A(n3279), .B(n2043), .ZN(n3358) );
  XOR2_X1 U4064 ( .A(n3357), .B(n3358), .Z(n3360) );
  XNOR2_X1 U4065 ( .A(n3361), .B(n3360), .ZN(n3285) );
  AND2_X1 U4066 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n4380) );
  AOI21_X1 U4067 ( .B1(n3889), .B2(n3909), .A(n4380), .ZN(n3282) );
  AOI22_X1 U4068 ( .A1(n3891), .A2(n3911), .B1(n3890), .B2(n3280), .ZN(n3281)
         );
  OAI211_X1 U4069 ( .C1(n3895), .C2(n3283), .A(n3282), .B(n3281), .ZN(n3284)
         );
  AOI21_X1 U4070 ( .B1(n3285), .B2(n3897), .A(n3284), .ZN(n3286) );
  INV_X1 U4071 ( .A(n3286), .ZN(U3228) );
  NAND2_X1 U4072 ( .A1(n3318), .A2(n3316), .ZN(n3469) );
  XNOR2_X1 U4073 ( .A(n3287), .B(n3469), .ZN(n3344) );
  AND2_X1 U4074 ( .A1(n3302), .A2(n3782), .ZN(n3288) );
  OR2_X1 U4075 ( .A1(n3288), .A2(n3325), .ZN(n3356) );
  OAI22_X1 U4076 ( .A1(n4106), .A2(n3289), .B1(n3785), .B2(n4476), .ZN(n3290)
         );
  AOI21_X1 U4077 ( .B1(n4012), .B2(n3908), .A(n3290), .ZN(n3293) );
  OAI22_X1 U4078 ( .A1(n3780), .A2(n3701), .B1(n4015), .B2(n3578), .ZN(n3291)
         );
  INV_X1 U4079 ( .A(n3291), .ZN(n3292) );
  OAI211_X1 U4080 ( .C1(n3356), .C2(n4164), .A(n3293), .B(n3292), .ZN(n3300)
         );
  INV_X1 U4081 ( .A(n3295), .ZN(n3296) );
  AOI21_X1 U4082 ( .B1(n3294), .B2(n3297), .A(n3296), .ZN(n3319) );
  XNOR2_X1 U4083 ( .A(n3319), .B(n3469), .ZN(n3298) );
  NAND2_X1 U4084 ( .A1(n3298), .A2(n4203), .ZN(n3348) );
  NOR2_X1 U4085 ( .A1(n3348), .A2(n4367), .ZN(n3299) );
  AOI211_X1 U4086 ( .C1(n4112), .C2(n3344), .A(n3300), .B(n3299), .ZN(n3301)
         );
  INV_X1 U4087 ( .A(n3301), .ZN(U3278) );
  OAI21_X1 U4088 ( .B1(n3303), .B2(n3372), .A(n3302), .ZN(n3569) );
  INV_X1 U4089 ( .A(REG0_REG_11__SCAN_IN), .ZN(n3311) );
  AOI21_X1 U4090 ( .B1(n3455), .B2(n3304), .A(n2067), .ZN(n3574) );
  AOI22_X1 U4091 ( .A1(n3907), .A2(n4283), .B1(n4295), .B2(n3374), .ZN(n3307)
         );
  XNOR2_X1 U4092 ( .A(n3294), .B(n3455), .ZN(n3305) );
  NAND2_X1 U4093 ( .A1(n3305), .A2(n4203), .ZN(n3306) );
  OAI211_X1 U4094 ( .C1(n3574), .C2(n4137), .A(n3307), .B(n3306), .ZN(n3566)
         );
  OAI22_X1 U4095 ( .A1(n3574), .A2(n3309), .B1(n3308), .B2(n4299), .ZN(n3310)
         );
  NOR2_X1 U4096 ( .A1(n3566), .A2(n3310), .ZN(n3313) );
  MUX2_X1 U4097 ( .A(n3311), .B(n3313), .S(n4529), .Z(n3312) );
  OAI21_X1 U4098 ( .B1(n3569), .B2(n4355), .A(n3312), .ZN(U3489) );
  MUX2_X1 U4099 ( .A(n3314), .B(n3313), .S(n4535), .Z(n3315) );
  OAI21_X1 U4100 ( .B1(n4292), .B2(n3569), .A(n3315), .ZN(U3529) );
  XNOR2_X1 U4101 ( .A(n3780), .B(n3588), .ZN(n3479) );
  INV_X1 U4102 ( .A(n3316), .ZN(n3317) );
  AOI21_X1 U4103 ( .B1(n3319), .B2(n3318), .A(n3317), .ZN(n3320) );
  XOR2_X1 U4104 ( .A(n3479), .B(n3320), .Z(n3323) );
  OAI22_X1 U4105 ( .A1(n3593), .A2(n4293), .B1(n4220), .B2(n3588), .ZN(n3321)
         );
  AOI21_X1 U4106 ( .B1(n4261), .B2(n3907), .A(n3321), .ZN(n3322) );
  OAI21_X1 U4107 ( .B1(n3323), .B2(n4159), .A(n3322), .ZN(n3380) );
  INV_X1 U4108 ( .A(n3380), .ZN(n3332) );
  XOR2_X1 U4109 ( .A(n3479), .B(n3324), .Z(n3381) );
  NOR2_X1 U4110 ( .A1(n3325), .A2(n3588), .ZN(n3326) );
  OR2_X1 U4111 ( .A1(n3327), .A2(n3326), .ZN(n3387) );
  INV_X1 U4112 ( .A(n3847), .ZN(n3328) );
  AOI22_X1 U4113 ( .A1(n4367), .A2(REG2_REG_13__SCAN_IN), .B1(n3328), .B2(
        n4486), .ZN(n3329) );
  OAI21_X1 U4114 ( .B1(n3387), .B2(n4164), .A(n3329), .ZN(n3330) );
  AOI21_X1 U4115 ( .B1(n3381), .B2(n4112), .A(n3330), .ZN(n3331) );
  OAI21_X1 U4116 ( .B1(n4367), .B2(n3332), .A(n3331), .ZN(U3277) );
  OAI22_X1 U4117 ( .A1(n4300), .A2(n4293), .B1(n4220), .B2(n3591), .ZN(n3333)
         );
  AOI21_X1 U4118 ( .B1(n4261), .B2(n3906), .A(n3333), .ZN(n3334) );
  OAI21_X1 U4119 ( .B1(n3335), .B2(n4159), .A(n3334), .ZN(n3336) );
  AOI21_X1 U4120 ( .B1(n3337), .B2(n4521), .A(n3336), .ZN(n3340) );
  MUX2_X1 U4121 ( .A(n3338), .B(n3340), .S(n4535), .Z(n3339) );
  OAI21_X1 U4122 ( .B1(n4292), .B2(n3343), .A(n3339), .ZN(U3532) );
  INV_X1 U4123 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3341) );
  MUX2_X1 U4124 ( .A(n3341), .B(n3340), .S(n4529), .Z(n3342) );
  OAI21_X1 U4125 ( .B1(n3343), .B2(n4355), .A(n3342), .ZN(U3495) );
  NAND2_X1 U4126 ( .A1(n3344), .A2(n4521), .ZN(n3350) );
  OR2_X1 U4127 ( .A1(n3745), .A2(n4299), .ZN(n3346) );
  NAND2_X1 U4128 ( .A1(n3782), .A2(n4295), .ZN(n3345) );
  OAI211_X1 U4129 ( .C1(n3780), .C2(n4293), .A(n3346), .B(n3345), .ZN(n3347)
         );
  INV_X1 U4130 ( .A(n3347), .ZN(n3349) );
  MUX2_X1 U4131 ( .A(n3351), .B(n3353), .S(n4535), .Z(n3352) );
  OAI21_X1 U4132 ( .B1(n4292), .B2(n3356), .A(n3352), .ZN(U3530) );
  INV_X1 U4133 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3354) );
  MUX2_X1 U4134 ( .A(n3354), .B(n3353), .S(n4529), .Z(n3355) );
  OAI21_X1 U4135 ( .B1(n3356), .B2(n4355), .A(n3355), .ZN(U3491) );
  NOR2_X1 U4136 ( .A1(n3358), .A2(n3357), .ZN(n3359) );
  AOI21_X2 U4137 ( .B1(n3361), .B2(n3360), .A(n3359), .ZN(n3744) );
  NAND2_X1 U4138 ( .A1(n3909), .A2(n3660), .ZN(n3363) );
  NAND2_X1 U4139 ( .A1(n2960), .A2(n3747), .ZN(n3362) );
  NAND2_X1 U4140 ( .A1(n3363), .A2(n3362), .ZN(n3364) );
  XNOR2_X1 U4141 ( .A(n3364), .B(n2043), .ZN(n3369) );
  NOR2_X1 U4142 ( .A1(n3679), .A2(n3365), .ZN(n3366) );
  AOI21_X1 U4143 ( .B1(n3669), .B2(n3909), .A(n3366), .ZN(n3367) );
  XNOR2_X1 U4144 ( .A(n3369), .B(n3367), .ZN(n3743) );
  INV_X1 U4145 ( .A(n3367), .ZN(n3368) );
  NAND2_X1 U4146 ( .A1(n3369), .A2(n3368), .ZN(n3370) );
  OAI22_X1 U4147 ( .A1(n3745), .A2(n3683), .B1(n3682), .B2(n3372), .ZN(n3371)
         );
  XNOR2_X1 U4148 ( .A(n3371), .B(n2043), .ZN(n3575) );
  OAI22_X1 U4149 ( .A1(n3745), .A2(n3680), .B1(n3679), .B2(n3372), .ZN(n3576)
         );
  XNOR2_X1 U4150 ( .A(n3575), .B(n3576), .ZN(n3373) );
  XNOR2_X1 U4151 ( .A(n3577), .B(n3373), .ZN(n3378) );
  AND2_X1 U4152 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4400) );
  AOI21_X1 U4153 ( .B1(n3889), .B2(n3907), .A(n4400), .ZN(n3376) );
  AOI22_X1 U4154 ( .A1(n3891), .A2(n3909), .B1(n3890), .B2(n3374), .ZN(n3375)
         );
  OAI211_X1 U4155 ( .C1(n3895), .C2(n3567), .A(n3376), .B(n3375), .ZN(n3377)
         );
  AOI21_X1 U4156 ( .B1(n3378), .B2(n3897), .A(n3377), .ZN(n3379) );
  INV_X1 U4157 ( .A(n3379), .ZN(U3233) );
  AOI21_X1 U4158 ( .B1(n4521), .B2(n3381), .A(n3380), .ZN(n3384) );
  MUX2_X1 U4159 ( .A(n3382), .B(n3384), .S(n4535), .Z(n3383) );
  OAI21_X1 U4160 ( .B1(n4292), .B2(n3387), .A(n3383), .ZN(U3531) );
  INV_X1 U4161 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3385) );
  MUX2_X1 U4162 ( .A(n3385), .B(n3384), .S(n4529), .Z(n3386) );
  OAI21_X1 U4163 ( .B1(n3387), .B2(n4355), .A(n3386), .ZN(U3493) );
  AOI22_X1 U4164 ( .A1(n3904), .A2(n4283), .B1(n2486), .B2(n4295), .ZN(n3388)
         );
  OAI211_X1 U4165 ( .C1(n3593), .C2(n4299), .A(n3389), .B(n3388), .ZN(n3390)
         );
  AOI21_X1 U4166 ( .B1(n3391), .B2(n4521), .A(n3390), .ZN(n3394) );
  MUX2_X1 U4167 ( .A(n3392), .B(n3394), .S(n4535), .Z(n3393) );
  OAI21_X1 U4168 ( .B1(n4292), .B2(n3397), .A(n3393), .ZN(U3533) );
  INV_X1 U4169 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3395) );
  MUX2_X1 U4170 ( .A(n3395), .B(n3394), .S(n4529), .Z(n3396) );
  OAI21_X1 U4171 ( .B1(n3397), .B2(n4355), .A(n3396), .ZN(U3497) );
  NAND2_X1 U4172 ( .A1(n2251), .A2(n4149), .ZN(n3466) );
  XNOR2_X1 U4173 ( .A(n3398), .B(n3466), .ZN(n3399) );
  NAND2_X1 U4174 ( .A1(n3399), .A2(n4203), .ZN(n4286) );
  XNOR2_X1 U4175 ( .A(n3400), .B(n3466), .ZN(n4289) );
  NAND2_X1 U4176 ( .A1(n4289), .A2(n4112), .ZN(n3408) );
  INV_X1 U4177 ( .A(n4194), .ZN(n3402) );
  INV_X1 U4178 ( .A(n4182), .ZN(n3401) );
  OAI21_X1 U4179 ( .B1(n3402), .B2(n3616), .A(n3401), .ZN(n4356) );
  INV_X1 U4180 ( .A(n4356), .ZN(n3406) );
  AOI22_X1 U4181 ( .A1(n4197), .A2(n4282), .B1(n4196), .B2(n4284), .ZN(n3404)
         );
  AOI22_X1 U4182 ( .A1(n4367), .A2(REG2_REG_17__SCAN_IN), .B1(n3812), .B2(
        n4486), .ZN(n3403) );
  OAI211_X1 U4183 ( .C1(n4287), .C2(n4202), .A(n3404), .B(n3403), .ZN(n3405)
         );
  AOI21_X1 U4184 ( .B1(n3406), .B2(n4490), .A(n3405), .ZN(n3407) );
  OAI211_X1 U4185 ( .C1(n4367), .C2(n4286), .A(n3408), .B(n3407), .ZN(U3273)
         );
  INV_X1 U4186 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4211) );
  NAND2_X1 U4187 ( .A1(n3409), .A2(REG2_REG_31__SCAN_IN), .ZN(n3412) );
  NAND2_X1 U4188 ( .A1(n3410), .A2(REG0_REG_31__SCAN_IN), .ZN(n3411) );
  OAI211_X1 U4189 ( .C1(n2311), .C2(n4211), .A(n3412), .B(n3411), .ZN(n3988)
         );
  INV_X1 U4190 ( .A(DATAI_30_), .ZN(n4696) );
  NOR2_X1 U4191 ( .A1(n2319), .A2(n4696), .ZN(n4218) );
  INV_X1 U4192 ( .A(n4218), .ZN(n3458) );
  OAI21_X1 U4193 ( .B1(n3702), .B2(n3414), .A(n3413), .ZN(n3542) );
  NOR3_X1 U4194 ( .A1(n3542), .A2(n4005), .A3(n3415), .ZN(n3441) );
  NAND2_X1 U4195 ( .A1(n3417), .A2(n3416), .ZN(n3437) );
  INV_X1 U4196 ( .A(n3437), .ZN(n3420) );
  NAND2_X1 U4197 ( .A1(n2333), .A2(DATAI_31_), .ZN(n3989) );
  NAND2_X1 U4198 ( .A1(n3988), .A2(n3989), .ZN(n3550) );
  OR2_X1 U4199 ( .A1(n3900), .A2(n3458), .ZN(n3418) );
  OAI211_X1 U4200 ( .C1(n3901), .C2(n3994), .A(n3550), .B(n3418), .ZN(n3436)
         );
  INV_X1 U4201 ( .A(n3436), .ZN(n3419) );
  OAI21_X1 U4202 ( .B1(n3420), .B2(n3542), .A(n3419), .ZN(n3546) );
  NAND2_X1 U4203 ( .A1(n3421), .A2(n3427), .ZN(n3530) );
  NAND2_X1 U4204 ( .A1(n3491), .A2(n3492), .ZN(n3426) );
  INV_X1 U4205 ( .A(n3493), .ZN(n3425) );
  INV_X1 U4206 ( .A(n3422), .ZN(n3424) );
  NAND3_X1 U4207 ( .A1(n3424), .A2(n3423), .A3(n2251), .ZN(n3495) );
  AOI211_X1 U4208 ( .C1(n3427), .C2(n3426), .A(n3425), .B(n3495), .ZN(n3529)
         );
  OAI21_X1 U4209 ( .B1(n3428), .B2(n3530), .A(n3529), .ZN(n3432) );
  INV_X1 U4210 ( .A(n3495), .ZN(n3431) );
  INV_X1 U4211 ( .A(n3429), .ZN(n3430) );
  NAND2_X1 U4212 ( .A1(n3431), .A2(n3430), .ZN(n3534) );
  NAND4_X1 U4213 ( .A1(n3432), .A2(n3536), .A3(n3535), .A4(n3534), .ZN(n3435)
         );
  INV_X1 U4214 ( .A(n3447), .ZN(n3433) );
  NAND2_X1 U4215 ( .A1(n3433), .A2(n3449), .ZN(n3539) );
  AOI21_X1 U4216 ( .B1(n3435), .B2(n3434), .A(n3539), .ZN(n3439) );
  NOR3_X1 U4217 ( .A1(n3437), .A2(n3538), .A3(n3436), .ZN(n3438) );
  OAI21_X1 U4218 ( .B1(n3439), .B2(n4023), .A(n3438), .ZN(n3440) );
  OAI21_X1 U4219 ( .B1(n3441), .B2(n3546), .A(n3440), .ZN(n3442) );
  OAI21_X1 U4220 ( .B1(n3988), .B2(n3458), .A(n3442), .ZN(n3557) );
  NAND2_X1 U4221 ( .A1(n3900), .A2(n3458), .ZN(n3547) );
  AOI21_X1 U4222 ( .B1(n3547), .B2(n3988), .A(n3989), .ZN(n3444) );
  NOR2_X1 U4223 ( .A1(n3444), .A2(n3443), .ZN(n3556) );
  NAND2_X1 U4224 ( .A1(n4022), .A2(n3445), .ZN(n4042) );
  INV_X1 U4225 ( .A(n4038), .ZN(n3446) );
  OR2_X1 U4226 ( .A1(n3447), .A2(n3446), .ZN(n4060) );
  NAND2_X1 U4227 ( .A1(n3449), .A2(n3448), .ZN(n4077) );
  NAND4_X1 U4228 ( .A1(n3453), .A2(n3452), .A3(n3451), .A4(n3450), .ZN(n3457)
         );
  NAND4_X1 U4229 ( .A1(n2637), .A2(n4205), .A3(n3455), .A4(n3515), .ZN(n3456)
         );
  NOR4_X1 U4230 ( .A1(n4077), .A2(n4100), .A3(n3457), .A4(n3456), .ZN(n3480)
         );
  XNOR2_X1 U4231 ( .A(n3900), .B(n3458), .ZN(n3461) );
  OR2_X1 U4232 ( .A1(n3988), .A2(n3989), .ZN(n3548) );
  NAND3_X1 U4233 ( .A1(n3548), .A2(n3550), .A3(n3459), .ZN(n3460) );
  NOR3_X1 U4234 ( .A1(n4515), .A2(n3461), .A3(n3460), .ZN(n3478) );
  INV_X1 U4235 ( .A(n3462), .ZN(n4074) );
  NOR2_X1 U4236 ( .A1(n4073), .A2(n4074), .ZN(n4111) );
  NAND2_X1 U4237 ( .A1(n2064), .A2(n3463), .ZN(n4129) );
  INV_X1 U4238 ( .A(n4129), .ZN(n3467) );
  NAND2_X1 U4239 ( .A1(n3465), .A2(n3464), .ZN(n4155) );
  NOR3_X1 U4240 ( .A1(n3467), .A2(n4155), .A3(n3466), .ZN(n3476) );
  NOR4_X1 U4241 ( .A1(n4174), .A2(n3470), .A3(n3469), .A4(n3468), .ZN(n3475)
         );
  NOR4_X1 U4242 ( .A1(n3473), .A2(n2320), .A3(n3472), .A4(n2977), .ZN(n3474)
         );
  AND4_X1 U4243 ( .A1(n4111), .A2(n3476), .A3(n3475), .A4(n3474), .ZN(n3477)
         );
  NAND4_X1 U4244 ( .A1(n3480), .A2(n3479), .A3(n3478), .A4(n3477), .ZN(n3481)
         );
  OR4_X1 U4245 ( .A1(n3482), .A2(n4042), .A3(n4060), .A4(n3481), .ZN(n3484) );
  XNOR2_X1 U4246 ( .A(n4237), .B(n4032), .ZN(n4019) );
  INV_X1 U4247 ( .A(n4019), .ZN(n4025) );
  NOR4_X1 U4248 ( .A1(n3484), .A2(n3483), .A3(n4005), .A4(n4025), .ZN(n3554)
         );
  INV_X1 U4249 ( .A(n3485), .ZN(n3541) );
  NOR2_X1 U4250 ( .A1(n2119), .A2(n3487), .ZN(n3488) );
  NAND4_X1 U4251 ( .A1(n3488), .A2(n2061), .A3(n3517), .A4(n3510), .ZN(n3489)
         );
  NAND2_X1 U4252 ( .A1(n3490), .A2(n3489), .ZN(n3524) );
  NAND4_X1 U4253 ( .A1(n2061), .A2(n3493), .A3(n3492), .A4(n3491), .ZN(n3494)
         );
  NOR2_X1 U4254 ( .A1(n3495), .A2(n3494), .ZN(n3523) );
  INV_X1 U4255 ( .A(n3496), .ZN(n3499) );
  OAI211_X1 U4256 ( .C1(n4359), .C2(n3499), .A(n3498), .B(n3497), .ZN(n3500)
         );
  NAND3_X1 U4257 ( .A1(n3502), .A2(n3501), .A3(n3500), .ZN(n3503) );
  NAND3_X1 U4258 ( .A1(n3505), .A2(n3504), .A3(n3503), .ZN(n3506) );
  NAND3_X1 U4259 ( .A1(n3508), .A2(n3507), .A3(n3506), .ZN(n3509) );
  NAND4_X1 U4260 ( .A1(n3512), .A2(n3511), .A3(n3510), .A4(n3509), .ZN(n3513)
         );
  NAND3_X1 U4261 ( .A1(n3515), .A2(n3514), .A3(n3513), .ZN(n3516) );
  NAND3_X1 U4262 ( .A1(n3518), .A2(n3517), .A3(n3516), .ZN(n3519) );
  NAND3_X1 U4263 ( .A1(n3521), .A2(n3520), .A3(n3519), .ZN(n3522) );
  AOI22_X1 U4264 ( .A1(n3529), .A2(n3524), .B1(n3523), .B2(n3522), .ZN(n3526)
         );
  OR4_X1 U4265 ( .A1(n3527), .A2(n2114), .A3(n3526), .A4(n3525), .ZN(n3533) );
  INV_X1 U4266 ( .A(n3528), .ZN(n3531) );
  OAI21_X1 U4267 ( .B1(n3531), .B2(n3530), .A(n3529), .ZN(n3532) );
  AND4_X1 U4268 ( .A1(n3535), .A2(n3534), .A3(n3533), .A4(n3532), .ZN(n3537)
         );
  OAI21_X1 U4269 ( .B1(n4073), .B2(n3537), .A(n3536), .ZN(n3540) );
  AOI211_X1 U4270 ( .C1(n3541), .C2(n3540), .A(n3539), .B(n3538), .ZN(n3543)
         );
  NOR2_X1 U4271 ( .A1(n3543), .A2(n3542), .ZN(n3545) );
  OAI211_X1 U4272 ( .C1(n3674), .C2(n3713), .A(n3545), .B(n3544), .ZN(n3552)
         );
  INV_X1 U4273 ( .A(n3546), .ZN(n3551) );
  NAND2_X1 U4274 ( .A1(n3548), .A2(n3547), .ZN(n3549) );
  AOI22_X1 U4275 ( .A1(n3552), .A2(n3551), .B1(n3550), .B2(n3549), .ZN(n3553)
         );
  MUX2_X1 U4276 ( .A(n3554), .B(n3553), .S(n2623), .Z(n3555) );
  AOI21_X1 U4277 ( .B1(n3557), .B2(n3556), .A(n3555), .ZN(n3558) );
  XNOR2_X1 U4278 ( .A(n3558), .B(n3982), .ZN(n3565) );
  NAND2_X1 U4279 ( .A1(n3560), .A2(n3559), .ZN(n3561) );
  OAI211_X1 U4280 ( .C1(n3562), .C2(n3564), .A(n3561), .B(B_REG_SCAN_IN), .ZN(
        n3563) );
  OAI21_X1 U4281 ( .B1(n3565), .B2(n3564), .A(n3563), .ZN(U3239) );
  NAND2_X1 U4282 ( .A1(n3566), .A2(n4187), .ZN(n3573) );
  OAI22_X1 U4283 ( .A1(n4187), .A2(n3568), .B1(n3567), .B2(n4476), .ZN(n3571)
         );
  NOR2_X1 U4284 ( .A1(n3569), .A2(n4164), .ZN(n3570) );
  AOI211_X1 U4285 ( .C1(n4012), .C2(n3909), .A(n3571), .B(n3570), .ZN(n3572)
         );
  OAI211_X1 U4286 ( .C1(n3574), .C2(n4147), .A(n3573), .B(n3572), .ZN(U3279)
         );
  OAI22_X1 U4287 ( .A1(n3580), .A2(n3683), .B1(n3682), .B2(n3578), .ZN(n3579)
         );
  XNOR2_X1 U4288 ( .A(n3579), .B(n2068), .ZN(n3586) );
  INV_X1 U4289 ( .A(n3586), .ZN(n3583) );
  OR2_X1 U4290 ( .A1(n3580), .A2(n3680), .ZN(n3582) );
  NAND2_X1 U4291 ( .A1(n3660), .A2(n3782), .ZN(n3581) );
  NAND2_X1 U4292 ( .A1(n3582), .A2(n3581), .ZN(n3584) );
  NAND2_X1 U4293 ( .A1(n3583), .A2(n3584), .ZN(n3776) );
  INV_X1 U4294 ( .A(n3584), .ZN(n3585) );
  OAI22_X1 U4295 ( .A1(n3780), .A2(n3683), .B1(n3682), .B2(n3588), .ZN(n3587)
         );
  XNOR2_X1 U4296 ( .A(n3587), .B(n3675), .ZN(n3842) );
  OAI22_X1 U4297 ( .A1(n3780), .A2(n3680), .B1(n3679), .B2(n3588), .ZN(n3841)
         );
  NAND2_X1 U4298 ( .A1(n3590), .A2(n3589), .ZN(n3605) );
  OAI22_X1 U4299 ( .A1(n3593), .A2(n3683), .B1(n3682), .B2(n3591), .ZN(n3592)
         );
  XNOR2_X1 U4300 ( .A(n3592), .B(n2043), .ZN(n3599) );
  OR2_X1 U4301 ( .A1(n3593), .A2(n3680), .ZN(n3595) );
  NAND2_X1 U4302 ( .A1(n3660), .A2(n3726), .ZN(n3594) );
  NAND2_X1 U4303 ( .A1(n3595), .A2(n3594), .ZN(n3598) );
  OAI22_X1 U4304 ( .A1(n4300), .A2(n3683), .B1(n3682), .B2(n3596), .ZN(n3597)
         );
  XNOR2_X1 U4305 ( .A(n2043), .B(n3597), .ZN(n3606) );
  OR2_X1 U4306 ( .A1(n3720), .A2(n3606), .ZN(n3601) );
  OR2_X1 U4307 ( .A1(n3606), .A2(n3721), .ZN(n3600) );
  OAI21_X1 U4308 ( .B1(n3605), .B2(n3601), .A(n3600), .ZN(n3602) );
  INV_X1 U4309 ( .A(n3602), .ZN(n3798) );
  OR2_X1 U4310 ( .A1(n4300), .A2(n3680), .ZN(n3604) );
  NAND2_X1 U4311 ( .A1(n3660), .A2(n2486), .ZN(n3603) );
  NAND2_X1 U4312 ( .A1(n3798), .A2(n3887), .ZN(n3610) );
  AND2_X1 U4313 ( .A1(n3606), .A2(n3721), .ZN(n3607) );
  OAI22_X1 U4314 ( .A1(n4287), .A2(n3680), .B1(n3679), .B2(n3608), .ZN(n3612)
         );
  OAI22_X1 U4315 ( .A1(n4287), .A2(n3683), .B1(n3682), .B2(n3608), .ZN(n3609)
         );
  XNOR2_X1 U4316 ( .A(n3609), .B(n3675), .ZN(n3611) );
  INV_X1 U4317 ( .A(n3611), .ZN(n3614) );
  INV_X1 U4318 ( .A(n3612), .ZN(n3613) );
  OAI22_X1 U4319 ( .A1(n4294), .A2(n3683), .B1(n3682), .B2(n3616), .ZN(n3617)
         );
  XNOR2_X1 U4320 ( .A(n3617), .B(n2043), .ZN(n3809) );
  OR2_X1 U4321 ( .A1(n4294), .A2(n3680), .ZN(n3619) );
  NAND2_X1 U4322 ( .A1(n3660), .A2(n4282), .ZN(n3618) );
  NAND2_X1 U4323 ( .A1(n3619), .A2(n3618), .ZN(n3810) );
  NOR2_X1 U4324 ( .A1(n3809), .A2(n3810), .ZN(n3862) );
  OAI22_X1 U4325 ( .A1(n4156), .A2(n3683), .B1(n3682), .B2(n4181), .ZN(n3620)
         );
  XNOR2_X1 U4326 ( .A(n3620), .B(n3675), .ZN(n3624) );
  INV_X1 U4327 ( .A(n3624), .ZN(n3622) );
  OAI22_X1 U4328 ( .A1(n4156), .A2(n3680), .B1(n3679), .B2(n4181), .ZN(n3623)
         );
  INV_X1 U4329 ( .A(n3623), .ZN(n3621) );
  NAND2_X1 U4330 ( .A1(n3622), .A2(n3621), .ZN(n3865) );
  INV_X1 U4331 ( .A(n3865), .ZN(n3626) );
  NAND2_X1 U4332 ( .A1(n3809), .A2(n3810), .ZN(n3863) );
  NAND2_X1 U4333 ( .A1(n3624), .A2(n3623), .ZN(n3866) );
  AND2_X1 U4334 ( .A1(n3863), .A2(n3866), .ZN(n3625) );
  OR2_X1 U4335 ( .A1(n3626), .A2(n3625), .ZN(n3753) );
  OAI22_X1 U4336 ( .A1(n3835), .A2(n3680), .B1(n3679), .B2(n4162), .ZN(n3631)
         );
  NAND2_X1 U4337 ( .A1(n4176), .A2(n3660), .ZN(n3628) );
  NAND2_X1 U4338 ( .A1(n2960), .A2(n3758), .ZN(n3627) );
  NAND2_X1 U4339 ( .A1(n3628), .A2(n3627), .ZN(n3629) );
  XNOR2_X1 U4340 ( .A(n3629), .B(n3675), .ZN(n3632) );
  XOR2_X1 U4341 ( .A(n3631), .B(n3632), .Z(n3755) );
  NAND2_X1 U4342 ( .A1(n3754), .A2(n3630), .ZN(n3634) );
  NAND2_X1 U4343 ( .A1(n3634), .A2(n3633), .ZN(n3829) );
  OAI22_X1 U4344 ( .A1(n4120), .A2(n3683), .B1(n3682), .B2(n4140), .ZN(n3635)
         );
  XNOR2_X1 U4345 ( .A(n3635), .B(n3675), .ZN(n3636) );
  OAI22_X1 U4346 ( .A1(n4120), .A2(n3680), .B1(n3679), .B2(n4140), .ZN(n3637)
         );
  NAND2_X1 U4347 ( .A1(n3636), .A2(n3637), .ZN(n3830) );
  INV_X1 U4348 ( .A(n3636), .ZN(n3639) );
  INV_X1 U4349 ( .A(n3637), .ZN(n3638) );
  NAND2_X1 U4350 ( .A1(n3639), .A2(n3638), .ZN(n3831) );
  OAI22_X1 U4351 ( .A1(n4133), .A2(n3683), .B1(n3682), .B2(n4115), .ZN(n3640)
         );
  XNOR2_X1 U4352 ( .A(n3640), .B(n3675), .ZN(n3769) );
  OAI22_X1 U4353 ( .A1(n4133), .A2(n3680), .B1(n3679), .B2(n4115), .ZN(n3768)
         );
  NOR2_X1 U4354 ( .A1(n3769), .A2(n3768), .ZN(n3642) );
  NAND2_X1 U4355 ( .A1(n3769), .A2(n3768), .ZN(n3641) );
  OAI22_X1 U4356 ( .A1(n4265), .A2(n3683), .B1(n3682), .B2(n4095), .ZN(n3643)
         );
  XNOR2_X1 U4357 ( .A(n3643), .B(n3675), .ZN(n3650) );
  OAI22_X1 U4358 ( .A1(n4265), .A2(n3680), .B1(n3679), .B2(n4095), .ZN(n3649)
         );
  XNOR2_X1 U4359 ( .A(n3650), .B(n3649), .ZN(n3853) );
  NAND2_X1 U4360 ( .A1(n4243), .A2(n3660), .ZN(n3646) );
  NAND2_X1 U4361 ( .A1(n2960), .A2(n3644), .ZN(n3645) );
  NAND2_X1 U4362 ( .A1(n3646), .A2(n3645), .ZN(n3647) );
  XNOR2_X1 U4363 ( .A(n3647), .B(n2068), .ZN(n3653) );
  NOR2_X1 U4364 ( .A1(n3679), .A2(n4083), .ZN(n3648) );
  AOI21_X1 U4365 ( .B1(n4243), .B2(n3669), .A(n3648), .ZN(n3652) );
  XNOR2_X1 U4366 ( .A(n3653), .B(n3652), .ZN(n3735) );
  NOR2_X1 U4367 ( .A1(n3650), .A2(n3649), .ZN(n3736) );
  NOR2_X1 U4368 ( .A1(n3735), .A2(n3736), .ZN(n3651) );
  NAND2_X1 U4369 ( .A1(n3734), .A2(n3651), .ZN(n3733) );
  NOR2_X1 U4370 ( .A1(n3653), .A2(n3652), .ZN(n3656) );
  OAI22_X1 U4371 ( .A1(n4050), .A2(n3680), .B1(n3679), .B2(n3823), .ZN(n3658)
         );
  NAND2_X1 U4372 ( .A1(n3733), .A2(n3654), .ZN(n3820) );
  OAI22_X1 U4373 ( .A1(n4050), .A2(n3683), .B1(n3682), .B2(n3823), .ZN(n3655)
         );
  XNOR2_X1 U4374 ( .A(n3655), .B(n3675), .ZN(n3822) );
  INV_X1 U4375 ( .A(n3656), .ZN(n3657) );
  NAND2_X1 U4376 ( .A1(n3733), .A2(n3657), .ZN(n3659) );
  NAND2_X1 U4377 ( .A1(n4063), .A2(n3660), .ZN(n3662) );
  NAND2_X1 U4378 ( .A1(n2960), .A2(n4233), .ZN(n3661) );
  NAND2_X1 U4379 ( .A1(n3662), .A2(n3661), .ZN(n3663) );
  XNOR2_X1 U4380 ( .A(n3663), .B(n2068), .ZN(n3666) );
  NOR2_X1 U4381 ( .A1(n3679), .A2(n4045), .ZN(n3664) );
  AOI21_X1 U4382 ( .B1(n4063), .B2(n3669), .A(n3664), .ZN(n3665) );
  NAND2_X1 U4383 ( .A1(n3666), .A2(n3665), .ZN(n3790) );
  NOR2_X1 U4384 ( .A1(n3666), .A2(n3665), .ZN(n3791) );
  OAI22_X1 U4385 ( .A1(n4237), .A2(n3683), .B1(n3682), .B2(n4032), .ZN(n3667)
         );
  XNOR2_X1 U4386 ( .A(n3667), .B(n2068), .ZN(n3673) );
  INV_X1 U4387 ( .A(n3673), .ZN(n3671) );
  NOR2_X1 U4388 ( .A1(n3683), .A2(n4032), .ZN(n3668) );
  AOI21_X1 U4389 ( .B1(n4046), .B2(n3669), .A(n3668), .ZN(n3672) );
  INV_X1 U4390 ( .A(n3672), .ZN(n3670) );
  NAND2_X1 U4391 ( .A1(n3671), .A2(n3670), .ZN(n3875) );
  AND2_X1 U4392 ( .A1(n3673), .A2(n3672), .ZN(n3874) );
  OAI22_X1 U4393 ( .A1(n3674), .A2(n3680), .B1(n4221), .B2(n3679), .ZN(n3678)
         );
  OAI22_X1 U4394 ( .A1(n3674), .A2(n3683), .B1(n4221), .B2(n3682), .ZN(n3676)
         );
  XNOR2_X1 U4395 ( .A(n3676), .B(n3675), .ZN(n3677) );
  XOR2_X1 U4396 ( .A(n3678), .B(n3677), .Z(n3711) );
  AOI22_X1 U4397 ( .A1(n3712), .A2(n3711), .B1(n3678), .B2(n3677), .ZN(n3688)
         );
  OAI22_X1 U4398 ( .A1(n3684), .A2(n3680), .B1(n3679), .B2(n3700), .ZN(n3681)
         );
  XNOR2_X1 U4399 ( .A(n3681), .B(n2043), .ZN(n3686) );
  OAI22_X1 U4400 ( .A1(n3684), .A2(n3683), .B1(n3682), .B2(n3700), .ZN(n3685)
         );
  XNOR2_X1 U4401 ( .A(n3686), .B(n3685), .ZN(n3687) );
  XNOR2_X1 U4402 ( .A(n3688), .B(n3687), .ZN(n3696) );
  NAND2_X1 U4403 ( .A1(n3901), .A2(n3889), .ZN(n3693) );
  OR2_X1 U4404 ( .A1(n3699), .A2(n3895), .ZN(n3692) );
  NAND2_X1 U4405 ( .A1(n3890), .A2(n3689), .ZN(n3691) );
  NAND2_X1 U4406 ( .A1(U3149), .A2(REG3_REG_28__SCAN_IN), .ZN(n3690) );
  NAND4_X1 U4407 ( .A1(n3693), .A2(n3692), .A3(n3691), .A4(n3690), .ZN(n3694)
         );
  AOI21_X1 U4408 ( .B1(n4028), .B2(n3891), .A(n3694), .ZN(n3695) );
  OAI21_X1 U4409 ( .B1(n3696), .B2(n3884), .A(n3695), .ZN(U3217) );
  INV_X1 U4410 ( .A(n3697), .ZN(n3708) );
  INV_X1 U4411 ( .A(REG2_REG_28__SCAN_IN), .ZN(n3698) );
  OAI22_X1 U4412 ( .A1(n3699), .A2(n4476), .B1(n3698), .B2(n4187), .ZN(n3704)
         );
  OAI22_X1 U4413 ( .A1(n3702), .A2(n3701), .B1(n3700), .B2(n4015), .ZN(n3703)
         );
  AOI211_X1 U4414 ( .C1(n4012), .C2(n4028), .A(n3704), .B(n3703), .ZN(n3705)
         );
  OAI21_X1 U4415 ( .B1(n3706), .B2(n4164), .A(n3705), .ZN(n3707) );
  AOI21_X1 U4416 ( .B1(n3708), .B2(n4187), .A(n3707), .ZN(n3709) );
  OAI21_X1 U4417 ( .B1(n3710), .B2(n4210), .A(n3709), .ZN(U3262) );
  XNOR2_X1 U4418 ( .A(n3712), .B(n3711), .ZN(n3719) );
  NAND2_X1 U4419 ( .A1(U3149), .A2(REG3_REG_27__SCAN_IN), .ZN(n3715) );
  NAND2_X1 U4420 ( .A1(n3890), .A2(n3713), .ZN(n3714) );
  OAI211_X1 U4421 ( .C1(n4237), .C2(n3856), .A(n3715), .B(n3714), .ZN(n3716)
         );
  AOI21_X1 U4422 ( .B1(n3889), .B2(n4224), .A(n3716), .ZN(n3718) );
  INV_X1 U4423 ( .A(n3895), .ZN(n3878) );
  NAND2_X1 U4424 ( .A1(n4011), .A2(n3878), .ZN(n3717) );
  OAI211_X1 U4425 ( .C1(n3719), .C2(n3884), .A(n3718), .B(n3717), .ZN(U3211)
         );
  INV_X1 U4426 ( .A(n3720), .ZN(n3722) );
  NAND2_X1 U4427 ( .A1(n3722), .A2(n3721), .ZN(n3723) );
  XNOR2_X1 U4428 ( .A(n3605), .B(n3723), .ZN(n3731) );
  NOR2_X1 U4429 ( .A1(n4660), .A2(STATE_REG_SCAN_IN), .ZN(n4427) );
  INV_X1 U4430 ( .A(n4427), .ZN(n3724) );
  OAI21_X1 U4431 ( .B1(n3857), .B2(n4300), .A(n3724), .ZN(n3725) );
  INV_X1 U4432 ( .A(n3725), .ZN(n3728) );
  AOI22_X1 U4433 ( .A1(n3891), .A2(n3906), .B1(n3890), .B2(n3726), .ZN(n3727)
         );
  OAI211_X1 U4434 ( .C1(n3895), .C2(n3729), .A(n3728), .B(n3727), .ZN(n3730)
         );
  AOI21_X1 U4435 ( .B1(n3731), .B2(n3897), .A(n3730), .ZN(n3732) );
  INV_X1 U4436 ( .A(n3732), .ZN(U3212) );
  INV_X1 U4437 ( .A(n3734), .ZN(n3851) );
  OAI21_X1 U4438 ( .B1(n3851), .B2(n3736), .A(n3735), .ZN(n3737) );
  NAND3_X1 U4439 ( .A1(n3733), .A2(n3737), .A3(n3897), .ZN(n3741) );
  NOR2_X1 U4440 ( .A1(n4265), .A2(n3856), .ZN(n3739) );
  OAI22_X1 U4441 ( .A1(n4050), .A2(n3857), .B1(n3881), .B2(n4083), .ZN(n3738)
         );
  AOI211_X1 U4442 ( .C1(REG3_REG_23__SCAN_IN), .C2(U3149), .A(n3739), .B(n3738), .ZN(n3740) );
  OAI211_X1 U4443 ( .C1(n3895), .C2(n4085), .A(n3741), .B(n3740), .ZN(U3213)
         );
  OAI211_X1 U4444 ( .C1(n3744), .C2(n3743), .A(n3742), .B(n3897), .ZN(n3752)
         );
  NAND2_X1 U4445 ( .A1(REG3_REG_10__SCAN_IN), .A2(U3149), .ZN(n4384) );
  OAI21_X1 U4446 ( .B1(n3857), .B2(n3745), .A(n4384), .ZN(n3746) );
  INV_X1 U4447 ( .A(n3746), .ZN(n3751) );
  AOI22_X1 U4448 ( .A1(n3891), .A2(n3910), .B1(n3890), .B2(n3747), .ZN(n3750)
         );
  OR2_X1 U4449 ( .A1(n3895), .A2(n3748), .ZN(n3749) );
  NAND4_X1 U4450 ( .A1(n3752), .A2(n3751), .A3(n3750), .A4(n3749), .ZN(U3214)
         );
  AND2_X1 U4451 ( .A1(n3754), .A2(n3753), .ZN(n3756) );
  XNOR2_X1 U4452 ( .A(n3756), .B(n3755), .ZN(n3762) );
  NAND2_X1 U4453 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n3981) );
  OAI21_X1 U4454 ( .B1(n3857), .B2(n4120), .A(n3981), .ZN(n3757) );
  INV_X1 U4455 ( .A(n3757), .ZN(n3760) );
  AOI22_X1 U4456 ( .A1(n3891), .A2(n4284), .B1(n3890), .B2(n3758), .ZN(n3759)
         );
  OAI211_X1 U4457 ( .C1(n3895), .C2(n4165), .A(n3760), .B(n3759), .ZN(n3761)
         );
  AOI21_X1 U4458 ( .B1(n3762), .B2(n3897), .A(n3761), .ZN(n3763) );
  INV_X1 U4459 ( .A(n3763), .ZN(U3216) );
  AOI22_X1 U4460 ( .A1(n3891), .A2(n4262), .B1(n3890), .B2(n4260), .ZN(n3765)
         );
  NAND2_X1 U4461 ( .A1(n4116), .A2(n3889), .ZN(n3764) );
  OAI211_X1 U4462 ( .C1(STATE_REG_SCAN_IN), .C2(n3766), .A(n3765), .B(n3764), 
        .ZN(n3773) );
  XNOR2_X1 U4463 ( .A(n3769), .B(n3768), .ZN(n3770) );
  XNOR2_X1 U4464 ( .A(n3767), .B(n3770), .ZN(n3771) );
  NOR2_X1 U4465 ( .A1(n3771), .A2(n3884), .ZN(n3772) );
  AOI211_X1 U4466 ( .C1(n4117), .C2(n3878), .A(n3773), .B(n3772), .ZN(n3774)
         );
  INV_X1 U4467 ( .A(n3774), .ZN(U3220) );
  INV_X1 U4468 ( .A(n3776), .ZN(n3778) );
  NOR2_X1 U4469 ( .A1(n3778), .A2(n3777), .ZN(n3779) );
  XNOR2_X1 U4470 ( .A(n3775), .B(n3779), .ZN(n3787) );
  NAND2_X1 U4471 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4404) );
  OAI21_X1 U4472 ( .B1(n3857), .B2(n3780), .A(n4404), .ZN(n3781) );
  INV_X1 U4473 ( .A(n3781), .ZN(n3784) );
  AOI22_X1 U4474 ( .A1(n3891), .A2(n3908), .B1(n3890), .B2(n3782), .ZN(n3783)
         );
  OAI211_X1 U4475 ( .C1(n3895), .C2(n3785), .A(n3784), .B(n3783), .ZN(n3786)
         );
  AOI21_X1 U4476 ( .B1(n3787), .B2(n3897), .A(n3786), .ZN(n3788) );
  INV_X1 U4477 ( .A(n3788), .ZN(U3221) );
  NOR2_X1 U4478 ( .A1(n3791), .A2(n2229), .ZN(n3792) );
  XNOR2_X1 U4479 ( .A(n3789), .B(n3792), .ZN(n3797) );
  INV_X1 U4480 ( .A(n3793), .ZN(n4047) );
  OAI22_X1 U4481 ( .A1(n4050), .A2(n3856), .B1(STATE_REG_SCAN_IN), .B2(n4542), 
        .ZN(n3795) );
  OAI22_X1 U4482 ( .A1(n4237), .A2(n3857), .B1(n3881), .B2(n4045), .ZN(n3794)
         );
  AOI211_X1 U4483 ( .C1(n4047), .C2(n3878), .A(n3795), .B(n3794), .ZN(n3796)
         );
  OAI21_X1 U4484 ( .B1(n3797), .B2(n3884), .A(n3796), .ZN(U3222) );
  INV_X1 U4485 ( .A(n3886), .ZN(n3799) );
  OAI21_X1 U4486 ( .B1(n3799), .B2(n3887), .A(n3798), .ZN(n3801) );
  XNOR2_X1 U4487 ( .A(n3801), .B(n3800), .ZN(n3806) );
  NAND2_X1 U4488 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4443) );
  OAI21_X1 U4489 ( .B1(n3857), .B2(n4294), .A(n4443), .ZN(n3802) );
  INV_X1 U4490 ( .A(n3802), .ZN(n3804) );
  AOI22_X1 U4491 ( .A1(n3891), .A2(n2487), .B1(n3890), .B2(n4296), .ZN(n3803)
         );
  OAI211_X1 U4492 ( .C1(n3895), .C2(n4198), .A(n3804), .B(n3803), .ZN(n3805)
         );
  AOI21_X1 U4493 ( .B1(n3806), .B2(n3897), .A(n3805), .ZN(n3807) );
  INV_X1 U4494 ( .A(n3807), .ZN(U3223) );
  XOR2_X1 U4495 ( .A(n3810), .B(n3809), .Z(n3811) );
  XNOR2_X1 U4496 ( .A(n3808), .B(n3811), .ZN(n3817) );
  INV_X1 U4497 ( .A(n3812), .ZN(n3815) );
  AND2_X1 U4498 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4457) );
  AOI21_X1 U4499 ( .B1(n3889), .B2(n4284), .A(n4457), .ZN(n3814) );
  AOI22_X1 U4500 ( .A1(n3891), .A2(n3904), .B1(n3890), .B2(n4282), .ZN(n3813)
         );
  OAI211_X1 U4501 ( .C1(n3895), .C2(n3815), .A(n3814), .B(n3813), .ZN(n3816)
         );
  AOI21_X1 U4502 ( .B1(n3817), .B2(n3897), .A(n3816), .ZN(n3818) );
  INV_X1 U4503 ( .A(n3818), .ZN(U3225) );
  NAND2_X1 U4504 ( .A1(n3819), .A2(n3820), .ZN(n3821) );
  XOR2_X1 U4505 ( .A(n3822), .B(n3821), .Z(n3827) );
  OAI22_X1 U4506 ( .A1(n4067), .A2(n3856), .B1(STATE_REG_SCAN_IN), .B2(n4698), 
        .ZN(n3825) );
  OAI22_X1 U4507 ( .A1(n4246), .A2(n3857), .B1(n3881), .B2(n3823), .ZN(n3824)
         );
  AOI211_X1 U4508 ( .C1(n4064), .C2(n3878), .A(n3825), .B(n3824), .ZN(n3826)
         );
  OAI21_X1 U4509 ( .B1(n3827), .B2(n3884), .A(n3826), .ZN(U3226) );
  NOR2_X1 U4510 ( .A1(n3828), .A2(n2205), .ZN(n3833) );
  AOI21_X1 U4511 ( .B1(n3831), .B2(n3830), .A(n3829), .ZN(n3832) );
  OAI21_X1 U4512 ( .B1(n3833), .B2(n3832), .A(n3897), .ZN(n3839) );
  NAND2_X1 U4513 ( .A1(n3890), .A2(n4131), .ZN(n3834) );
  OAI21_X1 U4514 ( .B1(n3835), .B2(n3856), .A(n3834), .ZN(n3837) );
  OAI22_X1 U4515 ( .A1(n3857), .A2(n4133), .B1(STATE_REG_SCAN_IN), .B2(n4669), 
        .ZN(n3836) );
  NOR2_X1 U4516 ( .A1(n3837), .A2(n3836), .ZN(n3838) );
  OAI211_X1 U4517 ( .C1(n3895), .C2(n4141), .A(n3839), .B(n3838), .ZN(U3230)
         );
  XNOR2_X1 U4518 ( .A(n3842), .B(n3841), .ZN(n3843) );
  XNOR2_X1 U4519 ( .A(n3840), .B(n3843), .ZN(n3849) );
  NOR2_X1 U4520 ( .A1(STATE_REG_SCAN_IN), .A2(n2452), .ZN(n4417) );
  AOI21_X1 U4521 ( .B1(n3889), .B2(n3905), .A(n4417), .ZN(n3846) );
  AOI22_X1 U4522 ( .A1(n3891), .A2(n3907), .B1(n3890), .B2(n3844), .ZN(n3845)
         );
  OAI211_X1 U4523 ( .C1(n3895), .C2(n3847), .A(n3846), .B(n3845), .ZN(n3848)
         );
  AOI21_X1 U4524 ( .B1(n3849), .B2(n3897), .A(n3848), .ZN(n3850) );
  INV_X1 U4525 ( .A(n3850), .ZN(U3231) );
  AOI21_X1 U4526 ( .B1(n3853), .B2(n3852), .A(n3851), .ZN(n3861) );
  INV_X1 U4527 ( .A(n3854), .ZN(n4098) );
  OAI22_X1 U4528 ( .A1(n3856), .A2(n4133), .B1(STATE_REG_SCAN_IN), .B2(n3855), 
        .ZN(n3859) );
  OAI22_X1 U4529 ( .A1(n4067), .A2(n3857), .B1(n3881), .B2(n4095), .ZN(n3858)
         );
  AOI211_X1 U4530 ( .C1(n4098), .C2(n3878), .A(n3859), .B(n3858), .ZN(n3860)
         );
  OAI21_X1 U4531 ( .B1(n3861), .B2(n3884), .A(n3860), .ZN(U3232) );
  OR2_X1 U4532 ( .A1(n3808), .A2(n3862), .ZN(n3864) );
  NAND2_X1 U4533 ( .A1(n3864), .A2(n3863), .ZN(n3868) );
  NAND2_X1 U4534 ( .A1(n3866), .A2(n3865), .ZN(n3867) );
  XNOR2_X1 U4535 ( .A(n3868), .B(n3867), .ZN(n3872) );
  AND2_X1 U4536 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4467) );
  AOI21_X1 U4537 ( .B1(n3889), .B2(n4176), .A(n4467), .ZN(n3870) );
  AOI22_X1 U4538 ( .A1(n3891), .A2(n4195), .B1(n3890), .B2(n4175), .ZN(n3869)
         );
  OAI211_X1 U4539 ( .C1(n3895), .C2(n4184), .A(n3870), .B(n3869), .ZN(n3871)
         );
  AOI21_X1 U4540 ( .B1(n3872), .B2(n3897), .A(n3871), .ZN(n3873) );
  INV_X1 U4541 ( .A(n3873), .ZN(U3235) );
  NAND2_X1 U4542 ( .A1(n2227), .A2(n3875), .ZN(n3876) );
  XNOR2_X1 U4543 ( .A(n3877), .B(n3876), .ZN(n3885) );
  AOI22_X1 U4544 ( .A1(n4063), .A2(n3891), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n3880) );
  NAND2_X1 U4545 ( .A1(n4033), .A2(n3878), .ZN(n3879) );
  OAI211_X1 U4546 ( .C1(n3881), .C2(n4032), .A(n3880), .B(n3879), .ZN(n3882)
         );
  AOI21_X1 U4547 ( .B1(n4028), .B2(n3889), .A(n3882), .ZN(n3883) );
  OAI21_X1 U4548 ( .B1(n3885), .B2(n3884), .A(n3883), .ZN(U3237) );
  NAND2_X1 U4549 ( .A1(n3886), .A2(n3798), .ZN(n3888) );
  XNOR2_X1 U4550 ( .A(n3888), .B(n3887), .ZN(n3898) );
  AND2_X1 U4551 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4437) );
  AOI21_X1 U4552 ( .B1(n3889), .B2(n3904), .A(n4437), .ZN(n3893) );
  AOI22_X1 U4553 ( .A1(n3891), .A2(n3905), .B1(n3890), .B2(n2486), .ZN(n3892)
         );
  OAI211_X1 U4554 ( .C1(n3895), .C2(n3894), .A(n3893), .B(n3892), .ZN(n3896)
         );
  AOI21_X1 U4555 ( .B1(n3898), .B2(n3897), .A(n3896), .ZN(n3899) );
  INV_X1 U4556 ( .A(n3899), .ZN(U3238) );
  MUX2_X1 U4557 ( .A(DATAO_REG_31__SCAN_IN), .B(n3988), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4558 ( .A(DATAO_REG_30__SCAN_IN), .B(n3900), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4559 ( .A(DATAO_REG_29__SCAN_IN), .B(n3901), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4560 ( .A(DATAO_REG_28__SCAN_IN), .B(n4224), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4561 ( .A(DATAO_REG_27__SCAN_IN), .B(n4028), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4562 ( .A(DATAO_REG_26__SCAN_IN), .B(n4046), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4563 ( .A(DATAO_REG_25__SCAN_IN), .B(n4063), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4564 ( .A(DATAO_REG_24__SCAN_IN), .B(n4234), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4565 ( .A(n4243), .B(DATAO_REG_23__SCAN_IN), .S(n3903), .Z(U3573)
         );
  MUX2_X1 U4566 ( .A(n4116), .B(DATAO_REG_22__SCAN_IN), .S(n3903), .Z(U3572)
         );
  MUX2_X1 U4567 ( .A(n3902), .B(DATAO_REG_21__SCAN_IN), .S(n3903), .Z(U3571)
         );
  MUX2_X1 U4568 ( .A(n4262), .B(DATAO_REG_20__SCAN_IN), .S(n3903), .Z(U3570)
         );
  MUX2_X1 U4569 ( .A(n4176), .B(DATAO_REG_19__SCAN_IN), .S(n3903), .Z(U3569)
         );
  MUX2_X1 U4570 ( .A(DATAO_REG_18__SCAN_IN), .B(n4284), .S(U4043), .Z(U3568)
         );
  MUX2_X1 U4571 ( .A(DATAO_REG_17__SCAN_IN), .B(n4195), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4572 ( .A(DATAO_REG_16__SCAN_IN), .B(n3904), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4573 ( .A(DATAO_REG_15__SCAN_IN), .B(n2487), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U4574 ( .A(DATAO_REG_14__SCAN_IN), .B(n3905), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4575 ( .A(DATAO_REG_13__SCAN_IN), .B(n3906), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4576 ( .A(DATAO_REG_12__SCAN_IN), .B(n3907), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4577 ( .A(DATAO_REG_11__SCAN_IN), .B(n3908), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4578 ( .A(DATAO_REG_10__SCAN_IN), .B(n3909), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4579 ( .A(DATAO_REG_9__SCAN_IN), .B(n3910), .S(U4043), .Z(U3559) );
  MUX2_X1 U4580 ( .A(DATAO_REG_8__SCAN_IN), .B(n3911), .S(U4043), .Z(U3558) );
  MUX2_X1 U4581 ( .A(DATAO_REG_7__SCAN_IN), .B(n3912), .S(U4043), .Z(U3557) );
  MUX2_X1 U4582 ( .A(DATAO_REG_6__SCAN_IN), .B(n3913), .S(U4043), .Z(U3556) );
  MUX2_X1 U4583 ( .A(DATAO_REG_5__SCAN_IN), .B(n3914), .S(U4043), .Z(U3555) );
  MUX2_X1 U4584 ( .A(DATAO_REG_4__SCAN_IN), .B(n3915), .S(U4043), .Z(U3554) );
  MUX2_X1 U4585 ( .A(DATAO_REG_3__SCAN_IN), .B(n2959), .S(U4043), .Z(U3553) );
  MUX2_X1 U4586 ( .A(DATAO_REG_2__SCAN_IN), .B(n3916), .S(U4043), .Z(U3552) );
  MUX2_X1 U4587 ( .A(DATAO_REG_1__SCAN_IN), .B(n3917), .S(U4043), .Z(U3551) );
  MUX2_X1 U4588 ( .A(DATAO_REG_0__SCAN_IN), .B(n2852), .S(U4043), .Z(U3550) );
  INV_X1 U4589 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4530) );
  NAND3_X1 U4590 ( .A1(n4470), .A2(IR_REG_0__SCAN_IN), .A3(n4530), .ZN(n3926)
         );
  AOI21_X1 U4591 ( .B1(n4530), .B2(n3918), .A(n3921), .ZN(n3920) );
  MUX2_X1 U4592 ( .A(n3921), .B(n3920), .S(n3919), .Z(n3922) );
  AOI22_X1 U4593 ( .A1(n3923), .A2(n3922), .B1(REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n3925) );
  NAND2_X1 U4594 ( .A1(n4468), .A2(ADDR_REG_0__SCAN_IN), .ZN(n3924) );
  NAND3_X1 U4595 ( .A1(n3926), .A2(n3925), .A3(n3924), .ZN(U3240) );
  OAI211_X1 U4596 ( .C1(n3930), .C2(n3929), .A(n4470), .B(n3928), .ZN(n3936)
         );
  OAI211_X1 U4597 ( .C1(n2776), .C2(n3933), .A(n4413), .B(n3932), .ZN(n3935)
         );
  AOI22_X1 U4598 ( .A1(n4468), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3934) );
  NAND4_X1 U4599 ( .A1(n3937), .A2(n3936), .A3(n3935), .A4(n3934), .ZN(U3241)
         );
  INV_X1 U4600 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3938) );
  MUX2_X1 U4601 ( .A(REG2_REG_19__SCAN_IN), .B(n3938), .S(n4360), .Z(n3953) );
  INV_X1 U4602 ( .A(n3954), .ZN(n4498) );
  INV_X1 U4603 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3939) );
  AOI22_X1 U4604 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4498), .B1(n3954), .B2(
        n3939), .ZN(n4466) );
  NOR2_X1 U4605 ( .A1(n4499), .A2(REG2_REG_17__SCAN_IN), .ZN(n3940) );
  AOI21_X1 U4606 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4499), .A(n3940), .ZN(n4455) );
  INV_X1 U4607 ( .A(n4503), .ZN(n4432) );
  NOR2_X1 U4608 ( .A1(n4412), .A2(n4505), .ZN(n4411) );
  NAND2_X1 U4609 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3957), .ZN(n3945) );
  INV_X1 U4610 ( .A(n3957), .ZN(n4507) );
  AOI22_X1 U4611 ( .A1(REG2_REG_11__SCAN_IN), .A2(n3957), .B1(n4507), .B2(
        n3568), .ZN(n4396) );
  NAND2_X1 U4612 ( .A1(n3958), .A2(REG2_REG_9__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4613 ( .A1(n3958), .A2(REG2_REG_9__SCAN_IN), .B1(n2372), .B2(n4510), .ZN(n4376) );
  NAND2_X1 U4614 ( .A1(n4376), .A2(n4375), .ZN(n4374) );
  NAND2_X1 U4615 ( .A1(n3942), .A2(n4374), .ZN(n3943) );
  NAND2_X1 U4616 ( .A1(n3963), .A2(n3943), .ZN(n3944) );
  INV_X1 U4617 ( .A(n3963), .ZN(n4508) );
  XNOR2_X1 U4618 ( .A(n3943), .B(n4508), .ZN(n4383) );
  NAND2_X1 U4619 ( .A1(n3967), .A2(n3946), .ZN(n3947) );
  XNOR2_X1 U4620 ( .A(n3946), .B(n4506), .ZN(n4403) );
  NOR2_X1 U4621 ( .A1(n4432), .A2(n3948), .ZN(n3949) );
  NOR2_X1 U4622 ( .A1(n2466), .A2(n4425), .ZN(n4424) );
  NOR2_X1 U4623 ( .A1(n3949), .A2(n4424), .ZN(n4435) );
  NAND2_X1 U4624 ( .A1(REG2_REG_15__SCAN_IN), .A2(n3955), .ZN(n3950) );
  OAI21_X1 U4625 ( .B1(REG2_REG_15__SCAN_IN), .B2(n3955), .A(n3950), .ZN(n4434) );
  INV_X1 U4626 ( .A(n3974), .ZN(n4501) );
  NAND2_X1 U4627 ( .A1(n3951), .A2(n4501), .ZN(n3952) );
  INV_X1 U4628 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4444) );
  NAND2_X1 U4629 ( .A1(n3952), .A2(n4445), .ZN(n4453) );
  NAND2_X1 U4630 ( .A1(n4455), .A2(n4453), .ZN(n4454) );
  AOI22_X1 U4631 ( .A1(REG1_REG_18__SCAN_IN), .A2(n3954), .B1(n4498), .B2(
        n3978), .ZN(n4472) );
  NOR2_X1 U4632 ( .A1(n4499), .A2(REG1_REG_17__SCAN_IN), .ZN(n3977) );
  NAND2_X1 U4633 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3955), .ZN(n3973) );
  AOI22_X1 U4634 ( .A1(REG1_REG_15__SCAN_IN), .A2(n3955), .B1(n4502), .B2(
        n3392), .ZN(n4440) );
  NAND2_X1 U4635 ( .A1(REG1_REG_13__SCAN_IN), .A2(n3956), .ZN(n3970) );
  AOI22_X1 U4636 ( .A1(REG1_REG_13__SCAN_IN), .A2(n3956), .B1(n4505), .B2(
        n3382), .ZN(n4421) );
  NAND2_X1 U4637 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3957), .ZN(n3966) );
  AOI22_X1 U4638 ( .A1(REG1_REG_11__SCAN_IN), .A2(n3957), .B1(n4507), .B2(
        n3314), .ZN(n4393) );
  NAND2_X1 U4639 ( .A1(n3958), .A2(REG1_REG_9__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U4640 ( .A1(n3958), .A2(REG1_REG_9__SCAN_IN), .B1(n2371), .B2(n4510), .ZN(n4373) );
  INV_X1 U4641 ( .A(n3960), .ZN(n3961) );
  NAND2_X1 U4642 ( .A1(n3963), .A2(n3964), .ZN(n3965) );
  XNOR2_X1 U4643 ( .A(n3964), .B(n4508), .ZN(n4388) );
  NAND2_X1 U4644 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4388), .ZN(n4387) );
  NAND2_X1 U4645 ( .A1(n3967), .A2(n3968), .ZN(n3969) );
  NAND2_X1 U4646 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4408), .ZN(n4407) );
  NAND2_X1 U4647 ( .A1(n4503), .A2(n3971), .ZN(n3972) );
  NAND2_X1 U4648 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4429), .ZN(n4428) );
  NAND2_X1 U4649 ( .A1(n3972), .A2(n4428), .ZN(n4439) );
  NAND2_X1 U4650 ( .A1(n4440), .A2(n4439), .ZN(n4438) );
  NOR2_X1 U4651 ( .A1(n3974), .A2(n3975), .ZN(n3976) );
  AOI22_X1 U4652 ( .A1(n4499), .A2(n4290), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4463), .ZN(n4458) );
  NOR2_X1 U4653 ( .A1(n4459), .A2(n4458), .ZN(n4460) );
  MUX2_X1 U4654 ( .A(n4277), .B(REG1_REG_19__SCAN_IN), .S(n4360), .Z(n3979) );
  NAND2_X1 U4655 ( .A1(n4468), .A2(ADDR_REG_19__SCAN_IN), .ZN(n3980) );
  OAI211_X1 U4656 ( .C1(n4475), .C2(n3982), .A(n3981), .B(n3980), .ZN(n3983)
         );
  AOI21_X1 U4657 ( .B1(n3984), .B2(n4470), .A(n3983), .ZN(n3985) );
  OAI21_X1 U4658 ( .B1(n3986), .B2(n4464), .A(n3985), .ZN(U3259) );
  NOR2_X2 U4659 ( .A1(n4215), .A2(n4218), .ZN(n4214) );
  XNOR2_X1 U4660 ( .A(n4214), .B(n3989), .ZN(n4311) );
  NAND2_X1 U4661 ( .A1(n3988), .A2(n3987), .ZN(n4216) );
  OAI21_X1 U4662 ( .B1(n3989), .B2(n4220), .A(n4216), .ZN(n4308) );
  NAND2_X1 U4663 ( .A1(n4106), .A2(n4308), .ZN(n3991) );
  NAND2_X1 U4664 ( .A1(n4367), .A2(REG2_REG_31__SCAN_IN), .ZN(n3990) );
  OAI211_X1 U4665 ( .C1(n4311), .C2(n4164), .A(n3991), .B(n3990), .ZN(U3260)
         );
  INV_X1 U4666 ( .A(n3992), .ZN(n4003) );
  INV_X1 U4667 ( .A(REG2_REG_29__SCAN_IN), .ZN(n3993) );
  OAI22_X1 U4668 ( .A1(n4015), .A2(n3994), .B1(n3993), .B2(n4187), .ZN(n3995)
         );
  AOI21_X1 U4669 ( .B1(n4224), .B2(n4012), .A(n3995), .ZN(n4002) );
  INV_X1 U4670 ( .A(n3996), .ZN(n4000) );
  OAI22_X1 U4671 ( .A1(n3998), .A2(n4164), .B1(n3997), .B2(n4476), .ZN(n3999)
         );
  OAI21_X1 U4672 ( .B1(n4000), .B2(n3999), .A(n4187), .ZN(n4001) );
  OAI211_X1 U4673 ( .C1(n4003), .C2(n4210), .A(n4002), .B(n4001), .ZN(U3354)
         );
  XNOR2_X1 U4674 ( .A(n4004), .B(n4005), .ZN(n4226) );
  NAND2_X1 U4675 ( .A1(n4006), .A2(n4005), .ZN(n4007) );
  AOI21_X1 U4676 ( .B1(n4008), .B2(n4007), .A(n4159), .ZN(n4222) );
  INV_X1 U4677 ( .A(n4031), .ZN(n4010) );
  OAI21_X1 U4678 ( .B1(n4010), .B2(n4221), .A(n4009), .ZN(n4318) );
  NOR2_X1 U4679 ( .A1(n4318), .A2(n4164), .ZN(n4017) );
  AOI22_X1 U4680 ( .A1(n4224), .A2(n4196), .B1(n4011), .B2(n4486), .ZN(n4014)
         );
  AOI22_X1 U4681 ( .A1(n4046), .A2(n4012), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4367), .ZN(n4013) );
  OAI211_X1 U4682 ( .C1(n4221), .C2(n4015), .A(n4014), .B(n4013), .ZN(n4016)
         );
  AOI211_X1 U4683 ( .C1(n4222), .C2(n4187), .A(n4017), .B(n4016), .ZN(n4018)
         );
  OAI21_X1 U4684 ( .B1(n4226), .B2(n4210), .A(n4018), .ZN(U3263) );
  XNOR2_X1 U4685 ( .A(n4020), .B(n4019), .ZN(n4230) );
  INV_X1 U4686 ( .A(n4230), .ZN(n4037) );
  INV_X1 U4687 ( .A(n4021), .ZN(n4024) );
  OAI21_X1 U4688 ( .B1(n4024), .B2(n4023), .A(n4022), .ZN(n4026) );
  XNOR2_X1 U4689 ( .A(n4026), .B(n4025), .ZN(n4030) );
  OAI22_X1 U4690 ( .A1(n4246), .A2(n4299), .B1(n4032), .B2(n4220), .ZN(n4027)
         );
  AOI21_X1 U4691 ( .B1(n4028), .B2(n4283), .A(n4027), .ZN(n4029) );
  OAI21_X1 U4692 ( .B1(n4030), .B2(n4159), .A(n4029), .ZN(n4229) );
  OAI21_X1 U4693 ( .B1(n4043), .B2(n4032), .A(n4031), .ZN(n4322) );
  AOI22_X1 U4694 ( .A1(n4033), .A2(n4486), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4367), .ZN(n4034) );
  OAI21_X1 U4695 ( .B1(n4322), .B2(n4164), .A(n4034), .ZN(n4035) );
  AOI21_X1 U4696 ( .B1(n4229), .B2(n4187), .A(n4035), .ZN(n4036) );
  OAI21_X1 U4697 ( .B1(n4037), .B2(n4210), .A(n4036), .ZN(U3264) );
  NAND2_X1 U4698 ( .A1(n4021), .A2(n4038), .ZN(n4039) );
  XNOR2_X1 U4699 ( .A(n4039), .B(n4042), .ZN(n4040) );
  NAND2_X1 U4700 ( .A1(n4040), .A2(n4203), .ZN(n4236) );
  XNOR2_X1 U4701 ( .A(n4041), .B(n4042), .ZN(n4239) );
  NAND2_X1 U4702 ( .A1(n4239), .A2(n4112), .ZN(n4054) );
  INV_X1 U4703 ( .A(n4043), .ZN(n4044) );
  OAI21_X1 U4704 ( .B1(n4061), .B2(n4045), .A(n4044), .ZN(n4326) );
  INV_X1 U4705 ( .A(n4326), .ZN(n4052) );
  AOI22_X1 U4706 ( .A1(n4046), .A2(n4196), .B1(n4197), .B2(n4233), .ZN(n4049)
         );
  AOI22_X1 U4707 ( .A1(n4047), .A2(n4486), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4367), .ZN(n4048) );
  OAI211_X1 U4708 ( .C1(n4050), .C2(n4202), .A(n4049), .B(n4048), .ZN(n4051)
         );
  AOI21_X1 U4709 ( .B1(n4052), .B2(n4490), .A(n4051), .ZN(n4053) );
  OAI211_X1 U4710 ( .C1(n4367), .C2(n4236), .A(n4054), .B(n4053), .ZN(U3265)
         );
  XOR2_X1 U4711 ( .A(n4060), .B(n4055), .Z(n4056) );
  NAND2_X1 U4712 ( .A1(n4056), .A2(n4203), .ZN(n4245) );
  NAND2_X1 U4713 ( .A1(n4058), .A2(n4057), .ZN(n4059) );
  XOR2_X1 U4714 ( .A(n4060), .B(n4059), .Z(n4248) );
  NAND2_X1 U4715 ( .A1(n4248), .A2(n4112), .ZN(n4071) );
  AND2_X1 U4716 ( .A1(n4082), .A2(n4242), .ZN(n4062) );
  OR2_X1 U4717 ( .A1(n4062), .A2(n4061), .ZN(n4330) );
  INV_X1 U4718 ( .A(n4330), .ZN(n4069) );
  AOI22_X1 U4719 ( .A1(n4063), .A2(n4196), .B1(n4197), .B2(n4242), .ZN(n4066)
         );
  AOI22_X1 U4720 ( .A1(n4064), .A2(n4486), .B1(REG2_REG_24__SCAN_IN), .B2(
        n4367), .ZN(n4065) );
  OAI211_X1 U4721 ( .C1(n4067), .C2(n4202), .A(n4066), .B(n4065), .ZN(n4068)
         );
  AOI21_X1 U4722 ( .B1(n4069), .B2(n4490), .A(n4068), .ZN(n4070) );
  OAI211_X1 U4723 ( .C1(n4367), .C2(n4245), .A(n4071), .B(n4070), .ZN(U3266)
         );
  XOR2_X1 U4724 ( .A(n4077), .B(n4072), .Z(n4252) );
  INV_X1 U4725 ( .A(n4252), .ZN(n4090) );
  INV_X1 U4726 ( .A(n4073), .ZN(n4075) );
  AOI21_X1 U4727 ( .B1(n4108), .B2(n4075), .A(n4074), .ZN(n4091) );
  OAI21_X1 U4728 ( .B1(n4091), .B2(n4100), .A(n4076), .ZN(n4078) );
  XNOR2_X1 U4729 ( .A(n4078), .B(n4077), .ZN(n4081) );
  OAI22_X1 U4730 ( .A1(n4265), .A2(n4299), .B1(n4220), .B2(n4083), .ZN(n4079)
         );
  AOI21_X1 U4731 ( .B1(n4234), .B2(n4283), .A(n4079), .ZN(n4080) );
  OAI21_X1 U4732 ( .B1(n4081), .B2(n4159), .A(n4080), .ZN(n4251) );
  INV_X1 U4733 ( .A(n4097), .ZN(n4084) );
  OAI21_X1 U4734 ( .B1(n4084), .B2(n4083), .A(n4082), .ZN(n4334) );
  INV_X1 U4735 ( .A(n4085), .ZN(n4086) );
  AOI22_X1 U4736 ( .A1(n4086), .A2(n4486), .B1(n4367), .B2(
        REG2_REG_23__SCAN_IN), .ZN(n4087) );
  OAI21_X1 U4737 ( .B1(n4334), .B2(n4164), .A(n4087), .ZN(n4088) );
  AOI21_X1 U4738 ( .B1(n4251), .B2(n4187), .A(n4088), .ZN(n4089) );
  OAI21_X1 U4739 ( .B1(n4090), .B2(n4210), .A(n4089), .ZN(U3267) );
  XOR2_X1 U4740 ( .A(n4100), .B(n4091), .Z(n4094) );
  OAI22_X1 U4741 ( .A1(n4133), .A2(n4299), .B1(n4095), .B2(n4220), .ZN(n4092)
         );
  AOI21_X1 U4742 ( .B1(n4243), .B2(n4283), .A(n4092), .ZN(n4093) );
  OAI21_X1 U4743 ( .B1(n4094), .B2(n4159), .A(n4093), .ZN(n4256) );
  OR2_X1 U4744 ( .A1(n4113), .A2(n4095), .ZN(n4096) );
  NAND2_X1 U4745 ( .A1(n4097), .A2(n4096), .ZN(n4338) );
  AOI22_X1 U4746 ( .A1(n4367), .A2(REG2_REG_22__SCAN_IN), .B1(n4098), .B2(
        n4486), .ZN(n4099) );
  OAI21_X1 U4747 ( .B1(n4338), .B2(n4164), .A(n4099), .ZN(n4105) );
  NOR2_X1 U4748 ( .A1(n4101), .A2(n4100), .ZN(n4255) );
  INV_X1 U4749 ( .A(n4102), .ZN(n4103) );
  NOR3_X1 U4750 ( .A1(n4255), .A2(n4103), .A3(n4210), .ZN(n4104) );
  AOI211_X1 U4751 ( .C1(n4106), .C2(n4256), .A(n4105), .B(n4104), .ZN(n4107)
         );
  INV_X1 U4752 ( .A(n4107), .ZN(U3268) );
  XNOR2_X1 U4753 ( .A(n4108), .B(n4111), .ZN(n4109) );
  NAND2_X1 U4754 ( .A1(n4109), .A2(n4203), .ZN(n4264) );
  XOR2_X1 U4755 ( .A(n4111), .B(n4110), .Z(n4267) );
  NAND2_X1 U4756 ( .A1(n4267), .A2(n4112), .ZN(n4124) );
  INV_X1 U4757 ( .A(n4113), .ZN(n4114) );
  OAI21_X1 U4758 ( .B1(n4138), .B2(n4115), .A(n4114), .ZN(n4342) );
  INV_X1 U4759 ( .A(n4342), .ZN(n4122) );
  AOI22_X1 U4760 ( .A1(n4116), .A2(n4196), .B1(n4197), .B2(n4260), .ZN(n4119)
         );
  AOI22_X1 U4761 ( .A1(n4367), .A2(REG2_REG_21__SCAN_IN), .B1(n4117), .B2(
        n4486), .ZN(n4118) );
  OAI211_X1 U4762 ( .C1(n4120), .C2(n4202), .A(n4119), .B(n4118), .ZN(n4121)
         );
  AOI21_X1 U4763 ( .B1(n4122), .B2(n4490), .A(n4121), .ZN(n4123) );
  OAI211_X1 U4764 ( .C1(n4367), .C2(n4264), .A(n4124), .B(n4123), .ZN(U3269)
         );
  XOR2_X1 U4765 ( .A(n4129), .B(n4125), .Z(n4270) );
  INV_X1 U4766 ( .A(n4126), .ZN(n4127) );
  NAND2_X1 U4767 ( .A1(n4128), .A2(n4127), .ZN(n4130) );
  XNOR2_X1 U4768 ( .A(n4130), .B(n4129), .ZN(n4135) );
  AOI22_X1 U4769 ( .A1(n4176), .A2(n4261), .B1(n4131), .B2(n4295), .ZN(n4132)
         );
  OAI21_X1 U4770 ( .B1(n4133), .B2(n4293), .A(n4132), .ZN(n4134) );
  AOI21_X1 U4771 ( .B1(n4135), .B2(n4203), .A(n4134), .ZN(n4136) );
  OAI21_X1 U4772 ( .B1(n4270), .B2(n4137), .A(n4136), .ZN(n4271) );
  NAND2_X1 U4773 ( .A1(n4271), .A2(n4187), .ZN(n4146) );
  INV_X1 U4774 ( .A(n4138), .ZN(n4139) );
  OAI21_X1 U4775 ( .B1(n2079), .B2(n4140), .A(n4139), .ZN(n4346) );
  INV_X1 U4776 ( .A(n4346), .ZN(n4144) );
  INV_X1 U4777 ( .A(REG2_REG_20__SCAN_IN), .ZN(n4142) );
  OAI22_X1 U4778 ( .A1(n4106), .A2(n4142), .B1(n4141), .B2(n4476), .ZN(n4143)
         );
  AOI21_X1 U4779 ( .B1(n4144), .B2(n4490), .A(n4143), .ZN(n4145) );
  OAI211_X1 U4780 ( .C1(n4270), .C2(n4147), .A(n4146), .B(n4145), .ZN(U3270)
         );
  XNOR2_X1 U4781 ( .A(n4148), .B(n4155), .ZN(n4276) );
  INV_X1 U4782 ( .A(n4276), .ZN(n4169) );
  NAND2_X1 U4783 ( .A1(n4150), .A2(n4149), .ZN(n4173) );
  INV_X1 U4784 ( .A(n4151), .ZN(n4153) );
  OAI21_X1 U4785 ( .B1(n4173), .B2(n4153), .A(n4152), .ZN(n4154) );
  XOR2_X1 U4786 ( .A(n4155), .B(n4154), .Z(n4160) );
  OAI22_X1 U4787 ( .A1(n4156), .A2(n4299), .B1(n4220), .B2(n4162), .ZN(n4157)
         );
  AOI21_X1 U4788 ( .B1(n4262), .B2(n4283), .A(n4157), .ZN(n4158) );
  OAI21_X1 U4789 ( .B1(n4160), .B2(n4159), .A(n4158), .ZN(n4275) );
  INV_X1 U4790 ( .A(n4180), .ZN(n4163) );
  OAI21_X1 U4791 ( .B1(n4163), .B2(n4162), .A(n4161), .ZN(n4350) );
  NOR2_X1 U4792 ( .A1(n4350), .A2(n4164), .ZN(n4167) );
  OAI22_X1 U4793 ( .A1(n4187), .A2(n3938), .B1(n4165), .B2(n4476), .ZN(n4166)
         );
  AOI211_X1 U4794 ( .C1(n4275), .C2(n4187), .A(n4167), .B(n4166), .ZN(n4168)
         );
  OAI21_X1 U4795 ( .B1(n4169), .B2(n4210), .A(n4168), .ZN(U3271) );
  OAI21_X1 U4796 ( .B1(n4171), .B2(n4174), .A(n4170), .ZN(n4172) );
  INV_X1 U4797 ( .A(n4172), .ZN(n4281) );
  XOR2_X1 U4798 ( .A(n4174), .B(n4173), .Z(n4179) );
  AOI22_X1 U4799 ( .A1(n4176), .A2(n4283), .B1(n4175), .B2(n4295), .ZN(n4177)
         );
  OAI21_X1 U4800 ( .B1(n4294), .B2(n4299), .A(n4177), .ZN(n4178) );
  AOI21_X1 U4801 ( .B1(n4179), .B2(n4203), .A(n4178), .ZN(n4280) );
  INV_X1 U4802 ( .A(n4280), .ZN(n4188) );
  OAI211_X1 U4803 ( .C1(n4182), .C2(n4181), .A(n4180), .B(n4302), .ZN(n4279)
         );
  NOR2_X1 U4804 ( .A1(n4279), .A2(n4183), .ZN(n4186) );
  OAI22_X1 U4805 ( .A1(n4106), .A2(n3939), .B1(n4184), .B2(n4476), .ZN(n4185)
         );
  AOI211_X1 U4806 ( .C1(n4188), .C2(n4187), .A(n4186), .B(n4185), .ZN(n4189)
         );
  OAI21_X1 U4807 ( .B1(n4281), .B2(n4210), .A(n4189), .ZN(U3272) );
  AOI21_X1 U4808 ( .B1(n4205), .B2(n4191), .A(n4190), .ZN(n4192) );
  INV_X1 U4809 ( .A(n4192), .ZN(n4307) );
  NAND2_X1 U4810 ( .A1(n2051), .A2(n4296), .ZN(n4193) );
  AND2_X1 U4811 ( .A1(n4194), .A2(n4193), .ZN(n4303) );
  AOI22_X1 U4812 ( .A1(n4197), .A2(n4296), .B1(n4196), .B2(n4195), .ZN(n4201)
         );
  INV_X1 U4813 ( .A(n4198), .ZN(n4199) );
  AOI22_X1 U4814 ( .A1(n4367), .A2(REG2_REG_16__SCAN_IN), .B1(n4199), .B2(
        n4486), .ZN(n4200) );
  OAI211_X1 U4815 ( .C1(n4300), .C2(n4202), .A(n4201), .B(n4200), .ZN(n4208)
         );
  OAI211_X1 U4816 ( .C1(n4206), .C2(n4205), .A(n4204), .B(n4203), .ZN(n4304)
         );
  NOR2_X1 U4817 ( .A1(n4304), .A2(n4367), .ZN(n4207) );
  AOI211_X1 U4818 ( .C1(n4303), .C2(n4490), .A(n4208), .B(n4207), .ZN(n4209)
         );
  OAI21_X1 U4819 ( .B1(n4307), .B2(n4210), .A(n4209), .ZN(U3274) );
  NOR2_X1 U4820 ( .A1(n4535), .A2(n4211), .ZN(n4212) );
  AOI21_X1 U4821 ( .B1(n4535), .B2(n4308), .A(n4212), .ZN(n4213) );
  OAI21_X1 U4822 ( .B1(n4311), .B2(n4292), .A(n4213), .ZN(U3549) );
  AOI21_X1 U4823 ( .B1(n4218), .B2(n4215), .A(n4214), .ZN(n4368) );
  INV_X1 U4824 ( .A(n4368), .ZN(n4314) );
  INV_X1 U4825 ( .A(n4216), .ZN(n4217) );
  AOI21_X1 U4826 ( .B1(n4218), .B2(n4295), .A(n4217), .ZN(n4370) );
  MUX2_X1 U4827 ( .A(n4370), .B(n2714), .S(n4533), .Z(n4219) );
  OAI21_X1 U4828 ( .B1(n4314), .B2(n4292), .A(n4219), .ZN(U3548) );
  OAI22_X1 U4829 ( .A1(n4237), .A2(n4299), .B1(n4221), .B2(n4220), .ZN(n4223)
         );
  AOI211_X1 U4830 ( .C1(n4283), .C2(n4224), .A(n4223), .B(n4222), .ZN(n4225)
         );
  OAI21_X1 U4831 ( .B1(n4226), .B2(n4306), .A(n4225), .ZN(n4315) );
  MUX2_X1 U4832 ( .A(REG1_REG_27__SCAN_IN), .B(n4315), .S(n4535), .Z(n4227) );
  INV_X1 U4833 ( .A(n4227), .ZN(n4228) );
  OAI21_X1 U4834 ( .B1(n4292), .B2(n4318), .A(n4228), .ZN(U3545) );
  AOI21_X1 U4835 ( .B1(n4230), .B2(n4521), .A(n4229), .ZN(n4319) );
  MUX2_X1 U4836 ( .A(n4231), .B(n4319), .S(n4535), .Z(n4232) );
  OAI21_X1 U4837 ( .B1(n4292), .B2(n4322), .A(n4232), .ZN(U3544) );
  AOI22_X1 U4838 ( .A1(n4234), .A2(n4261), .B1(n4233), .B2(n4295), .ZN(n4235)
         );
  OAI211_X1 U4839 ( .C1(n4237), .C2(n4293), .A(n4236), .B(n4235), .ZN(n4238)
         );
  AOI21_X1 U4840 ( .B1(n4239), .B2(n4521), .A(n4238), .ZN(n4323) );
  MUX2_X1 U4841 ( .A(n4240), .B(n4323), .S(n4535), .Z(n4241) );
  OAI21_X1 U4842 ( .B1(n4292), .B2(n4326), .A(n4241), .ZN(U3543) );
  AOI22_X1 U4843 ( .A1(n4243), .A2(n4261), .B1(n4295), .B2(n4242), .ZN(n4244)
         );
  OAI211_X1 U4844 ( .C1(n4246), .C2(n4293), .A(n4245), .B(n4244), .ZN(n4247)
         );
  AOI21_X1 U4845 ( .B1(n4248), .B2(n4521), .A(n4247), .ZN(n4327) );
  MUX2_X1 U4846 ( .A(n4249), .B(n4327), .S(n4535), .Z(n4250) );
  OAI21_X1 U4847 ( .B1(n4292), .B2(n4330), .A(n4250), .ZN(U3542) );
  AOI21_X1 U4848 ( .B1(n4252), .B2(n4521), .A(n4251), .ZN(n4331) );
  MUX2_X1 U4849 ( .A(n4253), .B(n4331), .S(n4535), .Z(n4254) );
  OAI21_X1 U4850 ( .B1(n4292), .B2(n4334), .A(n4254), .ZN(U3541) );
  NOR2_X1 U4851 ( .A1(n4255), .A2(n4306), .ZN(n4257) );
  AOI21_X1 U4852 ( .B1(n4257), .B2(n4102), .A(n4256), .ZN(n4335) );
  MUX2_X1 U4853 ( .A(n4258), .B(n4335), .S(n4535), .Z(n4259) );
  OAI21_X1 U4854 ( .B1(n4292), .B2(n4338), .A(n4259), .ZN(U3540) );
  AOI22_X1 U4855 ( .A1(n4262), .A2(n4261), .B1(n4260), .B2(n4295), .ZN(n4263)
         );
  OAI211_X1 U4856 ( .C1(n4265), .C2(n4293), .A(n4264), .B(n4263), .ZN(n4266)
         );
  AOI21_X1 U4857 ( .B1(n4267), .B2(n4521), .A(n4266), .ZN(n4339) );
  MUX2_X1 U4858 ( .A(n4268), .B(n4339), .S(n4535), .Z(n4269) );
  OAI21_X1 U4859 ( .B1(n4292), .B2(n4342), .A(n4269), .ZN(U3539) );
  INV_X1 U4860 ( .A(n4270), .ZN(n4272) );
  AOI21_X1 U4861 ( .B1(n4519), .B2(n4272), .A(n4271), .ZN(n4343) );
  MUX2_X1 U4862 ( .A(n4273), .B(n4343), .S(n4535), .Z(n4274) );
  OAI21_X1 U4863 ( .B1(n4292), .B2(n4346), .A(n4274), .ZN(U3538) );
  AOI21_X1 U4864 ( .B1(n4276), .B2(n4521), .A(n4275), .ZN(n4347) );
  MUX2_X1 U4865 ( .A(n4277), .B(n4347), .S(n4535), .Z(n4278) );
  OAI21_X1 U4866 ( .B1(n4292), .B2(n4350), .A(n4278), .ZN(U3537) );
  OAI211_X1 U4867 ( .C1(n4281), .C2(n4306), .A(n4280), .B(n4279), .ZN(n4351)
         );
  MUX2_X1 U4868 ( .A(REG1_REG_18__SCAN_IN), .B(n4351), .S(n4535), .Z(U3536) );
  AOI22_X1 U4869 ( .A1(n4284), .A2(n4283), .B1(n4295), .B2(n4282), .ZN(n4285)
         );
  OAI211_X1 U4870 ( .C1(n4287), .C2(n4299), .A(n4286), .B(n4285), .ZN(n4288)
         );
  AOI21_X1 U4871 ( .B1(n4289), .B2(n4521), .A(n4288), .ZN(n4352) );
  MUX2_X1 U4872 ( .A(n4290), .B(n4352), .S(n4535), .Z(n4291) );
  OAI21_X1 U4873 ( .B1(n4292), .B2(n4356), .A(n4291), .ZN(U3535) );
  OR2_X1 U4874 ( .A1(n4294), .A2(n4293), .ZN(n4298) );
  NAND2_X1 U4875 ( .A1(n4296), .A2(n4295), .ZN(n4297) );
  OAI211_X1 U4876 ( .C1(n4300), .C2(n4299), .A(n4298), .B(n4297), .ZN(n4301)
         );
  AOI21_X1 U4877 ( .B1(n4303), .B2(n4302), .A(n4301), .ZN(n4305) );
  OAI211_X1 U4878 ( .C1(n4307), .C2(n4306), .A(n4305), .B(n4304), .ZN(n4357)
         );
  MUX2_X1 U4879 ( .A(REG1_REG_16__SCAN_IN), .B(n4357), .S(n4535), .Z(U3534) );
  NAND2_X1 U4880 ( .A1(n4529), .A2(n4308), .ZN(n4310) );
  NAND2_X1 U4881 ( .A1(n4527), .A2(REG0_REG_31__SCAN_IN), .ZN(n4309) );
  OAI211_X1 U4882 ( .C1(n4311), .C2(n4355), .A(n4310), .B(n4309), .ZN(U3517)
         );
  INV_X1 U4883 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4312) );
  MUX2_X1 U4884 ( .A(n4370), .B(n4312), .S(n4527), .Z(n4313) );
  OAI21_X1 U4885 ( .B1(n4314), .B2(n4355), .A(n4313), .ZN(U3516) );
  MUX2_X1 U4886 ( .A(REG0_REG_27__SCAN_IN), .B(n4315), .S(n4529), .Z(n4316) );
  INV_X1 U4887 ( .A(n4316), .ZN(n4317) );
  OAI21_X1 U4888 ( .B1(n4318), .B2(n4355), .A(n4317), .ZN(U3513) );
  INV_X1 U4889 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4320) );
  MUX2_X1 U4890 ( .A(n4320), .B(n4319), .S(n4529), .Z(n4321) );
  OAI21_X1 U4891 ( .B1(n4322), .B2(n4355), .A(n4321), .ZN(U3512) );
  INV_X1 U4892 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4324) );
  MUX2_X1 U4893 ( .A(n4324), .B(n4323), .S(n4529), .Z(n4325) );
  OAI21_X1 U4894 ( .B1(n4326), .B2(n4355), .A(n4325), .ZN(U3511) );
  INV_X1 U4895 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4328) );
  MUX2_X1 U4896 ( .A(n4328), .B(n4327), .S(n4529), .Z(n4329) );
  OAI21_X1 U4897 ( .B1(n4330), .B2(n4355), .A(n4329), .ZN(U3510) );
  INV_X1 U4898 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4332) );
  MUX2_X1 U4899 ( .A(n4332), .B(n4331), .S(n4529), .Z(n4333) );
  OAI21_X1 U4900 ( .B1(n4334), .B2(n4355), .A(n4333), .ZN(U3509) );
  INV_X1 U4901 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4336) );
  MUX2_X1 U4902 ( .A(n4336), .B(n4335), .S(n4529), .Z(n4337) );
  OAI21_X1 U4903 ( .B1(n4338), .B2(n4355), .A(n4337), .ZN(U3508) );
  INV_X1 U4904 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4340) );
  MUX2_X1 U4905 ( .A(n4340), .B(n4339), .S(n4529), .Z(n4341) );
  OAI21_X1 U4906 ( .B1(n4342), .B2(n4355), .A(n4341), .ZN(U3507) );
  INV_X1 U4907 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4344) );
  MUX2_X1 U4908 ( .A(n4344), .B(n4343), .S(n4529), .Z(n4345) );
  OAI21_X1 U4909 ( .B1(n4346), .B2(n4355), .A(n4345), .ZN(U3506) );
  INV_X1 U4910 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4348) );
  MUX2_X1 U4911 ( .A(n4348), .B(n4347), .S(n4529), .Z(n4349) );
  OAI21_X1 U4912 ( .B1(n4350), .B2(n4355), .A(n4349), .ZN(U3505) );
  MUX2_X1 U4913 ( .A(REG0_REG_18__SCAN_IN), .B(n4351), .S(n4529), .Z(U3503) );
  MUX2_X1 U4914 ( .A(n4353), .B(n4352), .S(n4529), .Z(n4354) );
  OAI21_X1 U4915 ( .B1(n4356), .B2(n4355), .A(n4354), .ZN(U3501) );
  MUX2_X1 U4916 ( .A(REG0_REG_16__SCAN_IN), .B(n4357), .S(n4529), .Z(U3499) );
  MUX2_X1 U4917 ( .A(DATAI_30_), .B(n4358), .S(STATE_REG_SCAN_IN), .Z(U3322)
         );
  MUX2_X1 U4918 ( .A(DATAI_21_), .B(n4359), .S(STATE_REG_SCAN_IN), .Z(U3331)
         );
  MUX2_X1 U4919 ( .A(DATAI_20_), .B(n2651), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U4920 ( .A(n4360), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4921 ( .A(DATAI_8_), .B(n2091), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U4922 ( .A(n4362), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U4923 ( .A(n4363), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U4924 ( .A(n2105), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U4925 ( .A(DATAI_4_), .B(n4364), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4926 ( .A(n4365), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4927 ( .A(n4366), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  AOI22_X1 U4928 ( .A1(n4368), .A2(n4490), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4367), .ZN(n4369) );
  OAI211_X1 U4929 ( .C1(n4373), .C2(n4372), .A(n4470), .B(n4371), .ZN(n4378)
         );
  OAI211_X1 U4930 ( .C1(n4376), .C2(n4375), .A(n4413), .B(n4374), .ZN(n4377)
         );
  OAI211_X1 U4931 ( .C1(n4475), .C2(n4510), .A(n4378), .B(n4377), .ZN(n4379)
         );
  AOI211_X1 U4932 ( .C1(n4468), .C2(ADDR_REG_9__SCAN_IN), .A(n4380), .B(n4379), 
        .ZN(n4381) );
  INV_X1 U4933 ( .A(n4381), .ZN(U3249) );
  OAI211_X1 U4934 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4383), .A(n4413), .B(n4382), .ZN(n4385) );
  NAND2_X1 U4935 ( .A1(n4385), .A2(n4384), .ZN(n4386) );
  AOI21_X1 U4936 ( .B1(n4468), .B2(ADDR_REG_10__SCAN_IN), .A(n4386), .ZN(n4390) );
  OAI211_X1 U4937 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4388), .A(n4470), .B(n4387), .ZN(n4389) );
  OAI211_X1 U4938 ( .C1(n4475), .C2(n4508), .A(n4390), .B(n4389), .ZN(U3250)
         );
  OAI211_X1 U4939 ( .C1(n4393), .C2(n4392), .A(n4470), .B(n4391), .ZN(n4398)
         );
  OAI211_X1 U4940 ( .C1(n4396), .C2(n4395), .A(n4413), .B(n4394), .ZN(n4397)
         );
  OAI211_X1 U4941 ( .C1(n4475), .C2(n4507), .A(n4398), .B(n4397), .ZN(n4399)
         );
  AOI211_X1 U4942 ( .C1(n4468), .C2(ADDR_REG_11__SCAN_IN), .A(n4400), .B(n4399), .ZN(n4401) );
  INV_X1 U4943 ( .A(n4401), .ZN(U3251) );
  OAI211_X1 U4944 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4403), .A(n4413), .B(n4402), .ZN(n4405) );
  NAND2_X1 U4945 ( .A1(n4405), .A2(n4404), .ZN(n4406) );
  AOI21_X1 U4946 ( .B1(n4468), .B2(ADDR_REG_12__SCAN_IN), .A(n4406), .ZN(n4410) );
  OAI211_X1 U4947 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4408), .A(n4470), .B(n4407), .ZN(n4409) );
  OAI211_X1 U4948 ( .C1(n4475), .C2(n4506), .A(n4410), .B(n4409), .ZN(U3252)
         );
  AOI21_X1 U4949 ( .B1(n4412), .B2(n4505), .A(n4411), .ZN(n4416) );
  OAI21_X1 U4950 ( .B1(n4416), .B2(n4415), .A(n4413), .ZN(n4414) );
  AOI21_X1 U4951 ( .B1(n4416), .B2(n4415), .A(n4414), .ZN(n4418) );
  AOI211_X1 U4952 ( .C1(n4468), .C2(ADDR_REG_13__SCAN_IN), .A(n4418), .B(n4417), .ZN(n4423) );
  OAI211_X1 U4953 ( .C1(n4421), .C2(n4420), .A(n4470), .B(n4419), .ZN(n4422)
         );
  OAI211_X1 U4954 ( .C1(n4475), .C2(n4505), .A(n4423), .B(n4422), .ZN(U3253)
         );
  AOI211_X1 U4955 ( .C1(n2466), .C2(n4425), .A(n4424), .B(n4464), .ZN(n4426)
         );
  AOI211_X1 U4956 ( .C1(n4468), .C2(ADDR_REG_14__SCAN_IN), .A(n4427), .B(n4426), .ZN(n4431) );
  OAI211_X1 U4957 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4429), .A(n4470), .B(n4428), .ZN(n4430) );
  OAI211_X1 U4958 ( .C1(n4475), .C2(n4432), .A(n4431), .B(n4430), .ZN(U3254)
         );
  AOI211_X1 U4959 ( .C1(n4435), .C2(n4434), .A(n4433), .B(n4464), .ZN(n4436)
         );
  AOI211_X1 U4960 ( .C1(n4468), .C2(ADDR_REG_15__SCAN_IN), .A(n4437), .B(n4436), .ZN(n4442) );
  OAI211_X1 U4961 ( .C1(n4440), .C2(n4439), .A(n4470), .B(n4438), .ZN(n4441)
         );
  OAI211_X1 U4962 ( .C1(n4475), .C2(n4502), .A(n4442), .B(n4441), .ZN(U3255)
         );
  INV_X1 U4963 ( .A(n4443), .ZN(n4448) );
  AOI221_X1 U4964 ( .B1(n4446), .B2(n4445), .C1(n4444), .C2(n4445), .A(n4464), 
        .ZN(n4447) );
  AOI211_X1 U4965 ( .C1(n4468), .C2(ADDR_REG_16__SCAN_IN), .A(n4448), .B(n4447), .ZN(n4452) );
  OAI221_X1 U4966 ( .B1(n4450), .B2(REG1_REG_16__SCAN_IN), .C1(n4450), .C2(
        n4449), .A(n4470), .ZN(n4451) );
  OAI211_X1 U4967 ( .C1(n4475), .C2(n4501), .A(n4452), .B(n4451), .ZN(U3256)
         );
  AOI221_X1 U4968 ( .B1(n4455), .B2(n4454), .C1(n4453), .C2(n4454), .A(n4464), 
        .ZN(n4456) );
  AOI211_X1 U4969 ( .C1(n4468), .C2(ADDR_REG_17__SCAN_IN), .A(n4457), .B(n4456), .ZN(n4462) );
  OAI221_X1 U4970 ( .B1(n4460), .B2(n4459), .C1(n4460), .C2(n4458), .A(n4470), 
        .ZN(n4461) );
  OAI211_X1 U4971 ( .C1(n4475), .C2(n4463), .A(n4462), .B(n4461), .ZN(U3257)
         );
  OAI211_X1 U4972 ( .C1(n4472), .C2(n4471), .A(n4470), .B(n4469), .ZN(n4473)
         );
  OAI211_X1 U4973 ( .C1(n4475), .C2(n4498), .A(n4474), .B(n4473), .ZN(U3258)
         );
  OAI22_X1 U4974 ( .A1(n4106), .A2(n4478), .B1(n4477), .B2(n4476), .ZN(n4479)
         );
  INV_X1 U4975 ( .A(n4479), .ZN(n4484) );
  INV_X1 U4976 ( .A(n4480), .ZN(n4482) );
  AOI22_X1 U4977 ( .A1(n4482), .A2(n4491), .B1(n4490), .B2(n4481), .ZN(n4483)
         );
  OAI211_X1 U4978 ( .C1(n4367), .C2(n4485), .A(n4484), .B(n4483), .ZN(U3282)
         );
  AOI22_X1 U4979 ( .A1(n4367), .A2(REG2_REG_3__SCAN_IN), .B1(n4486), .B2(n4680), .ZN(n4494) );
  INV_X1 U4980 ( .A(n4487), .ZN(n4492) );
  INV_X1 U4981 ( .A(n4488), .ZN(n4489) );
  AOI22_X1 U4982 ( .A1(n4492), .A2(n4491), .B1(n4490), .B2(n4489), .ZN(n4493)
         );
  OAI211_X1 U4983 ( .C1(n4367), .C2(n4495), .A(n4494), .B(n4493), .ZN(U3287)
         );
  AND2_X1 U4984 ( .A1(D_REG_31__SCAN_IN), .A2(n4496), .ZN(U3291) );
  AND2_X1 U4985 ( .A1(D_REG_30__SCAN_IN), .A2(n4496), .ZN(U3292) );
  AND2_X1 U4986 ( .A1(D_REG_29__SCAN_IN), .A2(n4496), .ZN(U3293) );
  AND2_X1 U4987 ( .A1(D_REG_28__SCAN_IN), .A2(n4496), .ZN(U3294) );
  AND2_X1 U4988 ( .A1(D_REG_27__SCAN_IN), .A2(n4496), .ZN(U3295) );
  AND2_X1 U4989 ( .A1(D_REG_26__SCAN_IN), .A2(n4496), .ZN(U3296) );
  AND2_X1 U4990 ( .A1(D_REG_25__SCAN_IN), .A2(n4496), .ZN(U3297) );
  AND2_X1 U4991 ( .A1(D_REG_24__SCAN_IN), .A2(n4496), .ZN(U3298) );
  AND2_X1 U4992 ( .A1(D_REG_23__SCAN_IN), .A2(n4496), .ZN(U3299) );
  AND2_X1 U4993 ( .A1(D_REG_22__SCAN_IN), .A2(n4496), .ZN(U3300) );
  AND2_X1 U4994 ( .A1(D_REG_21__SCAN_IN), .A2(n4496), .ZN(U3301) );
  AND2_X1 U4995 ( .A1(D_REG_20__SCAN_IN), .A2(n4496), .ZN(U3302) );
  AND2_X1 U4996 ( .A1(D_REG_19__SCAN_IN), .A2(n4496), .ZN(U3303) );
  AND2_X1 U4997 ( .A1(D_REG_18__SCAN_IN), .A2(n4496), .ZN(U3304) );
  AND2_X1 U4998 ( .A1(D_REG_17__SCAN_IN), .A2(n4496), .ZN(U3305) );
  AND2_X1 U4999 ( .A1(D_REG_16__SCAN_IN), .A2(n4496), .ZN(U3306) );
  AND2_X1 U5000 ( .A1(D_REG_15__SCAN_IN), .A2(n4496), .ZN(U3307) );
  AND2_X1 U5001 ( .A1(D_REG_14__SCAN_IN), .A2(n4496), .ZN(U3308) );
  AND2_X1 U5002 ( .A1(D_REG_13__SCAN_IN), .A2(n4496), .ZN(U3309) );
  AND2_X1 U5003 ( .A1(D_REG_12__SCAN_IN), .A2(n4496), .ZN(U3310) );
  AND2_X1 U5004 ( .A1(D_REG_11__SCAN_IN), .A2(n4496), .ZN(U3311) );
  AND2_X1 U5005 ( .A1(D_REG_10__SCAN_IN), .A2(n4496), .ZN(U3312) );
  AND2_X1 U5006 ( .A1(D_REG_9__SCAN_IN), .A2(n4496), .ZN(U3313) );
  AND2_X1 U5007 ( .A1(D_REG_8__SCAN_IN), .A2(n4496), .ZN(U3314) );
  AND2_X1 U5008 ( .A1(D_REG_7__SCAN_IN), .A2(n4496), .ZN(U3315) );
  AND2_X1 U5009 ( .A1(D_REG_6__SCAN_IN), .A2(n4496), .ZN(U3316) );
  AND2_X1 U5010 ( .A1(D_REG_5__SCAN_IN), .A2(n4496), .ZN(U3317) );
  AND2_X1 U5011 ( .A1(D_REG_4__SCAN_IN), .A2(n4496), .ZN(U3318) );
  AND2_X1 U5012 ( .A1(D_REG_3__SCAN_IN), .A2(n4496), .ZN(U3319) );
  AND2_X1 U5013 ( .A1(D_REG_2__SCAN_IN), .A2(n4496), .ZN(U3320) );
  AOI21_X1 U5014 ( .B1(U3149), .B2(n2547), .A(n4497), .ZN(U3329) );
  INV_X1 U5015 ( .A(DATAI_18_), .ZN(n4625) );
  AOI22_X1 U5016 ( .A1(STATE_REG_SCAN_IN), .A2(n4498), .B1(n4625), .B2(U3149), 
        .ZN(U3334) );
  OAI22_X1 U5017 ( .A1(U3149), .A2(n4499), .B1(DATAI_17_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4500) );
  INV_X1 U5018 ( .A(n4500), .ZN(U3335) );
  INV_X1 U5019 ( .A(DATAI_16_), .ZN(n4689) );
  AOI22_X1 U5020 ( .A1(STATE_REG_SCAN_IN), .A2(n4501), .B1(n4689), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U5021 ( .A1(STATE_REG_SCAN_IN), .A2(n4502), .B1(n4681), .B2(U3149), 
        .ZN(U3337) );
  OAI22_X1 U5022 ( .A1(U3149), .A2(n4503), .B1(DATAI_14_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4504) );
  INV_X1 U5023 ( .A(n4504), .ZN(U3338) );
  AOI22_X1 U5024 ( .A1(STATE_REG_SCAN_IN), .A2(n4505), .B1(n2461), .B2(U3149), 
        .ZN(U3339) );
  INV_X1 U5025 ( .A(DATAI_12_), .ZN(n4657) );
  AOI22_X1 U5026 ( .A1(STATE_REG_SCAN_IN), .A2(n4506), .B1(n4657), .B2(U3149), 
        .ZN(U3340) );
  INV_X1 U5027 ( .A(DATAI_11_), .ZN(n4700) );
  AOI22_X1 U5028 ( .A1(STATE_REG_SCAN_IN), .A2(n4507), .B1(n4700), .B2(U3149), 
        .ZN(U3341) );
  INV_X1 U5029 ( .A(DATAI_10_), .ZN(n4635) );
  AOI22_X1 U5030 ( .A1(STATE_REG_SCAN_IN), .A2(n4508), .B1(n4635), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5031 ( .A(DATAI_9_), .ZN(n4509) );
  AOI22_X1 U5032 ( .A1(STATE_REG_SCAN_IN), .A2(n4510), .B1(n4509), .B2(U3149), 
        .ZN(U3343) );
  INV_X1 U5033 ( .A(n4511), .ZN(n4514) );
  INV_X1 U5034 ( .A(n4512), .ZN(n4513) );
  AOI211_X1 U5035 ( .C1(n4519), .C2(n4515), .A(n4514), .B(n4513), .ZN(n4531)
         );
  AOI22_X1 U5036 ( .A1(n4529), .A2(n4531), .B1(n2302), .B2(n4527), .ZN(U3467)
         );
  INV_X1 U5037 ( .A(n4516), .ZN(n4518) );
  AOI211_X1 U5038 ( .C1(n4520), .C2(n4519), .A(n4518), .B(n4517), .ZN(n4532)
         );
  AOI22_X1 U5039 ( .A1(n4529), .A2(n4532), .B1(n2336), .B2(n4527), .ZN(U3475)
         );
  NAND3_X1 U5040 ( .A1(n4523), .A2(n4522), .A3(n4521), .ZN(n4524) );
  INV_X1 U5041 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4528) );
  AOI22_X1 U5042 ( .A1(n4529), .A2(n4534), .B1(n4528), .B2(n4527), .ZN(U3481)
         );
  AOI22_X1 U5043 ( .A1(n4535), .A2(n4531), .B1(n4530), .B2(n4533), .ZN(U3518)
         );
  AOI22_X1 U5044 ( .A1(n4535), .A2(n4532), .B1(n2337), .B2(n4533), .ZN(U3522)
         );
  AOI22_X1 U5045 ( .A1(n4535), .A2(n4534), .B1(n2400), .B2(n4533), .ZN(U3525)
         );
  AOI22_X1 U5046 ( .A1(STATE_REG_SCAN_IN), .A2(IR_REG_0__SCAN_IN), .B1(
        DATAI_0_), .B2(U3149), .ZN(n4722) );
  AOI22_X1 U5047 ( .A1(n4537), .A2(keyinput_g0), .B1(n4635), .B2(keyinput_g21), 
        .ZN(n4536) );
  OAI221_X1 U5048 ( .B1(n4537), .B2(keyinput_g0), .C1(n4635), .C2(keyinput_g21), .A(n4536), .ZN(n4546) );
  AOI22_X1 U5049 ( .A1(n2608), .A2(keyinput_g3), .B1(keyinput_g18), .B2(n2461), 
        .ZN(n4538) );
  OAI221_X1 U5050 ( .B1(n2608), .B2(keyinput_g3), .C1(n2461), .C2(keyinput_g18), .A(n4538), .ZN(n4545) );
  AOI22_X1 U5051 ( .A1(n4540), .A2(keyinput_g10), .B1(keyinput_g19), .B2(n4657), .ZN(n4539) );
  OAI221_X1 U5052 ( .B1(n4540), .B2(keyinput_g10), .C1(n4657), .C2(
        keyinput_g19), .A(n4539), .ZN(n4544) );
  AOI22_X1 U5053 ( .A1(n4542), .A2(keyinput_g45), .B1(keyinput_g6), .B2(n4658), 
        .ZN(n4541) );
  OAI221_X1 U5054 ( .B1(n4542), .B2(keyinput_g45), .C1(n4658), .C2(keyinput_g6), .A(n4541), .ZN(n4543) );
  NOR4_X1 U5055 ( .A1(n4546), .A2(n4545), .A3(n4544), .A4(n4543), .ZN(n4579)
         );
  AOI22_X1 U5056 ( .A1(n2545), .A2(keyinput_g9), .B1(n4660), .B2(keyinput_g35), 
        .ZN(n4547) );
  OAI221_X1 U5057 ( .B1(n2545), .B2(keyinput_g9), .C1(n4660), .C2(keyinput_g35), .A(n4547), .ZN(n4555) );
  XNOR2_X1 U5058 ( .A(n4669), .B(keyinput_g53), .ZN(n4554) );
  XNOR2_X1 U5059 ( .A(keyinput_g54), .B(n2452), .ZN(n4553) );
  XNOR2_X1 U5060 ( .A(DATAI_1_), .B(keyinput_g30), .ZN(n4551) );
  XNOR2_X1 U5061 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_g57), .ZN(n4550) );
  XNOR2_X1 U5062 ( .A(DATAI_0_), .B(keyinput_g31), .ZN(n4549) );
  XNOR2_X1 U5063 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_g56), .ZN(n4548) );
  NAND4_X1 U5064 ( .A1(n4551), .A2(n4550), .A3(n4549), .A4(n4548), .ZN(n4552)
         );
  NOR4_X1 U5065 ( .A1(n4555), .A2(n4554), .A3(n4553), .A4(n4552), .ZN(n4578)
         );
  INV_X1 U5066 ( .A(DATAI_2_), .ZN(n4557) );
  AOI22_X1 U5067 ( .A1(n4680), .A2(keyinput_g38), .B1(keyinput_g29), .B2(n4557), .ZN(n4556) );
  OAI221_X1 U5068 ( .B1(n4680), .B2(keyinput_g38), .C1(n4557), .C2(
        keyinput_g29), .A(n4556), .ZN(n4565) );
  AOI22_X1 U5069 ( .A1(n2547), .A2(keyinput_g8), .B1(keyinput_g13), .B2(n4625), 
        .ZN(n4558) );
  OAI221_X1 U5070 ( .B1(n2547), .B2(keyinput_g8), .C1(n4625), .C2(keyinput_g13), .A(n4558), .ZN(n4564) );
  XNOR2_X1 U5071 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_g61), .ZN(n4562) );
  XNOR2_X1 U5072 ( .A(REG3_REG_17__SCAN_IN), .B(keyinput_g48), .ZN(n4561) );
  XNOR2_X1 U5073 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_g63), .ZN(n4560) );
  XNOR2_X1 U5074 ( .A(keyinput_g25), .B(DATAI_6_), .ZN(n4559) );
  NAND4_X1 U5075 ( .A1(n4562), .A2(n4561), .A3(n4560), .A4(n4559), .ZN(n4563)
         );
  NOR3_X1 U5076 ( .A1(n4565), .A2(n4564), .A3(n4563), .ZN(n4577) );
  AOI22_X1 U5077 ( .A1(n4700), .A2(keyinput_g20), .B1(n4685), .B2(keyinput_g39), .ZN(n4566) );
  OAI221_X1 U5078 ( .B1(n4700), .B2(keyinput_g20), .C1(n4685), .C2(
        keyinput_g39), .A(n4566), .ZN(n4575) );
  AOI22_X1 U5079 ( .A1(n4636), .A2(keyinput_g7), .B1(n4701), .B2(keyinput_g37), 
        .ZN(n4567) );
  OAI221_X1 U5080 ( .B1(n4636), .B2(keyinput_g7), .C1(n4701), .C2(keyinput_g37), .A(n4567), .ZN(n4574) );
  INV_X1 U5081 ( .A(DATAI_7_), .ZN(n4688) );
  AOI22_X1 U5082 ( .A1(n4688), .A2(keyinput_g24), .B1(n4569), .B2(keyinput_g26), .ZN(n4568) );
  OAI221_X1 U5083 ( .B1(n4688), .B2(keyinput_g24), .C1(n4569), .C2(
        keyinput_g26), .A(n4568), .ZN(n4573) );
  XNOR2_X1 U5084 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_g52), .ZN(n4571) );
  XNOR2_X1 U5085 ( .A(keyinput_g27), .B(DATAI_4_), .ZN(n4570) );
  NAND2_X1 U5086 ( .A1(n4571), .A2(n4570), .ZN(n4572) );
  NOR4_X1 U5087 ( .A1(n4575), .A2(n4574), .A3(n4573), .A4(n4572), .ZN(n4576)
         );
  NAND4_X1 U5088 ( .A1(n4579), .A2(n4578), .A3(n4577), .A4(n4576), .ZN(n4720)
         );
  AOI22_X1 U5089 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput_g42), .B1(DATAI_17_), 
        .B2(keyinput_g14), .ZN(n4580) );
  OAI221_X1 U5090 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput_g42), .C1(DATAI_17_), .C2(keyinput_g14), .A(n4580), .ZN(n4587) );
  AOI22_X1 U5091 ( .A1(DATAI_20_), .A2(keyinput_g11), .B1(DATAI_26_), .B2(
        keyinput_g5), .ZN(n4581) );
  OAI221_X1 U5092 ( .B1(DATAI_20_), .B2(keyinput_g11), .C1(DATAI_26_), .C2(
        keyinput_g5), .A(n4581), .ZN(n4586) );
  AOI22_X1 U5093 ( .A1(REG3_REG_9__SCAN_IN), .A2(keyinput_g51), .B1(
        IR_REG_0__SCAN_IN), .B2(keyinput_g55), .ZN(n4582) );
  OAI221_X1 U5094 ( .B1(REG3_REG_9__SCAN_IN), .B2(keyinput_g51), .C1(
        IR_REG_0__SCAN_IN), .C2(keyinput_g55), .A(n4582), .ZN(n4585) );
  AOI22_X1 U5095 ( .A1(REG3_REG_4__SCAN_IN), .A2(keyinput_g50), .B1(
        REG3_REG_12__SCAN_IN), .B2(keyinput_g44), .ZN(n4583) );
  OAI221_X1 U5096 ( .B1(REG3_REG_4__SCAN_IN), .B2(keyinput_g50), .C1(
        REG3_REG_12__SCAN_IN), .C2(keyinput_g44), .A(n4583), .ZN(n4584) );
  NOR4_X1 U5097 ( .A1(n4587), .A2(n4586), .A3(n4585), .A4(n4584), .ZN(n4614)
         );
  XOR2_X1 U5098 ( .A(U3149), .B(keyinput_g32), .Z(n4594) );
  AOI22_X1 U5099 ( .A1(DATAI_19_), .A2(keyinput_g12), .B1(n4681), .B2(
        keyinput_g16), .ZN(n4588) );
  OAI221_X1 U5100 ( .B1(DATAI_19_), .B2(keyinput_g12), .C1(n4681), .C2(
        keyinput_g16), .A(n4588), .ZN(n4593) );
  AOI22_X1 U5101 ( .A1(DATAI_27_), .A2(keyinput_g4), .B1(REG3_REG_24__SCAN_IN), 
        .B2(keyinput_g49), .ZN(n4589) );
  OAI221_X1 U5102 ( .B1(DATAI_27_), .B2(keyinput_g4), .C1(REG3_REG_24__SCAN_IN), .C2(keyinput_g49), .A(n4589), .ZN(n4592) );
  AOI22_X1 U5103 ( .A1(REG3_REG_23__SCAN_IN), .A2(keyinput_g36), .B1(
        REG3_REG_28__SCAN_IN), .B2(keyinput_g40), .ZN(n4590) );
  OAI221_X1 U5104 ( .B1(REG3_REG_23__SCAN_IN), .B2(keyinput_g36), .C1(
        REG3_REG_28__SCAN_IN), .C2(keyinput_g40), .A(n4590), .ZN(n4591) );
  NOR4_X1 U5105 ( .A1(n4594), .A2(n4593), .A3(n4592), .A4(n4591), .ZN(n4613)
         );
  AOI22_X1 U5106 ( .A1(REG3_REG_16__SCAN_IN), .A2(keyinput_g46), .B1(
        REG3_REG_21__SCAN_IN), .B2(keyinput_g43), .ZN(n4595) );
  OAI221_X1 U5107 ( .B1(REG3_REG_16__SCAN_IN), .B2(keyinput_g46), .C1(
        REG3_REG_21__SCAN_IN), .C2(keyinput_g43), .A(n4595), .ZN(n4602) );
  AOI22_X1 U5108 ( .A1(DATAI_9_), .A2(keyinput_g22), .B1(REG3_REG_27__SCAN_IN), 
        .B2(keyinput_g34), .ZN(n4596) );
  OAI221_X1 U5109 ( .B1(DATAI_9_), .B2(keyinput_g22), .C1(REG3_REG_27__SCAN_IN), .C2(keyinput_g34), .A(n4596), .ZN(n4601) );
  AOI22_X1 U5110 ( .A1(DATAI_29_), .A2(keyinput_g2), .B1(REG3_REG_8__SCAN_IN), 
        .B2(keyinput_g41), .ZN(n4597) );
  OAI221_X1 U5111 ( .B1(DATAI_29_), .B2(keyinput_g2), .C1(REG3_REG_8__SCAN_IN), 
        .C2(keyinput_g41), .A(n4597), .ZN(n4600) );
  AOI22_X1 U5112 ( .A1(DATAI_30_), .A2(keyinput_g1), .B1(DATAI_16_), .B2(
        keyinput_g15), .ZN(n4598) );
  OAI221_X1 U5113 ( .B1(DATAI_30_), .B2(keyinput_g1), .C1(DATAI_16_), .C2(
        keyinput_g15), .A(n4598), .ZN(n4599) );
  NOR4_X1 U5114 ( .A1(n4602), .A2(n4601), .A3(n4600), .A4(n4599), .ZN(n4612)
         );
  AOI22_X1 U5115 ( .A1(REG3_REG_7__SCAN_IN), .A2(keyinput_g33), .B1(
        IR_REG_7__SCAN_IN), .B2(keyinput_g62), .ZN(n4603) );
  OAI221_X1 U5116 ( .B1(REG3_REG_7__SCAN_IN), .B2(keyinput_g33), .C1(
        IR_REG_7__SCAN_IN), .C2(keyinput_g62), .A(n4603), .ZN(n4610) );
  AOI22_X1 U5117 ( .A1(DATAI_8_), .A2(keyinput_g23), .B1(DATAI_14_), .B2(
        keyinput_g17), .ZN(n4604) );
  OAI221_X1 U5118 ( .B1(DATAI_8_), .B2(keyinput_g23), .C1(DATAI_14_), .C2(
        keyinput_g17), .A(n4604), .ZN(n4609) );
  AOI22_X1 U5119 ( .A1(REG3_REG_5__SCAN_IN), .A2(keyinput_g47), .B1(
        IR_REG_5__SCAN_IN), .B2(keyinput_g60), .ZN(n4605) );
  OAI221_X1 U5120 ( .B1(REG3_REG_5__SCAN_IN), .B2(keyinput_g47), .C1(
        IR_REG_5__SCAN_IN), .C2(keyinput_g60), .A(n4605), .ZN(n4608) );
  AOI22_X1 U5121 ( .A1(IR_REG_4__SCAN_IN), .A2(keyinput_g59), .B1(
        IR_REG_3__SCAN_IN), .B2(keyinput_g58), .ZN(n4606) );
  OAI221_X1 U5122 ( .B1(IR_REG_4__SCAN_IN), .B2(keyinput_g59), .C1(
        IR_REG_3__SCAN_IN), .C2(keyinput_g58), .A(n4606), .ZN(n4607) );
  NOR4_X1 U5123 ( .A1(n4610), .A2(n4609), .A3(n4608), .A4(n4607), .ZN(n4611)
         );
  NAND4_X1 U5124 ( .A1(n4614), .A2(n4613), .A3(n4612), .A4(n4611), .ZN(n4719)
         );
  AOI22_X1 U5125 ( .A1(REG3_REG_1__SCAN_IN), .A2(keyinput_f42), .B1(
        REG3_REG_4__SCAN_IN), .B2(keyinput_f50), .ZN(n4615) );
  OAI221_X1 U5126 ( .B1(REG3_REG_1__SCAN_IN), .B2(keyinput_f42), .C1(
        REG3_REG_4__SCAN_IN), .C2(keyinput_f50), .A(n4615), .ZN(n4622) );
  AOI22_X1 U5127 ( .A1(DATAI_17_), .A2(keyinput_f14), .B1(DATAI_20_), .B2(
        keyinput_f11), .ZN(n4616) );
  OAI221_X1 U5128 ( .B1(DATAI_17_), .B2(keyinput_f14), .C1(DATAI_20_), .C2(
        keyinput_f11), .A(n4616), .ZN(n4621) );
  AOI22_X1 U5129 ( .A1(DATAI_8_), .A2(keyinput_f23), .B1(DATAI_14_), .B2(
        keyinput_f17), .ZN(n4617) );
  OAI221_X1 U5130 ( .B1(DATAI_8_), .B2(keyinput_f23), .C1(DATAI_14_), .C2(
        keyinput_f17), .A(n4617), .ZN(n4620) );
  AOI22_X1 U5131 ( .A1(REG3_REG_9__SCAN_IN), .A2(keyinput_f51), .B1(
        REG3_REG_13__SCAN_IN), .B2(keyinput_f54), .ZN(n4618) );
  OAI221_X1 U5132 ( .B1(REG3_REG_9__SCAN_IN), .B2(keyinput_f51), .C1(
        REG3_REG_13__SCAN_IN), .C2(keyinput_f54), .A(n4618), .ZN(n4619) );
  NOR4_X1 U5133 ( .A1(n4622), .A2(n4621), .A3(n4620), .A4(n4619), .ZN(n4653)
         );
  INV_X1 U5134 ( .A(DATAI_19_), .ZN(n4623) );
  XOR2_X1 U5135 ( .A(n4623), .B(keyinput_f12), .Z(n4631) );
  AOI22_X1 U5136 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput_f52), .B1(n4625), 
        .B2(keyinput_f13), .ZN(n4624) );
  OAI221_X1 U5137 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput_f52), .C1(n4625), 
        .C2(keyinput_f13), .A(n4624), .ZN(n4630) );
  AOI22_X1 U5138 ( .A1(DATAI_31_), .A2(keyinput_f0), .B1(DATAI_21_), .B2(
        keyinput_f10), .ZN(n4626) );
  OAI221_X1 U5139 ( .B1(DATAI_31_), .B2(keyinput_f0), .C1(DATAI_21_), .C2(
        keyinput_f10), .A(n4626), .ZN(n4629) );
  AOI22_X1 U5140 ( .A1(REG3_REG_23__SCAN_IN), .A2(keyinput_f36), .B1(
        REG3_REG_28__SCAN_IN), .B2(keyinput_f40), .ZN(n4627) );
  OAI221_X1 U5141 ( .B1(REG3_REG_23__SCAN_IN), .B2(keyinput_f36), .C1(
        REG3_REG_28__SCAN_IN), .C2(keyinput_f40), .A(n4627), .ZN(n4628) );
  NOR4_X1 U5142 ( .A1(n4631), .A2(n4630), .A3(n4629), .A4(n4628), .ZN(n4652)
         );
  AOI22_X1 U5143 ( .A1(REG3_REG_21__SCAN_IN), .A2(keyinput_f43), .B1(
        REG3_REG_27__SCAN_IN), .B2(keyinput_f34), .ZN(n4632) );
  OAI221_X1 U5144 ( .B1(REG3_REG_21__SCAN_IN), .B2(keyinput_f43), .C1(
        REG3_REG_27__SCAN_IN), .C2(keyinput_f34), .A(n4632), .ZN(n4641) );
  AOI22_X1 U5145 ( .A1(DATAI_9_), .A2(keyinput_f22), .B1(IR_REG_8__SCAN_IN), 
        .B2(keyinput_f63), .ZN(n4633) );
  OAI221_X1 U5146 ( .B1(DATAI_9_), .B2(keyinput_f22), .C1(IR_REG_8__SCAN_IN), 
        .C2(keyinput_f63), .A(n4633), .ZN(n4640) );
  AOI22_X1 U5147 ( .A1(n4636), .A2(keyinput_f7), .B1(n4635), .B2(keyinput_f21), 
        .ZN(n4634) );
  OAI221_X1 U5148 ( .B1(n4636), .B2(keyinput_f7), .C1(n4635), .C2(keyinput_f21), .A(n4634), .ZN(n4639) );
  AOI22_X1 U5149 ( .A1(REG3_REG_16__SCAN_IN), .A2(keyinput_f46), .B1(n2608), 
        .B2(keyinput_f3), .ZN(n4637) );
  OAI221_X1 U5150 ( .B1(REG3_REG_16__SCAN_IN), .B2(keyinput_f46), .C1(n2608), 
        .C2(keyinput_f3), .A(n4637), .ZN(n4638) );
  NOR4_X1 U5151 ( .A1(n4641), .A2(n4640), .A3(n4639), .A4(n4638), .ZN(n4651)
         );
  AOI22_X1 U5152 ( .A1(DATAI_1_), .A2(keyinput_f30), .B1(DATAI_2_), .B2(
        keyinput_f29), .ZN(n4642) );
  OAI221_X1 U5153 ( .B1(DATAI_1_), .B2(keyinput_f30), .C1(DATAI_2_), .C2(
        keyinput_f29), .A(n4642), .ZN(n4649) );
  AOI22_X1 U5154 ( .A1(DATAI_6_), .A2(keyinput_f25), .B1(IR_REG_6__SCAN_IN), 
        .B2(keyinput_f61), .ZN(n4643) );
  OAI221_X1 U5155 ( .B1(DATAI_6_), .B2(keyinput_f25), .C1(IR_REG_6__SCAN_IN), 
        .C2(keyinput_f61), .A(n4643), .ZN(n4648) );
  AOI22_X1 U5156 ( .A1(DATAI_5_), .A2(keyinput_f26), .B1(IR_REG_5__SCAN_IN), 
        .B2(keyinput_f60), .ZN(n4644) );
  OAI221_X1 U5157 ( .B1(DATAI_5_), .B2(keyinput_f26), .C1(IR_REG_5__SCAN_IN), 
        .C2(keyinput_f60), .A(n4644), .ZN(n4647) );
  AOI22_X1 U5158 ( .A1(DATAI_4_), .A2(keyinput_f27), .B1(IR_REG_3__SCAN_IN), 
        .B2(keyinput_f58), .ZN(n4645) );
  OAI221_X1 U5159 ( .B1(DATAI_4_), .B2(keyinput_f27), .C1(IR_REG_3__SCAN_IN), 
        .C2(keyinput_f58), .A(n4645), .ZN(n4646) );
  NOR4_X1 U5160 ( .A1(n4649), .A2(n4648), .A3(n4647), .A4(n4646), .ZN(n4650)
         );
  NAND4_X1 U5161 ( .A1(n4653), .A2(n4652), .A3(n4651), .A4(n4650), .ZN(n4713)
         );
  AOI22_X1 U5162 ( .A1(n4655), .A2(keyinput_f47), .B1(keyinput_f9), .B2(n2545), 
        .ZN(n4654) );
  OAI221_X1 U5163 ( .B1(n4655), .B2(keyinput_f47), .C1(n2545), .C2(keyinput_f9), .A(n4654), .ZN(n4667) );
  AOI22_X1 U5164 ( .A1(n4658), .A2(keyinput_f6), .B1(keyinput_f19), .B2(n4657), 
        .ZN(n4656) );
  OAI221_X1 U5165 ( .B1(n4658), .B2(keyinput_f6), .C1(n4657), .C2(keyinput_f19), .A(n4656), .ZN(n4666) );
  AOI22_X1 U5166 ( .A1(n4661), .A2(keyinput_f2), .B1(n4660), .B2(keyinput_f35), 
        .ZN(n4659) );
  OAI221_X1 U5167 ( .B1(n4661), .B2(keyinput_f2), .C1(n4660), .C2(keyinput_f35), .A(n4659), .ZN(n4665) );
  XNOR2_X1 U5168 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_f56), .ZN(n4663) );
  XNOR2_X1 U5169 ( .A(REG3_REG_25__SCAN_IN), .B(keyinput_f45), .ZN(n4662) );
  NAND2_X1 U5170 ( .A1(n4663), .A2(n4662), .ZN(n4664) );
  NOR4_X1 U5171 ( .A1(n4667), .A2(n4666), .A3(n4665), .A4(n4664), .ZN(n4711)
         );
  INV_X1 U5172 ( .A(REG3_REG_8__SCAN_IN), .ZN(n4670) );
  AOI22_X1 U5173 ( .A1(n4670), .A2(keyinput_f41), .B1(n4669), .B2(keyinput_f53), .ZN(n4668) );
  OAI221_X1 U5174 ( .B1(n4670), .B2(keyinput_f41), .C1(n4669), .C2(
        keyinput_f53), .A(n4668), .ZN(n4678) );
  XNOR2_X1 U5175 ( .A(IR_REG_4__SCAN_IN), .B(keyinput_f59), .ZN(n4674) );
  XNOR2_X1 U5176 ( .A(REG3_REG_12__SCAN_IN), .B(keyinput_f44), .ZN(n4673) );
  XNOR2_X1 U5177 ( .A(DATAI_0_), .B(keyinput_f31), .ZN(n4672) );
  XNOR2_X1 U5178 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_f55), .ZN(n4671) );
  NAND4_X1 U5179 ( .A1(n4674), .A2(n4673), .A3(n4672), .A4(n4671), .ZN(n4677)
         );
  XNOR2_X1 U5180 ( .A(U3149), .B(keyinput_f32), .ZN(n4676) );
  XNOR2_X1 U5181 ( .A(keyinput_f18), .B(n2461), .ZN(n4675) );
  NOR4_X1 U5182 ( .A1(n4678), .A2(n4677), .A3(n4676), .A4(n4675), .ZN(n4710)
         );
  AOI22_X1 U5183 ( .A1(n4681), .A2(keyinput_f16), .B1(n4680), .B2(keyinput_f38), .ZN(n4679) );
  OAI221_X1 U5184 ( .B1(n4681), .B2(keyinput_f16), .C1(n4680), .C2(
        keyinput_f38), .A(n4679), .ZN(n4693) );
  AOI22_X1 U5185 ( .A1(n2396), .A2(keyinput_f33), .B1(keyinput_f4), .B2(n4683), 
        .ZN(n4682) );
  OAI221_X1 U5186 ( .B1(n2396), .B2(keyinput_f33), .C1(n4683), .C2(keyinput_f4), .A(n4682), .ZN(n4692) );
  AOI22_X1 U5187 ( .A1(n4686), .A2(keyinput_f48), .B1(n4685), .B2(keyinput_f39), .ZN(n4684) );
  OAI221_X1 U5188 ( .B1(n4686), .B2(keyinput_f48), .C1(n4685), .C2(
        keyinput_f39), .A(n4684), .ZN(n4691) );
  AOI22_X1 U5189 ( .A1(n4689), .A2(keyinput_f15), .B1(keyinput_f24), .B2(n4688), .ZN(n4687) );
  OAI221_X1 U5190 ( .B1(n4689), .B2(keyinput_f15), .C1(n4688), .C2(
        keyinput_f24), .A(n4687), .ZN(n4690) );
  NOR4_X1 U5191 ( .A1(n4693), .A2(n4692), .A3(n4691), .A4(n4690), .ZN(n4709)
         );
  AOI22_X1 U5192 ( .A1(n4696), .A2(keyinput_f1), .B1(n4695), .B2(keyinput_f5), 
        .ZN(n4694) );
  OAI221_X1 U5193 ( .B1(n4696), .B2(keyinput_f1), .C1(n4695), .C2(keyinput_f5), 
        .A(n4694), .ZN(n4707) );
  AOI22_X1 U5194 ( .A1(n2547), .A2(keyinput_f8), .B1(n4698), .B2(keyinput_f49), 
        .ZN(n4697) );
  OAI221_X1 U5195 ( .B1(n2547), .B2(keyinput_f8), .C1(n4698), .C2(keyinput_f49), .A(n4697), .ZN(n4706) );
  AOI22_X1 U5196 ( .A1(n4701), .A2(keyinput_f37), .B1(keyinput_f20), .B2(n4700), .ZN(n4699) );
  OAI221_X1 U5197 ( .B1(n4701), .B2(keyinput_f37), .C1(n4700), .C2(
        keyinput_f20), .A(n4699), .ZN(n4705) );
  XNOR2_X1 U5198 ( .A(IR_REG_7__SCAN_IN), .B(keyinput_f62), .ZN(n4703) );
  XNOR2_X1 U5199 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_f57), .ZN(n4702) );
  NAND2_X1 U5200 ( .A1(n4703), .A2(n4702), .ZN(n4704) );
  NOR4_X1 U5201 ( .A1(n4707), .A2(n4706), .A3(n4705), .A4(n4704), .ZN(n4708)
         );
  NAND4_X1 U5202 ( .A1(n4711), .A2(n4710), .A3(n4709), .A4(n4708), .ZN(n4712)
         );
  OAI22_X1 U5203 ( .A1(DATAI_3_), .A2(keyinput_f28), .B1(n4713), .B2(n4712), 
        .ZN(n4715) );
  INV_X1 U5204 ( .A(keyinput_g28), .ZN(n4714) );
  NAND2_X1 U5205 ( .A1(n4715), .A2(n4714), .ZN(n4717) );
  OAI211_X1 U5206 ( .C1(n4715), .C2(keyinput_f28), .A(DATAI_3_), .B(
        keyinput_g28), .ZN(n4716) );
  OAI21_X1 U5207 ( .B1(DATAI_3_), .B2(n4717), .A(n4716), .ZN(n4718) );
  OAI21_X1 U5208 ( .B1(n4720), .B2(n4719), .A(n4718), .ZN(n4721) );
  XOR2_X1 U5209 ( .A(n4722), .B(n4721), .Z(U3352) );
  CLKBUF_X1 U2291 ( .A(n2958), .Z(n3660) );
endmodule

