

module b14_C_gen_AntiSAT_k_128_2 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, 
        keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, 
        keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, 
        keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, 
        keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, 
        keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, 
        keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, 
        keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, 
        keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, 
        keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, 
        keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, 
        keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, 
        keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, 
        keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, 
        keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, 
        keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, 
        keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, 
        keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, 
        keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, 
        keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, 
        keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, 
        keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, 
        keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, 
        keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, 
        keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, 
        keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, 
        keyinput_g63, U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, 
        U3344, U3343, U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, 
        U3334, U3333, U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, 
        U3324, U3323, U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, 
        U3316, U3315, U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, 
        U3306, U3305, U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, 
        U3296, U3295, U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, 
        U3475, U3477, U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, 
        U3495, U3497, U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, 
        U3510, U3511, U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, 
        U3520, U3521, U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, 
        U3530, U3531, U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, 
        U3540, U3541, U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, 
        U3290, U3289, U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, 
        U3280, U3279, U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, 
        U3270, U3269, U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, 
        U3261, U3260, U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, 
        U3251, U3250, U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, 
        U3241, U3240, U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, 
        U3558, U3559, U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, 
        U3568, U3569, U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, 
        U3578, U3579, U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, 
        U3233, U3232, U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, 
        U3223, U3222, U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, 
        U3213, U3212, U3211, U3210, U3149, U3148, U4043 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput_f0, keyinput_f1, keyinput_f2,
         keyinput_f3, keyinput_f4, keyinput_f5, keyinput_f6, keyinput_f7,
         keyinput_f8, keyinput_f9, keyinput_f10, keyinput_f11, keyinput_f12,
         keyinput_f13, keyinput_f14, keyinput_f15, keyinput_f16, keyinput_f17,
         keyinput_f18, keyinput_f19, keyinput_f20, keyinput_f21, keyinput_f22,
         keyinput_f23, keyinput_f24, keyinput_f25, keyinput_f26, keyinput_f27,
         keyinput_f28, keyinput_f29, keyinput_f30, keyinput_f31, keyinput_f32,
         keyinput_f33, keyinput_f34, keyinput_f35, keyinput_f36, keyinput_f37,
         keyinput_f38, keyinput_f39, keyinput_f40, keyinput_f41, keyinput_f42,
         keyinput_f43, keyinput_f44, keyinput_f45, keyinput_f46, keyinput_f47,
         keyinput_f48, keyinput_f49, keyinput_f50, keyinput_f51, keyinput_f52,
         keyinput_f53, keyinput_f54, keyinput_f55, keyinput_f56, keyinput_f57,
         keyinput_f58, keyinput_f59, keyinput_f60, keyinput_f61, keyinput_f62,
         keyinput_f63, keyinput_g0, keyinput_g1, keyinput_g2, keyinput_g3,
         keyinput_g4, keyinput_g5, keyinput_g6, keyinput_g7, keyinput_g8,
         keyinput_g9, keyinput_g10, keyinput_g11, keyinput_g12, keyinput_g13,
         keyinput_g14, keyinput_g15, keyinput_g16, keyinput_g17, keyinput_g18,
         keyinput_g19, keyinput_g20, keyinput_g21, keyinput_g22, keyinput_g23,
         keyinput_g24, keyinput_g25, keyinput_g26, keyinput_g27, keyinput_g28,
         keyinput_g29, keyinput_g30, keyinput_g31, keyinput_g32, keyinput_g33,
         keyinput_g34, keyinput_g35, keyinput_g36, keyinput_g37, keyinput_g38,
         keyinput_g39, keyinput_g40, keyinput_g41, keyinput_g42, keyinput_g43,
         keyinput_g44, keyinput_g45, keyinput_g46, keyinput_g47, keyinput_g48,
         keyinput_g49, keyinput_g50, keyinput_g51, keyinput_g52, keyinput_g53,
         keyinput_g54, keyinput_g55, keyinput_g56, keyinput_g57, keyinput_g58,
         keyinput_g59, keyinput_g60, keyinput_g61, keyinput_g62, keyinput_g63;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751;

  NAND2_X1 U2283 ( .A1(n4069), .A2(n3781), .ZN(n2720) );
  AND2_X1 U2284 ( .A1(n2260), .A2(n2258), .ZN(n3761) );
  INV_X1 U2285 ( .A(n2765), .ZN(n2738) );
  NAND2_X1 U2286 ( .A1(n2104), .A2(n2053), .ZN(n4090) );
  INV_X1 U2287 ( .A(n2896), .ZN(n2902) );
  INV_X2 U2288 ( .A(n2509), .ZN(n3783) );
  AOI21_X1 U2289 ( .B1(n4398), .B2(n3034), .A(n3033), .ZN(n3138) );
  NAND4_X2 U2290 ( .A1(n2340), .A2(n2339), .A3(n2338), .A4(n2337), .ZN(n3965)
         );
  XNOR2_X2 U2291 ( .A(n2297), .B(IR_REG_30__SCAN_IN), .ZN(n2962) );
  NAND2_X2 U2292 ( .A1(n2686), .A2(n2685), .ZN(n2942) );
  NOR2_X2 U2293 ( .A1(n4494), .A2(n4493), .ZN(n4495) );
  NOR2_X2 U2294 ( .A1(n4485), .A2(n4028), .ZN(n4494) );
  INV_X1 U2295 ( .A(n2509), .ZN(n2041) );
  INV_X2 U2296 ( .A(n2791), .ZN(n2886) );
  NAND2_X1 U2297 ( .A1(n4474), .A2(n4025), .ZN(n4027) );
  NAND2_X1 U2298 ( .A1(n2643), .A2(n3799), .ZN(n3501) );
  NAND2_X1 U2299 ( .A1(n4095), .A2(n4083), .ZN(n4082) );
  NAND2_X1 U2300 ( .A1(n3435), .A2(n3434), .ZN(n3433) );
  AOI21_X1 U2301 ( .B1(n2196), .B2(n2195), .A(n2194), .ZN(n3435) );
  NAND2_X1 U2302 ( .A1(n2100), .A2(n2098), .ZN(n4409) );
  NAND2_X2 U2303 ( .A1(n3100), .A2(n4511), .ZN(n4514) );
  XNOR2_X1 U2304 ( .A(n3032), .B(n2113), .ZN(n3000) );
  AND2_X1 U2305 ( .A1(n2115), .A2(n2114), .ZN(n3045) );
  OR2_X1 U2306 ( .A1(n3064), .A2(n2116), .ZN(n2115) );
  NAND2_X2 U2307 ( .A1(n2348), .A2(n2347), .ZN(n3966) );
  AND2_X1 U2308 ( .A1(n3066), .A2(REG1_REG_4__SCAN_IN), .ZN(n3064) );
  AND3_X1 U2309 ( .A1(n2346), .A2(n2345), .A3(n2344), .ZN(n2347) );
  NAND2_X2 U2310 ( .A1(n2198), .A2(n2199), .ZN(n2527) );
  INV_X1 U2311 ( .A(n2621), .ZN(n2627) );
  NAND2_X1 U2312 ( .A1(n3015), .A2(n2995), .ZN(n2997) );
  AND2_X1 U2313 ( .A1(n2102), .A2(n2101), .ZN(n2271) );
  AND4_X1 U2314 ( .A1(n2280), .A2(n2279), .A3(n2278), .A4(n2277), .ZN(n2281)
         );
  INV_X1 U2315 ( .A(IR_REG_6__SCAN_IN), .ZN(n4693) );
  NOR2_X1 U2316 ( .A1(IR_REG_2__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2102)
         );
  INV_X1 U2317 ( .A(IR_REG_7__SCAN_IN), .ZN(n2416) );
  NAND2_X1 U2318 ( .A1(n2295), .A2(n2294), .ZN(n2042) );
  XNOR2_X2 U2319 ( .A(n2357), .B(IR_REG_2__SCAN_IN), .ZN(n4402) );
  AOI21_X1 U2320 ( .B1(n4072), .B2(n2594), .A(n2593), .ZN(n4060) );
  NAND2_X1 U2321 ( .A1(n2289), .A2(n2256), .ZN(n2292) );
  AND2_X1 U2322 ( .A1(n2603), .A2(n2602), .ZN(n3754) );
  OR2_X1 U2323 ( .A1(n3634), .A2(n2457), .ZN(n2603) );
  NAND2_X1 U2324 ( .A1(n4440), .A2(REG2_REG_12__SCAN_IN), .ZN(n4439) );
  AOI21_X1 U2325 ( .B1(n4093), .B2(n2584), .A(n2583), .ZN(n4072) );
  INV_X1 U2326 ( .A(n3736), .ZN(n2217) );
  NOR2_X1 U2327 ( .A1(n2047), .A2(n2207), .ZN(n2206) );
  INV_X1 U2328 ( .A(n2218), .ZN(n2207) );
  NAND2_X1 U2329 ( .A1(n3022), .A2(n2137), .ZN(n2136) );
  NAND2_X1 U2330 ( .A1(n4402), .A2(REG2_REG_2__SCAN_IN), .ZN(n2137) );
  NAND2_X1 U2331 ( .A1(n4408), .A2(n4013), .ZN(n4015) );
  AND2_X1 U2332 ( .A1(n3917), .A2(n2109), .ZN(n2108) );
  OR2_X1 U2333 ( .A1(n2110), .A2(n2654), .ZN(n2109) );
  NAND2_X1 U2334 ( .A1(n3914), .A2(n3791), .ZN(n2110) );
  NAND2_X1 U2335 ( .A1(n2506), .A2(n4317), .ZN(n2507) );
  NOR2_X1 U2336 ( .A1(n3883), .A2(n2124), .ZN(n2123) );
  INV_X1 U2337 ( .A(n3795), .ZN(n2124) );
  NAND2_X1 U2338 ( .A1(n3122), .A2(n3718), .ZN(n3813) );
  AND2_X1 U2339 ( .A1(n2043), .A2(n2290), .ZN(n2256) );
  NOR2_X1 U2340 ( .A1(IR_REG_14__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2279)
         );
  NOR2_X1 U2341 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2278)
         );
  NOR2_X1 U2342 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2277)
         );
  INV_X1 U2343 ( .A(n2558), .ZN(n2557) );
  INV_X1 U2344 ( .A(n2962), .ZN(n2199) );
  NAND2_X1 U2345 ( .A1(n2041), .A2(REG0_REG_1__SCAN_IN), .ZN(n2254) );
  INV_X1 U2346 ( .A(n3622), .ZN(n2873) );
  OR2_X1 U2347 ( .A1(n2960), .A2(n2962), .ZN(n2509) );
  INV_X1 U2348 ( .A(n2730), .ZN(n2370) );
  XNOR2_X1 U2349 ( .A(n2136), .B(n2996), .ZN(n3983) );
  INV_X1 U2350 ( .A(n4537), .ZN(n4009) );
  NAND2_X1 U2351 ( .A1(n4409), .A2(n4410), .ZN(n4408) );
  NOR2_X1 U2352 ( .A1(n2144), .A2(n2145), .ZN(n2143) );
  AND2_X1 U2353 ( .A1(n2082), .A2(n2074), .ZN(n4093) );
  NAND2_X1 U2354 ( .A1(n4109), .A2(n2574), .ZN(n2082) );
  NAND2_X1 U2355 ( .A1(n2445), .A2(n2444), .ZN(n3371) );
  NAND2_X1 U2356 ( .A1(n3336), .A2(n2443), .ZN(n2445) );
  NAND2_X1 U2357 ( .A1(n2662), .A2(IR_REG_28__SCAN_IN), .ZN(n2294) );
  NOR3_X1 U2358 ( .A1(n4082), .A2(n4061), .A3(n2924), .ZN(n2724) );
  OR2_X1 U2359 ( .A1(n2911), .A2(n2636), .ZN(n4330) );
  NAND2_X1 U2360 ( .A1(n2289), .A2(n2255), .ZN(n2666) );
  NAND2_X1 U2361 ( .A1(n3998), .A2(n4439), .ZN(n4452) );
  NOR2_X1 U2362 ( .A1(n4462), .A2(n2487), .ZN(n4461) );
  AND2_X1 U2363 ( .A1(n2188), .A2(n2063), .ZN(n2718) );
  INV_X1 U2364 ( .A(n2212), .ZN(n2210) );
  NAND2_X1 U2365 ( .A1(n2841), .A2(n2842), .ZN(n2218) );
  NAND2_X1 U2366 ( .A1(n3522), .A2(n2262), .ZN(n2261) );
  INV_X1 U2367 ( .A(n3521), .ZN(n2262) );
  NAND2_X1 U2368 ( .A1(n3520), .A2(n2263), .ZN(n2260) );
  NAND2_X1 U2369 ( .A1(n2828), .A2(n3521), .ZN(n2263) );
  NAND2_X1 U2370 ( .A1(n2099), .A2(REG2_REG_8__SCAN_IN), .ZN(n2162) );
  INV_X1 U2371 ( .A(n2162), .ZN(n2155) );
  INV_X1 U2372 ( .A(n2146), .ZN(n2144) );
  AND2_X1 U2373 ( .A1(n2655), .A2(n4073), .ZN(n3923) );
  OAI21_X1 U2374 ( .B1(n4149), .B2(n2166), .A(n2565), .ZN(n2165) );
  OAI21_X1 U2375 ( .B1(n2470), .B2(n2192), .A(n2264), .ZN(n2191) );
  AND2_X1 U2376 ( .A1(n2374), .A2(n2358), .ZN(n2376) );
  OR2_X1 U2377 ( .A1(n2375), .A2(n3206), .ZN(n2179) );
  OR2_X1 U2378 ( .A1(n2691), .A2(n2956), .ZN(n2732) );
  NAND2_X1 U2379 ( .A1(n4167), .A2(n4144), .ZN(n2094) );
  INV_X1 U2380 ( .A(IR_REG_26__SCAN_IN), .ZN(n2257) );
  INV_X1 U2381 ( .A(IR_REG_25__SCAN_IN), .ZN(n2288) );
  OAI21_X1 U2382 ( .B1(n2681), .B2(IR_REG_22__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2688) );
  NAND2_X1 U2383 ( .A1(n2532), .A2(n2531), .ZN(n2621) );
  INV_X1 U2384 ( .A(IR_REG_18__SCAN_IN), .ZN(n2531) );
  INV_X1 U2385 ( .A(n2530), .ZN(n2532) );
  NAND2_X1 U2386 ( .A1(n3746), .A2(n2247), .ZN(n2244) );
  NOR2_X1 U2387 ( .A1(n3745), .A2(n2246), .ZN(n2245) );
  NAND2_X1 U2388 ( .A1(n2237), .A2(n2235), .ZN(n2234) );
  INV_X1 U2389 ( .A(n2240), .ZN(n2235) );
  NAND2_X1 U2390 ( .A1(n2066), .A2(n2236), .ZN(n2232) );
  INV_X1 U2391 ( .A(n2237), .ZN(n2236) );
  INV_X1 U2392 ( .A(n3965), .ZN(n3122) );
  AND2_X1 U2393 ( .A1(n2916), .A2(n2732), .ZN(n2896) );
  NOR2_X1 U2394 ( .A1(n3761), .A2(n3682), .ZN(n2838) );
  NAND2_X1 U2395 ( .A1(n3762), .A2(n3764), .ZN(n2837) );
  NAND2_X1 U2396 ( .A1(n2242), .A2(n2248), .ZN(n2241) );
  INV_X1 U2397 ( .A(n2882), .ZN(n2242) );
  NAND2_X1 U2398 ( .A1(n2738), .A2(n2737), .ZN(n2741) );
  AOI21_X1 U2399 ( .B1(n3395), .B2(n2225), .A(n2224), .ZN(n2223) );
  INV_X1 U2400 ( .A(n3394), .ZN(n2225) );
  INV_X1 U2401 ( .A(n3395), .ZN(n2226) );
  NAND2_X1 U2402 ( .A1(n3725), .A2(n2068), .ZN(n2201) );
  NAND2_X1 U2403 ( .A1(n2303), .A2(REG3_REG_10__SCAN_IN), .ZN(n2459) );
  INV_X1 U2404 ( .A(n2447), .ZN(n2303) );
  OR2_X1 U2405 ( .A1(n2459), .A2(n2458), .ZN(n2472) );
  NAND2_X1 U2406 ( .A1(n2575), .A2(REG3_REG_25__SCAN_IN), .ZN(n2585) );
  OR2_X1 U2407 ( .A1(n2585), .A2(n3750), .ZN(n2596) );
  NOR2_X1 U2408 ( .A1(n3628), .A2(n2953), .ZN(n2685) );
  AND4_X1 U2409 ( .A1(n2414), .A2(n2413), .A3(n2412), .A4(n2411), .ZN(n3354)
         );
  AOI21_X1 U2410 ( .B1(n3983), .B2(REG2_REG_3__SCAN_IN), .A(n2057), .ZN(n2988)
         );
  AND2_X1 U2411 ( .A1(n2999), .A2(n4400), .ZN(n2116) );
  INV_X1 U2412 ( .A(n4398), .ZN(n2113) );
  NOR2_X1 U2413 ( .A1(n2160), .A2(n2158), .ZN(n2157) );
  INV_X1 U2414 ( .A(n4412), .ZN(n2158) );
  NAND2_X1 U2415 ( .A1(n4418), .A2(n4016), .ZN(n4428) );
  NAND2_X1 U2416 ( .A1(n4428), .A2(n4429), .ZN(n4427) );
  XNOR2_X1 U2417 ( .A(n3997), .B(n4532), .ZN(n4440) );
  OR2_X1 U2418 ( .A1(n4008), .A2(REG2_REG_13__SCAN_IN), .ZN(n2146) );
  OR2_X1 U2419 ( .A1(n4469), .A2(n2135), .ZN(n2134) );
  AND2_X1 U2420 ( .A1(n4007), .A2(REG2_REG_15__SCAN_IN), .ZN(n2135) );
  NAND2_X1 U2421 ( .A1(n4489), .A2(n2153), .ZN(n2152) );
  NAND2_X1 U2422 ( .A1(n4528), .A2(n2499), .ZN(n2153) );
  OR2_X1 U2423 ( .A1(n4200), .A2(n2107), .ZN(n2104) );
  INV_X1 U2424 ( .A(n2108), .ZN(n2107) );
  AOI21_X1 U2425 ( .B1(n2108), .B2(n2044), .A(n2106), .ZN(n2105) );
  AOI22_X1 U2426 ( .A1(n4157), .A2(n2545), .B1(n4167), .B2(n4193), .ZN(n4150)
         );
  OR2_X1 U2427 ( .A1(n3595), .A2(n3790), .ZN(n4200) );
  NOR2_X1 U2428 ( .A1(n2042), .A2(n2538), .ZN(n4184) );
  INV_X1 U2429 ( .A(n2170), .ZN(n2169) );
  NAND2_X1 U2430 ( .A1(n2080), .A2(n2079), .ZN(n2081) );
  OAI21_X1 U2431 ( .B1(n2061), .B2(n2171), .A(n4228), .ZN(n2170) );
  INV_X1 U2432 ( .A(n3793), .ZN(n2122) );
  AND2_X1 U2433 ( .A1(n2120), .A2(n3889), .ZN(n2119) );
  NAND2_X1 U2434 ( .A1(n2121), .A2(n3793), .ZN(n2120) );
  AND2_X1 U2435 ( .A1(n3909), .A2(n3911), .ZN(n3889) );
  NOR2_X1 U2436 ( .A1(n3572), .A2(n3889), .ZN(n3571) );
  NAND2_X1 U2437 ( .A1(n2645), .A2(n2123), .ZN(n3507) );
  NAND2_X1 U2438 ( .A1(n3542), .A2(n3478), .ZN(n2195) );
  AND2_X1 U2439 ( .A1(n3956), .A2(n3448), .ZN(n2194) );
  INV_X1 U2440 ( .A(n3477), .ZN(n2196) );
  NAND2_X1 U2441 ( .A1(n2193), .A2(n2470), .ZN(n3384) );
  INV_X1 U2442 ( .A(n3382), .ZN(n2193) );
  INV_X1 U2443 ( .A(n3959), .ZN(n3332) );
  OR2_X1 U2444 ( .A1(n3286), .A2(n2426), .ZN(n3336) );
  NAND2_X1 U2445 ( .A1(n2174), .A2(n2175), .ZN(n3244) );
  NAND2_X1 U2446 ( .A1(n2177), .A2(n2052), .ZN(n2175) );
  NAND2_X1 U2447 ( .A1(n3146), .A2(n2176), .ZN(n2174) );
  NAND2_X1 U2448 ( .A1(n2179), .A2(n2392), .ZN(n2177) );
  OAI21_X1 U2449 ( .B1(n3238), .B2(n3224), .A(n3826), .ZN(n3242) );
  NAND2_X1 U2450 ( .A1(n2661), .A2(n2660), .ZN(n4225) );
  NOR2_X1 U2451 ( .A1(n2509), .A2(n2367), .ZN(n2132) );
  NAND2_X1 U2452 ( .A1(n2042), .A2(n4403), .ZN(n2087) );
  NAND2_X1 U2453 ( .A1(n2089), .A2(DATAI_1_), .ZN(n2088) );
  AND2_X1 U2454 ( .A1(n2908), .A2(n2969), .ZN(n3098) );
  OR2_X1 U2455 ( .A1(n4051), .A2(n2924), .ZN(n2096) );
  NAND2_X1 U2456 ( .A1(n4060), .A2(n2604), .ZN(n2188) );
  NAND2_X1 U2457 ( .A1(n4150), .A2(n4149), .ZN(n4283) );
  AND4_X1 U2458 ( .A1(n2491), .A2(n2490), .A3(n2489), .A4(n2488), .ZN(n3584)
         );
  INV_X1 U2459 ( .A(n4225), .ZN(n4302) );
  AND2_X1 U2460 ( .A1(n3103), .A2(n2636), .ZN(n4231) );
  INV_X1 U2461 ( .A(n2737), .ZN(n3112) );
  INV_X1 U2462 ( .A(n2909), .ZN(n3099) );
  NAND2_X1 U2463 ( .A1(n2954), .A2(n2684), .ZN(n2968) );
  NAND2_X1 U2464 ( .A1(n2942), .A2(n4525), .ZN(n3095) );
  AND2_X1 U2465 ( .A1(n2256), .A2(n2296), .ZN(n2255) );
  AND4_X1 U2466 ( .A1(n2286), .A2(n2285), .A3(n2284), .A4(n2283), .ZN(n2287)
         );
  NOR2_X1 U2467 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2286)
         );
  NOR2_X1 U2468 ( .A1(IR_REG_21__SCAN_IN), .A2(IR_REG_24__SCAN_IN), .ZN(n2285)
         );
  INV_X1 U2469 ( .A(IR_REG_9__SCAN_IN), .ZN(n2272) );
  AND2_X1 U2470 ( .A1(n2572), .A2(n2571), .ZN(n3676) );
  OR2_X1 U2471 ( .A1(n3705), .A2(n2457), .ZN(n2572) );
  NAND2_X1 U2472 ( .A1(n2200), .A2(n2199), .ZN(n2364) );
  INV_X1 U2473 ( .A(n3546), .ZN(n3958) );
  NAND2_X1 U2474 ( .A1(n2986), .A2(n2987), .ZN(n3022) );
  NAND2_X1 U2475 ( .A1(n2139), .A2(n2138), .ZN(n4462) );
  OR2_X1 U2476 ( .A1(n4452), .A2(n2142), .ZN(n2138) );
  INV_X1 U2477 ( .A(n2141), .ZN(n2140) );
  NOR2_X1 U2478 ( .A1(n4471), .A2(n4470), .ZN(n4469) );
  XNOR2_X1 U2479 ( .A(n2134), .B(n2133), .ZN(n4481) );
  NAND2_X1 U2480 ( .A1(n4481), .A2(n4479), .ZN(n4480) );
  NAND2_X1 U2481 ( .A1(n4490), .A2(n4488), .ZN(n4489) );
  NAND2_X1 U2482 ( .A1(n2151), .A2(n4450), .ZN(n2150) );
  NAND2_X1 U2483 ( .A1(n2152), .A2(n4501), .ZN(n2151) );
  AOI21_X1 U2484 ( .B1(n4503), .B2(ADDR_REG_18__SCAN_IN), .A(n4502), .ZN(n2149) );
  NOR2_X1 U2485 ( .A1(n2152), .A2(n4501), .ZN(n4500) );
  AND2_X1 U2486 ( .A1(n2991), .A2(n2990), .ZN(n4505) );
  AOI21_X1 U2487 ( .B1(n4046), .B2(n4554), .A(n2674), .ZN(n2717) );
  OAI211_X1 U2488 ( .C1(n2188), .C2(n3905), .A(n2185), .B(n2183), .ZN(n3619)
         );
  OR2_X1 U2489 ( .A1(n3905), .A2(n2063), .ZN(n2185) );
  NAND2_X1 U2490 ( .A1(n2188), .A2(n2184), .ZN(n2183) );
  AND2_X1 U2491 ( .A1(n3905), .A2(n2063), .ZN(n2184) );
  INV_X1 U2492 ( .A(n2181), .ZN(n2180) );
  OAI21_X1 U2493 ( .B1(n2187), .B2(n4560), .A(n2186), .ZN(n2181) );
  NAND2_X1 U2494 ( .A1(n4560), .A2(REG0_REG_28__SCAN_IN), .ZN(n2186) );
  NAND2_X1 U2495 ( .A1(n4562), .A2(n4554), .ZN(n2182) );
  OAI21_X1 U2496 ( .B1(n2049), .B2(n3613), .A(n2725), .ZN(n3608) );
  NAND2_X1 U2497 ( .A1(n2130), .A2(n4251), .ZN(n4350) );
  AOI211_X1 U2498 ( .C1(n4319), .C2(n4250), .A(n4249), .B(n4248), .ZN(n4251)
         );
  OR2_X1 U2499 ( .A1(n4252), .A2(n4315), .ZN(n2130) );
  INV_X1 U2500 ( .A(n2954), .ZN(n3628) );
  NAND2_X1 U2501 ( .A1(n2289), .A2(n2117), .ZN(n2965) );
  AND2_X1 U2502 ( .A1(n2255), .A2(n2118), .ZN(n2117) );
  INV_X1 U2503 ( .A(IR_REG_29__SCAN_IN), .ZN(n2118) );
  INV_X1 U2504 ( .A(IR_REG_31__SCAN_IN), .ZN(n2964) );
  NOR2_X1 U2505 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_11__SCAN_IN), .ZN(n2280)
         );
  AND2_X1 U2506 ( .A1(REG3_REG_3__SCAN_IN), .A2(REG3_REG_4__SCAN_IN), .ZN(
        n2333) );
  NOR2_X1 U2507 ( .A1(n2472), .A2(n4681), .ZN(n2325) );
  OR2_X1 U2508 ( .A1(n2566), .A2(n3706), .ZN(n2576) );
  AND2_X1 U2509 ( .A1(n2325), .A2(REG3_REG_13__SCAN_IN), .ZN(n2324) );
  OR2_X1 U2510 ( .A1(n4112), .A2(n4258), .ZN(n4073) );
  AND2_X1 U2511 ( .A1(n2512), .A2(REG3_REG_18__SCAN_IN), .ZN(n2524) );
  INV_X1 U2512 ( .A(n3572), .ZN(n2080) );
  NOR2_X1 U2513 ( .A1(n2171), .A2(n3889), .ZN(n2079) );
  INV_X1 U2514 ( .A(n2123), .ZN(n2121) );
  AND2_X1 U2515 ( .A1(n3487), .A2(n3469), .ZN(n3840) );
  AND2_X1 U2516 ( .A1(n2376), .A2(n2052), .ZN(n2176) );
  NAND2_X1 U2517 ( .A1(n2730), .A2(n2366), .ZN(n3806) );
  INV_X1 U2518 ( .A(n2732), .ZN(n3101) );
  INV_X1 U2519 ( .A(n3403), .ZN(n2801) );
  INV_X1 U2520 ( .A(n3191), .ZN(n3249) );
  NAND3_X1 U2521 ( .A1(n2112), .A2(n3112), .A3(n3118), .ZN(n3113) );
  NOR2_X1 U2522 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_18__SCAN_IN), .ZN(n2283)
         );
  NOR2_X1 U2523 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_23__SCAN_IN), .ZN(n2284)
         );
  NAND2_X1 U2524 ( .A1(n2627), .A2(n2623), .ZN(n2681) );
  NAND2_X1 U2525 ( .A1(n2520), .A2(n2519), .ZN(n2530) );
  AND2_X1 U2526 ( .A1(n2282), .A2(n2281), .ZN(n2520) );
  NAND2_X1 U2527 ( .A1(n2779), .A2(n2203), .ZN(n2202) );
  NOR2_X1 U2528 ( .A1(n3185), .A2(n2204), .ZN(n2203) );
  OAI22_X1 U2529 ( .A1(n3584), .A2(n2765), .B1(n2791), .B2(n3557), .ZN(n3521)
         );
  XNOR2_X1 U2530 ( .A(n2762), .B(n2902), .ZN(n2766) );
  NAND2_X1 U2531 ( .A1(n2761), .A2(n2760), .ZN(n2762) );
  NAND2_X1 U2532 ( .A1(n2217), .A2(n2077), .ZN(n2212) );
  NAND2_X1 U2533 ( .A1(n3703), .A2(n2248), .ZN(n2240) );
  AOI21_X1 U2534 ( .B1(n2241), .B2(n2239), .A(n2238), .ZN(n2237) );
  INV_X1 U2535 ( .A(n3703), .ZN(n2239) );
  AND2_X1 U2536 ( .A1(n2882), .A2(n2881), .ZN(n2238) );
  OR2_X1 U2537 ( .A1(n2317), .A2(n4605), .ZN(n2497) );
  NOR2_X1 U2538 ( .A1(n3343), .A2(n2250), .ZN(n2249) );
  INV_X1 U2539 ( .A(n2252), .ZN(n2250) );
  NAND2_X1 U2540 ( .A1(n3299), .A2(n3298), .ZN(n2252) );
  NAND2_X1 U2541 ( .A1(n3297), .A2(n2253), .ZN(n2251) );
  OR2_X1 U2542 ( .A1(n3299), .A2(n3298), .ZN(n2253) );
  AND2_X1 U2543 ( .A1(n2086), .A2(n2085), .ZN(n3092) );
  NAND2_X1 U2544 ( .A1(n2042), .A2(IR_REG_0__SCAN_IN), .ZN(n2085) );
  NAND2_X1 U2545 ( .A1(n2089), .A2(DATAI_0_), .ZN(n2086) );
  NOR2_X1 U2546 ( .A1(n2300), .A2(n2359), .ZN(n2200) );
  INV_X1 U2547 ( .A(n2209), .ZN(n2208) );
  OAI21_X1 U2548 ( .B1(n2062), .B2(n2047), .A(n2855), .ZN(n2209) );
  OR2_X1 U2549 ( .A1(n2547), .A2(n2546), .ZN(n2558) );
  INV_X1 U2550 ( .A(REG3_REG_11__SCAN_IN), .ZN(n2458) );
  OAI22_X1 U2551 ( .A1(n2730), .A2(n2791), .B1(n2901), .B2(n2734), .ZN(n2733)
         );
  NAND2_X1 U2552 ( .A1(n2071), .A2(n2218), .ZN(n2213) );
  NOR2_X1 U2553 ( .A1(n2259), .A2(n2831), .ZN(n2258) );
  INV_X1 U2554 ( .A(n2261), .ZN(n2259) );
  NAND2_X1 U2555 ( .A1(n2832), .A2(n2831), .ZN(n3762) );
  NAND2_X1 U2556 ( .A1(n2324), .A2(REG3_REG_14__SCAN_IN), .ZN(n2486) );
  OR2_X1 U2557 ( .A1(n2731), .A2(n4395), .ZN(n2916) );
  AND4_X1 U2558 ( .A1(n2331), .A2(n2330), .A3(n2329), .A4(n2328), .ZN(n3542)
         );
  OR2_X1 U2559 ( .A1(n2457), .A2(n3719), .ZN(n2339) );
  INV_X1 U2560 ( .A(IR_REG_5__SCAN_IN), .ZN(n2388) );
  NOR2_X1 U2561 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_4__SCAN_IN), .ZN(n2270)
         );
  INV_X1 U2562 ( .A(IR_REG_8__SCAN_IN), .ZN(n4655) );
  NAND2_X1 U2563 ( .A1(n3992), .A2(n2162), .ZN(n2159) );
  NAND2_X1 U2564 ( .A1(n4011), .A2(n2099), .ZN(n2098) );
  NAND2_X1 U2565 ( .A1(n4010), .A2(REG1_REG_8__SCAN_IN), .ZN(n2100) );
  AOI21_X1 U2566 ( .B1(n2155), .B2(n2157), .A(n2069), .ZN(n2154) );
  INV_X1 U2567 ( .A(n2157), .ZN(n2156) );
  NAND2_X1 U2568 ( .A1(n4430), .A2(n3996), .ZN(n3997) );
  NAND2_X1 U2569 ( .A1(n4427), .A2(n4017), .ZN(n4019) );
  AOI21_X1 U2570 ( .B1(n2143), .B2(n4448), .A(n2078), .ZN(n2141) );
  OR2_X1 U2571 ( .A1(n4448), .A2(n4022), .ZN(n2142) );
  INV_X1 U2572 ( .A(n3893), .ZN(n2103) );
  OAI22_X1 U2573 ( .A1(n4150), .A2(n2163), .B1(n2164), .B2(n2268), .ZN(n4109)
         );
  NAND2_X1 U2574 ( .A1(n2167), .A2(n2556), .ZN(n2163) );
  INV_X1 U2575 ( .A(n2165), .ZN(n2164) );
  OAI21_X1 U2576 ( .B1(n4200), .B2(n3791), .A(n3914), .ZN(n4155) );
  NAND2_X1 U2577 ( .A1(n3569), .A2(n3911), .ZN(n3595) );
  NAND2_X1 U2578 ( .A1(n3433), .A2(n2494), .ZN(n3509) );
  NAND2_X1 U2579 ( .A1(n3458), .A2(n3541), .ZN(n2482) );
  INV_X1 U2580 ( .A(n2191), .ZN(n2190) );
  AND2_X1 U2581 ( .A1(n3799), .A2(n3839), .ZN(n3881) );
  INV_X1 U2582 ( .A(n2432), .ZN(n2302) );
  OAI21_X1 U2583 ( .B1(n3277), .B2(n2640), .A(n3823), .ZN(n3352) );
  OAI22_X1 U2584 ( .A1(n3244), .A2(n2407), .B1(n3963), .B2(n3191), .ZN(n3286)
         );
  NAND2_X1 U2585 ( .A1(n2125), .A2(n3818), .ZN(n3277) );
  NAND2_X1 U2586 ( .A1(n3242), .A2(n3825), .ZN(n2125) );
  AND2_X1 U2587 ( .A1(n2639), .A2(n3823), .ZN(n3888) );
  AND2_X1 U2588 ( .A1(n2377), .A2(REG3_REG_6__SCAN_IN), .ZN(n2409) );
  OAI21_X1 U2589 ( .B1(n3212), .B2(n2638), .A(n3816), .ZN(n3238) );
  NAND2_X1 U2590 ( .A1(n3162), .A2(n3812), .ZN(n3212) );
  AND4_X1 U2591 ( .A1(n2385), .A2(n2384), .A3(n2383), .A4(n2382), .ZN(n3716)
         );
  NAND2_X1 U2592 ( .A1(n3146), .A2(n2376), .ZN(n2178) );
  NAND2_X1 U2593 ( .A1(n3163), .A2(n3885), .ZN(n3162) );
  NAND2_X1 U2594 ( .A1(n3110), .A2(n2371), .ZN(n3147) );
  NAND2_X1 U2595 ( .A1(n3113), .A2(n3806), .ZN(n3151) );
  NAND2_X1 U2596 ( .A1(n3151), .A2(n3880), .ZN(n3150) );
  INV_X1 U2597 ( .A(n2300), .ZN(n2198) );
  NAND2_X1 U2598 ( .A1(n3783), .A2(REG0_REG_2__SCAN_IN), .ZN(n2355) );
  NAND2_X1 U2599 ( .A1(n3112), .A2(n3118), .ZN(n3801) );
  NOR2_X1 U2600 ( .A1(n2051), .A2(n4245), .ZN(n4242) );
  AND2_X1 U2601 ( .A1(n3614), .A2(n2722), .ZN(n2187) );
  INV_X1 U2602 ( .A(n2887), .ZN(n4083) );
  AND2_X1 U2603 ( .A1(n4110), .A2(n4258), .ZN(n4095) );
  NAND2_X1 U2604 ( .A1(n2093), .A2(n2092), .ZN(n2091) );
  INV_X1 U2605 ( .A(n2094), .ZN(n2093) );
  NOR2_X1 U2606 ( .A1(n4184), .A2(n2708), .ZN(n2092) );
  NOR2_X1 U2607 ( .A1(n4131), .A2(n4268), .ZN(n4110) );
  NOR3_X1 U2608 ( .A1(n4210), .A2(n4184), .A3(n4287), .ZN(n4159) );
  NOR2_X1 U2609 ( .A1(n4210), .A2(n4184), .ZN(n4181) );
  NAND2_X1 U2610 ( .A1(n4232), .A2(n2522), .ZN(n4230) );
  OR2_X1 U2611 ( .A1(n4230), .A2(n3652), .ZN(n4210) );
  OR2_X1 U2612 ( .A1(n3573), .A2(n3685), .ZN(n3597) );
  NOR2_X1 U2613 ( .A1(n3597), .A2(n4317), .ZN(n4232) );
  NAND2_X1 U2614 ( .A1(n3480), .A2(n2097), .ZN(n3573) );
  NOR2_X1 U2615 ( .A1(n3767), .A2(n3526), .ZN(n2097) );
  INV_X1 U2616 ( .A(n3515), .ZN(n3767) );
  NAND2_X1 U2617 ( .A1(n3480), .A2(n3557), .ZN(n3510) );
  AND2_X1 U2618 ( .A1(n3492), .A2(n3478), .ZN(n3480) );
  NOR2_X1 U2619 ( .A1(n3491), .A2(n3497), .ZN(n3492) );
  OR2_X1 U2620 ( .A1(n3385), .A2(n3455), .ZN(n3491) );
  NAND2_X1 U2621 ( .A1(n3372), .A2(n3423), .ZN(n3385) );
  INV_X1 U2622 ( .A(n3643), .ZN(n3423) );
  AND2_X1 U2623 ( .A1(n3361), .A2(n2801), .ZN(n3372) );
  AND4_X1 U2624 ( .A1(n2422), .A2(n2421), .A3(n2420), .A4(n2419), .ZN(n3406)
         );
  INV_X1 U2625 ( .A(n3353), .ZN(n3363) );
  OR2_X1 U2626 ( .A1(n3281), .A2(n3321), .ZN(n3362) );
  NOR2_X1 U2627 ( .A1(n3362), .A2(n3363), .ZN(n3361) );
  INV_X1 U2628 ( .A(n3289), .ZN(n3230) );
  OR2_X1 U2629 ( .A1(n3217), .A2(n3718), .ZN(n3231) );
  NOR2_X1 U2630 ( .A1(n3231), .A2(n3230), .ZN(n3250) );
  NOR2_X1 U2631 ( .A1(n3268), .A2(n3157), .ZN(n3167) );
  INV_X1 U2632 ( .A(n3165), .ZN(n3260) );
  NAND2_X1 U2633 ( .A1(n2734), .A2(n3092), .ZN(n3157) );
  INV_X1 U2634 ( .A(n4288), .ZN(n4333) );
  INV_X1 U2635 ( .A(n4330), .ZN(n4318) );
  AND3_X1 U2636 ( .A1(n2705), .A2(n2704), .A3(n2908), .ZN(n2712) );
  AND2_X1 U2637 ( .A1(n2050), .A2(n2293), .ZN(n2662) );
  AND2_X1 U2638 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2293)
         );
  NAND2_X1 U2639 ( .A1(n2292), .A2(n2291), .ZN(n2663) );
  INV_X1 U2640 ( .A(IR_REG_20__SCAN_IN), .ZN(n2633) );
  NAND2_X1 U2641 ( .A1(n2632), .A2(IR_REG_31__SCAN_IN), .ZN(n2634) );
  AND2_X1 U2642 ( .A1(n2313), .A2(n2312), .ZN(n4007) );
  INV_X1 U2643 ( .A(IR_REG_3__SCAN_IN), .ZN(n4626) );
  NAND2_X1 U2644 ( .A1(n3747), .A2(n2244), .ZN(n2243) );
  NAND2_X1 U2645 ( .A1(n2211), .A2(n2212), .ZN(n3650) );
  NAND2_X1 U2646 ( .A1(n2214), .A2(n2062), .ZN(n2211) );
  NAND2_X1 U2647 ( .A1(n2222), .A2(n3395), .ZN(n3413) );
  NAND2_X1 U2648 ( .A1(n3393), .A2(n3394), .ZN(n2222) );
  NAND2_X1 U2649 ( .A1(n2233), .A2(n2237), .ZN(n3674) );
  NAND2_X1 U2650 ( .A1(n2945), .A2(n2240), .ZN(n2233) );
  XNOR2_X1 U2651 ( .A(n2775), .B(n2776), .ZN(n3177) );
  AND2_X1 U2652 ( .A1(n2215), .A2(n2219), .ZN(n3695) );
  NAND2_X1 U2653 ( .A1(n2838), .A2(n2837), .ZN(n2215) );
  OAI21_X1 U2654 ( .B1(n2945), .B2(n2882), .A(n2881), .ZN(n3702) );
  INV_X1 U2655 ( .A(n3092), .ZN(n3118) );
  OR2_X1 U2656 ( .A1(n2933), .A2(n2920), .ZN(n3753) );
  NAND2_X1 U2657 ( .A1(n2221), .A2(n2220), .ZN(n3443) );
  AOI22_X1 U2658 ( .A1(n2227), .A2(n2230), .B1(n2223), .B2(n2226), .ZN(n2220)
         );
  NAND2_X1 U2659 ( .A1(n2201), .A2(n2060), .ZN(n3621) );
  NAND2_X1 U2660 ( .A1(n2214), .A2(n2213), .ZN(n3738) );
  AND2_X1 U2661 ( .A1(n2582), .A2(n2581), .ZN(n4272) );
  OR2_X1 U2662 ( .A1(n3675), .A2(n2457), .ZN(n2582) );
  OR2_X1 U2663 ( .A1(n2933), .A2(n2926), .ZN(n3751) );
  AOI21_X1 U2664 ( .B1(n3674), .B2(n3671), .A(n3672), .ZN(n3749) );
  INV_X1 U2665 ( .A(n3759), .ZN(n3775) );
  INV_X1 U2666 ( .A(n3754), .ZN(n4079) );
  NAND2_X1 U2667 ( .A1(n2591), .A2(n2590), .ZN(n4097) );
  INV_X1 U2668 ( .A(n4272), .ZN(n4112) );
  INV_X1 U2669 ( .A(n3676), .ZN(n4260) );
  INV_X1 U2670 ( .A(n4140), .ZN(n4269) );
  OAI211_X1 U2671 ( .C1(n2527), .C2(n4306), .A(n2537), .B(n2536), .ZN(n4289)
         );
  OAI211_X1 U2672 ( .C1(n4214), .C2(n2457), .A(n2529), .B(n2528), .ZN(n4222)
         );
  INV_X1 U2673 ( .A(n4323), .ZN(n3953) );
  INV_X1 U2674 ( .A(n3584), .ZN(n3955) );
  INV_X1 U2675 ( .A(n3542), .ZN(n3956) );
  NAND4_X1 U2676 ( .A1(n2453), .A2(n2452), .A3(n2451), .A4(n2450), .ZN(n3959)
         );
  INV_X1 U2677 ( .A(n3406), .ZN(n3961) );
  INV_X1 U2678 ( .A(n3354), .ZN(n3962) );
  NAND2_X1 U2679 ( .A1(n3970), .A2(n2985), .ZN(n3969) );
  AOI22_X1 U2680 ( .A1(n3063), .A2(REG2_REG_4__SCAN_IN), .B1(n4400), .B2(n2989), .ZN(n3050) );
  INV_X1 U2681 ( .A(n3046), .ZN(n2114) );
  INV_X1 U2682 ( .A(n2115), .ZN(n3047) );
  AOI22_X1 U2683 ( .A1(n3029), .A2(REG2_REG_6__SCAN_IN), .B1(n4398), .B2(n3028), .ZN(n3031) );
  NAND2_X1 U2684 ( .A1(n2159), .A2(n2157), .ZN(n4411) );
  NAND2_X1 U2685 ( .A1(n4431), .A2(n4432), .ZN(n4430) );
  XNOR2_X1 U2686 ( .A(n4019), .B(n4532), .ZN(n4445) );
  NOR2_X1 U2687 ( .A1(n4461), .A2(n4000), .ZN(n4471) );
  NAND2_X1 U2688 ( .A1(n2147), .A2(n2146), .ZN(n3999) );
  OR2_X1 U2689 ( .A1(n4452), .A2(n4448), .ZN(n2147) );
  NOR2_X1 U2690 ( .A1(n4484), .A2(REG1_REG_16__SCAN_IN), .ZN(n4485) );
  XNOR2_X1 U2691 ( .A(n4027), .B(n4026), .ZN(n4484) );
  NAND2_X1 U2692 ( .A1(n4480), .A2(n4003), .ZN(n4488) );
  INV_X1 U2693 ( .A(n2134), .ZN(n4002) );
  NAND2_X1 U2694 ( .A1(n2104), .A2(n2105), .ZN(n4106) );
  INV_X1 U2695 ( .A(n4268), .ZN(n4116) );
  NAND2_X1 U2696 ( .A1(n4283), .A2(n2556), .ZN(n4121) );
  INV_X1 U2697 ( .A(n4300), .ZN(n4193) );
  NAND2_X1 U2698 ( .A1(n2168), .A2(n2172), .ZN(n4229) );
  NAND2_X1 U2699 ( .A1(n2173), .A2(n2061), .ZN(n2168) );
  NAND2_X1 U2700 ( .A1(n3507), .A2(n3793), .ZN(n3570) );
  INV_X1 U2701 ( .A(n3685), .ZN(n4329) );
  NAND2_X1 U2702 ( .A1(n2645), .A2(n3795), .ZN(n3506) );
  AND4_X1 U2703 ( .A1(n2321), .A2(n2320), .A3(n2319), .A4(n2318), .ZN(n4334)
         );
  NAND2_X1 U2704 ( .A1(n3384), .A2(n2471), .ZN(n3490) );
  AND4_X1 U2705 ( .A1(n2464), .A2(n2463), .A3(n2462), .A4(n2461), .ZN(n3546)
         );
  OR2_X1 U2706 ( .A1(n3095), .A2(n2922), .ZN(n4511) );
  OR2_X1 U2707 ( .A1(n2527), .A2(n4563), .ZN(n2368) );
  NOR2_X1 U2708 ( .A1(n2054), .A2(n2132), .ZN(n2131) );
  OR2_X1 U2709 ( .A1(n2457), .A2(n3062), .ZN(n2369) );
  INV_X1 U2710 ( .A(n4048), .ZN(n4186) );
  AND2_X1 U2711 ( .A1(n4514), .A2(n4318), .ZN(n4185) );
  INV_X1 U2712 ( .A(n2750), .ZN(n3967) );
  OAI21_X1 U2713 ( .B1(n3619), .B2(n4315), .A(n2187), .ZN(n2727) );
  INV_X1 U2714 ( .A(REG0_REG_27__SCAN_IN), .ZN(n2128) );
  NAND2_X1 U2715 ( .A1(n2968), .A2(n2967), .ZN(n4524) );
  NAND2_X1 U2716 ( .A1(n2965), .A2(IR_REG_31__SCAN_IN), .ZN(n2297) );
  MUX2_X1 U2717 ( .A(IR_REG_31__SCAN_IN), .B(n2298), .S(IR_REG_29__SCAN_IN), 
        .Z(n2299) );
  AND2_X1 U2718 ( .A1(n2677), .A2(n2050), .ZN(n2954) );
  NAND2_X1 U2719 ( .A1(n2690), .A2(IR_REG_31__SCAN_IN), .ZN(n2682) );
  AND2_X1 U2720 ( .A1(n2972), .A2(STATE_REG_SCAN_IN), .ZN(n4525) );
  INV_X1 U2721 ( .A(n2636), .ZN(n2956) );
  XNOR2_X1 U2722 ( .A(n2631), .B(IR_REG_19__SCAN_IN), .ZN(n4395) );
  INV_X1 U2723 ( .A(n4007), .ZN(n4530) );
  INV_X1 U2724 ( .A(n4018), .ZN(n4532) );
  OR2_X1 U2725 ( .A1(n2442), .A2(n2441), .ZN(n4537) );
  AND2_X1 U2726 ( .A1(n2423), .A2(n2418), .ZN(n4397) );
  NOR2_X1 U2727 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_1__SCAN_IN), .ZN(n2356)
         );
  NAND2_X1 U2728 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2365)
         );
  INV_X1 U2729 ( .A(n2148), .ZN(n4509) );
  OAI21_X1 U2730 ( .B1(n4500), .B2(n2150), .A(n2149), .ZN(n2148) );
  OR2_X1 U2731 ( .A1(n4054), .A2(n4328), .ZN(n2715) );
  NAND2_X1 U2732 ( .A1(n2084), .A2(n2083), .ZN(U3545) );
  AOI22_X1 U2733 ( .A1(n4352), .A2(n4253), .B1(REG1_REG_27__SCAN_IN), .B2(
        n4567), .ZN(n2083) );
  NAND2_X1 U2734 ( .A1(n4350), .A2(n4569), .ZN(n2084) );
  OR2_X1 U2735 ( .A1(n4054), .A2(n4389), .ZN(n2710) );
  OAI21_X1 U2736 ( .B1(n3619), .B2(n2182), .A(n2180), .ZN(n2728) );
  AOI21_X1 U2737 ( .B1(n4352), .B2(n4351), .A(n2127), .ZN(n2126) );
  NAND2_X1 U2738 ( .A1(n4350), .A2(n4562), .ZN(n2129) );
  INV_X2 U2739 ( .A(n2360), .ZN(n2457) );
  AND2_X1 U2740 ( .A1(n2288), .A2(n2257), .ZN(n2043) );
  NAND2_X1 U2741 ( .A1(n2271), .A2(n2270), .ZN(n2386) );
  OR2_X1 U2742 ( .A1(n2654), .A2(n2111), .ZN(n2044) );
  AND4_X1 U2743 ( .A1(n2388), .A2(n4655), .A3(n2416), .A4(n4693), .ZN(n2045)
         );
  AND2_X1 U2744 ( .A1(n2793), .A2(n3186), .ZN(n2046) );
  INV_X1 U2745 ( .A(n2734), .ZN(n2366) );
  OR2_X1 U2746 ( .A1(n3649), .A2(n2210), .ZN(n2047) );
  NAND2_X1 U2747 ( .A1(n2202), .A2(n3186), .ZN(n3314) );
  INV_X1 U2748 ( .A(n3786), .ZN(n2089) );
  AND2_X1 U2749 ( .A1(n2159), .A2(n2161), .ZN(n2048) );
  INV_X1 U2750 ( .A(n4026), .ZN(n2133) );
  INV_X1 U2751 ( .A(n2901), .ZN(n2759) );
  NOR2_X1 U2752 ( .A1(n4082), .A2(n4061), .ZN(n2049) );
  AND4_X1 U2753 ( .A1(n2355), .A2(n2354), .A3(n2353), .A4(n2352), .ZN(n2750)
         );
  NAND2_X1 U2754 ( .A1(n2289), .A2(n2043), .ZN(n2050) );
  OR3_X1 U2755 ( .A1(n4082), .A2(n4061), .A3(n2096), .ZN(n2051) );
  XNOR2_X1 U2756 ( .A(n2634), .B(n2633), .ZN(n2636) );
  NAND2_X1 U2757 ( .A1(n3716), .A2(n3289), .ZN(n2052) );
  AND2_X1 U2758 ( .A1(n2962), .A2(n2960), .ZN(n2360) );
  AND2_X1 U2759 ( .A1(n2351), .A2(n2350), .ZN(n4401) );
  AND2_X1 U2760 ( .A1(n2943), .A2(n2877), .ZN(n2945) );
  AND2_X1 U2761 ( .A1(n2299), .A2(n2965), .ZN(n2960) );
  AND2_X1 U2762 ( .A1(n2105), .A2(n2103), .ZN(n2053) );
  AND2_X1 U2763 ( .A1(n2361), .A2(REG2_REG_0__SCAN_IN), .ZN(n2054) );
  AND2_X1 U2764 ( .A1(n4399), .A2(REG1_REG_5__SCAN_IN), .ZN(n2055) );
  AND2_X1 U2765 ( .A1(n2271), .A2(n2270), .ZN(n2197) );
  OR2_X1 U2766 ( .A1(n2945), .A2(n2241), .ZN(n2056) );
  AND2_X1 U2767 ( .A1(n2136), .A2(n4401), .ZN(n2057) );
  NAND2_X1 U2768 ( .A1(n3960), .A2(n3403), .ZN(n2058) );
  INV_X1 U2769 ( .A(IR_REG_27__SCAN_IN), .ZN(n2290) );
  NAND2_X1 U2770 ( .A1(n3953), .A2(n3685), .ZN(n2059) );
  XNOR2_X1 U2771 ( .A(n2682), .B(IR_REG_24__SCAN_IN), .ZN(n2686) );
  INV_X1 U2772 ( .A(n3415), .ZN(n2224) );
  INV_X1 U2773 ( .A(n2886), .ZN(n2919) );
  OR2_X1 U2774 ( .A1(n2871), .A2(n3659), .ZN(n2060) );
  AND2_X1 U2775 ( .A1(n2507), .A2(n2059), .ZN(n2061) );
  AND2_X1 U2776 ( .A1(n2213), .A2(n2217), .ZN(n2062) );
  NAND2_X1 U2777 ( .A1(n2251), .A2(n2249), .ZN(n3341) );
  OR2_X1 U2778 ( .A1(n3754), .A2(n4247), .ZN(n2063) );
  OR2_X1 U2779 ( .A1(n3660), .A2(n2870), .ZN(n2064) );
  OAI21_X1 U2780 ( .B1(n3443), .B2(n3444), .A(n3445), .ZN(n3520) );
  AND2_X1 U2781 ( .A1(n2173), .A2(n2059), .ZN(n2065) );
  INV_X1 U2782 ( .A(n3914), .ZN(n2111) );
  AND2_X1 U2783 ( .A1(n2245), .A2(n2234), .ZN(n2066) );
  INV_X1 U2784 ( .A(n3879), .ZN(n2106) );
  AND2_X1 U2785 ( .A1(n3693), .A2(n3692), .ZN(n2067) );
  INV_X1 U2786 ( .A(n3671), .ZN(n2246) );
  NAND2_X1 U2787 ( .A1(n2081), .A2(n2169), .ZN(n4227) );
  INV_X1 U2788 ( .A(n3526), .ZN(n3557) );
  INV_X1 U2789 ( .A(n2090), .ZN(n4146) );
  NOR3_X1 U2790 ( .A1(n4210), .A2(n2094), .A3(n4184), .ZN(n2090) );
  NOR2_X1 U2791 ( .A1(n4210), .A2(n2091), .ZN(n2095) );
  INV_X1 U2792 ( .A(n2556), .ZN(n2166) );
  AND2_X1 U2793 ( .A1(n2064), .A2(n3728), .ZN(n2068) );
  NAND2_X1 U2794 ( .A1(n2621), .A2(IR_REG_31__SCAN_IN), .ZN(n2631) );
  INV_X1 U2795 ( .A(n4206), .ZN(n4320) );
  AND3_X1 U2796 ( .A1(n2518), .A2(n2517), .A3(n2516), .ZN(n4206) );
  INV_X1 U2797 ( .A(n2172), .ZN(n2171) );
  NAND2_X1 U2798 ( .A1(n2070), .A2(n2507), .ZN(n2172) );
  INV_X1 U2799 ( .A(n2268), .ZN(n2167) );
  AND2_X1 U2800 ( .A1(n4009), .A2(REG2_REG_9__SCAN_IN), .ZN(n2069) );
  INV_X1 U2801 ( .A(n3672), .ZN(n2247) );
  NOR2_X1 U2802 ( .A1(n2506), .A2(n4317), .ZN(n2070) );
  OR2_X1 U2803 ( .A1(n2216), .A2(n2067), .ZN(n2071) );
  OR2_X1 U2804 ( .A1(n2227), .A2(n2223), .ZN(n2072) );
  OR2_X1 U2805 ( .A1(n4334), .A2(n3515), .ZN(n2073) );
  NAND2_X1 U2806 ( .A1(n3676), .A2(n4116), .ZN(n2074) );
  INV_X1 U2807 ( .A(n2471), .ZN(n2192) );
  AND2_X1 U2808 ( .A1(n2232), .A2(n2243), .ZN(n2075) );
  AND2_X1 U2809 ( .A1(n2873), .A2(n2060), .ZN(n2076) );
  INV_X1 U2810 ( .A(IR_REG_28__SCAN_IN), .ZN(n2296) );
  NAND2_X1 U2811 ( .A1(n2372), .A2(n2373), .ZN(n3146) );
  AND2_X1 U2812 ( .A1(n2178), .A2(n2179), .ZN(n3205) );
  NAND2_X1 U2813 ( .A1(n2251), .A2(n2252), .ZN(n3340) );
  AND2_X1 U2814 ( .A1(n2846), .A2(n2845), .ZN(n2077) );
  NAND2_X1 U2815 ( .A1(n3802), .A2(n3806), .ZN(n2637) );
  INV_X1 U2816 ( .A(n4022), .ZN(n2145) );
  AND2_X1 U2817 ( .A1(n2145), .A2(n2144), .ZN(n2078) );
  INV_X1 U2818 ( .A(n2219), .ZN(n2216) );
  NAND2_X1 U2819 ( .A1(n2836), .A2(n2835), .ZN(n2219) );
  AND4_X1 U2820 ( .A1(n2254), .A2(n2364), .A3(n2362), .A4(n2363), .ZN(n2730)
         );
  NAND2_X1 U2821 ( .A1(n3228), .A2(n4540), .ZN(n4554) );
  INV_X1 U2822 ( .A(n2292), .ZN(n2664) );
  INV_X1 U2823 ( .A(n2161), .ZN(n2160) );
  INV_X1 U2824 ( .A(n4029), .ZN(n4528) );
  INV_X1 U2825 ( .A(IR_REG_0__SCAN_IN), .ZN(n2101) );
  NAND2_X1 U2826 ( .A1(n4396), .A2(n4513), .ZN(n2161) );
  INV_X1 U2827 ( .A(n4396), .ZN(n2099) );
  XNOR2_X1 U2828 ( .A(n3992), .B(n4396), .ZN(n3993) );
  NAND2_X1 U2829 ( .A1(n2637), .A2(n3108), .ZN(n3110) );
  INV_X1 U2830 ( .A(n3147), .ZN(n2372) );
  NAND2_X1 U2831 ( .A1(n4227), .A2(n2523), .ZN(n4176) );
  AND4_X2 U2832 ( .A1(n2197), .A2(n2281), .A3(n2287), .A4(n2045), .ZN(n2289)
         );
  INV_X1 U2833 ( .A(n2289), .ZN(n2678) );
  NAND2_X1 U2834 ( .A1(n2666), .A2(IR_REG_31__SCAN_IN), .ZN(n2298) );
  AND2_X2 U2835 ( .A1(n2088), .A2(n2087), .ZN(n2734) );
  INV_X1 U2836 ( .A(n2095), .ZN(n4131) );
  INV_X1 U2837 ( .A(n2271), .ZN(n2341) );
  INV_X1 U2838 ( .A(n2637), .ZN(n2112) );
  NOR2_X2 U2839 ( .A1(n3045), .A2(n2055), .ZN(n3032) );
  OAI21_X1 U2840 ( .B1(n2645), .B2(n2122), .A(n2119), .ZN(n3569) );
  NAND2_X1 U2841 ( .A1(n2129), .A2(n2126), .ZN(U3513) );
  NOR2_X1 U2842 ( .A1(n4562), .A2(n2128), .ZN(n2127) );
  NAND3_X1 U2843 ( .A1(n2369), .A2(n2368), .A3(n2131), .ZN(n2737) );
  AOI21_X1 U2844 ( .B1(n4452), .B2(n2143), .A(n2140), .ZN(n2139) );
  OAI21_X1 U2845 ( .B1(n3992), .B2(n2156), .A(n2154), .ZN(n3994) );
  AOI21_X1 U2846 ( .B1(n3138), .B2(n3137), .A(n3136), .ZN(n4011) );
  OAI21_X1 U2847 ( .B1(n4090), .B2(n2656), .A(n3852), .ZN(n4067) );
  OAI21_X2 U2848 ( .B1(n3328), .B2(n3836), .A(n3822), .ZN(n3370) );
  INV_X1 U2849 ( .A(n3571), .ZN(n2173) );
  NAND2_X1 U2850 ( .A1(n3382), .A2(n2471), .ZN(n2189) );
  NAND2_X1 U2851 ( .A1(n2189), .A2(n2190), .ZN(n2483) );
  AND2_X1 U2852 ( .A1(n2197), .A2(n2045), .ZN(n2282) );
  NAND2_X1 U2853 ( .A1(n2201), .A2(n2076), .ZN(n2943) );
  NAND2_X1 U2854 ( .A1(n3725), .A2(n3728), .ZN(n3658) );
  NAND2_X1 U2855 ( .A1(n2202), .A2(n2046), .ZN(n3315) );
  NAND2_X1 U2856 ( .A1(n2779), .A2(n2778), .ZN(n3184) );
  INV_X1 U2857 ( .A(n2778), .ZN(n2204) );
  NAND2_X1 U2858 ( .A1(n2205), .A2(n2208), .ZN(n3726) );
  NAND3_X1 U2859 ( .A1(n2838), .A2(n2206), .A3(n2837), .ZN(n2205) );
  NAND3_X1 U2860 ( .A1(n2838), .A2(n2837), .A3(n2218), .ZN(n2214) );
  NAND2_X1 U2861 ( .A1(n3393), .A2(n2072), .ZN(n2221) );
  AOI21_X1 U2862 ( .B1(n3395), .B2(n2229), .A(n2228), .ZN(n2227) );
  INV_X1 U2863 ( .A(n3414), .ZN(n2228) );
  NOR2_X1 U2864 ( .A1(n3394), .A2(n3415), .ZN(n2229) );
  NAND2_X1 U2865 ( .A1(n3395), .A2(n2224), .ZN(n2230) );
  NAND2_X1 U2866 ( .A1(n2945), .A2(n2066), .ZN(n2231) );
  NAND2_X1 U2867 ( .A1(n2231), .A2(n2075), .ZN(n3633) );
  INV_X1 U2868 ( .A(n2881), .ZN(n2248) );
  NAND2_X1 U2869 ( .A1(n2289), .A2(n2288), .ZN(n2675) );
  NAND2_X1 U2870 ( .A1(n2260), .A2(n2261), .ZN(n2832) );
  NAND2_X1 U2871 ( .A1(n2370), .A2(n2734), .ZN(n3802) );
  OAI22_X2 U2872 ( .A1(n3371), .A2(n2455), .B1(n3332), .B2(n3423), .ZN(n3382)
         );
  XNOR2_X1 U2873 ( .A(n2733), .B(n2896), .ZN(n2745) );
  AND2_X1 U2874 ( .A1(n2553), .A2(n2552), .ZN(n4292) );
  OR2_X1 U2875 ( .A1(n3458), .A2(n3541), .ZN(n2264) );
  AND4_X1 U2876 ( .A1(n2503), .A2(n2502), .A3(n2501), .A4(n2500), .ZN(n4332)
         );
  INV_X1 U2877 ( .A(n4332), .ZN(n2506) );
  INV_X1 U2878 ( .A(n3458), .ZN(n3957) );
  AND4_X1 U2879 ( .A1(n2478), .A2(n2477), .A3(n2476), .A4(n2475), .ZN(n3458)
         );
  OR2_X2 U2880 ( .A1(n2901), .A2(n4231), .ZN(n2765) );
  OR2_X1 U2881 ( .A1(n2942), .A2(n4563), .ZN(n2265) );
  OR2_X1 U2882 ( .A1(n3608), .A2(n4328), .ZN(n2266) );
  OR2_X1 U2883 ( .A1(n3608), .A2(n4389), .ZN(n2267) );
  AND2_X2 U2884 ( .A1(n2712), .A2(n2909), .ZN(n4569) );
  AND2_X2 U2885 ( .A1(n2712), .A2(n3099), .ZN(n4562) );
  NAND2_X1 U2886 ( .A1(n2757), .A2(n2756), .ZN(n3076) );
  AND2_X1 U2887 ( .A1(n4269), .A2(n2708), .ZN(n2268) );
  OR2_X1 U2888 ( .A1(n2791), .A2(n3156), .ZN(n2269) );
  NAND2_X1 U2889 ( .A1(n3966), .A2(n2783), .ZN(n2761) );
  INV_X1 U2890 ( .A(n3317), .ZN(n2793) );
  INV_X1 U2891 ( .A(n4221), .ZN(n2522) );
  AND2_X1 U2892 ( .A1(n3208), .A2(n3161), .ZN(n2358) );
  NOR2_X1 U2893 ( .A1(n2947), .A2(n2944), .ZN(n2877) );
  NOR2_X1 U2894 ( .A1(n2497), .A2(n2496), .ZN(n2512) );
  INV_X1 U2895 ( .A(n2576), .ZN(n2575) );
  INV_X1 U2896 ( .A(n2960), .ZN(n2300) );
  NAND2_X1 U2897 ( .A1(n4206), .A2(n2522), .ZN(n2523) );
  AND2_X1 U2898 ( .A1(REG3_REG_8__SCAN_IN), .A2(REG3_REG_9__SCAN_IN), .ZN(
        n2301) );
  INV_X1 U2899 ( .A(IR_REG_17__SCAN_IN), .ZN(n2519) );
  INV_X1 U2900 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4681) );
  AND2_X1 U2901 ( .A1(n2333), .A2(REG3_REG_5__SCAN_IN), .ZN(n2377) );
  NAND2_X1 U2902 ( .A1(n3315), .A2(n2796), .ZN(n3297) );
  OR2_X1 U2903 ( .A1(n2854), .A2(n2853), .ZN(n2855) );
  OR2_X1 U2904 ( .A1(n2486), .A2(n2315), .ZN(n2317) );
  AND2_X2 U2905 ( .A1(n2962), .A2(n2300), .ZN(n2361) );
  AND2_X1 U2906 ( .A1(n2742), .A2(n2265), .ZN(n2735) );
  NAND2_X1 U2907 ( .A1(n4161), .A2(n2555), .ZN(n2556) );
  OR2_X1 U2908 ( .A1(n3955), .A2(n3526), .ZN(n2494) );
  INV_X1 U2909 ( .A(n3881), .ZN(n2470) );
  NAND2_X1 U2910 ( .A1(n2302), .A2(n2301), .ZN(n2447) );
  INV_X1 U2911 ( .A(n3603), .ZN(n4317) );
  OR3_X1 U2912 ( .A1(n2465), .A2(IR_REG_12__SCAN_IN), .A3(n2273), .ZN(n2322)
         );
  NAND2_X1 U2913 ( .A1(n2409), .A2(REG3_REG_7__SCAN_IN), .ZN(n2432) );
  NAND2_X1 U2914 ( .A1(n2557), .A2(REG3_REG_23__SCAN_IN), .ZN(n2566) );
  AND2_X1 U2915 ( .A1(n2524), .A2(REG3_REG_19__SCAN_IN), .ZN(n2533) );
  OR2_X1 U2916 ( .A1(n2754), .A2(n2753), .ZN(n2755) );
  OR2_X1 U2917 ( .A1(n2968), .A2(D_REG_1__SCAN_IN), .ZN(n3096) );
  OR2_X1 U2918 ( .A1(n3609), .A2(n2457), .ZN(n2612) );
  NAND2_X1 U2919 ( .A1(n2736), .A2(n2735), .ZN(n3006) );
  INV_X1 U2920 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4605) );
  OR2_X1 U2921 ( .A1(n2605), .A2(n2927), .ZN(n4053) );
  AND2_X1 U2922 ( .A1(n2646), .A2(n4202), .ZN(n4173) );
  INV_X1 U2923 ( .A(n4185), .ZN(n4166) );
  INV_X1 U2924 ( .A(n4331), .ZN(n4319) );
  OR2_X1 U2925 ( .A1(n2968), .A2(D_REG_0__SCAN_IN), .ZN(n2707) );
  INV_X1 U2926 ( .A(n4132), .ZN(n2708) );
  INV_X1 U2927 ( .A(n2555), .ZN(n4144) );
  INV_X1 U2928 ( .A(n3541), .ZN(n3497) );
  OR2_X1 U2929 ( .A1(n2968), .A2(n2703), .ZN(n2908) );
  INV_X1 U2930 ( .A(n3753), .ZN(n3766) );
  INV_X1 U2931 ( .A(n3751), .ZN(n3769) );
  NAND2_X1 U2932 ( .A1(n2533), .A2(REG3_REG_20__SCAN_IN), .ZN(n2547) );
  AND2_X1 U2933 ( .A1(n2596), .A2(n2586), .ZN(n4084) );
  AND2_X1 U2934 ( .A1(n2612), .A2(n2611), .ZN(n4049) );
  AND2_X1 U2935 ( .A1(n2564), .A2(n2563), .ZN(n4140) );
  AND4_X1 U2936 ( .A1(n2309), .A2(n2308), .A3(n2307), .A4(n2306), .ZN(n4323)
         );
  AND2_X1 U2937 ( .A1(n2976), .A2(n2975), .ZN(n2991) );
  AND2_X1 U2938 ( .A1(n2991), .A2(n3944), .ZN(n4450) );
  AND2_X1 U2939 ( .A1(n3782), .A2(n3780), .ZN(n3905) );
  NAND2_X1 U2940 ( .A1(n2644), .A2(n3797), .ZN(n3908) );
  INV_X1 U2941 ( .A(n4218), .ZN(n4237) );
  INV_X1 U2942 ( .A(n4213), .ZN(n4517) );
  AND2_X1 U2943 ( .A1(n2707), .A2(n2706), .ZN(n2909) );
  INV_X1 U2944 ( .A(n4389), .ZN(n4351) );
  AND2_X1 U2945 ( .A1(n3943), .A2(n2731), .ZN(n4552) );
  XNOR2_X1 U2946 ( .A(n2629), .B(n2622), .ZN(n2691) );
  AND2_X1 U2947 ( .A1(n2469), .A2(n2479), .ZN(n4533) );
  AND2_X1 U2948 ( .A1(n2976), .A2(n2974), .ZN(n4503) );
  NOR2_X1 U2949 ( .A1(n2938), .A2(n2937), .ZN(n2939) );
  AND2_X1 U2950 ( .A1(n2934), .A2(n3056), .ZN(n3773) );
  OR2_X1 U2951 ( .A1(n2933), .A2(n2914), .ZN(n3759) );
  INV_X1 U2952 ( .A(n4049), .ZN(n4250) );
  NAND2_X1 U2953 ( .A1(n2544), .A2(n2543), .ZN(n4300) );
  INV_X1 U2954 ( .A(n4334), .ZN(n3954) );
  INV_X1 U2955 ( .A(n4450), .ZN(n4499) );
  OR2_X1 U2956 ( .A1(n4233), .A2(n4547), .ZN(n4213) );
  AND2_X1 U2957 ( .A1(n2715), .A2(n2714), .ZN(n2716) );
  NAND2_X1 U2958 ( .A1(n4569), .A2(n4231), .ZN(n4328) );
  INV_X1 U2959 ( .A(n4569), .ZN(n4567) );
  AND2_X1 U2960 ( .A1(n2710), .A2(n2709), .ZN(n2711) );
  NAND2_X1 U2961 ( .A1(n4562), .A2(n4231), .ZN(n4389) );
  INV_X1 U2962 ( .A(n4562), .ZN(n4560) );
  INV_X1 U2963 ( .A(n2686), .ZN(n3629) );
  INV_X1 U2964 ( .A(n4008), .ZN(n4531) );
  AND2_X1 U2965 ( .A1(n2406), .A2(n2415), .ZN(n4398) );
  NAND2_X1 U2966 ( .A1(n2282), .A2(n2272), .ZN(n2465) );
  INV_X1 U2967 ( .A(n2280), .ZN(n2273) );
  NOR2_X1 U2968 ( .A1(n2322), .A2(IR_REG_13__SCAN_IN), .ZN(n2492) );
  INV_X1 U2969 ( .A(IR_REG_14__SCAN_IN), .ZN(n2274) );
  NAND2_X1 U2970 ( .A1(n2492), .A2(n2274), .ZN(n2275) );
  NAND2_X1 U2971 ( .A1(n2275), .A2(IR_REG_31__SCAN_IN), .ZN(n2311) );
  INV_X1 U2972 ( .A(IR_REG_15__SCAN_IN), .ZN(n2310) );
  NAND2_X1 U2973 ( .A1(n2311), .A2(n2310), .ZN(n2313) );
  NAND2_X1 U2974 ( .A1(n2313), .A2(IR_REG_31__SCAN_IN), .ZN(n2276) );
  XNOR2_X1 U2975 ( .A(n2276), .B(IR_REG_16__SCAN_IN), .ZN(n4026) );
  NAND2_X1 U2976 ( .A1(n2290), .A2(n2964), .ZN(n2291) );
  NAND2_X1 U2977 ( .A1(n2663), .A2(n2296), .ZN(n2295) );
  NAND2_X4 U2978 ( .A1(n2295), .A2(n2294), .ZN(n3786) );
  MUX2_X1 U2979 ( .A(DATAI_16_), .B(n4026), .S(n2042), .Z(n3685) );
  NAND2_X1 U2980 ( .A1(n3783), .A2(REG0_REG_16__SCAN_IN), .ZN(n2309) );
  INV_X1 U2981 ( .A(n2361), .ZN(n2343) );
  OR2_X1 U2982 ( .A1(n2343), .A2(n4479), .ZN(n2308) );
  INV_X1 U2983 ( .A(REG3_REG_15__SCAN_IN), .ZN(n2315) );
  NAND2_X1 U2984 ( .A1(n2317), .A2(n4605), .ZN(n2304) );
  NAND2_X1 U2985 ( .A1(n2497), .A2(n2304), .ZN(n3688) );
  OR2_X1 U2986 ( .A1(n2457), .A2(n3688), .ZN(n2307) );
  INV_X1 U2987 ( .A(REG1_REG_16__SCAN_IN), .ZN(n2305) );
  OR2_X1 U2988 ( .A1(n2527), .A2(n2305), .ZN(n2306) );
  INV_X1 U2989 ( .A(DATAI_15_), .ZN(n4672) );
  OR2_X1 U2990 ( .A1(n2311), .A2(n2310), .ZN(n2312) );
  MUX2_X1 U2991 ( .A(n4672), .B(n4530), .S(n3786), .Z(n3515) );
  NAND2_X1 U2992 ( .A1(n3783), .A2(REG0_REG_15__SCAN_IN), .ZN(n2321) );
  INV_X1 U2993 ( .A(REG2_REG_15__SCAN_IN), .ZN(n2314) );
  OR2_X1 U2994 ( .A1(n2343), .A2(n2314), .ZN(n2320) );
  NAND2_X1 U2995 ( .A1(n2486), .A2(n2315), .ZN(n2316) );
  NAND2_X1 U2996 ( .A1(n2317), .A2(n2316), .ZN(n3772) );
  OR2_X1 U2997 ( .A1(n2457), .A2(n3772), .ZN(n2319) );
  INV_X1 U2998 ( .A(REG1_REG_15__SCAN_IN), .ZN(n3587) );
  OR2_X1 U2999 ( .A1(n2527), .A2(n3587), .ZN(n2318) );
  INV_X1 U3000 ( .A(DATAI_13_), .ZN(n4691) );
  NAND2_X1 U3001 ( .A1(n2322), .A2(IR_REG_31__SCAN_IN), .ZN(n2323) );
  XNOR2_X1 U3002 ( .A(n2323), .B(IR_REG_13__SCAN_IN), .ZN(n4008) );
  MUX2_X1 U3003 ( .A(n4691), .B(n4531), .S(n2042), .Z(n3478) );
  INV_X1 U3004 ( .A(n3478), .ZN(n3448) );
  NAND2_X1 U3005 ( .A1(n3783), .A2(REG0_REG_13__SCAN_IN), .ZN(n2331) );
  INV_X1 U3006 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4449) );
  OR2_X1 U3007 ( .A1(n2343), .A2(n4449), .ZN(n2330) );
  INV_X1 U3008 ( .A(n2324), .ZN(n2484) );
  INV_X1 U3009 ( .A(n2325), .ZN(n2474) );
  INV_X1 U3010 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2326) );
  NAND2_X1 U3011 ( .A1(n2474), .A2(n2326), .ZN(n2327) );
  NAND2_X1 U3012 ( .A1(n2484), .A2(n2327), .ZN(n3481) );
  OR2_X1 U3013 ( .A1(n2457), .A2(n3481), .ZN(n2329) );
  INV_X1 U3014 ( .A(REG1_REG_13__SCAN_IN), .ZN(n3535) );
  OR2_X1 U3015 ( .A1(n2527), .A2(n3535), .ZN(n2328) );
  INV_X1 U3016 ( .A(REG1_REG_4__SCAN_IN), .ZN(n2332) );
  OR2_X1 U3017 ( .A1(n2527), .A2(n2332), .ZN(n2340) );
  INV_X1 U3018 ( .A(n2333), .ZN(n2379) );
  INV_X1 U3019 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2334) );
  INV_X1 U3020 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3123) );
  NAND2_X1 U3021 ( .A1(n2334), .A2(n3123), .ZN(n2335) );
  NAND2_X1 U3022 ( .A1(n2379), .A2(n2335), .ZN(n3719) );
  NAND2_X1 U3023 ( .A1(n2361), .A2(REG2_REG_4__SCAN_IN), .ZN(n2338) );
  INV_X1 U3024 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2336) );
  OR2_X1 U3025 ( .A1(n2509), .A2(n2336), .ZN(n2337) );
  NAND2_X1 U3026 ( .A1(n2341), .A2(IR_REG_31__SCAN_IN), .ZN(n2349) );
  NAND2_X1 U3027 ( .A1(n2349), .A2(n4626), .ZN(n2351) );
  NAND2_X1 U3028 ( .A1(n2351), .A2(IR_REG_31__SCAN_IN), .ZN(n2342) );
  XNOR2_X1 U3029 ( .A(n2342), .B(IR_REG_4__SCAN_IN), .ZN(n4400) );
  MUX2_X1 U3030 ( .A(DATAI_4_), .B(n4400), .S(n3786), .Z(n3718) );
  INV_X1 U3031 ( .A(n3718), .ZN(n3218) );
  NAND2_X1 U3032 ( .A1(n3965), .A2(n3218), .ZN(n3816) );
  NAND2_X1 U3033 ( .A1(n3813), .A2(n3816), .ZN(n2374) );
  INV_X1 U3034 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3982) );
  OR2_X1 U3035 ( .A1(n2343), .A2(n3982), .ZN(n2348) );
  NAND2_X1 U3036 ( .A1(n3783), .A2(REG0_REG_3__SCAN_IN), .ZN(n2346) );
  OR2_X1 U3037 ( .A1(n2457), .A2(REG3_REG_3__SCAN_IN), .ZN(n2345) );
  INV_X1 U3038 ( .A(REG1_REG_3__SCAN_IN), .ZN(n3172) );
  OR2_X1 U3039 ( .A1(n2527), .A2(n3172), .ZN(n2344) );
  INV_X1 U3040 ( .A(n3966), .ZN(n3079) );
  OR2_X1 U3041 ( .A1(n2349), .A2(n4626), .ZN(n2350) );
  MUX2_X1 U3042 ( .A(DATAI_3_), .B(n4401), .S(n3786), .Z(n3165) );
  NAND2_X1 U3043 ( .A1(n3079), .A2(n3260), .ZN(n3208) );
  INV_X1 U3044 ( .A(REG1_REG_2__SCAN_IN), .ZN(n2993) );
  OR2_X1 U3045 ( .A1(n2527), .A2(n2993), .ZN(n2354) );
  NAND2_X1 U3046 ( .A1(n2360), .A2(REG3_REG_2__SCAN_IN), .ZN(n2353) );
  NAND2_X1 U3047 ( .A1(n2361), .A2(REG2_REG_2__SCAN_IN), .ZN(n2352) );
  OR2_X1 U3048 ( .A1(n2356), .A2(n2964), .ZN(n2357) );
  MUX2_X1 U3049 ( .A(DATAI_2_), .B(n4402), .S(n3786), .Z(n3268) );
  INV_X1 U3050 ( .A(n3268), .ZN(n3156) );
  NAND2_X1 U3051 ( .A1(n2750), .A2(n3156), .ZN(n3161) );
  NAND2_X1 U3052 ( .A1(n2750), .A2(n3268), .ZN(n3807) );
  NAND2_X1 U3053 ( .A1(n3967), .A2(n3156), .ZN(n3810) );
  AND2_X2 U3054 ( .A1(n3807), .A2(n3810), .ZN(n3880) );
  INV_X1 U3055 ( .A(n3880), .ZN(n2373) );
  INV_X1 U3056 ( .A(REG1_REG_1__SCAN_IN), .ZN(n2359) );
  NAND2_X1 U3057 ( .A1(n2360), .A2(REG3_REG_1__SCAN_IN), .ZN(n2363) );
  NAND2_X1 U3058 ( .A1(n2361), .A2(REG2_REG_1__SCAN_IN), .ZN(n2362) );
  XNOR2_X2 U3059 ( .A(n2365), .B(IR_REG_1__SCAN_IN), .ZN(n4403) );
  INV_X1 U3060 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3062) );
  INV_X1 U3061 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2367) );
  INV_X1 U3062 ( .A(REG1_REG_0__SCAN_IN), .ZN(n4563) );
  AND2_X1 U3063 ( .A1(n2737), .A2(n3118), .ZN(n3108) );
  NAND2_X1 U3064 ( .A1(n2370), .A2(n2366), .ZN(n2371) );
  INV_X1 U3065 ( .A(n2374), .ZN(n2375) );
  NAND2_X1 U3066 ( .A1(n3966), .A2(n3165), .ZN(n3206) );
  NAND2_X1 U3067 ( .A1(n3965), .A2(n3718), .ZN(n3225) );
  NAND2_X1 U3068 ( .A1(n3783), .A2(REG0_REG_5__SCAN_IN), .ZN(n2385) );
  INV_X1 U3069 ( .A(REG1_REG_5__SCAN_IN), .ZN(n3313) );
  OR2_X1 U3070 ( .A1(n2527), .A2(n3313), .ZN(n2384) );
  INV_X1 U3071 ( .A(n2377), .ZN(n2395) );
  INV_X1 U3072 ( .A(REG3_REG_5__SCAN_IN), .ZN(n2378) );
  NAND2_X1 U3073 ( .A1(n2379), .A2(n2378), .ZN(n2380) );
  NAND2_X1 U3074 ( .A1(n2395), .A2(n2380), .ZN(n3233) );
  OR2_X1 U3075 ( .A1(n2457), .A2(n3233), .ZN(n2383) );
  INV_X1 U3076 ( .A(REG2_REG_5__SCAN_IN), .ZN(n2381) );
  OR2_X1 U3077 ( .A1(n2343), .A2(n2381), .ZN(n2382) );
  INV_X1 U3078 ( .A(n3716), .ZN(n3964) );
  INV_X1 U3079 ( .A(DATAI_5_), .ZN(n2390) );
  NAND2_X1 U3080 ( .A1(n2386), .A2(IR_REG_31__SCAN_IN), .ZN(n2387) );
  MUX2_X1 U3081 ( .A(n2387), .B(IR_REG_31__SCAN_IN), .S(n2388), .Z(n2389) );
  NAND2_X1 U3082 ( .A1(n2197), .A2(n2388), .ZN(n2404) );
  NAND2_X1 U3083 ( .A1(n2389), .A2(n2404), .ZN(n3052) );
  MUX2_X1 U3084 ( .A(n2390), .B(n3052), .S(n3786), .Z(n3289) );
  NAND2_X1 U3085 ( .A1(n3964), .A2(n3230), .ZN(n2391) );
  AND2_X1 U3086 ( .A1(n3225), .A2(n2391), .ZN(n2392) );
  NAND2_X1 U3087 ( .A1(n2361), .A2(REG2_REG_6__SCAN_IN), .ZN(n2402) );
  INV_X1 U3088 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2393) );
  OR2_X1 U3089 ( .A1(n2509), .A2(n2393), .ZN(n2401) );
  INV_X1 U3090 ( .A(n2409), .ZN(n2397) );
  INV_X1 U3091 ( .A(REG3_REG_6__SCAN_IN), .ZN(n2394) );
  NAND2_X1 U3092 ( .A1(n2395), .A2(n2394), .ZN(n2396) );
  NAND2_X1 U3093 ( .A1(n2397), .A2(n2396), .ZN(n3251) );
  OR2_X1 U3094 ( .A1(n2457), .A2(n3251), .ZN(n2400) );
  INV_X1 U3095 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2398) );
  OR2_X1 U3096 ( .A1(n2527), .A2(n2398), .ZN(n2399) );
  NAND4_X1 U3097 ( .A1(n2402), .A2(n2401), .A3(n2400), .A4(n2399), .ZN(n3963)
         );
  NAND2_X1 U3098 ( .A1(n2404), .A2(IR_REG_31__SCAN_IN), .ZN(n2403) );
  MUX2_X1 U3099 ( .A(n2403), .B(IR_REG_31__SCAN_IN), .S(n4693), .Z(n2406) );
  INV_X1 U3100 ( .A(n2404), .ZN(n2405) );
  NAND2_X1 U3101 ( .A1(n2405), .A2(n4693), .ZN(n2415) );
  MUX2_X1 U3102 ( .A(DATAI_6_), .B(n4398), .S(n3786), .Z(n3191) );
  AND2_X1 U3103 ( .A1(n3963), .A2(n3191), .ZN(n2407) );
  NAND2_X1 U3104 ( .A1(n3783), .A2(REG0_REG_7__SCAN_IN), .ZN(n2414) );
  INV_X1 U3105 ( .A(REG2_REG_7__SCAN_IN), .ZN(n2408) );
  OR2_X1 U3106 ( .A1(n2343), .A2(n2408), .ZN(n2413) );
  OAI21_X1 U3107 ( .B1(n2409), .B2(REG3_REG_7__SCAN_IN), .A(n2432), .ZN(n3324)
         );
  OR2_X1 U3108 ( .A1(n2457), .A2(n3324), .ZN(n2412) );
  INV_X1 U3109 ( .A(REG1_REG_7__SCAN_IN), .ZN(n2410) );
  OR2_X1 U3110 ( .A1(n2527), .A2(n2410), .ZN(n2411) );
  NAND2_X1 U3111 ( .A1(n2415), .A2(IR_REG_31__SCAN_IN), .ZN(n2417) );
  NAND2_X1 U3112 ( .A1(n2417), .A2(n2416), .ZN(n2423) );
  OR2_X1 U3113 ( .A1(n2417), .A2(n2416), .ZN(n2418) );
  MUX2_X1 U3114 ( .A(DATAI_7_), .B(n4397), .S(n3786), .Z(n3321) );
  NAND2_X1 U3115 ( .A1(n3354), .A2(n3321), .ZN(n2639) );
  INV_X1 U3116 ( .A(n3321), .ZN(n2792) );
  NAND2_X1 U3117 ( .A1(n3962), .A2(n2792), .ZN(n3823) );
  NAND2_X1 U3118 ( .A1(n3783), .A2(REG0_REG_8__SCAN_IN), .ZN(n2422) );
  INV_X1 U3119 ( .A(REG1_REG_8__SCAN_IN), .ZN(n4012) );
  OR2_X1 U3120 ( .A1(n2527), .A2(n4012), .ZN(n2421) );
  INV_X1 U3121 ( .A(REG3_REG_8__SCAN_IN), .ZN(n2431) );
  XNOR2_X1 U3122 ( .A(n2432), .B(n2431), .ZN(n4512) );
  OR2_X1 U3123 ( .A1(n2457), .A2(n4512), .ZN(n2420) );
  INV_X1 U3124 ( .A(REG2_REG_8__SCAN_IN), .ZN(n4513) );
  OR2_X1 U3125 ( .A1(n2343), .A2(n4513), .ZN(n2419) );
  INV_X1 U3126 ( .A(DATAI_8_), .ZN(n2425) );
  NAND2_X1 U3127 ( .A1(n2423), .A2(IR_REG_31__SCAN_IN), .ZN(n2424) );
  XNOR2_X1 U3128 ( .A(n2424), .B(n4655), .ZN(n4396) );
  MUX2_X1 U3129 ( .A(n2425), .B(n4396), .S(n2042), .Z(n3353) );
  AND2_X1 U3130 ( .A1(n3406), .A2(n3353), .ZN(n2429) );
  OR2_X1 U3131 ( .A1(n3888), .A2(n2429), .ZN(n2426) );
  NAND2_X1 U3132 ( .A1(n3962), .A2(n3321), .ZN(n3350) );
  NAND2_X1 U3133 ( .A1(n3961), .A2(n3363), .ZN(n2427) );
  AND2_X1 U3134 ( .A1(n3350), .A2(n2427), .ZN(n2428) );
  OR2_X1 U3135 ( .A1(n2429), .A2(n2428), .ZN(n3335) );
  NAND2_X1 U3136 ( .A1(n3783), .A2(REG0_REG_9__SCAN_IN), .ZN(n2439) );
  INV_X1 U3137 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2430) );
  OAI21_X1 U3138 ( .B1(n2432), .B2(n2431), .A(n2430), .ZN(n2433) );
  NAND2_X1 U3139 ( .A1(n2433), .A2(n2447), .ZN(n3346) );
  OR2_X1 U3140 ( .A1(n2457), .A2(n3346), .ZN(n2438) );
  INV_X1 U3141 ( .A(REG1_REG_9__SCAN_IN), .ZN(n2434) );
  OR2_X1 U3142 ( .A1(n2527), .A2(n2434), .ZN(n2437) );
  INV_X1 U3143 ( .A(REG2_REG_9__SCAN_IN), .ZN(n2435) );
  OR2_X1 U3144 ( .A1(n2343), .A2(n2435), .ZN(n2436) );
  NAND4_X1 U3145 ( .A1(n2439), .A2(n2438), .A3(n2437), .A4(n2436), .ZN(n3960)
         );
  NOR2_X1 U3146 ( .A1(n2282), .A2(n2964), .ZN(n2440) );
  MUX2_X1 U3147 ( .A(n2964), .B(n2440), .S(IR_REG_9__SCAN_IN), .Z(n2442) );
  INV_X1 U31480 ( .A(n2465), .ZN(n2441) );
  MUX2_X1 U31490 ( .A(DATAI_9_), .B(n4009), .S(n3786), .Z(n3403) );
  AND2_X1 U3150 ( .A1(n3335), .A2(n2058), .ZN(n2443) );
  INV_X1 U3151 ( .A(n3960), .ZN(n3302) );
  NAND2_X1 U3152 ( .A1(n3302), .A2(n2801), .ZN(n2444) );
  NAND2_X1 U3153 ( .A1(n3783), .A2(REG0_REG_10__SCAN_IN), .ZN(n2453) );
  INV_X1 U3154 ( .A(REG1_REG_10__SCAN_IN), .ZN(n2446) );
  OR2_X1 U3155 ( .A1(n2527), .A2(n2446), .ZN(n2452) );
  INV_X1 U3156 ( .A(REG3_REG_10__SCAN_IN), .ZN(n4666) );
  NAND2_X1 U3157 ( .A1(n2447), .A2(n4666), .ZN(n2448) );
  NAND2_X1 U3158 ( .A1(n2459), .A2(n2448), .ZN(n3644) );
  OR2_X1 U3159 ( .A1(n2457), .A2(n3644), .ZN(n2451) );
  INV_X1 U3160 ( .A(REG2_REG_10__SCAN_IN), .ZN(n2449) );
  OR2_X1 U3161 ( .A1(n2343), .A2(n2449), .ZN(n2450) );
  NAND2_X1 U3162 ( .A1(n2465), .A2(IR_REG_31__SCAN_IN), .ZN(n2454) );
  XNOR2_X1 U3163 ( .A(n2454), .B(IR_REG_10__SCAN_IN), .ZN(n4014) );
  MUX2_X1 U3164 ( .A(DATAI_10_), .B(n4014), .S(n3786), .Z(n3643) );
  NOR2_X1 U3165 ( .A1(n3959), .A2(n3643), .ZN(n2455) );
  NAND2_X1 U3166 ( .A1(n3783), .A2(REG0_REG_11__SCAN_IN), .ZN(n2464) );
  INV_X1 U3167 ( .A(REG1_REG_11__SCAN_IN), .ZN(n2456) );
  OR2_X1 U3168 ( .A1(n2527), .A2(n2456), .ZN(n2463) );
  NAND2_X1 U3169 ( .A1(n2459), .A2(n2458), .ZN(n2460) );
  NAND2_X1 U3170 ( .A1(n2472), .A2(n2460), .ZN(n3399) );
  OR2_X1 U3171 ( .A1(n2457), .A2(n3399), .ZN(n2462) );
  INV_X1 U3172 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3387) );
  OR2_X1 U3173 ( .A1(n2343), .A2(n3387), .ZN(n2461) );
  OR2_X1 U3174 ( .A1(n2465), .A2(IR_REG_10__SCAN_IN), .ZN(n2466) );
  NAND2_X1 U3175 ( .A1(n2466), .A2(IR_REG_31__SCAN_IN), .ZN(n2468) );
  INV_X1 U3176 ( .A(IR_REG_11__SCAN_IN), .ZN(n2467) );
  OR2_X1 U3177 ( .A1(n2468), .A2(n2467), .ZN(n2469) );
  NAND2_X1 U3178 ( .A1(n2468), .A2(n2467), .ZN(n2479) );
  MUX2_X1 U3179 ( .A(DATAI_11_), .B(n4533), .S(n3786), .Z(n3455) );
  NAND2_X1 U3180 ( .A1(n3546), .A2(n3455), .ZN(n3799) );
  INV_X1 U3181 ( .A(n3455), .ZN(n2815) );
  NAND2_X1 U3182 ( .A1(n3958), .A2(n2815), .ZN(n3839) );
  NAND2_X1 U3183 ( .A1(n3546), .A2(n2815), .ZN(n2471) );
  NAND2_X1 U3184 ( .A1(n3783), .A2(REG0_REG_12__SCAN_IN), .ZN(n2478) );
  INV_X1 U3185 ( .A(REG2_REG_12__SCAN_IN), .ZN(n3495) );
  OR2_X1 U3186 ( .A1(n2343), .A2(n3495), .ZN(n2477) );
  NAND2_X1 U3187 ( .A1(n2472), .A2(n4681), .ZN(n2473) );
  NAND2_X1 U3188 ( .A1(n2474), .A2(n2473), .ZN(n3494) );
  OR2_X1 U3189 ( .A1(n2457), .A2(n3494), .ZN(n2476) );
  INV_X1 U3190 ( .A(REG1_REG_12__SCAN_IN), .ZN(n3554) );
  OR2_X1 U3191 ( .A1(n2527), .A2(n3554), .ZN(n2475) );
  INV_X1 U3192 ( .A(DATAI_12_), .ZN(n2481) );
  NAND2_X1 U3193 ( .A1(n2479), .A2(IR_REG_31__SCAN_IN), .ZN(n2480) );
  XNOR2_X1 U3194 ( .A(n2480), .B(IR_REG_12__SCAN_IN), .ZN(n4018) );
  MUX2_X1 U3195 ( .A(n2481), .B(n4532), .S(n2042), .Z(n3541) );
  NAND2_X1 U3196 ( .A1(n2483), .A2(n2482), .ZN(n3477) );
  NAND2_X1 U3197 ( .A1(n3783), .A2(REG0_REG_14__SCAN_IN), .ZN(n2491) );
  INV_X1 U3198 ( .A(REG1_REG_14__SCAN_IN), .ZN(n3566) );
  OR2_X1 U3199 ( .A1(n2527), .A2(n3566), .ZN(n2490) );
  INV_X1 U3200 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4573) );
  NAND2_X1 U3201 ( .A1(n2484), .A2(n4573), .ZN(n2485) );
  NAND2_X1 U3202 ( .A1(n2486), .A2(n2485), .ZN(n3529) );
  OR2_X1 U3203 ( .A1(n2457), .A2(n3529), .ZN(n2489) );
  INV_X1 U3204 ( .A(REG2_REG_14__SCAN_IN), .ZN(n2487) );
  OR2_X1 U3205 ( .A1(n2343), .A2(n2487), .ZN(n2488) );
  OR2_X1 U3206 ( .A1(n2492), .A2(n2964), .ZN(n2493) );
  XNOR2_X1 U3207 ( .A(n2493), .B(IR_REG_14__SCAN_IN), .ZN(n4022) );
  MUX2_X1 U3208 ( .A(DATAI_14_), .B(n4022), .S(n3786), .Z(n3526) );
  NAND2_X1 U3209 ( .A1(n3584), .A2(n3526), .ZN(n3795) );
  NAND2_X1 U32100 ( .A1(n3955), .A2(n3557), .ZN(n3792) );
  NAND2_X1 U32110 ( .A1(n3795), .A2(n3792), .ZN(n3434) );
  NAND2_X1 U32120 ( .A1(n3509), .A2(n2073), .ZN(n2495) );
  OAI21_X1 U32130 ( .B1(n3767), .B2(n3954), .A(n2495), .ZN(n3572) );
  NAND2_X1 U32140 ( .A1(n4323), .A2(n3685), .ZN(n3909) );
  NAND2_X1 U32150 ( .A1(n3953), .A2(n4329), .ZN(n3911) );
  NAND2_X1 U32160 ( .A1(n3783), .A2(REG0_REG_17__SCAN_IN), .ZN(n2503) );
  INV_X1 U32170 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4326) );
  OR2_X1 U32180 ( .A1(n2527), .A2(n4326), .ZN(n2502) );
  INV_X1 U32190 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2496) );
  INV_X1 U32200 ( .A(n2512), .ZN(n2514) );
  NAND2_X1 U32210 ( .A1(n2497), .A2(n2496), .ZN(n2498) );
  NAND2_X1 U32220 ( .A1(n2514), .A2(n2498), .ZN(n3698) );
  OR2_X1 U32230 ( .A1(n3698), .A2(n2457), .ZN(n2501) );
  INV_X1 U32240 ( .A(REG2_REG_17__SCAN_IN), .ZN(n2499) );
  OR2_X1 U32250 ( .A1(n2343), .A2(n2499), .ZN(n2500) );
  INV_X1 U32260 ( .A(DATAI_17_), .ZN(n2505) );
  OR2_X1 U32270 ( .A1(n2520), .A2(n2964), .ZN(n2504) );
  XNOR2_X1 U32280 ( .A(n2504), .B(IR_REG_17__SCAN_IN), .ZN(n4029) );
  MUX2_X1 U32290 ( .A(n2505), .B(n4528), .S(n3786), .Z(n3603) );
  INV_X1 U32300 ( .A(REG0_REG_18__SCAN_IN), .ZN(n2508) );
  OR2_X1 U32310 ( .A1(n2509), .A2(n2508), .ZN(n2511) );
  INV_X1 U32320 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4031) );
  OR2_X1 U32330 ( .A1(n2527), .A2(n4031), .ZN(n2510) );
  AND2_X1 U32340 ( .A1(n2511), .A2(n2510), .ZN(n2518) );
  INV_X1 U32350 ( .A(n2524), .ZN(n2525) );
  INV_X1 U32360 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2513) );
  NAND2_X1 U32370 ( .A1(n2514), .A2(n2513), .ZN(n2515) );
  NAND2_X1 U32380 ( .A1(n2525), .A2(n2515), .ZN(n4234) );
  OR2_X1 U32390 ( .A1(n4234), .A2(n2457), .ZN(n2517) );
  NAND2_X1 U32400 ( .A1(n2361), .A2(REG2_REG_18__SCAN_IN), .ZN(n2516) );
  NAND2_X1 U32410 ( .A1(n2530), .A2(IR_REG_31__SCAN_IN), .ZN(n2521) );
  XNOR2_X1 U32420 ( .A(n2521), .B(IR_REG_18__SCAN_IN), .ZN(n4006) );
  MUX2_X1 U32430 ( .A(DATAI_18_), .B(n4006), .S(n3786), .Z(n4221) );
  NAND2_X1 U32440 ( .A1(n4206), .A2(n4221), .ZN(n4201) );
  NAND2_X1 U32450 ( .A1(n4320), .A2(n2522), .ZN(n4202) );
  NAND2_X1 U32460 ( .A1(n4201), .A2(n4202), .ZN(n4228) );
  INV_X1 U32470 ( .A(n2533), .ZN(n2534) );
  INV_X1 U32480 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4665) );
  NAND2_X1 U32490 ( .A1(n2525), .A2(n4665), .ZN(n2526) );
  NAND2_X1 U32500 ( .A1(n2534), .A2(n2526), .ZN(n4214) );
  AOI22_X1 U32510 ( .A1(n2361), .A2(REG2_REG_19__SCAN_IN), .B1(n3783), .B2(
        REG0_REG_19__SCAN_IN), .ZN(n2529) );
  INV_X1 U32520 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4310) );
  OR2_X1 U32530 ( .A1(n2527), .A2(n4310), .ZN(n2528) );
  MUX2_X1 U32540 ( .A(DATAI_19_), .B(n4395), .S(n2042), .Z(n3652) );
  OR2_X1 U32550 ( .A1(n4222), .A2(n3652), .ZN(n3867) );
  INV_X1 U32560 ( .A(n3867), .ZN(n4177) );
  INV_X1 U32570 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4306) );
  INV_X1 U32580 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4571) );
  NAND2_X1 U32590 ( .A1(n2534), .A2(n4571), .ZN(n2535) );
  NAND2_X1 U32600 ( .A1(n2547), .A2(n2535), .ZN(n4187) );
  OR2_X1 U32610 ( .A1(n4187), .A2(n2457), .ZN(n2537) );
  AOI22_X1 U32620 ( .A1(n2361), .A2(REG2_REG_20__SCAN_IN), .B1(n3783), .B2(
        REG0_REG_20__SCAN_IN), .ZN(n2536) );
  INV_X1 U32630 ( .A(DATAI_20_), .ZN(n2538) );
  NAND2_X1 U32640 ( .A1(n4289), .A2(n4184), .ZN(n3873) );
  NAND2_X1 U32650 ( .A1(n4222), .A2(n3652), .ZN(n4178) );
  OAI211_X1 U32660 ( .C1(n4176), .C2(n4177), .A(n3873), .B(n4178), .ZN(n2539)
         );
  INV_X1 U32670 ( .A(n4289), .ZN(n3664) );
  INV_X1 U32680 ( .A(n4184), .ZN(n4297) );
  NAND2_X1 U32690 ( .A1(n3664), .A2(n4297), .ZN(n3874) );
  NAND2_X1 U32700 ( .A1(n2539), .A2(n3874), .ZN(n4157) );
  XNOR2_X1 U32710 ( .A(n2547), .B(REG3_REG_21__SCAN_IN), .ZN(n4163) );
  NAND2_X1 U32720 ( .A1(n2360), .A2(n4163), .ZN(n2544) );
  INV_X1 U32730 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4295) );
  NAND2_X1 U32740 ( .A1(n3783), .A2(REG0_REG_21__SCAN_IN), .ZN(n2541) );
  NAND2_X1 U32750 ( .A1(n2361), .A2(REG2_REG_21__SCAN_IN), .ZN(n2540) );
  OAI211_X1 U32760 ( .C1(n2527), .C2(n4295), .A(n2541), .B(n2540), .ZN(n2542)
         );
  INV_X1 U32770 ( .A(n2542), .ZN(n2543) );
  NAND2_X1 U32780 ( .A1(n2089), .A2(DATAI_21_), .ZN(n4167) );
  INV_X1 U32790 ( .A(n4167), .ZN(n4287) );
  NAND2_X1 U32800 ( .A1(n4300), .A2(n4287), .ZN(n2545) );
  INV_X1 U32810 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3665) );
  INV_X1 U32820 ( .A(REG3_REG_22__SCAN_IN), .ZN(n3623) );
  OAI21_X1 U32830 ( .B1(n2547), .B2(n3665), .A(n3623), .ZN(n2548) );
  NAND2_X1 U32840 ( .A1(REG3_REG_21__SCAN_IN), .A2(REG3_REG_22__SCAN_IN), .ZN(
        n2546) );
  AND2_X1 U32850 ( .A1(n2548), .A2(n2558), .ZN(n4147) );
  NAND2_X1 U32860 ( .A1(n2360), .A2(n4147), .ZN(n2553) );
  INV_X1 U32870 ( .A(REG1_REG_22__SCAN_IN), .ZN(n4285) );
  NAND2_X1 U32880 ( .A1(n3783), .A2(REG0_REG_22__SCAN_IN), .ZN(n2550) );
  NAND2_X1 U32890 ( .A1(n2361), .A2(REG2_REG_22__SCAN_IN), .ZN(n2549) );
  OAI211_X1 U32900 ( .C1(n2527), .C2(n4285), .A(n2550), .B(n2549), .ZN(n2551)
         );
  INV_X1 U32910 ( .A(n2551), .ZN(n2552) );
  INV_X1 U32920 ( .A(DATAI_22_), .ZN(n2554) );
  NOR2_X1 U32930 ( .A1(n3786), .A2(n2554), .ZN(n2555) );
  NAND2_X1 U32940 ( .A1(n4292), .A2(n2555), .ZN(n4125) );
  INV_X1 U32950 ( .A(n4292), .ZN(n4161) );
  NAND2_X1 U32960 ( .A1(n4161), .A2(n4144), .ZN(n2652) );
  NAND2_X1 U32970 ( .A1(n4125), .A2(n2652), .ZN(n4149) );
  INV_X1 U32980 ( .A(REG3_REG_23__SCAN_IN), .ZN(n4682) );
  NAND2_X1 U32990 ( .A1(n2558), .A2(n4682), .ZN(n2559) );
  NAND2_X1 U33000 ( .A1(n2566), .A2(n2559), .ZN(n4133) );
  OR2_X1 U33010 ( .A1(n4133), .A2(n2457), .ZN(n2564) );
  INV_X1 U33020 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4279) );
  NAND2_X1 U33030 ( .A1(n2361), .A2(REG2_REG_23__SCAN_IN), .ZN(n2561) );
  NAND2_X1 U33040 ( .A1(n3783), .A2(REG0_REG_23__SCAN_IN), .ZN(n2560) );
  OAI211_X1 U33050 ( .C1(n4279), .C2(n2527), .A(n2561), .B(n2560), .ZN(n2562)
         );
  INV_X1 U33060 ( .A(n2562), .ZN(n2563) );
  NAND2_X1 U33070 ( .A1(n2089), .A2(DATAI_23_), .ZN(n4132) );
  NAND2_X1 U33080 ( .A1(n4140), .A2(n4132), .ZN(n2565) );
  INV_X1 U33090 ( .A(REG3_REG_24__SCAN_IN), .ZN(n3706) );
  NAND2_X1 U33100 ( .A1(n2566), .A2(n3706), .ZN(n2567) );
  NAND2_X1 U33110 ( .A1(n2576), .A2(n2567), .ZN(n3705) );
  INV_X1 U33120 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4275) );
  NAND2_X1 U33130 ( .A1(n2361), .A2(REG2_REG_24__SCAN_IN), .ZN(n2569) );
  NAND2_X1 U33140 ( .A1(n3783), .A2(REG0_REG_24__SCAN_IN), .ZN(n2568) );
  OAI211_X1 U33150 ( .C1(n4275), .C2(n2527), .A(n2569), .B(n2568), .ZN(n2570)
         );
  INV_X1 U33160 ( .A(n2570), .ZN(n2571) );
  INV_X1 U33170 ( .A(DATAI_24_), .ZN(n2573) );
  NOR2_X1 U33180 ( .A1(n2042), .A2(n2573), .ZN(n4268) );
  NAND2_X1 U33190 ( .A1(n4260), .A2(n4268), .ZN(n2574) );
  INV_X1 U33200 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4603) );
  NAND2_X1 U33210 ( .A1(n2576), .A2(n4603), .ZN(n2577) );
  NAND2_X1 U33220 ( .A1(n2585), .A2(n2577), .ZN(n3675) );
  INV_X1 U33230 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4266) );
  NAND2_X1 U33240 ( .A1(n2361), .A2(REG2_REG_25__SCAN_IN), .ZN(n2579) );
  NAND2_X1 U33250 ( .A1(n3783), .A2(REG0_REG_25__SCAN_IN), .ZN(n2578) );
  OAI211_X1 U33260 ( .C1(n4266), .C2(n2527), .A(n2579), .B(n2578), .ZN(n2580)
         );
  INV_X1 U33270 ( .A(n2580), .ZN(n2581) );
  NAND2_X1 U33280 ( .A1(n2089), .A2(DATAI_25_), .ZN(n4258) );
  NAND2_X1 U33290 ( .A1(n4272), .A2(n4258), .ZN(n2584) );
  NOR2_X1 U33300 ( .A1(n4272), .A2(n4258), .ZN(n2583) );
  INV_X1 U33310 ( .A(REG3_REG_26__SCAN_IN), .ZN(n3750) );
  NAND2_X1 U33320 ( .A1(n2585), .A2(n3750), .ZN(n2586) );
  NAND2_X1 U33330 ( .A1(n2360), .A2(n4084), .ZN(n2591) );
  INV_X1 U33340 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4256) );
  NAND2_X1 U33350 ( .A1(n2361), .A2(REG2_REG_26__SCAN_IN), .ZN(n2588) );
  NAND2_X1 U33360 ( .A1(n3783), .A2(REG0_REG_26__SCAN_IN), .ZN(n2587) );
  OAI211_X1 U33370 ( .C1(n4256), .C2(n2527), .A(n2588), .B(n2587), .ZN(n2589)
         );
  INV_X1 U33380 ( .A(n2589), .ZN(n2590) );
  INV_X1 U33390 ( .A(DATAI_26_), .ZN(n2592) );
  NOR2_X1 U33400 ( .A1(n2042), .A2(n2592), .ZN(n2887) );
  NAND2_X1 U33410 ( .A1(n4097), .A2(n2887), .ZN(n2594) );
  NOR2_X1 U33420 ( .A1(n4097), .A2(n2887), .ZN(n2593) );
  INV_X1 U33430 ( .A(n2596), .ZN(n2595) );
  NAND2_X1 U33440 ( .A1(n2595), .A2(REG3_REG_27__SCAN_IN), .ZN(n2605) );
  INV_X1 U33450 ( .A(REG3_REG_27__SCAN_IN), .ZN(n4586) );
  NAND2_X1 U33460 ( .A1(n2596), .A2(n4586), .ZN(n2597) );
  NAND2_X1 U33470 ( .A1(n2605), .A2(n2597), .ZN(n3634) );
  INV_X1 U33480 ( .A(REG1_REG_27__SCAN_IN), .ZN(n2600) );
  NAND2_X1 U33490 ( .A1(n2361), .A2(REG2_REG_27__SCAN_IN), .ZN(n2599) );
  NAND2_X1 U33500 ( .A1(n3783), .A2(REG0_REG_27__SCAN_IN), .ZN(n2598) );
  OAI211_X1 U33510 ( .C1(n2600), .C2(n2527), .A(n2599), .B(n2598), .ZN(n2601)
         );
  INV_X1 U33520 ( .A(n2601), .ZN(n2602) );
  NAND2_X1 U3353 ( .A1(n2089), .A2(DATAI_27_), .ZN(n4247) );
  NAND2_X1 U33540 ( .A1(n3754), .A2(n4247), .ZN(n2604) );
  INV_X1 U3355 ( .A(REG3_REG_28__SCAN_IN), .ZN(n2927) );
  NAND2_X1 U3356 ( .A1(n2605), .A2(n2927), .ZN(n2606) );
  NAND2_X1 U3357 ( .A1(n4053), .A2(n2606), .ZN(n3609) );
  INV_X1 U3358 ( .A(REG1_REG_28__SCAN_IN), .ZN(n2609) );
  NAND2_X1 U3359 ( .A1(n2361), .A2(REG2_REG_28__SCAN_IN), .ZN(n2608) );
  NAND2_X1 U3360 ( .A1(n3783), .A2(REG0_REG_28__SCAN_IN), .ZN(n2607) );
  OAI211_X1 U3361 ( .C1(n2609), .C2(n2527), .A(n2608), .B(n2607), .ZN(n2610)
         );
  INV_X1 U3362 ( .A(n2610), .ZN(n2611) );
  INV_X1 U3363 ( .A(DATAI_28_), .ZN(n2613) );
  NOR2_X1 U3364 ( .A1(n2042), .A2(n2613), .ZN(n2924) );
  NAND2_X1 U3365 ( .A1(n4049), .A2(n2924), .ZN(n3782) );
  INV_X1 U3366 ( .A(n2924), .ZN(n3613) );
  NAND2_X1 U3367 ( .A1(n4250), .A2(n3613), .ZN(n3780) );
  OAI22_X1 U3368 ( .A1(n2718), .A2(n3905), .B1(n4049), .B2(n3613), .ZN(n2620)
         );
  OR2_X1 U3369 ( .A1(n4053), .A2(n2457), .ZN(n2618) );
  INV_X1 U3370 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2713) );
  NAND2_X1 U3371 ( .A1(n2361), .A2(REG2_REG_29__SCAN_IN), .ZN(n2615) );
  NAND2_X1 U3372 ( .A1(n2041), .A2(REG0_REG_29__SCAN_IN), .ZN(n2614) );
  OAI211_X1 U3373 ( .C1(n2713), .C2(n2527), .A(n2615), .B(n2614), .ZN(n2616)
         );
  INV_X1 U3374 ( .A(n2616), .ZN(n2617) );
  NAND2_X1 U3375 ( .A1(n2618), .A2(n2617), .ZN(n3951) );
  INV_X1 U3376 ( .A(DATAI_29_), .ZN(n2619) );
  NOR2_X1 U3377 ( .A1(n3786), .A2(n2619), .ZN(n4051) );
  XNOR2_X1 U3378 ( .A(n3951), .B(n4051), .ZN(n3904) );
  XNOR2_X1 U3379 ( .A(n2620), .B(n3904), .ZN(n4046) );
  NOR2_X1 U3380 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2626)
         );
  INV_X1 U3381 ( .A(IR_REG_21__SCAN_IN), .ZN(n2622) );
  AND2_X1 U3382 ( .A1(n2626), .A2(n2622), .ZN(n2623) );
  NAND2_X1 U3383 ( .A1(n2681), .A2(IR_REG_31__SCAN_IN), .ZN(n2625) );
  INV_X1 U3384 ( .A(IR_REG_22__SCAN_IN), .ZN(n2624) );
  XNOR2_X1 U3385 ( .A(n2625), .B(n2624), .ZN(n2731) );
  INV_X1 U3386 ( .A(n2731), .ZN(n4393) );
  NAND2_X1 U3387 ( .A1(n2627), .A2(n2626), .ZN(n2628) );
  NAND2_X1 U3388 ( .A1(n2628), .A2(IR_REG_31__SCAN_IN), .ZN(n2629) );
  INV_X1 U3389 ( .A(IR_REG_19__SCAN_IN), .ZN(n2630) );
  NAND2_X1 U3390 ( .A1(n2631), .A2(n2630), .ZN(n2632) );
  XNOR2_X1 U3391 ( .A(n4393), .B(n2732), .ZN(n2635) );
  INV_X1 U3392 ( .A(n4395), .ZN(n4036) );
  NAND2_X1 U3393 ( .A1(n2635), .A2(n4036), .ZN(n3228) );
  AND2_X1 U3394 ( .A1(n2636), .A2(n4395), .ZN(n3943) );
  INV_X1 U3395 ( .A(n4552), .ZN(n4540) );
  INV_X1 U3396 ( .A(n4051), .ZN(n3778) );
  NAND2_X1 U3397 ( .A1(n2731), .A2(n2691), .ZN(n2911) );
  NAND2_X1 U3398 ( .A1(n3150), .A2(n3807), .ZN(n3163) );
  NAND2_X1 U3399 ( .A1(n3079), .A2(n3165), .ZN(n3812) );
  NAND2_X1 U3400 ( .A1(n3966), .A2(n3260), .ZN(n3809) );
  AND2_X1 U3401 ( .A1(n3812), .A2(n3809), .ZN(n3885) );
  INV_X1 U3402 ( .A(n3813), .ZN(n2638) );
  AND2_X1 U3403 ( .A1(n3964), .A2(n3289), .ZN(n3224) );
  NAND2_X1 U3404 ( .A1(n3716), .A2(n3230), .ZN(n3826) );
  NAND2_X1 U3405 ( .A1(n3963), .A2(n3249), .ZN(n3825) );
  INV_X1 U3406 ( .A(n3963), .ZN(n3290) );
  NAND2_X1 U3407 ( .A1(n3290), .A2(n3191), .ZN(n3818) );
  INV_X1 U3408 ( .A(n2639), .ZN(n2640) );
  NAND2_X1 U3409 ( .A1(n3406), .A2(n3363), .ZN(n3821) );
  NAND2_X1 U3410 ( .A1(n3352), .A2(n3821), .ZN(n2641) );
  NAND2_X1 U3411 ( .A1(n3961), .A2(n3353), .ZN(n3824) );
  NAND2_X1 U3412 ( .A1(n2641), .A2(n3824), .ZN(n3328) );
  AND2_X1 U3413 ( .A1(n3960), .A2(n2801), .ZN(n3836) );
  NAND2_X1 U3414 ( .A1(n3302), .A2(n3403), .ZN(n3822) );
  NAND2_X1 U3415 ( .A1(n3959), .A2(n3423), .ZN(n3838) );
  NAND2_X1 U3416 ( .A1(n3370), .A2(n3838), .ZN(n2642) );
  NAND2_X1 U3417 ( .A1(n3332), .A2(n3643), .ZN(n3833) );
  NAND2_X1 U3418 ( .A1(n2642), .A2(n3833), .ZN(n3381) );
  NAND2_X1 U3419 ( .A1(n3381), .A2(n3839), .ZN(n2643) );
  NAND2_X1 U3420 ( .A1(n3957), .A2(n3541), .ZN(n3487) );
  NAND2_X1 U3421 ( .A1(n3956), .A2(n3478), .ZN(n3469) );
  NAND2_X1 U3422 ( .A1(n3501), .A2(n3840), .ZN(n2644) );
  NOR2_X1 U3423 ( .A1(n3957), .A2(n3541), .ZN(n3488) );
  NOR2_X1 U3424 ( .A1(n3956), .A2(n3478), .ZN(n3470) );
  AOI21_X1 U3425 ( .B1(n3840), .B2(n3488), .A(n3470), .ZN(n3797) );
  INV_X1 U3426 ( .A(n3434), .ZN(n3882) );
  NAND2_X1 U3427 ( .A1(n3908), .A2(n3882), .ZN(n2645) );
  NAND2_X1 U3428 ( .A1(n4334), .A2(n3767), .ZN(n3794) );
  NAND2_X1 U3429 ( .A1(n3954), .A2(n3515), .ZN(n3793) );
  NAND2_X1 U3430 ( .A1(n3794), .A2(n3793), .ZN(n3883) );
  AND2_X1 U3431 ( .A1(n2506), .A2(n3603), .ZN(n3790) );
  NAND2_X1 U3432 ( .A1(n4289), .A2(n4297), .ZN(n2650) );
  INV_X1 U3433 ( .A(n3652), .ZN(n4211) );
  NAND2_X1 U3434 ( .A1(n4222), .A2(n4211), .ZN(n2646) );
  NAND2_X1 U3435 ( .A1(n2650), .A2(n4173), .ZN(n3791) );
  INV_X1 U3436 ( .A(n4173), .ZN(n2648) );
  NAND2_X1 U3437 ( .A1(n4332), .A2(n4317), .ZN(n4199) );
  AND2_X1 U3438 ( .A1(n4201), .A2(n4199), .ZN(n2647) );
  OAI22_X1 U3439 ( .A1(n2648), .A2(n2647), .B1(n4211), .B2(n4222), .ZN(n4172)
         );
  NOR2_X1 U3440 ( .A1(n4289), .A2(n4297), .ZN(n2649) );
  OR2_X1 U3441 ( .A1(n4172), .A2(n2649), .ZN(n2651) );
  NAND2_X1 U3442 ( .A1(n2651), .A2(n2650), .ZN(n3914) );
  OR2_X1 U3443 ( .A1(n4300), .A2(n4167), .ZN(n3895) );
  AND2_X1 U3444 ( .A1(n4125), .A2(n3895), .ZN(n3915) );
  INV_X1 U3445 ( .A(n3915), .ZN(n2654) );
  NAND2_X1 U3446 ( .A1(n4269), .A2(n4132), .ZN(n3878) );
  AND2_X1 U3447 ( .A1(n3878), .A2(n2652), .ZN(n3848) );
  AND2_X1 U3448 ( .A1(n4300), .A2(n4167), .ZN(n4122) );
  NAND2_X1 U3449 ( .A1(n4125), .A2(n4122), .ZN(n2653) );
  AND2_X1 U3450 ( .A1(n3848), .A2(n2653), .ZN(n3917) );
  NAND2_X1 U3451 ( .A1(n4140), .A2(n2708), .ZN(n3879) );
  NOR2_X1 U3452 ( .A1(n4260), .A2(n4116), .ZN(n3893) );
  OR2_X1 U3453 ( .A1(n4097), .A2(n4083), .ZN(n2655) );
  INV_X1 U3454 ( .A(n3923), .ZN(n2656) );
  NAND2_X1 U3455 ( .A1(n4112), .A2(n4258), .ZN(n3860) );
  NAND2_X1 U3456 ( .A1(n4260), .A2(n4116), .ZN(n4089) );
  NAND2_X1 U3457 ( .A1(n3860), .A2(n4089), .ZN(n4074) );
  AND2_X1 U34580 ( .A1(n4097), .A2(n4083), .ZN(n3925) );
  AOI21_X1 U34590 ( .B1(n3923), .B2(n4074), .A(n3925), .ZN(n3852) );
  XNOR2_X1 U3460 ( .A(n4079), .B(n4247), .ZN(n4066) );
  OR2_X2 U3461 ( .A1(n4067), .A2(n4066), .ZN(n4069) );
  INV_X1 U3462 ( .A(n4247), .ZN(n4061) );
  NAND2_X1 U3463 ( .A1(n3754), .A2(n4061), .ZN(n3781) );
  INV_X1 U3464 ( .A(n3782), .ZN(n2657) );
  AOI21_X1 U3465 ( .B1(n2720), .B2(n3780), .A(n2657), .ZN(n2659) );
  INV_X1 U3466 ( .A(n3904), .ZN(n2658) );
  XNOR2_X1 U34670 ( .A(n2659), .B(n2658), .ZN(n2672) );
  NAND2_X1 U3468 ( .A1(n4393), .A2(n4395), .ZN(n2661) );
  INV_X1 U34690 ( .A(n2691), .ZN(n4394) );
  NAND2_X1 U3470 ( .A1(n4394), .A2(n2956), .ZN(n2660) );
  NOR2_X1 U34710 ( .A1(n2663), .A2(n2662), .ZN(n3007) );
  NOR2_X1 U3472 ( .A1(n2664), .A2(n2964), .ZN(n2665) );
  MUX2_X1 U34730 ( .A(n2964), .B(n2665), .S(IR_REG_28__SCAN_IN), .Z(n2668) );
  INV_X1 U3474 ( .A(n2666), .ZN(n2667) );
  OR2_X1 U34750 ( .A1(n2668), .A2(n2667), .ZN(n3008) );
  NAND2_X1 U3476 ( .A1(n4393), .A2(n4394), .ZN(n2912) );
  INV_X1 U34770 ( .A(n2912), .ZN(n2973) );
  NAND2_X1 U3478 ( .A1(n3008), .A2(n2973), .ZN(n4331) );
  AOI21_X1 U34790 ( .B1(B_REG_SCAN_IN), .B2(n3007), .A(n4331), .ZN(n4041) );
  INV_X1 U3480 ( .A(REG1_REG_30__SCAN_IN), .ZN(n2671) );
  NAND2_X1 U34810 ( .A1(n2361), .A2(REG2_REG_30__SCAN_IN), .ZN(n2670) );
  NAND2_X1 U3482 ( .A1(n3783), .A2(REG0_REG_30__SCAN_IN), .ZN(n2669) );
  OAI211_X1 U34830 ( .C1(n2527), .C2(n2671), .A(n2670), .B(n2669), .ZN(n3950)
         );
  AOI22_X2 U3484 ( .A1(n2672), .A2(n4225), .B1(n4041), .B2(n3950), .ZN(n4052)
         );
  NOR2_X2 U34850 ( .A1(n3008), .A2(n2912), .ZN(n4288) );
  NAND2_X1 U3486 ( .A1(n4250), .A2(n4288), .ZN(n2673) );
  OAI211_X1 U34870 ( .C1(n3778), .C2(n4330), .A(n4052), .B(n2673), .ZN(n2674)
         );
  NAND2_X1 U3488 ( .A1(n2675), .A2(IR_REG_31__SCAN_IN), .ZN(n2676) );
  MUX2_X1 U34890 ( .A(IR_REG_31__SCAN_IN), .B(n2676), .S(IR_REG_26__SCAN_IN), 
        .Z(n2677) );
  NAND2_X1 U3490 ( .A1(n2678), .A2(IR_REG_31__SCAN_IN), .ZN(n2679) );
  MUX2_X1 U34910 ( .A(IR_REG_31__SCAN_IN), .B(n2679), .S(IR_REG_25__SCAN_IN), 
        .Z(n2680) );
  NAND2_X1 U3492 ( .A1(n2680), .A2(n2675), .ZN(n2953) );
  NAND2_X1 U34930 ( .A1(n2953), .A2(B_REG_SCAN_IN), .ZN(n2683) );
  INV_X1 U3494 ( .A(IR_REG_23__SCAN_IN), .ZN(n2687) );
  NAND2_X1 U34950 ( .A1(n2688), .A2(n2687), .ZN(n2690) );
  MUX2_X1 U3496 ( .A(n2683), .B(B_REG_SCAN_IN), .S(n2686), .Z(n2684) );
  NAND2_X1 U34970 ( .A1(n3628), .A2(n2953), .ZN(n2969) );
  NAND2_X1 U3498 ( .A1(n3096), .A2(n2969), .ZN(n2705) );
  OR2_X1 U34990 ( .A1(n2688), .A2(n2687), .ZN(n2689) );
  NAND2_X1 U3500 ( .A1(n2690), .A2(n2689), .ZN(n2972) );
  NAND2_X1 U35010 ( .A1(n4552), .A2(n2691), .ZN(n2922) );
  AND2_X1 U3502 ( .A1(n2636), .A2(n4036), .ZN(n2910) );
  OR2_X1 U35030 ( .A1(n2912), .A2(n2910), .ZN(n3093) );
  NAND2_X1 U3504 ( .A1(n2922), .A2(n3093), .ZN(n2692) );
  NOR2_X1 U35050 ( .A1(n3095), .A2(n2692), .ZN(n2704) );
  NOR4_X1 U35060 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_19__SCAN_IN), .A3(
        D_REG_20__SCAN_IN), .A4(D_REG_21__SCAN_IN), .ZN(n2696) );
  NOR4_X1 U35070 ( .A1(D_REG_16__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_15__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n2695) );
  NOR4_X1 U35080 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_31__SCAN_IN), .ZN(n2694) );
  NOR4_X1 U35090 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_23__SCAN_IN), .A3(
        D_REG_24__SCAN_IN), .A4(D_REG_25__SCAN_IN), .ZN(n2693) );
  NAND4_X1 U35100 ( .A1(n2696), .A2(n2695), .A3(n2694), .A4(n2693), .ZN(n2702)
         );
  NOR2_X1 U35110 ( .A1(D_REG_2__SCAN_IN), .A2(D_REG_3__SCAN_IN), .ZN(n2700) );
  NOR4_X1 U35120 ( .A1(D_REG_29__SCAN_IN), .A2(D_REG_30__SCAN_IN), .A3(
        D_REG_4__SCAN_IN), .A4(D_REG_5__SCAN_IN), .ZN(n2699) );
  NOR4_X1 U35130 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_11__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2698) );
  NOR4_X1 U35140 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_7__SCAN_IN), .A3(
        D_REG_8__SCAN_IN), .A4(D_REG_9__SCAN_IN), .ZN(n2697) );
  NAND4_X1 U35150 ( .A1(n2700), .A2(n2699), .A3(n2698), .A4(n2697), .ZN(n2701)
         );
  NOR2_X1 U35160 ( .A1(n2702), .A2(n2701), .ZN(n2703) );
  NAND2_X1 U35170 ( .A1(n3629), .A2(n3628), .ZN(n2706) );
  NAND2_X1 U35180 ( .A1(n3167), .A2(n3260), .ZN(n3217) );
  NAND2_X1 U35190 ( .A1(n3250), .A2(n3249), .ZN(n3281) );
  OAI21_X1 U35200 ( .B1(n2724), .B2(n3778), .A(n2051), .ZN(n4054) );
  INV_X1 U35210 ( .A(n2911), .ZN(n3103) );
  NAND2_X1 U35220 ( .A1(n4560), .A2(REG0_REG_29__SCAN_IN), .ZN(n2709) );
  OAI21_X1 U35230 ( .B1(n2717), .B2(n4560), .A(n2711), .ZN(U3515) );
  NAND2_X1 U35240 ( .A1(n4567), .A2(REG1_REG_29__SCAN_IN), .ZN(n2714) );
  OAI21_X1 U35250 ( .B1(n2717), .B2(n4567), .A(n2716), .ZN(U3547) );
  INV_X1 U35260 ( .A(n4554), .ZN(n4315) );
  OAI22_X1 U35270 ( .A1(n3754), .A2(n4333), .B1(n4330), .B2(n3613), .ZN(n2719)
         );
  AOI21_X1 U35280 ( .B1(n4319), .B2(n3951), .A(n2719), .ZN(n2722) );
  XNOR2_X1 U35290 ( .A(n2720), .B(n3905), .ZN(n2721) );
  NAND2_X1 U35300 ( .A1(n2721), .A2(n4225), .ZN(n3614) );
  MUX2_X1 U35310 ( .A(REG1_REG_28__SCAN_IN), .B(n2727), .S(n4569), .Z(n2723)
         );
  INV_X1 U35320 ( .A(n2723), .ZN(n2726) );
  INV_X1 U35330 ( .A(n2724), .ZN(n2725) );
  NAND2_X1 U35340 ( .A1(n2726), .A2(n2266), .ZN(U3546) );
  INV_X1 U35350 ( .A(n2728), .ZN(n2729) );
  NAND2_X1 U35360 ( .A1(n2729), .A2(n2267), .ZN(U3514) );
  NAND2_X2 U35370 ( .A1(n2942), .A2(n3101), .ZN(n2791) );
  NAND2_X4 U35380 ( .A1(n2942), .A2(n2732), .ZN(n2901) );
  OAI22_X1 U35390 ( .A1(n2730), .A2(n2765), .B1(n2791), .B2(n2734), .ZN(n2746)
         );
  XNOR2_X1 U35400 ( .A(n2745), .B(n2746), .ZN(n3086) );
  INV_X1 U35410 ( .A(n2791), .ZN(n2783) );
  NAND2_X1 U35420 ( .A1(n2737), .A2(n2783), .ZN(n2736) );
  NAND2_X1 U35430 ( .A1(n2759), .A2(n3118), .ZN(n2742) );
  INV_X1 U35440 ( .A(n2942), .ZN(n2739) );
  AOI22_X1 U35450 ( .A1(n2783), .A2(n3118), .B1(n2739), .B2(IR_REG_0__SCAN_IN), 
        .ZN(n2740) );
  NAND2_X1 U35460 ( .A1(n2741), .A2(n2740), .ZN(n3005) );
  NAND2_X1 U35470 ( .A1(n3006), .A2(n3005), .ZN(n2744) );
  NAND2_X1 U35480 ( .A1(n2742), .A2(n2896), .ZN(n2743) );
  NAND2_X1 U35490 ( .A1(n2744), .A2(n2743), .ZN(n3085) );
  NAND2_X1 U35500 ( .A1(n3086), .A2(n3085), .ZN(n2749) );
  INV_X1 U35510 ( .A(n2745), .ZN(n2747) );
  NAND2_X1 U35520 ( .A1(n2747), .A2(n2746), .ZN(n2748) );
  NAND2_X1 U35530 ( .A1(n2749), .A2(n2748), .ZN(n3075) );
  INV_X1 U35540 ( .A(n3075), .ZN(n2757) );
  OAI22_X1 U35550 ( .A1(n2750), .A2(n2791), .B1(n2901), .B2(n3156), .ZN(n2751)
         );
  XNOR2_X1 U35560 ( .A(n2751), .B(n2896), .ZN(n2754) );
  OAI21_X1 U35570 ( .B1(n2750), .B2(n2765), .A(n2269), .ZN(n2752) );
  INV_X1 U35580 ( .A(n2752), .ZN(n2753) );
  NAND2_X1 U35590 ( .A1(n2754), .A2(n2753), .ZN(n2758) );
  NAND2_X1 U35600 ( .A1(n2755), .A2(n2758), .ZN(n3078) );
  INV_X1 U35610 ( .A(n3078), .ZN(n2756) );
  NAND2_X1 U35620 ( .A1(n3076), .A2(n2758), .ZN(n3127) );
  NAND2_X1 U35630 ( .A1(n2759), .A2(n3165), .ZN(n2760) );
  NOR2_X1 U35640 ( .A1(n2791), .A2(n3260), .ZN(n2763) );
  AOI21_X1 U35650 ( .B1(n2738), .B2(n3966), .A(n2763), .ZN(n2767) );
  XNOR2_X1 U35660 ( .A(n2766), .B(n2767), .ZN(n3128) );
  NAND2_X1 U35670 ( .A1(n3127), .A2(n3128), .ZN(n3126) );
  OAI22_X1 U35680 ( .A1(n3122), .A2(n2791), .B1(n2901), .B2(n3218), .ZN(n2764)
         );
  XNOR2_X1 U35690 ( .A(n2764), .B(n2896), .ZN(n2770) );
  OAI22_X1 U35700 ( .A1(n3122), .A2(n2765), .B1(n2919), .B2(n3218), .ZN(n2771)
         );
  XNOR2_X1 U35710 ( .A(n2770), .B(n2771), .ZN(n3712) );
  INV_X1 U35720 ( .A(n2766), .ZN(n2768) );
  NAND2_X1 U35730 ( .A1(n2768), .A2(n2767), .ZN(n3711) );
  AND2_X1 U35740 ( .A1(n3712), .A2(n3711), .ZN(n2769) );
  NAND2_X1 U35750 ( .A1(n3126), .A2(n2769), .ZN(n3713) );
  INV_X1 U35760 ( .A(n2770), .ZN(n2772) );
  NAND2_X1 U35770 ( .A1(n2772), .A2(n2771), .ZN(n2773) );
  NAND2_X1 U35780 ( .A1(n3713), .A2(n2773), .ZN(n3176) );
  OAI22_X1 U35790 ( .A1(n3716), .A2(n2919), .B1(n2901), .B2(n3289), .ZN(n2774)
         );
  XNOR2_X1 U35800 ( .A(n2774), .B(n2896), .ZN(n2775) );
  OAI22_X1 U35810 ( .A1(n3716), .A2(n2765), .B1(n2919), .B2(n3289), .ZN(n2776)
         );
  NAND2_X1 U3582 ( .A1(n3176), .A2(n3177), .ZN(n2779) );
  INV_X1 U3583 ( .A(n2775), .ZN(n2777) );
  NAND2_X1 U3584 ( .A1(n2777), .A2(n2776), .ZN(n2778) );
  NAND2_X1 U3585 ( .A1(n3963), .A2(n2783), .ZN(n2781) );
  NAND2_X1 U3586 ( .A1(n2759), .A2(n3191), .ZN(n2780) );
  NAND2_X1 U3587 ( .A1(n2781), .A2(n2780), .ZN(n2782) );
  XNOR2_X1 U3588 ( .A(n2782), .B(n2902), .ZN(n2786) );
  NAND2_X1 U3589 ( .A1(n2738), .A2(n3963), .ZN(n2785) );
  NAND2_X1 U3590 ( .A1(n2783), .A2(n3191), .ZN(n2784) );
  NAND2_X1 U3591 ( .A1(n2785), .A2(n2784), .ZN(n2787) );
  AND2_X1 U3592 ( .A1(n2786), .A2(n2787), .ZN(n3185) );
  INV_X1 U3593 ( .A(n2786), .ZN(n2789) );
  INV_X1 U3594 ( .A(n2787), .ZN(n2788) );
  NAND2_X1 U3595 ( .A1(n2789), .A2(n2788), .ZN(n3186) );
  OAI22_X1 U3596 ( .A1(n3354), .A2(n2919), .B1(n2901), .B2(n2792), .ZN(n2790)
         );
  XNOR2_X1 U3597 ( .A(n2790), .B(n2902), .ZN(n2795) );
  OAI22_X1 U3598 ( .A1(n3354), .A2(n2765), .B1(n2919), .B2(n2792), .ZN(n2794)
         );
  XNOR2_X1 U3599 ( .A(n2795), .B(n2794), .ZN(n3317) );
  NAND2_X1 U3600 ( .A1(n2795), .A2(n2794), .ZN(n2796) );
  OAI22_X1 U3601 ( .A1(n3406), .A2(n2765), .B1(n2919), .B2(n3353), .ZN(n3298)
         );
  OAI22_X1 U3602 ( .A1(n3406), .A2(n2919), .B1(n2901), .B2(n3353), .ZN(n2797)
         );
  XNOR2_X1 U3603 ( .A(n2797), .B(n2902), .ZN(n3299) );
  NAND2_X1 U3604 ( .A1(n3960), .A2(n2783), .ZN(n2799) );
  NAND2_X1 U3605 ( .A1(n2759), .A2(n3403), .ZN(n2798) );
  NAND2_X1 U3606 ( .A1(n2799), .A2(n2798), .ZN(n2800) );
  XNOR2_X1 U3607 ( .A(n2800), .B(n2896), .ZN(n2808) );
  NOR2_X1 U3608 ( .A1(n2919), .A2(n2801), .ZN(n2802) );
  AOI21_X1 U3609 ( .B1(n2738), .B2(n3960), .A(n2802), .ZN(n2807) );
  XNOR2_X1 U3610 ( .A(n2808), .B(n2807), .ZN(n3343) );
  NAND2_X1 U3611 ( .A1(n3959), .A2(n2783), .ZN(n2804) );
  NAND2_X1 U3612 ( .A1(n2759), .A2(n3643), .ZN(n2803) );
  NAND2_X1 U3613 ( .A1(n2804), .A2(n2803), .ZN(n2805) );
  XNOR2_X1 U3614 ( .A(n2805), .B(n2902), .ZN(n2812) );
  NOR2_X1 U3615 ( .A1(n2919), .A2(n3423), .ZN(n2806) );
  AOI21_X1 U3616 ( .B1(n2738), .B2(n3959), .A(n2806), .ZN(n2810) );
  XNOR2_X1 U3617 ( .A(n2812), .B(n2810), .ZN(n3641) );
  NAND2_X1 U3618 ( .A1(n2808), .A2(n2807), .ZN(n3639) );
  AND2_X1 U3619 ( .A1(n3641), .A2(n3639), .ZN(n2809) );
  NAND2_X1 U3620 ( .A1(n3341), .A2(n2809), .ZN(n3640) );
  INV_X1 U3621 ( .A(n2810), .ZN(n2811) );
  NAND2_X1 U3622 ( .A1(n2812), .A2(n2811), .ZN(n2813) );
  NAND2_X1 U3623 ( .A1(n3640), .A2(n2813), .ZN(n3393) );
  OAI22_X1 U3624 ( .A1(n3546), .A2(n2919), .B1(n2901), .B2(n2815), .ZN(n2814)
         );
  XNOR2_X1 U3625 ( .A(n2814), .B(n2896), .ZN(n2817) );
  NOR2_X1 U3626 ( .A1(n2919), .A2(n2815), .ZN(n2816) );
  AOI21_X1 U3627 ( .B1(n3958), .B2(n2738), .A(n2816), .ZN(n2818) );
  NAND2_X1 U3628 ( .A1(n2817), .A2(n2818), .ZN(n3394) );
  INV_X1 U3629 ( .A(n2817), .ZN(n2820) );
  INV_X1 U3630 ( .A(n2818), .ZN(n2819) );
  NAND2_X1 U3631 ( .A1(n2820), .A2(n2819), .ZN(n3395) );
  OAI22_X1 U3632 ( .A1(n3458), .A2(n2919), .B1(n2901), .B2(n3541), .ZN(n2821)
         );
  XNOR2_X1 U3633 ( .A(n2821), .B(n2902), .ZN(n3415) );
  OAI22_X1 U3634 ( .A1(n3458), .A2(n2765), .B1(n2791), .B2(n3541), .ZN(n3414)
         );
  OAI22_X1 U3635 ( .A1(n3542), .A2(n2791), .B1(n2901), .B2(n3478), .ZN(n2822)
         );
  XNOR2_X1 U3636 ( .A(n2822), .B(n2902), .ZN(n2823) );
  OAI22_X1 U3637 ( .A1(n3542), .A2(n2765), .B1(n2791), .B2(n3478), .ZN(n2824)
         );
  AND2_X1 U3638 ( .A1(n2823), .A2(n2824), .ZN(n3444) );
  INV_X1 U3639 ( .A(n2823), .ZN(n2826) );
  INV_X1 U3640 ( .A(n2824), .ZN(n2825) );
  NAND2_X1 U3641 ( .A1(n2826), .A2(n2825), .ZN(n3445) );
  OAI22_X1 U3642 ( .A1(n3584), .A2(n2791), .B1(n2901), .B2(n3557), .ZN(n2827)
         );
  XNOR2_X1 U3643 ( .A(n2827), .B(n2896), .ZN(n3522) );
  INV_X1 U3644 ( .A(n3522), .ZN(n2828) );
  OAI22_X1 U3645 ( .A1(n4334), .A2(n2919), .B1(n2901), .B2(n3515), .ZN(n2829)
         );
  XNOR2_X1 U3646 ( .A(n2829), .B(n2896), .ZN(n2831) );
  OAI22_X1 U3647 ( .A1(n4323), .A2(n2791), .B1(n2901), .B2(n4329), .ZN(n2830)
         );
  XNOR2_X1 U3648 ( .A(n2830), .B(n2902), .ZN(n2833) );
  OAI22_X1 U3649 ( .A1(n4323), .A2(n2765), .B1(n2791), .B2(n4329), .ZN(n2834)
         );
  XNOR2_X1 U3650 ( .A(n2833), .B(n2834), .ZN(n3682) );
  OAI22_X1 U3651 ( .A1(n4334), .A2(n2765), .B1(n2791), .B2(n3515), .ZN(n3764)
         );
  INV_X1 U3652 ( .A(n2833), .ZN(n2836) );
  INV_X1 U3653 ( .A(n2834), .ZN(n2835) );
  OAI22_X1 U3654 ( .A1(n4332), .A2(n2791), .B1(n2901), .B2(n3603), .ZN(n2839)
         );
  XNOR2_X1 U3655 ( .A(n2839), .B(n2896), .ZN(n3693) );
  NOR2_X1 U3656 ( .A1(n2791), .A2(n3603), .ZN(n2840) );
  AOI21_X1 U3657 ( .B1(n2506), .B2(n2738), .A(n2840), .ZN(n3692) );
  INV_X1 U3658 ( .A(n3693), .ZN(n2842) );
  INV_X1 U3659 ( .A(n3692), .ZN(n2841) );
  OAI22_X1 U3660 ( .A1(n4206), .A2(n2791), .B1(n2901), .B2(n2522), .ZN(n2843)
         );
  XNOR2_X1 U3661 ( .A(n2843), .B(n2896), .ZN(n2848) );
  INV_X1 U3662 ( .A(n2848), .ZN(n2846) );
  NOR2_X1 U3663 ( .A1(n2791), .A2(n2522), .ZN(n2844) );
  AOI21_X1 U3664 ( .B1(n4320), .B2(n2738), .A(n2844), .ZN(n2847) );
  INV_X1 U3665 ( .A(n2847), .ZN(n2845) );
  AND2_X1 U3666 ( .A1(n2848), .A2(n2847), .ZN(n3736) );
  AOI22_X1 U3667 ( .A1(n4222), .A2(n2738), .B1(n2886), .B2(n3652), .ZN(n2852)
         );
  NAND2_X1 U3668 ( .A1(n4222), .A2(n2783), .ZN(n2850) );
  NAND2_X1 U3669 ( .A1(n2759), .A2(n3652), .ZN(n2849) );
  NAND2_X1 U3670 ( .A1(n2850), .A2(n2849), .ZN(n2851) );
  XNOR2_X1 U3671 ( .A(n2851), .B(n2902), .ZN(n2854) );
  XOR2_X1 U3672 ( .A(n2852), .B(n2854), .Z(n3649) );
  INV_X1 U3673 ( .A(n2852), .ZN(n2853) );
  NAND2_X1 U3674 ( .A1(n4289), .A2(n2886), .ZN(n2857) );
  NAND2_X1 U3675 ( .A1(n2759), .A2(n4184), .ZN(n2856) );
  NAND2_X1 U3676 ( .A1(n2857), .A2(n2856), .ZN(n2858) );
  XNOR2_X1 U3677 ( .A(n2858), .B(n2902), .ZN(n2861) );
  NAND2_X1 U3678 ( .A1(n4289), .A2(n2738), .ZN(n2860) );
  NAND2_X1 U3679 ( .A1(n2886), .A2(n4184), .ZN(n2859) );
  NAND2_X1 U3680 ( .A1(n2860), .A2(n2859), .ZN(n2862) );
  NAND2_X1 U3681 ( .A1(n2861), .A2(n2862), .ZN(n3727) );
  NAND2_X1 U3682 ( .A1(n3726), .A2(n3727), .ZN(n3725) );
  INV_X1 U3683 ( .A(n2861), .ZN(n2864) );
  INV_X1 U3684 ( .A(n2862), .ZN(n2863) );
  NAND2_X1 U3685 ( .A1(n2864), .A2(n2863), .ZN(n3728) );
  NAND2_X1 U3686 ( .A1(n4300), .A2(n2886), .ZN(n2866) );
  NAND2_X1 U3687 ( .A1(n2759), .A2(n4287), .ZN(n2865) );
  NAND2_X1 U3688 ( .A1(n2866), .A2(n2865), .ZN(n2867) );
  XNOR2_X1 U3689 ( .A(n2867), .B(n2902), .ZN(n3660) );
  NAND2_X1 U3690 ( .A1(n4300), .A2(n2738), .ZN(n2869) );
  NAND2_X1 U3691 ( .A1(n2886), .A2(n4287), .ZN(n2868) );
  NAND2_X1 U3692 ( .A1(n2869), .A2(n2868), .ZN(n2870) );
  INV_X1 U3693 ( .A(n3660), .ZN(n2871) );
  INV_X1 U3694 ( .A(n2870), .ZN(n3659) );
  OAI22_X1 U3695 ( .A1(n4292), .A2(n2919), .B1(n2901), .B2(n4144), .ZN(n2872)
         );
  XNOR2_X1 U3696 ( .A(n2872), .B(n2902), .ZN(n2876) );
  OAI22_X1 U3697 ( .A1(n4292), .A2(n2765), .B1(n2791), .B2(n4144), .ZN(n2875)
         );
  XNOR2_X1 U3698 ( .A(n2876), .B(n2875), .ZN(n3622) );
  OAI22_X1 U3699 ( .A1(n4140), .A2(n2791), .B1(n2901), .B2(n4132), .ZN(n2874)
         );
  XNOR2_X1 U3700 ( .A(n2874), .B(n2902), .ZN(n2879) );
  OAI22_X1 U3701 ( .A1(n4140), .A2(n2765), .B1(n2791), .B2(n4132), .ZN(n2878)
         );
  XNOR2_X1 U3702 ( .A(n2879), .B(n2878), .ZN(n2947) );
  NOR2_X1 U3703 ( .A1(n2876), .A2(n2875), .ZN(n2944) );
  AND2_X1 U3704 ( .A1(n2879), .A2(n2878), .ZN(n2882) );
  OAI22_X1 U3705 ( .A1(n3676), .A2(n2765), .B1(n2791), .B2(n4116), .ZN(n2881)
         );
  OAI22_X1 U3706 ( .A1(n3676), .A2(n2791), .B1(n2901), .B2(n4116), .ZN(n2880)
         );
  XOR2_X1 U3707 ( .A(n2902), .B(n2880), .Z(n3703) );
  OAI22_X1 U3708 ( .A1(n4272), .A2(n2791), .B1(n2901), .B2(n4258), .ZN(n2883)
         );
  XNOR2_X1 U3709 ( .A(n2883), .B(n2902), .ZN(n2885) );
  OAI22_X1 U3710 ( .A1(n4272), .A2(n2765), .B1(n2791), .B2(n4258), .ZN(n2884)
         );
  OR2_X1 U3711 ( .A1(n2885), .A2(n2884), .ZN(n3671) );
  AND2_X1 U3712 ( .A1(n2885), .A2(n2884), .ZN(n3672) );
  NAND2_X1 U3713 ( .A1(n4097), .A2(n2886), .ZN(n2889) );
  NAND2_X1 U3714 ( .A1(n2759), .A2(n2887), .ZN(n2888) );
  NAND2_X1 U3715 ( .A1(n2889), .A2(n2888), .ZN(n2890) );
  XNOR2_X1 U3716 ( .A(n2890), .B(n2896), .ZN(n2895) );
  INV_X1 U3717 ( .A(n2895), .ZN(n2893) );
  NOR2_X1 U3718 ( .A1(n2791), .A2(n4083), .ZN(n2891) );
  AOI21_X1 U3719 ( .B1(n4097), .B2(n2738), .A(n2891), .ZN(n2894) );
  INV_X1 U3720 ( .A(n2894), .ZN(n2892) );
  NAND2_X1 U3721 ( .A1(n2893), .A2(n2892), .ZN(n3746) );
  AND2_X1 U3722 ( .A1(n2895), .A2(n2894), .ZN(n3745) );
  OAI22_X1 U3723 ( .A1(n3754), .A2(n2791), .B1(n4247), .B2(n2901), .ZN(n2897)
         );
  XNOR2_X1 U3724 ( .A(n2897), .B(n2896), .ZN(n2898) );
  OAI22_X1 U3725 ( .A1(n3754), .A2(n2765), .B1(n4247), .B2(n2791), .ZN(n2900)
         );
  XNOR2_X1 U3726 ( .A(n2898), .B(n2900), .ZN(n3632) );
  INV_X1 U3727 ( .A(n2898), .ZN(n2899) );
  AOI22_X1 U3728 ( .A1(n3633), .A2(n3632), .B1(n2900), .B2(n2899), .ZN(n2907)
         );
  OAI22_X1 U3729 ( .A1(n4049), .A2(n2765), .B1(n2791), .B2(n3613), .ZN(n2905)
         );
  OAI22_X1 U3730 ( .A1(n4049), .A2(n2919), .B1(n2901), .B2(n3613), .ZN(n2903)
         );
  XNOR2_X1 U3731 ( .A(n2903), .B(n2902), .ZN(n2904) );
  XOR2_X1 U3732 ( .A(n2905), .B(n2904), .Z(n2906) );
  XNOR2_X1 U3733 ( .A(n2907), .B(n2906), .ZN(n2915) );
  NAND3_X1 U3734 ( .A1(n3098), .A2(n2909), .A3(n3096), .ZN(n2933) );
  OR2_X1 U3735 ( .A1(n2911), .A2(n2910), .ZN(n2913) );
  NAND2_X1 U3736 ( .A1(n2913), .A2(n2912), .ZN(n2929) );
  OR2_X1 U3737 ( .A1(n3095), .A2(n2929), .ZN(n2914) );
  NAND2_X1 U3738 ( .A1(n2915), .A2(n3775), .ZN(n2940) );
  INV_X1 U3739 ( .A(n2916), .ZN(n2917) );
  NAND2_X1 U3740 ( .A1(n4525), .A2(n2917), .ZN(n2918) );
  NOR2_X1 U3741 ( .A1(n2919), .A2(n2918), .ZN(n3945) );
  NAND2_X1 U3742 ( .A1(n3945), .A2(n3008), .ZN(n2920) );
  OR2_X1 U3743 ( .A1(n3095), .A2(n4330), .ZN(n2921) );
  OR2_X1 U3744 ( .A1(n2933), .A2(n2921), .ZN(n2923) );
  NAND2_X1 U3745 ( .A1(n2923), .A2(n4511), .ZN(n3768) );
  AOI22_X1 U3746 ( .A1(n3951), .A2(n3766), .B1(n2924), .B2(n3768), .ZN(n2925)
         );
  INV_X1 U3747 ( .A(n2925), .ZN(n2938) );
  INV_X1 U3748 ( .A(n3008), .ZN(n4392) );
  NAND2_X1 U3749 ( .A1(n3945), .A2(n4392), .ZN(n2926) );
  OAI22_X1 U3750 ( .A1(n3754), .A2(n3751), .B1(STATE_REG_SCAN_IN), .B2(n2927), 
        .ZN(n2928) );
  INV_X1 U3751 ( .A(n2928), .ZN(n2936) );
  NAND2_X1 U3752 ( .A1(n2929), .A2(n4330), .ZN(n2930) );
  NAND2_X1 U3753 ( .A1(n2933), .A2(n2930), .ZN(n2931) );
  NAND2_X1 U3754 ( .A1(n2931), .A2(n3093), .ZN(n3057) );
  NAND2_X1 U3755 ( .A1(n2942), .A2(n2972), .ZN(n2932) );
  OAI21_X1 U3756 ( .B1(n3057), .B2(n2932), .A(STATE_REG_SCAN_IN), .ZN(n2934)
         );
  NAND2_X1 U3757 ( .A1(n2933), .A2(n3945), .ZN(n3056) );
  OR2_X1 U3758 ( .A1(n3609), .A2(n3773), .ZN(n2935) );
  NAND2_X1 U3759 ( .A1(n2936), .A2(n2935), .ZN(n2937) );
  NAND2_X1 U3760 ( .A1(n2940), .A2(n2939), .ZN(U3217) );
  INV_X1 U3761 ( .A(n4525), .ZN(n2941) );
  OR2_X1 U3762 ( .A1(n2942), .A2(n2941), .ZN(n3952) );
  INV_X2 U3763 ( .A(n3952), .ZN(U4043) );
  INV_X2 U3764 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3765 ( .A(n2943), .ZN(n3620) );
  OR2_X1 U3766 ( .A1(n3620), .A2(n2944), .ZN(n2946) );
  AOI211_X1 U3767 ( .C1(n2947), .C2(n2946), .A(n3759), .B(n2945), .ZN(n2951)
         );
  NOR2_X1 U3768 ( .A1(n3773), .A2(n4133), .ZN(n2950) );
  OAI22_X1 U3769 ( .A1(n4292), .A2(n3751), .B1(STATE_REG_SCAN_IN), .B2(n4682), 
        .ZN(n2949) );
  INV_X1 U3770 ( .A(n3768), .ZN(n3752) );
  OAI22_X1 U3771 ( .A1(n3676), .A2(n3753), .B1(n3752), .B2(n4132), .ZN(n2948)
         );
  OR4_X1 U3772 ( .A1(n2951), .A2(n2950), .A3(n2949), .A4(n2948), .ZN(U3213) );
  NAND2_X1 U3773 ( .A1(U3149), .A2(DATAI_25_), .ZN(n2952) );
  OAI21_X1 U3774 ( .B1(n2953), .B2(U3149), .A(n2952), .ZN(U3327) );
  NAND2_X1 U3775 ( .A1(n2954), .A2(STATE_REG_SCAN_IN), .ZN(n2955) );
  OAI21_X1 U3776 ( .B1(STATE_REG_SCAN_IN), .B2(n2592), .A(n2955), .ZN(U3326)
         );
  NAND2_X1 U3777 ( .A1(n2956), .A2(STATE_REG_SCAN_IN), .ZN(n2957) );
  OAI21_X1 U3778 ( .B1(STATE_REG_SCAN_IN), .B2(n2538), .A(n2957), .ZN(U3332)
         );
  INV_X1 U3779 ( .A(DATAI_27_), .ZN(n2959) );
  NAND2_X1 U3780 ( .A1(n3007), .A2(STATE_REG_SCAN_IN), .ZN(n2958) );
  OAI21_X1 U3781 ( .B1(STATE_REG_SCAN_IN), .B2(n2959), .A(n2958), .ZN(U3325)
         );
  NAND2_X1 U3782 ( .A1(n2960), .A2(STATE_REG_SCAN_IN), .ZN(n2961) );
  OAI21_X1 U3783 ( .B1(STATE_REG_SCAN_IN), .B2(n2619), .A(n2961), .ZN(U3323)
         );
  INV_X1 U3784 ( .A(DATAI_30_), .ZN(n4574) );
  NAND2_X1 U3785 ( .A1(n2962), .A2(STATE_REG_SCAN_IN), .ZN(n2963) );
  OAI21_X1 U3786 ( .B1(STATE_REG_SCAN_IN), .B2(n4574), .A(n2963), .ZN(U3322)
         );
  INV_X1 U3787 ( .A(DATAI_31_), .ZN(n4679) );
  OR4_X1 U3788 ( .A1(n2965), .A2(IR_REG_30__SCAN_IN), .A3(n2964), .A4(U3149), 
        .ZN(n2966) );
  OAI21_X1 U3789 ( .B1(STATE_REG_SCAN_IN), .B2(n4679), .A(n2966), .ZN(U3321)
         );
  INV_X1 U3790 ( .A(n3095), .ZN(n2967) );
  INV_X1 U3791 ( .A(D_REG_1__SCAN_IN), .ZN(n2971) );
  INV_X1 U3792 ( .A(n2969), .ZN(n2970) );
  AOI22_X1 U3793 ( .A1(n4524), .A2(n2971), .B1(n2970), .B2(n4525), .ZN(U3459)
         );
  OR2_X1 U3794 ( .A1(n2972), .A2(U3149), .ZN(n3948) );
  NAND2_X1 U3795 ( .A1(n3095), .A2(n3948), .ZN(n2976) );
  AOI21_X1 U3796 ( .B1(n2973), .B2(n2972), .A(n2042), .ZN(n2975) );
  INV_X1 U3797 ( .A(n2975), .ZN(n2974) );
  NOR2_X1 U3798 ( .A1(n4503), .A2(U4043), .ZN(U3148) );
  INV_X1 U3799 ( .A(n2991), .ZN(n2980) );
  INV_X1 U3800 ( .A(REG2_REG_0__SCAN_IN), .ZN(n2977) );
  AOI21_X1 U3801 ( .B1(n3007), .B2(n2977), .A(n3008), .ZN(n3010) );
  OAI21_X1 U3802 ( .B1(REG1_REG_0__SCAN_IN), .B2(n3007), .A(n3010), .ZN(n2978)
         );
  MUX2_X1 U3803 ( .A(n2978), .B(n3010), .S(IR_REG_0__SCAN_IN), .Z(n2979) );
  OAI22_X1 U3804 ( .A1(n2980), .A2(n2979), .B1(STATE_REG_SCAN_IN), .B2(n3062), 
        .ZN(n2982) );
  INV_X1 U3805 ( .A(n3007), .ZN(n2990) );
  INV_X1 U3806 ( .A(n4505), .ZN(n3044) );
  NOR3_X1 U3807 ( .A1(n3044), .A2(REG1_REG_0__SCAN_IN), .A3(n2101), .ZN(n2981)
         );
  AOI211_X1 U3808 ( .C1(n4503), .C2(ADDR_REG_0__SCAN_IN), .A(n2982), .B(n2981), 
        .ZN(n2983) );
  INV_X1 U3809 ( .A(n2983), .ZN(U3240) );
  INV_X1 U3810 ( .A(n3052), .ZN(n4399) );
  INV_X1 U3811 ( .A(REG2_REG_2__SCAN_IN), .ZN(n3018) );
  INV_X1 U3812 ( .A(n4402), .ZN(n3014) );
  MUX2_X1 U3813 ( .A(REG2_REG_2__SCAN_IN), .B(n3018), .S(n4402), .Z(n2987) );
  INV_X1 U3814 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2984) );
  MUX2_X1 U3815 ( .A(REG2_REG_1__SCAN_IN), .B(n2984), .S(n4403), .Z(n3970) );
  AND2_X1 U3816 ( .A1(REG2_REG_0__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2985)
         );
  NAND2_X1 U3817 ( .A1(n4403), .A2(REG2_REG_1__SCAN_IN), .ZN(n3019) );
  NAND2_X1 U3818 ( .A1(n3969), .A2(n3019), .ZN(n2986) );
  XNOR2_X1 U3819 ( .A(n2988), .B(n4400), .ZN(n3063) );
  INV_X1 U3820 ( .A(n2988), .ZN(n2989) );
  MUX2_X1 U3821 ( .A(REG2_REG_5__SCAN_IN), .B(n2381), .S(n3052), .Z(n3049) );
  NOR2_X1 U3822 ( .A1(n3050), .A2(n3049), .ZN(n3048) );
  AOI21_X1 U3823 ( .B1(n4399), .B2(REG2_REG_5__SCAN_IN), .A(n3048), .ZN(n3027)
         );
  XNOR2_X1 U3824 ( .A(n3027), .B(n4398), .ZN(n3029) );
  XNOR2_X1 U3825 ( .A(n3029), .B(REG2_REG_6__SCAN_IN), .ZN(n3004) );
  NOR2_X1 U3826 ( .A1(n3008), .A2(n2990), .ZN(n3944) );
  NAND2_X1 U3827 ( .A1(n2991), .A2(n3008), .ZN(n4510) );
  INV_X1 U3828 ( .A(n4510), .ZN(n3979) );
  NAND2_X1 U3829 ( .A1(n4503), .A2(ADDR_REG_6__SCAN_IN), .ZN(n2992) );
  NAND2_X1 U3830 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3189) );
  NAND2_X1 U3831 ( .A1(n2992), .A2(n3189), .ZN(n3002) );
  XNOR2_X1 U3832 ( .A(n4402), .B(n2993), .ZN(n3017) );
  XNOR2_X1 U3833 ( .A(n4403), .B(n2359), .ZN(n3974) );
  AND2_X1 U3834 ( .A1(REG1_REG_0__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n3973)
         );
  NAND2_X1 U3835 ( .A1(n3974), .A2(n3973), .ZN(n3972) );
  NAND2_X1 U3836 ( .A1(n4403), .A2(REG1_REG_1__SCAN_IN), .ZN(n2994) );
  NAND2_X1 U3837 ( .A1(n3972), .A2(n2994), .ZN(n3016) );
  NAND2_X1 U3838 ( .A1(n3017), .A2(n3016), .ZN(n3015) );
  NAND2_X1 U3839 ( .A1(n4402), .A2(REG1_REG_2__SCAN_IN), .ZN(n2995) );
  INV_X1 U3840 ( .A(n4401), .ZN(n2996) );
  XNOR2_X1 U3841 ( .A(n2997), .B(n2996), .ZN(n3981) );
  NAND2_X1 U3842 ( .A1(n3981), .A2(REG1_REG_3__SCAN_IN), .ZN(n3980) );
  NAND2_X1 U3843 ( .A1(n2997), .A2(n4401), .ZN(n2998) );
  NAND2_X1 U3844 ( .A1(n3980), .A2(n2998), .ZN(n2999) );
  INV_X1 U3845 ( .A(n4400), .ZN(n3070) );
  XNOR2_X1 U3846 ( .A(n2999), .B(n3070), .ZN(n3066) );
  XNOR2_X1 U3847 ( .A(n3052), .B(n3313), .ZN(n3046) );
  NOR2_X1 U3848 ( .A1(n3000), .A2(n2398), .ZN(n3033) );
  AOI211_X1 U3849 ( .C1(n2398), .C2(n3000), .A(n3044), .B(n3033), .ZN(n3001)
         );
  AOI211_X1 U3850 ( .C1(n3979), .C2(n4398), .A(n3002), .B(n3001), .ZN(n3003)
         );
  OAI21_X1 U3851 ( .B1(n3004), .B2(n4499), .A(n3003), .ZN(U3246) );
  XNOR2_X1 U3852 ( .A(n3006), .B(n3005), .ZN(n3059) );
  NOR2_X1 U3853 ( .A1(n3008), .A2(n3007), .ZN(n3012) );
  INV_X1 U3854 ( .A(n3944), .ZN(n3009) );
  NAND2_X1 U3855 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3968) );
  OAI22_X1 U3856 ( .A1(IR_REG_0__SCAN_IN), .A2(n3010), .B1(n3009), .B2(n3968), 
        .ZN(n3011) );
  AOI211_X1 U3857 ( .C1(n3059), .C2(n3012), .A(n3952), .B(n3011), .ZN(n3071)
         );
  AOI22_X1 U3858 ( .A1(n4503), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3013) );
  OAI21_X1 U3859 ( .B1(n4510), .B2(n3014), .A(n3013), .ZN(n3026) );
  OAI211_X1 U3860 ( .C1(n3017), .C2(n3016), .A(n4505), .B(n3015), .ZN(n3024)
         );
  MUX2_X1 U3861 ( .A(n3018), .B(REG2_REG_2__SCAN_IN), .S(n4402), .Z(n3020) );
  NAND3_X1 U3862 ( .A1(n3020), .A2(n3969), .A3(n3019), .ZN(n3021) );
  NAND3_X1 U3863 ( .A1(n4450), .A2(n3022), .A3(n3021), .ZN(n3023) );
  NAND2_X1 U3864 ( .A1(n3024), .A2(n3023), .ZN(n3025) );
  OR3_X1 U3865 ( .A1(n3071), .A2(n3026), .A3(n3025), .ZN(U3242) );
  INV_X1 U3866 ( .A(n3027), .ZN(n3028) );
  MUX2_X1 U3867 ( .A(n2408), .B(REG2_REG_7__SCAN_IN), .S(n4397), .Z(n3030) );
  NOR2_X1 U3868 ( .A1(n3031), .A2(n3030), .ZN(n3140) );
  AOI211_X1 U3869 ( .C1(n3031), .C2(n3030), .A(n4499), .B(n3140), .ZN(n3043)
         );
  INV_X1 U3870 ( .A(n3032), .ZN(n3034) );
  INV_X1 U3871 ( .A(n4397), .ZN(n3040) );
  AND2_X1 U3872 ( .A1(n3040), .A2(n2410), .ZN(n3136) );
  INV_X1 U3873 ( .A(n3136), .ZN(n3035) );
  NAND2_X1 U3874 ( .A1(n4397), .A2(REG1_REG_7__SCAN_IN), .ZN(n3137) );
  NAND2_X1 U3875 ( .A1(n3035), .A2(n3137), .ZN(n3037) );
  OAI21_X1 U3876 ( .B1(n3138), .B2(n3037), .A(n4505), .ZN(n3036) );
  AOI21_X1 U3877 ( .B1(n3138), .B2(n3037), .A(n3036), .ZN(n3042) );
  INV_X1 U3878 ( .A(REG3_REG_7__SCAN_IN), .ZN(n3038) );
  NOR2_X1 U3879 ( .A1(n3038), .A2(STATE_REG_SCAN_IN), .ZN(n3318) );
  AOI21_X1 U3880 ( .B1(n4503), .B2(ADDR_REG_7__SCAN_IN), .A(n3318), .ZN(n3039)
         );
  OAI21_X1 U3881 ( .B1(n4510), .B2(n3040), .A(n3039), .ZN(n3041) );
  OR3_X1 U3882 ( .A1(n3043), .A2(n3042), .A3(n3041), .ZN(U3247) );
  AOI211_X1 U3883 ( .C1(n3047), .C2(n3046), .A(n3045), .B(n3044), .ZN(n3055)
         );
  AOI211_X1 U3884 ( .C1(n3050), .C2(n3049), .A(n3048), .B(n4499), .ZN(n3054)
         );
  NOR2_X1 U3885 ( .A1(STATE_REG_SCAN_IN), .A2(n2378), .ZN(n3178) );
  AOI21_X1 U3886 ( .B1(n4503), .B2(ADDR_REG_5__SCAN_IN), .A(n3178), .ZN(n3051)
         );
  OAI21_X1 U3887 ( .B1(n4510), .B2(n3052), .A(n3051), .ZN(n3053) );
  OR3_X1 U3888 ( .A1(n3055), .A2(n3054), .A3(n3053), .ZN(U3245) );
  INV_X1 U3889 ( .A(n3056), .ZN(n3058) );
  NOR3_X1 U3890 ( .A1(n3058), .A2(n3057), .A3(n3095), .ZN(n3087) );
  OAI22_X1 U3891 ( .A1(n2730), .A2(n3753), .B1(n3759), .B2(n3059), .ZN(n3060)
         );
  AOI21_X1 U3892 ( .B1(n3118), .B2(n3768), .A(n3060), .ZN(n3061) );
  OAI21_X1 U3893 ( .B1(n3087), .B2(n3062), .A(n3061), .ZN(U3229) );
  XOR2_X1 U3894 ( .A(REG2_REG_4__SCAN_IN), .B(n3063), .Z(n3073) );
  INV_X1 U3895 ( .A(n3064), .ZN(n3065) );
  OAI211_X1 U3896 ( .C1(REG1_REG_4__SCAN_IN), .C2(n3066), .A(n4505), .B(n3065), 
        .ZN(n3069) );
  NAND2_X1 U3897 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n3715) );
  INV_X1 U3898 ( .A(n3715), .ZN(n3067) );
  AOI21_X1 U3899 ( .B1(n4503), .B2(ADDR_REG_4__SCAN_IN), .A(n3067), .ZN(n3068)
         );
  OAI211_X1 U3900 ( .C1(n4510), .C2(n3070), .A(n3069), .B(n3068), .ZN(n3072)
         );
  AOI211_X1 U3901 ( .C1(n4450), .C2(n3073), .A(n3072), .B(n3071), .ZN(n3074)
         );
  INV_X1 U3902 ( .A(n3074), .ZN(U3244) );
  INV_X1 U3903 ( .A(n3076), .ZN(n3077) );
  AOI21_X1 U3904 ( .B1(n3075), .B2(n3078), .A(n3077), .ZN(n3084) );
  OAI22_X1 U3905 ( .A1(n3079), .A2(n3753), .B1(n3751), .B2(n2730), .ZN(n3082)
         );
  INV_X1 U3906 ( .A(REG3_REG_2__SCAN_IN), .ZN(n3080) );
  NOR2_X1 U3907 ( .A1(n3087), .A2(n3080), .ZN(n3081) );
  AOI211_X1 U3908 ( .C1(n3268), .C2(n3768), .A(n3082), .B(n3081), .ZN(n3083)
         );
  OAI21_X1 U3909 ( .B1(n3084), .B2(n3759), .A(n3083), .ZN(U3234) );
  XNOR2_X1 U3910 ( .A(n3085), .B(n3086), .ZN(n3091) );
  OAI22_X1 U3911 ( .A1(n3112), .A2(n3751), .B1(n3753), .B2(n2750), .ZN(n3089)
         );
  INV_X1 U3912 ( .A(REG3_REG_1__SCAN_IN), .ZN(n3197) );
  NOR2_X1 U3913 ( .A1(n3087), .A2(n3197), .ZN(n3088) );
  AOI211_X1 U3914 ( .C1(n2366), .C2(n3768), .A(n3089), .B(n3088), .ZN(n3090)
         );
  OAI21_X1 U3915 ( .B1(n3091), .B2(n3759), .A(n3090), .ZN(U3219) );
  NAND2_X1 U3916 ( .A1(n2737), .A2(n3092), .ZN(n3803) );
  AND2_X1 U3917 ( .A1(n3801), .A2(n3803), .ZN(n4541) );
  INV_X1 U3918 ( .A(n3093), .ZN(n3094) );
  NOR2_X1 U3919 ( .A1(n3095), .A2(n3094), .ZN(n3097) );
  NAND4_X1 U3920 ( .A1(n3099), .A2(n3098), .A3(n3097), .A4(n3096), .ZN(n3100)
         );
  NAND2_X1 U3921 ( .A1(n3101), .A2(n4395), .ZN(n3227) );
  INV_X1 U3922 ( .A(n3227), .ZN(n3102) );
  NAND2_X1 U3923 ( .A1(n4514), .A2(n3102), .ZN(n3248) );
  NAND2_X1 U3924 ( .A1(n3118), .A2(n3103), .ZN(n4538) );
  AOI21_X1 U3925 ( .B1(n4302), .B2(n3228), .A(n4541), .ZN(n3104) );
  AOI21_X1 U3926 ( .B1(n4319), .B2(n2370), .A(n3104), .ZN(n4539) );
  OAI21_X1 U3927 ( .B1(n3943), .B2(n4538), .A(n4539), .ZN(n3105) );
  INV_X1 U3928 ( .A(n4511), .ZN(n4188) );
  AOI22_X1 U3929 ( .A1(n3105), .A2(n4514), .B1(REG3_REG_0__SCAN_IN), .B2(n4188), .ZN(n3107) );
  NAND2_X1 U3930 ( .A1(n4523), .A2(REG2_REG_0__SCAN_IN), .ZN(n3106) );
  OAI211_X1 U3931 ( .C1(n4541), .C2(n3248), .A(n3107), .B(n3106), .ZN(U3290)
         );
  OR2_X1 U3932 ( .A1(n3108), .A2(n2637), .ZN(n3109) );
  NAND2_X1 U3933 ( .A1(n3110), .A2(n3109), .ZN(n3198) );
  INV_X1 U3934 ( .A(n3198), .ZN(n3117) );
  AOI22_X1 U3935 ( .A1(n3967), .A2(n4319), .B1(n4318), .B2(n2366), .ZN(n3111)
         );
  OAI21_X1 U3936 ( .B1(n3112), .B2(n4333), .A(n3111), .ZN(n3116) );
  INV_X1 U3937 ( .A(n3113), .ZN(n3114) );
  AOI21_X1 U3938 ( .B1(n2637), .B2(n3801), .A(n3114), .ZN(n3115) );
  OAI22_X1 U3939 ( .A1(n3115), .A2(n4302), .B1(n3228), .B2(n3198), .ZN(n3199)
         );
  AOI211_X1 U3940 ( .C1(n4552), .C2(n3117), .A(n3116), .B(n3199), .ZN(n3135)
         );
  NAND2_X1 U3941 ( .A1(n3118), .A2(n2366), .ZN(n3119) );
  NAND2_X1 U3942 ( .A1(n3157), .A2(n3119), .ZN(n3204) );
  OAI22_X1 U3943 ( .A1(n4328), .A2(n3204), .B1(n4569), .B2(n2359), .ZN(n3120)
         );
  INV_X1 U3944 ( .A(n3120), .ZN(n3121) );
  OAI21_X1 U3945 ( .B1(n3135), .B2(n4567), .A(n3121), .ZN(U3519) );
  OAI22_X1 U3946 ( .A1(n2750), .A2(n3751), .B1(n3753), .B2(n3122), .ZN(n3125)
         );
  INV_X1 U3947 ( .A(n3773), .ZN(n3757) );
  MUX2_X1 U3948 ( .A(U3149), .B(n3757), .S(n3123), .Z(n3124) );
  AOI211_X1 U3949 ( .C1(n3165), .C2(n3768), .A(n3125), .B(n3124), .ZN(n3131)
         );
  OAI21_X1 U3950 ( .B1(n3128), .B2(n3127), .A(n3126), .ZN(n3129) );
  NAND2_X1 U3951 ( .A1(n3129), .A2(n3775), .ZN(n3130) );
  NAND2_X1 U3952 ( .A1(n3131), .A2(n3130), .ZN(U3215) );
  INV_X1 U3953 ( .A(REG0_REG_1__SCAN_IN), .ZN(n3132) );
  OAI22_X1 U3954 ( .A1(n4389), .A2(n3204), .B1(n4562), .B2(n3132), .ZN(n3133)
         );
  INV_X1 U3955 ( .A(n3133), .ZN(n3134) );
  OAI21_X1 U3956 ( .B1(n3135), .B2(n4560), .A(n3134), .ZN(U3469) );
  XNOR2_X1 U3957 ( .A(n4011), .B(n4396), .ZN(n4010) );
  XOR2_X1 U3958 ( .A(REG1_REG_8__SCAN_IN), .B(n4010), .Z(n3139) );
  NAND2_X1 U3959 ( .A1(n3139), .A2(n4505), .ZN(n3145) );
  AOI21_X1 U3960 ( .B1(REG2_REG_7__SCAN_IN), .B2(n4397), .A(n3140), .ZN(n3992)
         );
  XNOR2_X1 U3961 ( .A(REG2_REG_8__SCAN_IN), .B(n3993), .ZN(n3141) );
  NAND2_X1 U3962 ( .A1(n4450), .A2(n3141), .ZN(n3142) );
  NAND2_X1 U3963 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3301) );
  NAND2_X1 U3964 ( .A1(n3142), .A2(n3301), .ZN(n3143) );
  AOI21_X1 U3965 ( .B1(n4503), .B2(ADDR_REG_8__SCAN_IN), .A(n3143), .ZN(n3144)
         );
  OAI211_X1 U3966 ( .C1(n4510), .C2(n4396), .A(n3145), .B(n3144), .ZN(U3248)
         );
  NAND2_X1 U3967 ( .A1(n3147), .A2(n3880), .ZN(n3148) );
  NAND2_X1 U3968 ( .A1(n3146), .A2(n3148), .ZN(n3270) );
  AOI22_X1 U3969 ( .A1(n3966), .A2(n4319), .B1(n3268), .B2(n4318), .ZN(n3149)
         );
  OAI21_X1 U3970 ( .B1(n2730), .B2(n4333), .A(n3149), .ZN(n3155) );
  INV_X1 U3971 ( .A(n3228), .ZN(n3359) );
  NAND2_X1 U3972 ( .A1(n3270), .A2(n3359), .ZN(n3154) );
  OAI21_X1 U3973 ( .B1(n3880), .B2(n3151), .A(n3150), .ZN(n3152) );
  NAND2_X1 U3974 ( .A1(n3152), .A2(n4225), .ZN(n3153) );
  NAND2_X1 U3975 ( .A1(n3154), .A2(n3153), .ZN(n3267) );
  AOI211_X1 U3976 ( .C1(n4552), .C2(n3270), .A(n3155), .B(n3267), .ZN(n3160)
         );
  XNOR2_X1 U3977 ( .A(n3157), .B(n3156), .ZN(n3269) );
  AOI22_X1 U3978 ( .A1(n4351), .A2(n3269), .B1(REG0_REG_2__SCAN_IN), .B2(n4560), .ZN(n3158) );
  OAI21_X1 U3979 ( .B1(n3160), .B2(n4560), .A(n3158), .ZN(U3471) );
  INV_X1 U3980 ( .A(n4328), .ZN(n4253) );
  AOI22_X1 U3981 ( .A1(n4253), .A2(n3269), .B1(REG1_REG_2__SCAN_IN), .B2(n4567), .ZN(n3159) );
  OAI21_X1 U3982 ( .B1(n3160), .B2(n4567), .A(n3159), .ZN(U3520) );
  NAND2_X1 U3983 ( .A1(n3146), .A2(n3161), .ZN(n3207) );
  XNOR2_X1 U3984 ( .A(n3207), .B(n3885), .ZN(n3266) );
  OAI21_X1 U3985 ( .B1(n3885), .B2(n3163), .A(n3162), .ZN(n3164) );
  AOI22_X1 U3986 ( .A1(n3164), .A2(n4225), .B1(n4288), .B2(n3967), .ZN(n3261)
         );
  AOI22_X1 U3987 ( .A1(n3965), .A2(n4319), .B1(n4318), .B2(n3165), .ZN(n3166)
         );
  OAI211_X1 U3988 ( .C1(n4315), .C2(n3266), .A(n3261), .B(n3166), .ZN(n3174)
         );
  OR2_X1 U3989 ( .A1(n3167), .A2(n3260), .ZN(n3168) );
  NAND2_X1 U3990 ( .A1(n3168), .A2(n3217), .ZN(n3257) );
  INV_X1 U3991 ( .A(REG0_REG_3__SCAN_IN), .ZN(n3169) );
  OAI22_X1 U3992 ( .A1(n4389), .A2(n3257), .B1(n4562), .B2(n3169), .ZN(n3170)
         );
  AOI21_X1 U3993 ( .B1(n3174), .B2(n4562), .A(n3170), .ZN(n3171) );
  INV_X1 U3994 ( .A(n3171), .ZN(U3473) );
  OAI22_X1 U3995 ( .A1(n4328), .A2(n3257), .B1(n4569), .B2(n3172), .ZN(n3173)
         );
  AOI21_X1 U3996 ( .B1(n3174), .B2(n4569), .A(n3173), .ZN(n3175) );
  INV_X1 U3997 ( .A(n3175), .ZN(U3521) );
  XOR2_X1 U3998 ( .A(n3176), .B(n3177), .Z(n3182) );
  AOI21_X1 U3999 ( .B1(n3766), .B2(n3963), .A(n3178), .ZN(n3180) );
  AOI22_X1 U4000 ( .A1(n3769), .A2(n3965), .B1(n3768), .B2(n3230), .ZN(n3179)
         );
  OAI211_X1 U4001 ( .C1(n3773), .C2(n3233), .A(n3180), .B(n3179), .ZN(n3181)
         );
  AOI21_X1 U4002 ( .B1(n3182), .B2(n3775), .A(n3181), .ZN(n3183) );
  INV_X1 U4003 ( .A(n3183), .ZN(U3224) );
  INV_X1 U4004 ( .A(n3185), .ZN(n3187) );
  NAND2_X1 U4005 ( .A1(n3187), .A2(n3186), .ZN(n3188) );
  XNOR2_X1 U4006 ( .A(n3184), .B(n3188), .ZN(n3195) );
  OAI21_X1 U4007 ( .B1(n3753), .B2(n3354), .A(n3189), .ZN(n3190) );
  INV_X1 U4008 ( .A(n3190), .ZN(n3193) );
  AOI22_X1 U4009 ( .A1(n3769), .A2(n3964), .B1(n3768), .B2(n3191), .ZN(n3192)
         );
  OAI211_X1 U4010 ( .C1(n3773), .C2(n3251), .A(n3193), .B(n3192), .ZN(n3194)
         );
  AOI21_X1 U4011 ( .B1(n3195), .B2(n3775), .A(n3194), .ZN(n3196) );
  INV_X1 U4012 ( .A(n3196), .ZN(U3236) );
  NAND2_X1 U4013 ( .A1(n4514), .A2(n4036), .ZN(n4233) );
  INV_X1 U4014 ( .A(n4231), .ZN(n4547) );
  AND2_X1 U4015 ( .A1(n4514), .A2(n4319), .ZN(n4162) );
  OAI22_X1 U4016 ( .A1(n3248), .A2(n3198), .B1(n3197), .B2(n4511), .ZN(n3201)
         );
  MUX2_X1 U4017 ( .A(REG2_REG_1__SCAN_IN), .B(n3199), .S(n4514), .Z(n3200) );
  AOI211_X1 U4018 ( .C1(n4162), .C2(n3967), .A(n3201), .B(n3200), .ZN(n3203)
         );
  NAND2_X1 U4019 ( .A1(n4514), .A2(n4288), .ZN(n4048) );
  AOI22_X1 U4020 ( .A1(n4186), .A2(n2737), .B1(n4185), .B2(n2366), .ZN(n3202)
         );
  OAI211_X1 U4021 ( .C1(n4213), .C2(n3204), .A(n3203), .B(n3202), .ZN(U3289)
         );
  NAND2_X1 U4022 ( .A1(n3207), .A2(n3206), .ZN(n3209) );
  NAND2_X1 U4023 ( .A1(n3209), .A2(n3208), .ZN(n3210) );
  NAND2_X1 U4024 ( .A1(n3210), .A2(n2375), .ZN(n3211) );
  AND2_X1 U4025 ( .A1(n3205), .A2(n3211), .ZN(n4546) );
  INV_X1 U4026 ( .A(n4546), .ZN(n3223) );
  XOR2_X1 U4027 ( .A(n2375), .B(n3212), .Z(n3216) );
  AOI22_X1 U4028 ( .A1(n3966), .A2(n4288), .B1(n3718), .B2(n4318), .ZN(n3213)
         );
  OAI21_X1 U4029 ( .B1(n3716), .B2(n4331), .A(n3213), .ZN(n3214) );
  AOI21_X1 U4030 ( .B1(n4546), .B2(n3359), .A(n3214), .ZN(n3215) );
  OAI21_X1 U4031 ( .B1(n3216), .B2(n4302), .A(n3215), .ZN(n4544) );
  INV_X1 U4032 ( .A(n3217), .ZN(n3219) );
  OAI211_X1 U4033 ( .C1(n3219), .C2(n3218), .A(n4231), .B(n3231), .ZN(n4543)
         );
  OAI22_X1 U4034 ( .A1(n4543), .A2(n4395), .B1(n4511), .B2(n3719), .ZN(n3220)
         );
  OAI21_X1 U4035 ( .B1(n4544), .B2(n3220), .A(n4514), .ZN(n3222) );
  NAND2_X1 U4036 ( .A1(n4523), .A2(REG2_REG_4__SCAN_IN), .ZN(n3221) );
  OAI211_X1 U4037 ( .C1(n3223), .C2(n3248), .A(n3222), .B(n3221), .ZN(U3286)
         );
  INV_X1 U4038 ( .A(n3224), .ZN(n3815) );
  AND2_X1 U4039 ( .A1(n3815), .A2(n3826), .ZN(n3863) );
  NAND2_X1 U4040 ( .A1(n3205), .A2(n3225), .ZN(n3226) );
  XOR2_X1 U4041 ( .A(n3863), .B(n3226), .Z(n3294) );
  NAND2_X1 U4042 ( .A1(n3228), .A2(n3227), .ZN(n3229) );
  NAND2_X1 U40430 ( .A1(n4514), .A2(n3229), .ZN(n4218) );
  AND2_X1 U4044 ( .A1(n3231), .A2(n3230), .ZN(n3232) );
  NOR2_X1 U4045 ( .A1(n3250), .A2(n3232), .ZN(n3310) );
  AOI22_X1 U4046 ( .A1(n4186), .A2(n3965), .B1(n4162), .B2(n3963), .ZN(n3236)
         );
  INV_X1 U4047 ( .A(n3233), .ZN(n3234) );
  AOI22_X1 U4048 ( .A1(n4523), .A2(REG2_REG_5__SCAN_IN), .B1(n3234), .B2(n4188), .ZN(n3235) );
  OAI211_X1 U4049 ( .C1(n3289), .C2(n4166), .A(n3236), .B(n3235), .ZN(n3237)
         );
  AOI21_X1 U4050 ( .B1(n4517), .B2(n3310), .A(n3237), .ZN(n3241) );
  XNOR2_X1 U4051 ( .A(n3238), .B(n3863), .ZN(n3239) );
  NOR2_X1 U4052 ( .A1(n3239), .A2(n4302), .ZN(n3291) );
  NAND2_X1 U4053 ( .A1(n3291), .A2(n4514), .ZN(n3240) );
  OAI211_X1 U4054 ( .C1(n3294), .C2(n4218), .A(n3241), .B(n3240), .ZN(U3285)
         );
  AND2_X1 U4055 ( .A1(n3818), .A2(n3825), .ZN(n3884) );
  XOR2_X1 U4056 ( .A(n3884), .B(n3242), .Z(n3247) );
  OAI22_X1 U4057 ( .A1(n3354), .A2(n4331), .B1(n4330), .B2(n3249), .ZN(n3243)
         );
  AOI21_X1 U4058 ( .B1(n4288), .B2(n3964), .A(n3243), .ZN(n3246) );
  XNOR2_X1 U4059 ( .A(n3244), .B(n3884), .ZN(n4553) );
  NAND2_X1 U4060 ( .A1(n4553), .A2(n3359), .ZN(n3245) );
  OAI211_X1 U4061 ( .C1(n3247), .C2(n4302), .A(n3246), .B(n3245), .ZN(n4550)
         );
  INV_X1 U4062 ( .A(n4550), .ZN(n3256) );
  INV_X1 U4063 ( .A(n4514), .ZN(n4404) );
  INV_X1 U4064 ( .A(n3248), .ZN(n4518) );
  INV_X1 U4065 ( .A(n3281), .ZN(n4548) );
  NOR2_X1 U4066 ( .A1(n3250), .A2(n3249), .ZN(n4549) );
  NOR3_X1 U4067 ( .A1(n4213), .A2(n4548), .A3(n4549), .ZN(n3254) );
  INV_X1 U4068 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3252) );
  OAI22_X1 U4069 ( .A1(n4514), .A2(n3252), .B1(n3251), .B2(n4511), .ZN(n3253)
         );
  AOI211_X1 U4070 ( .C1(n4553), .C2(n4518), .A(n3254), .B(n3253), .ZN(n3255)
         );
  OAI21_X1 U4071 ( .B1(n3256), .B2(n4404), .A(n3255), .ZN(U3284) );
  INV_X1 U4072 ( .A(n3257), .ZN(n3264) );
  OAI22_X1 U4073 ( .A1(n4514), .A2(n3982), .B1(REG3_REG_3__SCAN_IN), .B2(n4511), .ZN(n3258) );
  AOI21_X1 U4074 ( .B1(n4162), .B2(n3965), .A(n3258), .ZN(n3259) );
  OAI21_X1 U4075 ( .B1(n3260), .B2(n4166), .A(n3259), .ZN(n3263) );
  NOR2_X1 U4076 ( .A1(n3261), .A2(n4404), .ZN(n3262) );
  AOI211_X1 U4077 ( .C1(n3264), .C2(n4517), .A(n3263), .B(n3262), .ZN(n3265)
         );
  OAI21_X1 U4078 ( .B1(n4218), .B2(n3266), .A(n3265), .ZN(U3287) );
  MUX2_X1 U4079 ( .A(REG2_REG_2__SCAN_IN), .B(n3267), .S(n4514), .Z(n3276) );
  AOI22_X1 U4080 ( .A1(n4186), .A2(n2370), .B1(n4185), .B2(n3268), .ZN(n3274)
         );
  NAND2_X1 U4081 ( .A1(n4517), .A2(n3269), .ZN(n3273) );
  AOI22_X1 U4082 ( .A1(n4518), .A2(n3270), .B1(REG3_REG_2__SCAN_IN), .B2(n4188), .ZN(n3272) );
  NAND2_X1 U4083 ( .A1(n4162), .A2(n3966), .ZN(n3271) );
  NAND4_X1 U4084 ( .A1(n3274), .A2(n3273), .A3(n3272), .A4(n3271), .ZN(n3275)
         );
  OR2_X1 U4085 ( .A1(n3276), .A2(n3275), .ZN(U3288) );
  XNOR2_X1 U4086 ( .A(n3277), .B(n3888), .ZN(n3280) );
  AOI22_X1 U4087 ( .A1(n3961), .A2(n4319), .B1(n4318), .B2(n3321), .ZN(n3278)
         );
  OAI21_X1 U4088 ( .B1(n3290), .B2(n4333), .A(n3278), .ZN(n3279) );
  AOI21_X1 U4089 ( .B1(n3280), .B2(n4225), .A(n3279), .ZN(n4559) );
  AOI21_X1 U4090 ( .B1(n3281), .B2(n3321), .A(n4547), .ZN(n3282) );
  NAND2_X1 U4091 ( .A1(n3282), .A2(n3362), .ZN(n4558) );
  INV_X1 U4092 ( .A(n4558), .ZN(n3285) );
  INV_X1 U4093 ( .A(n4233), .ZN(n3284) );
  OAI22_X1 U4094 ( .A1(n4514), .A2(n2408), .B1(n3324), .B2(n4511), .ZN(n3283)
         );
  AOI21_X1 U4095 ( .B1(n3285), .B2(n3284), .A(n3283), .ZN(n3288) );
  OR2_X1 U4096 ( .A1(n3286), .A2(n3888), .ZN(n4556) );
  NAND2_X1 U4097 ( .A1(n3286), .A2(n3888), .ZN(n4555) );
  NAND3_X1 U4098 ( .A1(n4556), .A2(n4555), .A3(n4237), .ZN(n3287) );
  OAI211_X1 U4099 ( .C1(n4559), .C2(n4523), .A(n3288), .B(n3287), .ZN(U3283)
         );
  OAI22_X1 U4100 ( .A1(n3290), .A2(n4331), .B1(n4330), .B2(n3289), .ZN(n3292)
         );
  AOI211_X1 U4101 ( .C1(n4288), .C2(n3965), .A(n3292), .B(n3291), .ZN(n3293)
         );
  OAI21_X1 U4102 ( .B1(n4315), .B2(n3294), .A(n3293), .ZN(n3309) );
  INV_X1 U4103 ( .A(n3309), .ZN(n3296) );
  AOI22_X1 U4104 ( .A1(n4351), .A2(n3310), .B1(REG0_REG_5__SCAN_IN), .B2(n4560), .ZN(n3295) );
  OAI21_X1 U4105 ( .B1(n3296), .B2(n4560), .A(n3295), .ZN(U3477) );
  XNOR2_X1 U4106 ( .A(n3299), .B(n3298), .ZN(n3300) );
  XNOR2_X1 U4107 ( .A(n3297), .B(n3300), .ZN(n3307) );
  OAI21_X1 U4108 ( .B1(n3753), .B2(n3302), .A(n3301), .ZN(n3303) );
  INV_X1 U4109 ( .A(n3303), .ZN(n3305) );
  AOI22_X1 U4110 ( .A1(n3769), .A2(n3962), .B1(n3768), .B2(n3363), .ZN(n3304)
         );
  OAI211_X1 U4111 ( .C1(n3773), .C2(n4512), .A(n3305), .B(n3304), .ZN(n3306)
         );
  AOI21_X1 U4112 ( .B1(n3307), .B2(n3775), .A(n3306), .ZN(n3308) );
  INV_X1 U4113 ( .A(n3308), .ZN(U3218) );
  NAND2_X1 U4114 ( .A1(n3309), .A2(n4569), .ZN(n3312) );
  NAND2_X1 U4115 ( .A1(n4253), .A2(n3310), .ZN(n3311) );
  OAI211_X1 U4116 ( .C1(n4569), .C2(n3313), .A(n3312), .B(n3311), .ZN(U3523)
         );
  INV_X1 U4117 ( .A(n3315), .ZN(n3316) );
  AOI211_X1 U4118 ( .C1(n3317), .C2(n3314), .A(n3759), .B(n3316), .ZN(n3326)
         );
  INV_X1 U4119 ( .A(n3318), .ZN(n3319) );
  OAI21_X1 U4120 ( .B1(n3753), .B2(n3406), .A(n3319), .ZN(n3320) );
  INV_X1 U4121 ( .A(n3320), .ZN(n3323) );
  AOI22_X1 U4122 ( .A1(n3769), .A2(n3963), .B1(n3768), .B2(n3321), .ZN(n3322)
         );
  OAI211_X1 U4123 ( .C1(n3773), .C2(n3324), .A(n3323), .B(n3322), .ZN(n3325)
         );
  OR2_X1 U4124 ( .A1(n3326), .A2(n3325), .ZN(U3210) );
  INV_X1 U4125 ( .A(n3836), .ZN(n3327) );
  AND2_X1 U4126 ( .A1(n3327), .A2(n3822), .ZN(n3864) );
  XOR2_X1 U4127 ( .A(n3864), .B(n3328), .Z(n3329) );
  NAND2_X1 U4128 ( .A1(n3329), .A2(n4225), .ZN(n3405) );
  INV_X1 U4129 ( .A(n3361), .ZN(n3330) );
  AOI21_X1 U4130 ( .B1(n3403), .B2(n3330), .A(n3372), .ZN(n3410) );
  INV_X1 U4131 ( .A(n4162), .ZN(n4192) );
  AOI22_X1 U4132 ( .A1(n4186), .A2(n3961), .B1(n4185), .B2(n3403), .ZN(n3331)
         );
  OAI21_X1 U4133 ( .B1(n3332), .B2(n4192), .A(n3331), .ZN(n3334) );
  OAI22_X1 U4134 ( .A1(n3346), .A2(n4511), .B1(n2435), .B2(n4514), .ZN(n3333)
         );
  AOI211_X1 U4135 ( .C1(n3410), .C2(n4517), .A(n3334), .B(n3333), .ZN(n3339)
         );
  NAND2_X1 U4136 ( .A1(n3336), .A2(n3335), .ZN(n3337) );
  XNOR2_X1 U4137 ( .A(n3337), .B(n3864), .ZN(n3408) );
  NAND2_X1 U4138 ( .A1(n3408), .A2(n4237), .ZN(n3338) );
  OAI211_X1 U4139 ( .C1(n3405), .C2(n4404), .A(n3339), .B(n3338), .ZN(U3281)
         );
  INV_X1 U4140 ( .A(n3341), .ZN(n3342) );
  AOI21_X1 U4141 ( .B1(n3343), .B2(n3340), .A(n3342), .ZN(n3349) );
  NOR2_X1 U4142 ( .A1(STATE_REG_SCAN_IN), .A2(n2430), .ZN(n4416) );
  AOI21_X1 U4143 ( .B1(n3766), .B2(n3959), .A(n4416), .ZN(n3345) );
  AOI22_X1 U4144 ( .A1(n3769), .A2(n3961), .B1(n3768), .B2(n3403), .ZN(n3344)
         );
  OAI211_X1 U4145 ( .C1(n3773), .C2(n3346), .A(n3345), .B(n3344), .ZN(n3347)
         );
  INV_X1 U4146 ( .A(n3347), .ZN(n3348) );
  OAI21_X1 U4147 ( .B1(n3349), .B2(n3759), .A(n3348), .ZN(U3228) );
  INV_X1 U4148 ( .A(REG0_REG_8__SCAN_IN), .ZN(n3366) );
  NAND2_X1 U4149 ( .A1(n4556), .A2(n3350), .ZN(n3351) );
  AND2_X1 U4150 ( .A1(n3821), .A2(n3824), .ZN(n3887) );
  XNOR2_X1 U4151 ( .A(n3351), .B(n3887), .ZN(n4519) );
  INV_X1 U4152 ( .A(n4519), .ZN(n3360) );
  XNOR2_X1 U4153 ( .A(n3352), .B(n3887), .ZN(n3357) );
  OAI22_X1 U4154 ( .A1(n3354), .A2(n4333), .B1(n3353), .B2(n4330), .ZN(n3355)
         );
  AOI21_X1 U4155 ( .B1(n4319), .B2(n3960), .A(n3355), .ZN(n3356) );
  OAI21_X1 U4156 ( .B1(n3357), .B2(n4302), .A(n3356), .ZN(n3358) );
  AOI21_X1 U4157 ( .B1(n3359), .B2(n4519), .A(n3358), .ZN(n4522) );
  OAI21_X1 U4158 ( .B1(n4540), .B2(n3360), .A(n4522), .ZN(n3367) );
  NAND2_X1 U4159 ( .A1(n3367), .A2(n4562), .ZN(n3365) );
  AOI21_X1 U4160 ( .B1(n3363), .B2(n3362), .A(n3361), .ZN(n4516) );
  NAND2_X1 U4161 ( .A1(n4516), .A2(n4351), .ZN(n3364) );
  OAI211_X1 U4162 ( .C1(n4562), .C2(n3366), .A(n3365), .B(n3364), .ZN(U3483)
         );
  NAND2_X1 U4163 ( .A1(n3367), .A2(n4569), .ZN(n3369) );
  NAND2_X1 U4164 ( .A1(n4516), .A2(n4253), .ZN(n3368) );
  OAI211_X1 U4165 ( .C1(n4569), .C2(n4012), .A(n3369), .B(n3368), .ZN(U3526)
         );
  AND2_X1 U4166 ( .A1(n3833), .A2(n3838), .ZN(n3868) );
  XOR2_X1 U4167 ( .A(n3868), .B(n3370), .Z(n3426) );
  NAND2_X1 U4168 ( .A1(n4514), .A2(n4225), .ZN(n4198) );
  XOR2_X1 U4169 ( .A(n3868), .B(n3371), .Z(n3428) );
  NAND2_X1 U4170 ( .A1(n3428), .A2(n4237), .ZN(n3380) );
  INV_X1 U4171 ( .A(n3372), .ZN(n3374) );
  INV_X1 U4172 ( .A(n3385), .ZN(n3373) );
  AOI21_X1 U4173 ( .B1(n3643), .B2(n3374), .A(n3373), .ZN(n3430) );
  AOI22_X1 U4174 ( .A1(n4186), .A2(n3960), .B1(n4185), .B2(n3643), .ZN(n3377)
         );
  INV_X1 U4175 ( .A(n3644), .ZN(n3375) );
  AOI22_X1 U4176 ( .A1(n4523), .A2(REG2_REG_10__SCAN_IN), .B1(n3375), .B2(
        n4188), .ZN(n3376) );
  OAI211_X1 U4177 ( .C1(n3546), .C2(n4192), .A(n3377), .B(n3376), .ZN(n3378)
         );
  AOI21_X1 U4178 ( .B1(n3430), .B2(n4517), .A(n3378), .ZN(n3379) );
  OAI211_X1 U4179 ( .C1(n3426), .C2(n4198), .A(n3380), .B(n3379), .ZN(U3280)
         );
  XNOR2_X1 U4180 ( .A(n3381), .B(n2470), .ZN(n3462) );
  NAND2_X1 U4181 ( .A1(n3382), .A2(n3881), .ZN(n3383) );
  NAND2_X1 U4182 ( .A1(n3384), .A2(n3383), .ZN(n3454) );
  NAND2_X1 U4183 ( .A1(n3385), .A2(n3455), .ZN(n3386) );
  NAND2_X1 U4184 ( .A1(n3491), .A2(n3386), .ZN(n3468) );
  OAI22_X1 U4185 ( .A1(n4514), .A2(n3387), .B1(n3399), .B2(n4511), .ZN(n3388)
         );
  AOI21_X1 U4186 ( .B1(n4162), .B2(n3957), .A(n3388), .ZN(n3390) );
  AOI22_X1 U4187 ( .A1(n4186), .A2(n3959), .B1(n4185), .B2(n3455), .ZN(n3389)
         );
  OAI211_X1 U4188 ( .C1(n3468), .C2(n4213), .A(n3390), .B(n3389), .ZN(n3391)
         );
  AOI21_X1 U4189 ( .B1(n3454), .B2(n4237), .A(n3391), .ZN(n3392) );
  OAI21_X1 U4190 ( .B1(n4198), .B2(n3462), .A(n3392), .ZN(U3279) );
  NAND2_X1 U4191 ( .A1(n3395), .A2(n3394), .ZN(n3396) );
  XNOR2_X1 U4192 ( .A(n3393), .B(n3396), .ZN(n3401) );
  AND2_X1 U4193 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4437) );
  AOI21_X1 U4194 ( .B1(n3766), .B2(n3957), .A(n4437), .ZN(n3398) );
  AOI22_X1 U4195 ( .A1(n3769), .A2(n3959), .B1(n3768), .B2(n3455), .ZN(n3397)
         );
  OAI211_X1 U4196 ( .C1(n3773), .C2(n3399), .A(n3398), .B(n3397), .ZN(n3400)
         );
  AOI21_X1 U4197 ( .B1(n3401), .B2(n3775), .A(n3400), .ZN(n3402) );
  INV_X1 U4198 ( .A(n3402), .ZN(U3233) );
  AOI22_X1 U4199 ( .A1(n3959), .A2(n4319), .B1(n4318), .B2(n3403), .ZN(n3404)
         );
  OAI211_X1 U4200 ( .C1(n3406), .C2(n4333), .A(n3405), .B(n3404), .ZN(n3407)
         );
  AOI21_X1 U4201 ( .B1(n3408), .B2(n4554), .A(n3407), .ZN(n3412) );
  AOI22_X1 U4202 ( .A1(n3410), .A2(n4253), .B1(REG1_REG_9__SCAN_IN), .B2(n4567), .ZN(n3409) );
  OAI21_X1 U4203 ( .B1(n3412), .B2(n4567), .A(n3409), .ZN(U3527) );
  AOI22_X1 U4204 ( .A1(n3410), .A2(n4351), .B1(REG0_REG_9__SCAN_IN), .B2(n4560), .ZN(n3411) );
  OAI21_X1 U4205 ( .B1(n3412), .B2(n4560), .A(n3411), .ZN(U3485) );
  XNOR2_X1 U4206 ( .A(n3415), .B(n3414), .ZN(n3416) );
  XNOR2_X1 U4207 ( .A(n3413), .B(n3416), .ZN(n3421) );
  NAND2_X1 U4208 ( .A1(REG3_REG_12__SCAN_IN), .A2(U3149), .ZN(n4441) );
  OAI21_X1 U4209 ( .B1(n3753), .B2(n3542), .A(n4441), .ZN(n3417) );
  INV_X1 U4210 ( .A(n3417), .ZN(n3419) );
  AOI22_X1 U4211 ( .A1(n3769), .A2(n3958), .B1(n3768), .B2(n3497), .ZN(n3418)
         );
  OAI211_X1 U4212 ( .C1(n3773), .C2(n3494), .A(n3419), .B(n3418), .ZN(n3420)
         );
  AOI21_X1 U4213 ( .B1(n3421), .B2(n3775), .A(n3420), .ZN(n3422) );
  INV_X1 U4214 ( .A(n3422), .ZN(U3221) );
  OAI22_X1 U4215 ( .A1(n3546), .A2(n4331), .B1(n4330), .B2(n3423), .ZN(n3424)
         );
  AOI21_X1 U4216 ( .B1(n4288), .B2(n3960), .A(n3424), .ZN(n3425) );
  OAI21_X1 U4217 ( .B1(n3426), .B2(n4302), .A(n3425), .ZN(n3427) );
  AOI21_X1 U4218 ( .B1(n4554), .B2(n3428), .A(n3427), .ZN(n3432) );
  AOI22_X1 U4219 ( .A1(n3430), .A2(n4253), .B1(REG1_REG_10__SCAN_IN), .B2(
        n4567), .ZN(n3429) );
  OAI21_X1 U4220 ( .B1(n3432), .B2(n4567), .A(n3429), .ZN(U3528) );
  AOI22_X1 U4221 ( .A1(n3430), .A2(n4351), .B1(REG0_REG_10__SCAN_IN), .B2(
        n4560), .ZN(n3431) );
  OAI21_X1 U4222 ( .B1(n3432), .B2(n4560), .A(n3431), .ZN(U3487) );
  XNOR2_X1 U4223 ( .A(n3908), .B(n3434), .ZN(n3560) );
  OAI21_X1 U4224 ( .B1(n3435), .B2(n3434), .A(n3433), .ZN(n3562) );
  NAND2_X1 U4225 ( .A1(n3562), .A2(n4237), .ZN(n3442) );
  OAI21_X1 U4226 ( .B1(n3480), .B2(n3557), .A(n3510), .ZN(n3568) );
  INV_X1 U4227 ( .A(n3568), .ZN(n3440) );
  AOI22_X1 U4228 ( .A1(n4186), .A2(n3956), .B1(n4185), .B2(n3526), .ZN(n3438)
         );
  INV_X1 U4229 ( .A(n3529), .ZN(n3436) );
  AOI22_X1 U4230 ( .A1(n4523), .A2(REG2_REG_14__SCAN_IN), .B1(n3436), .B2(
        n4188), .ZN(n3437) );
  OAI211_X1 U4231 ( .C1(n4334), .C2(n4192), .A(n3438), .B(n3437), .ZN(n3439)
         );
  AOI21_X1 U4232 ( .B1(n3440), .B2(n4517), .A(n3439), .ZN(n3441) );
  OAI211_X1 U4233 ( .C1(n3560), .C2(n4198), .A(n3442), .B(n3441), .ZN(U3276)
         );
  INV_X1 U4234 ( .A(n3444), .ZN(n3446) );
  NAND2_X1 U4235 ( .A1(n3446), .A2(n3445), .ZN(n3447) );
  XNOR2_X1 U4236 ( .A(n3443), .B(n3447), .ZN(n3452) );
  NOR2_X1 U4237 ( .A1(STATE_REG_SCAN_IN), .A2(n2326), .ZN(n4454) );
  AOI21_X1 U4238 ( .B1(n3766), .B2(n3955), .A(n4454), .ZN(n3450) );
  AOI22_X1 U4239 ( .A1(n3769), .A2(n3957), .B1(n3768), .B2(n3448), .ZN(n3449)
         );
  OAI211_X1 U4240 ( .C1(n3773), .C2(n3481), .A(n3450), .B(n3449), .ZN(n3451)
         );
  AOI21_X1 U4241 ( .B1(n3452), .B2(n3775), .A(n3451), .ZN(n3453) );
  INV_X1 U4242 ( .A(n3453), .ZN(U3231) );
  NAND2_X1 U4243 ( .A1(n3454), .A2(n4554), .ZN(n3461) );
  NAND2_X1 U4244 ( .A1(n3455), .A2(n4318), .ZN(n3457) );
  NAND2_X1 U4245 ( .A1(n3959), .A2(n4288), .ZN(n3456) );
  OAI211_X1 U4246 ( .C1(n3458), .C2(n4331), .A(n3457), .B(n3456), .ZN(n3459)
         );
  INV_X1 U4247 ( .A(n3459), .ZN(n3460) );
  OAI211_X1 U4248 ( .C1(n3462), .C2(n4302), .A(n3461), .B(n3460), .ZN(n3465)
         );
  MUX2_X1 U4249 ( .A(n3465), .B(REG0_REG_11__SCAN_IN), .S(n4560), .Z(n3463) );
  INV_X1 U4250 ( .A(n3463), .ZN(n3464) );
  OAI21_X1 U4251 ( .B1(n3468), .B2(n4389), .A(n3464), .ZN(U3489) );
  MUX2_X1 U4252 ( .A(REG1_REG_11__SCAN_IN), .B(n3465), .S(n4569), .Z(n3466) );
  INV_X1 U4253 ( .A(n3466), .ZN(n3467) );
  OAI21_X1 U4254 ( .B1(n4328), .B2(n3468), .A(n3467), .ZN(U3529) );
  OAI21_X1 U4255 ( .B1(n3501), .B2(n3488), .A(n3487), .ZN(n3472) );
  INV_X1 U4256 ( .A(n3469), .ZN(n3471) );
  OR2_X1 U4257 ( .A1(n3471), .A2(n3470), .ZN(n3476) );
  INV_X1 U4258 ( .A(n3476), .ZN(n3870) );
  XNOR2_X1 U4259 ( .A(n3472), .B(n3870), .ZN(n3475) );
  OAI22_X1 U4260 ( .A1(n3584), .A2(n4331), .B1(n4330), .B2(n3478), .ZN(n3473)
         );
  AOI21_X1 U4261 ( .B1(n4288), .B2(n3957), .A(n3473), .ZN(n3474) );
  OAI21_X1 U4262 ( .B1(n3475), .B2(n4302), .A(n3474), .ZN(n3533) );
  INV_X1 U4263 ( .A(n3533), .ZN(n3486) );
  XNOR2_X1 U4264 ( .A(n3477), .B(n3476), .ZN(n3534) );
  NOR2_X1 U4265 ( .A1(n3492), .A2(n3478), .ZN(n3479) );
  OR2_X1 U4266 ( .A1(n3480), .A2(n3479), .ZN(n3540) );
  INV_X1 U4267 ( .A(n3481), .ZN(n3482) );
  AOI22_X1 U4268 ( .A1(n4523), .A2(REG2_REG_13__SCAN_IN), .B1(n3482), .B2(
        n4188), .ZN(n3483) );
  OAI21_X1 U4269 ( .B1(n3540), .B2(n4213), .A(n3483), .ZN(n3484) );
  AOI21_X1 U4270 ( .B1(n3534), .B2(n4237), .A(n3484), .ZN(n3485) );
  OAI21_X1 U4271 ( .B1(n3486), .B2(n4404), .A(n3485), .ZN(U3277) );
  INV_X1 U4272 ( .A(n3487), .ZN(n3489) );
  OR2_X1 U4273 ( .A1(n3489), .A2(n3488), .ZN(n3500) );
  XNOR2_X1 U4274 ( .A(n3490), .B(n3500), .ZN(n3548) );
  AND2_X1 U4275 ( .A1(n3491), .A2(n3497), .ZN(n3493) );
  OR2_X1 U4276 ( .A1(n3493), .A2(n3492), .ZN(n3556) );
  OAI22_X1 U4277 ( .A1(n4514), .A2(n3495), .B1(n3494), .B2(n4511), .ZN(n3496)
         );
  AOI21_X1 U4278 ( .B1(n3497), .B2(n4185), .A(n3496), .ZN(n3499) );
  AOI22_X1 U4279 ( .A1(n4186), .A2(n3958), .B1(n4162), .B2(n3956), .ZN(n3498)
         );
  OAI211_X1 U4280 ( .C1(n3556), .C2(n4213), .A(n3499), .B(n3498), .ZN(n3504)
         );
  INV_X1 U4281 ( .A(n3500), .ZN(n3865) );
  XNOR2_X1 U4282 ( .A(n3501), .B(n3865), .ZN(n3502) );
  NAND2_X1 U4283 ( .A1(n3502), .A2(n4225), .ZN(n3545) );
  NOR2_X1 U4284 ( .A1(n3545), .A2(n4523), .ZN(n3503) );
  AOI211_X1 U4285 ( .C1(n4237), .C2(n3548), .A(n3504), .B(n3503), .ZN(n3505)
         );
  INV_X1 U4286 ( .A(n3505), .ZN(U3278) );
  AOI21_X1 U4287 ( .B1(n3506), .B2(n3883), .A(n4302), .ZN(n3508) );
  NAND2_X1 U4288 ( .A1(n3508), .A2(n3507), .ZN(n3583) );
  XNOR2_X1 U4289 ( .A(n3509), .B(n3883), .ZN(n3586) );
  NAND2_X1 U4290 ( .A1(n3586), .A2(n4237), .ZN(n3519) );
  INV_X1 U4291 ( .A(n3510), .ZN(n3511) );
  OAI21_X1 U4292 ( .B1(n3511), .B2(n3515), .A(n3573), .ZN(n3592) );
  INV_X1 U4293 ( .A(n3592), .ZN(n3517) );
  AOI22_X1 U4294 ( .A1(n4186), .A2(n3955), .B1(n4162), .B2(n3953), .ZN(n3514)
         );
  INV_X1 U4295 ( .A(n3772), .ZN(n3512) );
  AOI22_X1 U4296 ( .A1(n4523), .A2(REG2_REG_15__SCAN_IN), .B1(n3512), .B2(
        n4188), .ZN(n3513) );
  OAI211_X1 U4297 ( .C1(n3515), .C2(n4166), .A(n3514), .B(n3513), .ZN(n3516)
         );
  AOI21_X1 U4298 ( .B1(n3517), .B2(n4517), .A(n3516), .ZN(n3518) );
  OAI211_X1 U4299 ( .C1(n4404), .C2(n3583), .A(n3519), .B(n3518), .ZN(U3275)
         );
  XNOR2_X1 U4300 ( .A(n3522), .B(n3521), .ZN(n3523) );
  XNOR2_X1 U4301 ( .A(n3520), .B(n3523), .ZN(n3531) );
  NOR2_X1 U4302 ( .A1(n4573), .A2(STATE_REG_SCAN_IN), .ZN(n4464) );
  INV_X1 U4303 ( .A(n4464), .ZN(n3524) );
  OAI21_X1 U4304 ( .B1(n3753), .B2(n4334), .A(n3524), .ZN(n3525) );
  INV_X1 U4305 ( .A(n3525), .ZN(n3528) );
  AOI22_X1 U4306 ( .A1(n3769), .A2(n3956), .B1(n3768), .B2(n3526), .ZN(n3527)
         );
  OAI211_X1 U4307 ( .C1(n3773), .C2(n3529), .A(n3528), .B(n3527), .ZN(n3530)
         );
  AOI21_X1 U4308 ( .B1(n3531), .B2(n3775), .A(n3530), .ZN(n3532) );
  INV_X1 U4309 ( .A(n3532), .ZN(U3212) );
  AOI21_X1 U4310 ( .B1(n4554), .B2(n3534), .A(n3533), .ZN(n3537) );
  MUX2_X1 U4311 ( .A(n3535), .B(n3537), .S(n4569), .Z(n3536) );
  OAI21_X1 U4312 ( .B1(n4328), .B2(n3540), .A(n3536), .ZN(U3531) );
  INV_X1 U4313 ( .A(REG0_REG_13__SCAN_IN), .ZN(n3538) );
  MUX2_X1 U4314 ( .A(n3538), .B(n3537), .S(n4562), .Z(n3539) );
  OAI21_X1 U4315 ( .B1(n3540), .B2(n4389), .A(n3539), .ZN(U3493) );
  OAI22_X1 U4316 ( .A1(n3542), .A2(n4331), .B1(n4330), .B2(n3541), .ZN(n3543)
         );
  INV_X1 U4317 ( .A(n3543), .ZN(n3544) );
  OAI211_X1 U4318 ( .C1(n3546), .C2(n4333), .A(n3545), .B(n3544), .ZN(n3547)
         );
  INV_X1 U4319 ( .A(n3547), .ZN(n3550) );
  NAND2_X1 U4320 ( .A1(n3548), .A2(n4554), .ZN(n3549) );
  AND2_X1 U4321 ( .A1(n3550), .A2(n3549), .ZN(n3553) );
  INV_X1 U4322 ( .A(REG0_REG_12__SCAN_IN), .ZN(n3551) );
  MUX2_X1 U4323 ( .A(n3553), .B(n3551), .S(n4560), .Z(n3552) );
  OAI21_X1 U4324 ( .B1(n3556), .B2(n4389), .A(n3552), .ZN(U3491) );
  MUX2_X1 U4325 ( .A(n3554), .B(n3553), .S(n4569), .Z(n3555) );
  OAI21_X1 U4326 ( .B1(n4328), .B2(n3556), .A(n3555), .ZN(U3530) );
  INV_X1 U4327 ( .A(REG0_REG_14__SCAN_IN), .ZN(n3563) );
  OAI22_X1 U4328 ( .A1(n4334), .A2(n4331), .B1(n4330), .B2(n3557), .ZN(n3558)
         );
  AOI21_X1 U4329 ( .B1(n4288), .B2(n3956), .A(n3558), .ZN(n3559) );
  OAI21_X1 U4330 ( .B1(n3560), .B2(n4302), .A(n3559), .ZN(n3561) );
  AOI21_X1 U4331 ( .B1(n3562), .B2(n4554), .A(n3561), .ZN(n3565) );
  MUX2_X1 U4332 ( .A(n3563), .B(n3565), .S(n4562), .Z(n3564) );
  OAI21_X1 U4333 ( .B1(n3568), .B2(n4389), .A(n3564), .ZN(U3495) );
  MUX2_X1 U4334 ( .A(n3566), .B(n3565), .S(n4569), .Z(n3567) );
  OAI21_X1 U4335 ( .B1(n4328), .B2(n3568), .A(n3567), .ZN(U3532) );
  INV_X1 U4336 ( .A(n4514), .ZN(n4523) );
  OAI211_X1 U4337 ( .C1(n3570), .C2(n3889), .A(n3569), .B(n4225), .ZN(n4338)
         );
  AOI21_X1 U4338 ( .B1(n3889), .B2(n3572), .A(n3571), .ZN(n4341) );
  NAND2_X1 U4339 ( .A1(n4341), .A2(n4237), .ZN(n3581) );
  NAND2_X1 U4340 ( .A1(n3573), .A2(n3685), .ZN(n3574) );
  NAND2_X1 U4341 ( .A1(n3597), .A2(n3574), .ZN(n4339) );
  INV_X1 U4342 ( .A(n4339), .ZN(n3579) );
  AOI22_X1 U4343 ( .A1(n4186), .A2(n3954), .B1(n4162), .B2(n2506), .ZN(n3577)
         );
  INV_X1 U4344 ( .A(n3688), .ZN(n3575) );
  AOI22_X1 U4345 ( .A1(n4523), .A2(REG2_REG_16__SCAN_IN), .B1(n3575), .B2(
        n4188), .ZN(n3576) );
  OAI211_X1 U4346 ( .C1(n4329), .C2(n4166), .A(n3577), .B(n3576), .ZN(n3578)
         );
  AOI21_X1 U4347 ( .B1(n3579), .B2(n4517), .A(n3578), .ZN(n3580) );
  OAI211_X1 U4348 ( .C1(n4523), .C2(n4338), .A(n3581), .B(n3580), .ZN(U3274)
         );
  AOI22_X1 U4349 ( .A1(n3953), .A2(n4319), .B1(n4318), .B2(n3767), .ZN(n3582)
         );
  OAI211_X1 U4350 ( .C1(n3584), .C2(n4333), .A(n3583), .B(n3582), .ZN(n3585)
         );
  AOI21_X1 U4351 ( .B1(n3586), .B2(n4554), .A(n3585), .ZN(n3589) );
  MUX2_X1 U4352 ( .A(n3587), .B(n3589), .S(n4569), .Z(n3588) );
  OAI21_X1 U4353 ( .B1(n4328), .B2(n3592), .A(n3588), .ZN(U3533) );
  INV_X1 U4354 ( .A(REG0_REG_15__SCAN_IN), .ZN(n3590) );
  MUX2_X1 U4355 ( .A(n3590), .B(n3589), .S(n4562), .Z(n3591) );
  OAI21_X1 U4356 ( .B1(n3592), .B2(n4389), .A(n3591), .ZN(U3497) );
  INV_X1 U4357 ( .A(n3790), .ZN(n3593) );
  AND2_X1 U4358 ( .A1(n3593), .A2(n4199), .ZN(n3869) );
  INV_X1 U4359 ( .A(n3869), .ZN(n3594) );
  XNOR2_X1 U4360 ( .A(n3595), .B(n3594), .ZN(n3596) );
  NAND2_X1 U4361 ( .A1(n3596), .A2(n4225), .ZN(n4322) );
  XOR2_X1 U4362 ( .A(n3869), .B(n2065), .Z(n4325) );
  NAND2_X1 U4363 ( .A1(n4325), .A2(n4237), .ZN(n3607) );
  INV_X1 U4364 ( .A(n3597), .ZN(n3599) );
  INV_X1 U4365 ( .A(n4232), .ZN(n3598) );
  OAI21_X1 U4366 ( .B1(n3599), .B2(n3603), .A(n3598), .ZN(n4390) );
  INV_X1 U4367 ( .A(n4390), .ZN(n3605) );
  AOI22_X1 U4368 ( .A1(n4186), .A2(n3953), .B1(n4162), .B2(n4320), .ZN(n3602)
         );
  INV_X1 U4369 ( .A(n3698), .ZN(n3600) );
  AOI22_X1 U4370 ( .A1(n4523), .A2(REG2_REG_17__SCAN_IN), .B1(n3600), .B2(
        n4188), .ZN(n3601) );
  OAI211_X1 U4371 ( .C1(n3603), .C2(n4166), .A(n3602), .B(n3601), .ZN(n3604)
         );
  AOI21_X1 U4372 ( .B1(n3605), .B2(n4517), .A(n3604), .ZN(n3606) );
  OAI211_X1 U4373 ( .C1(n4523), .C2(n4322), .A(n3607), .B(n3606), .ZN(U3273)
         );
  INV_X1 U4374 ( .A(n3608), .ZN(n3617) );
  AOI22_X1 U4375 ( .A1(n4079), .A2(n4186), .B1(n4162), .B2(n3951), .ZN(n3612)
         );
  INV_X1 U4376 ( .A(n3609), .ZN(n3610) );
  AOI22_X1 U4377 ( .A1(n3610), .A2(n4188), .B1(REG2_REG_28__SCAN_IN), .B2(
        n4404), .ZN(n3611) );
  OAI211_X1 U4378 ( .C1(n3613), .C2(n4166), .A(n3612), .B(n3611), .ZN(n3616)
         );
  NOR2_X1 U4379 ( .A1(n3614), .A2(n4404), .ZN(n3615) );
  AOI211_X1 U4380 ( .C1(n4517), .C2(n3617), .A(n3616), .B(n3615), .ZN(n3618)
         );
  OAI21_X1 U4381 ( .B1(n3619), .B2(n4218), .A(n3618), .ZN(U3262) );
  AOI21_X1 U4382 ( .B1(n3622), .B2(n3621), .A(n3620), .ZN(n3627) );
  OAI22_X1 U4383 ( .A1(n3751), .A2(n4193), .B1(STATE_REG_SCAN_IN), .B2(n3623), 
        .ZN(n3625) );
  OAI22_X1 U4384 ( .A1(n3752), .A2(n4144), .B1(n4140), .B2(n3753), .ZN(n3624)
         );
  AOI211_X1 U4385 ( .C1(n3757), .C2(n4147), .A(n3625), .B(n3624), .ZN(n3626)
         );
  OAI21_X1 U4386 ( .B1(n3627), .B2(n3759), .A(n3626), .ZN(U3232) );
  INV_X1 U4387 ( .A(D_REG_0__SCAN_IN), .ZN(n3631) );
  AND2_X1 U4388 ( .A1(n4525), .A2(n3628), .ZN(n3630) );
  AOI22_X1 U4389 ( .A1(n4524), .A2(n3631), .B1(n3630), .B2(n3629), .ZN(U3458)
         );
  XNOR2_X1 U4390 ( .A(n3633), .B(n3632), .ZN(n3638) );
  INV_X1 U4391 ( .A(n3634), .ZN(n4062) );
  INV_X1 U4392 ( .A(n4097), .ZN(n4263) );
  OAI22_X1 U4393 ( .A1(n4263), .A2(n3751), .B1(STATE_REG_SCAN_IN), .B2(n4586), 
        .ZN(n3636) );
  OAI22_X1 U4394 ( .A1(n4049), .A2(n3753), .B1(n3752), .B2(n4247), .ZN(n3635)
         );
  AOI211_X1 U4395 ( .C1(n4062), .C2(n3757), .A(n3636), .B(n3635), .ZN(n3637)
         );
  OAI21_X1 U4396 ( .B1(n3638), .B2(n3759), .A(n3637), .ZN(U3211) );
  AND2_X1 U4397 ( .A1(n3341), .A2(n3639), .ZN(n3642) );
  OAI211_X1 U4398 ( .C1(n3642), .C2(n3641), .A(n3775), .B(n3640), .ZN(n3648)
         );
  NOR2_X1 U4399 ( .A1(STATE_REG_SCAN_IN), .A2(n4666), .ZN(n4425) );
  AOI21_X1 U4400 ( .B1(n3766), .B2(n3958), .A(n4425), .ZN(n3647) );
  AOI22_X1 U4401 ( .A1(n3769), .A2(n3960), .B1(n3768), .B2(n3643), .ZN(n3646)
         );
  OR2_X1 U4402 ( .A1(n3773), .A2(n3644), .ZN(n3645) );
  NAND4_X1 U4403 ( .A1(n3648), .A2(n3647), .A3(n3646), .A4(n3645), .ZN(U3214)
         );
  XNOR2_X1 U4404 ( .A(n3650), .B(n3649), .ZN(n3656) );
  NAND2_X1 U4405 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4035) );
  OAI21_X1 U4406 ( .B1(n3753), .B2(n3664), .A(n4035), .ZN(n3651) );
  INV_X1 U4407 ( .A(n3651), .ZN(n3654) );
  AOI22_X1 U4408 ( .A1(n3769), .A2(n4320), .B1(n3768), .B2(n3652), .ZN(n3653)
         );
  OAI211_X1 U4409 ( .C1(n3773), .C2(n4214), .A(n3654), .B(n3653), .ZN(n3655)
         );
  AOI21_X1 U4410 ( .B1(n3656), .B2(n3775), .A(n3655), .ZN(n3657) );
  INV_X1 U4411 ( .A(n3657), .ZN(U3216) );
  INV_X1 U4412 ( .A(n4163), .ZN(n3670) );
  XNOR2_X1 U4413 ( .A(n3660), .B(n3659), .ZN(n3661) );
  XNOR2_X1 U4414 ( .A(n3658), .B(n3661), .ZN(n3662) );
  NAND2_X1 U4415 ( .A1(n3662), .A2(n3775), .ZN(n3669) );
  NAND2_X1 U4416 ( .A1(n3768), .A2(n4287), .ZN(n3663) );
  OAI21_X1 U4417 ( .B1(n3664), .B2(n3751), .A(n3663), .ZN(n3667) );
  OAI22_X1 U4418 ( .A1(n4292), .A2(n3753), .B1(STATE_REG_SCAN_IN), .B2(n3665), 
        .ZN(n3666) );
  NOR2_X1 U4419 ( .A1(n3667), .A2(n3666), .ZN(n3668) );
  OAI211_X1 U4420 ( .C1(n3773), .C2(n3670), .A(n3669), .B(n3668), .ZN(U3220)
         );
  NOR2_X1 U4421 ( .A1(n2246), .A2(n3672), .ZN(n3673) );
  XNOR2_X1 U4422 ( .A(n3674), .B(n3673), .ZN(n3680) );
  INV_X1 U4423 ( .A(n3675), .ZN(n4098) );
  OAI22_X1 U4424 ( .A1(n3676), .A2(n3751), .B1(n3752), .B2(n4258), .ZN(n3678)
         );
  OAI22_X1 U4425 ( .A1(n4263), .A2(n3753), .B1(STATE_REG_SCAN_IN), .B2(n4603), 
        .ZN(n3677) );
  AOI211_X1 U4426 ( .C1(n4098), .C2(n3757), .A(n3678), .B(n3677), .ZN(n3679)
         );
  OAI21_X1 U4427 ( .B1(n3680), .B2(n3759), .A(n3679), .ZN(U3222) );
  OAI21_X1 U4428 ( .B1(n3761), .B2(n3764), .A(n3762), .ZN(n3681) );
  XOR2_X1 U4429 ( .A(n3682), .B(n3681), .Z(n3690) );
  NOR2_X1 U4430 ( .A1(n4605), .A2(STATE_REG_SCAN_IN), .ZN(n4483) );
  INV_X1 U4431 ( .A(n4483), .ZN(n3683) );
  OAI21_X1 U4432 ( .B1(n3753), .B2(n4332), .A(n3683), .ZN(n3684) );
  INV_X1 U4433 ( .A(n3684), .ZN(n3687) );
  AOI22_X1 U4434 ( .A1(n3769), .A2(n3954), .B1(n3768), .B2(n3685), .ZN(n3686)
         );
  OAI211_X1 U4435 ( .C1(n3773), .C2(n3688), .A(n3687), .B(n3686), .ZN(n3689)
         );
  AOI21_X1 U4436 ( .B1(n3690), .B2(n3775), .A(n3689), .ZN(n3691) );
  INV_X1 U4437 ( .A(n3691), .ZN(U3223) );
  XNOR2_X1 U4438 ( .A(n3693), .B(n3692), .ZN(n3694) );
  XNOR2_X1 U4439 ( .A(n3695), .B(n3694), .ZN(n3700) );
  AND2_X1 U4440 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4492) );
  AOI21_X1 U4441 ( .B1(n3766), .B2(n4320), .A(n4492), .ZN(n3697) );
  AOI22_X1 U4442 ( .A1(n3769), .A2(n3953), .B1(n3768), .B2(n4317), .ZN(n3696)
         );
  OAI211_X1 U4443 ( .C1(n3773), .C2(n3698), .A(n3697), .B(n3696), .ZN(n3699)
         );
  AOI21_X1 U4444 ( .B1(n3700), .B2(n3775), .A(n3699), .ZN(n3701) );
  INV_X1 U4445 ( .A(n3701), .ZN(U3225) );
  NAND2_X1 U4446 ( .A1(n2056), .A2(n3702), .ZN(n3704) );
  XNOR2_X1 U4447 ( .A(n3704), .B(n3703), .ZN(n3710) );
  INV_X1 U4448 ( .A(n3705), .ZN(n4113) );
  OAI22_X1 U4449 ( .A1(n4140), .A2(n3751), .B1(STATE_REG_SCAN_IN), .B2(n3706), 
        .ZN(n3708) );
  OAI22_X1 U4450 ( .A1(n4272), .A2(n3753), .B1(n3752), .B2(n4116), .ZN(n3707)
         );
  AOI211_X1 U4451 ( .C1(n4113), .C2(n3757), .A(n3708), .B(n3707), .ZN(n3709)
         );
  OAI21_X1 U4452 ( .B1(n3710), .B2(n3759), .A(n3709), .ZN(U3226) );
  AND2_X1 U4453 ( .A1(n3126), .A2(n3711), .ZN(n3714) );
  OAI211_X1 U4454 ( .C1(n3714), .C2(n3712), .A(n3775), .B(n3713), .ZN(n3723)
         );
  OAI21_X1 U4455 ( .B1(n3753), .B2(n3716), .A(n3715), .ZN(n3717) );
  INV_X1 U4456 ( .A(n3717), .ZN(n3722) );
  AOI22_X1 U4457 ( .A1(n3769), .A2(n3966), .B1(n3768), .B2(n3718), .ZN(n3721)
         );
  OR2_X1 U4458 ( .A1(n3773), .A2(n3719), .ZN(n3720) );
  NAND4_X1 U4459 ( .A1(n3723), .A2(n3722), .A3(n3721), .A4(n3720), .ZN(U3227)
         );
  INV_X1 U4460 ( .A(n3728), .ZN(n3724) );
  NOR2_X1 U4461 ( .A1(n3725), .A2(n3724), .ZN(n3730) );
  AOI21_X1 U4462 ( .B1(n3728), .B2(n3727), .A(n3726), .ZN(n3729) );
  OAI21_X1 U4463 ( .B1(n3730), .B2(n3729), .A(n3775), .ZN(n3735) );
  INV_X1 U4464 ( .A(n4222), .ZN(n4298) );
  NAND2_X1 U4465 ( .A1(n3768), .A2(n4184), .ZN(n3731) );
  OAI21_X1 U4466 ( .B1(n4298), .B2(n3751), .A(n3731), .ZN(n3733) );
  OAI22_X1 U4467 ( .A1(n3753), .A2(n4193), .B1(STATE_REG_SCAN_IN), .B2(n4571), 
        .ZN(n3732) );
  NOR2_X1 U4468 ( .A1(n3733), .A2(n3732), .ZN(n3734) );
  OAI211_X1 U4469 ( .C1(n3773), .C2(n4187), .A(n3735), .B(n3734), .ZN(U3230)
         );
  NOR2_X1 U4470 ( .A1(n2077), .A2(n3736), .ZN(n3737) );
  XNOR2_X1 U4471 ( .A(n3738), .B(n3737), .ZN(n3743) );
  NAND2_X1 U4472 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4498) );
  OAI21_X1 U4473 ( .B1(n3753), .B2(n4298), .A(n4498), .ZN(n3739) );
  INV_X1 U4474 ( .A(n3739), .ZN(n3741) );
  AOI22_X1 U4475 ( .A1(n3769), .A2(n2506), .B1(n3768), .B2(n4221), .ZN(n3740)
         );
  OAI211_X1 U4476 ( .C1(n3773), .C2(n4234), .A(n3741), .B(n3740), .ZN(n3742)
         );
  AOI21_X1 U4477 ( .B1(n3743), .B2(n3775), .A(n3742), .ZN(n3744) );
  INV_X1 U4478 ( .A(n3744), .ZN(U3235) );
  INV_X1 U4479 ( .A(n3745), .ZN(n3747) );
  NAND2_X1 U4480 ( .A1(n3747), .A2(n3746), .ZN(n3748) );
  XNOR2_X1 U4481 ( .A(n3749), .B(n3748), .ZN(n3760) );
  OAI22_X1 U4482 ( .A1(n4272), .A2(n3751), .B1(STATE_REG_SCAN_IN), .B2(n3750), 
        .ZN(n3756) );
  OAI22_X1 U4483 ( .A1(n3754), .A2(n3753), .B1(n3752), .B2(n4083), .ZN(n3755)
         );
  AOI211_X1 U4484 ( .C1(n4084), .C2(n3757), .A(n3756), .B(n3755), .ZN(n3758)
         );
  OAI21_X1 U4485 ( .B1(n3760), .B2(n3759), .A(n3758), .ZN(U3237) );
  INV_X1 U4486 ( .A(n3761), .ZN(n3763) );
  NAND2_X1 U4487 ( .A1(n3763), .A2(n3762), .ZN(n3765) );
  XNOR2_X1 U4488 ( .A(n3765), .B(n3764), .ZN(n3776) );
  AND2_X1 U4489 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4473) );
  AOI21_X1 U4490 ( .B1(n3766), .B2(n3953), .A(n4473), .ZN(n3771) );
  AOI22_X1 U4491 ( .A1(n3769), .A2(n3955), .B1(n3768), .B2(n3767), .ZN(n3770)
         );
  OAI211_X1 U4492 ( .C1(n3773), .C2(n3772), .A(n3771), .B(n3770), .ZN(n3774)
         );
  AOI21_X1 U4493 ( .B1(n3776), .B2(n3775), .A(n3774), .ZN(n3777) );
  INV_X1 U4494 ( .A(n3777), .ZN(U3238) );
  NAND2_X1 U4495 ( .A1(n3951), .A2(n3778), .ZN(n3779) );
  NAND2_X1 U4496 ( .A1(n3780), .A2(n3779), .ZN(n3926) );
  INV_X1 U4497 ( .A(n3926), .ZN(n3853) );
  NAND2_X1 U4498 ( .A1(n3782), .A2(n3781), .ZN(n3921) );
  NAND2_X1 U4499 ( .A1(n3853), .A2(n3921), .ZN(n3789) );
  INV_X1 U4500 ( .A(n3951), .ZN(n3788) );
  INV_X1 U4501 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4239) );
  NAND2_X1 U4502 ( .A1(n2361), .A2(REG2_REG_31__SCAN_IN), .ZN(n3785) );
  NAND2_X1 U4503 ( .A1(n2041), .A2(REG0_REG_31__SCAN_IN), .ZN(n3784) );
  OAI211_X1 U4504 ( .C1(n2527), .C2(n4239), .A(n3785), .B(n3784), .ZN(n4042)
         );
  NAND2_X1 U4505 ( .A1(n2089), .A2(DATAI_31_), .ZN(n4043) );
  NAND2_X1 U4506 ( .A1(n4042), .A2(n4043), .ZN(n3857) );
  NOR2_X1 U4507 ( .A1(n3786), .A2(n4574), .ZN(n4245) );
  INV_X1 U4508 ( .A(n4245), .ZN(n3931) );
  OR2_X1 U4509 ( .A1(n3950), .A2(n3931), .ZN(n3787) );
  NAND2_X1 U4510 ( .A1(n3857), .A2(n3787), .ZN(n3862) );
  AOI21_X1 U4511 ( .B1(n3788), .B2(n4051), .A(n3862), .ZN(n3922) );
  NAND2_X1 U4512 ( .A1(n3789), .A2(n3922), .ZN(n3927) );
  INV_X1 U4513 ( .A(n3927), .ZN(n3855) );
  NAND2_X1 U4514 ( .A1(n4079), .A2(n4247), .ZN(n3851) );
  NOR2_X1 U4515 ( .A1(n3893), .A2(n2106), .ZN(n3919) );
  NOR2_X1 U4516 ( .A1(n3791), .A2(n3790), .ZN(n3912) );
  INV_X1 U4517 ( .A(n3911), .ZN(n3844) );
  NAND2_X1 U4518 ( .A1(n3793), .A2(n3792), .ZN(n3800) );
  NAND2_X1 U4519 ( .A1(n3800), .A2(n3794), .ZN(n3906) );
  INV_X1 U4520 ( .A(n3840), .ZN(n3798) );
  NAND2_X1 U4521 ( .A1(n3795), .A2(n3794), .ZN(n3907) );
  INV_X1 U4522 ( .A(n3907), .ZN(n3796) );
  OAI211_X1 U4523 ( .C1(n3799), .C2(n3798), .A(n3797), .B(n3796), .ZN(n3842)
         );
  INV_X1 U4524 ( .A(n3800), .ZN(n3832) );
  INV_X1 U4525 ( .A(n3801), .ZN(n3804) );
  OAI211_X1 U4526 ( .C1(n4394), .C2(n3804), .A(n3803), .B(n3802), .ZN(n3805)
         );
  NAND3_X1 U4527 ( .A1(n3807), .A2(n3806), .A3(n3805), .ZN(n3808) );
  NAND3_X1 U4528 ( .A1(n3810), .A2(n3809), .A3(n3808), .ZN(n3811) );
  NAND3_X1 U4529 ( .A1(n3813), .A2(n3812), .A3(n3811), .ZN(n3814) );
  NAND4_X1 U4530 ( .A1(n3816), .A2(n3825), .A3(n3815), .A4(n3814), .ZN(n3817)
         );
  NAND3_X1 U4531 ( .A1(n3888), .A2(n3818), .A3(n3817), .ZN(n3819) );
  NAND3_X1 U4532 ( .A1(n3823), .A2(n3824), .A3(n3819), .ZN(n3820) );
  NAND3_X1 U4533 ( .A1(n3822), .A2(n3821), .A3(n3820), .ZN(n3831) );
  INV_X1 U4534 ( .A(n3823), .ZN(n3829) );
  INV_X1 U4535 ( .A(n3824), .ZN(n3828) );
  INV_X1 U4536 ( .A(n3825), .ZN(n3827) );
  NOR4_X1 U4537 ( .A1(n3829), .A2(n3828), .A3(n3827), .A4(n3826), .ZN(n3830)
         );
  AOI22_X1 U4538 ( .A1(n3832), .A2(n3831), .B1(n3830), .B2(n3906), .ZN(n3835)
         );
  INV_X1 U4539 ( .A(n3906), .ZN(n3834) );
  OAI22_X1 U4540 ( .A1(n3836), .A2(n3835), .B1(n3834), .B2(n3833), .ZN(n3837)
         );
  AND4_X1 U4541 ( .A1(n3840), .A2(n3839), .A3(n3838), .A4(n3837), .ZN(n3841)
         );
  AOI21_X1 U4542 ( .B1(n3906), .B2(n3842), .A(n3841), .ZN(n3843) );
  OAI21_X1 U4543 ( .B1(n3844), .B2(n3843), .A(n3909), .ZN(n3845) );
  AOI21_X1 U4544 ( .B1(n3912), .B2(n3845), .A(n2111), .ZN(n3846) );
  OAI21_X1 U4545 ( .B1(n4122), .B2(n3846), .A(n3915), .ZN(n3847) );
  NAND2_X1 U4546 ( .A1(n3848), .A2(n3847), .ZN(n3849) );
  NAND3_X1 U4547 ( .A1(n3923), .A2(n3919), .A3(n3849), .ZN(n3850) );
  NAND4_X1 U4548 ( .A1(n3853), .A2(n3852), .A3(n3851), .A4(n3850), .ZN(n3854)
         );
  NAND2_X1 U4549 ( .A1(n3855), .A2(n3854), .ZN(n3859) );
  NAND2_X1 U4550 ( .A1(n3950), .A2(n3931), .ZN(n3932) );
  OR2_X1 U4551 ( .A1(n4042), .A2(n4043), .ZN(n3856) );
  NAND2_X1 U4552 ( .A1(n3932), .A2(n3856), .ZN(n3861) );
  NAND2_X1 U4553 ( .A1(n3861), .A2(n3857), .ZN(n3858) );
  NAND2_X1 U4554 ( .A1(n3859), .A2(n3858), .ZN(n3942) );
  INV_X1 U4555 ( .A(n4066), .ZN(n3903) );
  NAND2_X1 U4556 ( .A1(n4073), .A2(n3860), .ZN(n4094) );
  INV_X1 U4557 ( .A(n4094), .ZN(n3900) );
  INV_X1 U4558 ( .A(n4149), .ZN(n3877) );
  NOR2_X1 U4559 ( .A1(n3862), .A2(n3861), .ZN(n3876) );
  INV_X1 U4560 ( .A(n4228), .ZN(n3866) );
  NAND4_X1 U4561 ( .A1(n3866), .A2(n3865), .A3(n3864), .A4(n3863), .ZN(n3872)
         );
  NAND2_X1 U4562 ( .A1(n3867), .A2(n4178), .ZN(n4204) );
  NAND4_X1 U4563 ( .A1(n3870), .A2(n4204), .A3(n3869), .A4(n3868), .ZN(n3871)
         );
  NOR2_X1 U4564 ( .A1(n3872), .A2(n3871), .ZN(n3875) );
  NAND2_X1 U4565 ( .A1(n3874), .A2(n3873), .ZN(n4179) );
  AND4_X1 U4566 ( .A1(n3877), .A2(n3876), .A3(n3875), .A4(n4179), .ZN(n3899)
         );
  NAND2_X1 U4567 ( .A1(n3879), .A2(n3878), .ZN(n4126) );
  NAND4_X1 U4568 ( .A1(n3882), .A2(n3881), .A3(n2375), .A4(n3880), .ZN(n3892)
         );
  INV_X1 U4569 ( .A(n3883), .ZN(n3886) );
  NAND4_X1 U4570 ( .A1(n2112), .A2(n3886), .A3(n3885), .A4(n3884), .ZN(n3891)
         );
  NAND4_X1 U4571 ( .A1(n3889), .A2(n3888), .A3(n4541), .A4(n3887), .ZN(n3890)
         );
  NOR4_X1 U4572 ( .A1(n4126), .A2(n3892), .A3(n3891), .A4(n3890), .ZN(n3898)
         );
  INV_X1 U4573 ( .A(n4089), .ZN(n3894) );
  OR2_X1 U4574 ( .A1(n3894), .A2(n3893), .ZN(n4108) );
  INV_X1 U4575 ( .A(n3895), .ZN(n4123) );
  NOR2_X1 U4576 ( .A1(n4123), .A2(n4122), .ZN(n4158) );
  INV_X1 U4577 ( .A(n4158), .ZN(n3896) );
  NOR2_X1 U4578 ( .A1(n4108), .A2(n3896), .ZN(n3897) );
  NAND4_X1 U4579 ( .A1(n3900), .A2(n3899), .A3(n3898), .A4(n3897), .ZN(n3901)
         );
  XNOR2_X1 U4580 ( .A(n4097), .B(n4083), .ZN(n4076) );
  NOR2_X1 U4581 ( .A1(n3901), .A2(n4076), .ZN(n3902) );
  AND4_X1 U4582 ( .A1(n3905), .A2(n3904), .A3(n3903), .A4(n3902), .ZN(n3937)
         );
  OAI21_X1 U4583 ( .B1(n3908), .B2(n3907), .A(n3906), .ZN(n3910) );
  NAND2_X1 U4584 ( .A1(n3910), .A2(n3909), .ZN(n3913) );
  NAND3_X1 U4585 ( .A1(n3913), .A2(n3912), .A3(n3911), .ZN(n3916) );
  NAND3_X1 U4586 ( .A1(n3916), .A2(n3915), .A3(n3914), .ZN(n3918) );
  NAND2_X1 U4587 ( .A1(n3918), .A2(n3917), .ZN(n3920) );
  AOI21_X1 U4588 ( .B1(n3920), .B2(n3919), .A(n4074), .ZN(n3930) );
  INV_X1 U4589 ( .A(n3921), .ZN(n3924) );
  NAND3_X1 U4590 ( .A1(n3924), .A2(n3923), .A3(n3922), .ZN(n3929) );
  NOR3_X1 U4591 ( .A1(n3926), .A2(n4066), .A3(n3925), .ZN(n3928) );
  OAI22_X1 U4592 ( .A1(n3930), .A2(n3929), .B1(n3928), .B2(n3927), .ZN(n3935)
         );
  OR2_X1 U4593 ( .A1(n4042), .A2(n3931), .ZN(n3934) );
  AOI21_X1 U4594 ( .B1(n3932), .B2(n4042), .A(n4043), .ZN(n3933) );
  AOI21_X1 U4595 ( .B1(n3935), .B2(n3934), .A(n3933), .ZN(n3936) );
  MUX2_X1 U4596 ( .A(n3937), .B(n3936), .S(n4394), .Z(n3938) );
  NOR2_X1 U4597 ( .A1(n3938), .A2(n2636), .ZN(n3940) );
  AOI21_X1 U4598 ( .B1(n2636), .B2(n3942), .A(n3940), .ZN(n3939) );
  MUX2_X1 U4599 ( .A(n3940), .B(n3939), .S(n4036), .Z(n3941) );
  AOI21_X1 U4600 ( .B1(n3943), .B2(n3942), .A(n3941), .ZN(n3949) );
  NAND2_X1 U4601 ( .A1(n3945), .A2(n3944), .ZN(n3946) );
  OAI211_X1 U4602 ( .C1(n4393), .C2(n3948), .A(n3946), .B(B_REG_SCAN_IN), .ZN(
        n3947) );
  OAI21_X1 U4603 ( .B1(n3949), .B2(n3948), .A(n3947), .ZN(U3239) );
  MUX2_X1 U4604 ( .A(DATAO_REG_31__SCAN_IN), .B(n4042), .S(U4043), .Z(U3581)
         );
  MUX2_X1 U4605 ( .A(DATAO_REG_30__SCAN_IN), .B(n3950), .S(U4043), .Z(U3580)
         );
  MUX2_X1 U4606 ( .A(DATAO_REG_29__SCAN_IN), .B(n3951), .S(U4043), .Z(U3579)
         );
  MUX2_X1 U4607 ( .A(DATAO_REG_28__SCAN_IN), .B(n4250), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U4608 ( .A(DATAO_REG_27__SCAN_IN), .B(n4079), .S(U4043), .Z(U3577)
         );
  MUX2_X1 U4609 ( .A(DATAO_REG_26__SCAN_IN), .B(n4097), .S(U4043), .Z(U3576)
         );
  MUX2_X1 U4610 ( .A(DATAO_REG_25__SCAN_IN), .B(n4112), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U4611 ( .A(DATAO_REG_24__SCAN_IN), .B(n4260), .S(U4043), .Z(U3574)
         );
  MUX2_X1 U4612 ( .A(n4269), .B(DATAO_REG_23__SCAN_IN), .S(n3952), .Z(U3573)
         );
  MUX2_X1 U4613 ( .A(DATAO_REG_22__SCAN_IN), .B(n4161), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U4614 ( .A(n4300), .B(DATAO_REG_21__SCAN_IN), .S(n3952), .Z(U3571)
         );
  MUX2_X1 U4615 ( .A(n4289), .B(DATAO_REG_20__SCAN_IN), .S(n3952), .Z(U3570)
         );
  MUX2_X1 U4616 ( .A(n4222), .B(DATAO_REG_19__SCAN_IN), .S(n3952), .Z(U3569)
         );
  MUX2_X1 U4617 ( .A(n4320), .B(DATAO_REG_18__SCAN_IN), .S(n3952), .Z(U3568)
         );
  MUX2_X1 U4618 ( .A(DATAO_REG_17__SCAN_IN), .B(n2506), .S(U4043), .Z(U3567)
         );
  MUX2_X1 U4619 ( .A(DATAO_REG_16__SCAN_IN), .B(n3953), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U4620 ( .A(DATAO_REG_15__SCAN_IN), .B(n3954), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U4621 ( .A(DATAO_REG_14__SCAN_IN), .B(n3955), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U4622 ( .A(DATAO_REG_13__SCAN_IN), .B(n3956), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U4623 ( .A(DATAO_REG_12__SCAN_IN), .B(n3957), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U4624 ( .A(DATAO_REG_11__SCAN_IN), .B(n3958), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U4625 ( .A(DATAO_REG_10__SCAN_IN), .B(n3959), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U4626 ( .A(DATAO_REG_9__SCAN_IN), .B(n3960), .S(U4043), .Z(U3559) );
  MUX2_X1 U4627 ( .A(DATAO_REG_8__SCAN_IN), .B(n3961), .S(U4043), .Z(U3558) );
  MUX2_X1 U4628 ( .A(DATAO_REG_7__SCAN_IN), .B(n3962), .S(U4043), .Z(U3557) );
  MUX2_X1 U4629 ( .A(DATAO_REG_6__SCAN_IN), .B(n3963), .S(U4043), .Z(U3556) );
  MUX2_X1 U4630 ( .A(DATAO_REG_5__SCAN_IN), .B(n3964), .S(U4043), .Z(U3555) );
  MUX2_X1 U4631 ( .A(DATAO_REG_4__SCAN_IN), .B(n3965), .S(U4043), .Z(U3554) );
  MUX2_X1 U4632 ( .A(DATAO_REG_3__SCAN_IN), .B(n3966), .S(U4043), .Z(U3553) );
  MUX2_X1 U4633 ( .A(DATAO_REG_2__SCAN_IN), .B(n3967), .S(U4043), .Z(U3552) );
  MUX2_X1 U4634 ( .A(DATAO_REG_1__SCAN_IN), .B(n2370), .S(U4043), .Z(U3551) );
  MUX2_X1 U4635 ( .A(DATAO_REG_0__SCAN_IN), .B(n2737), .S(U4043), .Z(U3550) );
  NAND2_X1 U4636 ( .A1(n3979), .A2(n4403), .ZN(n3978) );
  INV_X1 U4637 ( .A(n3968), .ZN(n3971) );
  OAI211_X1 U4638 ( .C1(n3971), .C2(n3970), .A(n4450), .B(n3969), .ZN(n3977)
         );
  OAI211_X1 U4639 ( .C1(n3974), .C2(n3973), .A(n4505), .B(n3972), .ZN(n3976)
         );
  AOI22_X1 U4640 ( .A1(n4503), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3975) );
  NAND4_X1 U4641 ( .A1(n3978), .A2(n3977), .A3(n3976), .A4(n3975), .ZN(U3241)
         );
  NAND2_X1 U4642 ( .A1(n3979), .A2(n4401), .ZN(n3988) );
  OAI211_X1 U4643 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3981), .A(n4505), .B(n3980), 
        .ZN(n3987) );
  AOI22_X1 U4644 ( .A1(n4503), .A2(ADDR_REG_3__SCAN_IN), .B1(
        REG3_REG_3__SCAN_IN), .B2(U3149), .ZN(n3986) );
  XNOR2_X1 U4645 ( .A(n3983), .B(n3982), .ZN(n3984) );
  NAND2_X1 U4646 ( .A1(n4450), .A2(n3984), .ZN(n3985) );
  NAND4_X1 U4647 ( .A1(n3988), .A2(n3987), .A3(n3986), .A4(n3985), .ZN(U3243)
         );
  INV_X1 U4648 ( .A(REG2_REG_19__SCAN_IN), .ZN(n3989) );
  MUX2_X1 U4649 ( .A(REG2_REG_19__SCAN_IN), .B(n3989), .S(n4395), .Z(n4005) );
  INV_X1 U4650 ( .A(n4006), .ZN(n4527) );
  INV_X1 U4651 ( .A(REG2_REG_18__SCAN_IN), .ZN(n3990) );
  AOI22_X1 U4652 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4527), .B1(n4006), .B2(
        n3990), .ZN(n4501) );
  NOR2_X1 U4653 ( .A1(n4029), .A2(REG2_REG_17__SCAN_IN), .ZN(n3991) );
  AOI21_X1 U4654 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4029), .A(n3991), .ZN(n4490) );
  NOR2_X1 U4655 ( .A1(n4449), .A2(n4531), .ZN(n4448) );
  NAND2_X1 U4656 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4533), .ZN(n3996) );
  INV_X1 U4657 ( .A(n4533), .ZN(n4435) );
  AOI22_X1 U4658 ( .A1(REG2_REG_11__SCAN_IN), .A2(n4533), .B1(n4435), .B2(
        n3387), .ZN(n4432) );
  AOI22_X1 U4659 ( .A1(n4009), .A2(REG2_REG_9__SCAN_IN), .B1(n2435), .B2(n4537), .ZN(n4412) );
  NAND2_X1 U4660 ( .A1(n4014), .A2(n3994), .ZN(n3995) );
  INV_X1 U4661 ( .A(n4014), .ZN(n4535) );
  XNOR2_X1 U4662 ( .A(n3994), .B(n4535), .ZN(n4421) );
  NAND2_X1 U4663 ( .A1(REG2_REG_10__SCAN_IN), .A2(n4421), .ZN(n4420) );
  NAND2_X1 U4664 ( .A1(n3995), .A2(n4420), .ZN(n4431) );
  NAND2_X1 U4665 ( .A1(n4018), .A2(n3997), .ZN(n3998) );
  NOR2_X1 U4666 ( .A1(n2145), .A2(n3999), .ZN(n4000) );
  NAND2_X1 U4667 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4007), .ZN(n4001) );
  OAI21_X1 U4668 ( .B1(REG2_REG_15__SCAN_IN), .B2(n4007), .A(n4001), .ZN(n4470) );
  NAND2_X1 U4669 ( .A1(n4002), .A2(n2133), .ZN(n4003) );
  INV_X1 U4670 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4479) );
  AOI21_X1 U4671 ( .B1(n4006), .B2(REG2_REG_18__SCAN_IN), .A(n4500), .ZN(n4004) );
  XOR2_X1 U4672 ( .A(n4005), .B(n4004), .Z(n4040) );
  AOI22_X1 U4673 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4006), .B1(n4527), .B2(
        n4031), .ZN(n4507) );
  NOR2_X1 U4674 ( .A1(n4029), .A2(REG1_REG_17__SCAN_IN), .ZN(n4030) );
  NAND2_X1 U4675 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4007), .ZN(n4025) );
  AOI22_X1 U4676 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4007), .B1(n4530), .B2(
        n3587), .ZN(n4476) );
  NAND2_X1 U4677 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4008), .ZN(n4021) );
  AOI22_X1 U4678 ( .A1(REG1_REG_13__SCAN_IN), .A2(n4008), .B1(n4531), .B2(
        n3535), .ZN(n4458) );
  NAND2_X1 U4679 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4533), .ZN(n4017) );
  AOI22_X1 U4680 ( .A1(REG1_REG_11__SCAN_IN), .A2(n4533), .B1(n4435), .B2(
        n2456), .ZN(n4429) );
  NAND2_X1 U4681 ( .A1(n4009), .A2(REG1_REG_9__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4682 ( .A1(n4009), .A2(REG1_REG_9__SCAN_IN), .B1(n2434), .B2(n4537), .ZN(n4410) );
  NAND2_X1 U4683 ( .A1(n4014), .A2(n4015), .ZN(n4016) );
  XNOR2_X1 U4684 ( .A(n4015), .B(n4535), .ZN(n4419) );
  NAND2_X1 U4685 ( .A1(REG1_REG_10__SCAN_IN), .A2(n4419), .ZN(n4418) );
  NAND2_X1 U4686 ( .A1(n4018), .A2(n4019), .ZN(n4020) );
  NAND2_X1 U4687 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4445), .ZN(n4444) );
  NAND2_X1 U4688 ( .A1(n4020), .A2(n4444), .ZN(n4457) );
  NAND2_X1 U4689 ( .A1(n4458), .A2(n4457), .ZN(n4456) );
  NAND2_X1 U4690 ( .A1(n4021), .A2(n4456), .ZN(n4023) );
  NAND2_X1 U4691 ( .A1(n4022), .A2(n4023), .ZN(n4024) );
  XNOR2_X1 U4692 ( .A(n4023), .B(n2145), .ZN(n4466) );
  NAND2_X1 U4693 ( .A1(REG1_REG_14__SCAN_IN), .A2(n4466), .ZN(n4465) );
  NAND2_X1 U4694 ( .A1(n4024), .A2(n4465), .ZN(n4475) );
  NAND2_X1 U4695 ( .A1(n4476), .A2(n4475), .ZN(n4474) );
  NOR2_X1 U4696 ( .A1(n4026), .A2(n4027), .ZN(n4028) );
  AOI22_X1 U4697 ( .A1(n4029), .A2(n4326), .B1(REG1_REG_17__SCAN_IN), .B2(
        n4528), .ZN(n4493) );
  NOR2_X1 U4698 ( .A1(n4030), .A2(n4495), .ZN(n4506) );
  NAND2_X1 U4699 ( .A1(n4507), .A2(n4506), .ZN(n4504) );
  OAI21_X1 U4700 ( .B1(n4031), .B2(n4527), .A(n4504), .ZN(n4033) );
  MUX2_X1 U4701 ( .A(n4310), .B(REG1_REG_19__SCAN_IN), .S(n4395), .Z(n4032) );
  XNOR2_X1 U4702 ( .A(n4033), .B(n4032), .ZN(n4038) );
  NAND2_X1 U4703 ( .A1(n4503), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4034) );
  OAI211_X1 U4704 ( .C1(n4510), .C2(n4036), .A(n4035), .B(n4034), .ZN(n4037)
         );
  AOI21_X1 U4705 ( .B1(n4038), .B2(n4505), .A(n4037), .ZN(n4039) );
  OAI21_X1 U4706 ( .B1(n4040), .B2(n4499), .A(n4039), .ZN(U3259) );
  XNOR2_X1 U4707 ( .A(n4242), .B(n4043), .ZN(n4346) );
  NAND2_X1 U4708 ( .A1(n4042), .A2(n4041), .ZN(n4243) );
  OAI21_X1 U4709 ( .B1(n4043), .B2(n4330), .A(n4243), .ZN(n4343) );
  NAND2_X1 U4710 ( .A1(n4514), .A2(n4343), .ZN(n4045) );
  NAND2_X1 U4711 ( .A1(n4523), .A2(REG2_REG_31__SCAN_IN), .ZN(n4044) );
  OAI211_X1 U4712 ( .C1(n4346), .C2(n4213), .A(n4045), .B(n4044), .ZN(U3260)
         );
  INV_X1 U4713 ( .A(n4046), .ZN(n4059) );
  INV_X1 U4714 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4047) );
  OAI22_X1 U4715 ( .A1(n4049), .A2(n4048), .B1(n4514), .B2(n4047), .ZN(n4050)
         );
  AOI21_X1 U4716 ( .B1(n4051), .B2(n4185), .A(n4050), .ZN(n4058) );
  INV_X1 U4717 ( .A(n4052), .ZN(n4056) );
  OAI22_X1 U4718 ( .A1(n4054), .A2(n4213), .B1(n4053), .B2(n4511), .ZN(n4055)
         );
  OAI21_X1 U4719 ( .B1(n4056), .B2(n4055), .A(n4514), .ZN(n4057) );
  OAI211_X1 U4720 ( .C1(n4059), .C2(n4218), .A(n4058), .B(n4057), .ZN(U3354)
         );
  XNOR2_X1 U4721 ( .A(n4060), .B(n4066), .ZN(n4252) );
  AOI21_X1 U4722 ( .B1(n4061), .B2(n4082), .A(n2049), .ZN(n4352) );
  AOI22_X1 U4723 ( .A1(n4250), .A2(n4162), .B1(n4186), .B2(n4097), .ZN(n4064)
         );
  AOI22_X1 U4724 ( .A1(n4062), .A2(n4188), .B1(REG2_REG_27__SCAN_IN), .B2(
        n4404), .ZN(n4063) );
  OAI211_X1 U4725 ( .C1(n4247), .C2(n4166), .A(n4064), .B(n4063), .ZN(n4065)
         );
  AOI21_X1 U4726 ( .B1(n4352), .B2(n4517), .A(n4065), .ZN(n4071) );
  NAND2_X1 U4727 ( .A1(n4067), .A2(n4066), .ZN(n4068) );
  AOI21_X1 U4728 ( .B1(n4069), .B2(n4068), .A(n4302), .ZN(n4248) );
  NAND2_X1 U4729 ( .A1(n4248), .A2(n4514), .ZN(n4070) );
  OAI211_X1 U4730 ( .C1(n4252), .C2(n4218), .A(n4071), .B(n4070), .ZN(U3263)
         );
  XNOR2_X1 U4731 ( .A(n4072), .B(n4076), .ZN(n4255) );
  INV_X1 U4732 ( .A(n4255), .ZN(n4088) );
  INV_X1 U4733 ( .A(n4090), .ZN(n4075) );
  OAI21_X1 U4734 ( .B1(n4075), .B2(n4074), .A(n4073), .ZN(n4077) );
  XNOR2_X1 U4735 ( .A(n4077), .B(n4076), .ZN(n4081) );
  OAI22_X1 U4736 ( .A1(n4272), .A2(n4333), .B1(n4083), .B2(n4330), .ZN(n4078)
         );
  AOI21_X1 U4737 ( .B1(n4079), .B2(n4319), .A(n4078), .ZN(n4080) );
  OAI21_X1 U4738 ( .B1(n4081), .B2(n4302), .A(n4080), .ZN(n4254) );
  OAI21_X1 U4739 ( .B1(n4095), .B2(n4083), .A(n4082), .ZN(n4356) );
  AOI22_X1 U4740 ( .A1(n4084), .A2(n4188), .B1(REG2_REG_26__SCAN_IN), .B2(
        n4404), .ZN(n4085) );
  OAI21_X1 U4741 ( .B1(n4356), .B2(n4213), .A(n4085), .ZN(n4086) );
  AOI21_X1 U4742 ( .B1(n4254), .B2(n4514), .A(n4086), .ZN(n4087) );
  OAI21_X1 U4743 ( .B1(n4088), .B2(n4218), .A(n4087), .ZN(U3264) );
  NAND2_X1 U4744 ( .A1(n4090), .A2(n4089), .ZN(n4091) );
  XNOR2_X1 U4745 ( .A(n4091), .B(n4094), .ZN(n4092) );
  NAND2_X1 U4746 ( .A1(n4092), .A2(n4225), .ZN(n4262) );
  XOR2_X1 U4747 ( .A(n4094), .B(n4093), .Z(n4265) );
  NAND2_X1 U4748 ( .A1(n4265), .A2(n4237), .ZN(n4104) );
  INV_X1 U4749 ( .A(n4095), .ZN(n4096) );
  OAI21_X1 U4750 ( .B1(n4110), .B2(n4258), .A(n4096), .ZN(n4360) );
  INV_X1 U4751 ( .A(n4360), .ZN(n4102) );
  AOI22_X1 U4752 ( .A1(n4097), .A2(n4162), .B1(n4186), .B2(n4260), .ZN(n4100)
         );
  AOI22_X1 U4753 ( .A1(n4098), .A2(n4188), .B1(REG2_REG_25__SCAN_IN), .B2(
        n4404), .ZN(n4099) );
  OAI211_X1 U4754 ( .C1(n4258), .C2(n4166), .A(n4100), .B(n4099), .ZN(n4101)
         );
  AOI21_X1 U4755 ( .B1(n4102), .B2(n4517), .A(n4101), .ZN(n4103) );
  OAI211_X1 U4756 ( .C1(n4523), .C2(n4262), .A(n4104), .B(n4103), .ZN(U3265)
         );
  INV_X1 U4757 ( .A(n4108), .ZN(n4105) );
  XNOR2_X1 U4758 ( .A(n4106), .B(n4105), .ZN(n4107) );
  NAND2_X1 U4759 ( .A1(n4107), .A2(n4225), .ZN(n4271) );
  XNOR2_X1 U4760 ( .A(n4109), .B(n4108), .ZN(n4274) );
  NAND2_X1 U4761 ( .A1(n4274), .A2(n4237), .ZN(n4120) );
  INV_X1 U4762 ( .A(n4110), .ZN(n4111) );
  OAI21_X1 U4763 ( .B1(n2095), .B2(n4116), .A(n4111), .ZN(n4364) );
  INV_X1 U4764 ( .A(n4364), .ZN(n4118) );
  AOI22_X1 U4765 ( .A1(n4112), .A2(n4162), .B1(n4186), .B2(n4269), .ZN(n4115)
         );
  AOI22_X1 U4766 ( .A1(n4523), .A2(REG2_REG_24__SCAN_IN), .B1(n4113), .B2(
        n4188), .ZN(n4114) );
  OAI211_X1 U4767 ( .C1(n4116), .C2(n4166), .A(n4115), .B(n4114), .ZN(n4117)
         );
  AOI21_X1 U4768 ( .B1(n4118), .B2(n4517), .A(n4117), .ZN(n4119) );
  OAI211_X1 U4769 ( .C1(n4523), .C2(n4271), .A(n4120), .B(n4119), .ZN(U3266)
         );
  XOR2_X1 U4770 ( .A(n4126), .B(n4121), .Z(n4278) );
  INV_X1 U4771 ( .A(n4278), .ZN(n4138) );
  INV_X1 U4772 ( .A(n4122), .ZN(n4124) );
  AOI21_X1 U4773 ( .B1(n4155), .B2(n4124), .A(n4123), .ZN(n4139) );
  OAI21_X1 U4774 ( .B1(n4139), .B2(n4149), .A(n4125), .ZN(n4127) );
  XNOR2_X1 U4775 ( .A(n4127), .B(n4126), .ZN(n4130) );
  OAI22_X1 U4776 ( .A1(n4292), .A2(n4333), .B1(n4330), .B2(n4132), .ZN(n4128)
         );
  AOI21_X1 U4777 ( .B1(n4260), .B2(n4319), .A(n4128), .ZN(n4129) );
  OAI21_X1 U4778 ( .B1(n4130), .B2(n4302), .A(n4129), .ZN(n4277) );
  OAI21_X1 U4779 ( .B1(n2090), .B2(n4132), .A(n4131), .ZN(n4368) );
  INV_X1 U4780 ( .A(n4133), .ZN(n4134) );
  AOI22_X1 U4781 ( .A1(n4523), .A2(REG2_REG_23__SCAN_IN), .B1(n4134), .B2(
        n4188), .ZN(n4135) );
  OAI21_X1 U4782 ( .B1(n4368), .B2(n4213), .A(n4135), .ZN(n4136) );
  AOI21_X1 U4783 ( .B1(n4277), .B2(n4514), .A(n4136), .ZN(n4137) );
  OAI21_X1 U4784 ( .B1(n4138), .B2(n4218), .A(n4137), .ZN(U3267) );
  XOR2_X1 U4785 ( .A(n4149), .B(n4139), .Z(n4143) );
  OAI22_X1 U4786 ( .A1(n4140), .A2(n4331), .B1(n4144), .B2(n4330), .ZN(n4141)
         );
  AOI21_X1 U4787 ( .B1(n4288), .B2(n4300), .A(n4141), .ZN(n4142) );
  OAI21_X1 U4788 ( .B1(n4143), .B2(n4302), .A(n4142), .ZN(n4282) );
  OR2_X1 U4789 ( .A1(n4159), .A2(n4144), .ZN(n4145) );
  NAND2_X1 U4790 ( .A1(n4146), .A2(n4145), .ZN(n4372) );
  AOI22_X1 U4791 ( .A1(n4523), .A2(REG2_REG_22__SCAN_IN), .B1(n4147), .B2(
        n4188), .ZN(n4148) );
  OAI21_X1 U4792 ( .B1(n4372), .B2(n4213), .A(n4148), .ZN(n4153) );
  NOR2_X1 U4793 ( .A1(n4150), .A2(n4149), .ZN(n4281) );
  INV_X1 U4794 ( .A(n4283), .ZN(n4151) );
  NOR3_X1 U4795 ( .A1(n4281), .A2(n4151), .A3(n4218), .ZN(n4152) );
  AOI211_X1 U4796 ( .C1(n4514), .C2(n4282), .A(n4153), .B(n4152), .ZN(n4154)
         );
  INV_X1 U4797 ( .A(n4154), .ZN(U3268) );
  XNOR2_X1 U4798 ( .A(n4155), .B(n4158), .ZN(n4156) );
  NAND2_X1 U4799 ( .A1(n4156), .A2(n4225), .ZN(n4291) );
  XOR2_X1 U4800 ( .A(n4158), .B(n4157), .Z(n4294) );
  NAND2_X1 U4801 ( .A1(n4294), .A2(n4237), .ZN(n4171) );
  INV_X1 U4802 ( .A(n4159), .ZN(n4160) );
  OAI21_X1 U4803 ( .B1(n4181), .B2(n4167), .A(n4160), .ZN(n4376) );
  INV_X1 U4804 ( .A(n4376), .ZN(n4169) );
  AOI22_X1 U4805 ( .A1(n4186), .A2(n4289), .B1(n4162), .B2(n4161), .ZN(n4165)
         );
  AOI22_X1 U4806 ( .A1(n4523), .A2(REG2_REG_21__SCAN_IN), .B1(n4163), .B2(
        n4188), .ZN(n4164) );
  OAI211_X1 U4807 ( .C1(n4167), .C2(n4166), .A(n4165), .B(n4164), .ZN(n4168)
         );
  AOI21_X1 U4808 ( .B1(n4169), .B2(n4517), .A(n4168), .ZN(n4170) );
  OAI211_X1 U4809 ( .C1(n4523), .C2(n4291), .A(n4171), .B(n4170), .ZN(U3269)
         );
  INV_X1 U4810 ( .A(n4200), .ZN(n4174) );
  AOI21_X1 U4811 ( .B1(n4174), .B2(n4173), .A(n4172), .ZN(n4175) );
  XNOR2_X1 U4812 ( .A(n4175), .B(n4179), .ZN(n4303) );
  AOI21_X1 U4813 ( .B1(n4176), .B2(n4178), .A(n4177), .ZN(n4180) );
  XNOR2_X1 U4814 ( .A(n4180), .B(n4179), .ZN(n4305) );
  NAND2_X1 U4815 ( .A1(n4305), .A2(n4237), .ZN(n4197) );
  INV_X1 U4816 ( .A(n4210), .ZN(n4183) );
  INV_X1 U4817 ( .A(n4181), .ZN(n4182) );
  OAI21_X1 U4818 ( .B1(n4183), .B2(n4297), .A(n4182), .ZN(n4380) );
  INV_X1 U4819 ( .A(n4380), .ZN(n4195) );
  AOI22_X1 U4820 ( .A1(n4186), .A2(n4222), .B1(n4185), .B2(n4184), .ZN(n4191)
         );
  INV_X1 U4821 ( .A(n4187), .ZN(n4189) );
  AOI22_X1 U4822 ( .A1(n4523), .A2(REG2_REG_20__SCAN_IN), .B1(n4189), .B2(
        n4188), .ZN(n4190) );
  OAI211_X1 U4823 ( .C1(n4193), .C2(n4192), .A(n4191), .B(n4190), .ZN(n4194)
         );
  AOI21_X1 U4824 ( .B1(n4195), .B2(n4517), .A(n4194), .ZN(n4196) );
  OAI211_X1 U4825 ( .C1(n4303), .C2(n4198), .A(n4197), .B(n4196), .ZN(U3270)
         );
  XOR2_X1 U4826 ( .A(n4204), .B(n4176), .Z(n4309) );
  INV_X1 U4827 ( .A(n4309), .ZN(n4219) );
  NAND2_X1 U4828 ( .A1(n4200), .A2(n4199), .ZN(n4220) );
  INV_X1 U4829 ( .A(n4201), .ZN(n4203) );
  OAI21_X1 U4830 ( .B1(n4220), .B2(n4203), .A(n4202), .ZN(n4205) );
  XNOR2_X1 U4831 ( .A(n4205), .B(n4204), .ZN(n4209) );
  OAI22_X1 U4832 ( .A1(n4206), .A2(n4333), .B1(n4330), .B2(n4211), .ZN(n4207)
         );
  AOI21_X1 U4833 ( .B1(n4289), .B2(n4319), .A(n4207), .ZN(n4208) );
  OAI21_X1 U4834 ( .B1(n4209), .B2(n4302), .A(n4208), .ZN(n4308) );
  INV_X1 U4835 ( .A(n4230), .ZN(n4212) );
  OAI21_X1 U4836 ( .B1(n4212), .B2(n4211), .A(n4210), .ZN(n4384) );
  NOR2_X1 U4837 ( .A1(n4384), .A2(n4213), .ZN(n4216) );
  OAI22_X1 U4838 ( .A1(n4514), .A2(n3989), .B1(n4214), .B2(n4511), .ZN(n4215)
         );
  AOI211_X1 U4839 ( .C1(n4308), .C2(n4514), .A(n4216), .B(n4215), .ZN(n4217)
         );
  OAI21_X1 U4840 ( .B1(n4219), .B2(n4218), .A(n4217), .ZN(U3271) );
  XOR2_X1 U4841 ( .A(n4228), .B(n4220), .Z(n4226) );
  AOI22_X1 U4842 ( .A1(n4222), .A2(n4319), .B1(n4221), .B2(n4318), .ZN(n4223)
         );
  OAI21_X1 U4843 ( .B1(n4332), .B2(n4333), .A(n4223), .ZN(n4224) );
  AOI21_X1 U4844 ( .B1(n4226), .B2(n4225), .A(n4224), .ZN(n4314) );
  OAI21_X1 U4845 ( .B1(n4229), .B2(n4228), .A(n4227), .ZN(n4312) );
  OAI211_X1 U4846 ( .C1(n4232), .C2(n2522), .A(n4231), .B(n4230), .ZN(n4313)
         );
  NOR2_X1 U4847 ( .A1(n4313), .A2(n4233), .ZN(n4236) );
  OAI22_X1 U4848 ( .A1(n4514), .A2(n3990), .B1(n4234), .B2(n4511), .ZN(n4235)
         );
  AOI211_X1 U4849 ( .C1(n4312), .C2(n4237), .A(n4236), .B(n4235), .ZN(n4238)
         );
  OAI21_X1 U4850 ( .B1(n4404), .B2(n4314), .A(n4238), .ZN(U3272) );
  NOR2_X1 U4851 ( .A1(n4569), .A2(n4239), .ZN(n4240) );
  AOI21_X1 U4852 ( .B1(n4569), .B2(n4343), .A(n4240), .ZN(n4241) );
  OAI21_X1 U4853 ( .B1(n4346), .B2(n4328), .A(n4241), .ZN(U3549) );
  AOI21_X1 U4854 ( .B1(n4245), .B2(n2051), .A(n4242), .ZN(n4405) );
  INV_X1 U4855 ( .A(n4405), .ZN(n4349) );
  INV_X1 U4856 ( .A(n4243), .ZN(n4244) );
  AOI21_X1 U4857 ( .B1(n4245), .B2(n4318), .A(n4244), .ZN(n4407) );
  MUX2_X1 U4858 ( .A(n2671), .B(n4407), .S(n4569), .Z(n4246) );
  OAI21_X1 U4859 ( .B1(n4349), .B2(n4328), .A(n4246), .ZN(U3548) );
  OAI22_X1 U4860 ( .A1(n4263), .A2(n4333), .B1(n4247), .B2(n4330), .ZN(n4249)
         );
  AOI21_X1 U4861 ( .B1(n4255), .B2(n4554), .A(n4254), .ZN(n4353) );
  MUX2_X1 U4862 ( .A(n4256), .B(n4353), .S(n4569), .Z(n4257) );
  OAI21_X1 U4863 ( .B1(n4328), .B2(n4356), .A(n4257), .ZN(U3544) );
  INV_X1 U4864 ( .A(n4258), .ZN(n4259) );
  AOI22_X1 U4865 ( .A1(n4260), .A2(n4288), .B1(n4259), .B2(n4318), .ZN(n4261)
         );
  OAI211_X1 U4866 ( .C1(n4263), .C2(n4331), .A(n4262), .B(n4261), .ZN(n4264)
         );
  AOI21_X1 U4867 ( .B1(n4265), .B2(n4554), .A(n4264), .ZN(n4357) );
  MUX2_X1 U4868 ( .A(n4266), .B(n4357), .S(n4569), .Z(n4267) );
  OAI21_X1 U4869 ( .B1(n4328), .B2(n4360), .A(n4267), .ZN(U3543) );
  AOI22_X1 U4870 ( .A1(n4269), .A2(n4288), .B1(n4318), .B2(n4268), .ZN(n4270)
         );
  OAI211_X1 U4871 ( .C1(n4272), .C2(n4331), .A(n4271), .B(n4270), .ZN(n4273)
         );
  AOI21_X1 U4872 ( .B1(n4274), .B2(n4554), .A(n4273), .ZN(n4361) );
  MUX2_X1 U4873 ( .A(n4275), .B(n4361), .S(n4569), .Z(n4276) );
  OAI21_X1 U4874 ( .B1(n4328), .B2(n4364), .A(n4276), .ZN(U3542) );
  AOI21_X1 U4875 ( .B1(n4278), .B2(n4554), .A(n4277), .ZN(n4365) );
  MUX2_X1 U4876 ( .A(n4279), .B(n4365), .S(n4569), .Z(n4280) );
  OAI21_X1 U4877 ( .B1(n4328), .B2(n4368), .A(n4280), .ZN(U3541) );
  NOR2_X1 U4878 ( .A1(n4281), .A2(n4315), .ZN(n4284) );
  AOI21_X1 U4879 ( .B1(n4284), .B2(n4283), .A(n4282), .ZN(n4369) );
  MUX2_X1 U4880 ( .A(n4285), .B(n4369), .S(n4569), .Z(n4286) );
  OAI21_X1 U4881 ( .B1(n4328), .B2(n4372), .A(n4286), .ZN(U3540) );
  AOI22_X1 U4882 ( .A1(n4289), .A2(n4288), .B1(n4287), .B2(n4318), .ZN(n4290)
         );
  OAI211_X1 U4883 ( .C1(n4292), .C2(n4331), .A(n4291), .B(n4290), .ZN(n4293)
         );
  AOI21_X1 U4884 ( .B1(n4294), .B2(n4554), .A(n4293), .ZN(n4373) );
  MUX2_X1 U4885 ( .A(n4295), .B(n4373), .S(n4569), .Z(n4296) );
  OAI21_X1 U4886 ( .B1(n4328), .B2(n4376), .A(n4296), .ZN(U3539) );
  OAI22_X1 U4887 ( .A1(n4298), .A2(n4333), .B1(n4297), .B2(n4330), .ZN(n4299)
         );
  AOI21_X1 U4888 ( .B1(n4319), .B2(n4300), .A(n4299), .ZN(n4301) );
  OAI21_X1 U4889 ( .B1(n4303), .B2(n4302), .A(n4301), .ZN(n4304) );
  AOI21_X1 U4890 ( .B1(n4305), .B2(n4554), .A(n4304), .ZN(n4377) );
  MUX2_X1 U4891 ( .A(n4306), .B(n4377), .S(n4569), .Z(n4307) );
  OAI21_X1 U4892 ( .B1(n4328), .B2(n4380), .A(n4307), .ZN(U3538) );
  AOI21_X1 U4893 ( .B1(n4309), .B2(n4554), .A(n4308), .ZN(n4381) );
  MUX2_X1 U4894 ( .A(n4310), .B(n4381), .S(n4569), .Z(n4311) );
  OAI21_X1 U4895 ( .B1(n4328), .B2(n4384), .A(n4311), .ZN(U3537) );
  INV_X1 U4896 ( .A(n4312), .ZN(n4316) );
  OAI211_X1 U4897 ( .C1(n4316), .C2(n4315), .A(n4314), .B(n4313), .ZN(n4385)
         );
  MUX2_X1 U4898 ( .A(REG1_REG_18__SCAN_IN), .B(n4385), .S(n4569), .Z(U3536) );
  AOI22_X1 U4899 ( .A1(n4320), .A2(n4319), .B1(n4318), .B2(n4317), .ZN(n4321)
         );
  OAI211_X1 U4900 ( .C1(n4323), .C2(n4333), .A(n4322), .B(n4321), .ZN(n4324)
         );
  AOI21_X1 U4901 ( .B1(n4325), .B2(n4554), .A(n4324), .ZN(n4386) );
  MUX2_X1 U4902 ( .A(n4326), .B(n4386), .S(n4569), .Z(n4327) );
  OAI21_X1 U4903 ( .B1(n4328), .B2(n4390), .A(n4327), .ZN(U3535) );
  OAI22_X1 U4904 ( .A1(n4332), .A2(n4331), .B1(n4330), .B2(n4329), .ZN(n4336)
         );
  NOR2_X1 U4905 ( .A1(n4334), .A2(n4333), .ZN(n4335) );
  NOR2_X1 U4906 ( .A1(n4336), .A2(n4335), .ZN(n4337) );
  OAI211_X1 U4907 ( .C1(n4547), .C2(n4339), .A(n4338), .B(n4337), .ZN(n4340)
         );
  AOI21_X1 U4908 ( .B1(n4341), .B2(n4554), .A(n4340), .ZN(n4342) );
  INV_X1 U4909 ( .A(n4342), .ZN(n4391) );
  MUX2_X1 U4910 ( .A(REG1_REG_16__SCAN_IN), .B(n4391), .S(n4569), .Z(U3534) );
  NAND2_X1 U4911 ( .A1(n4562), .A2(n4343), .ZN(n4345) );
  NAND2_X1 U4912 ( .A1(n4560), .A2(REG0_REG_31__SCAN_IN), .ZN(n4344) );
  OAI211_X1 U4913 ( .C1(n4346), .C2(n4389), .A(n4345), .B(n4344), .ZN(U3517)
         );
  INV_X1 U4914 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4347) );
  MUX2_X1 U4915 ( .A(n4347), .B(n4407), .S(n4562), .Z(n4348) );
  OAI21_X1 U4916 ( .B1(n4349), .B2(n4389), .A(n4348), .ZN(U3516) );
  INV_X1 U4917 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4354) );
  MUX2_X1 U4918 ( .A(n4354), .B(n4353), .S(n4562), .Z(n4355) );
  OAI21_X1 U4919 ( .B1(n4356), .B2(n4389), .A(n4355), .ZN(U3512) );
  INV_X1 U4920 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4358) );
  MUX2_X1 U4921 ( .A(n4358), .B(n4357), .S(n4562), .Z(n4359) );
  OAI21_X1 U4922 ( .B1(n4360), .B2(n4389), .A(n4359), .ZN(U3511) );
  INV_X1 U4923 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4362) );
  MUX2_X1 U4924 ( .A(n4362), .B(n4361), .S(n4562), .Z(n4363) );
  OAI21_X1 U4925 ( .B1(n4364), .B2(n4389), .A(n4363), .ZN(U3510) );
  INV_X1 U4926 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4366) );
  MUX2_X1 U4927 ( .A(n4366), .B(n4365), .S(n4562), .Z(n4367) );
  OAI21_X1 U4928 ( .B1(n4368), .B2(n4389), .A(n4367), .ZN(U3509) );
  INV_X1 U4929 ( .A(REG0_REG_22__SCAN_IN), .ZN(n4370) );
  MUX2_X1 U4930 ( .A(n4370), .B(n4369), .S(n4562), .Z(n4371) );
  OAI21_X1 U4931 ( .B1(n4372), .B2(n4389), .A(n4371), .ZN(U3508) );
  INV_X1 U4932 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4374) );
  MUX2_X1 U4933 ( .A(n4374), .B(n4373), .S(n4562), .Z(n4375) );
  OAI21_X1 U4934 ( .B1(n4376), .B2(n4389), .A(n4375), .ZN(U3507) );
  INV_X1 U4935 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4378) );
  MUX2_X1 U4936 ( .A(n4378), .B(n4377), .S(n4562), .Z(n4379) );
  OAI21_X1 U4937 ( .B1(n4380), .B2(n4389), .A(n4379), .ZN(U3506) );
  INV_X1 U4938 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4382) );
  MUX2_X1 U4939 ( .A(n4382), .B(n4381), .S(n4562), .Z(n4383) );
  OAI21_X1 U4940 ( .B1(n4384), .B2(n4389), .A(n4383), .ZN(U3505) );
  MUX2_X1 U4941 ( .A(REG0_REG_18__SCAN_IN), .B(n4385), .S(n4562), .Z(U3503) );
  INV_X1 U4942 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4387) );
  MUX2_X1 U4943 ( .A(n4387), .B(n4386), .S(n4562), .Z(n4388) );
  OAI21_X1 U4944 ( .B1(n4390), .B2(n4389), .A(n4388), .ZN(U3501) );
  MUX2_X1 U4945 ( .A(REG0_REG_16__SCAN_IN), .B(n4391), .S(n4562), .Z(U3499) );
  MUX2_X1 U4946 ( .A(n4392), .B(DATAI_28_), .S(U3149), .Z(U3324) );
  MUX2_X1 U4947 ( .A(DATAI_24_), .B(n2686), .S(STATE_REG_SCAN_IN), .Z(U3328)
         );
  MUX2_X1 U4948 ( .A(DATAI_22_), .B(n4393), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U4949 ( .A(DATAI_21_), .B(n4394), .S(STATE_REG_SCAN_IN), .Z(U3331)
         );
  MUX2_X1 U4950 ( .A(n4395), .B(DATAI_19_), .S(U3149), .Z(U3333) );
  MUX2_X1 U4951 ( .A(DATAI_8_), .B(n2099), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U4952 ( .A(n4397), .B(DATAI_7_), .S(U3149), .Z(U3345) );
  MUX2_X1 U4953 ( .A(n4398), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U4954 ( .A(n4399), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U4955 ( .A(DATAI_4_), .B(n4400), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U4956 ( .A(n4401), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U4957 ( .A(n4402), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U4958 ( .A(n4403), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  AOI22_X1 U4959 ( .A1(n4405), .A2(n4517), .B1(REG2_REG_30__SCAN_IN), .B2(
        n4404), .ZN(n4406) );
  OAI21_X1 U4960 ( .B1(n4523), .B2(n4407), .A(n4406), .ZN(U3261) );
  OAI211_X1 U4961 ( .C1(n4410), .C2(n4409), .A(n4505), .B(n4408), .ZN(n4414)
         );
  OAI211_X1 U4962 ( .C1(n4412), .C2(n2048), .A(n4450), .B(n4411), .ZN(n4413)
         );
  OAI211_X1 U4963 ( .C1(n4510), .C2(n4537), .A(n4414), .B(n4413), .ZN(n4415)
         );
  AOI211_X1 U4964 ( .C1(n4503), .C2(ADDR_REG_9__SCAN_IN), .A(n4416), .B(n4415), 
        .ZN(n4417) );
  INV_X1 U4965 ( .A(n4417), .ZN(U3249) );
  OAI211_X1 U4966 ( .C1(REG1_REG_10__SCAN_IN), .C2(n4419), .A(n4505), .B(n4418), .ZN(n4423) );
  OAI211_X1 U4967 ( .C1(REG2_REG_10__SCAN_IN), .C2(n4421), .A(n4450), .B(n4420), .ZN(n4422) );
  OAI211_X1 U4968 ( .C1(n4510), .C2(n4535), .A(n4423), .B(n4422), .ZN(n4424)
         );
  AOI211_X1 U4969 ( .C1(n4503), .C2(ADDR_REG_10__SCAN_IN), .A(n4425), .B(n4424), .ZN(n4426) );
  INV_X1 U4970 ( .A(n4426), .ZN(U3250) );
  OAI211_X1 U4971 ( .C1(n4429), .C2(n4428), .A(n4505), .B(n4427), .ZN(n4434)
         );
  OAI211_X1 U4972 ( .C1(n4432), .C2(n4431), .A(n4450), .B(n4430), .ZN(n4433)
         );
  OAI211_X1 U4973 ( .C1(n4510), .C2(n4435), .A(n4434), .B(n4433), .ZN(n4436)
         );
  AOI211_X1 U4974 ( .C1(n4503), .C2(ADDR_REG_11__SCAN_IN), .A(n4437), .B(n4436), .ZN(n4438) );
  INV_X1 U4975 ( .A(n4438), .ZN(U3251) );
  OAI211_X1 U4976 ( .C1(REG2_REG_12__SCAN_IN), .C2(n4440), .A(n4450), .B(n4439), .ZN(n4442) );
  NAND2_X1 U4977 ( .A1(n4442), .A2(n4441), .ZN(n4443) );
  AOI21_X1 U4978 ( .B1(n4503), .B2(ADDR_REG_12__SCAN_IN), .A(n4443), .ZN(n4447) );
  OAI211_X1 U4979 ( .C1(REG1_REG_12__SCAN_IN), .C2(n4445), .A(n4505), .B(n4444), .ZN(n4446) );
  OAI211_X1 U4980 ( .C1(n4510), .C2(n4532), .A(n4447), .B(n4446), .ZN(U3252)
         );
  AOI21_X1 U4981 ( .B1(n4449), .B2(n4531), .A(n4448), .ZN(n4453) );
  OAI21_X1 U4982 ( .B1(n4453), .B2(n4452), .A(n4450), .ZN(n4451) );
  AOI21_X1 U4983 ( .B1(n4453), .B2(n4452), .A(n4451), .ZN(n4455) );
  AOI211_X1 U4984 ( .C1(n4503), .C2(ADDR_REG_13__SCAN_IN), .A(n4455), .B(n4454), .ZN(n4460) );
  OAI211_X1 U4985 ( .C1(n4458), .C2(n4457), .A(n4505), .B(n4456), .ZN(n4459)
         );
  OAI211_X1 U4986 ( .C1(n4510), .C2(n4531), .A(n4460), .B(n4459), .ZN(U3253)
         );
  AOI211_X1 U4987 ( .C1(n2487), .C2(n4462), .A(n4461), .B(n4499), .ZN(n4463)
         );
  AOI211_X1 U4988 ( .C1(n4503), .C2(ADDR_REG_14__SCAN_IN), .A(n4464), .B(n4463), .ZN(n4468) );
  OAI211_X1 U4989 ( .C1(REG1_REG_14__SCAN_IN), .C2(n4466), .A(n4505), .B(n4465), .ZN(n4467) );
  OAI211_X1 U4990 ( .C1(n4510), .C2(n2145), .A(n4468), .B(n4467), .ZN(U3254)
         );
  AOI211_X1 U4991 ( .C1(n4471), .C2(n4470), .A(n4469), .B(n4499), .ZN(n4472)
         );
  AOI211_X1 U4992 ( .C1(n4503), .C2(ADDR_REG_15__SCAN_IN), .A(n4473), .B(n4472), .ZN(n4478) );
  OAI211_X1 U4993 ( .C1(n4476), .C2(n4475), .A(n4505), .B(n4474), .ZN(n4477)
         );
  OAI211_X1 U4994 ( .C1(n4510), .C2(n4530), .A(n4478), .B(n4477), .ZN(U3255)
         );
  AOI221_X1 U4995 ( .B1(n4481), .B2(n4480), .C1(n4479), .C2(n4480), .A(n4499), 
        .ZN(n4482) );
  AOI211_X1 U4996 ( .C1(n4503), .C2(ADDR_REG_16__SCAN_IN), .A(n4483), .B(n4482), .ZN(n4487) );
  OAI221_X1 U4997 ( .B1(n4485), .B2(REG1_REG_16__SCAN_IN), .C1(n4485), .C2(
        n4484), .A(n4505), .ZN(n4486) );
  OAI211_X1 U4998 ( .C1(n4510), .C2(n2133), .A(n4487), .B(n4486), .ZN(U3256)
         );
  AOI221_X1 U4999 ( .B1(n4490), .B2(n4489), .C1(n4488), .C2(n4489), .A(n4499), 
        .ZN(n4491) );
  AOI211_X1 U5000 ( .C1(n4503), .C2(ADDR_REG_17__SCAN_IN), .A(n4492), .B(n4491), .ZN(n4497) );
  OAI221_X1 U5001 ( .B1(n4495), .B2(n4494), .C1(n4495), .C2(n4493), .A(n4505), 
        .ZN(n4496) );
  OAI211_X1 U5002 ( .C1(n4510), .C2(n4528), .A(n4497), .B(n4496), .ZN(U3257)
         );
  INV_X1 U5003 ( .A(n4498), .ZN(n4502) );
  OAI211_X1 U5004 ( .C1(n4507), .C2(n4506), .A(n4505), .B(n4504), .ZN(n4508)
         );
  OAI211_X1 U5005 ( .C1(n4510), .C2(n4527), .A(n4509), .B(n4508), .ZN(U3258)
         );
  OAI22_X1 U5006 ( .A1(n4514), .A2(n4513), .B1(n4512), .B2(n4511), .ZN(n4515)
         );
  INV_X1 U5007 ( .A(n4515), .ZN(n4521) );
  AOI22_X1 U5008 ( .A1(n4519), .A2(n4518), .B1(n4517), .B2(n4516), .ZN(n4520)
         );
  OAI211_X1 U5009 ( .C1(n4523), .C2(n4522), .A(n4521), .B(n4520), .ZN(U3282)
         );
  AND2_X1 U5010 ( .A1(D_REG_31__SCAN_IN), .A2(n4524), .ZN(U3291) );
  AND2_X1 U5011 ( .A1(D_REG_30__SCAN_IN), .A2(n4524), .ZN(U3292) );
  AND2_X1 U5012 ( .A1(D_REG_29__SCAN_IN), .A2(n4524), .ZN(U3293) );
  AND2_X1 U5013 ( .A1(D_REG_28__SCAN_IN), .A2(n4524), .ZN(U3294) );
  AND2_X1 U5014 ( .A1(D_REG_27__SCAN_IN), .A2(n4524), .ZN(U3295) );
  AND2_X1 U5015 ( .A1(D_REG_26__SCAN_IN), .A2(n4524), .ZN(U3296) );
  AND2_X1 U5016 ( .A1(D_REG_25__SCAN_IN), .A2(n4524), .ZN(U3297) );
  AND2_X1 U5017 ( .A1(D_REG_24__SCAN_IN), .A2(n4524), .ZN(U3298) );
  AND2_X1 U5018 ( .A1(D_REG_23__SCAN_IN), .A2(n4524), .ZN(U3299) );
  AND2_X1 U5019 ( .A1(D_REG_22__SCAN_IN), .A2(n4524), .ZN(U3300) );
  AND2_X1 U5020 ( .A1(D_REG_21__SCAN_IN), .A2(n4524), .ZN(U3301) );
  AND2_X1 U5021 ( .A1(D_REG_20__SCAN_IN), .A2(n4524), .ZN(U3302) );
  AND2_X1 U5022 ( .A1(D_REG_19__SCAN_IN), .A2(n4524), .ZN(U3303) );
  AND2_X1 U5023 ( .A1(D_REG_18__SCAN_IN), .A2(n4524), .ZN(U3304) );
  AND2_X1 U5024 ( .A1(D_REG_17__SCAN_IN), .A2(n4524), .ZN(U3305) );
  AND2_X1 U5025 ( .A1(D_REG_16__SCAN_IN), .A2(n4524), .ZN(U3306) );
  AND2_X1 U5026 ( .A1(D_REG_15__SCAN_IN), .A2(n4524), .ZN(U3307) );
  AND2_X1 U5027 ( .A1(D_REG_14__SCAN_IN), .A2(n4524), .ZN(U3308) );
  AND2_X1 U5028 ( .A1(D_REG_13__SCAN_IN), .A2(n4524), .ZN(U3309) );
  AND2_X1 U5029 ( .A1(D_REG_12__SCAN_IN), .A2(n4524), .ZN(U3310) );
  AND2_X1 U5030 ( .A1(D_REG_11__SCAN_IN), .A2(n4524), .ZN(U3311) );
  AND2_X1 U5031 ( .A1(D_REG_10__SCAN_IN), .A2(n4524), .ZN(U3312) );
  AND2_X1 U5032 ( .A1(D_REG_9__SCAN_IN), .A2(n4524), .ZN(U3313) );
  AND2_X1 U5033 ( .A1(D_REG_8__SCAN_IN), .A2(n4524), .ZN(U3314) );
  AND2_X1 U5034 ( .A1(D_REG_7__SCAN_IN), .A2(n4524), .ZN(U3315) );
  AND2_X1 U5035 ( .A1(D_REG_6__SCAN_IN), .A2(n4524), .ZN(U3316) );
  AND2_X1 U5036 ( .A1(D_REG_5__SCAN_IN), .A2(n4524), .ZN(U3317) );
  AND2_X1 U5037 ( .A1(D_REG_4__SCAN_IN), .A2(n4524), .ZN(U3318) );
  AND2_X1 U5038 ( .A1(D_REG_3__SCAN_IN), .A2(n4524), .ZN(U3319) );
  AND2_X1 U5039 ( .A1(D_REG_2__SCAN_IN), .A2(n4524), .ZN(U3320) );
  INV_X1 U5040 ( .A(DATAI_23_), .ZN(n4601) );
  AOI21_X1 U5041 ( .B1(U3149), .B2(n4601), .A(n4525), .ZN(U3329) );
  INV_X1 U5042 ( .A(DATAI_18_), .ZN(n4526) );
  AOI22_X1 U5043 ( .A1(STATE_REG_SCAN_IN), .A2(n4527), .B1(n4526), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5044 ( .A1(STATE_REG_SCAN_IN), .A2(n4528), .B1(n2505), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5045 ( .A(DATAI_16_), .ZN(n4529) );
  AOI22_X1 U5046 ( .A1(STATE_REG_SCAN_IN), .A2(n2133), .B1(n4529), .B2(U3149), 
        .ZN(U3336) );
  AOI22_X1 U5047 ( .A1(STATE_REG_SCAN_IN), .A2(n4530), .B1(n4672), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5048 ( .A(DATAI_14_), .ZN(n4670) );
  AOI22_X1 U5049 ( .A1(STATE_REG_SCAN_IN), .A2(n2145), .B1(n4670), .B2(U3149), 
        .ZN(U3338) );
  AOI22_X1 U5050 ( .A1(STATE_REG_SCAN_IN), .A2(n4531), .B1(n4691), .B2(U3149), 
        .ZN(U3339) );
  AOI22_X1 U5051 ( .A1(STATE_REG_SCAN_IN), .A2(n4532), .B1(n2481), .B2(U3149), 
        .ZN(U3340) );
  OAI22_X1 U5052 ( .A1(U3149), .A2(n4533), .B1(DATAI_11_), .B2(
        STATE_REG_SCAN_IN), .ZN(n4534) );
  INV_X1 U5053 ( .A(n4534), .ZN(U3341) );
  INV_X1 U5054 ( .A(DATAI_10_), .ZN(n4743) );
  AOI22_X1 U5055 ( .A1(STATE_REG_SCAN_IN), .A2(n4535), .B1(n4743), .B2(U3149), 
        .ZN(U3342) );
  INV_X1 U5056 ( .A(DATAI_9_), .ZN(n4536) );
  AOI22_X1 U5057 ( .A1(STATE_REG_SCAN_IN), .A2(n4537), .B1(n4536), .B2(U3149), 
        .ZN(U3343) );
  OAI211_X1 U5058 ( .C1(n4541), .C2(n4540), .A(n4539), .B(n4538), .ZN(n4542)
         );
  INV_X1 U5059 ( .A(n4542), .ZN(n4564) );
  AOI22_X1 U5060 ( .A1(n4562), .A2(n4564), .B1(n2367), .B2(n4560), .ZN(U3467)
         );
  INV_X1 U5061 ( .A(n4543), .ZN(n4545) );
  AOI211_X1 U5062 ( .C1(n4546), .C2(n4552), .A(n4545), .B(n4544), .ZN(n4565)
         );
  AOI22_X1 U5063 ( .A1(n4562), .A2(n4565), .B1(n2336), .B2(n4560), .ZN(U3475)
         );
  NOR3_X1 U5064 ( .A1(n4549), .A2(n4548), .A3(n4547), .ZN(n4551) );
  AOI211_X1 U5065 ( .C1(n4553), .C2(n4552), .A(n4551), .B(n4550), .ZN(n4566)
         );
  AOI22_X1 U5066 ( .A1(n4562), .A2(n4566), .B1(n2393), .B2(n4560), .ZN(U3479)
         );
  NAND3_X1 U5067 ( .A1(n4556), .A2(n4555), .A3(n4554), .ZN(n4557) );
  AND3_X1 U5068 ( .A1(n4559), .A2(n4558), .A3(n4557), .ZN(n4568) );
  INV_X1 U5069 ( .A(REG0_REG_7__SCAN_IN), .ZN(n4561) );
  AOI22_X1 U5070 ( .A1(n4562), .A2(n4568), .B1(n4561), .B2(n4560), .ZN(U3481)
         );
  AOI22_X1 U5071 ( .A1(n4569), .A2(n4564), .B1(n4563), .B2(n4567), .ZN(U3518)
         );
  AOI22_X1 U5072 ( .A1(n4569), .A2(n4565), .B1(n2332), .B2(n4567), .ZN(U3522)
         );
  AOI22_X1 U5073 ( .A1(n4569), .A2(n4566), .B1(n2398), .B2(n4567), .ZN(U3524)
         );
  AOI22_X1 U5074 ( .A1(n4569), .A2(n4568), .B1(n2410), .B2(n4567), .ZN(U3525)
         );
  AOI22_X1 U5075 ( .A1(STATE_REG_SCAN_IN), .A2(IR_REG_0__SCAN_IN), .B1(
        DATAI_0_), .B2(U3149), .ZN(n4751) );
  AOI22_X1 U5076 ( .A1(n4571), .A2(keyinput_g53), .B1(keyinput_g51), .B2(n2430), .ZN(n4570) );
  OAI221_X1 U5077 ( .B1(n4571), .B2(keyinput_g53), .C1(n2430), .C2(
        keyinput_g51), .A(n4570), .ZN(n4581) );
  AOI22_X1 U5078 ( .A1(n4573), .A2(keyinput_g35), .B1(keyinput_g18), .B2(n4691), .ZN(n4572) );
  OAI221_X1 U5079 ( .B1(n4573), .B2(keyinput_g35), .C1(n4691), .C2(
        keyinput_g18), .A(n4572), .ZN(n4580) );
  XOR2_X1 U5080 ( .A(n4574), .B(keyinput_g1), .Z(n4578) );
  XNOR2_X1 U5081 ( .A(DATAI_0_), .B(keyinput_g31), .ZN(n4577) );
  XNOR2_X1 U5082 ( .A(DATAI_9_), .B(keyinput_g22), .ZN(n4576) );
  XNOR2_X1 U5083 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_g50), .ZN(n4575) );
  NAND4_X1 U5084 ( .A1(n4578), .A2(n4577), .A3(n4576), .A4(n4575), .ZN(n4579)
         );
  NOR3_X1 U5085 ( .A1(n4581), .A2(n4580), .A3(n4579), .ZN(n4615) );
  AOI22_X1 U5086 ( .A1(n2378), .A2(keyinput_g47), .B1(keyinput_g16), .B2(n4672), .ZN(n4582) );
  OAI221_X1 U5087 ( .B1(n2378), .B2(keyinput_g47), .C1(n4672), .C2(
        keyinput_g16), .A(n4582), .ZN(n4590) );
  AOI22_X1 U5088 ( .A1(DATAI_19_), .A2(keyinput_g12), .B1(IR_REG_8__SCAN_IN), 
        .B2(keyinput_g63), .ZN(n4583) );
  OAI221_X1 U5089 ( .B1(DATAI_19_), .B2(keyinput_g12), .C1(IR_REG_8__SCAN_IN), 
        .C2(keyinput_g63), .A(n4583), .ZN(n4589) );
  AOI22_X1 U5090 ( .A1(n4666), .A2(keyinput_g37), .B1(n4665), .B2(keyinput_g39), .ZN(n4584) );
  OAI221_X1 U5091 ( .B1(n4666), .B2(keyinput_g37), .C1(n4665), .C2(
        keyinput_g39), .A(n4584), .ZN(n4588) );
  INV_X1 U5092 ( .A(DATAI_25_), .ZN(n4673) );
  AOI22_X1 U5093 ( .A1(n4586), .A2(keyinput_g34), .B1(keyinput_g6), .B2(n4673), 
        .ZN(n4585) );
  OAI221_X1 U5094 ( .B1(n4586), .B2(keyinput_g34), .C1(n4673), .C2(keyinput_g6), .A(n4585), .ZN(n4587) );
  NOR4_X1 U5095 ( .A1(n4590), .A2(n4589), .A3(n4588), .A4(n4587), .ZN(n4614)
         );
  AOI22_X1 U5096 ( .A1(n2538), .A2(keyinput_g11), .B1(n3665), .B2(keyinput_g43), .ZN(n4591) );
  OAI221_X1 U5097 ( .B1(n2538), .B2(keyinput_g11), .C1(n3665), .C2(
        keyinput_g43), .A(n4591), .ZN(n4599) );
  AOI22_X1 U5098 ( .A1(n4681), .A2(keyinput_g44), .B1(n2326), .B2(keyinput_g54), .ZN(n4592) );
  OAI221_X1 U5099 ( .B1(n4681), .B2(keyinput_g44), .C1(n2326), .C2(
        keyinput_g54), .A(n4592), .ZN(n4598) );
  XNOR2_X1 U5100 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput_g33), .ZN(n4596) );
  XNOR2_X1 U5101 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_g42), .ZN(n4595) );
  XNOR2_X1 U5102 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_g38), .ZN(n4594) );
  XNOR2_X1 U5103 ( .A(keyinput_g27), .B(DATAI_4_), .ZN(n4593) );
  NAND4_X1 U5104 ( .A1(n4596), .A2(n4595), .A3(n4594), .A4(n4593), .ZN(n4597)
         );
  NOR3_X1 U5105 ( .A1(n4599), .A2(n4598), .A3(n4597), .ZN(n4613) );
  AOI22_X1 U5106 ( .A1(n2505), .A2(keyinput_g14), .B1(n4601), .B2(keyinput_g8), 
        .ZN(n4600) );
  OAI221_X1 U5107 ( .B1(n2505), .B2(keyinput_g14), .C1(n4601), .C2(keyinput_g8), .A(n4600), .ZN(n4611) );
  AOI22_X1 U5108 ( .A1(n4603), .A2(keyinput_g45), .B1(keyinput_g19), .B2(n2481), .ZN(n4602) );
  OAI221_X1 U5109 ( .B1(n4603), .B2(keyinput_g45), .C1(n2481), .C2(
        keyinput_g19), .A(n4602), .ZN(n4610) );
  AOI22_X1 U5110 ( .A1(n2619), .A2(keyinput_g2), .B1(n4605), .B2(keyinput_g46), 
        .ZN(n4604) );
  OAI221_X1 U5111 ( .B1(n2619), .B2(keyinput_g2), .C1(n4605), .C2(keyinput_g46), .A(n4604), .ZN(n4609) );
  XNOR2_X1 U5112 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_g61), .ZN(n4607) );
  XNOR2_X1 U5113 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_g56), .ZN(n4606) );
  NAND2_X1 U5114 ( .A1(n4607), .A2(n4606), .ZN(n4608) );
  NOR4_X1 U5115 ( .A1(n4611), .A2(n4610), .A3(n4609), .A4(n4608), .ZN(n4612)
         );
  NAND4_X1 U5116 ( .A1(n4615), .A2(n4614), .A3(n4613), .A4(n4612), .ZN(n4749)
         );
  AOI22_X1 U5117 ( .A1(DATAI_28_), .A2(keyinput_g3), .B1(REG3_REG_24__SCAN_IN), 
        .B2(keyinput_g49), .ZN(n4616) );
  OAI221_X1 U5118 ( .B1(DATAI_28_), .B2(keyinput_g3), .C1(REG3_REG_24__SCAN_IN), .C2(keyinput_g49), .A(n4616), .ZN(n4623) );
  AOI22_X1 U5119 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput_g52), .B1(
        REG3_REG_28__SCAN_IN), .B2(keyinput_g40), .ZN(n4617) );
  OAI221_X1 U5120 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput_g52), .C1(
        REG3_REG_28__SCAN_IN), .C2(keyinput_g40), .A(n4617), .ZN(n4622) );
  AOI22_X1 U5121 ( .A1(REG3_REG_17__SCAN_IN), .A2(keyinput_g48), .B1(
        IR_REG_0__SCAN_IN), .B2(keyinput_g55), .ZN(n4618) );
  OAI221_X1 U5122 ( .B1(REG3_REG_17__SCAN_IN), .B2(keyinput_g48), .C1(
        IR_REG_0__SCAN_IN), .C2(keyinput_g55), .A(n4618), .ZN(n4621) );
  AOI22_X1 U5123 ( .A1(DATAI_21_), .A2(keyinput_g10), .B1(DATAI_22_), .B2(
        keyinput_g9), .ZN(n4619) );
  OAI221_X1 U5124 ( .B1(DATAI_21_), .B2(keyinput_g10), .C1(DATAI_22_), .C2(
        keyinput_g9), .A(n4619), .ZN(n4620) );
  NOR4_X1 U5125 ( .A1(n4623), .A2(n4622), .A3(n4621), .A4(n4620), .ZN(n4652)
         );
  AOI22_X1 U5126 ( .A1(DATAI_3_), .A2(keyinput_g28), .B1(STATE_REG_SCAN_IN), 
        .B2(keyinput_g32), .ZN(n4624) );
  OAI221_X1 U5127 ( .B1(DATAI_3_), .B2(keyinput_g28), .C1(STATE_REG_SCAN_IN), 
        .C2(keyinput_g32), .A(n4624), .ZN(n4632) );
  AOI22_X1 U5128 ( .A1(DATAI_24_), .A2(keyinput_g7), .B1(DATAI_27_), .B2(
        keyinput_g4), .ZN(n4625) );
  OAI221_X1 U5129 ( .B1(DATAI_24_), .B2(keyinput_g7), .C1(DATAI_27_), .C2(
        keyinput_g4), .A(n4625), .ZN(n4631) );
  XNOR2_X1 U5130 ( .A(n4626), .B(keyinput_g58), .ZN(n4629) );
  XNOR2_X1 U5131 ( .A(n4682), .B(keyinput_g36), .ZN(n4628) );
  XNOR2_X1 U5132 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_g60), .ZN(n4627) );
  NAND3_X1 U5133 ( .A1(n4629), .A2(n4628), .A3(n4627), .ZN(n4630) );
  NOR3_X1 U5134 ( .A1(n4632), .A2(n4631), .A3(n4630), .ZN(n4651) );
  AOI22_X1 U5135 ( .A1(DATAI_1_), .A2(keyinput_g30), .B1(DATAI_2_), .B2(
        keyinput_g29), .ZN(n4633) );
  OAI221_X1 U5136 ( .B1(DATAI_1_), .B2(keyinput_g30), .C1(DATAI_2_), .C2(
        keyinput_g29), .A(n4633), .ZN(n4640) );
  AOI22_X1 U5137 ( .A1(REG3_REG_8__SCAN_IN), .A2(keyinput_g41), .B1(
        IR_REG_2__SCAN_IN), .B2(keyinput_g57), .ZN(n4634) );
  OAI221_X1 U5138 ( .B1(REG3_REG_8__SCAN_IN), .B2(keyinput_g41), .C1(
        IR_REG_2__SCAN_IN), .C2(keyinput_g57), .A(n4634), .ZN(n4639) );
  AOI22_X1 U5139 ( .A1(DATAI_31_), .A2(keyinput_g0), .B1(DATAI_26_), .B2(
        keyinput_g5), .ZN(n4635) );
  OAI221_X1 U5140 ( .B1(DATAI_31_), .B2(keyinput_g0), .C1(DATAI_26_), .C2(
        keyinput_g5), .A(n4635), .ZN(n4638) );
  AOI22_X1 U5141 ( .A1(DATAI_8_), .A2(keyinput_g23), .B1(DATAI_14_), .B2(
        keyinput_g17), .ZN(n4636) );
  OAI221_X1 U5142 ( .B1(DATAI_8_), .B2(keyinput_g23), .C1(DATAI_14_), .C2(
        keyinput_g17), .A(n4636), .ZN(n4637) );
  NOR4_X1 U5143 ( .A1(n4640), .A2(n4639), .A3(n4638), .A4(n4637), .ZN(n4650)
         );
  AOI22_X1 U5144 ( .A1(DATAI_6_), .A2(keyinput_g25), .B1(DATAI_7_), .B2(
        keyinput_g24), .ZN(n4641) );
  OAI221_X1 U5145 ( .B1(DATAI_6_), .B2(keyinput_g25), .C1(DATAI_7_), .C2(
        keyinput_g24), .A(n4641), .ZN(n4648) );
  AOI22_X1 U5146 ( .A1(DATAI_18_), .A2(keyinput_g13), .B1(DATAI_16_), .B2(
        keyinput_g15), .ZN(n4642) );
  OAI221_X1 U5147 ( .B1(DATAI_18_), .B2(keyinput_g13), .C1(DATAI_16_), .C2(
        keyinput_g15), .A(n4642), .ZN(n4647) );
  AOI22_X1 U5148 ( .A1(DATAI_11_), .A2(keyinput_g20), .B1(IR_REG_7__SCAN_IN), 
        .B2(keyinput_g62), .ZN(n4643) );
  OAI221_X1 U5149 ( .B1(DATAI_11_), .B2(keyinput_g20), .C1(IR_REG_7__SCAN_IN), 
        .C2(keyinput_g62), .A(n4643), .ZN(n4646) );
  AOI22_X1 U5150 ( .A1(DATAI_5_), .A2(keyinput_g26), .B1(IR_REG_4__SCAN_IN), 
        .B2(keyinput_g59), .ZN(n4644) );
  OAI221_X1 U5151 ( .B1(DATAI_5_), .B2(keyinput_g26), .C1(IR_REG_4__SCAN_IN), 
        .C2(keyinput_g59), .A(n4644), .ZN(n4645) );
  NOR4_X1 U5152 ( .A1(n4648), .A2(n4647), .A3(n4646), .A4(n4645), .ZN(n4649)
         );
  NAND4_X1 U5153 ( .A1(n4652), .A2(n4651), .A3(n4650), .A4(n4649), .ZN(n4748)
         );
  INV_X1 U5154 ( .A(DATAI_19_), .ZN(n4654) );
  AOI22_X1 U5155 ( .A1(n4654), .A2(keyinput_f12), .B1(U3149), .B2(keyinput_f32), .ZN(n4653) );
  OAI221_X1 U5156 ( .B1(n4654), .B2(keyinput_f12), .C1(U3149), .C2(
        keyinput_f32), .A(n4653), .ZN(n4663) );
  XNOR2_X1 U5157 ( .A(n4655), .B(keyinput_f63), .ZN(n4662) );
  XNOR2_X1 U5158 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput_f33), .ZN(n4659) );
  XNOR2_X1 U5159 ( .A(IR_REG_7__SCAN_IN), .B(keyinput_f62), .ZN(n4658) );
  XNOR2_X1 U5160 ( .A(REG3_REG_14__SCAN_IN), .B(keyinput_f35), .ZN(n4657) );
  XNOR2_X1 U5161 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_f42), .ZN(n4656) );
  NAND4_X1 U5162 ( .A1(n4659), .A2(n4658), .A3(n4657), .A4(n4656), .ZN(n4661)
         );
  XNOR2_X1 U5163 ( .A(keyinput_f5), .B(n2592), .ZN(n4660) );
  NOR4_X1 U5164 ( .A1(n4663), .A2(n4662), .A3(n4661), .A4(n4660), .ZN(n4705)
         );
  AOI22_X1 U5165 ( .A1(n4666), .A2(keyinput_f37), .B1(n4665), .B2(keyinput_f39), .ZN(n4664) );
  OAI221_X1 U5166 ( .B1(n4666), .B2(keyinput_f37), .C1(n4665), .C2(
        keyinput_f39), .A(n4664), .ZN(n4677) );
  INV_X1 U5167 ( .A(DATAI_6_), .ZN(n4668) );
  AOI22_X1 U5168 ( .A1(DATAI_20_), .A2(keyinput_f11), .B1(n4668), .B2(
        keyinput_f25), .ZN(n4667) );
  OAI221_X1 U5169 ( .B1(DATAI_20_), .B2(keyinput_f11), .C1(n4668), .C2(
        keyinput_f25), .A(n4667), .ZN(n4676) );
  AOI22_X1 U5170 ( .A1(n4670), .A2(keyinput_f17), .B1(n3665), .B2(keyinput_f43), .ZN(n4669) );
  OAI221_X1 U5171 ( .B1(n4670), .B2(keyinput_f17), .C1(n3665), .C2(
        keyinput_f43), .A(n4669), .ZN(n4675) );
  AOI22_X1 U5172 ( .A1(n4673), .A2(keyinput_f6), .B1(keyinput_f16), .B2(n4672), 
        .ZN(n4671) );
  OAI221_X1 U5173 ( .B1(n4673), .B2(keyinput_f6), .C1(n4672), .C2(keyinput_f16), .A(n4671), .ZN(n4674) );
  NOR4_X1 U5174 ( .A1(n4677), .A2(n4676), .A3(n4675), .A4(n4674), .ZN(n4704)
         );
  AOI22_X1 U5175 ( .A1(n4679), .A2(keyinput_f0), .B1(n2481), .B2(keyinput_f19), 
        .ZN(n4678) );
  OAI221_X1 U5176 ( .B1(n4679), .B2(keyinput_f0), .C1(n2481), .C2(keyinput_f19), .A(n4678), .ZN(n4689) );
  AOI22_X1 U5177 ( .A1(n4682), .A2(keyinput_f36), .B1(keyinput_f44), .B2(n4681), .ZN(n4680) );
  OAI221_X1 U5178 ( .B1(n4682), .B2(keyinput_f36), .C1(n4681), .C2(
        keyinput_f44), .A(n4680), .ZN(n4688) );
  XNOR2_X1 U5179 ( .A(IR_REG_3__SCAN_IN), .B(keyinput_f58), .ZN(n4686) );
  XNOR2_X1 U5180 ( .A(REG3_REG_3__SCAN_IN), .B(keyinput_f38), .ZN(n4685) );
  XNOR2_X1 U5181 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_f57), .ZN(n4684) );
  XNOR2_X1 U5182 ( .A(keyinput_f29), .B(DATAI_2_), .ZN(n4683) );
  NAND4_X1 U5183 ( .A1(n4686), .A2(n4685), .A3(n4684), .A4(n4683), .ZN(n4687)
         );
  NOR3_X1 U5184 ( .A1(n4689), .A2(n4688), .A3(n4687), .ZN(n4703) );
  AOI22_X1 U5185 ( .A1(n4691), .A2(keyinput_f18), .B1(n2619), .B2(keyinput_f2), 
        .ZN(n4690) );
  OAI221_X1 U5186 ( .B1(n4691), .B2(keyinput_f18), .C1(n2619), .C2(keyinput_f2), .A(n4690), .ZN(n4701) );
  INV_X1 U5187 ( .A(DATAI_4_), .ZN(n4694) );
  AOI22_X1 U5188 ( .A1(n4694), .A2(keyinput_f27), .B1(n4693), .B2(keyinput_f61), .ZN(n4692) );
  OAI221_X1 U5189 ( .B1(n4694), .B2(keyinput_f27), .C1(n4693), .C2(
        keyinput_f61), .A(n4692), .ZN(n4700) );
  XOR2_X1 U5190 ( .A(n2505), .B(keyinput_f14), .Z(n4698) );
  XNOR2_X1 U5191 ( .A(keyinput_f23), .B(DATAI_8_), .ZN(n4697) );
  XNOR2_X1 U5192 ( .A(DATAI_1_), .B(keyinput_f30), .ZN(n4696) );
  XNOR2_X1 U5193 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_f56), .ZN(n4695) );
  NAND4_X1 U5194 ( .A1(n4698), .A2(n4697), .A3(n4696), .A4(n4695), .ZN(n4699)
         );
  NOR3_X1 U5195 ( .A1(n4701), .A2(n4700), .A3(n4699), .ZN(n4702) );
  NAND4_X1 U5196 ( .A1(n4705), .A2(n4704), .A3(n4703), .A4(n4702), .ZN(n4742)
         );
  AOI22_X1 U5197 ( .A1(DATAI_22_), .A2(keyinput_f9), .B1(DATAI_28_), .B2(
        keyinput_f3), .ZN(n4706) );
  OAI221_X1 U5198 ( .B1(DATAI_22_), .B2(keyinput_f9), .C1(DATAI_28_), .C2(
        keyinput_f3), .A(n4706), .ZN(n4713) );
  AOI22_X1 U5199 ( .A1(DATAI_30_), .A2(keyinput_f1), .B1(REG3_REG_20__SCAN_IN), 
        .B2(keyinput_f53), .ZN(n4707) );
  OAI221_X1 U5200 ( .B1(DATAI_30_), .B2(keyinput_f1), .C1(REG3_REG_20__SCAN_IN), .C2(keyinput_f53), .A(n4707), .ZN(n4712) );
  AOI22_X1 U5201 ( .A1(DATAI_18_), .A2(keyinput_f13), .B1(REG3_REG_17__SCAN_IN), .B2(keyinput_f48), .ZN(n4708) );
  OAI221_X1 U5202 ( .B1(DATAI_18_), .B2(keyinput_f13), .C1(
        REG3_REG_17__SCAN_IN), .C2(keyinput_f48), .A(n4708), .ZN(n4711) );
  AOI22_X1 U5203 ( .A1(DATAI_21_), .A2(keyinput_f10), .B1(IR_REG_0__SCAN_IN), 
        .B2(keyinput_f55), .ZN(n4709) );
  OAI221_X1 U5204 ( .B1(DATAI_21_), .B2(keyinput_f10), .C1(IR_REG_0__SCAN_IN), 
        .C2(keyinput_f55), .A(n4709), .ZN(n4710) );
  NOR4_X1 U5205 ( .A1(n4713), .A2(n4712), .A3(n4711), .A4(n4710), .ZN(n4740)
         );
  XOR2_X1 U5206 ( .A(REG3_REG_28__SCAN_IN), .B(keyinput_f40), .Z(n4720) );
  AOI22_X1 U5207 ( .A1(DATAI_3_), .A2(keyinput_f28), .B1(REG3_REG_25__SCAN_IN), 
        .B2(keyinput_f45), .ZN(n4714) );
  OAI221_X1 U5208 ( .B1(DATAI_3_), .B2(keyinput_f28), .C1(REG3_REG_25__SCAN_IN), .C2(keyinput_f45), .A(n4714), .ZN(n4719) );
  AOI22_X1 U5209 ( .A1(REG3_REG_0__SCAN_IN), .A2(keyinput_f52), .B1(
        REG3_REG_24__SCAN_IN), .B2(keyinput_f49), .ZN(n4715) );
  OAI221_X1 U5210 ( .B1(REG3_REG_0__SCAN_IN), .B2(keyinput_f52), .C1(
        REG3_REG_24__SCAN_IN), .C2(keyinput_f49), .A(n4715), .ZN(n4718) );
  AOI22_X1 U5211 ( .A1(DATAI_24_), .A2(keyinput_f7), .B1(DATAI_27_), .B2(
        keyinput_f4), .ZN(n4716) );
  OAI221_X1 U5212 ( .B1(DATAI_24_), .B2(keyinput_f7), .C1(DATAI_27_), .C2(
        keyinput_f4), .A(n4716), .ZN(n4717) );
  NOR4_X1 U5213 ( .A1(n4720), .A2(n4719), .A3(n4718), .A4(n4717), .ZN(n4739)
         );
  AOI22_X1 U5214 ( .A1(DATAI_0_), .A2(keyinput_f31), .B1(REG3_REG_16__SCAN_IN), 
        .B2(keyinput_f46), .ZN(n4721) );
  OAI221_X1 U5215 ( .B1(DATAI_0_), .B2(keyinput_f31), .C1(REG3_REG_16__SCAN_IN), .C2(keyinput_f46), .A(n4721), .ZN(n4728) );
  AOI22_X1 U5216 ( .A1(DATAI_11_), .A2(keyinput_f20), .B1(REG3_REG_8__SCAN_IN), 
        .B2(keyinput_f41), .ZN(n4722) );
  OAI221_X1 U5217 ( .B1(DATAI_11_), .B2(keyinput_f20), .C1(REG3_REG_8__SCAN_IN), .C2(keyinput_f41), .A(n4722), .ZN(n4727) );
  AOI22_X1 U5218 ( .A1(REG3_REG_27__SCAN_IN), .A2(keyinput_f34), .B1(
        IR_REG_5__SCAN_IN), .B2(keyinput_f60), .ZN(n4723) );
  OAI221_X1 U5219 ( .B1(REG3_REG_27__SCAN_IN), .B2(keyinput_f34), .C1(
        IR_REG_5__SCAN_IN), .C2(keyinput_f60), .A(n4723), .ZN(n4726) );
  AOI22_X1 U5220 ( .A1(DATAI_23_), .A2(keyinput_f8), .B1(REG3_REG_4__SCAN_IN), 
        .B2(keyinput_f50), .ZN(n4724) );
  OAI221_X1 U5221 ( .B1(DATAI_23_), .B2(keyinput_f8), .C1(REG3_REG_4__SCAN_IN), 
        .C2(keyinput_f50), .A(n4724), .ZN(n4725) );
  NOR4_X1 U5222 ( .A1(n4728), .A2(n4727), .A3(n4726), .A4(n4725), .ZN(n4738)
         );
  AOI22_X1 U5223 ( .A1(DATAI_7_), .A2(keyinput_f24), .B1(IR_REG_4__SCAN_IN), 
        .B2(keyinput_f59), .ZN(n4729) );
  OAI221_X1 U5224 ( .B1(DATAI_7_), .B2(keyinput_f24), .C1(IR_REG_4__SCAN_IN), 
        .C2(keyinput_f59), .A(n4729), .ZN(n4736) );
  AOI22_X1 U5225 ( .A1(DATAI_16_), .A2(keyinput_f15), .B1(REG3_REG_13__SCAN_IN), .B2(keyinput_f54), .ZN(n4730) );
  OAI221_X1 U5226 ( .B1(DATAI_16_), .B2(keyinput_f15), .C1(
        REG3_REG_13__SCAN_IN), .C2(keyinput_f54), .A(n4730), .ZN(n4735) );
  AOI22_X1 U5227 ( .A1(DATAI_9_), .A2(keyinput_f22), .B1(REG3_REG_9__SCAN_IN), 
        .B2(keyinput_f51), .ZN(n4731) );
  OAI221_X1 U5228 ( .B1(DATAI_9_), .B2(keyinput_f22), .C1(REG3_REG_9__SCAN_IN), 
        .C2(keyinput_f51), .A(n4731), .ZN(n4734) );
  AOI22_X1 U5229 ( .A1(DATAI_5_), .A2(keyinput_f26), .B1(REG3_REG_5__SCAN_IN), 
        .B2(keyinput_f47), .ZN(n4732) );
  OAI221_X1 U5230 ( .B1(DATAI_5_), .B2(keyinput_f26), .C1(REG3_REG_5__SCAN_IN), 
        .C2(keyinput_f47), .A(n4732), .ZN(n4733) );
  NOR4_X1 U5231 ( .A1(n4736), .A2(n4735), .A3(n4734), .A4(n4733), .ZN(n4737)
         );
  NAND4_X1 U5232 ( .A1(n4740), .A2(n4739), .A3(n4738), .A4(n4737), .ZN(n4741)
         );
  OAI22_X1 U5233 ( .A1(keyinput_f21), .A2(n4743), .B1(n4742), .B2(n4741), .ZN(
        n4744) );
  OAI21_X1 U5234 ( .B1(n4744), .B2(keyinput_f21), .A(n4743), .ZN(n4746) );
  NAND3_X1 U5235 ( .A1(n4744), .A2(keyinput_g21), .A3(DATAI_10_), .ZN(n4745)
         );
  OAI21_X1 U5236 ( .B1(keyinput_g21), .B2(n4746), .A(n4745), .ZN(n4747) );
  OAI21_X1 U5237 ( .B1(n4749), .B2(n4748), .A(n4747), .ZN(n4750) );
  XOR2_X1 U5238 ( .A(n4751), .B(n4750), .Z(U3352) );
endmodule

