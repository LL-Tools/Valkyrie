

module b22_C_gen_AntiSAT_k_128_10 ( P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, 
        SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, 
        SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, 
        SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, 
        SI_0_, P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN, 
        P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN, 
        P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN, 
        P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN, 
        P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN, 
        P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN, 
        P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN, 
        P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN, 
        P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN, 
        P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN, P3_REG3_REG_0__SCAN_IN, 
        P3_REG3_REG_20__SCAN_IN, P3_REG3_REG_13__SCAN_IN, 
        P3_REG3_REG_22__SCAN_IN, P3_REG3_REG_11__SCAN_IN, 
        P3_REG3_REG_2__SCAN_IN, P3_REG3_REG_18__SCAN_IN, 
        P3_REG3_REG_6__SCAN_IN, P3_REG3_REG_26__SCAN_IN, 
        P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_ADDR_REG_0__SCAN_IN, 
        P3_ADDR_REG_1__SCAN_IN, P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN, 
        P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN, P3_ADDR_REG_6__SCAN_IN, 
        P3_ADDR_REG_7__SCAN_IN, P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, 
        P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, 
        P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, 
        P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, 
        P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, 
        P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, 
        P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, 
        P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, 
        P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, 
        P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, 
        P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, 
        P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, 
        P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, 
        P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, 
        P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, 
        P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, 
        P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, 
        P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, 
        P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, 
        P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, 
        P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, 
        P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, 
        P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN, 
        P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN, 
        P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN, 
        P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN, 
        P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN, 
        P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN, 
        P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN, 
        P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN, 
        P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN, 
        P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN, 
        P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN, 
        P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN, 
        P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN, 
        P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN, 
        P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN, 
        P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN, 
        P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN, 
        P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN, 
        P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN, 
        P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN, 
        P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN, 
        P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN, P2_RD_REG_SCAN_IN, 
        P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN, P3_IR_REG_1__SCAN_IN, 
        P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN, P3_IR_REG_4__SCAN_IN, 
        P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN, P3_IR_REG_7__SCAN_IN, 
        P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN, P3_IR_REG_10__SCAN_IN, 
        P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN, P3_IR_REG_13__SCAN_IN, 
        P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN, P3_IR_REG_16__SCAN_IN, 
        P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN, P3_IR_REG_19__SCAN_IN, 
        P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN, P3_IR_REG_22__SCAN_IN, 
        P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN, P3_IR_REG_25__SCAN_IN, 
        P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN, P3_IR_REG_28__SCAN_IN, 
        P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN, P3_IR_REG_31__SCAN_IN, 
        P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN, P3_D_REG_2__SCAN_IN, 
        P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN, P3_D_REG_5__SCAN_IN, 
        P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN, P3_D_REG_8__SCAN_IN, 
        P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN, P3_D_REG_11__SCAN_IN, 
        P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN, P3_D_REG_14__SCAN_IN, 
        P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN, P3_D_REG_17__SCAN_IN, 
        P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN, P3_D_REG_20__SCAN_IN, 
        P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN, P3_D_REG_23__SCAN_IN, 
        P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN, P3_D_REG_26__SCAN_IN, 
        P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN, P3_D_REG_29__SCAN_IN, 
        P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN, P3_REG0_REG_0__SCAN_IN, 
        P3_REG0_REG_1__SCAN_IN, P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN, 
        P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN, P3_REG0_REG_6__SCAN_IN, 
        P3_REG0_REG_7__SCAN_IN, P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN, 
        P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN, 
        P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN, 
        P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN, 
        P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN, 
        P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN, 
        P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN, 
        P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN, 
        P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN, 
        P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN, 
        P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN, 
        P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN, 
        P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN, P3_REG1_REG_2__SCAN_IN, 
        P3_REG1_REG_3__SCAN_IN, P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN, 
        P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN, P3_REG1_REG_8__SCAN_IN, 
        P3_REG1_REG_9__SCAN_IN, P3_REG1_REG_10__SCAN_IN, 
        P3_REG1_REG_11__SCAN_IN, P3_REG1_REG_12__SCAN_IN, 
        P3_REG1_REG_13__SCAN_IN, P3_REG1_REG_14__SCAN_IN, 
        P3_REG1_REG_15__SCAN_IN, P3_REG1_REG_16__SCAN_IN, 
        P3_REG1_REG_17__SCAN_IN, P3_REG1_REG_18__SCAN_IN, 
        P3_REG1_REG_19__SCAN_IN, P3_REG1_REG_20__SCAN_IN, 
        P3_REG1_REG_21__SCAN_IN, P3_REG1_REG_22__SCAN_IN, 
        P3_REG1_REG_23__SCAN_IN, P3_REG1_REG_24__SCAN_IN, 
        P3_REG1_REG_25__SCAN_IN, P3_REG1_REG_26__SCAN_IN, 
        P3_REG1_REG_27__SCAN_IN, P3_REG1_REG_28__SCAN_IN, 
        P3_REG1_REG_29__SCAN_IN, P3_REG1_REG_30__SCAN_IN, 
        P3_REG1_REG_31__SCAN_IN, P3_REG2_REG_0__SCAN_IN, 
        P3_REG2_REG_1__SCAN_IN, P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN, 
        P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN, P3_REG2_REG_6__SCAN_IN, 
        P3_REG2_REG_7__SCAN_IN, P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN, 
        P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN, 
        P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN, 
        P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN, 
        P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN, 
        P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN, 
        P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN, 
        P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN, 
        P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN, 
        P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN, 
        P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN, 
        P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN, 
        P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN, 
        P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN, 
        P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN, 
        P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN, 
        P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0, 
        keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5, 
        keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10, 
        keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15, 
        keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20, 
        keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25, 
        keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30, 
        keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35, 
        keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40, 
        keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45, 
        keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50, 
        keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55, 
        keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60, 
        keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1, 
        keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6, 
        keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11, 
        keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16, 
        keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21, 
        keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26, 
        keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31, 
        keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36, 
        keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41, 
        keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46, 
        keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51, 
        keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56, 
        keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61, 
        keyinput_g62, keyinput_g63, SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, 
        SUB_1596_U64, SUB_1596_U65, SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, 
        SUB_1596_U69, SUB_1596_U70, SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, 
        SUB_1596_U57, SUB_1596_U58, SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, 
        SUB_1596_U5, SUB_1596_U53, U29, U28, P1_U3355, P1_U3354, P1_U3353, 
        P1_U3352, P1_U3351, P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, 
        P1_U3345, P1_U3344, P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, 
        P1_U3338, P1_U3337, P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, 
        P1_U3331, P1_U3330, P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, 
        P1_U3324, P1_U3445, P1_U3446, P1_U3323, P1_U3322, P1_U3321, P1_U3320, 
        P1_U3319, P1_U3318, P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, 
        P1_U3312, P1_U3311, P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, 
        P1_U3305, P1_U3304, P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, 
        P1_U3298, P1_U3297, P1_U3296, P1_U3295, P1_U3294, P1_U3459, P1_U3462, 
        P1_U3465, P1_U3468, P1_U3471, P1_U3474, P1_U3477, P1_U3480, P1_U3483, 
        P1_U3486, P1_U3489, P1_U3492, P1_U3495, P1_U3498, P1_U3501, P1_U3504, 
        P1_U3507, P1_U3510, P1_U3513, P1_U3515, P1_U3516, P1_U3517, P1_U3518, 
        P1_U3519, P1_U3520, P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, 
        P1_U3526, P1_U3527, P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, 
        P1_U3533, P1_U3534, P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, 
        P1_U3540, P1_U3541, P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, 
        P1_U3547, P1_U3548, P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, 
        P1_U3554, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3293, 
        P1_U3292, P1_U3291, P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, 
        P1_U3285, P1_U3284, P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, 
        P1_U3278, P1_U3277, P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, 
        P1_U3271, P1_U3270, P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, 
        P1_U3356, P1_U3264, P1_U3263, P1_U3262, P1_U3261, P1_U3260, P1_U3259, 
        P1_U3258, P1_U3257, P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, 
        P1_U3251, P1_U3250, P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, 
        P1_U3244, P1_U3243, P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, 
        P1_U3565, P1_U3566, P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, 
        P1_U3572, P1_U3573, P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, 
        P1_U3579, P1_U3580, P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, 
        P1_U3586, P1_U3587, P1_U3588, P1_U3589, P1_U3590, P1_U3591, P1_U3242, 
        P1_U3241, P1_U3240, P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, 
        P1_U3234, P1_U3233, P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, 
        P1_U3227, P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, 
        P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, 
        P1_U3213, P1_U3086, P1_U3085, P1_U4016, P2_U3327, P2_U3326, P2_U3325, 
        P2_U3324, P2_U3323, P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, 
        P2_U3317, P2_U3316, P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, 
        P2_U3310, P2_U3309, P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, 
        P2_U3303, P2_U3302, P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, 
        P2_U3296, P2_U3416, P2_U3417, P2_U3295, P2_U3294, P2_U3293, P2_U3292, 
        P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287, P2_U3286, P2_U3285, 
        P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280, P2_U3279, P2_U3278, 
        P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273, P2_U3272, P2_U3271, 
        P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266, P2_U3430, P2_U3433, 
        P2_U3436, P2_U3439, P2_U3442, P2_U3445, P2_U3448, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3486, P2_U3487, P2_U3488, P2_U3489, 
        P2_U3490, P2_U3491, P2_U3492, P2_U3493, P2_U3494, P2_U3495, P2_U3496, 
        P2_U3497, P2_U3498, P2_U3499, P2_U3500, P2_U3501, P2_U3502, P2_U3503, 
        P2_U3504, P2_U3505, P2_U3506, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3265, 
        P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259, P2_U3258, 
        P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252, P2_U3251, 
        P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3531, P2_U3532, P2_U3533, P2_U3534, P2_U3535, 
        P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540, P2_U3541, P2_U3542, 
        P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547, P2_U3548, P2_U3549, 
        P2_U3550, P2_U3551, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3328, 
        P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3208, P2_U3207, 
        P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, 
        P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, 
        P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, 
        P2_U3185, P2_U3088, P2_U3087, P2_U3947, P3_U3295, P3_U3294, P3_U3293, 
        P3_U3292, P3_U3291, P3_U3290, P3_U3289, P3_U3288, P3_U3287, P3_U3286, 
        P3_U3285, P3_U3284, P3_U3283, P3_U3282, P3_U3281, P3_U3280, P3_U3279, 
        P3_U3278, P3_U3277, P3_U3276, P3_U3275, P3_U3274, P3_U3273, P3_U3272, 
        P3_U3271, P3_U3270, P3_U3269, P3_U3268, P3_U3267, P3_U3266, P3_U3265, 
        P3_U3264, P3_U3376, P3_U3377, P3_U3263, P3_U3262, P3_U3261, P3_U3260, 
        P3_U3259, P3_U3258, P3_U3257, P3_U3256, P3_U3255, P3_U3254, P3_U3253, 
        P3_U3252, P3_U3251, P3_U3250, P3_U3249, P3_U3248, P3_U3247, P3_U3246, 
        P3_U3245, P3_U3244, P3_U3243, P3_U3242, P3_U3241, P3_U3240, P3_U3239, 
        P3_U3238, P3_U3237, P3_U3236, P3_U3235, P3_U3234, P3_U3390, P3_U3393, 
        P3_U3396, P3_U3399, P3_U3402, P3_U3405, P3_U3408, P3_U3411, P3_U3414, 
        P3_U3417, P3_U3420, P3_U3423, P3_U3426, P3_U3429, P3_U3432, P3_U3435, 
        P3_U3438, P3_U3441, P3_U3444, P3_U3446, P3_U3447, P3_U3448, P3_U3449, 
        P3_U3450, P3_U3451, P3_U3452, P3_U3453, P3_U3454, P3_U3455, P3_U3456, 
        P3_U3457, P3_U3458, P3_U3459, P3_U3460, P3_U3461, P3_U3462, P3_U3463, 
        P3_U3464, P3_U3465, P3_U3466, P3_U3467, P3_U3468, P3_U3469, P3_U3470, 
        P3_U3471, P3_U3472, P3_U3473, P3_U3474, P3_U3475, P3_U3476, P3_U3477, 
        P3_U3478, P3_U3479, P3_U3480, P3_U3481, P3_U3482, P3_U3483, P3_U3484, 
        P3_U3485, P3_U3486, P3_U3487, P3_U3488, P3_U3489, P3_U3490, P3_U3233, 
        P3_U3232, P3_U3231, P3_U3230, P3_U3229, P3_U3228, P3_U3227, P3_U3226, 
        P3_U3225, P3_U3224, P3_U3223, P3_U3222, P3_U3221, P3_U3220, P3_U3219, 
        P3_U3218, P3_U3217, P3_U3216, P3_U3215, P3_U3214, P3_U3213, P3_U3212, 
        P3_U3211, P3_U3210, P3_U3209, P3_U3208, P3_U3207, P3_U3206, P3_U3205, 
        P3_U3204, P3_U3203, P3_U3202, P3_U3201, P3_U3200, P3_U3199, P3_U3198, 
        P3_U3197, P3_U3196, P3_U3195, P3_U3194, P3_U3193, P3_U3192, P3_U3191, 
        P3_U3190, P3_U3189, P3_U3188, P3_U3187, P3_U3186, P3_U3185, P3_U3184, 
        P3_U3183, P3_U3182, P3_U3491, P3_U3492, P3_U3493, P3_U3494, P3_U3495, 
        P3_U3496, P3_U3497, P3_U3498, P3_U3499, P3_U3500, P3_U3501, P3_U3502, 
        P3_U3503, P3_U3504, P3_U3505, P3_U3506, P3_U3507, P3_U3508, P3_U3509, 
        P3_U3510, P3_U3511, P3_U3512, P3_U3513, P3_U3514, P3_U3515, P3_U3516, 
        P3_U3517, P3_U3518, P3_U3519, P3_U3520, P3_U3521, P3_U3522, P3_U3296, 
        P3_U3181, P3_U3180, P3_U3179, P3_U3178, P3_U3177, P3_U3176, P3_U3175, 
        P3_U3174, P3_U3173, P3_U3172, P3_U3171, P3_U3170, P3_U3169, P3_U3168, 
        P3_U3167, P3_U3166, P3_U3165, P3_U3164, P3_U3163, P3_U3162, P3_U3161, 
        P3_U3160, P3_U3159, P3_U3158, P3_U3157, P3_U3156, P3_U3155, P3_U3154, 
        P3_U3153, P3_U3151, P3_U3150, P3_U3897 );
  input P3_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_, SI_28_, SI_27_, SI_26_,
         SI_25_, SI_24_, SI_23_, SI_22_, SI_21_, SI_20_, SI_19_, SI_18_,
         SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, SI_12_, SI_11_, SI_10_, SI_9_,
         SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, SI_3_, SI_2_, SI_1_, SI_0_,
         P3_RD_REG_SCAN_IN, P3_STATE_REG_SCAN_IN, P3_REG3_REG_7__SCAN_IN,
         P3_REG3_REG_27__SCAN_IN, P3_REG3_REG_14__SCAN_IN,
         P3_REG3_REG_23__SCAN_IN, P3_REG3_REG_10__SCAN_IN,
         P3_REG3_REG_3__SCAN_IN, P3_REG3_REG_19__SCAN_IN,
         P3_REG3_REG_28__SCAN_IN, P3_REG3_REG_8__SCAN_IN,
         P3_REG3_REG_1__SCAN_IN, P3_REG3_REG_21__SCAN_IN,
         P3_REG3_REG_12__SCAN_IN, P3_REG3_REG_25__SCAN_IN,
         P3_REG3_REG_16__SCAN_IN, P3_REG3_REG_5__SCAN_IN,
         P3_REG3_REG_17__SCAN_IN, P3_REG3_REG_24__SCAN_IN,
         P3_REG3_REG_4__SCAN_IN, P3_REG3_REG_9__SCAN_IN,
         P3_REG3_REG_0__SCAN_IN, P3_REG3_REG_20__SCAN_IN,
         P3_REG3_REG_13__SCAN_IN, P3_REG3_REG_22__SCAN_IN,
         P3_REG3_REG_11__SCAN_IN, P3_REG3_REG_2__SCAN_IN,
         P3_REG3_REG_18__SCAN_IN, P3_REG3_REG_6__SCAN_IN,
         P3_REG3_REG_26__SCAN_IN, P3_REG3_REG_15__SCAN_IN, P3_B_REG_SCAN_IN,
         P3_DATAO_REG_31__SCAN_IN, P3_DATAO_REG_30__SCAN_IN,
         P3_DATAO_REG_29__SCAN_IN, P3_DATAO_REG_28__SCAN_IN,
         P3_DATAO_REG_27__SCAN_IN, P3_DATAO_REG_26__SCAN_IN,
         P3_DATAO_REG_25__SCAN_IN, P3_DATAO_REG_24__SCAN_IN,
         P3_DATAO_REG_23__SCAN_IN, P3_DATAO_REG_22__SCAN_IN,
         P3_DATAO_REG_21__SCAN_IN, P3_DATAO_REG_20__SCAN_IN,
         P3_DATAO_REG_19__SCAN_IN, P3_DATAO_REG_18__SCAN_IN,
         P3_DATAO_REG_17__SCAN_IN, P3_DATAO_REG_16__SCAN_IN,
         P3_DATAO_REG_15__SCAN_IN, P3_DATAO_REG_14__SCAN_IN,
         P3_DATAO_REG_13__SCAN_IN, P3_DATAO_REG_12__SCAN_IN,
         P3_DATAO_REG_11__SCAN_IN, P3_DATAO_REG_10__SCAN_IN,
         P3_DATAO_REG_9__SCAN_IN, P3_DATAO_REG_8__SCAN_IN,
         P3_DATAO_REG_7__SCAN_IN, P3_DATAO_REG_6__SCAN_IN,
         P3_DATAO_REG_5__SCAN_IN, P3_DATAO_REG_4__SCAN_IN,
         P3_DATAO_REG_3__SCAN_IN, P3_DATAO_REG_2__SCAN_IN,
         P3_DATAO_REG_1__SCAN_IN, P3_DATAO_REG_0__SCAN_IN,
         P3_ADDR_REG_0__SCAN_IN, P3_ADDR_REG_1__SCAN_IN,
         P3_ADDR_REG_2__SCAN_IN, P3_ADDR_REG_3__SCAN_IN,
         P3_ADDR_REG_4__SCAN_IN, P3_ADDR_REG_5__SCAN_IN,
         P3_ADDR_REG_6__SCAN_IN, P3_ADDR_REG_7__SCAN_IN,
         P3_ADDR_REG_8__SCAN_IN, P3_ADDR_REG_9__SCAN_IN, P1_IR_REG_0__SCAN_IN,
         P1_IR_REG_1__SCAN_IN, P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN,
         P1_IR_REG_4__SCAN_IN, P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN,
         P1_IR_REG_7__SCAN_IN, P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN,
         P1_IR_REG_10__SCAN_IN, P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN,
         P1_IR_REG_13__SCAN_IN, P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN,
         P1_IR_REG_16__SCAN_IN, P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN,
         P1_IR_REG_19__SCAN_IN, P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN,
         P1_IR_REG_22__SCAN_IN, P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN,
         P1_IR_REG_25__SCAN_IN, P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN,
         P1_IR_REG_28__SCAN_IN, P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN,
         P1_IR_REG_31__SCAN_IN, P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN,
         P1_D_REG_2__SCAN_IN, P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN,
         P1_D_REG_5__SCAN_IN, P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN,
         P1_D_REG_8__SCAN_IN, P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN,
         P1_D_REG_11__SCAN_IN, P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN,
         P1_D_REG_14__SCAN_IN, P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN,
         P1_D_REG_17__SCAN_IN, P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN,
         P1_D_REG_20__SCAN_IN, P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN,
         P1_D_REG_23__SCAN_IN, P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN,
         P1_D_REG_26__SCAN_IN, P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN,
         P1_D_REG_29__SCAN_IN, P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN,
         P1_REG0_REG_0__SCAN_IN, P1_REG0_REG_1__SCAN_IN,
         P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN,
         P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN,
         P1_REG0_REG_6__SCAN_IN, P1_REG0_REG_7__SCAN_IN,
         P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN,
         P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN,
         P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN,
         P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN,
         P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN,
         P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN,
         P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN,
         P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN,
         P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN,
         P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN,
         P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN,
         P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN,
         P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN,
         P1_REG1_REG_2__SCAN_IN, P1_REG1_REG_3__SCAN_IN,
         P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN,
         P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN,
         P1_REG1_REG_8__SCAN_IN, P1_REG1_REG_9__SCAN_IN,
         P1_REG1_REG_10__SCAN_IN, P1_REG1_REG_11__SCAN_IN,
         P1_REG1_REG_12__SCAN_IN, P1_REG1_REG_13__SCAN_IN,
         P1_REG1_REG_14__SCAN_IN, P1_REG1_REG_15__SCAN_IN,
         P1_REG1_REG_16__SCAN_IN, P1_REG1_REG_17__SCAN_IN,
         P1_REG1_REG_18__SCAN_IN, P1_REG1_REG_19__SCAN_IN,
         P1_REG1_REG_20__SCAN_IN, P1_REG1_REG_21__SCAN_IN,
         P1_REG1_REG_22__SCAN_IN, P1_REG1_REG_23__SCAN_IN,
         P1_REG1_REG_24__SCAN_IN, P1_REG1_REG_25__SCAN_IN,
         P1_REG1_REG_26__SCAN_IN, P1_REG1_REG_27__SCAN_IN,
         P1_REG1_REG_28__SCAN_IN, P1_REG1_REG_29__SCAN_IN,
         P1_REG1_REG_30__SCAN_IN, P1_REG1_REG_31__SCAN_IN,
         P1_REG2_REG_0__SCAN_IN, P1_REG2_REG_1__SCAN_IN,
         P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN,
         P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN,
         P1_REG2_REG_6__SCAN_IN, P1_REG2_REG_7__SCAN_IN,
         P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN,
         P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN,
         P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN,
         P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN,
         P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN,
         P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN,
         P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN,
         P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN,
         P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN,
         P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN,
         P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN,
         P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN,
         P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN,
         P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN,
         P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN,
         P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN,
         P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN,
         P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN,
         P1_ADDR_REG_7__SCAN_IN, P1_ADDR_REG_6__SCAN_IN,
         P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN,
         P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN,
         P1_ADDR_REG_1__SCAN_IN, P1_ADDR_REG_0__SCAN_IN,
         P1_DATAO_REG_0__SCAN_IN, P1_DATAO_REG_1__SCAN_IN,
         P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_3__SCAN_IN,
         P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_5__SCAN_IN,
         P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_7__SCAN_IN,
         P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_9__SCAN_IN,
         P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_11__SCAN_IN,
         P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_13__SCAN_IN,
         P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_15__SCAN_IN,
         P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_17__SCAN_IN,
         P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_19__SCAN_IN,
         P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_21__SCAN_IN,
         P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_23__SCAN_IN,
         P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_25__SCAN_IN,
         P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_27__SCAN_IN,
         P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_29__SCAN_IN,
         P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN,
         P1_REG3_REG_15__SCAN_IN, P1_REG3_REG_26__SCAN_IN,
         P1_REG3_REG_6__SCAN_IN, P1_REG3_REG_18__SCAN_IN,
         P1_REG3_REG_2__SCAN_IN, P1_REG3_REG_11__SCAN_IN,
         P1_REG3_REG_22__SCAN_IN, P1_REG3_REG_13__SCAN_IN,
         P1_REG3_REG_20__SCAN_IN, P1_REG3_REG_0__SCAN_IN,
         P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN,
         P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN,
         P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN,
         P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN,
         P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN,
         P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN,
         P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN,
         P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN,
         P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN,
         P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN,
         P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN,
         P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN,
         P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN,
         P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN,
         P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN,
         P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN,
         P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN,
         P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN,
         P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN,
         P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN,
         P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN,
         P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN,
         P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN,
         P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN,
         P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN,
         P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN,
         P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN,
         P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN,
         P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN,
         P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN,
         P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN,
         P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN,
         P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN,
         P2_REG0_REG_3__SCAN_IN, P2_REG0_REG_4__SCAN_IN,
         P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN,
         P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN,
         P2_REG0_REG_9__SCAN_IN, P2_REG0_REG_10__SCAN_IN,
         P2_REG0_REG_11__SCAN_IN, P2_REG0_REG_12__SCAN_IN,
         P2_REG0_REG_13__SCAN_IN, P2_REG0_REG_14__SCAN_IN,
         P2_REG0_REG_15__SCAN_IN, P2_REG0_REG_16__SCAN_IN,
         P2_REG0_REG_17__SCAN_IN, P2_REG0_REG_18__SCAN_IN,
         P2_REG0_REG_19__SCAN_IN, P2_REG0_REG_20__SCAN_IN,
         P2_REG0_REG_21__SCAN_IN, P2_REG0_REG_22__SCAN_IN,
         P2_REG0_REG_23__SCAN_IN, P2_REG0_REG_24__SCAN_IN,
         P2_REG0_REG_25__SCAN_IN, P2_REG0_REG_26__SCAN_IN,
         P2_REG0_REG_27__SCAN_IN, P2_REG0_REG_28__SCAN_IN,
         P2_REG0_REG_29__SCAN_IN, P2_REG0_REG_30__SCAN_IN,
         P2_REG0_REG_31__SCAN_IN, P2_REG1_REG_0__SCAN_IN,
         P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN,
         P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN,
         P2_REG1_REG_5__SCAN_IN, P2_REG1_REG_6__SCAN_IN,
         P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN,
         P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN,
         P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN,
         P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN,
         P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN,
         P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN,
         P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN,
         P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN,
         P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN,
         P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN,
         P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN,
         P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN,
         P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN,
         P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN,
         P2_REG2_REG_3__SCAN_IN, P2_REG2_REG_4__SCAN_IN,
         P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN,
         P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN,
         P2_REG2_REG_9__SCAN_IN, P2_REG2_REG_10__SCAN_IN,
         P2_REG2_REG_11__SCAN_IN, P2_REG2_REG_12__SCAN_IN,
         P2_REG2_REG_13__SCAN_IN, P2_REG2_REG_14__SCAN_IN,
         P2_REG2_REG_15__SCAN_IN, P2_REG2_REG_16__SCAN_IN,
         P2_REG2_REG_17__SCAN_IN, P2_REG2_REG_18__SCAN_IN,
         P2_REG2_REG_19__SCAN_IN, P2_REG2_REG_20__SCAN_IN,
         P2_REG2_REG_21__SCAN_IN, P2_REG2_REG_22__SCAN_IN,
         P2_REG2_REG_23__SCAN_IN, P2_REG2_REG_24__SCAN_IN,
         P2_REG2_REG_25__SCAN_IN, P2_REG2_REG_26__SCAN_IN,
         P2_REG2_REG_27__SCAN_IN, P2_REG2_REG_28__SCAN_IN,
         P2_REG2_REG_29__SCAN_IN, P2_REG2_REG_30__SCAN_IN,
         P2_REG2_REG_31__SCAN_IN, P2_ADDR_REG_19__SCAN_IN,
         P2_ADDR_REG_18__SCAN_IN, P2_ADDR_REG_17__SCAN_IN,
         P2_ADDR_REG_16__SCAN_IN, P2_ADDR_REG_15__SCAN_IN,
         P2_ADDR_REG_14__SCAN_IN, P2_ADDR_REG_13__SCAN_IN,
         P2_ADDR_REG_12__SCAN_IN, P2_ADDR_REG_11__SCAN_IN,
         P2_ADDR_REG_10__SCAN_IN, P2_ADDR_REG_9__SCAN_IN,
         P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN,
         P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN,
         P2_ADDR_REG_4__SCAN_IN, P2_ADDR_REG_3__SCAN_IN,
         P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN,
         P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN,
         P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN,
         P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN,
         P2_DATAO_REG_5__SCAN_IN, P2_DATAO_REG_6__SCAN_IN,
         P2_DATAO_REG_7__SCAN_IN, P2_DATAO_REG_8__SCAN_IN,
         P2_DATAO_REG_9__SCAN_IN, P2_DATAO_REG_10__SCAN_IN,
         P2_DATAO_REG_11__SCAN_IN, P2_DATAO_REG_12__SCAN_IN,
         P2_DATAO_REG_13__SCAN_IN, P2_DATAO_REG_14__SCAN_IN,
         P2_DATAO_REG_15__SCAN_IN, P2_DATAO_REG_16__SCAN_IN,
         P2_DATAO_REG_17__SCAN_IN, P2_DATAO_REG_18__SCAN_IN,
         P2_DATAO_REG_19__SCAN_IN, P2_DATAO_REG_20__SCAN_IN,
         P2_DATAO_REG_21__SCAN_IN, P2_DATAO_REG_22__SCAN_IN,
         P2_DATAO_REG_23__SCAN_IN, P2_DATAO_REG_24__SCAN_IN,
         P2_DATAO_REG_25__SCAN_IN, P2_DATAO_REG_26__SCAN_IN,
         P2_DATAO_REG_27__SCAN_IN, P2_DATAO_REG_28__SCAN_IN,
         P2_DATAO_REG_29__SCAN_IN, P2_DATAO_REG_30__SCAN_IN,
         P2_DATAO_REG_31__SCAN_IN, P2_B_REG_SCAN_IN, P2_REG3_REG_15__SCAN_IN,
         P2_REG3_REG_26__SCAN_IN, P2_REG3_REG_6__SCAN_IN,
         P2_REG3_REG_18__SCAN_IN, P2_REG3_REG_2__SCAN_IN,
         P2_REG3_REG_11__SCAN_IN, P2_REG3_REG_22__SCAN_IN,
         P2_REG3_REG_13__SCAN_IN, P2_REG3_REG_20__SCAN_IN,
         P2_REG3_REG_0__SCAN_IN, P2_REG3_REG_9__SCAN_IN,
         P2_REG3_REG_4__SCAN_IN, P2_REG3_REG_24__SCAN_IN,
         P2_REG3_REG_17__SCAN_IN, P2_REG3_REG_5__SCAN_IN,
         P2_REG3_REG_16__SCAN_IN, P2_REG3_REG_25__SCAN_IN,
         P2_REG3_REG_12__SCAN_IN, P2_REG3_REG_21__SCAN_IN,
         P2_REG3_REG_1__SCAN_IN, P2_REG3_REG_8__SCAN_IN,
         P2_REG3_REG_28__SCAN_IN, P2_REG3_REG_19__SCAN_IN,
         P2_REG3_REG_3__SCAN_IN, P2_REG3_REG_10__SCAN_IN,
         P2_REG3_REG_23__SCAN_IN, P2_REG3_REG_14__SCAN_IN,
         P2_REG3_REG_27__SCAN_IN, P2_REG3_REG_7__SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_RD_REG_SCAN_IN, P2_WR_REG_SCAN_IN, P3_IR_REG_0__SCAN_IN,
         P3_IR_REG_1__SCAN_IN, P3_IR_REG_2__SCAN_IN, P3_IR_REG_3__SCAN_IN,
         P3_IR_REG_4__SCAN_IN, P3_IR_REG_5__SCAN_IN, P3_IR_REG_6__SCAN_IN,
         P3_IR_REG_7__SCAN_IN, P3_IR_REG_8__SCAN_IN, P3_IR_REG_9__SCAN_IN,
         P3_IR_REG_10__SCAN_IN, P3_IR_REG_11__SCAN_IN, P3_IR_REG_12__SCAN_IN,
         P3_IR_REG_13__SCAN_IN, P3_IR_REG_14__SCAN_IN, P3_IR_REG_15__SCAN_IN,
         P3_IR_REG_16__SCAN_IN, P3_IR_REG_17__SCAN_IN, P3_IR_REG_18__SCAN_IN,
         P3_IR_REG_19__SCAN_IN, P3_IR_REG_20__SCAN_IN, P3_IR_REG_21__SCAN_IN,
         P3_IR_REG_22__SCAN_IN, P3_IR_REG_23__SCAN_IN, P3_IR_REG_24__SCAN_IN,
         P3_IR_REG_25__SCAN_IN, P3_IR_REG_26__SCAN_IN, P3_IR_REG_27__SCAN_IN,
         P3_IR_REG_28__SCAN_IN, P3_IR_REG_29__SCAN_IN, P3_IR_REG_30__SCAN_IN,
         P3_IR_REG_31__SCAN_IN, P3_D_REG_0__SCAN_IN, P3_D_REG_1__SCAN_IN,
         P3_D_REG_2__SCAN_IN, P3_D_REG_3__SCAN_IN, P3_D_REG_4__SCAN_IN,
         P3_D_REG_5__SCAN_IN, P3_D_REG_6__SCAN_IN, P3_D_REG_7__SCAN_IN,
         P3_D_REG_8__SCAN_IN, P3_D_REG_9__SCAN_IN, P3_D_REG_10__SCAN_IN,
         P3_D_REG_11__SCAN_IN, P3_D_REG_12__SCAN_IN, P3_D_REG_13__SCAN_IN,
         P3_D_REG_14__SCAN_IN, P3_D_REG_15__SCAN_IN, P3_D_REG_16__SCAN_IN,
         P3_D_REG_17__SCAN_IN, P3_D_REG_18__SCAN_IN, P3_D_REG_19__SCAN_IN,
         P3_D_REG_20__SCAN_IN, P3_D_REG_21__SCAN_IN, P3_D_REG_22__SCAN_IN,
         P3_D_REG_23__SCAN_IN, P3_D_REG_24__SCAN_IN, P3_D_REG_25__SCAN_IN,
         P3_D_REG_26__SCAN_IN, P3_D_REG_27__SCAN_IN, P3_D_REG_28__SCAN_IN,
         P3_D_REG_29__SCAN_IN, P3_D_REG_30__SCAN_IN, P3_D_REG_31__SCAN_IN,
         P3_REG0_REG_0__SCAN_IN, P3_REG0_REG_1__SCAN_IN,
         P3_REG0_REG_2__SCAN_IN, P3_REG0_REG_3__SCAN_IN,
         P3_REG0_REG_4__SCAN_IN, P3_REG0_REG_5__SCAN_IN,
         P3_REG0_REG_6__SCAN_IN, P3_REG0_REG_7__SCAN_IN,
         P3_REG0_REG_8__SCAN_IN, P3_REG0_REG_9__SCAN_IN,
         P3_REG0_REG_10__SCAN_IN, P3_REG0_REG_11__SCAN_IN,
         P3_REG0_REG_12__SCAN_IN, P3_REG0_REG_13__SCAN_IN,
         P3_REG0_REG_14__SCAN_IN, P3_REG0_REG_15__SCAN_IN,
         P3_REG0_REG_16__SCAN_IN, P3_REG0_REG_17__SCAN_IN,
         P3_REG0_REG_18__SCAN_IN, P3_REG0_REG_19__SCAN_IN,
         P3_REG0_REG_20__SCAN_IN, P3_REG0_REG_21__SCAN_IN,
         P3_REG0_REG_22__SCAN_IN, P3_REG0_REG_23__SCAN_IN,
         P3_REG0_REG_24__SCAN_IN, P3_REG0_REG_25__SCAN_IN,
         P3_REG0_REG_26__SCAN_IN, P3_REG0_REG_27__SCAN_IN,
         P3_REG0_REG_28__SCAN_IN, P3_REG0_REG_29__SCAN_IN,
         P3_REG0_REG_30__SCAN_IN, P3_REG0_REG_31__SCAN_IN,
         P3_REG1_REG_0__SCAN_IN, P3_REG1_REG_1__SCAN_IN,
         P3_REG1_REG_2__SCAN_IN, P3_REG1_REG_3__SCAN_IN,
         P3_REG1_REG_4__SCAN_IN, P3_REG1_REG_5__SCAN_IN,
         P3_REG1_REG_6__SCAN_IN, P3_REG1_REG_7__SCAN_IN,
         P3_REG1_REG_8__SCAN_IN, P3_REG1_REG_9__SCAN_IN,
         P3_REG1_REG_10__SCAN_IN, P3_REG1_REG_11__SCAN_IN,
         P3_REG1_REG_12__SCAN_IN, P3_REG1_REG_13__SCAN_IN,
         P3_REG1_REG_14__SCAN_IN, P3_REG1_REG_15__SCAN_IN,
         P3_REG1_REG_16__SCAN_IN, P3_REG1_REG_17__SCAN_IN,
         P3_REG1_REG_18__SCAN_IN, P3_REG1_REG_19__SCAN_IN,
         P3_REG1_REG_20__SCAN_IN, P3_REG1_REG_21__SCAN_IN,
         P3_REG1_REG_22__SCAN_IN, P3_REG1_REG_23__SCAN_IN,
         P3_REG1_REG_24__SCAN_IN, P3_REG1_REG_25__SCAN_IN,
         P3_REG1_REG_26__SCAN_IN, P3_REG1_REG_27__SCAN_IN,
         P3_REG1_REG_28__SCAN_IN, P3_REG1_REG_29__SCAN_IN,
         P3_REG1_REG_30__SCAN_IN, P3_REG1_REG_31__SCAN_IN,
         P3_REG2_REG_0__SCAN_IN, P3_REG2_REG_1__SCAN_IN,
         P3_REG2_REG_2__SCAN_IN, P3_REG2_REG_3__SCAN_IN,
         P3_REG2_REG_4__SCAN_IN, P3_REG2_REG_5__SCAN_IN,
         P3_REG2_REG_6__SCAN_IN, P3_REG2_REG_7__SCAN_IN,
         P3_REG2_REG_8__SCAN_IN, P3_REG2_REG_9__SCAN_IN,
         P3_REG2_REG_10__SCAN_IN, P3_REG2_REG_11__SCAN_IN,
         P3_REG2_REG_12__SCAN_IN, P3_REG2_REG_13__SCAN_IN,
         P3_REG2_REG_14__SCAN_IN, P3_REG2_REG_15__SCAN_IN,
         P3_REG2_REG_16__SCAN_IN, P3_REG2_REG_17__SCAN_IN,
         P3_REG2_REG_18__SCAN_IN, P3_REG2_REG_19__SCAN_IN,
         P3_REG2_REG_20__SCAN_IN, P3_REG2_REG_21__SCAN_IN,
         P3_REG2_REG_22__SCAN_IN, P3_REG2_REG_23__SCAN_IN,
         P3_REG2_REG_24__SCAN_IN, P3_REG2_REG_25__SCAN_IN,
         P3_REG2_REG_26__SCAN_IN, P3_REG2_REG_27__SCAN_IN,
         P3_REG2_REG_28__SCAN_IN, P3_REG2_REG_29__SCAN_IN,
         P3_REG2_REG_30__SCAN_IN, P3_REG2_REG_31__SCAN_IN,
         P3_ADDR_REG_19__SCAN_IN, P3_ADDR_REG_18__SCAN_IN,
         P3_ADDR_REG_17__SCAN_IN, P3_ADDR_REG_16__SCAN_IN,
         P3_ADDR_REG_15__SCAN_IN, P3_ADDR_REG_14__SCAN_IN,
         P3_ADDR_REG_13__SCAN_IN, P3_ADDR_REG_12__SCAN_IN,
         P3_ADDR_REG_11__SCAN_IN, P3_ADDR_REG_10__SCAN_IN, keyinput_f0,
         keyinput_f1, keyinput_f2, keyinput_f3, keyinput_f4, keyinput_f5,
         keyinput_f6, keyinput_f7, keyinput_f8, keyinput_f9, keyinput_f10,
         keyinput_f11, keyinput_f12, keyinput_f13, keyinput_f14, keyinput_f15,
         keyinput_f16, keyinput_f17, keyinput_f18, keyinput_f19, keyinput_f20,
         keyinput_f21, keyinput_f22, keyinput_f23, keyinput_f24, keyinput_f25,
         keyinput_f26, keyinput_f27, keyinput_f28, keyinput_f29, keyinput_f30,
         keyinput_f31, keyinput_f32, keyinput_f33, keyinput_f34, keyinput_f35,
         keyinput_f36, keyinput_f37, keyinput_f38, keyinput_f39, keyinput_f40,
         keyinput_f41, keyinput_f42, keyinput_f43, keyinput_f44, keyinput_f45,
         keyinput_f46, keyinput_f47, keyinput_f48, keyinput_f49, keyinput_f50,
         keyinput_f51, keyinput_f52, keyinput_f53, keyinput_f54, keyinput_f55,
         keyinput_f56, keyinput_f57, keyinput_f58, keyinput_f59, keyinput_f60,
         keyinput_f61, keyinput_f62, keyinput_f63, keyinput_g0, keyinput_g1,
         keyinput_g2, keyinput_g3, keyinput_g4, keyinput_g5, keyinput_g6,
         keyinput_g7, keyinput_g8, keyinput_g9, keyinput_g10, keyinput_g11,
         keyinput_g12, keyinput_g13, keyinput_g14, keyinput_g15, keyinput_g16,
         keyinput_g17, keyinput_g18, keyinput_g19, keyinput_g20, keyinput_g21,
         keyinput_g22, keyinput_g23, keyinput_g24, keyinput_g25, keyinput_g26,
         keyinput_g27, keyinput_g28, keyinput_g29, keyinput_g30, keyinput_g31,
         keyinput_g32, keyinput_g33, keyinput_g34, keyinput_g35, keyinput_g36,
         keyinput_g37, keyinput_g38, keyinput_g39, keyinput_g40, keyinput_g41,
         keyinput_g42, keyinput_g43, keyinput_g44, keyinput_g45, keyinput_g46,
         keyinput_g47, keyinput_g48, keyinput_g49, keyinput_g50, keyinput_g51,
         keyinput_g52, keyinput_g53, keyinput_g54, keyinput_g55, keyinput_g56,
         keyinput_g57, keyinput_g58, keyinput_g59, keyinput_g60, keyinput_g61,
         keyinput_g62, keyinput_g63;
  output SUB_1596_U4, SUB_1596_U62, SUB_1596_U63, SUB_1596_U64, SUB_1596_U65,
         SUB_1596_U66, SUB_1596_U67, SUB_1596_U68, SUB_1596_U69, SUB_1596_U70,
         SUB_1596_U54, SUB_1596_U55, SUB_1596_U56, SUB_1596_U57, SUB_1596_U58,
         SUB_1596_U59, SUB_1596_U60, SUB_1596_U61, SUB_1596_U5, SUB_1596_U53,
         U29, U28, P1_U3355, P1_U3354, P1_U3353, P1_U3352, P1_U3351, P1_U3350,
         P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343,
         P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336,
         P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329,
         P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3445, P1_U3446,
         P1_U3323, P1_U3322, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317,
         P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310,
         P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303,
         P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296,
         P1_U3295, P1_U3294, P1_U3459, P1_U3462, P1_U3465, P1_U3468, P1_U3471,
         P1_U3474, P1_U3477, P1_U3480, P1_U3483, P1_U3486, P1_U3489, P1_U3492,
         P1_U3495, P1_U3498, P1_U3501, P1_U3504, P1_U3507, P1_U3510, P1_U3513,
         P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521,
         P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528,
         P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535,
         P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542,
         P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549,
         P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3555, P1_U3556,
         P1_U3557, P1_U3558, P1_U3559, P1_U3293, P1_U3292, P1_U3291, P1_U3290,
         P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283,
         P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276,
         P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269,
         P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3356, P1_U3264, P1_U3263,
         P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256,
         P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249,
         P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3560,
         P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567,
         P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574,
         P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581,
         P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3587, P1_U3588,
         P1_U3589, P1_U3590, P1_U3591, P1_U3242, P1_U3241, P1_U3240, P1_U3239,
         P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232,
         P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3086, P1_U3085,
         P1_U4016, P2_U3327, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322,
         P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315,
         P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308,
         P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301,
         P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3296, P2_U3416, P2_U3417,
         P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289,
         P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282,
         P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275,
         P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268,
         P2_U3267, P2_U3266, P2_U3430, P2_U3433, P2_U3436, P2_U3439, P2_U3442,
         P2_U3445, P2_U3448, P2_U3451, P2_U3454, P2_U3457, P2_U3460, P2_U3463,
         P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481, P2_U3484,
         P2_U3486, P2_U3487, P2_U3488, P2_U3489, P2_U3490, P2_U3491, P2_U3492,
         P2_U3493, P2_U3494, P2_U3495, P2_U3496, P2_U3497, P2_U3498, P2_U3499,
         P2_U3500, P2_U3501, P2_U3502, P2_U3503, P2_U3504, P2_U3505, P2_U3506,
         P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512, P2_U3513,
         P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519, P2_U3520,
         P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526, P2_U3527,
         P2_U3528, P2_U3529, P2_U3530, P2_U3265, P2_U3264, P2_U3263, P2_U3262,
         P2_U3261, P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255,
         P2_U3254, P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248,
         P2_U3247, P2_U3246, P2_U3245, P2_U3244, P2_U3243, P2_U3242, P2_U3241,
         P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234,
         P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227,
         P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220,
         P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3531,
         P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538,
         P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545,
         P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3552,
         P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558, P2_U3559,
         P2_U3560, P2_U3561, P2_U3562, P2_U3328, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204,
         P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197,
         P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190,
         P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3088, P2_U3087,
         P2_U3947, P3_U3295, P3_U3294, P3_U3293, P3_U3292, P3_U3291, P3_U3290,
         P3_U3289, P3_U3288, P3_U3287, P3_U3286, P3_U3285, P3_U3284, P3_U3283,
         P3_U3282, P3_U3281, P3_U3280, P3_U3279, P3_U3278, P3_U3277, P3_U3276,
         P3_U3275, P3_U3274, P3_U3273, P3_U3272, P3_U3271, P3_U3270, P3_U3269,
         P3_U3268, P3_U3267, P3_U3266, P3_U3265, P3_U3264, P3_U3376, P3_U3377,
         P3_U3263, P3_U3262, P3_U3261, P3_U3260, P3_U3259, P3_U3258, P3_U3257,
         P3_U3256, P3_U3255, P3_U3254, P3_U3253, P3_U3252, P3_U3251, P3_U3250,
         P3_U3249, P3_U3248, P3_U3247, P3_U3246, P3_U3245, P3_U3244, P3_U3243,
         P3_U3242, P3_U3241, P3_U3240, P3_U3239, P3_U3238, P3_U3237, P3_U3236,
         P3_U3235, P3_U3234, P3_U3390, P3_U3393, P3_U3396, P3_U3399, P3_U3402,
         P3_U3405, P3_U3408, P3_U3411, P3_U3414, P3_U3417, P3_U3420, P3_U3423,
         P3_U3426, P3_U3429, P3_U3432, P3_U3435, P3_U3438, P3_U3441, P3_U3444,
         P3_U3446, P3_U3447, P3_U3448, P3_U3449, P3_U3450, P3_U3451, P3_U3452,
         P3_U3453, P3_U3454, P3_U3455, P3_U3456, P3_U3457, P3_U3458, P3_U3459,
         P3_U3460, P3_U3461, P3_U3462, P3_U3463, P3_U3464, P3_U3465, P3_U3466,
         P3_U3467, P3_U3468, P3_U3469, P3_U3470, P3_U3471, P3_U3472, P3_U3473,
         P3_U3474, P3_U3475, P3_U3476, P3_U3477, P3_U3478, P3_U3479, P3_U3480,
         P3_U3481, P3_U3482, P3_U3483, P3_U3484, P3_U3485, P3_U3486, P3_U3487,
         P3_U3488, P3_U3489, P3_U3490, P3_U3233, P3_U3232, P3_U3231, P3_U3230,
         P3_U3229, P3_U3228, P3_U3227, P3_U3226, P3_U3225, P3_U3224, P3_U3223,
         P3_U3222, P3_U3221, P3_U3220, P3_U3219, P3_U3218, P3_U3217, P3_U3216,
         P3_U3215, P3_U3214, P3_U3213, P3_U3212, P3_U3211, P3_U3210, P3_U3209,
         P3_U3208, P3_U3207, P3_U3206, P3_U3205, P3_U3204, P3_U3203, P3_U3202,
         P3_U3201, P3_U3200, P3_U3199, P3_U3198, P3_U3197, P3_U3196, P3_U3195,
         P3_U3194, P3_U3193, P3_U3192, P3_U3191, P3_U3190, P3_U3189, P3_U3188,
         P3_U3187, P3_U3186, P3_U3185, P3_U3184, P3_U3183, P3_U3182, P3_U3491,
         P3_U3492, P3_U3493, P3_U3494, P3_U3495, P3_U3496, P3_U3497, P3_U3498,
         P3_U3499, P3_U3500, P3_U3501, P3_U3502, P3_U3503, P3_U3504, P3_U3505,
         P3_U3506, P3_U3507, P3_U3508, P3_U3509, P3_U3510, P3_U3511, P3_U3512,
         P3_U3513, P3_U3514, P3_U3515, P3_U3516, P3_U3517, P3_U3518, P3_U3519,
         P3_U3520, P3_U3521, P3_U3522, P3_U3296, P3_U3181, P3_U3180, P3_U3179,
         P3_U3178, P3_U3177, P3_U3176, P3_U3175, P3_U3174, P3_U3173, P3_U3172,
         P3_U3171, P3_U3170, P3_U3169, P3_U3168, P3_U3167, P3_U3166, P3_U3165,
         P3_U3164, P3_U3163, P3_U3162, P3_U3161, P3_U3160, P3_U3159, P3_U3158,
         P3_U3157, P3_U3156, P3_U3155, P3_U3154, P3_U3153, P3_U3151, P3_U3150,
         P3_U3897;
  wire   n6468, n6469, n6470, n6471, n6472, n6473, n6475, n6476, n6477, n6478,
         n6479, n6480, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253;

  NAND2_X1 U7216 ( .A1(n6929), .A2(n6926), .ZN(n13211) );
  AND2_X1 U7217 ( .A1(n10290), .A2(n10322), .ZN(n10370) );
  NAND2_X2 U7219 ( .A1(n9961), .A2(n9960), .ZN(n14789) );
  CLKBUF_X2 U7220 ( .A(n7563), .Z(n8055) );
  INV_X1 U7221 ( .A(n13536), .ZN(n13471) );
  BUF_X2 U7222 ( .A(n9115), .Z(n11688) );
  CLKBUF_X1 U7223 ( .A(n9853), .Z(n11516) );
  CLKBUF_X2 U7224 ( .A(n6476), .Z(n11470) );
  INV_X1 U7225 ( .A(n7754), .ZN(n7743) );
  NAND4_X1 U7226 ( .A1(n9618), .A2(n9617), .A3(n9616), .A4(n9615), .ZN(n13665)
         );
  NAND4_X2 U7227 ( .A1(n9568), .A2(n9567), .A3(n9566), .A4(n9565), .ZN(n14525)
         );
  INV_X1 U7228 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n8907) );
  INV_X1 U7229 ( .A(n11215), .ZN(n11554) );
  INV_X1 U7230 ( .A(P2_IR_REG_5__SCAN_IN), .ZN(n8515) );
  NOR2_X1 U7231 ( .A1(n14859), .A2(n14858), .ZN(n14857) );
  NOR2_X1 U7232 ( .A1(n12207), .A2(n12535), .ZN(n12206) );
  XNOR2_X1 U7233 ( .A(n8313), .B(n12247), .ZN(n12243) );
  NAND2_X1 U7234 ( .A1(n7933), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7934) );
  AND2_X1 U7235 ( .A1(n9107), .A2(n14755), .ZN(n14715) );
  OR2_X1 U7236 ( .A1(n8702), .A2(n6975), .ZN(n6974) );
  INV_X4 U7237 ( .A(n6508), .ZN(n11971) );
  AOI22_X1 U7238 ( .A1(n12083), .A2(n12026), .B1(n6907), .B2(n11955), .ZN(
        n11956) );
  OAI21_X1 U7239 ( .B1(n14880), .B2(n6955), .A(n6954), .ZN(n12149) );
  INV_X2 U7240 ( .A(n8899), .ZN(n9142) );
  NAND2_X1 U7241 ( .A1(n8669), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8670) );
  NOR2_X1 U7242 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n6947) );
  INV_X2 U7243 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n13075) );
  NAND2_X1 U7245 ( .A1(n13886), .A2(n13885), .ZN(n13884) );
  AND2_X1 U7246 ( .A1(n7071), .A2(n9569), .ZN(n14555) );
  XNOR2_X1 U7247 ( .A(n14148), .B(n6688), .ZN(n14189) );
  OAI21_X2 U7248 ( .B1(n8899), .B2(n13075), .A(n8898), .ZN(n14743) );
  OAI211_X1 U7249 ( .C1(n10845), .C2(n7011), .A(n10907), .B(n7008), .ZN(n11052) );
  NAND2_X1 U7250 ( .A1(n10768), .A2(n10767), .ZN(n14432) );
  NAND2_X1 U7251 ( .A1(n11319), .A2(n11318), .ZN(n13987) );
  NAND2_X1 U7252 ( .A1(n6977), .A2(n6973), .ZN(n13432) );
  NAND4_X1 U7253 ( .A1(n9637), .A2(n9636), .A3(n9635), .A4(n9634), .ZN(n13664)
         );
  INV_X1 U7254 ( .A(n13893), .ZN(n14531) );
  XNOR2_X1 U7255 ( .A(n8775), .B(n8774), .ZN(n11185) );
  NAND2_X1 U7256 ( .A1(n8728), .A2(n8727), .ZN(n14121) );
  INV_X2 U7258 ( .A(n13538), .ZN(n13485) );
  INV_X1 U7259 ( .A(n6487), .ZN(n11502) );
  XNOR2_X2 U7260 ( .A(n14198), .B(P2_ADDR_REG_7__SCAN_IN), .ZN(n15250) );
  NAND2_X2 U7261 ( .A1(n11908), .A2(n11907), .ZN(n13992) );
  OAI21_X2 U7262 ( .B1(n7474), .B2(n7337), .A(n7335), .ZN(n11908) );
  NOR2_X2 U7263 ( .A1(n14816), .A2(n8294), .ZN(n8295) );
  NAND2_X2 U7264 ( .A1(n6866), .A2(n14197), .ZN(n14198) );
  NAND2_X2 U7265 ( .A1(n8506), .A2(n8505), .ZN(n8520) );
  AND2_X2 U7266 ( .A1(n6941), .A2(n6940), .ZN(n8313) );
  NAND2_X2 U7267 ( .A1(n10677), .A2(n10676), .ZN(n10769) );
  XNOR2_X2 U7268 ( .A(n14141), .B(n14140), .ZN(n14183) );
  NAND2_X2 U7269 ( .A1(n6664), .A2(n6684), .ZN(n14141) );
  NAND2_X2 U7270 ( .A1(n14146), .A2(n14147), .ZN(n14148) );
  NOR2_X2 U7272 ( .A1(n10343), .A2(n15034), .ZN(n10342) );
  XNOR2_X2 U7273 ( .A(n8300), .B(n10341), .ZN(n10343) );
  OR2_X1 U7274 ( .A1(n9666), .A2(n14545), .ZN(n6469) );
  OR2_X1 U7275 ( .A1(n9666), .A2(n14545), .ZN(n14596) );
  XOR2_X2 U7278 ( .A(n14172), .B(P2_ADDR_REG_4__SCAN_IN), .Z(n15245) );
  NOR2_X2 U7279 ( .A1(n8301), .A2(n10342), .ZN(n14859) );
  NAND2_X2 U7280 ( .A1(n13950), .A2(n13949), .ZN(n13948) );
  NAND2_X2 U7281 ( .A1(n14112), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8772) );
  NOR2_X2 U7282 ( .A1(n7517), .A2(n7516), .ZN(n7518) );
  NAND2_X1 U7283 ( .A1(n11185), .A2(n14120), .ZN(n9853) );
  XNOR2_X2 U7284 ( .A(n8670), .B(P2_IR_REG_21__SCAN_IN), .ZN(n8931) );
  XNOR2_X2 U7285 ( .A(n8306), .B(n8266), .ZN(n12163) );
  INV_X1 U7286 ( .A(n8777), .ZN(n14120) );
  NOR2_X2 U7287 ( .A1(n14270), .A2(n14269), .ZN(n14268) );
  AOI21_X2 U7288 ( .B1(n14478), .B2(n14475), .A(n14232), .ZN(n14270) );
  AND2_X1 U7289 ( .A1(n8067), .A2(n8066), .ZN(n8081) );
  NAND2_X1 U7290 ( .A1(n13624), .A2(n13625), .ZN(n13623) );
  AOI21_X1 U7291 ( .B1(n6743), .B2(n14581), .A(n14028), .ZN(n6742) );
  OAI21_X1 U7292 ( .B1(n7947), .B2(n14949), .A(n12020), .ZN(n12291) );
  NAND2_X1 U7293 ( .A1(n11967), .A2(n11966), .ZN(n12109) );
  NAND2_X1 U7294 ( .A1(n11915), .A2(n11914), .ZN(n13921) );
  OAI22_X1 U7295 ( .A1(n12881), .A2(n6746), .B1(n12882), .B2(n6747), .ZN(
        n12889) );
  OAI22_X1 U7296 ( .A1(n7446), .A2(n6515), .B1(n12874), .B2(n12875), .ZN(
        n12881) );
  NAND2_X1 U7298 ( .A1(n10979), .A2(n10978), .ZN(n13648) );
  INV_X1 U7299 ( .A(n13662), .ZN(n10376) );
  NAND2_X1 U7300 ( .A1(n11575), .A2(n14515), .ZN(n14514) );
  INV_X1 U7301 ( .A(n13665), .ZN(n10192) );
  CLKBUF_X2 U7302 ( .A(P2_U3947), .Z(n6471) );
  XNOR2_X1 U7303 ( .A(n12754), .B(n13064), .ZN(n14701) );
  INV_X2 U7304 ( .A(n11228), .ZN(n14561) );
  NAND2_X1 U7305 ( .A1(n11221), .A2(n11222), .ZN(n11219) );
  XNOR2_X1 U7306 ( .A(n14525), .B(n14555), .ZN(n10151) );
  INV_X4 U7307 ( .A(n12772), .ZN(n12959) );
  CLKBUF_X1 U7308 ( .A(n11502), .Z(n6482) );
  INV_X1 U7309 ( .A(n13063), .ZN(n9188) );
  INV_X2 U7310 ( .A(n6477), .ZN(n12772) );
  INV_X2 U7311 ( .A(n9336), .ZN(n11628) );
  INV_X1 U7312 ( .A(n12740), .ZN(n9024) );
  AOI21_X1 U7313 ( .B1(P3_REG1_REG_4__SCAN_IN), .B2(n9185), .A(n9174), .ZN(
        n8291) );
  INV_X2 U7314 ( .A(n9335), .ZN(n11749) );
  BUF_X4 U7315 ( .A(n6520), .Z(n7625) );
  AND2_X2 U7316 ( .A1(n7754), .A2(n11361), .ZN(n7616) );
  INV_X1 U7317 ( .A(n10112), .ZN(n8231) );
  NAND2_X2 U7318 ( .A1(n11190), .A2(n9284), .ZN(n13539) );
  NAND2_X2 U7319 ( .A1(n7945), .A2(n6841), .ZN(n7754) );
  INV_X2 U7320 ( .A(n13806), .ZN(n11204) );
  NAND2_X1 U7321 ( .A1(n8931), .A2(n8952), .ZN(n9327) );
  NAND2_X2 U7322 ( .A1(n8743), .A2(n14121), .ZN(n11364) );
  NOR2_X1 U7323 ( .A1(n15022), .A2(n9219), .ZN(n9218) );
  INV_X4 U7324 ( .A(n11361), .ZN(n11543) );
  OR2_X1 U7325 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n8465) );
  NOR2_X4 U7326 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .ZN(
        n8247) );
  AOI211_X1 U7327 ( .C1(n14519), .C2(n14033), .A(n11925), .B(n11924), .ZN(
        n11926) );
  OR2_X1 U7328 ( .A1(n12993), .A2(n12989), .ZN(n12990) );
  AND2_X1 U7329 ( .A1(n7174), .A2(n7173), .ZN(n11992) );
  AOI21_X1 U7330 ( .B1(n12952), .B2(n12956), .A(n6763), .ZN(n12958) );
  NOR2_X1 U7331 ( .A1(n6627), .A2(n6626), .ZN(n6625) );
  AND2_X1 U7332 ( .A1(n13330), .A2(n13329), .ZN(n6675) );
  AND2_X1 U7333 ( .A1(n14029), .A2(n14392), .ZN(n6627) );
  NAND2_X1 U7334 ( .A1(n13623), .A2(n13491), .ZN(n13492) );
  XNOR2_X1 U7335 ( .A(n6704), .B(n13173), .ZN(n13335) );
  AOI21_X1 U7336 ( .B1(n7075), .B2(n14392), .A(n7072), .ZN(n14035) );
  OR2_X1 U7337 ( .A1(n13880), .A2(n13879), .ZN(n14059) );
  OAI211_X1 U7338 ( .C1(n8202), .C2(n8201), .A(n8227), .B(n6770), .ZN(n7306)
         );
  AND2_X1 U7339 ( .A1(n12287), .A2(n14983), .ZN(n7981) );
  AND2_X1 U7340 ( .A1(n8390), .A2(n8389), .ZN(n8402) );
  OR2_X1 U7341 ( .A1(n12910), .A2(n12909), .ZN(n12915) );
  NAND2_X1 U7342 ( .A1(n7043), .A2(n6492), .ZN(n13844) );
  AND2_X1 U7343 ( .A1(n8388), .A2(n8387), .ZN(n8389) );
  NAND2_X1 U7344 ( .A1(n11920), .A2(n11919), .ZN(n13878) );
  AND2_X1 U7345 ( .A1(n7965), .A2(n8196), .ZN(n7971) );
  OR2_X1 U7346 ( .A1(n13884), .A2(n7052), .ZN(n7043) );
  AOI21_X1 U7347 ( .B1(n6492), .B2(n7052), .A(n7045), .ZN(n7044) );
  AOI21_X1 U7348 ( .B1(n7006), .B2(n13592), .A(n7005), .ZN(n7004) );
  NAND2_X1 U7349 ( .A1(n11964), .A2(n11963), .ZN(n12046) );
  NAND2_X1 U7350 ( .A1(n13921), .A2(n13920), .ZN(n13919) );
  NAND2_X1 U7351 ( .A1(n12334), .A2(n12335), .ZN(n12333) );
  OR2_X1 U7352 ( .A1(n12311), .A2(n12312), .ZN(n12313) );
  OR2_X1 U7353 ( .A1(n12304), .A2(n11968), .ZN(n8196) );
  XNOR2_X1 U7354 ( .A(n11673), .B(n11662), .ZN(n12690) );
  NAND2_X1 U7355 ( .A1(n13943), .A2(n11897), .ZN(n13933) );
  OAI21_X1 U7356 ( .B1(n12362), .B2(n7869), .A(n7868), .ZN(n12351) );
  OR2_X1 U7357 ( .A1(n8283), .A2(n14893), .ZN(n6624) );
  NAND2_X2 U7358 ( .A1(n11620), .A2(n11619), .ZN(n13363) );
  NAND2_X2 U7359 ( .A1(n11389), .A2(n11388), .ZN(n14062) );
  NAND2_X1 U7360 ( .A1(n13289), .A2(n13288), .ZN(n13287) );
  NAND2_X1 U7361 ( .A1(n11661), .A2(n11660), .ZN(n13368) );
  NAND2_X1 U7362 ( .A1(n6967), .A2(n6965), .ZN(n13289) );
  OAI21_X1 U7363 ( .B1(n13306), .B2(n6710), .A(n6708), .ZN(n6713) );
  NAND2_X1 U7364 ( .A1(n14000), .A2(n11894), .ZN(n13976) );
  NAND2_X1 U7365 ( .A1(n7391), .A2(n7390), .ZN(n12371) );
  NAND2_X1 U7366 ( .A1(n12410), .A2(n7180), .ZN(n12395) );
  OR2_X1 U7367 ( .A1(n11096), .A2(n11905), .ZN(n14003) );
  NAND2_X1 U7368 ( .A1(n6864), .A2(n14462), .ZN(n14468) );
  AND2_X1 U7369 ( .A1(n10844), .A2(n10847), .ZN(n10845) );
  AOI21_X1 U7370 ( .B1(n12825), .B2(n7462), .A(n7458), .ZN(n12837) );
  OR2_X1 U7371 ( .A1(n13648), .A2(n13504), .ZN(n11297) );
  NAND2_X1 U7372 ( .A1(n10732), .A2(n10731), .ZN(n12842) );
  AND2_X1 U7373 ( .A1(n7294), .A2(n10539), .ZN(n7513) );
  NAND2_X1 U7374 ( .A1(n10683), .A2(n10682), .ZN(n10763) );
  NAND2_X1 U7375 ( .A1(n7730), .A2(n7729), .ZN(n12481) );
  NAND2_X1 U7376 ( .A1(n10171), .A2(n10170), .ZN(n10417) );
  XNOR2_X1 U7377 ( .A(n9349), .B(n9348), .ZN(n10970) );
  NAND2_X1 U7378 ( .A1(n6848), .A2(n6847), .ZN(n10142) );
  NAND2_X1 U7379 ( .A1(n14925), .A2(n8114), .ZN(n14913) );
  INV_X1 U7380 ( .A(n10077), .ZN(n6848) );
  AND2_X1 U7381 ( .A1(n10635), .A2(n7685), .ZN(n10807) );
  NAND2_X1 U7382 ( .A1(n6850), .A2(n6849), .ZN(n10077) );
  INV_X1 U7383 ( .A(n10052), .ZN(n6850) );
  NAND2_X1 U7384 ( .A1(n14914), .A2(n7388), .ZN(n10635) );
  NAND2_X1 U7385 ( .A1(n14916), .A2(n14915), .ZN(n14914) );
  AOI21_X1 U7386 ( .B1(n6913), .B2(n6498), .A(n6567), .ZN(n6912) );
  AND2_X1 U7387 ( .A1(n10661), .A2(n6914), .ZN(n6913) );
  NAND2_X1 U7388 ( .A1(n9788), .A2(n9787), .ZN(n12801) );
  NAND2_X1 U7389 ( .A1(n6662), .A2(n9404), .ZN(n9769) );
  CLKBUF_X1 U7390 ( .A(n12703), .Z(n14331) );
  NAND2_X1 U7391 ( .A1(n10150), .A2(n9671), .ZN(n9672) );
  AND2_X1 U7392 ( .A1(n10356), .A2(n7639), .ZN(n14930) );
  OAI21_X1 U7393 ( .B1(n10275), .B2(n6631), .A(n7637), .ZN(n10356) );
  NAND2_X1 U7394 ( .A1(n10152), .A2(n10151), .ZN(n10150) );
  NAND2_X1 U7395 ( .A1(n14514), .A2(n9670), .ZN(n10152) );
  INV_X2 U7396 ( .A(n14808), .ZN(n6470) );
  NAND2_X1 U7397 ( .A1(n8645), .A2(n8644), .ZN(n8658) );
  NAND2_X1 U7398 ( .A1(n6875), .A2(n6874), .ZN(n10306) );
  NAND2_X1 U7399 ( .A1(n9193), .A2(n9192), .ZN(n12776) );
  AND2_X1 U7400 ( .A1(n9293), .A2(n9292), .ZN(n9575) );
  AND2_X1 U7401 ( .A1(n7366), .A2(n8096), .ZN(n10120) );
  AND2_X2 U7402 ( .A1(n8421), .A2(n9889), .ZN(n15015) );
  AND2_X1 U7403 ( .A1(n8121), .A2(n8120), .ZN(n14912) );
  AND2_X1 U7404 ( .A1(n8087), .A2(n8100), .ZN(n14950) );
  AND4_X1 U7405 ( .A1(n7675), .A2(n7674), .A3(n7673), .A4(n7672), .ZN(n10521)
         );
  AND4_X1 U7406 ( .A1(n7662), .A2(n7661), .A3(n7660), .A4(n7659), .ZN(n12101)
         );
  AND4_X1 U7407 ( .A1(n7589), .A2(n7588), .A3(n7587), .A4(n7586), .ZN(n9992)
         );
  NAND2_X1 U7408 ( .A1(n6805), .A2(n6806), .ZN(n9552) );
  AND3_X1 U7409 ( .A1(n9603), .A2(n9602), .A3(n9601), .ZN(n11160) );
  XNOR2_X1 U7410 ( .A(n8291), .B(n9398), .ZN(n9386) );
  NAND2_X1 U7411 ( .A1(n9100), .A2(n9099), .ZN(n12759) );
  NAND4_X1 U7412 ( .A1(n9151), .A2(n9150), .A3(n9149), .A4(n9148), .ZN(n13063)
         );
  NAND4_X2 U7413 ( .A1(n9119), .A2(n9118), .A3(n9117), .A4(n9116), .ZN(n13064)
         );
  INV_X2 U7414 ( .A(n9853), .ZN(n11503) );
  BUF_X2 U7415 ( .A(n12976), .Z(n6477) );
  CLKBUF_X1 U7416 ( .A(n11447), .Z(n6486) );
  INV_X2 U7417 ( .A(n13539), .ZN(n9619) );
  NAND2_X1 U7418 ( .A1(n12721), .A2(n12720), .ZN(n12976) );
  OR2_X2 U7419 ( .A1(n13535), .A2(n13881), .ZN(n13538) );
  NAND4_X1 U7420 ( .A1(n8715), .A2(n8714), .A3(n8713), .A4(n8712), .ZN(n9437)
         );
  INV_X2 U7421 ( .A(n13535), .ZN(n13481) );
  NOR2_X2 U7422 ( .A1(n9327), .A2(n13253), .ZN(n12721) );
  NOR2_X1 U7423 ( .A1(n7557), .A2(n12015), .ZN(n6520) );
  NAND2_X2 U7424 ( .A1(n7754), .A2(n11543), .ZN(n8073) );
  XNOR2_X1 U7425 ( .A(n7932), .B(P3_IR_REG_22__SCAN_IN), .ZN(n9978) );
  NAND2_X1 U7426 ( .A1(n9115), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n8894) );
  INV_X4 U7427 ( .A(n11490), .ZN(n11547) );
  NAND2_X2 U7428 ( .A1(n8915), .A2(n8914), .ZN(n13253) );
  XNOR2_X1 U7429 ( .A(n7938), .B(n7937), .ZN(n9758) );
  XNOR2_X1 U7430 ( .A(n7555), .B(n12588), .ZN(n12015) );
  AND2_X2 U7431 ( .A1(n8711), .A2(n8710), .ZN(n9145) );
  OAI21_X2 U7432 ( .B1(n8527), .B2(n8500), .A(n8499), .ZN(n8538) );
  NAND2_X1 U7433 ( .A1(n7554), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7555) );
  NAND2_X1 U7434 ( .A1(n6745), .A2(n8668), .ZN(n12720) );
  AND2_X1 U7435 ( .A1(n8730), .A2(n9252), .ZN(n8483) );
  XNOR2_X1 U7436 ( .A(n14145), .B(n6868), .ZN(n14170) );
  INV_X1 U7437 ( .A(n11190), .ZN(n9940) );
  XNOR2_X1 U7438 ( .A(n8482), .B(P1_IR_REG_25__SCAN_IN), .ZN(n9253) );
  INV_X1 U7439 ( .A(n14127), .ZN(n9252) );
  AND2_X1 U7440 ( .A1(n14545), .A2(n11206), .ZN(n11190) );
  NOR2_X1 U7441 ( .A1(n7930), .A2(P3_IR_REG_19__SCAN_IN), .ZN(n7935) );
  NAND2_X1 U7442 ( .A1(n7014), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8482) );
  NAND2_X1 U7443 ( .A1(n13424), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8701) );
  XNOR2_X1 U7444 ( .A(n8917), .B(n8916), .ZN(n8952) );
  NOR2_X1 U7445 ( .A1(n8286), .A2(n9218), .ZN(n9046) );
  INV_X1 U7446 ( .A(n8703), .ZN(n8704) );
  XNOR2_X1 U7447 ( .A(n8722), .B(P1_IR_REG_21__SCAN_IN), .ZN(n14545) );
  XNOR2_X1 U7448 ( .A(n8719), .B(P1_IR_REG_22__SCAN_IN), .ZN(n14544) );
  NAND2_X1 U7449 ( .A1(n7536), .A2(n6550), .ZN(n7549) );
  MUX2_X1 U7450 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8726), .S(
        P1_IR_REG_27__SCAN_IN), .Z(n8728) );
  INV_X1 U7451 ( .A(n8718), .ZN(n8470) );
  NAND2_X1 U7452 ( .A1(n8718), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8719) );
  AND2_X1 U7453 ( .A1(n8516), .A2(n8515), .ZN(n8886) );
  NAND2_X1 U7454 ( .A1(n8491), .A2(SI_1_), .ZN(n8497) );
  NAND2_X2 U7455 ( .A1(n11543), .A2(P1_U3086), .ZN(n14124) );
  NAND2_X1 U7456 ( .A1(n8720), .A2(n8469), .ZN(n8718) );
  NOR2_X1 U7457 ( .A1(n8523), .A2(P2_IR_REG_4__SCAN_IN), .ZN(n8516) );
  AND4_X1 U7458 ( .A1(n6766), .A2(n7479), .A3(n6901), .A4(n7395), .ZN(n6765)
         );
  XNOR2_X1 U7459 ( .A(n7607), .B(n7609), .ZN(n9185) );
  NAND2_X1 U7460 ( .A1(n6982), .A2(n6981), .ZN(n9058) );
  INV_X2 U7461 ( .A(n8495), .ZN(n11361) );
  NOR2_X1 U7462 ( .A1(n7396), .A2(P3_IR_REG_26__SCAN_IN), .ZN(n7395) );
  AND3_X1 U7463 ( .A1(n8435), .A2(n8434), .A3(n8433), .ZN(n8885) );
  AND2_X1 U7464 ( .A1(n7483), .A2(P2_DATAO_REG_0__SCAN_IN), .ZN(n7578) );
  AND2_X1 U7465 ( .A1(n7524), .A2(n7680), .ZN(n6900) );
  AND2_X1 U7466 ( .A1(n6676), .A2(P3_ADDR_REG_0__SCAN_IN), .ZN(n14176) );
  INV_X1 U7467 ( .A(P2_IR_REG_30__SCAN_IN), .ZN(n8700) );
  NOR2_X1 U7468 ( .A1(P1_IR_REG_10__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n8781) );
  INV_X1 U7469 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n8784) );
  XNOR2_X1 U7470 ( .A(P3_ADDR_REG_1__SCAN_IN), .B(P1_ADDR_REG_1__SCAN_IN), 
        .ZN(n14175) );
  INV_X4 U7471 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3086) );
  NOR2_X1 U7472 ( .A1(P1_IR_REG_14__SCAN_IN), .A2(P1_IR_REG_8__SCAN_IN), .ZN(
        n8460) );
  NOR2_X1 U7473 ( .A1(P3_IR_REG_15__SCAN_IN), .A2(P3_IR_REG_13__SCAN_IN), .ZN(
        n7527) );
  NOR2_X1 U7474 ( .A1(P3_IR_REG_14__SCAN_IN), .A2(P3_IR_REG_10__SCAN_IN), .ZN(
        n7528) );
  INV_X1 U7475 ( .A(P1_IR_REG_13__SCAN_IN), .ZN(n8970) );
  XNOR2_X1 U7476 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .ZN(n7568) );
  INV_X4 U7477 ( .A(P3_STATE_REG_SCAN_IN), .ZN(P3_U3151) );
  INV_X1 U7478 ( .A(P3_IR_REG_6__SCAN_IN), .ZN(n7650) );
  INV_X1 U7479 ( .A(P3_IR_REG_5__SCAN_IN), .ZN(n7648) );
  NOR2_X1 U7480 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_3__SCAN_IN), .ZN(
        n7524) );
  INV_X1 U7481 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n8511) );
  NOR2_X1 U7482 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n11195) );
  INV_X4 U7483 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3088) );
  NAND2_X1 U7484 ( .A1(n7326), .A2(n7327), .ZN(n6472) );
  NAND2_X1 U7485 ( .A1(n7326), .A2(n7327), .ZN(n13843) );
  OR2_X1 U7486 ( .A1(n14257), .A2(P2_ADDR_REG_10__SCAN_IN), .ZN(n6873) );
  NAND2_X1 U7487 ( .A1(n7348), .A2(n7347), .ZN(n7346) );
  INV_X1 U7488 ( .A(n9593), .ZN(n6473) );
  AOI21_X2 U7489 ( .B1(n10417), .B2(n10416), .A(n10415), .ZN(n10426) );
  NOR2_X1 U7490 ( .A1(n12260), .A2(n6666), .ZN(n8315) );
  CLKBUF_X1 U7491 ( .A(n9594), .Z(n6475) );
  BUF_X2 U7492 ( .A(n9594), .Z(n6476) );
  NAND2_X1 U7493 ( .A1(n8777), .A2(n8776), .ZN(n9594) );
  NAND2_X1 U7494 ( .A1(n7341), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8775) );
  OAI22_X2 U7495 ( .A1(n13201), .A2(n13200), .B1(n13345), .B2(n13042), .ZN(
        n13187) );
  CLKBUF_X1 U7496 ( .A(n9669), .Z(n6478) );
  CLKBUF_X1 U7497 ( .A(n9669), .Z(n6479) );
  CLKBUF_X2 U7498 ( .A(n9669), .Z(n6480) );
  NAND3_X1 U7499 ( .A1(n6670), .A2(n6500), .A3(n9304), .ZN(n9669) );
  OAI222_X1 U7500 ( .A1(n14120), .A2(P1_U3086), .B1(n14119), .B2(n14118), .C1(
        n14117), .C2(n14124), .ZN(P1_U3325) );
  AOI21_X1 U7501 ( .B1(n7970), .B2(n6775), .A(n8205), .ZN(n6774) );
  MUX2_X1 U7503 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n14097), .S(n14613), .Z(
        P1_U3525) );
  OAI21_X1 U7504 ( .B1(n14030), .B2(n14541), .A(n6625), .ZN(n14097) );
  AOI21_X2 U7505 ( .B1(n13959), .B2(n13962), .A(n6518), .ZN(n13950) );
  AND4_X1 U7506 ( .A1(n7311), .A2(n7025), .A3(n8581), .A4(n9269), .ZN(n8720)
         );
  OR2_X1 U7507 ( .A1(n9593), .A2(n14617), .ZN(n9615) );
  BUF_X4 U7508 ( .A(n9030), .Z(n11123) );
  OAI21_X2 U7509 ( .B1(n13499), .B2(n7018), .A(n7016), .ZN(n13569) );
  NAND2_X2 U7510 ( .A1(n13500), .A2(n13501), .ZN(n13499) );
  NAND2_X2 U7511 ( .A1(n11209), .A2(n11213), .ZN(n11575) );
  NAND2_X2 U7512 ( .A1(n6669), .A2(n9667), .ZN(n11209) );
  OAI211_X2 U7513 ( .C1(n9846), .C2(n9624), .A(n9623), .B(n9622), .ZN(n11228)
         );
  NOR2_X1 U7514 ( .A1(n6486), .A2(n9305), .ZN(n9306) );
  XNOR2_X2 U7515 ( .A(n6667), .B(n11998), .ZN(n14030) );
  XNOR2_X2 U7516 ( .A(n8304), .B(n8346), .ZN(n14880) );
  NOR2_X2 U7517 ( .A1(n14857), .A2(n8303), .ZN(n8304) );
  AND2_X1 U7518 ( .A1(n8711), .A2(n8710), .ZN(n6484) );
  AND2_X1 U7519 ( .A1(n8711), .A2(n8710), .ZN(n6485) );
  NAND2_X2 U7520 ( .A1(n8543), .A2(n8464), .ZN(n8587) );
  NOR2_X4 U7521 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n8543) );
  NAND2_X1 U7522 ( .A1(n11185), .A2(n8777), .ZN(n11447) );
  OAI21_X2 U7523 ( .B1(n13992), .B2(n11910), .A(n11909), .ZN(n13974) );
  AND2_X1 U7525 ( .A1(n7754), .A2(n11361), .ZN(n6488) );
  AND3_X1 U7526 ( .A1(n13975), .A2(n11574), .A3(n7119), .ZN(n6490) );
  NAND2_X1 U7527 ( .A1(n7123), .A2(n7120), .ZN(n7119) );
  AND2_X1 U7528 ( .A1(n7106), .A2(n7103), .ZN(n7102) );
  NAND2_X1 U7529 ( .A1(n7107), .A2(n7105), .ZN(n7103) );
  AND2_X1 U7530 ( .A1(n14391), .A2(n11284), .ZN(n7106) );
  AOI21_X1 U7531 ( .B1(n6490), .B2(n7121), .A(n6568), .ZN(n7118) );
  NOR2_X1 U7532 ( .A1(n7123), .A2(n7122), .ZN(n7121) );
  INV_X1 U7533 ( .A(n11909), .ZN(n7122) );
  OAI21_X1 U7534 ( .B1(n7409), .B2(n6727), .A(n7419), .ZN(n6726) );
  NAND2_X1 U7535 ( .A1(P3_ADDR_REG_2__SCAN_IN), .A2(n6685), .ZN(n6684) );
  INV_X1 U7536 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6685) );
  AND2_X1 U7537 ( .A1(n6900), .A2(n6768), .ZN(n6767) );
  INV_X1 U7538 ( .A(n7034), .ZN(n10225) );
  NAND2_X1 U7539 ( .A1(n7039), .A2(n10373), .ZN(n7035) );
  AND3_X2 U7540 ( .A1(n7311), .A2(n8581), .A3(n8468), .ZN(n8477) );
  INV_X1 U7541 ( .A(n6513), .ZN(n8058) );
  OR2_X1 U7542 ( .A1(n12088), .A2(n11941), .ZN(n8160) );
  NOR2_X1 U7543 ( .A1(n11551), .A2(n11213), .ZN(n7080) );
  INV_X1 U7544 ( .A(n11297), .ZN(n7097) );
  INV_X1 U7545 ( .A(n7102), .ZN(n7098) );
  INV_X1 U7546 ( .A(n6514), .ZN(n7093) );
  AOI21_X1 U7547 ( .B1(n6795), .B2(n8123), .A(n6793), .ZN(n6792) );
  NAND2_X1 U7548 ( .A1(n8127), .A2(n8213), .ZN(n6793) );
  AOI21_X1 U7549 ( .B1(n7132), .B2(n7131), .A(n7130), .ZN(n7129) );
  AOI21_X1 U7550 ( .B1(n6789), .B2(n6791), .A(n14898), .ZN(n6788) );
  INV_X1 U7551 ( .A(n6792), .ZN(n6791) );
  AOI21_X1 U7552 ( .B1(n7118), .B2(n7116), .A(n7115), .ZN(n7114) );
  INV_X1 U7553 ( .A(n11341), .ZN(n7115) );
  NOR2_X1 U7554 ( .A1(n11342), .A2(n6490), .ZN(n7116) );
  NAND2_X1 U7555 ( .A1(n12870), .A2(n7447), .ZN(n7446) );
  NAND2_X1 U7556 ( .A1(n12874), .A2(n12875), .ZN(n7447) );
  OAI22_X1 U7557 ( .A1(n8165), .A2(n12416), .B1(n8167), .B2(n8164), .ZN(n6804)
         );
  AND2_X1 U7558 ( .A1(n12355), .A2(n12026), .ZN(n8181) );
  NAND2_X1 U7559 ( .A1(n6715), .A2(n6716), .ZN(n10534) );
  AOI21_X1 U7560 ( .B1(n6504), .B2(n6717), .A(n6600), .ZN(n6716) );
  AND2_X1 U7561 ( .A1(n8467), .A2(n8466), .ZN(n8468) );
  NOR2_X1 U7562 ( .A1(P1_IR_REG_16__SCAN_IN), .A2(P1_IR_REG_15__SCAN_IN), .ZN(
        n8467) );
  NOR2_X1 U7563 ( .A1(P1_IR_REG_18__SCAN_IN), .A2(P1_IR_REG_17__SCAN_IN), .ZN(
        n8466) );
  INV_X1 U7564 ( .A(n6726), .ZN(n6724) );
  INV_X1 U7565 ( .A(n8532), .ZN(n6650) );
  NAND2_X1 U7566 ( .A1(n14143), .A2(n14144), .ZN(n14145) );
  INV_X1 U7567 ( .A(n11970), .ZN(n6898) );
  NAND2_X1 U7568 ( .A1(n7306), .A2(n8203), .ZN(n7302) );
  AND2_X1 U7569 ( .A1(n8620), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n8294) );
  OR2_X1 U7570 ( .A1(n12317), .A2(n12071), .ZN(n8193) );
  NOR2_X1 U7571 ( .A1(n7847), .A2(n7393), .ZN(n7392) );
  INV_X1 U7572 ( .A(n7831), .ZN(n7393) );
  AOI21_X1 U7573 ( .B1(n7161), .B2(n7163), .A(n7159), .ZN(n7158) );
  NAND2_X1 U7574 ( .A1(n14913), .A2(n7161), .ZN(n7160) );
  INV_X1 U7575 ( .A(n8125), .ZN(n7159) );
  INV_X1 U7576 ( .A(n7500), .ZN(n6781) );
  NAND2_X1 U7577 ( .A1(n7216), .A2(n7215), .ZN(n7214) );
  INV_X1 U7578 ( .A(n9416), .ZN(n6696) );
  AND2_X1 U7579 ( .A1(n11574), .A2(n11895), .ZN(n7057) );
  NAND2_X1 U7580 ( .A1(n6888), .A2(n14426), .ZN(n10999) );
  OAI21_X1 U7581 ( .B1(n13933), .B2(n7061), .A(n7059), .ZN(n7069) );
  INV_X1 U7582 ( .A(n7062), .ZN(n7061) );
  AOI21_X1 U7583 ( .B1(n7062), .B2(n7060), .A(n6558), .ZN(n7059) );
  NAND2_X1 U7584 ( .A1(n11430), .A2(n11175), .ZN(n11457) );
  NOR2_X1 U7585 ( .A1(n8475), .A2(n8474), .ZN(n8476) );
  OR2_X1 U7586 ( .A1(n11421), .A2(n11420), .ZN(n11171) );
  NAND2_X1 U7587 ( .A1(n11167), .A2(n11166), .ZN(n11421) );
  AOI21_X1 U7588 ( .B1(n6736), .B2(n6738), .A(n6735), .ZN(n6734) );
  INV_X1 U7589 ( .A(n11073), .ZN(n6735) );
  INV_X1 U7590 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n8461) );
  INV_X1 U7591 ( .A(n8766), .ZN(n7416) );
  AND2_X1 U7592 ( .A1(n12018), .A2(n6897), .ZN(n6896) );
  OR2_X1 U7593 ( .A1(n12110), .A2(n6898), .ZN(n6897) );
  INV_X1 U7594 ( .A(n10668), .ZN(n6914) );
  NOR2_X1 U7595 ( .A1(n7908), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n7917) );
  AND2_X1 U7596 ( .A1(n9758), .A2(n9360), .ZN(n9547) );
  OR2_X1 U7597 ( .A1(n12586), .A2(n9496), .ZN(n9509) );
  AND4_X1 U7598 ( .A1(n7830), .A2(n7829), .A3(n7828), .A4(n7827), .ZN(n11941)
         );
  INV_X1 U7599 ( .A(n9226), .ZN(n8328) );
  OR2_X1 U7600 ( .A1(n9392), .A2(n7350), .ZN(n7349) );
  OR2_X1 U7601 ( .A1(n14819), .A2(n9393), .ZN(n7350) );
  NAND2_X1 U7602 ( .A1(n8254), .A2(n7352), .ZN(n7351) );
  INV_X1 U7603 ( .A(n14819), .ZN(n7352) );
  AOI21_X1 U7604 ( .B1(P3_REG2_REG_16__SCAN_IN), .B2(n12222), .A(n12214), .ZN(
        n8273) );
  NOR2_X1 U7605 ( .A1(n7903), .A2(n7385), .ZN(n7383) );
  OAI22_X1 U7606 ( .A1(n7903), .A2(n7382), .B1(n12330), .B2(n12121), .ZN(n7381) );
  NOR2_X1 U7607 ( .A1(n6594), .A2(n7369), .ZN(n7368) );
  INV_X1 U7608 ( .A(n7789), .ZN(n7369) );
  NAND2_X1 U7609 ( .A1(n7150), .A2(n7148), .ZN(n12442) );
  AOI21_X1 U7610 ( .B1(n7151), .B2(n7153), .A(n7149), .ZN(n7148) );
  INV_X1 U7611 ( .A(n14949), .ZN(n14961) );
  INV_X1 U7612 ( .A(n8073), .ZN(n8047) );
  NAND2_X1 U7613 ( .A1(n7824), .A2(n7823), .ZN(n12088) );
  OAI21_X1 U7614 ( .B1(n7914), .B2(n6825), .A(n6822), .ZN(n8045) );
  INV_X1 U7615 ( .A(n6826), .ZN(n6825) );
  AND2_X1 U7616 ( .A1(n6823), .A2(n6828), .ZN(n6822) );
  AOI21_X1 U7617 ( .B1(n6830), .B2(n8028), .A(n6829), .ZN(n6828) );
  NAND2_X1 U7618 ( .A1(n7553), .A2(n7554), .ZN(n7557) );
  MUX2_X1 U7619 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7550), .S(
        P3_IR_REG_29__SCAN_IN), .Z(n7553) );
  OAI21_X1 U7620 ( .B1(n7914), .B2(n7521), .A(n6833), .ZN(n8027) );
  INV_X1 U7621 ( .A(n7396), .ZN(n7394) );
  NAND2_X1 U7622 ( .A1(P1_DATAO_REG_14__SCAN_IN), .A2(n7299), .ZN(n7298) );
  INV_X1 U7623 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n7299) );
  NAND2_X1 U7624 ( .A1(n7740), .A2(n7738), .ZN(n7505) );
  OAI22_X1 U7625 ( .A1(n12637), .A2(n12636), .B1(n11658), .B2(n11657), .ZN(
        n11673) );
  NAND2_X1 U7626 ( .A1(n11721), .A2(n11720), .ZN(n12922) );
  AND2_X1 U7627 ( .A1(n12708), .A2(n6521), .ZN(n7266) );
  AOI21_X1 U7628 ( .B1(n7216), .B2(n7213), .A(n7212), .ZN(n7211) );
  NOR2_X1 U7629 ( .A1(n11886), .A2(n11884), .ZN(n7212) );
  NOR2_X1 U7630 ( .A1(n13173), .A2(n6523), .ZN(n7213) );
  NAND2_X1 U7631 ( .A1(n7202), .A2(n6526), .ZN(n13230) );
  XNOR2_X1 U7632 ( .A(n13358), .B(n12623), .ZN(n13231) );
  NAND2_X1 U7633 ( .A1(n11855), .A2(n11854), .ZN(n13247) );
  OR2_X1 U7634 ( .A1(n13363), .A2(n12691), .ZN(n11854) );
  NAND2_X1 U7635 ( .A1(n13368), .A2(n13046), .ZN(n7203) );
  AOI21_X1 U7636 ( .B1(n13273), .B2(n11878), .A(n6557), .ZN(n13269) );
  NAND2_X1 U7637 ( .A1(n13269), .A2(n13268), .ZN(n13267) );
  OR2_X1 U7638 ( .A1(n12830), .A2(n13055), .ZN(n7197) );
  NAND2_X1 U7640 ( .A1(n6953), .A2(n9774), .ZN(n9775) );
  NOR2_X1 U7641 ( .A1(n8931), .A2(n13026), .ZN(n8927) );
  NOR2_X1 U7642 ( .A1(n8937), .A2(n13435), .ZN(n14732) );
  NAND2_X1 U7643 ( .A1(n8441), .A2(n7480), .ZN(n8673) );
  NAND2_X1 U7644 ( .A1(n8449), .A2(n8443), .ZN(n8452) );
  AOI22_X1 U7645 ( .A1(n13485), .A2(n6480), .B1(n9619), .B2(n9667), .ZN(n9584)
         );
  INV_X1 U7646 ( .A(n7019), .ZN(n7017) );
  AOI22_X1 U7647 ( .A1(n13481), .A2(n9668), .B1(n9285), .B2(
        P1_REG1_REG_0__SCAN_IN), .ZN(n9293) );
  AND2_X1 U7648 ( .A1(n7125), .A2(n7124), .ZN(n11610) );
  NAND2_X1 U7649 ( .A1(n6503), .A2(n11537), .ZN(n7124) );
  NAND2_X1 U7650 ( .A1(n11550), .A2(n11549), .ZN(n13812) );
  NAND2_X1 U7651 ( .A1(n13847), .A2(n14527), .ZN(n7073) );
  NAND2_X1 U7652 ( .A1(n13828), .A2(n11902), .ZN(n11997) );
  NAND2_X1 U7653 ( .A1(n13905), .A2(n6877), .ZN(n13833) );
  NOR2_X1 U7654 ( .A1(n14038), .A2(n6879), .ZN(n6877) );
  XNOR2_X1 U7655 ( .A(n14049), .B(n13630), .ZN(n13860) );
  OAI21_X1 U7656 ( .B1(n10470), .B2(n7055), .A(n7053), .ZN(n10683) );
  INV_X1 U7657 ( .A(n7054), .ZN(n7053) );
  INV_X1 U7658 ( .A(n10222), .ZN(n7040) );
  NAND2_X1 U7659 ( .A1(n6887), .A2(n14555), .ZN(n10160) );
  INV_X1 U7660 ( .A(n14517), .ZN(n6887) );
  INV_X1 U7661 ( .A(n14024), .ZN(n6743) );
  OAI21_X1 U7662 ( .B1(P1_ADDR_REG_12__SCAN_IN), .B2(n14166), .A(n14165), .ZN(
        n14218) );
  OAI21_X1 U7663 ( .B1(n11012), .B2(n11006), .A(n11011), .ZN(n11013) );
  AOI21_X1 U7664 ( .B1(n11684), .B2(n11683), .A(n11682), .ZN(n12672) );
  NAND2_X1 U7665 ( .A1(n7210), .A2(n7216), .ZN(n6704) );
  NAND2_X1 U7666 ( .A1(n11479), .A2(n11478), .ZN(n14032) );
  INV_X1 U7667 ( .A(n13650), .ZN(n13626) );
  INV_X1 U7668 ( .A(n11241), .ZN(n11244) );
  AOI21_X1 U7669 ( .B1(n12802), .B2(n12803), .A(n6517), .ZN(n7449) );
  NAND2_X1 U7670 ( .A1(n7452), .A2(n7451), .ZN(n7450) );
  INV_X1 U7671 ( .A(n12803), .ZN(n7451) );
  INV_X1 U7672 ( .A(n12802), .ZN(n7452) );
  INV_X1 U7673 ( .A(n11287), .ZN(n7105) );
  NAND2_X1 U7674 ( .A1(n6846), .A2(n8098), .ZN(n6845) );
  NAND2_X1 U7675 ( .A1(n12832), .A2(n6590), .ZN(n7462) );
  INV_X1 U7676 ( .A(n7100), .ZN(n7099) );
  NAND2_X1 U7677 ( .A1(n7093), .A2(n11296), .ZN(n7091) );
  INV_X1 U7678 ( .A(n6761), .ZN(n6760) );
  OAI21_X1 U7679 ( .B1(n12844), .B2(n12843), .A(n6562), .ZN(n6761) );
  AND2_X1 U7680 ( .A1(n12843), .A2(n12844), .ZN(n6762) );
  INV_X1 U7681 ( .A(n11320), .ZN(n7123) );
  INV_X1 U7682 ( .A(n6789), .ZN(n6786) );
  INV_X1 U7683 ( .A(n6788), .ZN(n6787) );
  NAND2_X1 U7684 ( .A1(n11342), .A2(n6490), .ZN(n7110) );
  INV_X1 U7685 ( .A(n7114), .ZN(n7111) );
  NOR2_X1 U7686 ( .A1(n11340), .A2(n7118), .ZN(n7113) );
  OR2_X1 U7687 ( .A1(n8142), .A2(n6838), .ZN(n6837) );
  NAND2_X1 U7688 ( .A1(n6840), .A2(n6839), .ZN(n6838) );
  NAND2_X1 U7689 ( .A1(n8143), .A2(n8415), .ZN(n6839) );
  AND2_X1 U7690 ( .A1(n12882), .A2(n6747), .ZN(n6746) );
  INV_X1 U7691 ( .A(n12880), .ZN(n6747) );
  NAND2_X1 U7692 ( .A1(n6799), .A2(n6797), .ZN(n8184) );
  AND2_X1 U7693 ( .A1(n12363), .A2(n6798), .ZN(n6797) );
  NAND2_X1 U7694 ( .A1(n6801), .A2(n6800), .ZN(n6799) );
  AND2_X1 U7695 ( .A1(n8173), .A2(n8174), .ZN(n6798) );
  NAND2_X1 U7696 ( .A1(n7457), .A2(n7454), .ZN(n12908) );
  NAND2_X1 U7697 ( .A1(n7456), .A2(n7455), .ZN(n7454) );
  INV_X1 U7698 ( .A(n12903), .ZN(n7455) );
  OAI21_X1 U7699 ( .B1(n8192), .B2(n8191), .A(n8206), .ZN(n8198) );
  NOR2_X1 U7700 ( .A1(n11427), .A2(n11424), .ZN(n7137) );
  NAND2_X1 U7701 ( .A1(n11424), .A2(n11427), .ZN(n7136) );
  NAND2_X1 U7702 ( .A1(n7145), .A2(n11205), .ZN(n11499) );
  NAND2_X1 U7703 ( .A1(n11204), .A2(n11203), .ZN(n7145) );
  INV_X1 U7704 ( .A(n9348), .ZN(n9236) );
  NOR2_X1 U7705 ( .A1(n9126), .A2(n7423), .ZN(n7422) );
  INV_X1 U7706 ( .A(n8964), .ZN(n7423) );
  INV_X1 U7707 ( .A(n8825), .ZN(n7412) );
  INV_X1 U7708 ( .A(n12146), .ZN(n7344) );
  NAND2_X1 U7709 ( .A1(n11618), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n6831) );
  NAND2_X1 U7710 ( .A1(n7177), .A2(n7176), .ZN(n7175) );
  INV_X1 U7711 ( .A(P3_IR_REG_17__SCAN_IN), .ZN(n7177) );
  INV_X1 U7712 ( .A(P3_IR_REG_16__SCAN_IN), .ZN(n7176) );
  NAND2_X1 U7713 ( .A1(n12913), .A2(n12914), .ZN(n7465) );
  INV_X1 U7714 ( .A(n13231), .ZN(n6931) );
  INV_X1 U7715 ( .A(n7066), .ZN(n7060) );
  NOR2_X1 U7716 ( .A1(n11591), .A2(n7031), .ZN(n7030) );
  NOR2_X1 U7717 ( .A1(n10762), .A2(n7032), .ZN(n7031) );
  INV_X1 U7718 ( .A(n10764), .ZN(n7032) );
  NAND2_X1 U7719 ( .A1(n10535), .A2(n7436), .ZN(n7435) );
  OAI21_X1 U7720 ( .B1(n8495), .B2(n8502), .A(n8501), .ZN(n8503) );
  NAND2_X1 U7721 ( .A1(n8495), .A2(P1_DATAO_REG_3__SCAN_IN), .ZN(n8501) );
  NAND2_X1 U7722 ( .A1(n7556), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n7587) );
  NOR2_X1 U7723 ( .A1(n14976), .A2(n9221), .ZN(n9220) );
  NAND2_X1 U7724 ( .A1(n9058), .A2(P3_REG2_REG_2__SCAN_IN), .ZN(n8248) );
  OR2_X1 U7725 ( .A1(n14834), .A2(n8298), .ZN(n8300) );
  NOR2_X1 U7726 ( .A1(n7378), .A2(n6840), .ZN(n7375) );
  INV_X1 U7727 ( .A(n12451), .ZN(n7378) );
  INV_X1 U7728 ( .A(n7762), .ZN(n7377) );
  NOR2_X1 U7729 ( .A1(n12451), .A2(n7155), .ZN(n7154) );
  NAND2_X1 U7730 ( .A1(n8113), .A2(n8105), .ZN(n8110) );
  NAND2_X1 U7731 ( .A1(n12141), .A2(n9715), .ZN(n7366) );
  NAND2_X1 U7732 ( .A1(n8231), .A2(n8230), .ZN(n9546) );
  AND2_X1 U7733 ( .A1(n11067), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n7516) );
  INV_X1 U7734 ( .A(n7870), .ZN(n6815) );
  NOR2_X1 U7735 ( .A1(n7794), .A2(n7175), .ZN(n6922) );
  INV_X1 U7736 ( .A(n6820), .ZN(n6819) );
  OAI21_X1 U7737 ( .B1(n7791), .B2(n6821), .A(n7803), .ZN(n6820) );
  INV_X1 U7738 ( .A(n7508), .ZN(n6821) );
  NOR2_X1 U7739 ( .A1(n7289), .A2(n7292), .ZN(n7286) );
  NAND2_X1 U7740 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n7503), .ZN(n7504) );
  INV_X1 U7741 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n7501) );
  INV_X1 U7742 ( .A(n6780), .ZN(n6779) );
  OAI21_X1 U7743 ( .B1(n7693), .B2(n6781), .A(n7709), .ZN(n6780) );
  OR2_X1 U7744 ( .A1(n11621), .A2(n11622), .ZN(n7273) );
  NAND2_X1 U7745 ( .A1(n9328), .A2(n9327), .ZN(n9336) );
  NOR2_X1 U7746 ( .A1(n13327), .A2(n13331), .ZN(n6857) );
  AND2_X1 U7747 ( .A1(n6932), .A2(n6931), .ZN(n6930) );
  AND2_X1 U7748 ( .A1(n6934), .A2(n6931), .ZN(n6928) );
  NOR2_X1 U7749 ( .A1(n13247), .A2(n6936), .ZN(n6935) );
  INV_X1 U7750 ( .A(n6938), .ZN(n6936) );
  INV_X1 U7751 ( .A(n13044), .ZN(n12623) );
  INV_X1 U7752 ( .A(n13045), .ZN(n12691) );
  NOR2_X1 U7753 ( .A1(n7186), .A2(n6712), .ZN(n6711) );
  NOR2_X1 U7754 ( .A1(n12873), .A2(n13049), .ZN(n7186) );
  INV_X1 U7755 ( .A(n7187), .ZN(n6712) );
  INV_X1 U7756 ( .A(n13307), .ZN(n6709) );
  NOR2_X1 U7757 ( .A1(n11133), .A2(n7188), .ZN(n13306) );
  AND2_X1 U7758 ( .A1(n12851), .A2(n13051), .ZN(n7188) );
  INV_X1 U7759 ( .A(n10246), .ZN(n6943) );
  OR2_X1 U7760 ( .A1(n12842), .A2(n13053), .ZN(n10941) );
  NAND2_X1 U7761 ( .A1(n8441), .A2(n8916), .ZN(n8669) );
  INV_X1 U7762 ( .A(n14027), .ZN(n11570) );
  AND2_X1 U7763 ( .A1(n7063), .A2(n7065), .ZN(n7062) );
  XNOR2_X1 U7764 ( .A(n11572), .B(n11917), .ZN(n11916) );
  NAND2_X1 U7765 ( .A1(n14003), .A2(n11893), .ZN(n14000) );
  AND2_X1 U7766 ( .A1(n11591), .A2(n7317), .ZN(n7316) );
  OR2_X1 U7767 ( .A1(n11592), .A2(n7318), .ZN(n7317) );
  INV_X1 U7768 ( .A(n10770), .ZN(n7318) );
  AND2_X1 U7769 ( .A1(n11587), .A2(n10469), .ZN(n7056) );
  AOI21_X1 U7770 ( .B1(n10192), .B2(n14561), .A(n7323), .ZN(n7322) );
  NAND2_X1 U7771 ( .A1(n9255), .A2(n9254), .ZN(n9937) );
  INV_X1 U7772 ( .A(n7431), .ZN(n7430) );
  AOI21_X1 U7773 ( .B1(n7431), .B2(n7429), .A(n7428), .ZN(n7427) );
  INV_X1 U7774 ( .A(n11541), .ZN(n7428) );
  INV_X1 U7775 ( .A(n11480), .ZN(n7429) );
  OAI21_X1 U7776 ( .B1(n11476), .B2(n11477), .A(n11184), .ZN(n11481) );
  NAND2_X1 U7777 ( .A1(n11171), .A2(n7437), .ZN(n11430) );
  AND2_X1 U7778 ( .A1(n11174), .A2(n11170), .ZN(n7437) );
  INV_X1 U7779 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n11192) );
  OR2_X1 U7780 ( .A1(n10534), .A2(n10533), .ZN(n10700) );
  INV_X1 U7781 ( .A(n7435), .ZN(n7434) );
  AND2_X1 U7782 ( .A1(n8468), .A2(n9273), .ZN(n7025) );
  INV_X1 U7783 ( .A(n8477), .ZN(n9271) );
  NAND2_X1 U7784 ( .A1(n9933), .A2(SI_18_), .ZN(n6721) );
  INV_X1 U7785 ( .A(n9815), .ZN(n9816) );
  OR2_X1 U7786 ( .A1(n6726), .A2(n8960), .ZN(n6725) );
  AND2_X1 U7787 ( .A1(n9364), .A2(n9242), .ZN(n9362) );
  NAND2_X1 U7788 ( .A1(n8961), .A2(n8960), .ZN(n8965) );
  AOI21_X1 U7789 ( .B1(n8766), .B2(n7415), .A(n7414), .ZN(n7413) );
  INV_X1 U7790 ( .A(n8657), .ZN(n7415) );
  INV_X1 U7791 ( .A(n8768), .ZN(n7414) );
  INV_X1 U7792 ( .A(n7405), .ZN(n7404) );
  OAI21_X1 U7793 ( .B1(n8519), .B2(n7406), .A(n8556), .ZN(n7405) );
  INV_X1 U7794 ( .A(n8509), .ZN(n7406) );
  NAND2_X1 U7795 ( .A1(n8520), .A2(n8519), .ZN(n8522) );
  OR2_X1 U7796 ( .A1(n8497), .A2(n8618), .ZN(n8494) );
  INV_X1 U7797 ( .A(P3_ADDR_REG_4__SCAN_IN), .ZN(n6868) );
  INV_X1 U7798 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n14171) );
  INV_X1 U7799 ( .A(P3_ADDR_REG_3__SCAN_IN), .ZN(n14140) );
  OAI21_X1 U7800 ( .B1(P1_ADDR_REG_8__SCAN_IN), .B2(n14853), .A(n14157), .ZN(
        n14169) );
  AOI21_X1 U7801 ( .B1(n6896), .B2(n6898), .A(n6537), .ZN(n6894) );
  OR2_X1 U7802 ( .A1(n11949), .A2(n11948), .ZN(n11950) );
  NAND2_X1 U7803 ( .A1(n7732), .A2(n7731), .ZN(n7769) );
  AOI21_X1 U7804 ( .B1(n6904), .B2(n6903), .A(n6569), .ZN(n6902) );
  INV_X1 U7805 ( .A(n12077), .ZN(n6903) );
  NAND2_X1 U7806 ( .A1(n7303), .A2(n7301), .ZN(n7300) );
  AOI21_X1 U7807 ( .B1(n7306), .B2(n7304), .A(n8224), .ZN(n7303) );
  NAND2_X1 U7808 ( .A1(n7302), .A2(n8415), .ZN(n7301) );
  XNOR2_X1 U7809 ( .A(n8000), .B(P3_IR_REG_23__SCAN_IN), .ZN(n9495) );
  OAI21_X1 U7810 ( .B1(n7999), .B2(P3_IR_REG_22__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n8000) );
  AND4_X1 U7811 ( .A1(n7880), .A2(n7879), .A3(n7878), .A4(n7877), .ZN(n12026)
         );
  AND4_X1 U7812 ( .A1(n7846), .A2(n7845), .A3(n7844), .A4(n7843), .ZN(n11944)
         );
  AND4_X1 U7813 ( .A1(n7720), .A2(n7719), .A3(n7718), .A4(n7717), .ZN(n10861)
         );
  AND4_X1 U7814 ( .A1(n7603), .A2(n7602), .A3(n7601), .A4(n7600), .ZN(n10033)
         );
  NOR2_X1 U7815 ( .A1(n12605), .A2(n8003), .ZN(n9496) );
  NOR2_X1 U7816 ( .A1(n9046), .A2(n9045), .ZN(n9044) );
  OAI21_X1 U7817 ( .B1(n9067), .B2(n6958), .A(n6957), .ZN(n9174) );
  NAND2_X1 U7818 ( .A1(n6959), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n6958) );
  INV_X1 U7819 ( .A(n9175), .ZN(n6959) );
  OAI21_X1 U7820 ( .B1(n9063), .B2(n7361), .A(n7360), .ZN(n9178) );
  NAND2_X1 U7821 ( .A1(n7362), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7361) );
  INV_X1 U7822 ( .A(n9179), .ZN(n7362) );
  OR2_X1 U7823 ( .A1(n9392), .A2(n9393), .ZN(n7354) );
  OAI21_X1 U7824 ( .B1(n9386), .B2(n6961), .A(n6960), .ZN(n14816) );
  NAND2_X1 U7825 ( .A1(n6964), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n6961) );
  INV_X1 U7826 ( .A(n14817), .ZN(n6964) );
  OR2_X1 U7827 ( .A1(n9386), .A2(n9387), .ZN(n6963) );
  AND3_X1 U7828 ( .A1(n7351), .A2(n6589), .A3(n7349), .ZN(n8256) );
  NAND2_X1 U7829 ( .A1(n8269), .A2(n8356), .ZN(n8270) );
  OR2_X1 U7830 ( .A1(n12225), .A2(n12224), .ZN(n6941) );
  NOR2_X1 U7831 ( .A1(n12236), .A2(n12235), .ZN(n12241) );
  NOR2_X1 U7832 ( .A1(n12262), .A2(n12261), .ZN(n12260) );
  AND2_X1 U7833 ( .A1(n7917), .A2(n7547), .ZN(n7939) );
  AND2_X1 U7834 ( .A1(n12118), .A2(n12282), .ZN(n8401) );
  AND2_X1 U7835 ( .A1(n7967), .A2(n7966), .ZN(n7968) );
  NAND2_X1 U7836 ( .A1(n8223), .A2(n7387), .ZN(n7386) );
  AND2_X1 U7837 ( .A1(n12402), .A2(n8164), .ZN(n7180) );
  NAND2_X1 U7838 ( .A1(n12428), .A2(n8155), .ZN(n12412) );
  AOI21_X1 U7839 ( .B1(n7152), .B2(n7154), .A(n8150), .ZN(n7151) );
  INV_X1 U7840 ( .A(n7157), .ZN(n7152) );
  INV_X1 U7841 ( .A(n7154), .ZN(n7153) );
  NOR2_X1 U7842 ( .A1(n8145), .A2(n8143), .ZN(n7157) );
  AND2_X1 U7843 ( .A1(n7951), .A2(n8140), .ZN(n12473) );
  INV_X1 U7844 ( .A(n7167), .ZN(n7166) );
  AOI21_X1 U7845 ( .B1(n7165), .B2(n7167), .A(n8135), .ZN(n7164) );
  INV_X1 U7846 ( .A(n7170), .ZN(n7165) );
  AOI21_X1 U7847 ( .B1(n7373), .B2(n14898), .A(n6601), .ZN(n7372) );
  INV_X1 U7848 ( .A(n7701), .ZN(n7373) );
  INV_X1 U7849 ( .A(n10917), .ZN(n10922) );
  AND2_X1 U7850 ( .A1(n8134), .A2(n8138), .ZN(n10917) );
  NOR2_X1 U7851 ( .A1(n7171), .A2(n14898), .ZN(n7170) );
  INV_X1 U7852 ( .A(n8129), .ZN(n7171) );
  NOR2_X1 U7853 ( .A1(n10922), .A2(n7168), .ZN(n7167) );
  INV_X1 U7854 ( .A(n8131), .ZN(n7168) );
  NAND2_X1 U7855 ( .A1(n10805), .A2(n7701), .ZN(n14899) );
  NAND2_X1 U7856 ( .A1(n10807), .A2(n10806), .ZN(n10805) );
  NAND2_X1 U7857 ( .A1(n7980), .A2(n7979), .ZN(n14968) );
  INV_X1 U7858 ( .A(n9547), .ZN(n9508) );
  NAND2_X1 U7859 ( .A1(n7840), .A2(n7839), .ZN(n12518) );
  NAND2_X1 U7860 ( .A1(n7950), .A2(n8129), .ZN(n14896) );
  OR2_X1 U7861 ( .A1(n8418), .A2(n8417), .ZN(n9514) );
  INV_X1 U7862 ( .A(n9509), .ZN(n9889) );
  OR2_X1 U7863 ( .A1(n9978), .A2(n10112), .ZN(n14298) );
  INV_X1 U7864 ( .A(P3_IR_REG_28__SCAN_IN), .ZN(n7181) );
  NAND2_X1 U7865 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n14123), .ZN(n6832) );
  AND2_X2 U7866 ( .A1(n7308), .A2(n7307), .ZN(n7914) );
  NAND2_X1 U7867 ( .A1(n13439), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n7307) );
  INV_X1 U7868 ( .A(n7904), .ZN(n7309) );
  AND2_X1 U7869 ( .A1(n6767), .A2(n6528), .ZN(n7986) );
  NAND2_X1 U7870 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n10708), .ZN(n7514) );
  NAND2_X1 U7871 ( .A1(n7293), .A2(n6608), .ZN(n7294) );
  AND2_X1 U7872 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n7512), .ZN(n7848) );
  OAI21_X1 U7873 ( .B1(P2_DATAO_REG_18__SCAN_IN), .B2(n9829), .A(n7509), .ZN(
        n7834) );
  NAND2_X1 U7874 ( .A1(n6922), .A2(n6921), .ZN(n7930) );
  INV_X1 U7875 ( .A(P3_IR_REG_18__SCAN_IN), .ZN(n6921) );
  NAND2_X1 U7876 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n9251), .ZN(n7508) );
  NAND2_X1 U7877 ( .A1(n7297), .A2(n7295), .ZN(n7793) );
  NAND2_X1 U7878 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n7296), .ZN(n7295) );
  NAND2_X1 U7879 ( .A1(n7275), .A2(n7502), .ZN(n7740) );
  INV_X1 U7880 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n7499) );
  XNOR2_X1 U7881 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(P2_DATAO_REG_9__SCAN_IN), 
        .ZN(n7693) );
  NAND2_X1 U7882 ( .A1(n7498), .A2(n7497), .ZN(n7694) );
  INV_X1 U7883 ( .A(P3_IR_REG_7__SCAN_IN), .ZN(n7525) );
  OAI21_X1 U7884 ( .B1(n7647), .B2(n7493), .A(n7494), .ZN(n7664) );
  INV_X1 U7885 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n7487) );
  INV_X1 U7886 ( .A(n13055), .ZN(n14323) );
  INV_X1 U7887 ( .A(n9925), .ZN(n7258) );
  AND2_X1 U7888 ( .A1(n12698), .A2(n11631), .ZN(n7250) );
  INV_X1 U7889 ( .A(n12662), .ZN(n7249) );
  INV_X1 U7890 ( .A(n11736), .ZN(n7268) );
  INV_X1 U7891 ( .A(n7263), .ZN(n7262) );
  INV_X1 U7892 ( .A(n9481), .ZN(n7228) );
  AND2_X1 U7893 ( .A1(n9726), .A2(n7227), .ZN(n7226) );
  NAND2_X1 U7894 ( .A1(n7229), .A2(n9481), .ZN(n7227) );
  INV_X1 U7895 ( .A(n10392), .ZN(n7254) );
  AOI21_X1 U7896 ( .B1(n9925), .B2(n7257), .A(n7256), .ZN(n7255) );
  INV_X1 U7897 ( .A(n9922), .ZN(n7257) );
  INV_X1 U7898 ( .A(n9957), .ZN(n7256) );
  NAND2_X1 U7899 ( .A1(n10400), .A2(n10399), .ZN(n10496) );
  AND2_X1 U7900 ( .A1(n9157), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9198) );
  XOR2_X1 U7901 ( .A(n11750), .B(n12842), .Z(n11621) );
  INV_X1 U7902 ( .A(n6855), .ZN(n6852) );
  NOR2_X1 U7903 ( .A1(n13161), .A2(n6856), .ZN(n6855) );
  INV_X1 U7904 ( .A(n6857), .ZN(n6856) );
  NAND2_X1 U7905 ( .A1(n7211), .A2(n7207), .ZN(n7206) );
  NAND2_X1 U7906 ( .A1(n13022), .A2(n7214), .ZN(n7207) );
  INV_X1 U7907 ( .A(n7214), .ZN(n7209) );
  NAND2_X1 U7908 ( .A1(n6573), .A2(n7218), .ZN(n7216) );
  NAND2_X1 U7909 ( .A1(n6524), .A2(n11883), .ZN(n7217) );
  NAND2_X1 U7910 ( .A1(n13203), .A2(n13345), .ZN(n13202) );
  AOI22_X1 U7911 ( .A1(n13211), .A2(n13215), .B1(n12674), .B2(n13352), .ZN(
        n13201) );
  OR2_X1 U7912 ( .A1(n13352), .A2(n13043), .ZN(n11882) );
  XNOR2_X1 U7913 ( .A(n13352), .B(n13043), .ZN(n13215) );
  NAND2_X1 U7914 ( .A1(n11879), .A2(n12691), .ZN(n7201) );
  NAND2_X1 U7915 ( .A1(n11855), .A2(n13260), .ZN(n6934) );
  NAND2_X1 U7916 ( .A1(n6933), .A2(n11855), .ZN(n6932) );
  INV_X1 U7917 ( .A(n6935), .ZN(n6933) );
  OR2_X1 U7918 ( .A1(n13259), .A2(n13268), .ZN(n6937) );
  NAND2_X1 U7919 ( .A1(n6939), .A2(n13046), .ZN(n6938) );
  NOR2_X1 U7920 ( .A1(n13245), .A2(n7200), .ZN(n7199) );
  INV_X1 U7921 ( .A(n7203), .ZN(n7200) );
  NAND2_X1 U7922 ( .A1(n11877), .A2(n6700), .ZN(n13273) );
  NAND2_X1 U7923 ( .A1(n12688), .A2(n12879), .ZN(n6700) );
  AOI21_X1 U7924 ( .B1(n6968), .B2(n11139), .A(n6966), .ZN(n6965) );
  INV_X1 U7925 ( .A(n11848), .ZN(n6966) );
  NAND2_X1 U7926 ( .A1(n6860), .A2(n6859), .ZN(n13296) );
  NOR2_X1 U7927 ( .A1(n13016), .A2(n6969), .ZN(n6968) );
  INV_X1 U7928 ( .A(n11138), .ZN(n6969) );
  OR2_X1 U7929 ( .A1(n13308), .A2(n11139), .ZN(n6970) );
  OR2_X1 U7930 ( .A1(n13390), .A2(n13050), .ZN(n7187) );
  NAND2_X1 U7931 ( .A1(n13306), .A2(n13307), .ZN(n13305) );
  NAND2_X1 U7932 ( .A1(n11036), .A2(n13397), .ZN(n13313) );
  XNOR2_X1 U7933 ( .A(n14342), .B(n13054), .ZN(n14345) );
  INV_X1 U7934 ( .A(n10743), .ZN(n7196) );
  NOR2_X1 U7935 ( .A1(n14345), .A2(n7194), .ZN(n7193) );
  INV_X1 U7936 ( .A(n7197), .ZN(n7194) );
  NAND2_X1 U7937 ( .A1(n10131), .A2(n10130), .ZN(n12823) );
  NAND2_X1 U7938 ( .A1(n6691), .A2(n6497), .ZN(n6692) );
  AND2_X1 U7939 ( .A1(n10057), .A2(n10043), .ZN(n13005) );
  AND2_X1 U7940 ( .A1(n10044), .A2(n9790), .ZN(n13004) );
  NAND2_X1 U7941 ( .A1(n9791), .A2(n9767), .ZN(n13002) );
  NOR2_X1 U7942 ( .A1(n13002), .A2(n6948), .ZN(n6952) );
  INV_X1 U7943 ( .A(n9774), .ZN(n6948) );
  NAND2_X1 U7944 ( .A1(n9772), .A2(n9771), .ZN(n6953) );
  INV_X1 U7945 ( .A(n9417), .ZN(n6699) );
  NAND2_X1 U7946 ( .A1(n9197), .A2(n9203), .ZN(n9414) );
  NAND2_X1 U7947 ( .A1(n6689), .A2(n9141), .ZN(n9196) );
  INV_X1 U7948 ( .A(n14740), .ZN(n14352) );
  AND2_X1 U7949 ( .A1(n7480), .A2(n8674), .ZN(n7445) );
  OR2_X1 U7950 ( .A1(n8452), .A2(P2_IR_REG_25__SCAN_IN), .ZN(n8447) );
  NOR2_X1 U7951 ( .A1(n8669), .A2(P2_IR_REG_21__SCAN_IN), .ZN(n8664) );
  NAND2_X1 U7952 ( .A1(n6947), .A2(n8511), .ZN(n8529) );
  NAND2_X1 U7953 ( .A1(n13075), .A2(n7220), .ZN(n8535) );
  INV_X1 U7954 ( .A(P2_IR_REG_1__SCAN_IN), .ZN(n7220) );
  AND2_X1 U7955 ( .A1(n11769), .A2(n11768), .ZN(n11770) );
  NAND2_X1 U7956 ( .A1(n10459), .A2(n10458), .ZN(n11268) );
  INV_X1 U7957 ( .A(n10796), .ZN(n7010) );
  INV_X1 U7958 ( .A(n7007), .ZN(n7006) );
  OAI21_X1 U7959 ( .B1(n13510), .B2(n13592), .A(n13591), .ZN(n7007) );
  AOI21_X1 U7960 ( .B1(n7023), .B2(n11780), .A(n6494), .ZN(n7019) );
  NAND2_X1 U7961 ( .A1(n11492), .A2(n11491), .ZN(n13818) );
  OR2_X1 U7962 ( .A1(n14118), .A2(n11490), .ZN(n11492) );
  NAND2_X1 U7963 ( .A1(n6629), .A2(n6628), .ZN(n6653) );
  INV_X1 U7964 ( .A(n11923), .ZN(n6628) );
  INV_X1 U7965 ( .A(n11922), .ZN(n6629) );
  AOI21_X1 U7966 ( .B1(n7330), .B2(n13885), .A(n6564), .ZN(n7327) );
  NAND2_X1 U7967 ( .A1(n7329), .A2(n7328), .ZN(n7332) );
  INV_X1 U7968 ( .A(n13878), .ZN(n7329) );
  AND2_X1 U7969 ( .A1(n7331), .A2(n13860), .ZN(n7330) );
  INV_X1 U7970 ( .A(n7333), .ZN(n7331) );
  AND2_X1 U7971 ( .A1(n11393), .A2(n6744), .ZN(n7333) );
  AND2_X1 U7972 ( .A1(n13462), .A2(n11392), .ZN(n6744) );
  INV_X1 U7973 ( .A(n7332), .ZN(n13880) );
  OR2_X1 U7974 ( .A1(n11685), .A2(n11490), .ZN(n11393) );
  NOR2_X1 U7975 ( .A1(n7325), .A2(n13934), .ZN(n7324) );
  INV_X1 U7976 ( .A(n11916), .ZN(n13920) );
  NAND2_X1 U7977 ( .A1(n11311), .A2(n11310), .ZN(n13969) );
  NAND2_X1 U7978 ( .A1(n13975), .A2(n13976), .ZN(n7058) );
  INV_X1 U7979 ( .A(n7336), .ZN(n7335) );
  NAND2_X1 U7980 ( .A1(n10617), .A2(n10616), .ZN(n11273) );
  NAND2_X1 U7981 ( .A1(n10470), .A2(n7056), .ZN(n10614) );
  AOI21_X1 U7982 ( .B1(n7039), .B2(n7037), .A(n6552), .ZN(n7036) );
  OR2_X1 U7983 ( .A1(n11538), .A2(n13680), .ZN(n14008) );
  INV_X1 U7984 ( .A(n11581), .ZN(n7037) );
  NAND2_X1 U7985 ( .A1(n9672), .A2(n11219), .ZN(n9936) );
  NAND2_X1 U7986 ( .A1(n10153), .A2(n9678), .ZN(n9949) );
  NAND2_X1 U7987 ( .A1(n7046), .A2(n7051), .ZN(n13845) );
  NAND2_X1 U7988 ( .A1(n13884), .A2(n7049), .ZN(n7046) );
  NAND2_X1 U7989 ( .A1(n11113), .A2(n11112), .ZN(n14410) );
  AND3_X2 U7990 ( .A1(n9580), .A2(n9579), .A3(n9578), .ZN(n14550) );
  AND2_X1 U7991 ( .A1(n9665), .A2(n9664), .ZN(n9938) );
  INV_X1 U7992 ( .A(n14392), .ZN(n14542) );
  NOR2_X1 U7993 ( .A1(n11488), .A2(n7432), .ZN(n7431) );
  INV_X1 U7994 ( .A(n11485), .ZN(n7432) );
  INV_X1 U7995 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n8771) );
  AND2_X1 U7996 ( .A1(n8476), .A2(n7340), .ZN(n6876) );
  NAND2_X1 U7997 ( .A1(n7408), .A2(n15171), .ZN(n7407) );
  NAND2_X1 U7998 ( .A1(n11079), .A2(n11078), .ZN(n11166) );
  AND2_X1 U7999 ( .A1(n10962), .A2(n11060), .ZN(n11362) );
  NAND2_X1 U8000 ( .A1(n6674), .A2(n6673), .ZN(n10962) );
  INV_X1 U8001 ( .A(n11071), .ZN(n6674) );
  XNOR2_X1 U8002 ( .A(n9934), .B(n9933), .ZN(n11316) );
  NAND2_X1 U8003 ( .A1(n7439), .A2(n7438), .ZN(n9934) );
  NAND2_X1 U8004 ( .A1(n9820), .A2(n9821), .ZN(n7438) );
  NAND2_X1 U8005 ( .A1(n6720), .A2(SI_18_), .ZN(n7439) );
  AOI21_X1 U8006 ( .B1(n14182), .B2(n14181), .A(n14249), .ZN(n14185) );
  AOI22_X1 U8007 ( .A1(P3_ADDR_REG_13__SCAN_IN), .A2(n14217), .B1(n14218), 
        .B2(n14167), .ZN(n14222) );
  NAND2_X1 U8008 ( .A1(n6895), .A2(n11970), .ZN(n12017) );
  NAND2_X1 U8009 ( .A1(n7886), .A2(n7885), .ZN(n12031) );
  OR2_X1 U8010 ( .A1(n11942), .A2(n11941), .ZN(n11943) );
  OR2_X1 U8011 ( .A1(n8073), .A2(n8631), .ZN(n6806) );
  NAND2_X1 U8012 ( .A1(n7907), .A2(n7906), .ZN(n12317) );
  NAND2_X1 U8013 ( .A1(n7873), .A2(n7872), .ZN(n12355) );
  INV_X1 U8014 ( .A(n12115), .ZN(n14276) );
  NAND2_X1 U8015 ( .A1(n7782), .A2(n7781), .ZN(n14275) );
  INV_X1 U8016 ( .A(n11944), .ZN(n12126) );
  INV_X1 U8017 ( .A(n10580), .ZN(n12133) );
  XNOR2_X1 U8018 ( .A(n7633), .B(P3_IR_REG_5__SCAN_IN), .ZN(n9398) );
  OR2_X1 U8019 ( .A1(n14856), .A2(n14855), .ZN(n7348) );
  XNOR2_X1 U8020 ( .A(n7346), .B(n14877), .ZN(n14873) );
  NOR2_X1 U8021 ( .A1(n14874), .A2(n14873), .ZN(n14872) );
  XNOR2_X1 U8022 ( .A(n8270), .B(n12205), .ZN(n12198) );
  OR2_X1 U8023 ( .A1(n12234), .A2(n12233), .ZN(n7358) );
  INV_X1 U8024 ( .A(n8274), .ZN(n7357) );
  OAI21_X1 U8025 ( .B1(n12260), .B2(n6985), .A(n6984), .ZN(n6983) );
  AND2_X1 U8026 ( .A1(n12262), .A2(n12261), .ZN(n6985) );
  NOR2_X1 U8027 ( .A1(n6606), .A2(n6656), .ZN(n6655) );
  OAI21_X1 U8028 ( .B1(n14875), .B2(n12259), .A(n12258), .ZN(n6656) );
  OAI21_X1 U8029 ( .B1(n12234), .B2(n7356), .A(n7355), .ZN(n12250) );
  NAND2_X1 U8030 ( .A1(n7359), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7356) );
  INV_X1 U8031 ( .A(n12251), .ZN(n7359) );
  NOR2_X1 U8032 ( .A1(n8395), .A2(n8394), .ZN(n12286) );
  INV_X1 U8033 ( .A(n11977), .ZN(n8394) );
  NAND2_X1 U8034 ( .A1(n12282), .A2(n11164), .ZN(n7400) );
  NAND2_X1 U8035 ( .A1(n12286), .A2(n7401), .ZN(n11163) );
  NAND2_X1 U8036 ( .A1(n12283), .A2(n14983), .ZN(n7401) );
  AOI21_X1 U8037 ( .B1(n9059), .B2(n6488), .A(n7807), .ZN(n12575) );
  NAND2_X1 U8038 ( .A1(n15015), .A2(n15016), .ZN(n12583) );
  AND2_X1 U8039 ( .A1(n7995), .A2(n7994), .ZN(n12585) );
  AND2_X1 U8040 ( .A1(n7998), .A2(n7997), .ZN(n12587) );
  NAND2_X1 U8041 ( .A1(n11734), .A2(n11733), .ZN(n13339) );
  AOI21_X1 U8042 ( .B1(n12690), .B2(n12689), .A(n7481), .ZN(n12621) );
  INV_X1 U8043 ( .A(n6707), .ZN(n6706) );
  OAI21_X1 U8044 ( .B1(n12931), .B2(n9576), .A(n8892), .ZN(n6707) );
  NAND2_X1 U8045 ( .A1(n12679), .A2(n11645), .ZN(n12637) );
  AOI21_X1 U8046 ( .B1(n7238), .B2(n9693), .A(n7240), .ZN(n7239) );
  INV_X1 U8047 ( .A(n9470), .ZN(n7240) );
  NAND2_X1 U8048 ( .A1(n8899), .A2(n13441), .ZN(n8898) );
  NAND2_X1 U8049 ( .A1(n7231), .A2(n7233), .ZN(n11012) );
  AOI21_X1 U8050 ( .B1(n10498), .B2(n7235), .A(n7234), .ZN(n7233) );
  INV_X1 U8051 ( .A(n10568), .ZN(n7234) );
  INV_X1 U8052 ( .A(n12922), .ZN(n13345) );
  NAND2_X1 U8053 ( .A1(n7267), .A2(n7266), .ZN(n12707) );
  INV_X1 U8054 ( .A(n12983), .ZN(n12984) );
  NAND2_X1 U8055 ( .A1(n10593), .A2(n10594), .ZN(n10817) );
  INV_X1 U8056 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n7543) );
  AND2_X1 U8057 ( .A1(n13155), .A2(n14686), .ZN(n6633) );
  XNOR2_X1 U8058 ( .A(n13147), .B(n6634), .ZN(n13156) );
  INV_X1 U8059 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n6634) );
  OR2_X1 U8060 ( .A1(n11685), .A2(n12931), .ZN(n11687) );
  NAND2_X1 U8061 ( .A1(n10249), .A2(n10248), .ZN(n12830) );
  OAI21_X1 U8062 ( .B1(n13335), .B2(n13406), .A(n6703), .ZN(n13411) );
  AND2_X1 U8063 ( .A1(n13334), .A2(n13333), .ZN(n6703) );
  NAND2_X1 U8064 ( .A1(n8956), .A2(n8955), .ZN(n14735) );
  NOR2_X1 U8065 ( .A1(n8441), .A2(n8913), .ZN(n8914) );
  NAND2_X1 U8066 ( .A1(n9371), .A2(n8908), .ZN(n8915) );
  NAND2_X1 U8067 ( .A1(n6987), .A2(n6988), .ZN(n6993) );
  INV_X1 U8068 ( .A(n13898), .ZN(n14056) );
  NAND2_X1 U8069 ( .A1(n11330), .A2(n11329), .ZN(n14078) );
  OR2_X1 U8070 ( .A1(n9299), .A2(n9298), .ZN(n13650) );
  NAND2_X1 U8071 ( .A1(n6648), .A2(n6543), .ZN(n11612) );
  NAND2_X1 U8072 ( .A1(n11567), .A2(n11566), .ZN(n11609) );
  INV_X1 U8073 ( .A(n11563), .ZN(n11567) );
  NAND2_X1 U8074 ( .A1(n12001), .A2(n13819), .ZN(n14024) );
  NAND2_X1 U8075 ( .A1(n6653), .A2(n6668), .ZN(n6667) );
  NAND2_X1 U8076 ( .A1(n14032), .A2(n13654), .ZN(n6668) );
  NAND2_X1 U8077 ( .A1(n6653), .A2(n6652), .ZN(n14031) );
  NAND2_X1 U8078 ( .A1(n11922), .A2(n11923), .ZN(n6652) );
  NAND2_X1 U8079 ( .A1(n7074), .A2(n7073), .ZN(n7072) );
  XNOR2_X1 U8080 ( .A(n11997), .B(n11923), .ZN(n7075) );
  NAND2_X1 U8081 ( .A1(n13653), .A2(n14524), .ZN(n7074) );
  NAND2_X1 U8082 ( .A1(n10207), .A2(n10206), .ZN(n11259) );
  INV_X1 U8083 ( .A(P3_ADDR_REG_0__SCAN_IN), .ZN(n14177) );
  XNOR2_X1 U8084 ( .A(n14178), .B(n6679), .ZN(n15252) );
  INV_X1 U8085 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n6679) );
  XNOR2_X1 U8086 ( .A(n14185), .B(n6678), .ZN(n15251) );
  INV_X1 U8087 ( .A(n14184), .ZN(n6678) );
  NOR2_X1 U8088 ( .A1(n14210), .A2(n14209), .ZN(n14257) );
  INV_X1 U8089 ( .A(n14258), .ZN(n6872) );
  OAI21_X1 U8090 ( .B1(n14464), .B2(n14463), .A(P2_ADDR_REG_13__SCAN_IN), .ZN(
        n6864) );
  NOR2_X1 U8091 ( .A1(n14468), .A2(n14469), .ZN(n14467) );
  NAND2_X1 U8092 ( .A1(n7082), .A2(n11211), .ZN(n7081) );
  AOI21_X1 U8093 ( .B1(n11214), .B2(n7471), .A(n7080), .ZN(n7079) );
  AND2_X1 U8094 ( .A1(n11227), .A2(n11226), .ZN(n11232) );
  OR2_X1 U8095 ( .A1(n7142), .A2(n11248), .ZN(n7141) );
  INV_X1 U8096 ( .A(n11247), .ZN(n7142) );
  NAND2_X1 U8097 ( .A1(n6754), .A2(n6757), .ZN(n6753) );
  OAI21_X1 U8098 ( .B1(n12812), .B2(n12959), .A(n12811), .ZN(n12813) );
  INV_X1 U8099 ( .A(n12826), .ZN(n7461) );
  OR2_X1 U8100 ( .A1(n6590), .A2(n12832), .ZN(n7460) );
  NAND2_X1 U8101 ( .A1(n11272), .A2(n11269), .ZN(n7131) );
  NOR2_X1 U8102 ( .A1(n11272), .A2(n11269), .ZN(n7132) );
  AOI21_X1 U8103 ( .B1(n7102), .B2(n7104), .A(n7101), .ZN(n7100) );
  NOR2_X1 U8104 ( .A1(n7107), .A2(n7105), .ZN(n7104) );
  NOR2_X1 U8105 ( .A1(n6844), .A2(n6842), .ZN(n8112) );
  NAND2_X1 U8106 ( .A1(n6843), .A2(n10278), .ZN(n6842) );
  NAND2_X1 U8107 ( .A1(n8102), .A2(n8415), .ZN(n6843) );
  INV_X1 U8108 ( .A(n8130), .ZN(n6790) );
  AOI21_X1 U8109 ( .B1(n7094), .B2(n11288), .A(n7090), .ZN(n11300) );
  NOR2_X1 U8110 ( .A1(n7095), .A2(n6514), .ZN(n7094) );
  AOI21_X1 U8111 ( .B1(n6760), .B2(n6762), .A(n6570), .ZN(n6759) );
  INV_X1 U8112 ( .A(n8136), .ZN(n6784) );
  AOI21_X1 U8113 ( .B1(n7114), .B2(n7117), .A(n7113), .ZN(n7112) );
  NAND2_X1 U8114 ( .A1(n11340), .A2(n7118), .ZN(n7117) );
  NOR2_X1 U8115 ( .A1(n8146), .A2(n12451), .ZN(n6836) );
  OR2_X1 U8116 ( .A1(n6646), .A2(n11377), .ZN(n7089) );
  NAND2_X1 U8117 ( .A1(n6803), .A2(n6802), .ZN(n6801) );
  NAND2_X1 U8118 ( .A1(n8168), .A2(n8169), .ZN(n6802) );
  NAND2_X1 U8119 ( .A1(n6804), .A2(n12402), .ZN(n6803) );
  NOR2_X1 U8120 ( .A1(n12379), .A2(n8172), .ZN(n6800) );
  NAND2_X1 U8121 ( .A1(n6751), .A2(n6752), .ZN(n6750) );
  NOR2_X1 U8122 ( .A1(n6561), .A2(n6499), .ZN(n6748) );
  INV_X1 U8123 ( .A(n12902), .ZN(n7456) );
  INV_X1 U8124 ( .A(n8194), .ZN(n6775) );
  INV_X1 U8125 ( .A(n8196), .ZN(n7280) );
  INV_X1 U8126 ( .A(n10531), .ZN(n6718) );
  INV_X1 U8127 ( .A(n6592), .ZN(n6717) );
  AND2_X1 U8128 ( .A1(n7276), .A2(n7970), .ZN(n8206) );
  INV_X1 U8129 ( .A(n12300), .ZN(n7276) );
  OAI21_X1 U8130 ( .B1(n14912), .B2(n7163), .A(n10632), .ZN(n7162) );
  INV_X1 U8131 ( .A(n8121), .ZN(n7163) );
  INV_X1 U8132 ( .A(n9552), .ZN(n7583) );
  NAND2_X1 U8133 ( .A1(n7467), .A2(n7468), .ZN(n7466) );
  INV_X1 U8134 ( .A(n12914), .ZN(n7467) );
  AND2_X1 U8135 ( .A1(n12921), .A2(n7465), .ZN(n7463) );
  NAND2_X1 U8136 ( .A1(n12996), .A2(n9417), .ZN(n6698) );
  NOR2_X1 U8137 ( .A1(n13363), .A2(n6862), .ZN(n6861) );
  INV_X1 U8138 ( .A(n6863), .ZN(n6862) );
  AND2_X1 U8139 ( .A1(n7135), .A2(n7136), .ZN(n6672) );
  INV_X1 U8140 ( .A(n6737), .ZN(n6736) );
  OAI21_X1 U8141 ( .B1(n10703), .B2(n6738), .A(n7482), .ZN(n6737) );
  INV_X1 U8142 ( .A(n10960), .ZN(n6738) );
  INV_X1 U8143 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n8459) );
  INV_X1 U8144 ( .A(n7420), .ZN(n7419) );
  OAI21_X1 U8145 ( .B1(n7422), .B2(n7421), .A(n9231), .ZN(n7420) );
  INV_X1 U8146 ( .A(n9125), .ZN(n7421) );
  AND2_X1 U8147 ( .A1(n7410), .A2(n8824), .ZN(n7409) );
  NAND2_X1 U8148 ( .A1(n8658), .A2(n6531), .ZN(n7411) );
  INV_X1 U8149 ( .A(n11950), .ZN(n6906) );
  NAND2_X1 U8150 ( .A1(n6920), .A2(n6919), .ZN(n9716) );
  NAND2_X1 U8151 ( .A1(n6508), .A2(n9550), .ZN(n6919) );
  OR2_X1 U8152 ( .A1(n6508), .A2(n9551), .ZN(n6920) );
  NOR2_X1 U8153 ( .A1(n7305), .A2(n8415), .ZN(n7304) );
  INV_X1 U8154 ( .A(n8204), .ZN(n7305) );
  NAND2_X1 U8155 ( .A1(n7342), .A2(n7343), .ZN(n7345) );
  NOR2_X1 U8156 ( .A1(n8350), .A2(n8264), .ZN(n8265) );
  NOR2_X1 U8157 ( .A1(n8358), .A2(n12205), .ZN(n8359) );
  OAI21_X1 U8158 ( .B1(n12218), .B2(n12216), .A(n6659), .ZN(n12236) );
  INV_X1 U8159 ( .A(n12217), .ZN(n6659) );
  NAND2_X1 U8160 ( .A1(n12222), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n6940) );
  NAND2_X1 U8161 ( .A1(n7384), .A2(n7386), .ZN(n7382) );
  OR2_X1 U8162 ( .A1(n7887), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n7896) );
  NAND2_X1 U8163 ( .A1(n7961), .A2(n7960), .ZN(n12334) );
  OR2_X1 U8164 ( .A1(n8181), .A2(n12348), .ZN(n7959) );
  NOR2_X1 U8165 ( .A1(n6794), .A2(n8213), .ZN(n7371) );
  AND2_X1 U8166 ( .A1(n8114), .A2(n8119), .ZN(n14926) );
  NOR2_X1 U8167 ( .A1(n8015), .A2(n8014), .ZN(n8417) );
  AND2_X1 U8168 ( .A1(n6830), .A2(n6827), .ZN(n6826) );
  NAND2_X1 U8169 ( .A1(n7521), .A2(n6833), .ZN(n6827) );
  AND2_X1 U8170 ( .A1(n6832), .A2(n6831), .ZN(n6830) );
  AND2_X1 U8171 ( .A1(n6615), .A2(n6831), .ZN(n6829) );
  NAND2_X1 U8172 ( .A1(n6826), .A2(n6824), .ZN(n6823) );
  INV_X1 U8173 ( .A(n6833), .ZN(n6824) );
  INV_X1 U8174 ( .A(P3_IR_REG_27__SCAN_IN), .ZN(n7535) );
  NAND2_X1 U8175 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n6834), .ZN(n6833) );
  NAND2_X1 U8176 ( .A1(n7534), .A2(n7533), .ZN(n7396) );
  INV_X1 U8177 ( .A(P3_IR_REG_9__SCAN_IN), .ZN(n6769) );
  NAND2_X1 U8178 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n7510), .ZN(n7511) );
  AOI21_X1 U8179 ( .B1(n7426), .B2(n7425), .A(n6554), .ZN(n7424) );
  INV_X1 U8180 ( .A(n12969), .ZN(n7425) );
  INV_X1 U8181 ( .A(n12968), .ZN(n7426) );
  OR2_X1 U8182 ( .A1(n12963), .A2(n12962), .ZN(n12974) );
  NAND2_X1 U8183 ( .A1(n13339), .A2(n13041), .ZN(n7218) );
  OR2_X1 U8184 ( .A1(n13331), .A2(n11884), .ZN(n11859) );
  NOR2_X1 U8185 ( .A1(n13368), .A2(n12885), .ZN(n6863) );
  AND2_X1 U8186 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9146) );
  OAI21_X1 U8187 ( .B1(n8702), .B2(n8671), .A(n8672), .ZN(n6976) );
  OR2_X1 U8188 ( .A1(n8672), .A2(n8671), .ZN(n6975) );
  INV_X1 U8189 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n8456) );
  INV_X1 U8190 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n6946) );
  OR2_X1 U8191 ( .A1(n8906), .A2(n8905), .ZN(n7470) );
  NAND2_X1 U8192 ( .A1(n8886), .A2(n8885), .ZN(n8974) );
  OR2_X1 U8193 ( .A1(n8652), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n8694) );
  OR2_X1 U8194 ( .A1(n8637), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n8652) );
  AND2_X1 U8195 ( .A1(n11537), .A2(n7127), .ZN(n7126) );
  NAND2_X1 U8196 ( .A1(n11524), .A2(n11525), .ZN(n7127) );
  NAND2_X1 U8197 ( .A1(n7048), .A2(n7051), .ZN(n7047) );
  INV_X1 U8198 ( .A(n7049), .ZN(n7048) );
  INV_X1 U8199 ( .A(n13825), .ZN(n7045) );
  NOR2_X1 U8200 ( .A1(n11898), .A2(n7067), .ZN(n7066) );
  INV_X1 U8201 ( .A(n11913), .ZN(n7325) );
  NOR2_X1 U8202 ( .A1(n14078), .A2(n13969), .ZN(n6885) );
  INV_X1 U8203 ( .A(n11097), .ZN(n7337) );
  OAI21_X1 U8204 ( .B1(n7338), .B2(n7337), .A(n11905), .ZN(n7336) );
  AND2_X1 U8205 ( .A1(n11593), .A2(n10998), .ZN(n7338) );
  INV_X1 U8206 ( .A(n10613), .ZN(n7055) );
  OAI21_X1 U8207 ( .B1(n7056), .B2(n7055), .A(n11589), .ZN(n7054) );
  NAND2_X1 U8208 ( .A1(n6480), .A2(n14550), .ZN(n11213) );
  NOR2_X1 U8209 ( .A1(n13860), .A2(n7050), .ZN(n7049) );
  INV_X1 U8210 ( .A(n11899), .ZN(n7050) );
  AOI21_X1 U8211 ( .B1(n7030), .B2(n7032), .A(n6553), .ZN(n7028) );
  INV_X1 U8212 ( .A(n10304), .ZN(n6875) );
  NOR2_X1 U8213 ( .A1(n13519), .A2(n10160), .ZN(n9946) );
  INV_X1 U8214 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n8723) );
  NOR2_X1 U8215 ( .A1(P1_IR_REG_22__SCAN_IN), .A2(P1_IR_REG_23__SCAN_IN), .ZN(
        n7013) );
  NAND2_X1 U8216 ( .A1(n10704), .A2(n10703), .ZN(n10961) );
  OAI21_X1 U8217 ( .B1(P1_ADDR_REG_6__SCAN_IN), .B2(n14833), .A(n14152), .ZN(
        n14153) );
  OAI21_X1 U8218 ( .B1(P1_ADDR_REG_9__SCAN_IN), .B2(n14159), .A(n14158), .ZN(
        n14160) );
  OAI21_X1 U8219 ( .B1(P1_ADDR_REG_11__SCAN_IN), .B2(n14876), .A(n14164), .ZN(
        n14214) );
  INV_X1 U8220 ( .A(P3_REG3_REG_16__SCAN_IN), .ZN(n15210) );
  OAI21_X1 U8221 ( .B1(n10662), .B2(n6498), .A(n10661), .ZN(n10860) );
  NOR2_X1 U8222 ( .A1(n7715), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7732) );
  NOR2_X1 U8223 ( .A1(n12054), .A2(n6917), .ZN(n6916) );
  INV_X1 U8224 ( .A(n11934), .ZN(n6917) );
  AND2_X1 U8225 ( .A1(n7797), .A2(n15210), .ZN(n7808) );
  AND2_X1 U8226 ( .A1(n7670), .A2(n15058), .ZN(n7687) );
  INV_X1 U8227 ( .A(n12103), .ZN(n12440) );
  NAND2_X1 U8228 ( .A1(n7946), .A2(n8415), .ZN(n12100) );
  OR3_X1 U8229 ( .A1(n7769), .A2(P3_REG3_REG_14__SCAN_IN), .A3(
        P3_REG3_REG_13__SCAN_IN), .ZN(n7783) );
  NOR2_X1 U8230 ( .A1(n7783), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n7797) );
  OR2_X1 U8231 ( .A1(n7946), .A2(n8205), .ZN(n12103) );
  AND2_X1 U8232 ( .A1(n7922), .A2(n7921), .ZN(n11968) );
  AND4_X1 U8233 ( .A1(n7867), .A2(n7866), .A3(n7865), .A4(n7864), .ZN(n11953)
         );
  AND4_X1 U8234 ( .A1(n7858), .A2(n7857), .A3(n7856), .A4(n7855), .ZN(n11948)
         );
  AND4_X1 U8235 ( .A1(n7708), .A2(n7707), .A3(n7706), .A4(n7705), .ZN(n10580)
         );
  NOR2_X1 U8236 ( .A1(n9067), .A2(n15026), .ZN(n9066) );
  NOR2_X1 U8237 ( .A1(n9063), .A2(n9064), .ZN(n9062) );
  INV_X1 U8238 ( .A(n8300), .ZN(n8299) );
  AOI21_X1 U8239 ( .B1(n10335), .B2(n10338), .A(n10334), .ZN(n14863) );
  NAND2_X1 U8240 ( .A1(n14866), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7347) );
  NAND2_X1 U8241 ( .A1(n6956), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n6955) );
  INV_X1 U8242 ( .A(n12150), .ZN(n6956) );
  NOR2_X1 U8243 ( .A1(n14880), .A2(n14881), .ZN(n14879) );
  XNOR2_X1 U8244 ( .A(n7345), .B(n8655), .ZN(n12165) );
  OR3_X1 U8245 ( .A1(n12186), .A2(n12184), .A3(n12185), .ZN(n12187) );
  NAND2_X1 U8246 ( .A1(n6658), .A2(n6657), .ZN(n12201) );
  NAND2_X1 U8247 ( .A1(n8358), .A2(n12205), .ZN(n6657) );
  INV_X1 U8248 ( .A(n8359), .ZN(n6658) );
  NOR2_X1 U8249 ( .A1(n8363), .A2(n12241), .ZN(n8364) );
  OR2_X1 U8250 ( .A1(n12273), .A2(n7940), .ZN(n11976) );
  INV_X1 U8251 ( .A(n7925), .ZN(n7277) );
  AND2_X1 U8252 ( .A1(n8193), .A2(n12296), .ZN(n12312) );
  NAND2_X1 U8253 ( .A1(n12333), .A2(n7172), .ZN(n12294) );
  AND2_X1 U8254 ( .A1(n12326), .A2(n8188), .ZN(n7172) );
  NAND2_X1 U8255 ( .A1(n12395), .A2(n7178), .ZN(n12378) );
  NOR2_X1 U8256 ( .A1(n8170), .A2(n7179), .ZN(n7178) );
  INV_X1 U8257 ( .A(n8160), .ZN(n7179) );
  AOI21_X1 U8258 ( .B1(n12402), .B2(n7392), .A(n6502), .ZN(n7390) );
  OR2_X1 U8259 ( .A1(n7825), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7841) );
  OR2_X1 U8260 ( .A1(n12401), .A2(n12402), .ZN(n12399) );
  AND2_X1 U8261 ( .A1(n7954), .A2(n8155), .ZN(n12429) );
  AOI21_X1 U8262 ( .B1(n7377), .B2(n12451), .A(n6599), .ZN(n7376) );
  OR2_X1 U8263 ( .A1(n7702), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7715) );
  NAND2_X1 U8264 ( .A1(n14913), .A2(n14912), .ZN(n14911) );
  NOR2_X1 U8265 ( .A1(n10632), .A2(n7389), .ZN(n7388) );
  INV_X1 U8266 ( .A(n7669), .ZN(n7389) );
  NAND2_X1 U8267 ( .A1(n14914), .A2(n7669), .ZN(n10633) );
  OR2_X1 U8268 ( .A1(n7640), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7656) );
  NAND2_X1 U8269 ( .A1(n8101), .A2(n6632), .ZN(n6631) );
  INV_X1 U8270 ( .A(n14950), .ZN(n6632) );
  AOI21_X1 U8271 ( .B1(n10857), .B2(n6488), .A(n7895), .ZN(n12499) );
  NAND2_X1 U8272 ( .A1(n7852), .A2(n7851), .ZN(n11947) );
  INV_X1 U8273 ( .A(n6841), .ZN(n8316) );
  AND2_X1 U8274 ( .A1(n7985), .A2(n6510), .ZN(n8002) );
  AND2_X1 U8275 ( .A1(n6808), .A2(n6813), .ZN(n7884) );
  AOI21_X1 U8276 ( .B1(n6814), .B2(n6611), .A(n6609), .ZN(n6813) );
  OR2_X1 U8277 ( .A1(n7933), .A2(P3_IR_REG_21__SCAN_IN), .ZN(n7999) );
  NAND2_X1 U8278 ( .A1(n7935), .A2(n7937), .ZN(n7933) );
  INV_X1 U8279 ( .A(n6922), .ZN(n7835) );
  AOI21_X1 U8280 ( .B1(n6819), .B2(n6821), .A(n6610), .ZN(n6817) );
  NAND2_X1 U8281 ( .A1(n7505), .A2(n6506), .ZN(n7288) );
  OR2_X1 U8282 ( .A1(n7752), .A2(P3_IR_REG_13__SCAN_IN), .ZN(n7778) );
  AOI21_X1 U8283 ( .B1(n6779), .B2(n6781), .A(n6602), .ZN(n6777) );
  INV_X1 U8284 ( .A(n7526), .ZN(n6901) );
  INV_X1 U8285 ( .A(n7697), .ZN(n7723) );
  XNOR2_X1 U8286 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(P2_DATAO_REG_8__SCAN_IN), 
        .ZN(n7676) );
  XNOR2_X1 U8287 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .ZN(n7663) );
  INV_X1 U8288 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n7490) );
  XNOR2_X1 U8289 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(P2_DATAO_REG_5__SCAN_IN), 
        .ZN(n7630) );
  AOI21_X1 U8290 ( .B1(n7283), .B2(n7617), .A(n6565), .ZN(n7282) );
  INV_X1 U8291 ( .A(n7485), .ZN(n7283) );
  XNOR2_X1 U8292 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(P2_DATAO_REG_4__SCAN_IN), 
        .ZN(n7604) );
  NAND2_X1 U8293 ( .A1(n7230), .A2(n9476), .ZN(n7229) );
  INV_X1 U8294 ( .A(n9707), .ZN(n7230) );
  AOI21_X1 U8295 ( .B1(n7266), .B2(n7264), .A(n11724), .ZN(n7263) );
  INV_X1 U8296 ( .A(n12643), .ZN(n7264) );
  INV_X1 U8297 ( .A(n7273), .ZN(n7271) );
  AOI21_X1 U8298 ( .B1(n7273), .B2(n7270), .A(n6540), .ZN(n7269) );
  INV_X1 U8299 ( .A(n11019), .ZN(n7270) );
  OR2_X1 U8300 ( .A1(n9458), .A2(n9459), .ZN(n7242) );
  NOR2_X1 U8301 ( .A1(n9744), .A2(n9743), .ZN(n9794) );
  NAND2_X1 U8302 ( .A1(n9198), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n9744) );
  NAND2_X1 U8303 ( .A1(n7244), .A2(n7245), .ZN(n12680) );
  AOI21_X1 U8304 ( .B1(n7247), .B2(n7246), .A(n11638), .ZN(n7245) );
  INV_X1 U8305 ( .A(n7250), .ZN(n7246) );
  NOR2_X1 U8306 ( .A1(n7236), .A2(n10402), .ZN(n7232) );
  INV_X1 U8307 ( .A(n10498), .ZN(n7236) );
  INV_X1 U8308 ( .A(n10495), .ZN(n7235) );
  XNOR2_X1 U8309 ( .A(n9336), .B(n12732), .ZN(n9338) );
  NAND2_X1 U8310 ( .A1(n11749), .A2(n13067), .ZN(n9339) );
  AND2_X1 U8311 ( .A1(n9146), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9157) );
  AND2_X1 U8312 ( .A1(n12954), .A2(n12953), .ZN(n12955) );
  XNOR2_X1 U8313 ( .A(n12975), .B(n13164), .ZN(n12994) );
  NOR2_X1 U8314 ( .A1(n14646), .A2(n14645), .ZN(n14644) );
  NOR2_X1 U8315 ( .A1(n14678), .A2(n14679), .ZN(n14676) );
  NAND2_X1 U8316 ( .A1(n10483), .A2(n10482), .ZN(n10590) );
  OAI21_X1 U8317 ( .B1(n13131), .B2(n13136), .A(n13130), .ZN(n13144) );
  AND2_X1 U8318 ( .A1(n11742), .A2(n11728), .ZN(n13191) );
  XNOR2_X1 U8319 ( .A(n13339), .B(n13041), .ZN(n13189) );
  XNOR2_X1 U8320 ( .A(n12922), .B(n11856), .ZN(n13200) );
  AOI21_X1 U8321 ( .B1(n6932), .B2(n6928), .A(n6927), .ZN(n6926) );
  NOR2_X1 U8322 ( .A1(n13236), .A2(n13044), .ZN(n6927) );
  NAND2_X1 U8323 ( .A1(n13299), .A2(n6863), .ZN(n13263) );
  NAND2_X1 U8324 ( .A1(n13299), .A2(n13374), .ZN(n13276) );
  NAND2_X1 U8325 ( .A1(n13287), .A2(n11850), .ZN(n13275) );
  AOI21_X1 U8326 ( .B1(n6711), .B2(n6709), .A(n6559), .ZN(n6708) );
  INV_X1 U8327 ( .A(n6711), .ZN(n6710) );
  NOR2_X1 U8328 ( .A1(n10936), .A2(n10935), .ZN(n11037) );
  OR2_X1 U8329 ( .A1(n10747), .A2(n10746), .ZN(n10936) );
  NAND2_X1 U8330 ( .A1(n10745), .A2(n14356), .ZN(n10931) );
  INV_X1 U8331 ( .A(n7191), .ZN(n7190) );
  OAI21_X1 U8332 ( .B1(n14345), .B2(n7192), .A(n6556), .ZN(n7191) );
  NAND2_X1 U8333 ( .A1(n10742), .A2(n7197), .ZN(n7192) );
  XNOR2_X1 U8334 ( .A(n12842), .B(n10740), .ZN(n13010) );
  OR2_X1 U8335 ( .A1(n10064), .A2(n10500), .ZN(n10257) );
  NOR2_X1 U8336 ( .A1(n10722), .A2(n6943), .ZN(n6942) );
  NAND2_X1 U8337 ( .A1(n10254), .A2(n10741), .ZN(n14346) );
  AOI21_X1 U8338 ( .B1(n10072), .B2(n7184), .A(n6538), .ZN(n7183) );
  INV_X1 U8339 ( .A(n10041), .ZN(n7184) );
  NAND2_X1 U8340 ( .A1(n10040), .A2(n6532), .ZN(n6691) );
  OAI21_X1 U8341 ( .B1(n9772), .B2(n6951), .A(n6949), .ZN(n9793) );
  INV_X1 U8342 ( .A(n6952), .ZN(n6951) );
  AOI21_X1 U8343 ( .B1(n6952), .B2(n9770), .A(n6950), .ZN(n6949) );
  INV_X1 U8344 ( .A(n9791), .ZN(n6950) );
  OAI21_X1 U8345 ( .B1(n9155), .B2(n14712), .A(n6923), .ZN(n9187) );
  AOI21_X1 U8346 ( .B1(n14701), .B2(n6924), .A(n6525), .ZN(n6923) );
  INV_X1 U8347 ( .A(n9154), .ZN(n6924) );
  NAND2_X1 U8348 ( .A1(n9097), .A2(P1_DATAO_REG_2__SCAN_IN), .ZN(n7443) );
  NAND2_X1 U8349 ( .A1(n9035), .A2(n12732), .ZN(n9027) );
  NAND2_X1 U8350 ( .A1(n9020), .A2(n12995), .ZN(n9023) );
  NOR2_X1 U8351 ( .A1(n13253), .A2(n9329), .ZN(n9315) );
  AND2_X1 U8352 ( .A1(n9324), .A2(n8677), .ZN(n12711) );
  NAND2_X1 U8353 ( .A1(n11864), .A2(n11863), .ZN(n13327) );
  INV_X1 U8354 ( .A(n14768), .ZN(n13406) );
  INV_X1 U8355 ( .A(n14788), .ZN(n14774) );
  NAND2_X1 U8356 ( .A1(n14788), .A2(n12732), .ZN(n8930) );
  NOR2_X1 U8357 ( .A1(n8702), .A2(n6546), .ZN(n6977) );
  NAND2_X1 U8358 ( .A1(n8673), .A2(n6705), .ZN(n6973) );
  NOR2_X1 U8359 ( .A1(n8674), .A2(n8671), .ZN(n6705) );
  AND2_X1 U8360 ( .A1(n8442), .A2(n8456), .ZN(n8449) );
  INV_X1 U8361 ( .A(n8668), .ZN(n8442) );
  OR2_X1 U8362 ( .A1(n9212), .A2(P2_IR_REG_13__SCAN_IN), .ZN(n9354) );
  INV_X1 U8363 ( .A(n8535), .ZN(n7219) );
  NAND2_X1 U8364 ( .A1(n11378), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11395) );
  AOI21_X1 U8365 ( .B1(n13493), .B2(n13490), .A(n13533), .ZN(n7002) );
  INV_X1 U8366 ( .A(n7002), .ZN(n7000) );
  INV_X1 U8367 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n10180) );
  OR2_X1 U8368 ( .A1(n10606), .A2(n10605), .ZN(n10685) );
  INV_X1 U8369 ( .A(n13563), .ZN(n7005) );
  AND2_X1 U8370 ( .A1(n13480), .A2(n13478), .ZN(n13561) );
  AND2_X1 U8371 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_REG3_REG_3__SCAN_IN), 
        .ZN(n9633) );
  OR2_X1 U8372 ( .A1(n10989), .A2(n10988), .ZN(n11100) );
  NAND2_X1 U8373 ( .A1(P1_REG3_REG_24__SCAN_IN), .A2(n11396), .ZN(n11413) );
  AND2_X1 U8374 ( .A1(n13563), .A2(n13468), .ZN(n13591) );
  NAND2_X1 U8375 ( .A1(n13509), .A2(n13510), .ZN(n13590) );
  OAI21_X1 U8376 ( .B1(n13509), .B2(n13592), .A(n7006), .ZN(n13560) );
  OR2_X1 U8377 ( .A1(n10181), .A2(n10180), .ZN(n10209) );
  INV_X1 U8378 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n10208) );
  NAND2_X1 U8379 ( .A1(n6619), .A2(n6617), .ZN(n9294) );
  AOI21_X1 U8380 ( .B1(n9619), .B2(n9668), .A(n6618), .ZN(n6617) );
  NAND2_X1 U8381 ( .A1(n14526), .A2(n13485), .ZN(n6619) );
  NOR2_X1 U8382 ( .A1(n9284), .A2(n13671), .ZN(n6618) );
  AND2_X1 U8383 ( .A1(n11365), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11378) );
  NAND2_X1 U8384 ( .A1(n10461), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10606) );
  NAND2_X1 U8385 ( .A1(n10890), .A2(n10887), .ZN(n10908) );
  NOR2_X1 U8386 ( .A1(n11100), .A2(n11099), .ZN(n11101) );
  AND2_X1 U8387 ( .A1(n11101), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n11312) );
  NOR2_X1 U8388 ( .A1(n10775), .A2(n10774), .ZN(n10981) );
  AND2_X1 U8389 ( .A1(n11568), .A2(n11555), .ZN(n6649) );
  AND2_X1 U8390 ( .A1(n11558), .A2(n11559), .ZN(n6647) );
  NOR3_X1 U8391 ( .A1(n11603), .A2(n11998), .A3(n11602), .ZN(n11604) );
  AND4_X1 U8392 ( .A1(n11520), .A2(n11519), .A3(n11518), .A4(n11517), .ZN(
        n11569) );
  AND4_X1 U8393 ( .A1(n10986), .A2(n10985), .A3(n10984), .A4(n10983), .ZN(
        n13504) );
  NOR2_X1 U8394 ( .A1(n9594), .A2(n14533), .ZN(n6671) );
  OR2_X1 U8395 ( .A1(n8612), .A2(P1_IR_REG_6__SCAN_IN), .ZN(n8600) );
  XNOR2_X1 U8396 ( .A(n14032), .B(n13654), .ZN(n11923) );
  NAND2_X1 U8397 ( .A1(n11571), .A2(n13825), .ZN(n13842) );
  NAND2_X1 U8398 ( .A1(n13905), .A2(n14056), .ZN(n13883) );
  NAND2_X1 U8399 ( .A1(n13905), .A2(n6493), .ZN(n13864) );
  AND2_X1 U8400 ( .A1(n13903), .A2(n11918), .ZN(n7334) );
  NAND2_X1 U8401 ( .A1(n6572), .A2(n7070), .ZN(n7065) );
  NAND2_X1 U8402 ( .A1(n13933), .A2(n7066), .ZN(n7064) );
  NAND2_X1 U8403 ( .A1(n7064), .A2(n7062), .ZN(n13909) );
  NOR2_X1 U8404 ( .A1(n14062), .A2(n13922), .ZN(n13905) );
  NAND2_X1 U8405 ( .A1(n13983), .A2(n6881), .ZN(n13922) );
  NOR2_X1 U8406 ( .A1(n6886), .A2(n6883), .ZN(n6881) );
  NAND2_X1 U8407 ( .A1(n13983), .A2(n6885), .ZN(n13952) );
  NAND2_X1 U8408 ( .A1(n13983), .A2(n14083), .ZN(n13965) );
  NAND2_X1 U8409 ( .A1(n7474), .A2(n7338), .ZN(n11098) );
  AOI21_X1 U8410 ( .B1(n7316), .B2(n7318), .A(n6551), .ZN(n7314) );
  INV_X1 U8411 ( .A(n6888), .ZN(n14381) );
  NOR2_X1 U8412 ( .A1(n10623), .A2(n11273), .ZN(n10694) );
  OR2_X1 U8413 ( .A1(n10460), .A2(n11268), .ZN(n10623) );
  NOR2_X1 U8414 ( .A1(n10209), .A2(n10208), .ZN(n10228) );
  AND2_X1 U8415 ( .A1(n10228), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10461) );
  OR2_X1 U8416 ( .A1(n10369), .A2(n11259), .ZN(n10460) );
  NAND2_X1 U8417 ( .A1(n10370), .A2(n14589), .ZN(n10369) );
  NAND2_X1 U8418 ( .A1(n7041), .A2(n10222), .ZN(n10314) );
  NAND2_X1 U8419 ( .A1(n10285), .A2(n11581), .ZN(n7041) );
  NAND2_X1 U8420 ( .A1(n7321), .A2(n7319), .ZN(n10297) );
  NAND2_X1 U8421 ( .A1(n7320), .A2(n6522), .ZN(n7319) );
  INV_X1 U8422 ( .A(n7322), .ZN(n7320) );
  NAND2_X1 U8423 ( .A1(n7026), .A2(n11221), .ZN(n10216) );
  INV_X1 U8424 ( .A(n14023), .ZN(n14523) );
  NOR2_X1 U8425 ( .A1(n6469), .A2(n11204), .ZN(n13881) );
  INV_X1 U8426 ( .A(n14008), .ZN(n14524) );
  INV_X1 U8427 ( .A(n9945), .ZN(n12004) );
  NAND2_X1 U8428 ( .A1(n11308), .A2(n11307), .ZN(n14090) );
  NAND2_X1 U8429 ( .A1(n10470), .A2(n10469), .ZN(n10471) );
  AOI22_X1 U8430 ( .A1(n9599), .A2(n9017), .B1(n11317), .B2(n13689), .ZN(n7071) );
  INV_X1 U8431 ( .A(n8733), .ZN(n8734) );
  NAND2_X1 U8432 ( .A1(n9284), .A2(n8738), .ZN(n9301) );
  XNOR2_X1 U8433 ( .A(n11546), .B(n11545), .ZN(n12944) );
  OAI21_X1 U8434 ( .B1(n11481), .B2(n7430), .A(n7427), .ZN(n11546) );
  INV_X1 U8435 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n8774) );
  XNOR2_X1 U8436 ( .A(n11476), .B(n11477), .ZN(n11737) );
  XNOR2_X1 U8437 ( .A(n11457), .B(n11459), .ZN(n13431) );
  NAND2_X1 U8438 ( .A1(n8477), .A2(n8476), .ZN(n8479) );
  AND2_X1 U8439 ( .A1(n8476), .A2(n7077), .ZN(n7076) );
  AND2_X1 U8440 ( .A1(n11430), .A2(n11429), .ZN(n13434) );
  NAND2_X1 U8441 ( .A1(n11171), .A2(n11170), .ZN(n11172) );
  NAND2_X1 U8442 ( .A1(n8470), .A2(n11192), .ZN(n8484) );
  INV_X1 U8443 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n8469) );
  NAND2_X1 U8444 ( .A1(n7434), .A2(n10700), .ZN(n10701) );
  NAND2_X1 U8445 ( .A1(n10700), .A2(n10535), .ZN(n10537) );
  NAND2_X1 U8446 ( .A1(n14111), .A2(n9273), .ZN(n9272) );
  NOR2_X1 U8447 ( .A1(n9273), .A2(n14111), .ZN(n7144) );
  NAND2_X1 U8448 ( .A1(n6719), .A2(n6721), .ZN(n10532) );
  NAND2_X1 U8449 ( .A1(n6720), .A2(n6592), .ZN(n6719) );
  AND2_X1 U8450 ( .A1(n9130), .A2(n8972), .ZN(n10766) );
  NAND2_X1 U8451 ( .A1(n8965), .A2(n8964), .ZN(n9127) );
  OR2_X1 U8452 ( .A1(n8827), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n8828) );
  OAI21_X1 U8453 ( .B1(n8658), .B2(n7416), .A(n7413), .ZN(n8826) );
  NAND2_X1 U8454 ( .A1(n8641), .A2(n8640), .ZN(n8645) );
  NOR2_X1 U8455 ( .A1(n8600), .A2(P1_IR_REG_7__SCAN_IN), .ZN(n8603) );
  INV_X1 U8456 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n8602) );
  AOI21_X1 U8457 ( .B1(n7404), .B2(n7406), .A(n7403), .ZN(n7402) );
  INV_X1 U8458 ( .A(n8558), .ZN(n7403) );
  NAND2_X1 U8459 ( .A1(n8522), .A2(n8509), .ZN(n8557) );
  INV_X1 U8460 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n8464) );
  NAND2_X1 U8461 ( .A1(n8490), .A2(SI_0_), .ZN(n8532) );
  NAND2_X1 U8462 ( .A1(n8495), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n6731) );
  NAND2_X1 U8463 ( .A1(n14138), .A2(n6636), .ZN(n14174) );
  NAND2_X1 U8464 ( .A1(P3_ADDR_REG_1__SCAN_IN), .A2(n6637), .ZN(n6636) );
  INV_X1 U8465 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6637) );
  XOR2_X1 U8466 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(n14139), .Z(n14173) );
  XNOR2_X1 U8467 ( .A(n14170), .B(n14171), .ZN(n14172) );
  NAND2_X1 U8468 ( .A1(n14254), .A2(n14253), .ZN(n6866) );
  INV_X1 U8469 ( .A(n6635), .ZN(n14207) );
  AOI21_X1 U8470 ( .B1(n14256), .B2(P2_ADDR_REG_9__SCAN_IN), .A(n7477), .ZN(
        n14210) );
  AND2_X1 U8471 ( .A1(n14207), .A2(n14206), .ZN(n7477) );
  NAND2_X1 U8472 ( .A1(n14458), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n6871) );
  OR2_X1 U8473 ( .A1(n14458), .A2(P2_ADDR_REG_11__SCAN_IN), .ZN(n6870) );
  OAI21_X1 U8474 ( .B1(P3_ADDR_REG_14__SCAN_IN), .B2(n14225), .A(n14224), .ZN(
        n14230) );
  NAND2_X1 U8475 ( .A1(n6910), .A2(n6908), .ZN(n10875) );
  NAND2_X1 U8476 ( .A1(n6909), .A2(n6491), .ZN(n6908) );
  NAND2_X1 U8477 ( .A1(n6912), .A2(n6548), .ZN(n6909) );
  OAI21_X1 U8478 ( .B1(n6534), .B2(n6899), .A(n6891), .ZN(n6890) );
  INV_X1 U8479 ( .A(n6896), .ZN(n6892) );
  NAND2_X1 U8480 ( .A1(n11975), .A2(n6894), .ZN(n6893) );
  NAND2_X1 U8481 ( .A1(n12076), .A2(n11950), .ZN(n12040) );
  NAND2_X1 U8482 ( .A1(n14277), .A2(n11934), .ZN(n12053) );
  NAND2_X1 U8483 ( .A1(n6918), .A2(n6915), .ZN(n12060) );
  AND2_X1 U8484 ( .A1(n12061), .A2(n6496), .ZN(n6915) );
  AND2_X1 U8485 ( .A1(n6918), .A2(n6496), .ZN(n12062) );
  NAND2_X1 U8486 ( .A1(n11958), .A2(n11957), .ZN(n11959) );
  OR2_X1 U8487 ( .A1(n11945), .A2(n11944), .ZN(n11946) );
  NAND2_X1 U8488 ( .A1(n12078), .A2(n12077), .ZN(n12076) );
  NAND2_X1 U8489 ( .A1(n6911), .A2(n6912), .ZN(n10870) );
  NAND2_X1 U8490 ( .A1(n10662), .A2(n6913), .ZN(n6911) );
  NAND2_X1 U8491 ( .A1(n9518), .A2(n9889), .ZN(n12115) );
  NAND2_X1 U8492 ( .A1(n11965), .A2(n12071), .ZN(n11966) );
  NAND2_X1 U8493 ( .A1(n7916), .A2(n7915), .ZN(n12304) );
  AND2_X1 U8494 ( .A1(n9505), .A2(n9504), .ZN(n14286) );
  AND2_X1 U8495 ( .A1(n9507), .A2(n9506), .ZN(n14274) );
  INV_X1 U8496 ( .A(n11968), .ZN(n12119) );
  INV_X1 U8497 ( .A(n12026), .ZN(n12123) );
  INV_X1 U8498 ( .A(n11953), .ZN(n12124) );
  INV_X1 U8499 ( .A(n11948), .ZN(n12125) );
  INV_X1 U8500 ( .A(n11941), .ZN(n12127) );
  NAND4_X1 U8501 ( .A1(n7737), .A2(n7736), .A3(n7735), .A4(n7734), .ZN(n12131)
         );
  INV_X1 U8502 ( .A(n10861), .ZN(n12132) );
  INV_X1 U8503 ( .A(n12101), .ZN(n12136) );
  NAND4_X1 U8504 ( .A1(n7577), .A2(n7576), .A3(n7575), .A4(n7574), .ZN(n12144)
         );
  OR2_X1 U8505 ( .A1(n8245), .A2(n12586), .ZN(n12143) );
  XNOR2_X1 U8506 ( .A(n8330), .B(n8328), .ZN(n9217) );
  XNOR2_X1 U8507 ( .A(n7619), .B(P3_IR_REG_3__SCAN_IN), .ZN(n9072) );
  INV_X1 U8508 ( .A(n6963), .ZN(n9385) );
  INV_X1 U8509 ( .A(P3_ADDR_REG_6__SCAN_IN), .ZN(n14833) );
  AND2_X1 U8510 ( .A1(n7354), .A2(n7353), .ZN(n14820) );
  NAND2_X1 U8511 ( .A1(n7349), .A2(n7351), .ZN(n14818) );
  INV_X1 U8512 ( .A(n8292), .ZN(n6962) );
  NOR2_X1 U8513 ( .A1(n9896), .A2(n9895), .ZN(n9894) );
  INV_X1 U8514 ( .A(P3_ADDR_REG_8__SCAN_IN), .ZN(n14853) );
  XNOR2_X1 U8515 ( .A(n8259), .B(n6680), .ZN(n10332) );
  NOR2_X1 U8516 ( .A1(n12147), .A2(n12146), .ZN(n12145) );
  NOR2_X1 U8517 ( .A1(n14872), .A2(n8263), .ZN(n12147) );
  NOR2_X1 U8518 ( .A1(n12163), .A2(n14303), .ZN(n12162) );
  NOR2_X1 U8519 ( .A1(n12198), .A2(n12199), .ZN(n12197) );
  INV_X1 U8520 ( .A(n6941), .ZN(n12223) );
  NAND2_X1 U8521 ( .A1(n7365), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7364) );
  NAND2_X1 U8522 ( .A1(n8271), .A2(n7365), .ZN(n7363) );
  INV_X1 U8523 ( .A(n12215), .ZN(n7365) );
  AOI21_X1 U8524 ( .B1(n12592), .B2(n7616), .A(n8074), .ZN(n14288) );
  AND2_X1 U8525 ( .A1(n8049), .A2(n8048), .ZN(n14292) );
  INV_X1 U8526 ( .A(n12499), .ZN(n12330) );
  OAI21_X1 U8527 ( .B1(n12351), .B2(n7386), .A(n7384), .ZN(n12323) );
  NAND2_X1 U8528 ( .A1(n12395), .A2(n8160), .ZN(n12385) );
  NAND2_X1 U8529 ( .A1(n12410), .A2(n8164), .ZN(n12397) );
  OAI21_X1 U8530 ( .B1(n7952), .B2(n7153), .A(n7151), .ZN(n12444) );
  NAND2_X1 U8531 ( .A1(n7379), .A2(n7762), .ZN(n12452) );
  NAND2_X1 U8532 ( .A1(n12465), .A2(n12464), .ZN(n7379) );
  NAND2_X1 U8533 ( .A1(n7156), .A2(n8144), .ZN(n12450) );
  NAND2_X1 U8534 ( .A1(n7952), .A2(n7157), .ZN(n7156) );
  NAND2_X1 U8535 ( .A1(n7952), .A2(n7951), .ZN(n12463) );
  INV_X1 U8536 ( .A(n12458), .ZN(n12479) );
  NAND2_X1 U8537 ( .A1(n7169), .A2(n7167), .ZN(n10916) );
  NAND2_X1 U8538 ( .A1(n7950), .A2(n7170), .ZN(n7169) );
  NAND2_X1 U8539 ( .A1(n14899), .A2(n14898), .ZN(n14897) );
  NAND2_X1 U8540 ( .A1(n10640), .A2(n10113), .ZN(n14941) );
  NAND2_X1 U8541 ( .A1(n9889), .A2(n9888), .ZN(n14959) );
  NAND2_X1 U8542 ( .A1(n12479), .A2(n15016), .ZN(n14906) );
  AND2_X2 U8543 ( .A1(n9887), .A2(n8024), .ZN(n15038) );
  INV_X1 U8544 ( .A(n15038), .ZN(n15036) );
  INV_X1 U8545 ( .A(P3_REG0_REG_28__SCAN_IN), .ZN(n7399) );
  INV_X1 U8546 ( .A(n12031), .ZN(n12554) );
  AOI21_X1 U8547 ( .B1(n8958), .B2(n7616), .A(n7796), .ZN(n12579) );
  NAND2_X1 U8548 ( .A1(n8279), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12586) );
  INV_X1 U8549 ( .A(P3_IR_REG_29__SCAN_IN), .ZN(n7551) );
  XNOR2_X1 U8550 ( .A(n8045), .B(n8036), .ZN(n12597) );
  OAI21_X1 U8551 ( .B1(n8027), .B2(n8028), .A(n6832), .ZN(n8035) );
  INV_X1 U8552 ( .A(n8316), .ZN(n12602) );
  XNOR2_X1 U8553 ( .A(n8027), .B(n7523), .ZN(n12601) );
  MUX2_X1 U8554 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7982), .S(
        P3_IR_REG_26__SCAN_IN), .Z(n7983) );
  INV_X1 U8555 ( .A(n8002), .ZN(n10899) );
  NAND2_X1 U8556 ( .A1(n7848), .A2(n7861), .ZN(n6812) );
  NAND2_X1 U8557 ( .A1(n7513), .A2(n7861), .ZN(n6811) );
  OR2_X1 U8558 ( .A1(n7848), .A2(n7513), .ZN(n7862) );
  XNOR2_X1 U8559 ( .A(n7837), .B(n7836), .ZN(n9360) );
  INV_X1 U8560 ( .A(SI_17_), .ZN(n15072) );
  NAND2_X1 U8561 ( .A1(n6818), .A2(n7508), .ZN(n7804) );
  NAND2_X1 U8562 ( .A1(n7793), .A2(n7791), .ZN(n6818) );
  INV_X1 U8563 ( .A(SI_16_), .ZN(n15144) );
  INV_X1 U8564 ( .A(n8312), .ZN(n12222) );
  INV_X1 U8565 ( .A(SI_15_), .ZN(n15194) );
  INV_X1 U8566 ( .A(n8310), .ZN(n12205) );
  INV_X1 U8567 ( .A(n12193), .ZN(n8692) );
  NAND2_X1 U8568 ( .A1(n7505), .A2(n6505), .ZN(n7290) );
  NAND2_X1 U8569 ( .A1(n7287), .A2(P2_DATAO_REG_13__SCAN_IN), .ZN(n7291) );
  INV_X1 U8570 ( .A(SI_12_), .ZN(n15174) );
  INV_X1 U8571 ( .A(SI_11_), .ZN(n15209) );
  NAND2_X1 U8572 ( .A1(n6778), .A2(n7500), .ZN(n7710) );
  NAND2_X1 U8573 ( .A1(n7694), .A2(n7693), .ZN(n6778) );
  NOR2_X1 U8574 ( .A1(n7608), .A2(n7526), .ZN(n7679) );
  XNOR2_X1 U8575 ( .A(n7651), .B(n7650), .ZN(n8620) );
  NAND2_X1 U8576 ( .A1(n7486), .A2(n7485), .ZN(n7618) );
  NAND3_X1 U8577 ( .A1(n7570), .A2(P3_IR_REG_2__SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n6982) );
  MUX2_X1 U8578 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7569), .S(
        P3_IR_REG_1__SCAN_IN), .Z(n7571) );
  NAND2_X1 U8579 ( .A1(P3_IR_REG_0__SCAN_IN), .A2(P3_IR_REG_31__SCAN_IN), .ZN(
        n7569) );
  INV_X1 U8580 ( .A(n7224), .ZN(n9727) );
  AOI21_X1 U8581 ( .B1(n9698), .B2(n7225), .A(n7228), .ZN(n7224) );
  INV_X1 U8582 ( .A(n7229), .ZN(n7225) );
  OAI21_X1 U8583 ( .B1(n9923), .B2(n7258), .A(n7255), .ZN(n10393) );
  NAND2_X1 U8584 ( .A1(n7248), .A2(n7247), .ZN(n12628) );
  AND2_X1 U8585 ( .A1(n7248), .A2(n6529), .ZN(n12630) );
  NAND2_X1 U8586 ( .A1(n7249), .A2(n7250), .ZN(n7248) );
  AOI21_X1 U8587 ( .B1(n7261), .B2(n7265), .A(n6571), .ZN(n7260) );
  INV_X1 U8588 ( .A(n7226), .ZN(n7222) );
  AOI21_X1 U8589 ( .B1(n7226), .B2(n7228), .A(n6533), .ZN(n7221) );
  NAND2_X1 U8590 ( .A1(n11986), .A2(n11985), .ZN(n11984) );
  NAND2_X1 U8591 ( .A1(n10497), .A2(n10498), .ZN(n10569) );
  NAND2_X1 U8592 ( .A1(n10496), .A2(n10495), .ZN(n10497) );
  INV_X1 U8593 ( .A(n7272), .ZN(n12653) );
  OAI21_X1 U8594 ( .B1(n14325), .B2(n7271), .A(n7269), .ZN(n7272) );
  NAND2_X1 U8595 ( .A1(n11029), .A2(n11028), .ZN(n12851) );
  AND2_X1 U8596 ( .A1(n7242), .A2(n7243), .ZN(n9694) );
  NAND2_X1 U8597 ( .A1(n7242), .A2(n7241), .ZN(n9692) );
  NAND2_X1 U8598 ( .A1(n9923), .A2(n9922), .ZN(n9924) );
  NAND2_X1 U8599 ( .A1(n9924), .A2(n9925), .ZN(n9958) );
  INV_X1 U8600 ( .A(n12830), .ZN(n10741) );
  INV_X1 U8601 ( .A(n11672), .ZN(n11662) );
  OR2_X1 U8602 ( .A1(n10391), .A2(n10390), .ZN(n7252) );
  NOR2_X1 U8603 ( .A1(n12662), .A2(n11632), .ZN(n12699) );
  NAND2_X1 U8604 ( .A1(n14325), .A2(n11019), .ZN(n7274) );
  OAI21_X1 U8605 ( .B1(n9323), .B2(n9313), .A(n14706), .ZN(n12703) );
  NAND2_X1 U8606 ( .A1(n12993), .A2(n12987), .ZN(n12992) );
  OR2_X1 U8607 ( .A1(n8686), .A2(n8685), .ZN(n8758) );
  AOI21_X1 U8608 ( .B1(n14660), .B2(n13083), .A(n13082), .ZN(n13101) );
  AND2_X1 U8609 ( .A1(n8997), .A2(n8996), .ZN(n9079) );
  AND2_X1 U8610 ( .A1(n13124), .A2(n13123), .ZN(n13125) );
  AOI21_X1 U8611 ( .B1(n10009), .B2(n13120), .A(n13119), .ZN(n14695) );
  XOR2_X1 U8612 ( .A(n10730), .B(n10590), .Z(n10484) );
  NAND2_X1 U8613 ( .A1(n10817), .A2(n6614), .ZN(n10819) );
  NAND2_X1 U8614 ( .A1(n6852), .A2(n6858), .ZN(n6851) );
  AND2_X1 U8615 ( .A1(n11740), .A2(P2_REG3_REG_28__SCAN_IN), .ZN(n11887) );
  NAND2_X1 U8616 ( .A1(n7209), .A2(n11885), .ZN(n7208) );
  OAI21_X1 U8617 ( .B1(n7211), .B2(n11885), .A(n7206), .ZN(n7205) );
  NAND2_X1 U8618 ( .A1(n11700), .A2(n11699), .ZN(n13352) );
  AND2_X1 U8619 ( .A1(n7202), .A2(n7201), .ZN(n13232) );
  NAND2_X1 U8620 ( .A1(n6925), .A2(n6932), .ZN(n13227) );
  OR2_X1 U8621 ( .A1(n13259), .A2(n6934), .ZN(n6925) );
  NAND2_X1 U8622 ( .A1(n6937), .A2(n6938), .ZN(n13246) );
  NAND2_X1 U8623 ( .A1(n13267), .A2(n7203), .ZN(n13244) );
  NAND2_X1 U8624 ( .A1(n6970), .A2(n6968), .ZN(n11849) );
  NAND2_X1 U8625 ( .A1(n13305), .A2(n7187), .ZN(n11876) );
  NAND2_X1 U8626 ( .A1(n11132), .A2(n11131), .ZN(n13390) );
  NAND2_X1 U8627 ( .A1(n10930), .A2(n10929), .ZN(n13404) );
  NAND2_X1 U8628 ( .A1(n7195), .A2(n7197), .ZN(n14344) );
  AND2_X1 U8629 ( .A1(n7195), .A2(n7193), .ZN(n14343) );
  NAND2_X1 U8630 ( .A1(n7196), .A2(n7198), .ZN(n7195) );
  NAND2_X1 U8631 ( .A1(n6944), .A2(n10246), .ZN(n10721) );
  NAND2_X1 U8632 ( .A1(n10040), .A2(n10039), .ZN(n7185) );
  NAND2_X1 U8633 ( .A1(n6953), .A2(n6952), .ZN(n9792) );
  AOI21_X1 U8634 ( .B1(n9416), .B2(n9415), .A(n6699), .ZN(n6697) );
  NAND2_X1 U8635 ( .A1(n9155), .A2(n9154), .ZN(n14700) );
  INV_X1 U8636 ( .A(n14721), .ZN(n14341) );
  INV_X1 U8637 ( .A(n13282), .ZN(n14725) );
  NAND2_X1 U8638 ( .A1(n12732), .A2(n14743), .ZN(n8928) );
  INV_X1 U8639 ( .A(n14743), .ZN(n9441) );
  OR2_X1 U8640 ( .A1(n14731), .A2(n9313), .ZN(n14721) );
  INV_X1 U8641 ( .A(n13304), .ZN(n14727) );
  NAND2_X1 U8642 ( .A1(n9105), .A2(n14706), .ZN(n13316) );
  AND2_X1 U8643 ( .A1(n9319), .A2(n8940), .ZN(n14736) );
  NAND2_X1 U8644 ( .A1(n8673), .A2(n8445), .ZN(n13435) );
  NAND2_X1 U8645 ( .A1(n8667), .A2(n8666), .ZN(n6745) );
  NAND2_X1 U8646 ( .A1(n8665), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8666) );
  OAI21_X1 U8647 ( .B1(n8664), .B2(n8671), .A(P2_IR_REG_22__SCAN_IN), .ZN(
        n8667) );
  NAND2_X1 U8648 ( .A1(n8909), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8917) );
  INV_X1 U8649 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n8564) );
  INV_X1 U8650 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n8531) );
  INV_X1 U8651 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n8537) );
  NAND2_X1 U8652 ( .A1(n8536), .A2(n8535), .ZN(n13069) );
  NAND2_X1 U8653 ( .A1(n10846), .A2(n10845), .ZN(n10890) );
  NAND2_X1 U8654 ( .A1(n6991), .A2(n6986), .ZN(n13518) );
  NAND2_X1 U8655 ( .A1(n6993), .A2(n6992), .ZN(n6991) );
  INV_X1 U8656 ( .A(n6994), .ZN(n6990) );
  NAND2_X1 U8657 ( .A1(n7015), .A2(n11822), .ZN(n13552) );
  AND2_X1 U8658 ( .A1(n10909), .A2(n10906), .ZN(n10907) );
  NOR2_X1 U8659 ( .A1(n7011), .A2(n7010), .ZN(n7009) );
  NAND2_X1 U8660 ( .A1(n7023), .A2(n7021), .ZN(n7018) );
  NAND2_X1 U8661 ( .A1(n7017), .A2(n7021), .ZN(n7016) );
  INV_X1 U8662 ( .A(n13571), .ZN(n7021) );
  INV_X1 U8663 ( .A(n7022), .ZN(n13570) );
  OAI21_X1 U8664 ( .B1(n13499), .B2(n7020), .A(n7019), .ZN(n7022) );
  NAND2_X1 U8665 ( .A1(n6993), .A2(n9586), .ZN(n6995) );
  AND2_X1 U8666 ( .A1(n6995), .A2(n6989), .ZN(n9650) );
  INV_X1 U8667 ( .A(n9651), .ZN(n6989) );
  AND2_X1 U8668 ( .A1(n9867), .A2(n9868), .ZN(n6665) );
  XNOR2_X1 U8669 ( .A(n7024), .B(n11785), .ZN(n13638) );
  NAND2_X1 U8670 ( .A1(n13499), .A2(n11781), .ZN(n7024) );
  OR3_X1 U8671 ( .A1(n11498), .A2(n11497), .A3(n11496), .ZN(n13814) );
  NAND4_X1 U8672 ( .A1(n11456), .A2(n11455), .A3(n11454), .A4(n11453), .ZN(
        n13847) );
  AND2_X1 U8673 ( .A1(n11522), .A2(n11521), .ZN(n14027) );
  NAND2_X1 U8674 ( .A1(n7332), .A2(n7330), .ZN(n13859) );
  NAND2_X1 U8675 ( .A1(n13884), .A2(n11899), .ZN(n13858) );
  NAND2_X1 U8676 ( .A1(n13919), .A2(n11918), .ZN(n13904) );
  NAND2_X1 U8677 ( .A1(n13933), .A2(n13934), .ZN(n7068) );
  NAND2_X1 U8678 ( .A1(n13948), .A2(n11913), .ZN(n13929) );
  NAND2_X1 U8679 ( .A1(n7058), .A2(n11895), .ZN(n13961) );
  NAND2_X1 U8680 ( .A1(n11091), .A2(n11090), .ZN(n14409) );
  NAND2_X1 U8681 ( .A1(n10970), .A2(n11547), .ZN(n10973) );
  NAND2_X1 U8682 ( .A1(n7029), .A2(n10764), .ZN(n10969) );
  NAND2_X1 U8683 ( .A1(n10763), .A2(n10762), .ZN(n7029) );
  NAND2_X1 U8684 ( .A1(n10769), .A2(n11592), .ZN(n7315) );
  NAND2_X1 U8685 ( .A1(n10614), .A2(n10613), .ZN(n10681) );
  OAI21_X1 U8686 ( .B1(n10285), .B2(n7038), .A(n7036), .ZN(n10374) );
  NAND2_X1 U8687 ( .A1(n9936), .A2(n9935), .ZN(n10193) );
  NAND2_X1 U8688 ( .A1(n13893), .A2(n9944), .ZN(n14534) );
  INV_X1 U8689 ( .A(n14555), .ZN(n10164) );
  INV_X1 U8690 ( .A(n14534), .ZN(n14398) );
  NOR2_X1 U8691 ( .A1(n14531), .A2(n11539), .ZN(n14520) );
  INV_X1 U8692 ( .A(n13989), .ZN(n14519) );
  AND2_X2 U8693 ( .A1(n9687), .A2(n9686), .ZN(n14630) );
  INV_X1 U8694 ( .A(n6742), .ZN(n6626) );
  NAND2_X1 U8695 ( .A1(n14036), .A2(n6654), .ZN(n14098) );
  AND2_X1 U8696 ( .A1(n14035), .A2(n14034), .ZN(n6654) );
  NAND2_X1 U8697 ( .A1(n11542), .A2(n11489), .ZN(n14118) );
  NAND2_X1 U8698 ( .A1(n7433), .A2(n7431), .ZN(n11542) );
  NAND2_X1 U8699 ( .A1(n7433), .A2(n11485), .ZN(n11487) );
  NAND2_X1 U8700 ( .A1(n8727), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8724) );
  NAND2_X1 U8701 ( .A1(n7407), .A2(n11166), .ZN(n11082) );
  XNOR2_X1 U8702 ( .A(n11363), .B(P2_DATAO_REG_22__SCAN_IN), .ZN(n14132) );
  INV_X1 U8703 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n8786) );
  AND2_X1 U8704 ( .A1(n8660), .A2(n8649), .ZN(n13769) );
  INV_X1 U8705 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n8605) );
  INV_X1 U8706 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n8584) );
  INV_X1 U8707 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n8592) );
  NAND2_X1 U8708 ( .A1(n15252), .A2(n15253), .ZN(n14179) );
  NAND2_X1 U8709 ( .A1(n15251), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n14186) );
  XNOR2_X1 U8710 ( .A(n14194), .B(n6867), .ZN(n14254) );
  INV_X1 U8711 ( .A(P2_ADDR_REG_6__SCAN_IN), .ZN(n6867) );
  XNOR2_X1 U8712 ( .A(n14207), .B(n6865), .ZN(n14256) );
  INV_X1 U8713 ( .A(n14206), .ZN(n6865) );
  AND2_X1 U8714 ( .A1(n6638), .A2(n6639), .ZN(n14473) );
  NOR2_X1 U8715 ( .A1(n14473), .A2(n14472), .ZN(n14471) );
  INV_X1 U8716 ( .A(n7348), .ZN(n14854) );
  INV_X1 U8717 ( .A(n7358), .ZN(n12232) );
  OAI21_X1 U8718 ( .B1(n12264), .B2(n14893), .A(n6542), .ZN(P3_U3200) );
  AND2_X1 U8719 ( .A1(n7358), .A2(n7357), .ZN(n12252) );
  AND2_X1 U8720 ( .A1(n12282), .A2(n10361), .ZN(n8399) );
  OAI21_X1 U8721 ( .B1(n11992), .B2(n8422), .A(n8427), .ZN(P3_U3456) );
  OAI21_X1 U8722 ( .B1(n12275), .B2(n12583), .A(n8425), .ZN(n8426) );
  AOI21_X1 U8723 ( .B1(n11163), .B2(n15015), .A(n7397), .ZN(n11165) );
  NAND2_X1 U8724 ( .A1(n7400), .A2(n7398), .ZN(n7397) );
  OR2_X1 U8725 ( .A1(n15015), .A2(n7399), .ZN(n7398) );
  MUX2_X1 U8726 ( .A(n12539), .B(n12538), .S(n15015), .Z(n12540) );
  NAND2_X1 U8727 ( .A1(n9698), .A2(n9476), .ZN(n9708) );
  INV_X1 U8728 ( .A(n6642), .ZN(n6641) );
  OAI21_X1 U8729 ( .B1(n13345), .B2(n12719), .A(n12718), .ZN(n6642) );
  AOI21_X1 U8730 ( .B1(n13156), .B2(n14692), .A(n6633), .ZN(n13157) );
  NAND2_X1 U8731 ( .A1(n6702), .A2(n6605), .ZN(P2_U3495) );
  NAND2_X1 U8732 ( .A1(n13411), .A2(n14797), .ZN(n6702) );
  INV_X1 U8733 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6701) );
  AND2_X1 U8734 ( .A1(n13498), .A2(n6621), .ZN(n6620) );
  NAND2_X1 U8735 ( .A1(n14038), .A2(n13647), .ZN(n6621) );
  INV_X1 U8736 ( .A(n6993), .ZN(n9643) );
  OR2_X1 U8737 ( .A1(n11615), .A2(n11614), .ZN(n6660) );
  NAND2_X1 U8738 ( .A1(n6741), .A2(n6739), .ZN(P1_U3557) );
  OR2_X1 U8739 ( .A1(n14630), .A2(n6740), .ZN(n6739) );
  NAND2_X1 U8740 ( .A1(n14097), .A2(n14630), .ZN(n6741) );
  INV_X1 U8741 ( .A(P1_REG1_REG_29__SCAN_IN), .ZN(n6740) );
  NOR2_X1 U8742 ( .A1(n14459), .A2(n14458), .ZN(n14457) );
  AND2_X1 U8743 ( .A1(n6873), .A2(n6872), .ZN(n14459) );
  NOR2_X1 U8744 ( .A1(n15041), .A2(n15040), .ZN(n15243) );
  AND2_X1 U8745 ( .A1(n7253), .A2(n7252), .ZN(n6489) );
  INV_X1 U8746 ( .A(n12873), .ZN(n6859) );
  INV_X1 U8747 ( .A(n9620), .ZN(n9846) );
  AND2_X2 U8748 ( .A1(n11364), .A2(n11361), .ZN(n9599) );
  NAND2_X1 U8749 ( .A1(n10873), .A2(n10872), .ZN(n6491) );
  AND2_X1 U8750 ( .A1(n13846), .A2(n7047), .ZN(n6492) );
  NAND2_X1 U8751 ( .A1(n7367), .A2(n7557), .ZN(n7585) );
  INV_X2 U8752 ( .A(n7585), .ZN(n7556) );
  INV_X1 U8753 ( .A(n13934), .ZN(n7067) );
  AND2_X1 U8754 ( .A1(n14056), .A2(n13873), .ZN(n6493) );
  NAND2_X1 U8755 ( .A1(n11641), .A2(n11640), .ZN(n13380) );
  INV_X1 U8756 ( .A(n13885), .ZN(n7328) );
  AND3_X1 U8757 ( .A1(n6901), .A2(n6766), .A3(n6900), .ZN(n7697) );
  NAND2_X1 U8758 ( .A1(n14132), .A2(n11364), .ZN(n11572) );
  INV_X1 U8759 ( .A(n11572), .ZN(n6886) );
  AND2_X1 U8760 ( .A1(n11785), .A2(n13637), .ZN(n6494) );
  NOR3_X1 U8761 ( .A1(n12379), .A2(n12398), .A3(n8220), .ZN(n6495) );
  NAND2_X1 U8762 ( .A1(n11937), .A2(n11936), .ZN(n6496) );
  NAND2_X1 U8763 ( .A1(n11119), .A2(n11118), .ZN(n12873) );
  AND2_X1 U8764 ( .A1(n7183), .A2(n6545), .ZN(n6497) );
  INV_X1 U8765 ( .A(n8247), .ZN(n7570) );
  OR2_X1 U8766 ( .A1(n10658), .A2(n10660), .ZN(n6498) );
  AND2_X1 U8767 ( .A1(n12899), .A2(n6580), .ZN(n6499) );
  OR2_X1 U8768 ( .A1(n9853), .A2(n7312), .ZN(n6500) );
  NAND2_X1 U8769 ( .A1(n7255), .A2(n7254), .ZN(n6501) );
  NOR2_X1 U8770 ( .A1(n12392), .A2(n11944), .ZN(n6502) );
  NAND2_X1 U8771 ( .A1(n11523), .A2(n6582), .ZN(n6503) );
  AND2_X1 U8772 ( .A1(n6721), .A2(n6718), .ZN(n6504) );
  AND2_X1 U8773 ( .A1(n7504), .A2(n7292), .ZN(n6505) );
  AND2_X1 U8774 ( .A1(n6505), .A2(P1_DATAO_REG_13__SCAN_IN), .ZN(n6506) );
  NAND2_X1 U8775 ( .A1(n11461), .A2(n11460), .ZN(n14038) );
  AND2_X1 U8776 ( .A1(n7474), .A2(n10998), .ZN(n6507) );
  INV_X1 U8777 ( .A(n7861), .ZN(n6814) );
  AND2_X1 U8778 ( .A1(n7992), .A2(n7991), .ZN(n8787) );
  INV_X1 U8779 ( .A(n14545), .ZN(n7146) );
  AND2_X2 U8780 ( .A1(n9549), .A2(n9548), .ZN(n6508) );
  INV_X1 U8781 ( .A(n12976), .ZN(n12932) );
  INV_X1 U8782 ( .A(P3_IR_REG_4__SCAN_IN), .ZN(n7607) );
  NAND2_X1 U8783 ( .A1(n13267), .A2(n7199), .ZN(n7202) );
  NAND2_X1 U8784 ( .A1(n8247), .A2(n7524), .ZN(n7608) );
  NOR2_X1 U8785 ( .A1(n8086), .A2(n8085), .ZN(n8207) );
  AND2_X1 U8786 ( .A1(n14289), .A2(n14291), .ZN(n6509) );
  AND2_X1 U8787 ( .A1(n8247), .A2(n6769), .ZN(n6766) );
  INV_X1 U8788 ( .A(n11910), .ZN(n7120) );
  NAND2_X1 U8789 ( .A1(n7986), .A2(n7394), .ZN(n6510) );
  INV_X1 U8790 ( .A(n11233), .ZN(n6874) );
  NAND2_X1 U8791 ( .A1(n7986), .A2(n7533), .ZN(n6511) );
  OR2_X1 U8792 ( .A1(n14072), .A2(n13917), .ZN(n6512) );
  AND2_X2 U8793 ( .A1(n12595), .A2(n12015), .ZN(n6513) );
  INV_X1 U8794 ( .A(n8058), .ZN(n8039) );
  NOR2_X1 U8795 ( .A1(n11298), .A2(n11551), .ZN(n6514) );
  AND2_X1 U8796 ( .A1(n12866), .A2(n12865), .ZN(n6515) );
  XNOR2_X1 U8797 ( .A(n13327), .B(n11865), .ZN(n13022) );
  AND2_X1 U8798 ( .A1(n12847), .A2(n12846), .ZN(n6516) );
  INV_X1 U8799 ( .A(n8441), .ZN(n8909) );
  OAI21_X1 U8800 ( .B1(n8410), .B2(n14949), .A(n8409), .ZN(n12272) );
  AND2_X1 U8801 ( .A1(n12796), .A2(n12795), .ZN(n6517) );
  NOR2_X1 U8802 ( .A1(n13969), .A2(n13978), .ZN(n6518) );
  AND2_X1 U8803 ( .A1(n13299), .A2(n6861), .ZN(n6519) );
  OAI21_X1 U8804 ( .B1(n12078), .B2(n6905), .A(n6902), .ZN(n6907) );
  AND4_X1 U8805 ( .A1(n7629), .A2(n7628), .A3(n7627), .A4(n7626), .ZN(n7638)
         );
  INV_X1 U8806 ( .A(n9599), .ZN(n11490) );
  INV_X1 U8807 ( .A(n11973), .ZN(n7281) );
  INV_X1 U8808 ( .A(n7052), .ZN(n7051) );
  NOR2_X1 U8809 ( .A1(n13873), .A2(n13887), .ZN(n7052) );
  NAND2_X1 U8810 ( .A1(n11712), .A2(n11711), .ZN(n6521) );
  OR2_X1 U8811 ( .A1(n10192), .A2(n14561), .ZN(n6522) );
  AND2_X1 U8812 ( .A1(n7218), .A2(n11883), .ZN(n6523) );
  NOR2_X1 U8813 ( .A1(n12922), .A2(n13042), .ZN(n6524) );
  INV_X1 U8814 ( .A(P3_ADDR_REG_2__SCAN_IN), .ZN(n14139) );
  INV_X1 U8815 ( .A(n12975), .ZN(n6858) );
  NAND2_X1 U8816 ( .A1(n12946), .A2(n12945), .ZN(n12975) );
  XNOR2_X1 U8817 ( .A(n11570), .B(n11569), .ZN(n11998) );
  INV_X1 U8818 ( .A(n8213), .ZN(n10806) );
  NAND2_X1 U8819 ( .A1(n11423), .A2(n11422), .ZN(n14049) );
  NAND2_X1 U8820 ( .A1(n11432), .A2(n11431), .ZN(n14043) );
  INV_X1 U8821 ( .A(n11574), .ZN(n13962) );
  INV_X1 U8822 ( .A(n8144), .ZN(n7155) );
  INV_X1 U8823 ( .A(n13253), .ZN(n12988) );
  AND2_X1 U8824 ( .A1(n12754), .A2(n9156), .ZN(n6525) );
  AND2_X1 U8825 ( .A1(n13231), .A2(n7201), .ZN(n6526) );
  OR3_X1 U8826 ( .A1(P3_IR_REG_2__SCAN_IN), .A2(P3_IR_REG_1__SCAN_IN), .A3(
        P3_IR_REG_0__SCAN_IN), .ZN(n6527) );
  INV_X1 U8827 ( .A(n14898), .ZN(n6794) );
  AND3_X1 U8828 ( .A1(n6766), .A2(n7479), .A3(n6901), .ZN(n6528) );
  NAND2_X1 U8829 ( .A1(n11634), .A2(n11635), .ZN(n6529) );
  AND2_X1 U8830 ( .A1(n12791), .A2(n13061), .ZN(n6530) );
  NOR2_X1 U8831 ( .A1(n7262), .A2(n12609), .ZN(n7261) );
  AND2_X1 U8832 ( .A1(n7413), .A2(n7412), .ZN(n6531) );
  INV_X1 U8833 ( .A(n13161), .ZN(n13324) );
  OAI21_X1 U8834 ( .B1(n14118), .B2(n12931), .A(n12930), .ZN(n13161) );
  AND2_X1 U8835 ( .A1(n10072), .A2(n10039), .ZN(n6532) );
  AND2_X1 U8836 ( .A1(n11859), .A2(n11858), .ZN(n13173) );
  INV_X1 U8837 ( .A(n13173), .ZN(n7215) );
  AND2_X1 U8838 ( .A1(n9730), .A2(n9729), .ZN(n6533) );
  NAND2_X1 U8839 ( .A1(n11739), .A2(n11738), .ZN(n13331) );
  AND2_X1 U8840 ( .A1(n6894), .A2(n6892), .ZN(n6534) );
  NOR2_X1 U8841 ( .A1(n12197), .A2(n8271), .ZN(n6535) );
  AND2_X1 U8842 ( .A1(n7267), .A2(n6521), .ZN(n6536) );
  INV_X1 U8843 ( .A(n12885), .ZN(n13374) );
  NAND2_X1 U8844 ( .A1(n11648), .A2(n11647), .ZN(n12885) );
  AND2_X1 U8845 ( .A1(n11972), .A2(n11973), .ZN(n6537) );
  AND2_X1 U8846 ( .A1(n14789), .A2(n13058), .ZN(n6538) );
  AND2_X1 U8847 ( .A1(n9553), .A2(n9716), .ZN(n6539) );
  AND2_X1 U8848 ( .A1(n11621), .A2(n11622), .ZN(n6540) );
  AND2_X1 U8849 ( .A1(n12333), .A2(n8188), .ZN(n6541) );
  AND3_X1 U8850 ( .A1(n6983), .A2(n12257), .A3(n6655), .ZN(n6542) );
  INV_X1 U8851 ( .A(n6796), .ZN(n6795) );
  AND2_X1 U8852 ( .A1(n11560), .A2(n6647), .ZN(n6543) );
  AND2_X1 U8853 ( .A1(n7064), .A2(n7065), .ZN(n6544) );
  NAND2_X1 U8854 ( .A1(n12810), .A2(n13057), .ZN(n6545) );
  NAND2_X1 U8855 ( .A1(n13905), .A2(n6878), .ZN(n6880) );
  AND2_X1 U8856 ( .A1(n8674), .A2(n8671), .ZN(n6546) );
  INV_X1 U8857 ( .A(n8960), .ZN(n6727) );
  AND2_X1 U8858 ( .A1(n14043), .A2(n13866), .ZN(n6547) );
  NAND2_X1 U8859 ( .A1(n10871), .A2(n12130), .ZN(n6548) );
  AND2_X1 U8860 ( .A1(n8125), .A2(n8126), .ZN(n10632) );
  INV_X1 U8861 ( .A(n7380), .ZN(n12311) );
  AOI21_X1 U8862 ( .B1(n12351), .B2(n7383), .A(n7381), .ZN(n7380) );
  AND2_X1 U8863 ( .A1(n6937), .A2(n6935), .ZN(n6549) );
  NAND4_X1 U8864 ( .A1(n7567), .A2(n7566), .A3(n7565), .A4(n7564), .ZN(n12142)
         );
  INV_X1 U8865 ( .A(n12142), .ZN(n6807) );
  AND2_X1 U8866 ( .A1(n7535), .A2(n7181), .ZN(n6550) );
  INV_X1 U8867 ( .A(n7385), .ZN(n7384) );
  OAI21_X1 U8868 ( .B1(n7386), .B2(n7881), .A(n7893), .ZN(n7385) );
  INV_X1 U8869 ( .A(n7473), .ZN(n7243) );
  NOR2_X1 U8870 ( .A1(n14432), .A2(n14394), .ZN(n6551) );
  NOR2_X1 U8871 ( .A1(n14579), .A2(n10376), .ZN(n6552) );
  NOR2_X1 U8872 ( .A1(n14432), .A2(n11283), .ZN(n6553) );
  NOR2_X1 U8873 ( .A1(n12951), .A2(n12950), .ZN(n6554) );
  AND2_X1 U8874 ( .A1(n7278), .A2(n8205), .ZN(n6555) );
  NAND2_X1 U8875 ( .A1(n14342), .A2(n13054), .ZN(n6556) );
  INV_X1 U8876 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n14111) );
  AND2_X1 U8877 ( .A1(n13374), .A2(n12692), .ZN(n6557) );
  AND2_X1 U8878 ( .A1(n14062), .A2(n13918), .ZN(n6558) );
  AND2_X1 U8879 ( .A1(n12873), .A2(n13049), .ZN(n6559) );
  INV_X1 U8880 ( .A(n11975), .ZN(n6899) );
  AND2_X1 U8881 ( .A1(n7440), .A2(n12757), .ZN(n6560) );
  AND2_X1 U8882 ( .A1(n12902), .A2(n12903), .ZN(n6561) );
  INV_X1 U8883 ( .A(n12913), .ZN(n7468) );
  INV_X1 U8884 ( .A(n8101), .ZN(n10278) );
  OR2_X1 U8885 ( .A1(n6516), .A2(n7453), .ZN(n6562) );
  INV_X1 U8886 ( .A(n6879), .ZN(n6878) );
  NAND2_X1 U8887 ( .A1(n6493), .A2(n13854), .ZN(n6879) );
  INV_X1 U8888 ( .A(n6883), .ZN(n6882) );
  NAND2_X1 U8889 ( .A1(n6885), .A2(n6884), .ZN(n6883) );
  OR2_X1 U8890 ( .A1(n7271), .A2(n12654), .ZN(n6563) );
  NOR2_X1 U8891 ( .A1(n13873), .A2(n13630), .ZN(n6564) );
  AND2_X1 U8892 ( .A1(n8542), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n6565) );
  INV_X1 U8893 ( .A(n6905), .ZN(n6904) );
  OR2_X1 U8894 ( .A1(n12041), .A2(n6906), .ZN(n6905) );
  INV_X1 U8895 ( .A(n7039), .ZN(n7038) );
  NOR2_X1 U8896 ( .A1(n10223), .A2(n7040), .ZN(n7039) );
  OR2_X1 U8897 ( .A1(n9350), .A2(n9237), .ZN(n6566) );
  NAND2_X1 U8898 ( .A1(n10666), .A2(n10667), .ZN(n6567) );
  NAND2_X1 U8899 ( .A1(n11328), .A2(n11327), .ZN(n6568) );
  AND2_X1 U8900 ( .A1(n11952), .A2(n11953), .ZN(n6569) );
  AND2_X1 U8901 ( .A1(n6516), .A2(n7453), .ZN(n6570) );
  AND2_X1 U8902 ( .A1(n11735), .A2(n7268), .ZN(n6571) );
  INV_X1 U8903 ( .A(n7023), .ZN(n7020) );
  OR2_X1 U8904 ( .A1(n11785), .A2(n13637), .ZN(n7023) );
  INV_X1 U8905 ( .A(n10887), .ZN(n7011) );
  INV_X1 U8906 ( .A(n12899), .ZN(n6751) );
  NAND2_X1 U8907 ( .A1(n11916), .A2(n6512), .ZN(n6572) );
  NAND2_X1 U8908 ( .A1(n13186), .A2(n7217), .ZN(n6573) );
  NAND2_X1 U8909 ( .A1(n12399), .A2(n7831), .ZN(n12386) );
  INV_X1 U8910 ( .A(n11444), .ZN(n7135) );
  AND2_X1 U8911 ( .A1(n7068), .A2(n6512), .ZN(n6574) );
  OR2_X1 U8912 ( .A1(n12455), .A2(n12439), .ZN(n8147) );
  AND2_X1 U8913 ( .A1(n7211), .A2(n13022), .ZN(n6575) );
  OR2_X1 U8914 ( .A1(n11250), .A2(n10224), .ZN(n6576) );
  INV_X1 U8915 ( .A(n11587), .ZN(n10619) );
  OR2_X1 U8916 ( .A1(n14205), .A2(n14204), .ZN(n6577) );
  OR2_X1 U8917 ( .A1(n14215), .A2(n14216), .ZN(n6578) );
  AND2_X1 U8918 ( .A1(n6855), .A2(n12975), .ZN(n6579) );
  AND2_X1 U8919 ( .A1(n12896), .A2(n12895), .ZN(n6580) );
  AND2_X1 U8920 ( .A1(n7013), .A2(n7012), .ZN(n6581) );
  OR2_X1 U8921 ( .A1(n11524), .A2(n11525), .ZN(n6582) );
  AND2_X1 U8922 ( .A1(n6899), .A2(n6896), .ZN(n6583) );
  AND2_X1 U8923 ( .A1(n6913), .A2(n6491), .ZN(n6584) );
  AND2_X1 U8924 ( .A1(n11829), .A2(n11822), .ZN(n6585) );
  OR2_X1 U8925 ( .A1(n11249), .A2(n11247), .ZN(n6586) );
  AND2_X1 U8926 ( .A1(n8189), .A2(n12295), .ZN(n12326) );
  AOI21_X1 U8927 ( .B1(n7419), .B2(n7421), .A(n6566), .ZN(n7417) );
  AND2_X1 U8928 ( .A1(n12970), .A2(n7424), .ZN(n6587) );
  AND2_X1 U8929 ( .A1(n7340), .A2(n8771), .ZN(n6588) );
  NAND2_X1 U8930 ( .A1(n8620), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n6589) );
  AND2_X1 U8931 ( .A1(n12829), .A2(n12828), .ZN(n6590) );
  AND2_X1 U8932 ( .A1(n12629), .A2(n6529), .ZN(n7247) );
  AND2_X1 U8933 ( .A1(n8723), .A2(n7077), .ZN(n7340) );
  INV_X1 U8934 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n9273) );
  INV_X1 U8935 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n7077) );
  INV_X1 U8936 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n8674) );
  INV_X1 U8937 ( .A(n13358), .ZN(n13236) );
  NAND2_X1 U8938 ( .A1(n11687), .A2(n11686), .ZN(n13358) );
  INV_X1 U8939 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n9269) );
  INV_X1 U8940 ( .A(P3_IR_REG_2__SCAN_IN), .ZN(n7593) );
  INV_X1 U8941 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n7012) );
  INV_X1 U8942 ( .A(n7266), .ZN(n7265) );
  INV_X1 U8943 ( .A(n12443), .ZN(n7149) );
  OR2_X2 U8944 ( .A1(n14382), .A2(n14391), .ZN(n7474) );
  INV_X1 U8945 ( .A(n7617), .ZN(n7284) );
  XNOR2_X1 U8946 ( .A(n14062), .B(n13918), .ZN(n13903) );
  INV_X1 U8947 ( .A(n13903), .ZN(n7063) );
  INV_X1 U8948 ( .A(n10341), .ZN(n6680) );
  AND2_X1 U8949 ( .A1(n13983), .A2(n6882), .ZN(n6591) );
  INV_X1 U8950 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6732) );
  OR2_X1 U8951 ( .A1(n9933), .A2(SI_18_), .ZN(n6592) );
  NOR2_X1 U8952 ( .A1(n13313), .A2(n13390), .ZN(n6860) );
  INV_X1 U8953 ( .A(n12464), .ZN(n6840) );
  AND2_X1 U8954 ( .A1(n7311), .A2(n8581), .ZN(n9247) );
  NAND2_X1 U8955 ( .A1(n7747), .A2(n7746), .ZN(n12465) );
  NAND2_X1 U8956 ( .A1(n7790), .A2(n7789), .ZN(n12425) );
  XNOR2_X1 U8957 ( .A(n7274), .B(n11621), .ZN(n11623) );
  NAND2_X1 U8958 ( .A1(n7370), .A2(n7372), .ZN(n10921) );
  NAND2_X1 U8959 ( .A1(n11098), .A2(n11097), .ZN(n11906) );
  NAND2_X1 U8960 ( .A1(n6691), .A2(n7183), .ZN(n10140) );
  NAND2_X1 U8961 ( .A1(n7185), .A2(n10041), .ZN(n10073) );
  NAND2_X1 U8962 ( .A1(n7315), .A2(n10770), .ZN(n10997) );
  INV_X1 U8963 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n8973) );
  INV_X1 U8964 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n7296) );
  AND2_X1 U8965 ( .A1(n8624), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n6593) );
  INV_X1 U8966 ( .A(n11277), .ZN(n7130) );
  NOR2_X1 U8967 ( .A1(n12579), .A2(n11936), .ZN(n6594) );
  NOR2_X1 U8968 ( .A1(n14879), .A2(n8305), .ZN(n6595) );
  NOR2_X1 U8969 ( .A1(n12162), .A2(n8307), .ZN(n6596) );
  AND2_X1 U8970 ( .A1(n6970), .A2(n11138), .ZN(n6597) );
  AND2_X1 U8971 ( .A1(n12076), .A2(n6904), .ZN(n6598) );
  NOR2_X1 U8972 ( .A1(n12455), .A2(n11930), .ZN(n6599) );
  AND2_X1 U8973 ( .A1(n10530), .A2(n15045), .ZN(n6600) );
  NOR2_X1 U8974 ( .A1(n8974), .A2(n7470), .ZN(n9243) );
  AND2_X1 U8975 ( .A1(n12133), .A2(n15017), .ZN(n6601) );
  NOR2_X1 U8976 ( .A1(n14346), .A2(n14342), .ZN(n10745) );
  AND2_X1 U8977 ( .A1(n7501), .A2(P1_DATAO_REG_10__SCAN_IN), .ZN(n6602) );
  INV_X1 U8978 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n9215) );
  INV_X1 U8979 ( .A(n12402), .ZN(n12398) );
  INV_X1 U8980 ( .A(P3_IR_REG_21__SCAN_IN), .ZN(n7931) );
  INV_X1 U8981 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n8665) );
  NOR2_X1 U8982 ( .A1(n7794), .A2(P3_IR_REG_16__SCAN_IN), .ZN(n6603) );
  NOR2_X1 U8983 ( .A1(n9978), .A2(n14969), .ZN(n6604) );
  NAND2_X2 U8984 ( .A1(n8927), .A2(n12720), .ZN(n9329) );
  NAND2_X1 U8985 ( .A1(n9283), .A2(n14532), .ZN(n13647) );
  INV_X1 U8986 ( .A(n14887), .ZN(n6984) );
  NAND2_X1 U8987 ( .A1(n10519), .A2(n10518), .ZN(n10662) );
  OR2_X1 U8988 ( .A1(n14797), .A2(n6701), .ZN(n6605) );
  NAND2_X1 U8989 ( .A1(n6692), .A2(n10139), .ZN(n10253) );
  NAND2_X1 U8990 ( .A1(n7160), .A2(n7158), .ZN(n10804) );
  OAI21_X1 U8991 ( .B1(n6696), .B2(n6695), .A(n6693), .ZN(n9802) );
  NAND2_X1 U8992 ( .A1(n9804), .A2(n9803), .ZN(n10040) );
  NAND2_X1 U8993 ( .A1(n14911), .A2(n8121), .ZN(n10631) );
  INV_X1 U8994 ( .A(n6697), .ZN(n9765) );
  NAND2_X1 U8995 ( .A1(n11352), .A2(n11351), .ZN(n14072) );
  INV_X1 U8996 ( .A(n14072), .ZN(n6884) );
  AND2_X1 U8997 ( .A1(n14846), .A2(n12263), .ZN(n6606) );
  OR2_X1 U8998 ( .A1(n9740), .A2(n9739), .ZN(n9923) );
  INV_X1 U8999 ( .A(n9923), .ZN(n7251) );
  AND2_X1 U9000 ( .A1(n7169), .A2(n8131), .ZN(n6607) );
  AND2_X1 U9001 ( .A1(n7511), .A2(n10557), .ZN(n6608) );
  AND2_X1 U9002 ( .A1(n10967), .A2(P2_DATAO_REG_22__SCAN_IN), .ZN(n6609) );
  AND2_X1 U9003 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n9370), .ZN(n6610) );
  INV_X1 U9004 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n9358) );
  AND2_X1 U9005 ( .A1(n6815), .A2(n7514), .ZN(n6611) );
  NAND2_X1 U9006 ( .A1(n8932), .A2(n13253), .ZN(n9328) );
  NAND2_X1 U9007 ( .A1(n7538), .A2(n7549), .ZN(n7945) );
  XNOR2_X1 U9008 ( .A(n8724), .B(n8771), .ZN(n8743) );
  INV_X1 U9009 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n6834) );
  XNOR2_X1 U9010 ( .A(n9270), .B(n9269), .ZN(n11206) );
  INV_X1 U9011 ( .A(n11206), .ZN(n7147) );
  AND2_X1 U9012 ( .A1(n9693), .A2(n7243), .ZN(n7241) );
  XNOR2_X1 U9013 ( .A(n8250), .B(n9072), .ZN(n9063) );
  NAND2_X1 U9014 ( .A1(n6690), .A2(n9138), .ZN(n14711) );
  NAND2_X1 U9015 ( .A1(n10061), .A2(n10060), .ZN(n12810) );
  INV_X1 U9016 ( .A(n12810), .ZN(n6847) );
  INV_X1 U9017 ( .A(n14789), .ZN(n6849) );
  NOR2_X1 U9018 ( .A1(n9066), .A2(n8289), .ZN(n6612) );
  NOR2_X1 U9019 ( .A1(n9062), .A2(n8251), .ZN(n6613) );
  OR2_X1 U9020 ( .A1(n10822), .A2(n10818), .ZN(n6614) );
  INV_X1 U9021 ( .A(n9459), .ZN(n9464) );
  AND2_X1 U9022 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n11180), .ZN(n6615) );
  AND2_X1 U9023 ( .A1(n6963), .A2(n6962), .ZN(n6616) );
  INV_X1 U9024 ( .A(SI_22_), .ZN(n6673) );
  INV_X1 U9025 ( .A(n12263), .ZN(n9134) );
  INV_X1 U9026 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n7289) );
  INV_X1 U9027 ( .A(P1_ADDR_REG_0__SCAN_IN), .ZN(n6676) );
  INV_X1 U9028 ( .A(P3_ADDR_REG_5__SCAN_IN), .ZN(n6688) );
  INV_X1 U9029 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n7312) );
  NAND2_X1 U9030 ( .A1(n8734), .A2(n9252), .ZN(n9663) );
  NAND2_X1 U9031 ( .A1(n13612), .A2(n13613), .ZN(n13611) );
  NAND2_X1 U9032 ( .A1(n11841), .A2(n11840), .ZN(n13451) );
  NAND2_X1 U9033 ( .A1(n11052), .A2(n11051), .ZN(n11772) );
  NAND2_X1 U9034 ( .A1(n6622), .A2(n6620), .ZN(P1_U3214) );
  NAND2_X1 U9035 ( .A1(n10426), .A2(n10425), .ZN(n10791) );
  NOR2_X2 U9036 ( .A1(n9294), .A2(n9575), .ZN(n9574) );
  NAND2_X1 U9037 ( .A1(n13494), .A2(n13626), .ZN(n6622) );
  INV_X1 U9038 ( .A(n9645), .ZN(n6988) );
  NAND2_X1 U9039 ( .A1(n13565), .A2(n13480), .ZN(n13624) );
  NAND2_X1 U9040 ( .A1(n9866), .A2(n6665), .ZN(n10171) );
  NAND2_X1 U9041 ( .A1(n13602), .A2(n13601), .ZN(n7015) );
  INV_X1 U9042 ( .A(n7513), .ZN(n6810) );
  NAND2_X1 U9043 ( .A1(n7300), .A2(n8228), .ZN(n8237) );
  NAND2_X1 U9044 ( .A1(n6623), .A2(n7484), .ZN(n7592) );
  OAI21_X1 U9045 ( .B1(n7486), .B2(n7284), .A(n7282), .ZN(n7606) );
  OAI21_X1 U9046 ( .B1(n8198), .B2(n8197), .A(n6555), .ZN(n6771) );
  NAND2_X1 U9047 ( .A1(n7505), .A2(n7504), .ZN(n7287) );
  NAND2_X1 U9048 ( .A1(n7568), .A2(n7578), .ZN(n6623) );
  NAND2_X1 U9049 ( .A1(n6764), .A2(n7298), .ZN(n7777) );
  NAND2_X1 U9050 ( .A1(n7310), .A2(n7309), .ZN(n7308) );
  NAND2_X1 U9051 ( .A1(n7519), .A2(n7520), .ZN(n7905) );
  XNOR2_X1 U9052 ( .A(n8403), .B(n8207), .ZN(n8410) );
  NAND3_X1 U9053 ( .A1(n6624), .A2(n8382), .A3(n8381), .ZN(P3_U3201) );
  AOI21_X1 U9054 ( .B1(P3_REG2_REG_4__SCAN_IN), .B2(n9185), .A(n9178), .ZN(
        n8253) );
  NOR2_X1 U9055 ( .A1(n8273), .A2(n12247), .ZN(n8274) );
  NOR2_X1 U9056 ( .A1(n9050), .A2(n8249), .ZN(n8250) );
  NOR2_X1 U9057 ( .A1(n14837), .A2(n6593), .ZN(n8259) );
  NOR2_X1 U9058 ( .A1(n10331), .A2(n8260), .ZN(n14856) );
  NAND2_X1 U9059 ( .A1(n8251), .A2(n7362), .ZN(n7360) );
  AOI21_X2 U9060 ( .B1(n13843), .B2(n13842), .A(n6547), .ZN(n13824) );
  OAI21_X2 U9061 ( .B1(n13974), .B2(n11912), .A(n11911), .ZN(n13959) );
  NAND2_X1 U9062 ( .A1(n14175), .A2(n14176), .ZN(n14138) );
  NAND2_X1 U9063 ( .A1(n14473), .A2(n14472), .ZN(n14227) );
  AOI21_X2 U9064 ( .B1(n14238), .B2(n14237), .A(n14268), .ZN(n14244) );
  NAND2_X1 U9065 ( .A1(n14464), .A2(n14463), .ZN(n14462) );
  OAI21_X1 U9066 ( .B1(n14255), .B2(P2_ADDR_REG_8__SCAN_IN), .A(n6577), .ZN(
        n6635) );
  NAND2_X1 U9067 ( .A1(n6630), .A2(n11994), .ZN(P3_U3488) );
  NAND2_X1 U9068 ( .A1(n11993), .A2(n7469), .ZN(n6630) );
  INV_X1 U9069 ( .A(n12272), .ZN(n7173) );
  OR2_X1 U9070 ( .A1(n10660), .A2(n10659), .ZN(n10661) );
  NAND2_X1 U9071 ( .A1(n6869), .A2(n6871), .ZN(n14215) );
  INV_X1 U9072 ( .A(n6677), .ZN(n14464) );
  NAND2_X1 U9073 ( .A1(n14174), .A2(n14173), .ZN(n6664) );
  NOR2_X1 U9074 ( .A1(n14477), .A2(n14476), .ZN(n14232) );
  AND2_X1 U9075 ( .A1(n14244), .A2(n14245), .ZN(n15039) );
  NAND2_X1 U9076 ( .A1(n14220), .A2(n14221), .ZN(n6638) );
  INV_X1 U9077 ( .A(n14467), .ZN(n6639) );
  NAND2_X1 U9078 ( .A1(n6722), .A2(n6640), .ZN(n6661) );
  NAND2_X1 U9079 ( .A1(n6650), .A2(n8496), .ZN(n6640) );
  NAND2_X1 U9080 ( .A1(n9347), .A2(n9129), .ZN(n9349) );
  NAND2_X1 U9081 ( .A1(n6643), .A2(n6641), .ZN(P2_U3212) );
  NAND2_X1 U9082 ( .A1(n12709), .A2(n14328), .ZN(n6643) );
  NAND3_X1 U9083 ( .A1(n6645), .A2(n6644), .A3(n7126), .ZN(n7125) );
  NAND2_X1 U9084 ( .A1(n11467), .A2(n11466), .ZN(n6644) );
  NAND2_X1 U9085 ( .A1(n11463), .A2(n11462), .ZN(n6645) );
  NAND2_X1 U9086 ( .A1(n11610), .A2(n6649), .ZN(n6648) );
  NAND2_X1 U9087 ( .A1(n9128), .A2(n15089), .ZN(n9347) );
  AOI21_X1 U9088 ( .B1(n7100), .B2(n7098), .A(n7097), .ZN(n7096) );
  NAND2_X1 U9089 ( .A1(n7108), .A2(n7112), .ZN(n11355) );
  NAND2_X1 U9090 ( .A1(n7418), .A2(n9125), .ZN(n9232) );
  NAND2_X1 U9091 ( .A1(n11409), .A2(n11408), .ZN(n11425) );
  NAND2_X1 U9092 ( .A1(n11446), .A2(n11445), .ZN(n11464) );
  NAND2_X1 U9093 ( .A1(n7088), .A2(n7087), .ZN(n7086) );
  AOI21_X1 U9094 ( .B1(n11376), .B2(n11375), .A(n11374), .ZN(n6646) );
  AOI21_X1 U9095 ( .B1(n7137), .B2(n7136), .A(n7135), .ZN(n7134) );
  INV_X1 U9096 ( .A(P3_ADDR_REG_19__SCAN_IN), .ZN(n8378) );
  INV_X1 U9097 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n13811) );
  INV_X1 U9098 ( .A(n11404), .ZN(n11407) );
  NAND2_X1 U9099 ( .A1(n7084), .A2(n7086), .ZN(n11404) );
  NAND2_X1 U9100 ( .A1(n8489), .A2(n8631), .ZN(n8496) );
  XNOR2_X2 U9101 ( .A(n14397), .B(n13656), .ZN(n14391) );
  INV_X1 U9102 ( .A(n7096), .ZN(n7095) );
  NAND2_X1 U9103 ( .A1(n7313), .A2(n7314), .ZN(n14382) );
  NAND2_X1 U9104 ( .A1(n10455), .A2(n10454), .ZN(n10620) );
  NAND2_X1 U9105 ( .A1(n6651), .A2(n10194), .ZN(n10284) );
  NOR2_X1 U9106 ( .A1(n9306), .A2(n6671), .ZN(n6670) );
  NAND2_X1 U9107 ( .A1(n10297), .A2(n10298), .ZN(n6651) );
  NAND2_X1 U9108 ( .A1(n8348), .A2(n8349), .ZN(n12153) );
  NAND2_X1 U9109 ( .A1(n9897), .A2(n8336), .ZN(n14841) );
  INV_X1 U9110 ( .A(n7539), .ZN(n7536) );
  NOR2_X1 U9111 ( .A1(n12169), .A2(n12168), .ZN(n12185) );
  NAND2_X1 U9112 ( .A1(n7542), .A2(n7541), .ZN(n6841) );
  NOR2_X1 U9113 ( .A1(n14883), .A2(n14884), .ZN(n14882) );
  OAI21_X1 U9114 ( .B1(n11617), .B2(n11616), .A(n6660), .ZN(P1_U3242) );
  NAND2_X1 U9115 ( .A1(n7111), .A2(n7110), .ZN(n7109) );
  NAND3_X1 U9116 ( .A1(n6661), .A2(n8493), .A3(n8494), .ZN(n8527) );
  NAND2_X1 U9117 ( .A1(n8354), .A2(n8353), .ZN(n12168) );
  NAND2_X1 U9118 ( .A1(n9819), .A2(n9818), .ZN(n9820) );
  INV_X1 U9119 ( .A(n9820), .ZN(n6720) );
  NAND2_X1 U9120 ( .A1(n6767), .A2(n6765), .ZN(n7539) );
  NOR2_X1 U9121 ( .A1(n12201), .A2(n12202), .ZN(n12200) );
  NAND2_X1 U9122 ( .A1(n9402), .A2(n12996), .ZN(n6662) );
  NAND2_X1 U9123 ( .A1(n6663), .A2(n14188), .ZN(n14191) );
  NAND2_X1 U9124 ( .A1(n15245), .A2(n15244), .ZN(n6663) );
  OAI22_X2 U9125 ( .A1(n14335), .A2(n10729), .B1(n14362), .B2(n13054), .ZN(
        n10934) );
  NAND2_X1 U9126 ( .A1(n10244), .A2(n10243), .ZN(n6944) );
  NAND2_X1 U9127 ( .A1(n13328), .A2(n6675), .ZN(n13410) );
  OAI21_X1 U9128 ( .B1(n14461), .B2(P2_ADDR_REG_12__SCAN_IN), .A(n6578), .ZN(
        n6677) );
  NAND2_X1 U9129 ( .A1(n9187), .A2(n9186), .ZN(n9190) );
  NOR4_X2 U9130 ( .A1(n8223), .A2(n12352), .A3(n8222), .A4(n8221), .ZN(n8226)
         );
  NAND2_X1 U9131 ( .A1(n7777), .A2(n7775), .ZN(n7297) );
  NAND2_X1 U9132 ( .A1(n8233), .A2(n8232), .ZN(n8234) );
  INV_X1 U9133 ( .A(n7905), .ZN(n7310) );
  NAND2_X1 U9134 ( .A1(n7764), .A2(n7763), .ZN(n6764) );
  NAND2_X1 U9135 ( .A1(n7492), .A2(n7491), .ZN(n7647) );
  NAND2_X1 U9136 ( .A1(n7664), .A2(n7663), .ZN(n7496) );
  NAND2_X1 U9137 ( .A1(n7606), .A2(n7604), .ZN(n7489) );
  XNOR2_X1 U9138 ( .A(n8309), .B(n8310), .ZN(n12207) );
  OAI21_X1 U9139 ( .B1(n13569), .B2(n13582), .A(n13581), .ZN(n13580) );
  NOR2_X1 U9140 ( .A1(n12263), .A2(n12523), .ZN(n6666) );
  NAND2_X1 U9141 ( .A1(n13492), .A2(n13493), .ZN(n13534) );
  INV_X1 U9142 ( .A(n9644), .ZN(n6987) );
  XNOR2_X2 U9143 ( .A(n10838), .B(n10794), .ZN(n10797) );
  NAND2_X2 U9144 ( .A1(n13451), .A2(n13450), .ZN(n13509) );
  INV_X1 U9145 ( .A(n9935), .ZN(n7323) );
  NAND3_X1 U9146 ( .A1(n9672), .A2(n6522), .A3(n11219), .ZN(n7321) );
  INV_X1 U9147 ( .A(n11580), .ZN(n10298) );
  INV_X1 U9148 ( .A(n6478), .ZN(n6669) );
  NAND2_X1 U9149 ( .A1(n7092), .A2(n7091), .ZN(n7090) );
  OAI21_X1 U9150 ( .B1(n11425), .B2(n7137), .A(n6672), .ZN(n11445) );
  NAND3_X1 U9151 ( .A1(n6723), .A2(n7417), .A3(n6725), .ZN(n9239) );
  NOR2_X2 U9152 ( .A1(n14200), .A2(n14201), .ZN(n14205) );
  INV_X1 U9153 ( .A(n7346), .ZN(n8262) );
  NOR2_X1 U9154 ( .A1(n9220), .A2(n6681), .ZN(n9052) );
  AND2_X1 U9155 ( .A1(n8247), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n6681) );
  AOI21_X1 U9156 ( .B1(n8263), .B2(n7344), .A(n8265), .ZN(n7343) );
  XNOR2_X2 U9157 ( .A(n8772), .B(P1_IR_REG_30__SCAN_IN), .ZN(n8777) );
  NAND2_X1 U9158 ( .A1(n7339), .A2(n6588), .ZN(n7341) );
  NAND2_X1 U9159 ( .A1(n6682), .A2(n6984), .ZN(n8382) );
  XNOR2_X1 U9160 ( .A(n8315), .B(n6683), .ZN(n6682) );
  INV_X1 U9161 ( .A(n8366), .ZN(n6683) );
  NAND2_X1 U9162 ( .A1(n13878), .A2(n7330), .ZN(n7326) );
  NAND2_X1 U9163 ( .A1(n8562), .A2(n8561), .ZN(n8574) );
  NAND2_X1 U9164 ( .A1(n8289), .A2(n6959), .ZN(n6957) );
  AOI21_X1 U9165 ( .B1(P3_REG1_REG_2__SCAN_IN), .B2(n9058), .A(n9044), .ZN(
        n8288) );
  NAND2_X1 U9166 ( .A1(n14841), .A2(n14842), .ZN(n8340) );
  NOR2_X2 U9167 ( .A1(n12178), .A2(n8308), .ZN(n8309) );
  NAND2_X1 U9168 ( .A1(n8305), .A2(n6956), .ZN(n6954) );
  NOR2_X1 U9169 ( .A1(n8306), .A2(n8266), .ZN(n8307) );
  AOI21_X1 U9170 ( .B1(n8328), .B2(n8284), .A(n8286), .ZN(n8285) );
  NOR2_X1 U9171 ( .A1(n12206), .A2(n8311), .ZN(n12225) );
  NOR2_X1 U9172 ( .A1(n15039), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n15041) );
  AND2_X2 U9173 ( .A1(n6687), .A2(n6686), .ZN(n14477) );
  NAND2_X1 U9174 ( .A1(n14227), .A2(n14228), .ZN(n6686) );
  INV_X1 U9175 ( .A(n14471), .ZN(n6687) );
  XNOR2_X1 U9176 ( .A(n14205), .B(n14204), .ZN(n14255) );
  NAND2_X1 U9177 ( .A1(n14711), .A2(n14712), .ZN(n6689) );
  NAND2_X1 U9178 ( .A1(n9137), .A2(n9136), .ZN(n6690) );
  AOI21_X1 U9179 ( .B1(n6694), .B2(n6698), .A(n6530), .ZN(n6693) );
  AND2_X1 U9180 ( .A1(n13001), .A2(n6699), .ZN(n6694) );
  NAND2_X1 U9181 ( .A1(n6698), .A2(n13001), .ZN(n6695) );
  AND3_X4 U9182 ( .A1(n8436), .A2(n7182), .A3(n8885), .ZN(n8441) );
  XNOR2_X2 U9184 ( .A(n13067), .B(n9021), .ZN(n12995) );
  AND2_X2 U9185 ( .A1(n8891), .A2(n6706), .ZN(n9021) );
  INV_X1 U9186 ( .A(n6713), .ZN(n13286) );
  NAND2_X1 U9187 ( .A1(n8520), .A2(n7404), .ZN(n6714) );
  NAND2_X1 U9188 ( .A1(n6714), .A2(n7402), .ZN(n8562) );
  NAND2_X1 U9189 ( .A1(n8574), .A2(n8573), .ZN(n8578) );
  NAND2_X1 U9190 ( .A1(n9820), .A2(n6504), .ZN(n6715) );
  AND2_X1 U9191 ( .A1(n8497), .A2(n8618), .ZN(n6722) );
  NAND2_X1 U9192 ( .A1(n7411), .A2(n6724), .ZN(n6723) );
  NAND2_X1 U9193 ( .A1(n7411), .A2(n7409), .ZN(n8961) );
  INV_X1 U9194 ( .A(P2_RD_REG_SCAN_IN), .ZN(n6729) );
  AND2_X4 U9195 ( .A1(n6730), .A2(n6728), .ZN(n8495) );
  NAND4_X1 U9196 ( .A1(n8378), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(n6729), .A4(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n6728) );
  NAND4_X1 U9197 ( .A1(n13811), .A2(n7543), .A3(P3_ADDR_REG_19__SCAN_IN), .A4(
        n14248), .ZN(n6730) );
  OAI21_X1 U9198 ( .B1(n8495), .B2(n6732), .A(n6731), .ZN(n8490) );
  NAND2_X1 U9199 ( .A1(n10704), .A2(n6736), .ZN(n6733) );
  NAND2_X1 U9200 ( .A1(n6733), .A2(n6734), .ZN(n11079) );
  NAND2_X1 U9201 ( .A1(n10961), .A2(n10960), .ZN(n11071) );
  NAND2_X1 U9202 ( .A1(n11393), .A2(n11392), .ZN(n13898) );
  NAND2_X1 U9203 ( .A1(n12889), .A2(n12890), .ZN(n12888) );
  NAND3_X1 U9204 ( .A1(n12894), .A2(n12893), .A3(n6750), .ZN(n6749) );
  NAND2_X1 U9205 ( .A1(n6749), .A2(n6748), .ZN(n7457) );
  INV_X1 U9206 ( .A(n6580), .ZN(n6752) );
  NAND2_X1 U9207 ( .A1(n6755), .A2(n6753), .ZN(n12815) );
  INV_X1 U9208 ( .A(n12807), .ZN(n6754) );
  NAND3_X1 U9209 ( .A1(n7448), .A2(n7450), .A3(n6756), .ZN(n6755) );
  NAND2_X1 U9210 ( .A1(n12807), .A2(n12806), .ZN(n6756) );
  INV_X1 U9211 ( .A(n12806), .ZN(n6757) );
  NAND2_X1 U9212 ( .A1(n12845), .A2(n6760), .ZN(n6758) );
  NAND2_X1 U9213 ( .A1(n6758), .A2(n6759), .ZN(n12856) );
  NAND3_X1 U9214 ( .A1(n6587), .A2(n12974), .A3(n12994), .ZN(n6763) );
  NAND3_X1 U9215 ( .A1(n7285), .A2(n7507), .A3(n7288), .ZN(n7764) );
  NOR2_X1 U9216 ( .A1(n7175), .A2(n7532), .ZN(n6768) );
  NAND3_X1 U9217 ( .A1(n6901), .A2(n6900), .A3(n8247), .ZN(n7695) );
  NAND3_X1 U9218 ( .A1(n6772), .A2(n8207), .A3(n6771), .ZN(n6770) );
  AND2_X1 U9219 ( .A1(n6773), .A2(n11974), .ZN(n6772) );
  OAI21_X1 U9220 ( .B1(n8198), .B2(n8195), .A(n6774), .ZN(n6773) );
  NAND2_X1 U9221 ( .A1(n7694), .A2(n6779), .ZN(n6776) );
  NAND2_X1 U9222 ( .A1(n6776), .A2(n6777), .ZN(n7722) );
  NAND2_X1 U9223 ( .A1(n6782), .A2(n6783), .ZN(n8141) );
  NAND2_X1 U9224 ( .A1(n8124), .A2(n6785), .ZN(n6782) );
  AOI21_X1 U9225 ( .B1(n6785), .B2(n6787), .A(n6784), .ZN(n6783) );
  AOI21_X1 U9226 ( .B1(n6788), .B2(n6786), .A(n8137), .ZN(n6785) );
  AOI21_X1 U9227 ( .B1(n6792), .B2(n6796), .A(n6790), .ZN(n6789) );
  NAND2_X1 U9228 ( .A1(n8122), .A2(n10632), .ZN(n6796) );
  AND2_X1 U9229 ( .A1(n7572), .A2(n7573), .ZN(n6805) );
  NAND2_X1 U9230 ( .A1(n6807), .A2(n9552), .ZN(n8093) );
  INV_X1 U9231 ( .A(n7848), .ZN(n6809) );
  NAND3_X1 U9232 ( .A1(n6810), .A2(n6809), .A3(n6611), .ZN(n6808) );
  NAND3_X1 U9233 ( .A1(n6812), .A2(n6811), .A3(n7514), .ZN(n7871) );
  NAND2_X1 U9234 ( .A1(n7793), .A2(n6819), .ZN(n6816) );
  NAND2_X1 U9235 ( .A1(n6816), .A2(n6817), .ZN(n7820) );
  OAI22_X1 U9236 ( .A1(n6835), .A2(n7149), .B1(n8415), .B2(n8152), .ZN(n8156)
         );
  AOI21_X1 U9237 ( .B1(n6837), .B2(n6836), .A(n8151), .ZN(n6835) );
  MUX2_X1 U9238 ( .A(P3_REG1_REG_1__SCAN_IN), .B(P3_REG2_REG_1__SCAN_IN), .S(
        n8316), .Z(n8330) );
  MUX2_X1 U9239 ( .A(n8329), .B(n9891), .S(n8316), .Z(n14810) );
  MUX2_X1 U9240 ( .A(P3_REG1_REG_2__SCAN_IN), .B(P3_REG2_REG_2__SCAN_IN), .S(
        n8316), .Z(n8327) );
  MUX2_X1 U9241 ( .A(P3_REG1_REG_3__SCAN_IN), .B(P3_REG2_REG_3__SCAN_IN), .S(
        n8316), .Z(n8326) );
  MUX2_X1 U9242 ( .A(P3_REG1_REG_12__SCAN_IN), .B(P3_REG2_REG_12__SCAN_IN), 
        .S(n8316), .Z(n8351) );
  MUX2_X1 U9243 ( .A(P3_REG1_REG_16__SCAN_IN), .B(P3_REG2_REG_16__SCAN_IN), 
        .S(n8316), .Z(n8360) );
  MUX2_X1 U9244 ( .A(n8366), .B(n8367), .S(n8316), .Z(n8368) );
  MUX2_X1 U9245 ( .A(n8355), .B(n8356), .S(n8316), .Z(n8357) );
  AOI21_X1 U9246 ( .B1(n6845), .B2(n8100), .A(n8099), .ZN(n6844) );
  NAND3_X1 U9247 ( .A1(n8095), .A2(n8094), .A3(n10120), .ZN(n6846) );
  NOR2_X2 U9248 ( .A1(n12732), .A2(n14743), .ZN(n9026) );
  NOR2_X2 U9249 ( .A1(n9780), .A2(n14781), .ZN(n9807) );
  OR2_X2 U9250 ( .A1(n9414), .A2(n12791), .ZN(n9780) );
  NOR2_X2 U9251 ( .A1(n14713), .A2(n12773), .ZN(n9197) );
  NOR2_X2 U9252 ( .A1(n10142), .A2(n12823), .ZN(n10254) );
  AND2_X1 U9253 ( .A1(n13190), .A2(n6857), .ZN(n13168) );
  OR2_X1 U9254 ( .A1(n13190), .A2(n12975), .ZN(n6853) );
  NAND2_X1 U9255 ( .A1(n13190), .A2(n11886), .ZN(n13178) );
  NAND2_X1 U9256 ( .A1(n13190), .A2(n6855), .ZN(n13167) );
  NAND3_X1 U9257 ( .A1(n6854), .A2(n6853), .A3(n6851), .ZN(n13162) );
  NAND2_X1 U9258 ( .A1(n13190), .A2(n6579), .ZN(n6854) );
  NOR2_X2 U9259 ( .A1(n10931), .A2(n13404), .ZN(n11036) );
  NAND3_X1 U9260 ( .A1(n13236), .A2(n6861), .A3(n13299), .ZN(n13238) );
  NOR2_X2 U9261 ( .A1(n14192), .A2(n14193), .ZN(n14194) );
  NAND3_X1 U9262 ( .A1(n6873), .A2(n6872), .A3(n6870), .ZN(n6869) );
  NOR2_X2 U9263 ( .A1(n10306), .A2(n11238), .ZN(n10290) );
  NAND2_X1 U9264 ( .A1(n8477), .A2(n6876), .ZN(n8727) );
  INV_X1 U9265 ( .A(n6880), .ZN(n13852) );
  NOR2_X2 U9266 ( .A1(n10999), .A2(n13648), .ZN(n11113) );
  NOR2_X2 U9267 ( .A1(n10771), .A2(n14432), .ZN(n6888) );
  NAND3_X1 U9268 ( .A1(n8231), .A2(n8230), .A3(n12587), .ZN(n9549) );
  NAND2_X1 U9269 ( .A1(n12109), .A2(n12110), .ZN(n6895) );
  OAI211_X1 U9270 ( .C1(n12109), .C2(n6893), .A(n6890), .B(n6889), .ZN(n11981)
         );
  NAND2_X1 U9271 ( .A1(n12109), .A2(n6583), .ZN(n6889) );
  NAND2_X1 U9272 ( .A1(n6899), .A2(n6894), .ZN(n6891) );
  INV_X1 U9273 ( .A(n6907), .ZN(n11954) );
  NAND2_X1 U9274 ( .A1(n10662), .A2(n6584), .ZN(n6910) );
  NAND2_X1 U9275 ( .A1(n14277), .A2(n6916), .ZN(n6918) );
  INV_X1 U9276 ( .A(n6918), .ZN(n12052) );
  NAND2_X1 U9277 ( .A1(n13259), .A2(n6930), .ZN(n6929) );
  INV_X1 U9278 ( .A(n13368), .ZN(n6939) );
  NAND2_X1 U9279 ( .A1(n6944), .A2(n6942), .ZN(n10724) );
  NOR2_X2 U9280 ( .A1(n8529), .A2(n6945), .ZN(n7182) );
  NAND4_X1 U9281 ( .A1(n8907), .A2(n8515), .A3(n8903), .A4(n6946), .ZN(n6945)
         );
  INV_X2 U9282 ( .A(P2_IR_REG_15__SCAN_IN), .ZN(n8903) );
  XNOR2_X2 U9283 ( .A(n8288), .B(n9072), .ZN(n9067) );
  NAND2_X1 U9284 ( .A1(n8292), .A2(n6964), .ZN(n6960) );
  NAND2_X1 U9285 ( .A1(n13308), .A2(n6968), .ZN(n6967) );
  NAND2_X2 U9286 ( .A1(n8677), .A2(n13432), .ZN(n8899) );
  NAND2_X2 U9287 ( .A1(n6974), .A2(n6976), .ZN(n8677) );
  NAND2_X2 U9288 ( .A1(n6972), .A2(n6971), .ZN(n9097) );
  NAND3_X1 U9289 ( .A1(n6977), .A2(n6973), .A3(n11361), .ZN(n6971) );
  NAND3_X1 U9290 ( .A1(n6974), .A2(n6976), .A3(n11361), .ZN(n6972) );
  NAND2_X1 U9291 ( .A1(n8307), .A2(n6980), .ZN(n6978) );
  OAI21_X2 U9292 ( .B1(n12163), .B2(n6979), .A(n6978), .ZN(n12178) );
  NAND2_X1 U9293 ( .A1(n6980), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n6979) );
  INV_X1 U9294 ( .A(n12179), .ZN(n6980) );
  NAND2_X1 U9295 ( .A1(n9058), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n8287) );
  OAI21_X1 U9296 ( .B1(n8247), .B2(n7805), .A(n7593), .ZN(n6981) );
  INV_X1 U9297 ( .A(P3_IR_REG_31__SCAN_IN), .ZN(n7805) );
  NAND2_X1 U9298 ( .A1(n9651), .A2(n6990), .ZN(n6986) );
  NOR2_X1 U9299 ( .A1(n6994), .A2(n9587), .ZN(n6992) );
  INV_X1 U9300 ( .A(n6995), .ZN(n9652) );
  AND2_X1 U9301 ( .A1(n9589), .A2(n9590), .ZN(n6994) );
  OAI211_X1 U9302 ( .C1(n13623), .C2(n7001), .A(n6998), .B(n6996), .ZN(n13549)
         );
  NAND2_X1 U9303 ( .A1(n13623), .A2(n6997), .ZN(n6996) );
  NOR2_X1 U9304 ( .A1(n7000), .A2(n13543), .ZN(n6997) );
  OAI22_X1 U9305 ( .A1(n7000), .A2(n6999), .B1(n13543), .B2(n7002), .ZN(n6998)
         );
  NOR2_X1 U9306 ( .A1(n13543), .A2(n13493), .ZN(n6999) );
  NAND2_X1 U9307 ( .A1(n13493), .A2(n13543), .ZN(n7001) );
  NAND2_X1 U9308 ( .A1(n7003), .A2(n7004), .ZN(n13479) );
  NAND2_X1 U9309 ( .A1(n13509), .A2(n7006), .ZN(n7003) );
  NAND2_X1 U9310 ( .A1(n10797), .A2(n10796), .ZN(n10846) );
  NAND2_X1 U9311 ( .A1(n10797), .A2(n7009), .ZN(n7008) );
  NAND2_X1 U9312 ( .A1(n8470), .A2(n7013), .ZN(n8481) );
  NAND2_X1 U9313 ( .A1(n8470), .A2(n6581), .ZN(n7014) );
  NAND2_X1 U9314 ( .A1(n7015), .A2(n6585), .ZN(n11839) );
  NAND3_X1 U9315 ( .A1(n7311), .A2(n7025), .A3(n8581), .ZN(n11199) );
  NAND2_X1 U9316 ( .A1(n10216), .A2(n10215), .ZN(n10218) );
  NAND2_X1 U9317 ( .A1(n9949), .A2(n11577), .ZN(n7026) );
  NAND2_X1 U9318 ( .A1(n10763), .A2(n7030), .ZN(n7027) );
  NAND2_X1 U9319 ( .A1(n7027), .A2(n7028), .ZN(n14390) );
  OAI211_X1 U9320 ( .C1(n10285), .C2(n7035), .A(n6576), .B(n7033), .ZN(n7034)
         );
  OR2_X1 U9321 ( .A1(n11585), .A2(n7036), .ZN(n7033) );
  NAND2_X1 U9322 ( .A1(n7042), .A2(n7044), .ZN(n11900) );
  NAND2_X1 U9323 ( .A1(n13884), .A2(n6492), .ZN(n7042) );
  NAND2_X1 U9324 ( .A1(n7058), .A2(n7057), .ZN(n13941) );
  INV_X1 U9325 ( .A(n7069), .ZN(n13886) );
  INV_X1 U9326 ( .A(n11898), .ZN(n7070) );
  NAND2_X1 U9327 ( .A1(n8477), .A2(n7076), .ZN(n8725) );
  NAND2_X1 U9328 ( .A1(n8725), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8726) );
  INV_X1 U9329 ( .A(n10151), .ZN(n11576) );
  XNOR2_X1 U9330 ( .A(n8472), .B(P1_IR_REG_24__SCAN_IN), .ZN(n8730) );
  AOI21_X2 U9331 ( .B1(n9575), .B2(n13536), .A(n9574), .ZN(n9645) );
  NAND2_X1 U9332 ( .A1(n11896), .A2(n13941), .ZN(n13943) );
  NAND2_X1 U9333 ( .A1(n11035), .A2(n11034), .ZN(n11136) );
  NAND2_X1 U9334 ( .A1(n9793), .A2(n13004), .ZN(n10045) );
  NAND2_X1 U9335 ( .A1(n10063), .A2(n10062), .ZN(n10128) );
  NAND2_X1 U9336 ( .A1(n10724), .A2(n10723), .ZN(n14335) );
  NAND2_X1 U9337 ( .A1(n8901), .A2(n8900), .ZN(n9028) );
  NAND2_X1 U9338 ( .A1(n11853), .A2(n11852), .ZN(n13259) );
  NAND2_X1 U9339 ( .A1(n7078), .A2(n11576), .ZN(n11220) );
  NAND2_X1 U9340 ( .A1(n7081), .A2(n7079), .ZN(n7078) );
  NAND2_X1 U9341 ( .A1(n11554), .A2(n11210), .ZN(n7082) );
  NAND3_X1 U9342 ( .A1(n11227), .A2(n11226), .A3(n11231), .ZN(n7083) );
  NAND2_X1 U9343 ( .A1(n7083), .A2(n11229), .ZN(n11230) );
  NAND2_X1 U9344 ( .A1(n7085), .A2(n11390), .ZN(n7084) );
  NAND2_X1 U9345 ( .A1(n7089), .A2(n11391), .ZN(n7085) );
  INV_X1 U9346 ( .A(n11391), .ZN(n7087) );
  INV_X1 U9347 ( .A(n7089), .ZN(n7088) );
  INV_X1 U9348 ( .A(n11294), .ZN(n7101) );
  NAND3_X1 U9349 ( .A1(n7096), .A2(n7099), .A3(n7093), .ZN(n7092) );
  INV_X1 U9350 ( .A(n11286), .ZN(n7107) );
  NAND2_X1 U9351 ( .A1(n11321), .A2(n7109), .ZN(n7108) );
  NAND2_X1 U9352 ( .A1(n11270), .A2(n7131), .ZN(n7128) );
  OAI21_X1 U9353 ( .B1(n11270), .B2(n7132), .A(n7131), .ZN(n11276) );
  NAND2_X1 U9354 ( .A1(n7128), .A2(n7129), .ZN(n11275) );
  NAND2_X1 U9355 ( .A1(n11425), .A2(n7136), .ZN(n7133) );
  NAND2_X1 U9356 ( .A1(n7133), .A2(n7134), .ZN(n11443) );
  OAI21_X1 U9357 ( .B1(n11235), .B2(n7139), .A(n7138), .ZN(n11241) );
  NAND2_X1 U9358 ( .A1(n11234), .A2(n11237), .ZN(n7138) );
  NOR2_X1 U9359 ( .A1(n11237), .A2(n11234), .ZN(n7139) );
  NAND3_X1 U9360 ( .A1(n11246), .A2(n11245), .A3(n6586), .ZN(n7140) );
  NAND2_X1 U9361 ( .A1(n7140), .A2(n7141), .ZN(n11253) );
  INV_X1 U9362 ( .A(n11201), .ZN(n9274) );
  NAND2_X1 U9363 ( .A1(n7143), .A2(n9272), .ZN(n11201) );
  NAND2_X1 U9364 ( .A1(n9271), .A2(n7144), .ZN(n7143) );
  MUX2_X1 U9365 ( .A(n7147), .B(n7146), .S(n11499), .Z(n11215) );
  NAND2_X1 U9366 ( .A1(n7952), .A2(n7151), .ZN(n7150) );
  INV_X1 U9367 ( .A(n7162), .ZN(n7161) );
  OAI21_X1 U9368 ( .B1(n7950), .B2(n7166), .A(n7164), .ZN(n12474) );
  NAND2_X1 U9369 ( .A1(n12277), .A2(n14983), .ZN(n7174) );
  NAND2_X1 U9370 ( .A1(n7697), .A2(n7479), .ZN(n7794) );
  NAND2_X1 U9371 ( .A1(n7536), .A2(n7535), .ZN(n7541) );
  INV_X1 U9372 ( .A(n7549), .ZN(n7552) );
  NAND2_X1 U9373 ( .A1(n7549), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7550) );
  AND2_X2 U9374 ( .A1(n7445), .A2(n8441), .ZN(n8702) );
  NAND2_X1 U9375 ( .A1(n7193), .A2(n10743), .ZN(n7189) );
  NAND3_X1 U9376 ( .A1(n7190), .A2(n13010), .A3(n7189), .ZN(n10942) );
  AND2_X1 U9377 ( .A1(n7190), .A2(n7189), .ZN(n10744) );
  INV_X1 U9378 ( .A(n10742), .ZN(n7198) );
  INV_X1 U9379 ( .A(n7202), .ZN(n13243) );
  NAND2_X1 U9380 ( .A1(n13199), .A2(n6575), .ZN(n7204) );
  OAI211_X1 U9381 ( .C1(n13199), .C2(n7208), .A(n7204), .B(n7205), .ZN(n13325)
         );
  NAND2_X1 U9382 ( .A1(n13199), .A2(n6523), .ZN(n7210) );
  OAI21_X1 U9383 ( .B1(n13199), .B2(n6524), .A(n11883), .ZN(n13188) );
  NAND2_X1 U9384 ( .A1(n8512), .A2(n7219), .ZN(n8523) );
  INV_X1 U9385 ( .A(n9698), .ZN(n7223) );
  OAI21_X1 U9386 ( .B1(n7223), .B2(n7222), .A(n7221), .ZN(n9740) );
  NAND2_X1 U9387 ( .A1(n10400), .A2(n7232), .ZN(n7231) );
  NAND2_X1 U9388 ( .A1(n7237), .A2(n7239), .ZN(n9699) );
  NAND2_X1 U9389 ( .A1(n9458), .A2(n7241), .ZN(n7237) );
  NOR2_X1 U9390 ( .A1(n7473), .A2(n9464), .ZN(n7238) );
  NAND2_X1 U9391 ( .A1(n12662), .A2(n7247), .ZN(n7244) );
  OAI21_X2 U9392 ( .B1(n7251), .B2(n6501), .A(n6489), .ZN(n10403) );
  NAND3_X1 U9393 ( .A1(n7255), .A2(n7258), .A3(n7254), .ZN(n7253) );
  NAND2_X1 U9394 ( .A1(n7259), .A2(n7260), .ZN(n11754) );
  NAND2_X1 U9395 ( .A1(n12644), .A2(n7261), .ZN(n7259) );
  OAI21_X1 U9396 ( .B1(n12644), .B2(n7265), .A(n7263), .ZN(n12610) );
  NAND2_X1 U9397 ( .A1(n12644), .A2(n12643), .ZN(n7267) );
  OAI22_X1 U9398 ( .A1(n14325), .A2(n6563), .B1(n7269), .B2(n12654), .ZN(
        n12652) );
  NAND2_X1 U9399 ( .A1(n7722), .A2(n7721), .ZN(n7275) );
  NOR2_X1 U9400 ( .A1(n7970), .A2(n7277), .ZN(n7926) );
  AOI21_X1 U9401 ( .B1(n7970), .B2(n7280), .A(n7279), .ZN(n7278) );
  NOR2_X1 U9402 ( .A1(n12022), .A2(n11973), .ZN(n7279) );
  XNOR2_X2 U9403 ( .A(n12022), .B(n7281), .ZN(n7970) );
  NAND2_X1 U9404 ( .A1(n7287), .A2(n7286), .ZN(n7285) );
  NAND2_X1 U9405 ( .A1(n7291), .A2(n7290), .ZN(n7748) );
  NAND2_X1 U9406 ( .A1(n7505), .A2(n7504), .ZN(n7506) );
  INV_X1 U9407 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n7292) );
  NAND2_X1 U9408 ( .A1(n7834), .A2(n7832), .ZN(n7293) );
  NAND2_X1 U9409 ( .A1(n7293), .A2(n7511), .ZN(n7512) );
  INV_X1 U9410 ( .A(n7294), .ZN(n7849) );
  NOR2_X4 U9411 ( .A1(n8587), .A2(n8465), .ZN(n8581) );
  NOR2_X2 U9412 ( .A1(n8463), .A2(n8462), .ZN(n7311) );
  NAND2_X1 U9413 ( .A1(n10769), .A2(n7316), .ZN(n7313) );
  NAND2_X1 U9414 ( .A1(n13948), .A2(n7324), .ZN(n11915) );
  NOR2_X1 U9415 ( .A1(n13880), .A2(n7333), .ZN(n13861) );
  NAND2_X1 U9416 ( .A1(n13919), .A2(n7334), .ZN(n11920) );
  INV_X1 U9417 ( .A(n8479), .ZN(n7339) );
  INV_X1 U9418 ( .A(n7341), .ZN(n8773) );
  NAND2_X1 U9419 ( .A1(n14872), .A2(n7344), .ZN(n7342) );
  INV_X1 U9420 ( .A(n7345), .ZN(n8267) );
  INV_X1 U9421 ( .A(n7354), .ZN(n9391) );
  INV_X1 U9422 ( .A(n8254), .ZN(n7353) );
  NAND2_X1 U9423 ( .A1(n8274), .A2(n7359), .ZN(n7355) );
  XNOR2_X1 U9424 ( .A(n8273), .B(n12247), .ZN(n12234) );
  OAI21_X1 U9425 ( .B1(n12198), .B2(n7364), .A(n7363), .ZN(n12214) );
  AOI21_X1 U9426 ( .B1(n8100), .B2(n7366), .A(n8205), .ZN(n8099) );
  INV_X1 U9427 ( .A(n12015), .ZN(n7367) );
  NAND2_X1 U9428 ( .A1(n12414), .A2(n7815), .ZN(n12415) );
  NAND2_X1 U9429 ( .A1(n7790), .A2(n7368), .ZN(n12414) );
  NAND2_X1 U9430 ( .A1(n10807), .A2(n7371), .ZN(n7370) );
  NAND2_X1 U9431 ( .A1(n12465), .A2(n7375), .ZN(n7374) );
  NAND2_X1 U9432 ( .A1(n7374), .A2(n7376), .ZN(n12436) );
  OAI21_X1 U9433 ( .B1(n12351), .B2(n7882), .A(n7881), .ZN(n12336) );
  NAND2_X1 U9434 ( .A1(n7882), .A2(n7881), .ZN(n7387) );
  NAND2_X1 U9435 ( .A1(n12401), .A2(n7392), .ZN(n7391) );
  NAND3_X1 U9436 ( .A1(n7407), .A2(n11080), .A3(n11166), .ZN(n11167) );
  NAND2_X1 U9437 ( .A1(n11079), .A2(n11077), .ZN(n7408) );
  NAND2_X1 U9438 ( .A1(n8658), .A2(n8657), .ZN(n8767) );
  NAND3_X1 U9439 ( .A1(n7413), .A2(n7416), .A3(n7412), .ZN(n7410) );
  NAND2_X1 U9440 ( .A1(n8965), .A2(n7422), .ZN(n7418) );
  NAND2_X1 U9441 ( .A1(n11481), .A2(n11480), .ZN(n7433) );
  INV_X1 U9442 ( .A(n10536), .ZN(n7436) );
  NAND2_X1 U9443 ( .A1(n12751), .A2(n12750), .ZN(n7442) );
  NAND3_X1 U9444 ( .A1(n12751), .A2(n12750), .A3(n7441), .ZN(n7440) );
  INV_X1 U9445 ( .A(n12758), .ZN(n7441) );
  NAND2_X1 U9446 ( .A1(n7442), .A2(n12758), .ZN(n12762) );
  OAI211_X2 U9447 ( .C1(n9019), .C2(n8899), .A(n7444), .B(n7443), .ZN(n12740)
         );
  NAND2_X1 U9448 ( .A1(n12932), .A2(n12740), .ZN(n12742) );
  NAND2_X1 U9449 ( .A1(n9018), .A2(n9017), .ZN(n7444) );
  OAI21_X1 U9450 ( .B1(n12798), .B2(n12797), .A(n7449), .ZN(n7448) );
  INV_X1 U9451 ( .A(n12848), .ZN(n7453) );
  NAND2_X1 U9452 ( .A1(n7462), .A2(n7461), .ZN(n7459) );
  OAI21_X1 U9453 ( .B1(n12827), .B2(n7459), .A(n7460), .ZN(n7458) );
  NAND2_X1 U9454 ( .A1(n12915), .A2(n7466), .ZN(n7464) );
  NAND2_X1 U9455 ( .A1(n7464), .A2(n7465), .ZN(n12919) );
  NAND2_X1 U9456 ( .A1(n7464), .A2(n7463), .ZN(n12926) );
  NAND2_X1 U9457 ( .A1(n12046), .A2(n12047), .ZN(n11967) );
  NAND2_X1 U9458 ( .A1(n6513), .A2(P3_REG1_REG_1__SCAN_IN), .ZN(n7565) );
  OR2_X1 U9459 ( .A1(n14031), .A2(n14541), .ZN(n14036) );
  NAND2_X1 U9460 ( .A1(n10114), .A2(n8096), .ZN(n14947) );
  NOR2_X1 U9461 ( .A1(n8257), .A2(n9894), .ZN(n14839) );
  NAND2_X1 U9462 ( .A1(n12378), .A2(n7956), .ZN(n12376) );
  NAND2_X1 U9463 ( .A1(n12932), .A2(n13067), .ZN(n12734) );
  OAI211_X1 U9464 ( .C1(n12731), .C2(n6477), .A(n12730), .B(n12729), .ZN(
        n12736) );
  INV_X1 U9465 ( .A(n9232), .ZN(n9128) );
  INV_X1 U9466 ( .A(n12889), .ZN(n12892) );
  INV_X1 U9467 ( .A(n8093), .ZN(n9551) );
  NAND2_X1 U9468 ( .A1(n9437), .A2(n9441), .ZN(n12731) );
  OAI21_X1 U9469 ( .B1(n10934), .B2(n10933), .A(n10932), .ZN(n11032) );
  INV_X1 U9470 ( .A(n11991), .ZN(n8711) );
  NAND2_X1 U9471 ( .A1(n7948), .A2(n9522), .ZN(n14967) );
  OAI211_X1 U9472 ( .C1(n8073), .C2(n9280), .A(n7582), .B(n7581), .ZN(n9522)
         );
  AOI21_X2 U9473 ( .B1(n10253), .B2(n10252), .A(n10251), .ZN(n10743) );
  NAND2_X1 U9474 ( .A1(n11992), .A2(n15038), .ZN(n11993) );
  CLKBUF_X3 U9475 ( .A(n9113), .Z(n11701) );
  OR2_X1 U9476 ( .A1(n15038), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n7469) );
  AND2_X2 U9477 ( .A1(n9890), .A2(n14959), .ZN(n14979) );
  INV_X2 U9478 ( .A(n14979), .ZN(n14977) );
  NAND2_X1 U9479 ( .A1(n9208), .A2(n14735), .ZN(n14795) );
  NAND2_X1 U9480 ( .A1(n12985), .A2(n12984), .ZN(n12993) );
  AND2_X1 U9481 ( .A1(n11213), .A2(n11215), .ZN(n7471) );
  AND2_X1 U9482 ( .A1(n11218), .A2(n11217), .ZN(n7472) );
  AND2_X1 U9483 ( .A1(n9463), .A2(n9462), .ZN(n7473) );
  OR2_X1 U9484 ( .A1(n12541), .A2(n12537), .ZN(n7475) );
  NOR2_X1 U9485 ( .A1(P2_IR_REG_29__SCAN_IN), .A2(P2_IR_REG_28__SCAN_IN), .ZN(
        n7476) );
  INV_X1 U9486 ( .A(P1_DATAO_REG_12__SCAN_IN), .ZN(n8889) );
  INV_X1 U9487 ( .A(n8350), .ZN(n12158) );
  INV_X1 U9488 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n8502) );
  INV_X1 U9489 ( .A(n13053), .ZN(n10740) );
  INV_X1 U9490 ( .A(SI_18_), .ZN(n9821) );
  INV_X1 U9491 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n12013) );
  AND2_X1 U9492 ( .A1(n14742), .A2(n13026), .ZN(n7478) );
  INV_X1 U9493 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n9246) );
  INV_X1 U9494 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n10761) );
  AND4_X1 U9495 ( .A1(n7528), .A2(n7527), .A3(n7749), .A4(n7724), .ZN(n7479)
         );
  INV_X1 U9496 ( .A(P3_REG3_REG_9__SCAN_IN), .ZN(n7686) );
  INV_X1 U9497 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n9251) );
  XNOR2_X1 U9498 ( .A(n9024), .B(n13066), .ZN(n9101) );
  INV_X1 U9499 ( .A(n15015), .ZN(n8422) );
  INV_X1 U9500 ( .A(n12071), .ZN(n12120) );
  AND3_X1 U9501 ( .A1(n7912), .A2(n7911), .A3(n7910), .ZN(n12071) );
  AND4_X1 U9502 ( .A1(n8440), .A2(n8439), .A3(n8438), .A4(n8437), .ZN(n7480)
         );
  AND2_X1 U9503 ( .A1(n11673), .A2(n11672), .ZN(n7481) );
  OR2_X1 U9504 ( .A1(n11072), .A2(SI_22_), .ZN(n7482) );
  INV_X1 U9505 ( .A(n8181), .ZN(n8175) );
  CLKBUF_X3 U9506 ( .A(n11215), .Z(n11551) );
  CLKBUF_X3 U9507 ( .A(n9619), .Z(n13442) );
  NAND2_X1 U9508 ( .A1(n13066), .A2(n6477), .ZN(n12741) );
  OAI21_X1 U9509 ( .B1(n12736), .B2(n12737), .A(n12735), .ZN(n12745) );
  AOI21_X1 U9510 ( .B1(n12776), .B2(n6477), .A(n12775), .ZN(n12782) );
  OAI21_X1 U9511 ( .B1(n12785), .B2(n12784), .A(n12783), .ZN(n12794) );
  INV_X1 U9512 ( .A(n12816), .ZN(n12817) );
  AOI21_X1 U9513 ( .B1(n12827), .B2(n12826), .A(n12824), .ZN(n12825) );
  OAI21_X1 U9514 ( .B1(n12853), .B2(n6477), .A(n12852), .ZN(n12854) );
  INV_X1 U9515 ( .A(n12890), .ZN(n12891) );
  INV_X1 U9516 ( .A(P3_IR_REG_22__SCAN_IN), .ZN(n7529) );
  INV_X1 U9517 ( .A(n13010), .ZN(n13012) );
  INV_X1 U9518 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7510) );
  INV_X1 U9519 ( .A(P2_IR_REG_3__SCAN_IN), .ZN(n8429) );
  INV_X1 U9520 ( .A(n8248), .ZN(n8249) );
  INV_X1 U9521 ( .A(P3_REG2_REG_12__SCAN_IN), .ZN(n8264) );
  INV_X1 U9522 ( .A(P3_IR_REG_24__SCAN_IN), .ZN(n7533) );
  INV_X1 U9523 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n8437) );
  OAI21_X1 U9524 ( .B1(n9832), .B2(n9836), .A(n9831), .ZN(n9833) );
  INV_X1 U9525 ( .A(n14550), .ZN(n9667) );
  NAND2_X1 U9526 ( .A1(n11457), .A2(n11177), .ZN(n11179) );
  INV_X1 U9527 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n8967) );
  NAND2_X1 U9528 ( .A1(n14183), .A2(n14142), .ZN(n14143) );
  OR2_X1 U9529 ( .A1(n8411), .A2(n8086), .ZN(n8067) );
  OAI221_X1 U9530 ( .B1(n9226), .B2(P3_REG2_REG_0__SCAN_IN), .C1(n9226), .C2(
        n8551), .A(n8246), .ZN(n9221) );
  AND2_X1 U9531 ( .A1(n8423), .A2(n9376), .ZN(n8085) );
  OR2_X1 U9532 ( .A1(n7964), .A2(n12312), .ZN(n7966) );
  INV_X1 U9533 ( .A(n12438), .ZN(n11936) );
  INV_X1 U9534 ( .A(n9758), .ZN(n8230) );
  INV_X1 U9535 ( .A(P3_IR_REG_25__SCAN_IN), .ZN(n7534) );
  INV_X1 U9536 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n7503) );
  INV_X1 U9537 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n9963) );
  OR2_X1 U9538 ( .A1(n12810), .A2(n13057), .ZN(n10139) );
  INV_X1 U9539 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n8672) );
  INV_X1 U9540 ( .A(n9833), .ZN(n9834) );
  INV_X1 U9541 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n10605) );
  OR2_X1 U9542 ( .A1(n9593), .A2(n9303), .ZN(n9304) );
  INV_X1 U9543 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n9850) );
  NAND2_X1 U9544 ( .A1(n11179), .A2(n11178), .ZN(n11476) );
  AND2_X1 U9545 ( .A1(SI_24_), .A2(n11077), .ZN(n11078) );
  NAND2_X1 U9546 ( .A1(n9233), .A2(n15194), .ZN(n9238) );
  INV_X1 U9547 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n8488) );
  XNOR2_X1 U9548 ( .A(n8375), .B(n8229), .ZN(n8233) );
  OR2_X1 U9549 ( .A1(n7896), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n7908) );
  INV_X1 U9550 ( .A(n8655), .ZN(n8266) );
  NOR2_X1 U9551 ( .A1(n12242), .A2(n8314), .ZN(n12262) );
  AND2_X1 U9552 ( .A1(n8160), .A2(n8166), .ZN(n12402) );
  INV_X1 U9553 ( .A(n9360), .ZN(n8375) );
  INV_X1 U9554 ( .A(n12473), .ZN(n12480) );
  INV_X1 U9555 ( .A(n12100), .ZN(n12437) );
  INV_X1 U9556 ( .A(P3_IR_REG_12__SCAN_IN), .ZN(n7749) );
  AND2_X1 U9557 ( .A1(n8564), .A2(P2_DATAO_REG_6__SCAN_IN), .ZN(n7493) );
  INV_X1 U9558 ( .A(n10402), .ZN(n10399) );
  OR2_X1 U9559 ( .A1(n9964), .A2(n9963), .ZN(n10064) );
  INV_X1 U9560 ( .A(n13215), .ZN(n11880) );
  INV_X1 U9561 ( .A(n14322), .ZN(n12710) );
  INV_X1 U9562 ( .A(n10745), .ZN(n14347) );
  OR2_X1 U9563 ( .A1(n10169), .A2(n10168), .ZN(n10170) );
  AND2_X1 U9564 ( .A1(n10414), .A2(n10413), .ZN(n10415) );
  INV_X1 U9565 ( .A(n13551), .ZN(n11829) );
  OR2_X1 U9566 ( .A1(n9838), .A2(n9837), .ZN(n9839) );
  AND2_X1 U9567 ( .A1(n10888), .A2(n10889), .ZN(n10887) );
  NAND2_X1 U9568 ( .A1(n11565), .A2(n11564), .ZN(n11566) );
  OR2_X1 U9569 ( .A1(n11332), .A2(n11331), .ZN(n11344) );
  OR2_X1 U9570 ( .A1(n10685), .A2(n10684), .ZN(n10775) );
  XNOR2_X1 U9571 ( .A(n14038), .B(n13847), .ZN(n11921) );
  INV_X1 U9572 ( .A(n11395), .ZN(n11396) );
  NOR2_X1 U9573 ( .A1(n9851), .A2(n9850), .ZN(n9869) );
  INV_X1 U9574 ( .A(n11575), .ZN(n14521) );
  OR2_X1 U9575 ( .A1(n9663), .A2(P1_D_REG_1__SCAN_IN), .ZN(n9255) );
  NAND2_X1 U9576 ( .A1(n8481), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8472) );
  NAND2_X1 U9577 ( .A1(n9240), .A2(n15144), .ZN(n9364) );
  INV_X1 U9578 ( .A(P1_IR_REG_5__SCAN_IN), .ZN(n8582) );
  NOR2_X1 U9579 ( .A1(n7841), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n7853) );
  INV_X1 U9580 ( .A(P3_REG3_REG_8__SCAN_IN), .ZN(n15058) );
  NAND2_X1 U9581 ( .A1(n11962), .A2(n12027), .ZN(n11963) );
  NAND2_X1 U9582 ( .A1(n7808), .A2(n12063), .ZN(n7825) );
  AND2_X1 U9583 ( .A1(n7853), .A2(n12079), .ZN(n7874) );
  NAND2_X1 U9584 ( .A1(n9511), .A2(n9510), .ZN(n14281) );
  AND2_X1 U9585 ( .A1(n7939), .A2(n15066), .ZN(n12273) );
  AOI21_X1 U9586 ( .B1(n8380), .B2(n14843), .A(n8379), .ZN(n8381) );
  NAND2_X1 U9587 ( .A1(n7687), .A2(n7686), .ZN(n7702) );
  NOR2_X1 U9588 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(P3_REG3_REG_4__SCAN_IN), 
        .ZN(n7623) );
  INV_X1 U9589 ( .A(n12585), .ZN(n8021) );
  OR2_X1 U9590 ( .A1(n15015), .A2(n8424), .ZN(n8425) );
  AND2_X1 U9591 ( .A1(n8416), .A2(n8076), .ZN(n14949) );
  INV_X1 U9592 ( .A(n8110), .ZN(n10353) );
  XNOR2_X1 U9593 ( .A(n7518), .B(n11086), .ZN(n7894) );
  NOR2_X1 U9594 ( .A1(n10257), .A2(n10255), .ZN(n10733) );
  OR2_X1 U9595 ( .A1(n11121), .A2(n11120), .ZN(n11141) );
  OR2_X1 U9596 ( .A1(n8953), .A2(n12720), .ZN(n13027) );
  AND2_X1 U9597 ( .A1(n11744), .A2(n11743), .ZN(n13181) );
  NOR2_X1 U9598 ( .A1(n11141), .A2(n12683), .ZN(n11649) );
  INV_X1 U9599 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10500) );
  AOI22_X1 U9600 ( .A1(n13040), .A2(n12710), .B1(n13163), .B2(n13038), .ZN(
        n11873) );
  NOR2_X2 U9601 ( .A1(n13202), .A2(n13339), .ZN(n13190) );
  AOI21_X1 U9602 ( .B1(n13404), .B2(n13052), .A(n11026), .ZN(n11030) );
  INV_X1 U9603 ( .A(n14345), .ZN(n14336) );
  NAND2_X1 U9604 ( .A1(n14736), .A2(n9315), .ZN(n14706) );
  NAND2_X1 U9605 ( .A1(n8702), .A2(n7476), .ZN(n13424) );
  INV_X1 U9606 ( .A(P2_IR_REG_24__SCAN_IN), .ZN(n8443) );
  AND2_X1 U9607 ( .A1(n13526), .A2(n13524), .ZN(n11811) );
  INV_X1 U9608 ( .A(n14394), .ZN(n11283) );
  NAND2_X1 U9609 ( .A1(n11812), .A2(n11814), .ZN(n11815) );
  NAND2_X1 U9610 ( .A1(n11048), .A2(n11050), .ZN(n11051) );
  INV_X1 U9611 ( .A(n13639), .ZN(n13617) );
  NAND2_X1 U9612 ( .A1(n9632), .A2(P1_STATE_REG_SCAN_IN), .ZN(n13644) );
  NOR2_X1 U9613 ( .A1(n11344), .A2(n11343), .ZN(n11365) );
  NAND2_X1 U9614 ( .A1(n11312), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n11332) );
  INV_X1 U9615 ( .A(P1_ADDR_REG_3__SCAN_IN), .ZN(n14142) );
  INV_X1 U9616 ( .A(n11921), .ZN(n13826) );
  INV_X1 U9617 ( .A(n13887), .ZN(n13630) );
  AND2_X1 U9618 ( .A1(n9939), .A2(n9938), .ZN(n9945) );
  INV_X1 U9619 ( .A(n11582), .ZN(n10313) );
  NAND2_X1 U9620 ( .A1(n9945), .A2(n13881), .ZN(n13989) );
  INV_X1 U9621 ( .A(n14606), .ZN(n14580) );
  INV_X1 U9622 ( .A(n13657), .ZN(n11285) );
  XNOR2_X1 U9623 ( .A(n8962), .B(n15174), .ZN(n8960) );
  INV_X1 U9624 ( .A(n14281), .ZN(n12104) );
  INV_X1 U9625 ( .A(n14286), .ZN(n12112) );
  AND2_X1 U9626 ( .A1(n7562), .A2(n7561), .ZN(n11973) );
  AND4_X1 U9627 ( .A1(n7892), .A2(n7891), .A3(n7890), .A4(n7889), .ZN(n12070)
         );
  NOR2_X1 U9628 ( .A1(n7656), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7670) );
  INV_X1 U9629 ( .A(n14906), .ZN(n14957) );
  INV_X1 U9630 ( .A(n14959), .ZN(n14973) );
  AND3_X1 U9631 ( .A1(n8412), .A2(n8017), .A3(n8418), .ZN(n9887) );
  INV_X1 U9632 ( .A(n14298), .ZN(n15016) );
  OR2_X1 U9633 ( .A1(n14968), .A2(n6604), .ZN(n14983) );
  INV_X1 U9634 ( .A(n9495), .ZN(n8279) );
  INV_X1 U9635 ( .A(P3_IR_REG_30__SCAN_IN), .ZN(n12588) );
  INV_X1 U9636 ( .A(P3_IR_REG_20__SCAN_IN), .ZN(n7937) );
  INV_X1 U9637 ( .A(P3_IR_REG_11__SCAN_IN), .ZN(n7724) );
  INV_X1 U9638 ( .A(P3_IR_REG_8__SCAN_IN), .ZN(n7680) );
  INV_X1 U9639 ( .A(n12705), .ZN(n14328) );
  INV_X1 U9640 ( .A(n8952), .ZN(n13026) );
  INV_X1 U9641 ( .A(n9145), .ZN(n11663) );
  INV_X1 U9642 ( .A(n14639), .ZN(n14686) );
  AND2_X1 U9643 ( .A1(n8684), .A2(n11867), .ZN(n14692) );
  INV_X1 U9644 ( .A(n9329), .ZN(n14714) );
  INV_X1 U9645 ( .A(n13189), .ZN(n13186) );
  INV_X1 U9646 ( .A(n13017), .ZN(n13288) );
  XNOR2_X1 U9647 ( .A(n12791), .B(n9773), .ZN(n13001) );
  NAND2_X1 U9648 ( .A1(n12935), .A2(n8918), .ZN(n14740) );
  INV_X1 U9649 ( .A(n14735), .ZN(n9312) );
  OR2_X1 U9650 ( .A1(n12723), .A2(n13026), .ZN(n14793) );
  NAND2_X1 U9651 ( .A1(n14793), .A2(n9328), .ZN(n14768) );
  AND2_X1 U9652 ( .A1(n14737), .A2(n8954), .ZN(n9208) );
  AND2_X1 U9653 ( .A1(n9318), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8940) );
  AND2_X1 U9654 ( .A1(n11061), .A2(n10965), .ZN(n11659) );
  AND2_X1 U9655 ( .A1(n8517), .A2(n8553), .ZN(n14652) );
  OR2_X1 U9656 ( .A1(n9301), .A2(n9300), .ZN(n11613) );
  OR2_X1 U9657 ( .A1(n11470), .A2(n13546), .ZN(n11473) );
  AND2_X1 U9658 ( .A1(n11372), .A2(n11371), .ZN(n11917) );
  INV_X1 U9659 ( .A(n13801), .ZN(n14504) );
  AND2_X1 U9660 ( .A1(n8842), .A2(n8841), .ZN(n14508) );
  INV_X1 U9661 ( .A(n14006), .ZN(n14527) );
  INV_X1 U9662 ( .A(n14015), .ZN(n14383) );
  OR2_X1 U9663 ( .A1(n9297), .A2(n14544), .ZN(n14606) );
  AND2_X1 U9664 ( .A1(n14023), .A2(n14585), .ZN(n14541) );
  INV_X1 U9665 ( .A(n14541), .ZN(n14609) );
  INV_X1 U9666 ( .A(n14585), .ZN(n14599) );
  XNOR2_X1 U9667 ( .A(n8485), .B(n8471), .ZN(n9277) );
  AND2_X1 U9668 ( .A1(n14210), .A2(n14209), .ZN(n14258) );
  AND2_X1 U9669 ( .A1(n8372), .A2(n8371), .ZN(n14869) );
  INV_X1 U9670 ( .A(n14274), .ZN(n12095) );
  AND2_X1 U9671 ( .A1(n8061), .A2(n8043), .ZN(n9376) );
  INV_X1 U9672 ( .A(n12070), .ZN(n12122) );
  INV_X1 U9673 ( .A(n14846), .ZN(n14878) );
  NAND2_X1 U9674 ( .A1(n8374), .A2(n12602), .ZN(n14887) );
  NAND2_X1 U9675 ( .A1(n8374), .A2(n8282), .ZN(n14893) );
  AND2_X1 U9676 ( .A1(n10639), .A2(n10638), .ZN(n15009) );
  INV_X1 U9677 ( .A(n14941), .ZN(n12486) );
  NAND2_X1 U9678 ( .A1(n15038), .A2(n15016), .ZN(n12537) );
  AND2_X1 U9679 ( .A1(n15009), .A2(n15008), .ZN(n15033) );
  INV_X1 U9680 ( .A(SI_19_), .ZN(n15045) );
  INV_X1 U9681 ( .A(SI_14_), .ZN(n15089) );
  NAND2_X1 U9682 ( .A1(n9451), .A2(P2_STATE_REG_SCAN_IN), .ZN(n14334) );
  NAND2_X1 U9683 ( .A1(n9326), .A2(n9325), .ZN(n12705) );
  OR2_X1 U9684 ( .A1(n10739), .A2(n10738), .ZN(n13053) );
  OR2_X1 U9685 ( .A1(n8683), .A2(n11867), .ZN(n14639) );
  OR2_X1 U9686 ( .A1(n9105), .A2(n12988), .ZN(n13282) );
  INV_X1 U9687 ( .A(n13316), .ZN(n14708) );
  OR2_X1 U9688 ( .A1(n14731), .A2(n9096), .ZN(n13304) );
  NAND2_X1 U9689 ( .A1(n9208), .A2(n9312), .ZN(n14808) );
  OR2_X1 U9690 ( .A1(n14738), .A2(n14732), .ZN(n14733) );
  INV_X1 U9691 ( .A(n14736), .ZN(n14738) );
  INV_X1 U9692 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n9374) );
  INV_X1 U9693 ( .A(P1_DATAO_REG_3__SCAN_IN), .ZN(n8542) );
  INV_X1 U9694 ( .A(n13969), .ZN(n14083) );
  INV_X1 U9695 ( .A(n13647), .ZN(n13636) );
  INV_X1 U9696 ( .A(n11569), .ZN(n13653) );
  INV_X1 U9697 ( .A(n11917), .ZN(n13936) );
  OR2_X1 U9698 ( .A1(n8839), .A2(n12002), .ZN(n13801) );
  OR2_X1 U9699 ( .A1(n8839), .A2(n13680), .ZN(n14501) );
  INV_X1 U9700 ( .A(n13812), .ZN(n14018) );
  AND2_X1 U9701 ( .A1(n12004), .A2(n14532), .ZN(n14388) );
  NAND2_X1 U9702 ( .A1(n13893), .A2(n9943), .ZN(n14015) );
  INV_X1 U9703 ( .A(n14630), .ZN(n14627) );
  AND3_X1 U9704 ( .A1(n14431), .A2(n14430), .A3(n14429), .ZN(n14453) );
  INV_X1 U9705 ( .A(n14613), .ZN(n14611) );
  AND2_X2 U9706 ( .A1(n9687), .A2(n9938), .ZN(n14613) );
  AND2_X1 U9707 ( .A1(n9277), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8738) );
  INV_X1 U9708 ( .A(n11089), .ZN(n10714) );
  INV_X1 U9709 ( .A(n12143), .ZN(P3_U3897) );
  INV_X1 U9710 ( .A(n13667), .ZN(P1_U4016) );
  INV_X1 U9711 ( .A(P3_REG1_REG_27__SCAN_IN), .ZN(n8025) );
  INV_X1 U9712 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n14125) );
  NOR2_X1 U9713 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(n6834), .ZN(n7521) );
  INV_X1 U9714 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n13439) );
  INV_X1 U9715 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n14131) );
  AOI22_X1 U9716 ( .A1(P2_DATAO_REG_25__SCAN_IN), .A2(P1_DATAO_REG_25__SCAN_IN), .B1(n13439), .B2(n14131), .ZN(n7904) );
  INV_X1 U9717 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n10967) );
  AOI22_X1 U9718 ( .A1(P2_DATAO_REG_19__SCAN_IN), .A2(n12013), .B1(
        P1_DATAO_REG_19__SCAN_IN), .B2(n7510), .ZN(n7832) );
  INV_X1 U9719 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n9824) );
  AOI22_X1 U9720 ( .A1(P2_DATAO_REG_18__SCAN_IN), .A2(n9829), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n9824), .ZN(n7818) );
  AOI22_X1 U9721 ( .A1(P2_DATAO_REG_16__SCAN_IN), .A2(n9246), .B1(
        P1_DATAO_REG_16__SCAN_IN), .B2(n9251), .ZN(n7791) );
  AOI22_X1 U9722 ( .A1(P2_DATAO_REG_15__SCAN_IN), .A2(n9358), .B1(
        P1_DATAO_REG_15__SCAN_IN), .B2(n7296), .ZN(n7775) );
  XNOR2_X1 U9723 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .ZN(n7763) );
  INV_X1 U9724 ( .A(P1_DATAO_REG_0__SCAN_IN), .ZN(n7483) );
  NAND2_X1 U9725 ( .A1(n8537), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n7484) );
  XNOR2_X1 U9726 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(P2_DATAO_REG_2__SCAN_IN), 
        .ZN(n7590) );
  NAND2_X1 U9727 ( .A1(n7592), .A2(n7590), .ZN(n7486) );
  NAND2_X1 U9728 ( .A1(n8531), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n7485) );
  XNOR2_X1 U9729 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(P2_DATAO_REG_3__SCAN_IN), 
        .ZN(n7617) );
  NAND2_X1 U9730 ( .A1(n7487), .A2(P2_DATAO_REG_4__SCAN_IN), .ZN(n7488) );
  NAND2_X1 U9731 ( .A1(n7489), .A2(n7488), .ZN(n7632) );
  NAND2_X1 U9732 ( .A1(n7632), .A2(n7630), .ZN(n7492) );
  NAND2_X1 U9733 ( .A1(n7490), .A2(P2_DATAO_REG_5__SCAN_IN), .ZN(n7491) );
  NAND2_X1 U9734 ( .A1(n8592), .A2(P1_DATAO_REG_6__SCAN_IN), .ZN(n7494) );
  NAND2_X1 U9735 ( .A1(n8584), .A2(P1_DATAO_REG_7__SCAN_IN), .ZN(n7495) );
  NAND2_X1 U9736 ( .A1(n7496), .A2(n7495), .ZN(n7678) );
  NAND2_X1 U9737 ( .A1(n7678), .A2(n7676), .ZN(n7498) );
  NAND2_X1 U9738 ( .A1(n8605), .A2(P1_DATAO_REG_8__SCAN_IN), .ZN(n7497) );
  NAND2_X1 U9739 ( .A1(n7499), .A2(P1_DATAO_REG_9__SCAN_IN), .ZN(n7500) );
  XNOR2_X1 U9740 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(P2_DATAO_REG_10__SCAN_IN), 
        .ZN(n7709) );
  XNOR2_X1 U9741 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(P2_DATAO_REG_11__SCAN_IN), 
        .ZN(n7721) );
  NAND2_X1 U9742 ( .A1(n8786), .A2(P1_DATAO_REG_11__SCAN_IN), .ZN(n7502) );
  XNOR2_X1 U9743 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .ZN(n7738) );
  NAND2_X1 U9744 ( .A1(n7292), .A2(n7506), .ZN(n7507) );
  INV_X1 U9745 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n9370) );
  AOI22_X1 U9746 ( .A1(P2_DATAO_REG_17__SCAN_IN), .A2(n9374), .B1(
        P1_DATAO_REG_17__SCAN_IN), .B2(n9370), .ZN(n7803) );
  NAND2_X1 U9747 ( .A1(n7818), .A2(n7820), .ZN(n7509) );
  INV_X1 U9748 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n10708) );
  AOI22_X1 U9749 ( .A1(P2_DATAO_REG_21__SCAN_IN), .A2(n10761), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(n10708), .ZN(n7861) );
  INV_X1 U9750 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n7515) );
  AOI22_X1 U9751 ( .A1(P2_DATAO_REG_22__SCAN_IN), .A2(P1_DATAO_REG_22__SCAN_IN), .B1(n10967), .B2(n7515), .ZN(n7870) );
  INV_X1 U9752 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n11067) );
  INV_X1 U9753 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n11070) );
  AOI22_X1 U9754 ( .A1(P2_DATAO_REG_23__SCAN_IN), .A2(P1_DATAO_REG_23__SCAN_IN), .B1(n11067), .B2(n11070), .ZN(n7883) );
  NOR2_X1 U9755 ( .A1(n7884), .A2(n7883), .ZN(n7517) );
  NAND2_X1 U9756 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n7518), .ZN(n7520) );
  INV_X1 U9757 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n11086) );
  INV_X1 U9758 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n11084) );
  NAND2_X1 U9759 ( .A1(n7894), .A2(n11084), .ZN(n7519) );
  INV_X1 U9760 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n13433) );
  INV_X1 U9761 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n14123) );
  AOI22_X1 U9762 ( .A1(P2_DATAO_REG_27__SCAN_IN), .A2(P1_DATAO_REG_27__SCAN_IN), .B1(n13433), .B2(n14123), .ZN(n7522) );
  INV_X1 U9763 ( .A(n7522), .ZN(n7523) );
  NAND4_X1 U9764 ( .A1(n7650), .A2(n7607), .A3(n7648), .A4(n7525), .ZN(n7526)
         );
  NOR2_X1 U9765 ( .A1(P3_IR_REG_18__SCAN_IN), .A2(P3_IR_REG_23__SCAN_IN), .ZN(
        n7531) );
  NOR2_X1 U9766 ( .A1(P3_IR_REG_20__SCAN_IN), .A2(P3_IR_REG_19__SCAN_IN), .ZN(
        n7530) );
  NAND4_X1 U9767 ( .A1(n7531), .A2(n7530), .A3(n7529), .A4(n7931), .ZN(n7532)
         );
  NAND2_X1 U9768 ( .A1(n7541), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7537) );
  MUX2_X1 U9769 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7537), .S(
        P3_IR_REG_28__SCAN_IN), .Z(n7538) );
  NAND2_X1 U9770 ( .A1(n7539), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7540) );
  MUX2_X1 U9771 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7540), .S(
        P3_IR_REG_27__SCAN_IN), .Z(n7542) );
  NAND2_X1 U9772 ( .A1(n12601), .A2(n7616), .ZN(n7545) );
  NAND2_X1 U9773 ( .A1(n8047), .A2(SI_27_), .ZN(n7544) );
  NAND2_X2 U9774 ( .A1(n7545), .A2(n7544), .ZN(n12022) );
  INV_X1 U9775 ( .A(P3_REG3_REG_5__SCAN_IN), .ZN(n7622) );
  NAND2_X1 U9776 ( .A1(n7623), .A2(n7622), .ZN(n7640) );
  INV_X1 U9777 ( .A(P3_REG3_REG_12__SCAN_IN), .ZN(n7731) );
  INV_X1 U9778 ( .A(P3_REG3_REG_17__SCAN_IN), .ZN(n12063) );
  INV_X1 U9779 ( .A(P3_REG3_REG_20__SCAN_IN), .ZN(n12079) );
  NOR2_X1 U9780 ( .A1(P3_REG3_REG_22__SCAN_IN), .A2(P3_REG3_REG_21__SCAN_IN), 
        .ZN(n7546) );
  NAND2_X1 U9781 ( .A1(n7874), .A2(n7546), .ZN(n7887) );
  NOR2_X1 U9782 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(P3_REG3_REG_26__SCAN_IN), 
        .ZN(n7547) );
  INV_X1 U9783 ( .A(P3_REG3_REG_26__SCAN_IN), .ZN(n15206) );
  INV_X1 U9784 ( .A(P3_REG3_REG_27__SCAN_IN), .ZN(n15048) );
  AOI21_X1 U9785 ( .B1(n7917), .B2(n15206), .A(n15048), .ZN(n7548) );
  OR2_X1 U9786 ( .A1(n7939), .A2(n7548), .ZN(n12288) );
  NAND2_X1 U9787 ( .A1(n7552), .A2(n7551), .ZN(n7554) );
  NAND2_X1 U9788 ( .A1(n12288), .A2(n7625), .ZN(n7562) );
  NAND2_X1 U9789 ( .A1(n7556), .A2(P3_REG2_REG_27__SCAN_IN), .ZN(n7560) );
  AND2_X2 U9790 ( .A1(n7557), .A2(n12015), .ZN(n7563) );
  NAND2_X1 U9791 ( .A1(n8055), .A2(P3_REG0_REG_27__SCAN_IN), .ZN(n7559) );
  INV_X1 U9792 ( .A(n7557), .ZN(n12595) );
  NAND2_X1 U9793 ( .A1(n8039), .A2(P3_REG1_REG_27__SCAN_IN), .ZN(n7558) );
  AND3_X1 U9794 ( .A1(n7560), .A2(n7559), .A3(n7558), .ZN(n7561) );
  INV_X1 U9795 ( .A(P3_REG2_REG_1__SCAN_IN), .ZN(n14976) );
  OR2_X1 U9796 ( .A1(n7585), .A2(n14976), .ZN(n7567) );
  NAND2_X1 U9797 ( .A1(n6520), .A2(P3_REG3_REG_1__SCAN_IN), .ZN(n7566) );
  NAND2_X1 U9798 ( .A1(n7563), .A2(P3_REG0_REG_1__SCAN_IN), .ZN(n7564) );
  INV_X1 U9799 ( .A(SI_1_), .ZN(n8631) );
  XNOR2_X1 U9800 ( .A(n7568), .B(n7578), .ZN(n8629) );
  NAND2_X1 U9801 ( .A1(n7616), .A2(n8629), .ZN(n7573) );
  NAND2_X2 U9802 ( .A1(n7571), .A2(n7570), .ZN(n9226) );
  NAND2_X1 U9803 ( .A1(n7743), .A2(n8328), .ZN(n7572) );
  NAND2_X1 U9804 ( .A1(n12142), .A2(n7583), .ZN(n8092) );
  NAND2_X1 U9805 ( .A1(n8092), .A2(n8093), .ZN(n14966) );
  NAND2_X1 U9806 ( .A1(n6513), .A2(P3_REG1_REG_0__SCAN_IN), .ZN(n7577) );
  NAND2_X1 U9807 ( .A1(n7625), .A2(P3_REG3_REG_0__SCAN_IN), .ZN(n7576) );
  NAND2_X1 U9808 ( .A1(n7556), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n7575) );
  NAND2_X1 U9809 ( .A1(n7563), .A2(P3_REG0_REG_0__SCAN_IN), .ZN(n7574) );
  INV_X1 U9810 ( .A(SI_0_), .ZN(n9280) );
  INV_X1 U9811 ( .A(n7578), .ZN(n7580) );
  NAND2_X1 U9812 ( .A1(n6732), .A2(P1_DATAO_REG_0__SCAN_IN), .ZN(n7579) );
  NAND2_X1 U9813 ( .A1(n7580), .A2(n7579), .ZN(n8550) );
  NAND2_X1 U9814 ( .A1(n7616), .A2(n8550), .ZN(n7582) );
  NAND2_X1 U9815 ( .A1(n7743), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n7581) );
  NAND2_X1 U9816 ( .A1(n12144), .A2(n9522), .ZN(n14960) );
  NAND2_X1 U9817 ( .A1(n14966), .A2(n14960), .ZN(n7584) );
  NAND2_X1 U9818 ( .A1(n6807), .A2(n7583), .ZN(n9550) );
  NAND2_X1 U9819 ( .A1(n7584), .A2(n9550), .ZN(n10119) );
  NAND2_X1 U9820 ( .A1(n6513), .A2(P3_REG1_REG_2__SCAN_IN), .ZN(n7589) );
  NAND2_X1 U9821 ( .A1(n7625), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n7588) );
  NAND2_X1 U9822 ( .A1(n7563), .A2(P3_REG0_REG_2__SCAN_IN), .ZN(n7586) );
  INV_X1 U9823 ( .A(n7590), .ZN(n7591) );
  XNOR2_X1 U9824 ( .A(n7592), .B(n7591), .ZN(n8617) );
  NAND2_X1 U9825 ( .A1(n7616), .A2(n8617), .ZN(n7595) );
  NAND2_X1 U9826 ( .A1(n7743), .A2(n9058), .ZN(n7594) );
  OAI211_X1 U9827 ( .C1(n8073), .C2(SI_2_), .A(n7595), .B(n7594), .ZN(n9715)
         );
  INV_X1 U9828 ( .A(n9715), .ZN(n10117) );
  NAND2_X1 U9829 ( .A1(n9992), .A2(n10117), .ZN(n8096) );
  INV_X1 U9830 ( .A(n9992), .ZN(n12141) );
  INV_X1 U9831 ( .A(n10120), .ZN(n7596) );
  NAND2_X1 U9832 ( .A1(n10119), .A2(n7596), .ZN(n7598) );
  NAND2_X1 U9833 ( .A1(n9992), .A2(n9715), .ZN(n7597) );
  NAND2_X1 U9834 ( .A1(n7598), .A2(n7597), .ZN(n10275) );
  NAND2_X1 U9835 ( .A1(n7563), .A2(P3_REG0_REG_4__SCAN_IN), .ZN(n7603) );
  NAND2_X1 U9836 ( .A1(n6513), .A2(P3_REG1_REG_4__SCAN_IN), .ZN(n7602) );
  AND2_X1 U9837 ( .A1(P3_REG3_REG_4__SCAN_IN), .A2(P3_REG3_REG_3__SCAN_IN), 
        .ZN(n7599) );
  OR2_X1 U9838 ( .A1(n7599), .A2(n7623), .ZN(n10382) );
  NAND2_X1 U9839 ( .A1(n7625), .A2(n10382), .ZN(n7601) );
  NAND2_X1 U9840 ( .A1(n7556), .A2(P3_REG2_REG_4__SCAN_IN), .ZN(n7600) );
  INV_X1 U9841 ( .A(n7604), .ZN(n7605) );
  XNOR2_X1 U9842 ( .A(n7606), .B(n7605), .ZN(n8635) );
  NAND2_X1 U9843 ( .A1(n6488), .A2(n8635), .ZN(n7611) );
  NAND2_X1 U9844 ( .A1(n7608), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7609) );
  NAND2_X1 U9845 ( .A1(n7743), .A2(n9185), .ZN(n7610) );
  OAI211_X1 U9846 ( .C1(n8073), .C2(SI_4_), .A(n7611), .B(n7610), .ZN(n10327)
         );
  INV_X1 U9847 ( .A(n10327), .ZN(n10383) );
  NAND2_X1 U9848 ( .A1(n10033), .A2(n10383), .ZN(n8109) );
  INV_X1 U9849 ( .A(n10033), .ZN(n12139) );
  NAND2_X1 U9850 ( .A1(n12139), .A2(n10327), .ZN(n8103) );
  NAND2_X1 U9851 ( .A1(n8109), .A2(n8103), .ZN(n8101) );
  NAND2_X1 U9852 ( .A1(n6513), .A2(P3_REG1_REG_3__SCAN_IN), .ZN(n7615) );
  NAND2_X1 U9853 ( .A1(n7625), .A2(n15067), .ZN(n7614) );
  NAND2_X1 U9854 ( .A1(n7556), .A2(P3_REG2_REG_3__SCAN_IN), .ZN(n7613) );
  NAND2_X1 U9855 ( .A1(n7563), .A2(P3_REG0_REG_3__SCAN_IN), .ZN(n7612) );
  NAND4_X1 U9856 ( .A1(n7615), .A2(n7614), .A3(n7613), .A4(n7612), .ZN(n12140)
         );
  XNOR2_X1 U9857 ( .A(n7618), .B(n7284), .ZN(n8633) );
  NAND2_X1 U9858 ( .A1(n6488), .A2(n8633), .ZN(n7621) );
  NAND2_X1 U9859 ( .A1(P3_IR_REG_31__SCAN_IN), .A2(n6527), .ZN(n7619) );
  INV_X1 U9860 ( .A(n9072), .ZN(n8632) );
  NAND2_X1 U9861 ( .A1(n7743), .A2(n8632), .ZN(n7620) );
  OAI211_X1 U9862 ( .C1(n8073), .C2(SI_3_), .A(n7621), .B(n7620), .ZN(n9989)
         );
  OR2_X1 U9863 ( .A1(n12140), .A2(n9989), .ZN(n8087) );
  NAND2_X1 U9864 ( .A1(n12140), .A2(n9989), .ZN(n8100) );
  INV_X1 U9865 ( .A(n9989), .ZN(n14991) );
  AND2_X1 U9866 ( .A1(n12140), .A2(n14991), .ZN(n10276) );
  NAND2_X1 U9867 ( .A1(n8101), .A2(n10276), .ZN(n7636) );
  NAND2_X1 U9868 ( .A1(n7563), .A2(P3_REG0_REG_5__SCAN_IN), .ZN(n7629) );
  NAND2_X1 U9869 ( .A1(n6513), .A2(P3_REG1_REG_5__SCAN_IN), .ZN(n7628) );
  OR2_X1 U9870 ( .A1(n7623), .A2(n7622), .ZN(n7624) );
  NAND2_X1 U9871 ( .A1(n7640), .A2(n7624), .ZN(n14939) );
  NAND2_X1 U9872 ( .A1(n7625), .A2(n14939), .ZN(n7627) );
  NAND2_X1 U9873 ( .A1(n7556), .A2(P3_REG2_REG_5__SCAN_IN), .ZN(n7626) );
  INV_X1 U9874 ( .A(n7638), .ZN(n12138) );
  INV_X1 U9875 ( .A(n7630), .ZN(n7631) );
  XNOR2_X1 U9876 ( .A(n7632), .B(n7631), .ZN(n8627) );
  NAND2_X1 U9877 ( .A1(n6488), .A2(n8627), .ZN(n7635) );
  NOR2_X1 U9878 ( .A1(n7608), .A2(P3_IR_REG_4__SCAN_IN), .ZN(n7649) );
  OR2_X1 U9879 ( .A1(n7649), .A2(n7805), .ZN(n7633) );
  INV_X1 U9880 ( .A(n9398), .ZN(n8626) );
  NAND2_X1 U9881 ( .A1(n7743), .A2(n8626), .ZN(n7634) );
  OAI211_X1 U9882 ( .C1(n8073), .C2(SI_5_), .A(n7635), .B(n7634), .ZN(n10364)
         );
  NAND2_X1 U9883 ( .A1(n12138), .A2(n10364), .ZN(n8113) );
  INV_X1 U9884 ( .A(n10364), .ZN(n14940) );
  NAND2_X1 U9885 ( .A1(n7638), .A2(n14940), .ZN(n8105) );
  OR2_X1 U9886 ( .A1(n10033), .A2(n10327), .ZN(n10352) );
  AND3_X1 U9887 ( .A1(n7636), .A2(n8110), .A3(n10352), .ZN(n7637) );
  NAND2_X1 U9888 ( .A1(n7638), .A2(n10364), .ZN(n7639) );
  NAND2_X1 U9889 ( .A1(n7563), .A2(P3_REG0_REG_6__SCAN_IN), .ZN(n7645) );
  NAND2_X1 U9890 ( .A1(n6513), .A2(P3_REG1_REG_6__SCAN_IN), .ZN(n7644) );
  NAND2_X1 U9891 ( .A1(n7640), .A2(P3_REG3_REG_6__SCAN_IN), .ZN(n7641) );
  AND2_X1 U9892 ( .A1(n7656), .A2(n7641), .ZN(n14938) );
  INV_X1 U9893 ( .A(n14938), .ZN(n12099) );
  NAND2_X1 U9894 ( .A1(n7625), .A2(n12099), .ZN(n7643) );
  NAND2_X1 U9895 ( .A1(n7556), .A2(P3_REG2_REG_6__SCAN_IN), .ZN(n7642) );
  NAND4_X1 U9896 ( .A1(n7645), .A2(n7644), .A3(n7643), .A4(n7642), .ZN(n12137)
         );
  INV_X1 U9897 ( .A(SI_6_), .ZN(n15225) );
  XNOR2_X1 U9898 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(P2_DATAO_REG_6__SCAN_IN), 
        .ZN(n7646) );
  XNOR2_X1 U9899 ( .A(n7647), .B(n7646), .ZN(n8619) );
  NAND2_X1 U9900 ( .A1(n7616), .A2(n8619), .ZN(n7653) );
  NAND2_X1 U9901 ( .A1(n7649), .A2(n7648), .ZN(n7665) );
  NAND2_X1 U9902 ( .A1(n7665), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7651) );
  INV_X1 U9903 ( .A(n8620), .ZN(n14826) );
  NAND2_X1 U9904 ( .A1(n7743), .A2(n14826), .ZN(n7652) );
  OAI211_X1 U9905 ( .C1(n8073), .C2(n15225), .A(n7653), .B(n7652), .ZN(n14996)
         );
  INV_X1 U9906 ( .A(n14996), .ZN(n7654) );
  NOR2_X1 U9907 ( .A1(n12137), .A2(n7654), .ZN(n8107) );
  INV_X1 U9908 ( .A(n8107), .ZN(n8114) );
  NAND2_X1 U9909 ( .A1(n12137), .A2(n7654), .ZN(n8119) );
  INV_X1 U9910 ( .A(n14926), .ZN(n14929) );
  NAND2_X1 U9911 ( .A1(n14930), .A2(n14929), .ZN(n14928) );
  NAND2_X1 U9912 ( .A1(n12137), .A2(n14996), .ZN(n7655) );
  NAND2_X1 U9913 ( .A1(n14928), .A2(n7655), .ZN(n14916) );
  NAND2_X1 U9914 ( .A1(n6513), .A2(P3_REG1_REG_7__SCAN_IN), .ZN(n7662) );
  AND2_X1 U9915 ( .A1(n7656), .A2(P3_REG3_REG_7__SCAN_IN), .ZN(n7657) );
  NOR2_X1 U9916 ( .A1(n7670), .A2(n7657), .ZN(n14924) );
  INV_X1 U9917 ( .A(n14924), .ZN(n7658) );
  NAND2_X1 U9918 ( .A1(n6520), .A2(n7658), .ZN(n7661) );
  NAND2_X1 U9919 ( .A1(n7556), .A2(P3_REG2_REG_7__SCAN_IN), .ZN(n7660) );
  NAND2_X1 U9920 ( .A1(n8055), .A2(P3_REG0_REG_7__SCAN_IN), .ZN(n7659) );
  XNOR2_X1 U9921 ( .A(n7664), .B(n7663), .ZN(n8570) );
  NAND2_X1 U9922 ( .A1(n6488), .A2(n8570), .ZN(n7668) );
  OAI21_X1 U9923 ( .B1(n7665), .B2(P3_IR_REG_6__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7666) );
  XNOR2_X1 U9924 ( .A(n7666), .B(P3_IR_REG_7__SCAN_IN), .ZN(n8321) );
  INV_X1 U9925 ( .A(n8321), .ZN(n9901) );
  NAND2_X1 U9926 ( .A1(n7743), .A2(n9901), .ZN(n7667) );
  OAI211_X1 U9927 ( .C1(n8073), .C2(SI_7_), .A(n7668), .B(n7667), .ZN(n10438)
         );
  INV_X1 U9928 ( .A(n10438), .ZN(n15001) );
  NAND2_X1 U9929 ( .A1(n12101), .A2(n15001), .ZN(n8121) );
  NAND2_X1 U9930 ( .A1(n12136), .A2(n10438), .ZN(n8120) );
  INV_X1 U9931 ( .A(n14912), .ZN(n14915) );
  NAND2_X1 U9932 ( .A1(n12136), .A2(n15001), .ZN(n7669) );
  NAND2_X1 U9933 ( .A1(n7563), .A2(P3_REG0_REG_8__SCAN_IN), .ZN(n7675) );
  NAND2_X1 U9934 ( .A1(n6513), .A2(P3_REG1_REG_8__SCAN_IN), .ZN(n7674) );
  NOR2_X1 U9935 ( .A1(n7670), .A2(n15058), .ZN(n7671) );
  OR2_X1 U9936 ( .A1(n7687), .A2(n7671), .ZN(n10653) );
  NAND2_X1 U9937 ( .A1(n7625), .A2(n10653), .ZN(n7673) );
  NAND2_X1 U9938 ( .A1(n7556), .A2(P3_REG2_REG_8__SCAN_IN), .ZN(n7672) );
  INV_X1 U9939 ( .A(SI_8_), .ZN(n8625) );
  INV_X1 U9940 ( .A(n7676), .ZN(n7677) );
  XNOR2_X1 U9941 ( .A(n7678), .B(n7677), .ZN(n8622) );
  NAND2_X1 U9942 ( .A1(n7616), .A2(n8622), .ZN(n7683) );
  OR2_X1 U9943 ( .A1(n7679), .A2(n7805), .ZN(n7681) );
  XNOR2_X1 U9944 ( .A(n7681), .B(n7680), .ZN(n8624) );
  INV_X1 U9945 ( .A(n8624), .ZN(n14845) );
  NAND2_X1 U9946 ( .A1(n7743), .A2(n14845), .ZN(n7682) );
  OAI211_X1 U9947 ( .C1(n8073), .C2(n8625), .A(n7683), .B(n7682), .ZN(n10649)
         );
  NAND2_X1 U9948 ( .A1(n10521), .A2(n10649), .ZN(n8125) );
  INV_X1 U9949 ( .A(n10521), .ZN(n12135) );
  INV_X1 U9950 ( .A(n10649), .ZN(n7684) );
  NAND2_X1 U9951 ( .A1(n12135), .A2(n7684), .ZN(n8126) );
  NAND2_X1 U9952 ( .A1(n10521), .A2(n7684), .ZN(n7685) );
  NAND2_X1 U9953 ( .A1(n6513), .A2(P3_REG1_REG_9__SCAN_IN), .ZN(n7692) );
  NAND2_X1 U9954 ( .A1(n7563), .A2(P3_REG0_REG_9__SCAN_IN), .ZN(n7691) );
  OR2_X1 U9955 ( .A1(n7687), .A2(n7686), .ZN(n7688) );
  NAND2_X1 U9956 ( .A1(n7702), .A2(n7688), .ZN(n10812) );
  NAND2_X1 U9957 ( .A1(n7625), .A2(n10812), .ZN(n7690) );
  NAND2_X1 U9958 ( .A1(n7556), .A2(P3_REG2_REG_9__SCAN_IN), .ZN(n7689) );
  NAND4_X1 U9959 ( .A1(n7692), .A2(n7691), .A3(n7690), .A4(n7689), .ZN(n12134)
         );
  XNOR2_X1 U9960 ( .A(n7694), .B(n7693), .ZN(n8568) );
  NAND2_X1 U9961 ( .A1(n6488), .A2(n8568), .ZN(n7700) );
  NAND2_X1 U9962 ( .A1(n7695), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7696) );
  MUX2_X1 U9963 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7696), .S(
        P3_IR_REG_9__SCAN_IN), .Z(n7698) );
  NAND2_X1 U9964 ( .A1(n7698), .A2(n7723), .ZN(n10341) );
  NAND2_X1 U9965 ( .A1(n7743), .A2(n10341), .ZN(n7699) );
  OAI211_X1 U9966 ( .C1(n8073), .C2(SI_9_), .A(n7700), .B(n7699), .ZN(n10811)
         );
  INV_X1 U9967 ( .A(n10811), .ZN(n10524) );
  XNOR2_X1 U9968 ( .A(n12134), .B(n10524), .ZN(n8213) );
  NAND2_X1 U9969 ( .A1(n12134), .A2(n10524), .ZN(n7701) );
  NAND2_X1 U9970 ( .A1(n7563), .A2(P3_REG0_REG_10__SCAN_IN), .ZN(n7708) );
  NAND2_X1 U9971 ( .A1(n6513), .A2(P3_REG1_REG_10__SCAN_IN), .ZN(n7707) );
  NAND2_X1 U9972 ( .A1(n7702), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n7703) );
  AND2_X1 U9973 ( .A1(n7715), .A2(n7703), .ZN(n14910) );
  INV_X1 U9974 ( .A(n14910), .ZN(n7704) );
  NAND2_X1 U9975 ( .A1(n6520), .A2(n7704), .ZN(n7706) );
  NAND2_X1 U9976 ( .A1(n7556), .A2(P3_REG2_REG_10__SCAN_IN), .ZN(n7705) );
  XNOR2_X1 U9977 ( .A(n7710), .B(n7709), .ZN(n8566) );
  NAND2_X1 U9978 ( .A1(n6488), .A2(n8566), .ZN(n7714) );
  NAND2_X1 U9979 ( .A1(n7723), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7712) );
  INV_X1 U9980 ( .A(P3_IR_REG_10__SCAN_IN), .ZN(n7711) );
  XNOR2_X1 U9981 ( .A(n7712), .B(n7711), .ZN(n14866) );
  NAND2_X1 U9982 ( .A1(n7743), .A2(n14866), .ZN(n7713) );
  OAI211_X1 U9983 ( .C1(n8073), .C2(SI_10_), .A(n7714), .B(n7713), .ZN(n14905)
         );
  INV_X1 U9984 ( .A(n14905), .ZN(n15017) );
  NAND2_X1 U9985 ( .A1(n10580), .A2(n15017), .ZN(n8132) );
  NAND2_X1 U9986 ( .A1(n12133), .A2(n14905), .ZN(n8131) );
  NAND2_X1 U9987 ( .A1(n8132), .A2(n8131), .ZN(n14898) );
  NAND2_X1 U9988 ( .A1(n7563), .A2(P3_REG0_REG_11__SCAN_IN), .ZN(n7720) );
  NAND2_X1 U9989 ( .A1(n8039), .A2(P3_REG1_REG_11__SCAN_IN), .ZN(n7719) );
  AND2_X1 U9990 ( .A1(n7715), .A2(P3_REG3_REG_11__SCAN_IN), .ZN(n7716) );
  OR2_X1 U9991 ( .A1(n7716), .A2(n7732), .ZN(n10831) );
  NAND2_X1 U9992 ( .A1(n7625), .A2(n10831), .ZN(n7718) );
  NAND2_X1 U9993 ( .A1(n7556), .A2(P3_REG2_REG_11__SCAN_IN), .ZN(n7717) );
  XNOR2_X1 U9994 ( .A(n7722), .B(n7721), .ZN(n8651) );
  NAND2_X1 U9995 ( .A1(n7616), .A2(n8651), .ZN(n7727) );
  OR2_X1 U9996 ( .A1(n7723), .A2(P3_IR_REG_10__SCAN_IN), .ZN(n7741) );
  NAND2_X1 U9997 ( .A1(n7741), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7725) );
  XNOR2_X1 U9998 ( .A(n7725), .B(n7724), .ZN(n14877) );
  NAND2_X1 U9999 ( .A1(n7743), .A2(n14877), .ZN(n7726) );
  OAI211_X1 U10000 ( .C1(n8073), .C2(SI_11_), .A(n7727), .B(n7726), .ZN(n10918) );
  NAND2_X1 U10001 ( .A1(n10861), .A2(n10918), .ZN(n7728) );
  NAND2_X1 U10002 ( .A1(n10921), .A2(n7728), .ZN(n7730) );
  INV_X1 U10003 ( .A(n10918), .ZN(n10834) );
  NAND2_X1 U10004 ( .A1(n12132), .A2(n10834), .ZN(n7729) );
  NAND2_X1 U10005 ( .A1(n7563), .A2(P3_REG0_REG_12__SCAN_IN), .ZN(n7737) );
  NAND2_X1 U10006 ( .A1(n6513), .A2(P3_REG1_REG_12__SCAN_IN), .ZN(n7736) );
  OR2_X1 U10007 ( .A1(n7732), .A2(n7731), .ZN(n7733) );
  NAND2_X1 U10008 ( .A1(n7769), .A2(n7733), .ZN(n12476) );
  NAND2_X1 U10009 ( .A1(n7625), .A2(n12476), .ZN(n7735) );
  NAND2_X1 U10010 ( .A1(n7556), .A2(P3_REG2_REG_12__SCAN_IN), .ZN(n7734) );
  INV_X1 U10011 ( .A(n7738), .ZN(n7739) );
  XNOR2_X1 U10012 ( .A(n7740), .B(n7739), .ZN(n8585) );
  NAND2_X1 U10013 ( .A1(n7616), .A2(n8585), .ZN(n7745) );
  NOR2_X1 U10014 ( .A1(n7741), .A2(P3_IR_REG_11__SCAN_IN), .ZN(n7750) );
  OR2_X1 U10015 ( .A1(n7750), .A2(n7805), .ZN(n7742) );
  XNOR2_X1 U10016 ( .A(n7742), .B(P3_IR_REG_12__SCAN_IN), .ZN(n8350) );
  NAND2_X1 U10017 ( .A1(n7743), .A2(n8350), .ZN(n7744) );
  OAI211_X1 U10018 ( .C1(n8073), .C2(n15174), .A(n7745), .B(n7744), .ZN(n10663) );
  INV_X1 U10019 ( .A(n10663), .ZN(n12475) );
  NOR2_X1 U10020 ( .A1(n12131), .A2(n12475), .ZN(n8143) );
  INV_X1 U10021 ( .A(n8143), .ZN(n7951) );
  NAND2_X1 U10022 ( .A1(n12131), .A2(n12475), .ZN(n8140) );
  NAND2_X1 U10023 ( .A1(n12481), .A2(n12480), .ZN(n7747) );
  NAND2_X1 U10024 ( .A1(n12131), .A2(n10663), .ZN(n7746) );
  XNOR2_X1 U10025 ( .A(n7748), .B(P1_DATAO_REG_13__SCAN_IN), .ZN(n8656) );
  NAND2_X1 U10026 ( .A1(n8656), .A2(n6488), .ZN(n7757) );
  NAND2_X1 U10027 ( .A1(n7750), .A2(n7749), .ZN(n7752) );
  NAND2_X1 U10028 ( .A1(n7752), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7751) );
  MUX2_X1 U10029 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7751), .S(
        P3_IR_REG_13__SCAN_IN), .Z(n7753) );
  NAND2_X1 U10030 ( .A1(n7753), .A2(n7778), .ZN(n8655) );
  OAI22_X1 U10031 ( .A1(n8073), .A2(SI_13_), .B1(n8266), .B2(n7754), .ZN(n7755) );
  INV_X1 U10032 ( .A(n7755), .ZN(n7756) );
  NAND2_X1 U10033 ( .A1(n7757), .A2(n7756), .ZN(n14299) );
  NAND2_X1 U10034 ( .A1(n8055), .A2(P3_REG0_REG_13__SCAN_IN), .ZN(n7761) );
  NAND2_X1 U10035 ( .A1(n8039), .A2(P3_REG1_REG_13__SCAN_IN), .ZN(n7760) );
  XNOR2_X1 U10036 ( .A(n7769), .B(P3_REG3_REG_13__SCAN_IN), .ZN(n12468) );
  NAND2_X1 U10037 ( .A1(n7625), .A2(n12468), .ZN(n7759) );
  NAND2_X1 U10038 ( .A1(n7556), .A2(P3_REG2_REG_13__SCAN_IN), .ZN(n7758) );
  NAND4_X1 U10039 ( .A1(n7761), .A2(n7760), .A3(n7759), .A4(n7758), .ZN(n12130) );
  OR2_X1 U10040 ( .A1(n14299), .A2(n12130), .ZN(n7953) );
  NAND2_X1 U10041 ( .A1(n14299), .A2(n12130), .ZN(n8144) );
  NAND2_X1 U10042 ( .A1(n7953), .A2(n8144), .ZN(n12464) );
  INV_X1 U10043 ( .A(n12130), .ZN(n10873) );
  OR2_X1 U10044 ( .A1(n14299), .A2(n10873), .ZN(n7762) );
  XNOR2_X1 U10045 ( .A(n7764), .B(n7763), .ZN(n8693) );
  NAND2_X1 U10046 ( .A1(n8693), .A2(n7616), .ZN(n7768) );
  NAND2_X1 U10047 ( .A1(n7778), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7765) );
  XNOR2_X1 U10048 ( .A(n7765), .B(P3_IR_REG_14__SCAN_IN), .ZN(n12193) );
  OAI22_X1 U10049 ( .A1(n8073), .A2(SI_14_), .B1(n12193), .B2(n7754), .ZN(
        n7766) );
  INV_X1 U10050 ( .A(n7766), .ZN(n7767) );
  NAND2_X1 U10051 ( .A1(n7768), .A2(n7767), .ZN(n12455) );
  NAND2_X1 U10052 ( .A1(n8055), .A2(P3_REG0_REG_14__SCAN_IN), .ZN(n7774) );
  NAND2_X1 U10053 ( .A1(n8039), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n7773) );
  OAI21_X1 U10054 ( .B1(n7769), .B2(P3_REG3_REG_13__SCAN_IN), .A(
        P3_REG3_REG_14__SCAN_IN), .ZN(n7770) );
  NAND2_X1 U10055 ( .A1(n7770), .A2(n7783), .ZN(n12456) );
  NAND2_X1 U10056 ( .A1(n7625), .A2(n12456), .ZN(n7772) );
  NAND2_X1 U10057 ( .A1(n7556), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n7771) );
  NAND4_X1 U10058 ( .A1(n7774), .A2(n7773), .A3(n7772), .A4(n7771), .ZN(n12439) );
  NAND2_X1 U10059 ( .A1(n12455), .A2(n12439), .ZN(n8148) );
  NAND2_X1 U10060 ( .A1(n8147), .A2(n8148), .ZN(n12451) );
  INV_X1 U10061 ( .A(n12439), .ZN(n11930) );
  INV_X1 U10062 ( .A(n7775), .ZN(n7776) );
  XNOR2_X1 U10063 ( .A(n7777), .B(n7776), .ZN(n8820) );
  NAND2_X1 U10064 ( .A1(n8820), .A2(n7616), .ZN(n7782) );
  OAI21_X1 U10065 ( .B1(n7778), .B2(P3_IR_REG_14__SCAN_IN), .A(
        P3_IR_REG_31__SCAN_IN), .ZN(n7779) );
  XNOR2_X1 U10066 ( .A(n7779), .B(P3_IR_REG_15__SCAN_IN), .ZN(n8310) );
  OAI22_X1 U10067 ( .A1(n8073), .A2(n15194), .B1(n7754), .B2(n12205), .ZN(
        n7780) );
  INV_X1 U10068 ( .A(n7780), .ZN(n7781) );
  AND2_X1 U10069 ( .A1(n7783), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n7784) );
  NOR2_X1 U10070 ( .A1(n7797), .A2(n7784), .ZN(n14287) );
  INV_X1 U10071 ( .A(n14287), .ZN(n12445) );
  NAND2_X1 U10072 ( .A1(n7625), .A2(n12445), .ZN(n7788) );
  NAND2_X1 U10073 ( .A1(n8055), .A2(P3_REG0_REG_15__SCAN_IN), .ZN(n7787) );
  NAND2_X1 U10074 ( .A1(n7556), .A2(P3_REG2_REG_15__SCAN_IN), .ZN(n7786) );
  NAND2_X1 U10075 ( .A1(n8039), .A2(P3_REG1_REG_15__SCAN_IN), .ZN(n7785) );
  NAND4_X1 U10076 ( .A1(n7788), .A2(n7787), .A3(n7786), .A4(n7785), .ZN(n12129) );
  XNOR2_X1 U10077 ( .A(n14275), .B(n12129), .ZN(n12443) );
  NAND2_X1 U10078 ( .A1(n12436), .A2(n7149), .ZN(n7790) );
  NAND2_X1 U10079 ( .A1(n14275), .A2(n12129), .ZN(n7789) );
  INV_X1 U10080 ( .A(n7791), .ZN(n7792) );
  XNOR2_X1 U10081 ( .A(n7793), .B(n7792), .ZN(n8958) );
  NAND2_X1 U10082 ( .A1(n7794), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7795) );
  XNOR2_X1 U10083 ( .A(n7795), .B(P3_IR_REG_16__SCAN_IN), .ZN(n8312) );
  OAI22_X1 U10084 ( .A1(n8073), .A2(n15144), .B1(n7754), .B2(n12222), .ZN(
        n7796) );
  NAND2_X1 U10085 ( .A1(n8055), .A2(P3_REG0_REG_16__SCAN_IN), .ZN(n7802) );
  NAND2_X1 U10086 ( .A1(n8039), .A2(P3_REG1_REG_16__SCAN_IN), .ZN(n7801) );
  NOR2_X1 U10087 ( .A1(n7797), .A2(n15210), .ZN(n7798) );
  OR2_X1 U10088 ( .A1(n7808), .A2(n7798), .ZN(n12431) );
  NAND2_X1 U10089 ( .A1(n7625), .A2(n12431), .ZN(n7800) );
  NAND2_X1 U10090 ( .A1(n7556), .A2(P3_REG2_REG_16__SCAN_IN), .ZN(n7799) );
  NAND4_X1 U10091 ( .A1(n7802), .A2(n7801), .A3(n7800), .A4(n7799), .ZN(n12438) );
  NAND2_X1 U10092 ( .A1(n12579), .A2(n11936), .ZN(n12413) );
  XOR2_X1 U10093 ( .A(n7804), .B(n7803), .Z(n9059) );
  OR2_X1 U10094 ( .A1(n6603), .A2(n7805), .ZN(n7806) );
  XNOR2_X1 U10095 ( .A(n7806), .B(P3_IR_REG_17__SCAN_IN), .ZN(n12247) );
  INV_X1 U10096 ( .A(n12247), .ZN(n9060) );
  OAI22_X1 U10097 ( .A1(n8073), .A2(n15072), .B1(n7754), .B2(n9060), .ZN(n7807) );
  NAND2_X1 U10098 ( .A1(n8055), .A2(P3_REG0_REG_17__SCAN_IN), .ZN(n7813) );
  NAND2_X1 U10099 ( .A1(n8039), .A2(P3_REG1_REG_17__SCAN_IN), .ZN(n7812) );
  OR2_X1 U10100 ( .A1(n7808), .A2(n12063), .ZN(n7809) );
  NAND2_X1 U10101 ( .A1(n7825), .A2(n7809), .ZN(n12420) );
  NAND2_X1 U10102 ( .A1(n7625), .A2(n12420), .ZN(n7811) );
  NAND2_X1 U10103 ( .A1(n7556), .A2(P3_REG2_REG_17__SCAN_IN), .ZN(n7810) );
  NAND4_X1 U10104 ( .A1(n7813), .A2(n7812), .A3(n7811), .A4(n7810), .ZN(n12128) );
  AND2_X1 U10105 ( .A1(n12575), .A2(n12128), .ZN(n8159) );
  INV_X1 U10106 ( .A(n8159), .ZN(n7814) );
  INV_X1 U10107 ( .A(n12575), .ZN(n7816) );
  INV_X1 U10108 ( .A(n12128), .ZN(n11940) );
  NAND2_X1 U10109 ( .A1(n7816), .A2(n11940), .ZN(n8164) );
  NAND2_X1 U10110 ( .A1(n7814), .A2(n8164), .ZN(n12416) );
  AND2_X1 U10111 ( .A1(n12413), .A2(n12416), .ZN(n7815) );
  NAND2_X1 U10112 ( .A1(n7816), .A2(n12128), .ZN(n7817) );
  NAND2_X1 U10113 ( .A1(n12415), .A2(n7817), .ZN(n12401) );
  INV_X1 U10114 ( .A(n7818), .ZN(n7819) );
  XNOR2_X1 U10115 ( .A(n7820), .B(n7819), .ZN(n9133) );
  NAND2_X1 U10116 ( .A1(n9133), .A2(n6488), .ZN(n7824) );
  NAND2_X1 U10117 ( .A1(n7835), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7821) );
  XNOR2_X1 U10118 ( .A(n7821), .B(P3_IR_REG_18__SCAN_IN), .ZN(n12263) );
  OAI22_X1 U10119 ( .A1(n8073), .A2(n9821), .B1(n7754), .B2(n9134), .ZN(n7822)
         );
  INV_X1 U10120 ( .A(n7822), .ZN(n7823) );
  NAND2_X1 U10121 ( .A1(n8055), .A2(P3_REG0_REG_18__SCAN_IN), .ZN(n7830) );
  NAND2_X1 U10122 ( .A1(n8039), .A2(P3_REG1_REG_18__SCAN_IN), .ZN(n7829) );
  NAND2_X1 U10123 ( .A1(n7825), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n7826) );
  NAND2_X1 U10124 ( .A1(n7841), .A2(n7826), .ZN(n12405) );
  NAND2_X1 U10125 ( .A1(n7625), .A2(n12405), .ZN(n7828) );
  NAND2_X1 U10126 ( .A1(n7556), .A2(P3_REG2_REG_18__SCAN_IN), .ZN(n7827) );
  NAND2_X1 U10127 ( .A1(n12088), .A2(n11941), .ZN(n8166) );
  OR2_X1 U10128 ( .A1(n12088), .A2(n12127), .ZN(n7831) );
  INV_X1 U10129 ( .A(n7832), .ZN(n7833) );
  XNOR2_X1 U10130 ( .A(n7834), .B(n7833), .ZN(n9359) );
  NAND2_X1 U10131 ( .A1(n9359), .A2(n7616), .ZN(n7840) );
  NAND2_X1 U10132 ( .A1(n7930), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7837) );
  INV_X1 U10133 ( .A(P3_IR_REG_19__SCAN_IN), .ZN(n7836) );
  OAI22_X1 U10134 ( .A1(n8073), .A2(n15045), .B1(n7754), .B2(n9360), .ZN(n7838) );
  INV_X1 U10135 ( .A(n7838), .ZN(n7839) );
  NAND2_X1 U10136 ( .A1(n8055), .A2(P3_REG0_REG_19__SCAN_IN), .ZN(n7846) );
  NAND2_X1 U10137 ( .A1(n8039), .A2(P3_REG1_REG_19__SCAN_IN), .ZN(n7845) );
  AND2_X1 U10138 ( .A1(n7841), .A2(P3_REG3_REG_19__SCAN_IN), .ZN(n7842) );
  OR2_X1 U10139 ( .A1(n7842), .A2(n7853), .ZN(n12390) );
  NAND2_X1 U10140 ( .A1(n7625), .A2(n12390), .ZN(n7844) );
  NAND2_X1 U10141 ( .A1(n7556), .A2(P3_REG2_REG_19__SCAN_IN), .ZN(n7843) );
  NOR2_X1 U10142 ( .A1(n12518), .A2(n12126), .ZN(n7847) );
  INV_X1 U10143 ( .A(n12518), .ZN(n12392) );
  NOR2_X1 U10144 ( .A1(n7849), .A2(n7848), .ZN(n7850) );
  XNOR2_X1 U10145 ( .A(n7850), .B(P2_DATAO_REG_20__SCAN_IN), .ZN(n9757) );
  NAND2_X1 U10146 ( .A1(n9757), .A2(n7616), .ZN(n7852) );
  NAND2_X1 U10147 ( .A1(n8047), .A2(SI_20_), .ZN(n7851) );
  NAND2_X1 U10148 ( .A1(n8039), .A2(P3_REG1_REG_20__SCAN_IN), .ZN(n7858) );
  NAND2_X1 U10149 ( .A1(n8055), .A2(P3_REG0_REG_20__SCAN_IN), .ZN(n7857) );
  NOR2_X1 U10150 ( .A1(n7853), .A2(n12079), .ZN(n7854) );
  OR2_X1 U10151 ( .A1(n7874), .A2(n7854), .ZN(n12374) );
  NAND2_X1 U10152 ( .A1(n7625), .A2(n12374), .ZN(n7856) );
  NAND2_X1 U10153 ( .A1(n7556), .A2(P3_REG2_REG_20__SCAN_IN), .ZN(n7855) );
  XNOR2_X1 U10154 ( .A(n11947), .B(n11948), .ZN(n12379) );
  NAND2_X1 U10155 ( .A1(n12371), .A2(n12379), .ZN(n7860) );
  NAND2_X1 U10156 ( .A1(n11947), .A2(n12125), .ZN(n7859) );
  NAND2_X1 U10157 ( .A1(n7860), .A2(n7859), .ZN(n12362) );
  XNOR2_X1 U10158 ( .A(n7862), .B(n6814), .ZN(n9763) );
  INV_X1 U10159 ( .A(SI_21_), .ZN(n9761) );
  NOR2_X1 U10160 ( .A1(n8073), .A2(n9761), .ZN(n7863) );
  AOI21_X2 U10161 ( .B1(n9763), .B2(n7616), .A(n7863), .ZN(n12562) );
  NAND2_X1 U10162 ( .A1(n8055), .A2(P3_REG0_REG_21__SCAN_IN), .ZN(n7867) );
  NAND2_X1 U10163 ( .A1(n8039), .A2(P3_REG1_REG_21__SCAN_IN), .ZN(n7866) );
  INV_X1 U10164 ( .A(P3_REG3_REG_21__SCAN_IN), .ZN(n15192) );
  XNOR2_X1 U10165 ( .A(n7874), .B(n15192), .ZN(n12366) );
  NAND2_X1 U10166 ( .A1(n7625), .A2(n12366), .ZN(n7865) );
  NAND2_X1 U10167 ( .A1(n7556), .A2(P3_REG2_REG_21__SCAN_IN), .ZN(n7864) );
  NOR2_X1 U10168 ( .A1(n12562), .A2(n11953), .ZN(n7869) );
  NAND2_X1 U10169 ( .A1(n12562), .A2(n11953), .ZN(n7868) );
  XNOR2_X1 U10170 ( .A(n7871), .B(n7870), .ZN(n9977) );
  NAND2_X1 U10171 ( .A1(n9977), .A2(n7616), .ZN(n7873) );
  NAND2_X1 U10172 ( .A1(n8047), .A2(SI_22_), .ZN(n7872) );
  NAND2_X1 U10173 ( .A1(n8055), .A2(P3_REG0_REG_22__SCAN_IN), .ZN(n7880) );
  NAND2_X1 U10174 ( .A1(n8039), .A2(P3_REG1_REG_22__SCAN_IN), .ZN(n7879) );
  NAND2_X1 U10175 ( .A1(n7874), .A2(n15192), .ZN(n7875) );
  NAND2_X1 U10176 ( .A1(n7875), .A2(P3_REG3_REG_22__SCAN_IN), .ZN(n7876) );
  NAND2_X1 U10177 ( .A1(n7876), .A2(n7887), .ZN(n12356) );
  NAND2_X1 U10178 ( .A1(n7625), .A2(n12356), .ZN(n7878) );
  NAND2_X1 U10179 ( .A1(n7556), .A2(P3_REG2_REG_22__SCAN_IN), .ZN(n7877) );
  NOR2_X1 U10180 ( .A1(n12355), .A2(n12123), .ZN(n7882) );
  NAND2_X1 U10181 ( .A1(n12355), .A2(n12123), .ZN(n7881) );
  XNOR2_X1 U10182 ( .A(n7884), .B(n7883), .ZN(n10387) );
  NAND2_X1 U10183 ( .A1(n10387), .A2(n7616), .ZN(n7886) );
  NAND2_X1 U10184 ( .A1(n8047), .A2(SI_23_), .ZN(n7885) );
  NAND2_X1 U10185 ( .A1(n7887), .A2(P3_REG3_REG_23__SCAN_IN), .ZN(n7888) );
  NAND2_X1 U10186 ( .A1(n7896), .A2(n7888), .ZN(n12342) );
  NAND2_X1 U10187 ( .A1(n12342), .A2(n7625), .ZN(n7892) );
  NAND2_X1 U10188 ( .A1(n8039), .A2(P3_REG1_REG_23__SCAN_IN), .ZN(n7891) );
  NAND2_X1 U10189 ( .A1(n8055), .A2(P3_REG0_REG_23__SCAN_IN), .ZN(n7890) );
  NAND2_X1 U10190 ( .A1(n7556), .A2(P3_REG2_REG_23__SCAN_IN), .ZN(n7889) );
  XNOR2_X1 U10191 ( .A(n12031), .B(n12070), .ZN(n8223) );
  NAND2_X1 U10192 ( .A1(n12031), .A2(n12122), .ZN(n7893) );
  XOR2_X1 U10193 ( .A(n11084), .B(n7894), .Z(n10857) );
  INV_X1 U10194 ( .A(SI_24_), .ZN(n15171) );
  NOR2_X1 U10195 ( .A1(n8073), .A2(n15171), .ZN(n7895) );
  INV_X1 U10196 ( .A(P3_REG1_REG_24__SCAN_IN), .ZN(n7902) );
  NAND2_X1 U10197 ( .A1(n7896), .A2(P3_REG3_REG_24__SCAN_IN), .ZN(n7897) );
  NAND2_X1 U10198 ( .A1(n7908), .A2(n7897), .ZN(n12069) );
  NAND2_X1 U10199 ( .A1(n12069), .A2(n7625), .ZN(n7901) );
  NAND2_X1 U10200 ( .A1(n7556), .A2(P3_REG2_REG_24__SCAN_IN), .ZN(n7899) );
  NAND2_X1 U10201 ( .A1(n8055), .A2(P3_REG0_REG_24__SCAN_IN), .ZN(n7898) );
  AND2_X1 U10202 ( .A1(n7899), .A2(n7898), .ZN(n7900) );
  OAI211_X1 U10203 ( .C1(n7902), .C2(n8058), .A(n7901), .B(n7900), .ZN(n12121)
         );
  INV_X1 U10204 ( .A(n12121), .ZN(n12027) );
  NOR2_X1 U10205 ( .A1(n12499), .A2(n12027), .ZN(n7903) );
  XNOR2_X1 U10206 ( .A(n7905), .B(n7904), .ZN(n10898) );
  NAND2_X1 U10207 ( .A1(n10898), .A2(n7616), .ZN(n7907) );
  NAND2_X1 U10208 ( .A1(n8047), .A2(SI_25_), .ZN(n7906) );
  AND2_X1 U10209 ( .A1(n7908), .A2(P3_REG3_REG_25__SCAN_IN), .ZN(n7909) );
  OR2_X1 U10210 ( .A1(n7909), .A2(n7917), .ZN(n12318) );
  NAND2_X1 U10211 ( .A1(n12318), .A2(n7625), .ZN(n7912) );
  AOI22_X1 U10212 ( .A1(n8055), .A2(P3_REG0_REG_25__SCAN_IN), .B1(n8039), .B2(
        P3_REG1_REG_25__SCAN_IN), .ZN(n7911) );
  NAND2_X1 U10213 ( .A1(n7556), .A2(P3_REG2_REG_25__SCAN_IN), .ZN(n7910) );
  NAND2_X1 U10214 ( .A1(n12317), .A2(n12071), .ZN(n12296) );
  NAND2_X1 U10215 ( .A1(n12317), .A2(n12120), .ZN(n12299) );
  AOI22_X1 U10216 ( .A1(P2_DATAO_REG_26__SCAN_IN), .A2(
        P1_DATAO_REG_26__SCAN_IN), .B1(n6834), .B2(n14125), .ZN(n7913) );
  XNOR2_X1 U10217 ( .A(n7914), .B(n7913), .ZN(n12604) );
  NAND2_X1 U10218 ( .A1(n12604), .A2(n6488), .ZN(n7916) );
  NAND2_X1 U10219 ( .A1(n8047), .A2(SI_26_), .ZN(n7915) );
  XNOR2_X1 U10220 ( .A(n7917), .B(n15206), .ZN(n12305) );
  NAND2_X1 U10221 ( .A1(n12305), .A2(n7625), .ZN(n7922) );
  NAND2_X1 U10222 ( .A1(n7556), .A2(P3_REG2_REG_26__SCAN_IN), .ZN(n7920) );
  NAND2_X1 U10223 ( .A1(n8039), .A2(P3_REG1_REG_26__SCAN_IN), .ZN(n7919) );
  NAND2_X1 U10224 ( .A1(n8055), .A2(P3_REG0_REG_26__SCAN_IN), .ZN(n7918) );
  AND3_X1 U10225 ( .A1(n7920), .A2(n7919), .A3(n7918), .ZN(n7921) );
  NAND2_X1 U10226 ( .A1(n12304), .A2(n12119), .ZN(n7923) );
  AND2_X1 U10227 ( .A1(n12299), .A2(n7923), .ZN(n7925) );
  NAND2_X1 U10228 ( .A1(n12313), .A2(n7925), .ZN(n7924) );
  OR2_X1 U10229 ( .A1(n12304), .A2(n12119), .ZN(n7927) );
  AND2_X1 U10230 ( .A1(n7924), .A2(n7927), .ZN(n7929) );
  OAI21_X2 U10231 ( .B1(n12311), .B2(n12312), .A(n7926), .ZN(n8390) );
  OR2_X1 U10232 ( .A1(n7970), .A2(n7927), .ZN(n8383) );
  NAND2_X1 U10233 ( .A1(n8390), .A2(n8383), .ZN(n7928) );
  AOI21_X1 U10234 ( .B1(n7970), .B2(n7929), .A(n7928), .ZN(n7947) );
  NAND2_X1 U10235 ( .A1(n7999), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7932) );
  NAND2_X1 U10236 ( .A1(n9978), .A2(n8375), .ZN(n8416) );
  INV_X1 U10237 ( .A(n7935), .ZN(n7936) );
  NAND2_X1 U10238 ( .A1(n7936), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7938) );
  NAND2_X1 U10239 ( .A1(n10112), .A2(n8230), .ZN(n8076) );
  INV_X1 U10240 ( .A(P3_REG3_REG_28__SCAN_IN), .ZN(n15066) );
  NOR2_X1 U10241 ( .A1(n7939), .A2(n15066), .ZN(n7940) );
  NAND2_X1 U10242 ( .A1(n8055), .A2(P3_REG0_REG_28__SCAN_IN), .ZN(n7943) );
  NAND2_X1 U10243 ( .A1(n8039), .A2(P3_REG1_REG_28__SCAN_IN), .ZN(n7942) );
  NAND2_X1 U10244 ( .A1(n7556), .A2(P3_REG2_REG_28__SCAN_IN), .ZN(n7941) );
  NAND3_X1 U10245 ( .A1(n7943), .A2(n7942), .A3(n7941), .ZN(n7944) );
  AOI21_X1 U10246 ( .B1(n11976), .B2(n7625), .A(n7944), .ZN(n8407) );
  INV_X1 U10247 ( .A(n8407), .ZN(n12118) );
  INV_X1 U10248 ( .A(n7945), .ZN(n8373) );
  NAND2_X1 U10249 ( .A1(n8373), .A2(n8316), .ZN(n8281) );
  NAND2_X1 U10250 ( .A1(n8281), .A2(n7754), .ZN(n7946) );
  AND2_X2 U10251 ( .A1(n9978), .A2(n10112), .ZN(n8415) );
  INV_X2 U10252 ( .A(n8415), .ZN(n8205) );
  AOI22_X1 U10253 ( .A1(n12118), .A2(n12437), .B1(n12440), .B2(n12119), .ZN(
        n12020) );
  INV_X1 U10254 ( .A(n12144), .ZN(n7948) );
  INV_X1 U10255 ( .A(n14967), .ZN(n7949) );
  NAND2_X1 U10256 ( .A1(n7949), .A2(n8092), .ZN(n9555) );
  NAND2_X1 U10257 ( .A1(n9555), .A2(n8093), .ZN(n10115) );
  NAND2_X1 U10258 ( .A1(n10115), .A2(n10120), .ZN(n10114) );
  NAND2_X1 U10259 ( .A1(n14947), .A2(n14950), .ZN(n14946) );
  NAND2_X1 U10260 ( .A1(n14946), .A2(n8087), .ZN(n10273) );
  NAND2_X1 U10261 ( .A1(n10273), .A2(n10278), .ZN(n10272) );
  NAND2_X1 U10262 ( .A1(n10272), .A2(n8109), .ZN(n10351) );
  NAND2_X1 U10263 ( .A1(n10351), .A2(n10353), .ZN(n10350) );
  NAND2_X1 U10264 ( .A1(n10350), .A2(n8105), .ZN(n14927) );
  NAND2_X1 U10265 ( .A1(n14927), .A2(n14926), .ZN(n14925) );
  NAND2_X1 U10266 ( .A1(n12134), .A2(n10811), .ZN(n8128) );
  NAND2_X1 U10267 ( .A1(n10804), .A2(n8128), .ZN(n7950) );
  INV_X1 U10268 ( .A(n12134), .ZN(n10579) );
  NAND2_X1 U10269 ( .A1(n10579), .A2(n10524), .ZN(n8129) );
  NAND2_X1 U10270 ( .A1(n10861), .A2(n10834), .ZN(n8134) );
  NAND2_X1 U10271 ( .A1(n12132), .A2(n10918), .ZN(n8138) );
  NAND2_X1 U10272 ( .A1(n12474), .A2(n12473), .ZN(n7952) );
  INV_X1 U10273 ( .A(n7953), .ZN(n8145) );
  INV_X1 U10274 ( .A(n12129), .ZN(n11932) );
  NAND2_X1 U10275 ( .A1(n14275), .A2(n11932), .ZN(n8153) );
  NAND2_X1 U10276 ( .A1(n12442), .A2(n8153), .ZN(n12430) );
  AND2_X1 U10277 ( .A1(n12579), .A2(n12438), .ZN(n8158) );
  INV_X1 U10278 ( .A(n8158), .ZN(n7954) );
  INV_X1 U10279 ( .A(n12579), .ZN(n12057) );
  NAND2_X1 U10280 ( .A1(n12057), .A2(n11936), .ZN(n8155) );
  NAND2_X1 U10281 ( .A1(n12430), .A2(n12429), .ZN(n12428) );
  INV_X1 U10282 ( .A(n12416), .ZN(n12411) );
  NAND2_X1 U10283 ( .A1(n12412), .A2(n12411), .ZN(n12410) );
  OR2_X1 U10284 ( .A1(n12518), .A2(n11944), .ZN(n8163) );
  INV_X1 U10285 ( .A(n8163), .ZN(n8170) );
  NAND2_X1 U10286 ( .A1(n12518), .A2(n11944), .ZN(n12377) );
  INV_X1 U10287 ( .A(n12379), .ZN(n7955) );
  AND2_X1 U10288 ( .A1(n12377), .A2(n7955), .ZN(n7956) );
  OR2_X1 U10289 ( .A1(n11947), .A2(n11948), .ZN(n7957) );
  NAND2_X1 U10290 ( .A1(n12376), .A2(n7957), .ZN(n12361) );
  NOR2_X1 U10291 ( .A1(n12562), .A2(n12124), .ZN(n8178) );
  INV_X1 U10292 ( .A(n8178), .ZN(n12347) );
  AND2_X1 U10293 ( .A1(n12347), .A2(n8175), .ZN(n7958) );
  NAND2_X1 U10294 ( .A1(n12361), .A2(n7958), .ZN(n7961) );
  AND2_X1 U10295 ( .A1(n12562), .A2(n12124), .ZN(n8177) );
  INV_X1 U10296 ( .A(n8177), .ZN(n12348) );
  NOR2_X1 U10297 ( .A1(n12355), .A2(n12026), .ZN(n8180) );
  INV_X1 U10298 ( .A(n8180), .ZN(n8176) );
  AND2_X1 U10299 ( .A1(n7959), .A2(n8176), .ZN(n7960) );
  INV_X1 U10300 ( .A(n8223), .ZN(n12335) );
  NAND2_X1 U10301 ( .A1(n12554), .A2(n12122), .ZN(n8188) );
  NAND2_X1 U10302 ( .A1(n12499), .A2(n12121), .ZN(n8189) );
  NAND2_X1 U10303 ( .A1(n12330), .A2(n12027), .ZN(n12295) );
  NAND2_X1 U10304 ( .A1(n12304), .A2(n11968), .ZN(n8194) );
  AND2_X1 U10305 ( .A1(n12296), .A2(n8194), .ZN(n7963) );
  AND2_X1 U10306 ( .A1(n12295), .A2(n7963), .ZN(n7962) );
  NAND2_X1 U10307 ( .A1(n12294), .A2(n7962), .ZN(n7969) );
  INV_X1 U10308 ( .A(n7963), .ZN(n7964) );
  AND2_X1 U10309 ( .A1(n7969), .A2(n7966), .ZN(n7965) );
  AND2_X1 U10310 ( .A1(n7970), .A2(n8196), .ZN(n7967) );
  NAND2_X1 U10311 ( .A1(n7969), .A2(n7968), .ZN(n8397) );
  OAI21_X1 U10312 ( .B1(n7971), .B2(n7970), .A(n8397), .ZN(n12287) );
  NAND2_X1 U10313 ( .A1(n9978), .A2(n9758), .ZN(n7972) );
  NAND2_X1 U10314 ( .A1(n7972), .A2(n8375), .ZN(n7973) );
  NAND2_X1 U10315 ( .A1(n7973), .A2(n8231), .ZN(n7976) );
  NOR2_X1 U10316 ( .A1(n10112), .A2(n8230), .ZN(n7974) );
  OR2_X1 U10317 ( .A1(n7974), .A2(n9978), .ZN(n7975) );
  NAND2_X1 U10318 ( .A1(n7976), .A2(n7975), .ZN(n9513) );
  AND2_X1 U10319 ( .A1(n14298), .A2(n9547), .ZN(n7977) );
  NAND2_X1 U10320 ( .A1(n9513), .A2(n7977), .ZN(n7980) );
  NOR2_X1 U10321 ( .A1(n9758), .A2(n8375), .ZN(n7978) );
  AND2_X1 U10322 ( .A1(n9978), .A2(n7978), .ZN(n8018) );
  INV_X1 U10323 ( .A(n8018), .ZN(n7979) );
  NAND2_X1 U10324 ( .A1(n9758), .A2(n8375), .ZN(n14969) );
  NOR2_X1 U10325 ( .A1(n12291), .A2(n7981), .ZN(n12538) );
  NAND2_X1 U10326 ( .A1(n6510), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7982) );
  NAND2_X1 U10327 ( .A1(n7983), .A2(n7539), .ZN(n12605) );
  INV_X1 U10328 ( .A(n12605), .ZN(n7992) );
  NAND2_X1 U10329 ( .A1(n6511), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7984) );
  MUX2_X1 U10330 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7984), .S(
        P3_IR_REG_25__SCAN_IN), .Z(n7985) );
  INV_X1 U10331 ( .A(n7986), .ZN(n7987) );
  NAND2_X1 U10332 ( .A1(n7987), .A2(P3_IR_REG_31__SCAN_IN), .ZN(n7988) );
  MUX2_X1 U10333 ( .A(P3_IR_REG_31__SCAN_IN), .B(n7988), .S(
        P3_IR_REG_24__SCAN_IN), .Z(n7989) );
  NAND2_X1 U10334 ( .A1(n7989), .A2(n6511), .ZN(n10855) );
  XNOR2_X1 U10335 ( .A(n10855), .B(P3_B_REG_SCAN_IN), .ZN(n7990) );
  NAND2_X1 U10336 ( .A1(n10899), .A2(n7990), .ZN(n7991) );
  INV_X1 U10337 ( .A(P3_D_REG_1__SCAN_IN), .ZN(n7993) );
  NAND2_X1 U10338 ( .A1(n8787), .A2(n7993), .ZN(n7995) );
  NAND2_X1 U10339 ( .A1(n12605), .A2(n10899), .ZN(n7994) );
  INV_X1 U10340 ( .A(P3_D_REG_0__SCAN_IN), .ZN(n7996) );
  NAND2_X1 U10341 ( .A1(n8787), .A2(n7996), .ZN(n7998) );
  NAND2_X1 U10342 ( .A1(n12605), .A2(n10855), .ZN(n7997) );
  NAND2_X1 U10343 ( .A1(n12585), .A2(n12587), .ZN(n8412) );
  INV_X1 U10344 ( .A(n10855), .ZN(n8001) );
  NAND2_X1 U10345 ( .A1(n8002), .A2(n8001), .ZN(n8003) );
  INV_X1 U10346 ( .A(n8787), .ZN(n8015) );
  NOR2_X1 U10347 ( .A1(P3_D_REG_17__SCAN_IN), .A2(P3_D_REG_22__SCAN_IN), .ZN(
        n8007) );
  NOR4_X1 U10348 ( .A1(P3_D_REG_2__SCAN_IN), .A2(P3_D_REG_8__SCAN_IN), .A3(
        P3_D_REG_25__SCAN_IN), .A4(P3_D_REG_20__SCAN_IN), .ZN(n8006) );
  NOR4_X1 U10349 ( .A1(P3_D_REG_29__SCAN_IN), .A2(P3_D_REG_10__SCAN_IN), .A3(
        P3_D_REG_31__SCAN_IN), .A4(P3_D_REG_14__SCAN_IN), .ZN(n8005) );
  NOR4_X1 U10350 ( .A1(P3_D_REG_19__SCAN_IN), .A2(P3_D_REG_18__SCAN_IN), .A3(
        P3_D_REG_27__SCAN_IN), .A4(P3_D_REG_24__SCAN_IN), .ZN(n8004) );
  NAND4_X1 U10351 ( .A1(n8007), .A2(n8006), .A3(n8005), .A4(n8004), .ZN(n8013)
         );
  NOR4_X1 U10352 ( .A1(P3_D_REG_9__SCAN_IN), .A2(P3_D_REG_16__SCAN_IN), .A3(
        P3_D_REG_15__SCAN_IN), .A4(P3_D_REG_30__SCAN_IN), .ZN(n8011) );
  NOR4_X1 U10353 ( .A1(P3_D_REG_11__SCAN_IN), .A2(P3_D_REG_21__SCAN_IN), .A3(
        P3_D_REG_12__SCAN_IN), .A4(P3_D_REG_26__SCAN_IN), .ZN(n8010) );
  NOR4_X1 U10354 ( .A1(P3_D_REG_3__SCAN_IN), .A2(P3_D_REG_5__SCAN_IN), .A3(
        P3_D_REG_4__SCAN_IN), .A4(P3_D_REG_7__SCAN_IN), .ZN(n8009) );
  NOR4_X1 U10355 ( .A1(P3_D_REG_13__SCAN_IN), .A2(P3_D_REG_28__SCAN_IN), .A3(
        P3_D_REG_23__SCAN_IN), .A4(P3_D_REG_6__SCAN_IN), .ZN(n8008) );
  NAND4_X1 U10356 ( .A1(n8011), .A2(n8010), .A3(n8009), .A4(n8008), .ZN(n8012)
         );
  NOR2_X1 U10357 ( .A1(n8013), .A2(n8012), .ZN(n8014) );
  NOR2_X1 U10358 ( .A1(n9509), .A2(n8417), .ZN(n8017) );
  INV_X1 U10359 ( .A(n12587), .ZN(n8016) );
  NAND2_X1 U10360 ( .A1(n8021), .A2(n8016), .ZN(n8418) );
  OR2_X1 U10361 ( .A1(n8415), .A2(n8018), .ZN(n9883) );
  NAND2_X1 U10362 ( .A1(n8415), .A2(n9508), .ZN(n9886) );
  AND2_X1 U10363 ( .A1(n9883), .A2(n9886), .ZN(n8023) );
  NAND2_X1 U10364 ( .A1(n9978), .A2(n9360), .ZN(n8019) );
  OAI21_X1 U10365 ( .B1(n14298), .B2(n8230), .A(n8019), .ZN(n8020) );
  AOI21_X1 U10366 ( .B1(n8020), .B2(n9508), .A(n8415), .ZN(n8022) );
  MUX2_X1 U10367 ( .A(n8023), .B(n8022), .S(n8021), .Z(n8024) );
  MUX2_X1 U10368 ( .A(n8025), .B(n12538), .S(n15038), .Z(n8026) );
  INV_X1 U10369 ( .A(n12022), .ZN(n12541) );
  NAND2_X1 U10370 ( .A1(n8026), .A2(n7475), .ZN(P3_U3486) );
  NOR2_X1 U10371 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n14123), .ZN(n8028) );
  INV_X1 U10372 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n11180) );
  INV_X1 U10373 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n11618) );
  AOI22_X1 U10374 ( .A1(P2_DATAO_REG_28__SCAN_IN), .A2(n11180), .B1(
        P1_DATAO_REG_28__SCAN_IN), .B2(n11618), .ZN(n8029) );
  INV_X1 U10375 ( .A(n8029), .ZN(n8030) );
  XNOR2_X1 U10376 ( .A(n8035), .B(n8030), .ZN(n12599) );
  NAND2_X1 U10377 ( .A1(n12599), .A2(n6488), .ZN(n8032) );
  NAND2_X1 U10378 ( .A1(n8047), .A2(SI_28_), .ZN(n8031) );
  NAND2_X2 U10379 ( .A1(n8032), .A2(n8031), .ZN(n12282) );
  NAND2_X1 U10380 ( .A1(n12282), .A2(n8407), .ZN(n8199) );
  NAND2_X1 U10381 ( .A1(n12022), .A2(n11973), .ZN(n8396) );
  NAND2_X1 U10382 ( .A1(n8199), .A2(n8396), .ZN(n8082) );
  INV_X1 U10383 ( .A(n8082), .ZN(n8033) );
  NAND2_X1 U10384 ( .A1(n8397), .A2(n8033), .ZN(n8034) );
  OR2_X2 U10385 ( .A1(n12282), .A2(n8407), .ZN(n8200) );
  NAND2_X1 U10386 ( .A1(n8034), .A2(n8200), .ZN(n8411) );
  INV_X1 U10387 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n11186) );
  INV_X1 U10388 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n11189) );
  OAI22_X1 U10389 ( .A1(n11186), .A2(P1_DATAO_REG_29__SCAN_IN), .B1(n11189), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n8044) );
  INV_X1 U10390 ( .A(n8044), .ZN(n8036) );
  NAND2_X1 U10391 ( .A1(n12597), .A2(n7616), .ZN(n8038) );
  NAND2_X1 U10392 ( .A1(n8047), .A2(SI_29_), .ZN(n8037) );
  NAND2_X1 U10393 ( .A1(n8038), .A2(n8037), .ZN(n8423) );
  NAND2_X1 U10394 ( .A1(n12273), .A2(n7625), .ZN(n8061) );
  NAND2_X1 U10395 ( .A1(n8055), .A2(P3_REG0_REG_29__SCAN_IN), .ZN(n8042) );
  NAND2_X1 U10396 ( .A1(n8039), .A2(P3_REG1_REG_29__SCAN_IN), .ZN(n8041) );
  NAND2_X1 U10397 ( .A1(n7556), .A2(P3_REG2_REG_29__SCAN_IN), .ZN(n8040) );
  AND3_X1 U10398 ( .A1(n8042), .A2(n8041), .A3(n8040), .ZN(n8043) );
  NOR2_X1 U10399 ( .A1(n8423), .A2(n9376), .ZN(n8086) );
  OAI22_X1 U10400 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n11189), .B1(n8045), 
        .B2(n8044), .ZN(n8069) );
  INV_X1 U10401 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n11990) );
  INV_X1 U10402 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n14117) );
  AOI22_X1 U10403 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(
        P1_DATAO_REG_30__SCAN_IN), .B1(n11990), .B2(n14117), .ZN(n8046) );
  XNOR2_X1 U10404 ( .A(n8069), .B(n8046), .ZN(n12014) );
  NAND2_X1 U10405 ( .A1(n12014), .A2(n7616), .ZN(n8049) );
  NAND2_X1 U10406 ( .A1(n8047), .A2(SI_30_), .ZN(n8048) );
  INV_X1 U10407 ( .A(n14292), .ZN(n8063) );
  INV_X1 U10408 ( .A(P3_REG2_REG_30__SCAN_IN), .ZN(n8052) );
  NAND2_X1 U10409 ( .A1(n8055), .A2(P3_REG0_REG_30__SCAN_IN), .ZN(n8051) );
  NAND2_X1 U10410 ( .A1(n6513), .A2(P3_REG1_REG_30__SCAN_IN), .ZN(n8050) );
  OAI211_X1 U10411 ( .C1(n8052), .C2(n7585), .A(n8051), .B(n8050), .ZN(n8053)
         );
  INV_X1 U10412 ( .A(n8053), .ZN(n8054) );
  NAND2_X1 U10413 ( .A1(n8061), .A2(n8054), .ZN(n12117) );
  INV_X1 U10414 ( .A(n12117), .ZN(n8406) );
  NAND2_X1 U10415 ( .A1(n8063), .A2(n8406), .ZN(n8204) );
  INV_X1 U10416 ( .A(P3_REG1_REG_31__SCAN_IN), .ZN(n14290) );
  NAND2_X1 U10417 ( .A1(n7556), .A2(P3_REG2_REG_31__SCAN_IN), .ZN(n8057) );
  NAND2_X1 U10418 ( .A1(n8055), .A2(P3_REG0_REG_31__SCAN_IN), .ZN(n8056) );
  OAI211_X1 U10419 ( .C1(n14290), .C2(n8058), .A(n8057), .B(n8056), .ZN(n8059)
         );
  INV_X1 U10420 ( .A(n8059), .ZN(n8060) );
  NAND2_X1 U10421 ( .A1(n8061), .A2(n8060), .ZN(n12267) );
  INV_X1 U10422 ( .A(n12267), .ZN(n8062) );
  NAND2_X1 U10423 ( .A1(n8063), .A2(n8062), .ZN(n8064) );
  NAND2_X1 U10424 ( .A1(n8204), .A2(n8064), .ZN(n8065) );
  NOR2_X1 U10425 ( .A1(n8085), .A2(n8065), .ZN(n8066) );
  NAND2_X1 U10426 ( .A1(P2_DATAO_REG_30__SCAN_IN), .A2(n11990), .ZN(n8068) );
  AOI22_X1 U10427 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n14117), .B1(n8069), 
        .B2(n8068), .ZN(n8072) );
  INV_X1 U10428 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n8070) );
  INV_X1 U10429 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n8709) );
  AOI22_X1 U10430 ( .A1(P2_DATAO_REG_31__SCAN_IN), .A2(
        P1_DATAO_REG_31__SCAN_IN), .B1(n8070), .B2(n8709), .ZN(n8071) );
  XOR2_X1 U10431 ( .A(n8072), .B(n8071), .Z(n12592) );
  NOR2_X1 U10432 ( .A1(n8073), .A2(n15074), .ZN(n8074) );
  AND2_X1 U10433 ( .A1(n12267), .A2(n8375), .ZN(n8077) );
  NAND2_X1 U10434 ( .A1(n14292), .A2(n12117), .ZN(n8203) );
  AOI22_X1 U10435 ( .A1(n14288), .A2(n8375), .B1(n8077), .B2(n8203), .ZN(n8080) );
  AOI211_X1 U10436 ( .C1(n12267), .C2(n8203), .A(n8375), .B(n14288), .ZN(n8075) );
  AOI211_X1 U10437 ( .C1(n8077), .C2(n14288), .A(n8076), .B(n8075), .ZN(n8079)
         );
  NAND2_X1 U10438 ( .A1(n14288), .A2(n12267), .ZN(n8228) );
  NAND3_X1 U10439 ( .A1(n8081), .A2(n9360), .A3(n8228), .ZN(n8078) );
  OAI211_X1 U10440 ( .C1(n8081), .C2(n8080), .A(n8079), .B(n8078), .ZN(n8236)
         );
  NAND2_X1 U10441 ( .A1(n8082), .A2(n8200), .ZN(n8083) );
  MUX2_X1 U10442 ( .A(n8083), .B(n8200), .S(n8205), .Z(n8084) );
  AND2_X1 U10443 ( .A1(n8207), .A2(n8084), .ZN(n8202) );
  MUX2_X1 U10444 ( .A(n8086), .B(n8085), .S(n8205), .Z(n8201) );
  INV_X1 U10445 ( .A(n14275), .ZN(n12584) );
  AOI21_X1 U10446 ( .B1(n12584), .B2(n12129), .A(n8158), .ZN(n8152) );
  INV_X1 U10447 ( .A(n8087), .ZN(n8102) );
  INV_X1 U10448 ( .A(n9522), .ZN(n10108) );
  NAND2_X1 U10449 ( .A1(n12144), .A2(n10108), .ZN(n8208) );
  AOI211_X1 U10450 ( .C1(n10112), .C2(n8208), .A(n8415), .B(n9551), .ZN(n8091)
         );
  INV_X1 U10451 ( .A(n8208), .ZN(n8089) );
  INV_X1 U10452 ( .A(n9978), .ZN(n8088) );
  NOR3_X1 U10453 ( .A1(n14966), .A2(n8089), .A3(n8088), .ZN(n8090) );
  OAI22_X1 U10454 ( .A1(n8091), .A2(n8090), .B1(n10112), .B2(n14967), .ZN(
        n8095) );
  MUX2_X1 U10455 ( .A(n8093), .B(n8092), .S(n8205), .Z(n8094) );
  INV_X1 U10456 ( .A(n8096), .ZN(n8097) );
  OAI21_X1 U10457 ( .B1(n8102), .B2(n8097), .A(n8205), .ZN(n8098) );
  INV_X1 U10458 ( .A(n8103), .ZN(n8104) );
  NOR3_X1 U10459 ( .A1(n8112), .A2(n8104), .A3(n8110), .ZN(n8108) );
  INV_X1 U10460 ( .A(n8105), .ZN(n8106) );
  NOR3_X1 U10461 ( .A1(n8108), .A2(n8107), .A3(n8106), .ZN(n8118) );
  INV_X1 U10462 ( .A(n8109), .ZN(n8111) );
  NOR3_X1 U10463 ( .A1(n8112), .A2(n8111), .A3(n8110), .ZN(n8116) );
  NAND2_X1 U10464 ( .A1(n8119), .A2(n8113), .ZN(n8115) );
  OAI21_X1 U10465 ( .B1(n8116), .B2(n8115), .A(n8114), .ZN(n8117) );
  MUX2_X1 U10466 ( .A(n8118), .B(n8117), .S(n8205), .Z(n8124) );
  OAI21_X1 U10467 ( .B1(n8205), .B2(n8119), .A(n14912), .ZN(n8123) );
  MUX2_X1 U10468 ( .A(n8121), .B(n8120), .S(n8205), .Z(n8122) );
  MUX2_X1 U10469 ( .A(n8126), .B(n8125), .S(n8205), .Z(n8127) );
  MUX2_X1 U10470 ( .A(n8129), .B(n8128), .S(n8205), .Z(n8130) );
  MUX2_X1 U10471 ( .A(n8132), .B(n8131), .S(n8205), .Z(n8133) );
  NAND2_X1 U10472 ( .A1(n8133), .A2(n10917), .ZN(n8137) );
  INV_X1 U10473 ( .A(n8134), .ZN(n8135) );
  OAI21_X1 U10474 ( .B1(n8143), .B2(n8135), .A(n8205), .ZN(n8136) );
  AOI21_X1 U10475 ( .B1(n8140), .B2(n8138), .A(n8205), .ZN(n8139) );
  AOI21_X1 U10476 ( .B1(n8141), .B2(n8140), .A(n8139), .ZN(n8142) );
  MUX2_X1 U10477 ( .A(n7155), .B(n8145), .S(n8205), .Z(n8146) );
  INV_X1 U10478 ( .A(n8147), .ZN(n8150) );
  INV_X1 U10479 ( .A(n8148), .ZN(n8149) );
  MUX2_X1 U10480 ( .A(n8150), .B(n8149), .S(n8205), .Z(n8151) );
  AOI21_X1 U10481 ( .B1(n8155), .B2(n8153), .A(n8205), .ZN(n8154) );
  AOI21_X1 U10482 ( .B1(n8156), .B2(n8155), .A(n8154), .ZN(n8157) );
  AOI21_X1 U10483 ( .B1(n8158), .B2(n8415), .A(n8157), .ZN(n8165) );
  NAND2_X1 U10484 ( .A1(n8166), .A2(n8159), .ZN(n8161) );
  AND3_X1 U10485 ( .A1(n8161), .A2(n8415), .A3(n8160), .ZN(n8162) );
  AND2_X1 U10486 ( .A1(n8163), .A2(n8162), .ZN(n8167) );
  NAND3_X1 U10487 ( .A1(n12377), .A2(n8205), .A3(n8166), .ZN(n8169) );
  INV_X1 U10488 ( .A(n8167), .ZN(n8168) );
  INV_X1 U10489 ( .A(n12377), .ZN(n8171) );
  MUX2_X1 U10490 ( .A(n8171), .B(n8170), .S(n8205), .Z(n8172) );
  XNOR2_X1 U10491 ( .A(n12562), .B(n11953), .ZN(n12363) );
  NAND3_X1 U10492 ( .A1(n11947), .A2(n11948), .A3(n8205), .ZN(n8174) );
  INV_X1 U10493 ( .A(n11947), .ZN(n12566) );
  NAND3_X1 U10494 ( .A1(n12566), .A2(n8415), .A3(n12125), .ZN(n8173) );
  NAND2_X1 U10495 ( .A1(n8176), .A2(n8175), .ZN(n12352) );
  MUX2_X1 U10496 ( .A(n8178), .B(n8177), .S(n8205), .Z(n8179) );
  NOR2_X1 U10497 ( .A1(n12352), .A2(n8179), .ZN(n8183) );
  MUX2_X1 U10498 ( .A(n8181), .B(n8180), .S(n8415), .Z(n8182) );
  AOI211_X1 U10499 ( .C1(n8184), .C2(n8183), .A(n8182), .B(n8223), .ZN(n8186)
         );
  NOR3_X1 U10500 ( .A1(n12554), .A2(n12122), .A3(n8205), .ZN(n8185) );
  OAI21_X1 U10501 ( .B1(n8186), .B2(n8185), .A(n12326), .ZN(n8187) );
  NAND2_X1 U10502 ( .A1(n8187), .A2(n12312), .ZN(n8192) );
  AOI21_X1 U10503 ( .B1(n8189), .B2(n8188), .A(n8415), .ZN(n8190) );
  MUX2_X1 U10504 ( .A(n8415), .B(n8190), .S(n12295), .Z(n8191) );
  NAND2_X1 U10505 ( .A1(n8196), .A2(n8194), .ZN(n12300) );
  INV_X1 U10506 ( .A(n8193), .ZN(n8195) );
  INV_X1 U10507 ( .A(n12296), .ZN(n8197) );
  AND2_X2 U10508 ( .A1(n8200), .A2(n8199), .ZN(n11974) );
  AND2_X1 U10509 ( .A1(n8203), .A2(n8204), .ZN(n8227) );
  NOR2_X1 U10510 ( .A1(n14288), .A2(n12267), .ZN(n8224) );
  NAND2_X1 U10511 ( .A1(n8237), .A2(n9547), .ZN(n8235) );
  NAND4_X1 U10512 ( .A1(n8207), .A2(n11974), .A3(n12312), .A4(n8206), .ZN(
        n8222) );
  AND2_X1 U10513 ( .A1(n14967), .A2(n8208), .ZN(n9519) );
  NAND4_X1 U10514 ( .A1(n10353), .A2(n14912), .A3(n10632), .A4(n9519), .ZN(
        n8209) );
  NOR2_X1 U10515 ( .A1(n8209), .A2(n14898), .ZN(n8215) );
  NAND3_X1 U10516 ( .A1(n10278), .A2(n10120), .A3(n14926), .ZN(n8212) );
  INV_X1 U10517 ( .A(n14966), .ZN(n8210) );
  NAND2_X1 U10518 ( .A1(n8210), .A2(n14950), .ZN(n8211) );
  NOR2_X1 U10519 ( .A1(n8212), .A2(n8211), .ZN(n8214) );
  NAND4_X1 U10520 ( .A1(n8215), .A2(n8214), .A3(n8213), .A4(n10917), .ZN(n8216) );
  NOR2_X1 U10521 ( .A1(n8216), .A2(n12480), .ZN(n8217) );
  NAND2_X1 U10522 ( .A1(n6840), .A2(n8217), .ZN(n8218) );
  NOR2_X1 U10523 ( .A1(n12451), .A2(n8218), .ZN(n8219) );
  NAND4_X1 U10524 ( .A1(n12411), .A2(n12429), .A3(n8219), .A4(n12443), .ZN(
        n8220) );
  XNOR2_X1 U10525 ( .A(n12518), .B(n12126), .ZN(n12387) );
  NAND4_X1 U10526 ( .A1(n12326), .A2(n6495), .A3(n12387), .A4(n12363), .ZN(
        n8221) );
  INV_X1 U10527 ( .A(n8224), .ZN(n8225) );
  NAND4_X1 U10528 ( .A1(n8228), .A2(n8227), .A3(n8226), .A4(n8225), .ZN(n8229)
         );
  INV_X1 U10529 ( .A(n9546), .ZN(n8232) );
  NAND3_X1 U10530 ( .A1(n8236), .A2(n8235), .A3(n8234), .ZN(n8239) );
  NOR2_X1 U10531 ( .A1(n8237), .A2(n14969), .ZN(n8238) );
  AND2_X1 U10532 ( .A1(n9495), .A2(P3_STATE_REG_SCAN_IN), .ZN(n8240) );
  OAI21_X1 U10533 ( .B1(n8239), .B2(n8238), .A(n8240), .ZN(n8244) );
  NOR4_X1 U10534 ( .A1(n12103), .A2(n7945), .A3(n9509), .A4(n9508), .ZN(n8242)
         );
  INV_X1 U10535 ( .A(n8240), .ZN(n10388) );
  OAI21_X1 U10536 ( .B1(n10388), .B2(n9978), .A(P3_B_REG_SCAN_IN), .ZN(n8241)
         );
  OR2_X1 U10537 ( .A1(n8242), .A2(n8241), .ZN(n8243) );
  NAND2_X1 U10538 ( .A1(n8244), .A2(n8243), .ZN(P3_U3296) );
  INV_X1 U10539 ( .A(n9496), .ZN(n8245) );
  INV_X1 U10540 ( .A(P3_REG2_REG_17__SCAN_IN), .ZN(n12233) );
  INV_X1 U10541 ( .A(P3_REG2_REG_15__SCAN_IN), .ZN(n12199) );
  INV_X1 U10542 ( .A(n14877), .ZN(n8346) );
  INV_X1 U10543 ( .A(P3_IR_REG_0__SCAN_IN), .ZN(n8551) );
  NAND2_X1 U10544 ( .A1(n8247), .A2(P3_REG2_REG_0__SCAN_IN), .ZN(n8246) );
  OAI21_X1 U10545 ( .B1(P3_REG2_REG_2__SCAN_IN), .B2(n9058), .A(n8248), .ZN(
        n9051) );
  NOR2_X1 U10546 ( .A1(n9052), .A2(n9051), .ZN(n9050) );
  NOR2_X1 U10547 ( .A1(n9072), .A2(n8250), .ZN(n8251) );
  INV_X1 U10548 ( .A(P3_REG2_REG_3__SCAN_IN), .ZN(n9064) );
  NAND2_X1 U10549 ( .A1(P3_REG2_REG_4__SCAN_IN), .A2(n9185), .ZN(n8252) );
  OAI21_X1 U10550 ( .B1(P3_REG2_REG_4__SCAN_IN), .B2(n9185), .A(n8252), .ZN(
        n9179) );
  NOR2_X1 U10551 ( .A1(n9398), .A2(n8253), .ZN(n8254) );
  INV_X1 U10552 ( .A(P3_REG2_REG_5__SCAN_IN), .ZN(n9393) );
  XNOR2_X1 U10553 ( .A(n8253), .B(n9398), .ZN(n9392) );
  NAND2_X1 U10554 ( .A1(P3_REG2_REG_6__SCAN_IN), .A2(n8620), .ZN(n8255) );
  OAI21_X1 U10555 ( .B1(P3_REG2_REG_6__SCAN_IN), .B2(n8620), .A(n8255), .ZN(
        n14819) );
  NOR2_X1 U10556 ( .A1(n8321), .A2(n8256), .ZN(n8257) );
  INV_X1 U10557 ( .A(P3_REG2_REG_7__SCAN_IN), .ZN(n9896) );
  XNOR2_X1 U10558 ( .A(n8256), .B(n8321), .ZN(n9895) );
  NAND2_X1 U10559 ( .A1(P3_REG2_REG_8__SCAN_IN), .A2(n8624), .ZN(n8258) );
  OAI21_X1 U10560 ( .B1(P3_REG2_REG_8__SCAN_IN), .B2(n8624), .A(n8258), .ZN(
        n14838) );
  NOR2_X1 U10561 ( .A1(n14839), .A2(n14838), .ZN(n14837) );
  NOR2_X1 U10562 ( .A1(n6680), .A2(n8259), .ZN(n8260) );
  INV_X1 U10563 ( .A(P3_REG2_REG_9__SCAN_IN), .ZN(n10333) );
  NOR2_X1 U10564 ( .A1(n10333), .A2(n10332), .ZN(n10331) );
  NAND2_X1 U10565 ( .A1(P3_REG2_REG_10__SCAN_IN), .A2(n14866), .ZN(n8261) );
  OAI21_X1 U10566 ( .B1(P3_REG2_REG_10__SCAN_IN), .B2(n14866), .A(n8261), .ZN(
        n14855) );
  NOR2_X1 U10567 ( .A1(n8346), .A2(n8262), .ZN(n8263) );
  INV_X1 U10568 ( .A(P3_REG2_REG_11__SCAN_IN), .ZN(n14874) );
  AOI22_X1 U10569 ( .A1(P3_REG2_REG_12__SCAN_IN), .A2(n8350), .B1(n12158), 
        .B2(n8264), .ZN(n12146) );
  NOR2_X1 U10570 ( .A1(n8266), .A2(n8267), .ZN(n8268) );
  INV_X1 U10571 ( .A(P3_REG2_REG_13__SCAN_IN), .ZN(n12166) );
  NOR2_X1 U10572 ( .A1(n12166), .A2(n12165), .ZN(n12164) );
  NOR2_X1 U10573 ( .A1(n8268), .A2(n12164), .ZN(n12182) );
  NAND2_X1 U10574 ( .A1(n8692), .A2(P3_REG2_REG_14__SCAN_IN), .ZN(n8356) );
  OAI21_X1 U10575 ( .B1(n8692), .B2(P3_REG2_REG_14__SCAN_IN), .A(n8356), .ZN(
        n12181) );
  NOR2_X1 U10576 ( .A1(n12182), .A2(n12181), .ZN(n12180) );
  INV_X1 U10577 ( .A(n12180), .ZN(n8269) );
  AND2_X1 U10578 ( .A1(n12205), .A2(n8270), .ZN(n8271) );
  INV_X1 U10579 ( .A(P3_REG2_REG_16__SCAN_IN), .ZN(n8272) );
  AOI22_X1 U10580 ( .A1(P3_REG2_REG_16__SCAN_IN), .A2(n8312), .B1(n12222), 
        .B2(n8272), .ZN(n12215) );
  NAND2_X1 U10581 ( .A1(P3_REG2_REG_18__SCAN_IN), .A2(n9134), .ZN(n8275) );
  OAI21_X1 U10582 ( .B1(P3_REG2_REG_18__SCAN_IN), .B2(n9134), .A(n8275), .ZN(
        n12251) );
  INV_X1 U10583 ( .A(n8275), .ZN(n8276) );
  NOR2_X1 U10584 ( .A1(n12250), .A2(n8276), .ZN(n8278) );
  INV_X1 U10585 ( .A(P3_REG2_REG_19__SCAN_IN), .ZN(n8277) );
  MUX2_X1 U10586 ( .A(P3_REG2_REG_19__SCAN_IN), .B(n8277), .S(n9360), .Z(n8367) );
  XNOR2_X1 U10587 ( .A(n8278), .B(n8367), .ZN(n8283) );
  NAND2_X1 U10588 ( .A1(n10388), .A2(n9509), .ZN(n8371) );
  NAND2_X1 U10589 ( .A1(n8279), .A2(n8415), .ZN(n8280) );
  AND2_X1 U10590 ( .A1(n8280), .A2(n7754), .ZN(n8370) );
  AND2_X1 U10591 ( .A1(n8371), .A2(n8370), .ZN(n8374) );
  INV_X1 U10592 ( .A(n8281), .ZN(n8282) );
  INV_X1 U10593 ( .A(P3_REG1_REG_7__SCAN_IN), .ZN(n15030) );
  NAND2_X1 U10594 ( .A1(P3_REG1_REG_0__SCAN_IN), .A2(n8551), .ZN(n8284) );
  NOR2_X1 U10595 ( .A1(P3_IR_REG_1__SCAN_IN), .A2(n8284), .ZN(n8286) );
  INV_X1 U10596 ( .A(P3_REG1_REG_1__SCAN_IN), .ZN(n15022) );
  INV_X1 U10597 ( .A(n8285), .ZN(n9219) );
  OAI21_X1 U10598 ( .B1(P3_REG1_REG_2__SCAN_IN), .B2(n9058), .A(n8287), .ZN(
        n9045) );
  NOR2_X1 U10599 ( .A1(n9072), .A2(n8288), .ZN(n8289) );
  INV_X1 U10600 ( .A(P3_REG1_REG_3__SCAN_IN), .ZN(n15026) );
  NAND2_X1 U10601 ( .A1(P3_REG1_REG_4__SCAN_IN), .A2(n9185), .ZN(n8290) );
  OAI21_X1 U10602 ( .B1(P3_REG1_REG_4__SCAN_IN), .B2(n9185), .A(n8290), .ZN(
        n9175) );
  NOR2_X1 U10603 ( .A1(n9398), .A2(n8291), .ZN(n8292) );
  INV_X1 U10604 ( .A(P3_REG1_REG_5__SCAN_IN), .ZN(n9387) );
  NAND2_X1 U10605 ( .A1(P3_REG1_REG_6__SCAN_IN), .A2(n8620), .ZN(n8293) );
  OAI21_X1 U10606 ( .B1(P3_REG1_REG_6__SCAN_IN), .B2(n8620), .A(n8293), .ZN(
        n14817) );
  XNOR2_X1 U10607 ( .A(n8295), .B(n8321), .ZN(n9903) );
  NOR2_X1 U10608 ( .A1(n15030), .A2(n9903), .ZN(n9902) );
  NOR2_X1 U10609 ( .A1(n8321), .A2(n8295), .ZN(n8296) );
  NOR2_X1 U10610 ( .A1(n9902), .A2(n8296), .ZN(n14836) );
  NAND2_X1 U10611 ( .A1(P3_REG1_REG_8__SCAN_IN), .A2(n8624), .ZN(n8297) );
  OAI21_X1 U10612 ( .B1(P3_REG1_REG_8__SCAN_IN), .B2(n8624), .A(n8297), .ZN(
        n14835) );
  NOR2_X1 U10613 ( .A1(n14836), .A2(n14835), .ZN(n14834) );
  INV_X1 U10614 ( .A(n8297), .ZN(n8298) );
  NOR2_X1 U10615 ( .A1(n6680), .A2(n8299), .ZN(n8301) );
  INV_X1 U10616 ( .A(P3_REG1_REG_9__SCAN_IN), .ZN(n15034) );
  NAND2_X1 U10617 ( .A1(P3_REG1_REG_10__SCAN_IN), .A2(n14866), .ZN(n8302) );
  OAI21_X1 U10618 ( .B1(P3_REG1_REG_10__SCAN_IN), .B2(n14866), .A(n8302), .ZN(
        n14858) );
  INV_X1 U10619 ( .A(n8302), .ZN(n8303) );
  INV_X1 U10620 ( .A(P3_REG1_REG_11__SCAN_IN), .ZN(n14881) );
  NOR2_X1 U10621 ( .A1(n8346), .A2(n8304), .ZN(n8305) );
  INV_X1 U10622 ( .A(P3_REG1_REG_12__SCAN_IN), .ZN(n14307) );
  AOI22_X1 U10623 ( .A1(P3_REG1_REG_12__SCAN_IN), .A2(n8350), .B1(n12158), 
        .B2(n14307), .ZN(n12150) );
  AOI21_X2 U10624 ( .B1(P3_REG1_REG_12__SCAN_IN), .B2(n12158), .A(n12149), 
        .ZN(n8306) );
  INV_X1 U10625 ( .A(P3_REG1_REG_13__SCAN_IN), .ZN(n14303) );
  NAND2_X1 U10626 ( .A1(n8692), .A2(P3_REG1_REG_14__SCAN_IN), .ZN(n8355) );
  OAI21_X1 U10627 ( .B1(n8692), .B2(P3_REG1_REG_14__SCAN_IN), .A(n8355), .ZN(
        n12179) );
  INV_X1 U10628 ( .A(n8355), .ZN(n8308) );
  NOR2_X1 U10629 ( .A1(n8310), .A2(n8309), .ZN(n8311) );
  INV_X1 U10630 ( .A(P3_REG1_REG_15__SCAN_IN), .ZN(n12535) );
  INV_X1 U10631 ( .A(P3_REG1_REG_16__SCAN_IN), .ZN(n12531) );
  AOI22_X1 U10632 ( .A1(P3_REG1_REG_16__SCAN_IN), .A2(n8312), .B1(n12222), 
        .B2(n12531), .ZN(n12224) );
  INV_X1 U10633 ( .A(P3_REG1_REG_17__SCAN_IN), .ZN(n12527) );
  NOR2_X1 U10634 ( .A1(n12243), .A2(n12527), .ZN(n12242) );
  NOR2_X1 U10635 ( .A1(n12247), .A2(n8313), .ZN(n8314) );
  INV_X1 U10636 ( .A(P3_REG1_REG_18__SCAN_IN), .ZN(n12523) );
  AOI22_X1 U10637 ( .A1(P3_REG1_REG_18__SCAN_IN), .A2(n12263), .B1(n9134), 
        .B2(n12523), .ZN(n12261) );
  XNOR2_X1 U10638 ( .A(n8375), .B(P3_REG1_REG_19__SCAN_IN), .ZN(n8366) );
  INV_X1 U10639 ( .A(P3_REG2_REG_18__SCAN_IN), .ZN(n8317) );
  MUX2_X1 U10640 ( .A(n8317), .B(n12523), .S(n12602), .Z(n12254) );
  MUX2_X1 U10641 ( .A(P3_REG2_REG_17__SCAN_IN), .B(P3_REG1_REG_17__SCAN_IN), 
        .S(n12602), .Z(n8361) );
  AND2_X1 U10642 ( .A1(n8361), .A2(n9060), .ZN(n8363) );
  AND2_X1 U10643 ( .A1(n8360), .A2(n12222), .ZN(n12216) );
  MUX2_X1 U10644 ( .A(P3_REG2_REG_13__SCAN_IN), .B(P3_REG1_REG_13__SCAN_IN), 
        .S(n12602), .Z(n8318) );
  NOR2_X1 U10645 ( .A1(n8318), .A2(n8655), .ZN(n12186) );
  MUX2_X1 U10646 ( .A(n12181), .B(n12179), .S(n12602), .Z(n12184) );
  XNOR2_X1 U10647 ( .A(n8318), .B(n8655), .ZN(n12169) );
  NAND2_X1 U10648 ( .A1(n8351), .A2(n12158), .ZN(n8354) );
  MUX2_X1 U10649 ( .A(n14874), .B(n14881), .S(n12602), .Z(n8347) );
  NAND2_X1 U10650 ( .A1(n8347), .A2(n8346), .ZN(n8349) );
  INV_X1 U10651 ( .A(P3_REG2_REG_10__SCAN_IN), .ZN(n14904) );
  INV_X1 U10652 ( .A(P3_REG1_REG_10__SCAN_IN), .ZN(n8319) );
  MUX2_X1 U10653 ( .A(n14904), .B(n8319), .S(n12602), .Z(n8343) );
  INV_X1 U10654 ( .A(n14866), .ZN(n8344) );
  AND2_X1 U10655 ( .A1(n8343), .A2(n8344), .ZN(n8345) );
  MUX2_X1 U10656 ( .A(n10333), .B(n15034), .S(n12602), .Z(n8341) );
  INV_X1 U10657 ( .A(n8341), .ZN(n8320) );
  NAND2_X1 U10658 ( .A1(n8320), .A2(n10341), .ZN(n10335) );
  MUX2_X1 U10659 ( .A(P3_REG2_REG_8__SCAN_IN), .B(P3_REG1_REG_8__SCAN_IN), .S(
        n12602), .Z(n8337) );
  XNOR2_X1 U10660 ( .A(n8337), .B(n14845), .ZN(n14842) );
  MUX2_X1 U10661 ( .A(n9896), .B(n15030), .S(n12602), .Z(n8322) );
  NAND2_X1 U10662 ( .A1(n8322), .A2(n8321), .ZN(n8336) );
  XNOR2_X1 U10663 ( .A(n8322), .B(n9901), .ZN(n9899) );
  MUX2_X1 U10664 ( .A(P3_REG2_REG_6__SCAN_IN), .B(P3_REG1_REG_6__SCAN_IN), .S(
        n12602), .Z(n8323) );
  OR2_X1 U10665 ( .A1(n8323), .A2(n8620), .ZN(n8335) );
  XNOR2_X1 U10666 ( .A(n8323), .B(n14826), .ZN(n14823) );
  MUX2_X1 U10667 ( .A(n9393), .B(n9387), .S(n12602), .Z(n8324) );
  NAND2_X1 U10668 ( .A1(n8324), .A2(n9398), .ZN(n8334) );
  XNOR2_X1 U10669 ( .A(n8324), .B(n8626), .ZN(n9390) );
  MUX2_X1 U10670 ( .A(P3_REG2_REG_4__SCAN_IN), .B(P3_REG1_REG_4__SCAN_IN), .S(
        n12602), .Z(n8325) );
  OR2_X1 U10671 ( .A1(n8325), .A2(n9185), .ZN(n8333) );
  XOR2_X1 U10672 ( .A(n9185), .B(n8325), .Z(n9172) );
  OR2_X1 U10673 ( .A1(n8326), .A2(n8632), .ZN(n8332) );
  XNOR2_X1 U10674 ( .A(n8326), .B(n9072), .ZN(n9075) );
  OR2_X1 U10675 ( .A1(n8327), .A2(n9058), .ZN(n8331) );
  XOR2_X1 U10676 ( .A(n9058), .B(n8327), .Z(n9041) );
  INV_X1 U10677 ( .A(P3_REG2_REG_0__SCAN_IN), .ZN(n9891) );
  INV_X1 U10678 ( .A(P3_REG1_REG_0__SCAN_IN), .ZN(n8329) );
  AND2_X1 U10679 ( .A1(n14810), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n14813) );
  NAND2_X1 U10680 ( .A1(n9217), .A2(n14813), .ZN(n9216) );
  OAI21_X1 U10681 ( .B1(n8330), .B2(n9226), .A(n9216), .ZN(n9042) );
  NAND2_X1 U10682 ( .A1(n9041), .A2(n9042), .ZN(n9040) );
  NAND2_X1 U10683 ( .A1(n8331), .A2(n9040), .ZN(n9074) );
  NAND2_X1 U10684 ( .A1(n9075), .A2(n9074), .ZN(n9073) );
  NAND2_X1 U10685 ( .A1(n8332), .A2(n9073), .ZN(n9171) );
  NAND2_X1 U10686 ( .A1(n9172), .A2(n9171), .ZN(n9170) );
  NAND2_X1 U10687 ( .A1(n8333), .A2(n9170), .ZN(n9389) );
  NAND2_X1 U10688 ( .A1(n9390), .A2(n9389), .ZN(n9388) );
  NAND2_X1 U10689 ( .A1(n8334), .A2(n9388), .ZN(n14824) );
  NAND2_X1 U10690 ( .A1(n14823), .A2(n14824), .ZN(n14822) );
  NAND2_X1 U10691 ( .A1(n8335), .A2(n14822), .ZN(n9898) );
  NAND2_X1 U10692 ( .A1(n9899), .A2(n9898), .ZN(n9897) );
  INV_X1 U10693 ( .A(n8337), .ZN(n8338) );
  NAND2_X1 U10694 ( .A1(n8338), .A2(n14845), .ZN(n8339) );
  NAND2_X1 U10695 ( .A1(n8340), .A2(n8339), .ZN(n10338) );
  AND2_X1 U10696 ( .A1(n8341), .A2(n6680), .ZN(n10334) );
  INV_X1 U10697 ( .A(n8345), .ZN(n8342) );
  OAI21_X1 U10698 ( .B1(n8344), .B2(n8343), .A(n8342), .ZN(n14864) );
  NOR2_X1 U10699 ( .A1(n14863), .A2(n14864), .ZN(n14862) );
  NOR2_X1 U10700 ( .A1(n8345), .A2(n14862), .ZN(n14883) );
  OAI21_X1 U10701 ( .B1(n8347), .B2(n8346), .A(n8349), .ZN(n14884) );
  INV_X1 U10702 ( .A(n14882), .ZN(n8348) );
  INV_X1 U10703 ( .A(n12153), .ZN(n8352) );
  XNOR2_X1 U10704 ( .A(n8351), .B(n8350), .ZN(n12154) );
  NAND2_X1 U10705 ( .A1(n8352), .A2(n12154), .ZN(n8353) );
  NAND2_X1 U10706 ( .A1(n12187), .A2(n8357), .ZN(n8358) );
  MUX2_X1 U10707 ( .A(P3_REG2_REG_15__SCAN_IN), .B(P3_REG1_REG_15__SCAN_IN), 
        .S(n12602), .Z(n12202) );
  NOR2_X1 U10708 ( .A1(n8359), .A2(n12200), .ZN(n12218) );
  NOR2_X1 U10709 ( .A1(n8360), .A2(n12222), .ZN(n12217) );
  NOR2_X1 U10710 ( .A1(n8361), .A2(n9060), .ZN(n8362) );
  OR2_X1 U10711 ( .A1(n8363), .A2(n8362), .ZN(n12235) );
  XNOR2_X1 U10712 ( .A(n9134), .B(n8364), .ZN(n12255) );
  NAND2_X1 U10713 ( .A1(n12254), .A2(n12255), .ZN(n12253) );
  NAND2_X1 U10714 ( .A1(n12263), .A2(n8364), .ZN(n8365) );
  NAND2_X1 U10715 ( .A1(n12253), .A2(n8365), .ZN(n8369) );
  XNOR2_X1 U10716 ( .A(n8369), .B(n8368), .ZN(n8380) );
  NOR2_X2 U10717 ( .A1(n12143), .A2(n8373), .ZN(n14843) );
  INV_X1 U10718 ( .A(n8370), .ZN(n8372) );
  INV_X1 U10719 ( .A(n14869), .ZN(n14875) );
  MUX2_X1 U10720 ( .A(n8374), .B(P3_U3897), .S(n8373), .Z(n14846) );
  NAND2_X1 U10721 ( .A1(n14846), .A2(n8375), .ZN(n8377) );
  NAND2_X1 U10722 ( .A1(P3_REG3_REG_19__SCAN_IN), .A2(P3_U3151), .ZN(n8376) );
  OAI211_X1 U10723 ( .C1(n8378), .C2(n14875), .A(n8377), .B(n8376), .ZN(n8379)
         );
  OR2_X1 U10724 ( .A1(n12022), .A2(n7281), .ZN(n8384) );
  AND2_X1 U10725 ( .A1(n8384), .A2(n8383), .ZN(n8387) );
  NAND2_X1 U10726 ( .A1(n8390), .A2(n8387), .ZN(n8385) );
  NAND2_X1 U10727 ( .A1(n8385), .A2(n11974), .ZN(n8386) );
  NAND2_X1 U10728 ( .A1(n8386), .A2(n14961), .ZN(n8391) );
  INV_X1 U10729 ( .A(n11974), .ZN(n8388) );
  NOR2_X1 U10730 ( .A1(n8391), .A2(n8402), .ZN(n8395) );
  OR2_X1 U10731 ( .A1(n9376), .A2(n12100), .ZN(n8393) );
  NAND2_X1 U10732 ( .A1(n7281), .A2(n12440), .ZN(n8392) );
  AND2_X1 U10733 ( .A1(n8393), .A2(n8392), .ZN(n11977) );
  NAND2_X1 U10734 ( .A1(n8397), .A2(n8396), .ZN(n8398) );
  XNOR2_X1 U10735 ( .A(n8398), .B(n11974), .ZN(n12283) );
  MUX2_X1 U10736 ( .A(P3_REG1_REG_28__SCAN_IN), .B(n11163), .S(n15038), .Z(
        n8400) );
  INV_X1 U10737 ( .A(n12537), .ZN(n10361) );
  OR2_X1 U10738 ( .A1(n8400), .A2(n8399), .ZN(P3_U3487) );
  NOR2_X1 U10739 ( .A1(n8402), .A2(n8401), .ZN(n8403) );
  INV_X1 U10740 ( .A(P3_B_REG_SCAN_IN), .ZN(n8404) );
  NOR2_X1 U10741 ( .A1(n7945), .A2(n8404), .ZN(n8405) );
  OR2_X1 U10742 ( .A1(n12100), .A2(n8405), .ZN(n12265) );
  OAI22_X1 U10743 ( .A1(n8407), .A2(n12103), .B1(n12265), .B2(n8406), .ZN(
        n8408) );
  INV_X1 U10744 ( .A(n8408), .ZN(n8409) );
  XOR2_X1 U10745 ( .A(n8411), .B(n8207), .Z(n12277) );
  INV_X1 U10746 ( .A(n8412), .ZN(n8414) );
  INV_X1 U10747 ( .A(n8417), .ZN(n8413) );
  NAND2_X1 U10748 ( .A1(n8414), .A2(n8413), .ZN(n9517) );
  NAND2_X1 U10749 ( .A1(n8415), .A2(n9547), .ZN(n9502) );
  OR2_X1 U10750 ( .A1(n8416), .A2(n9546), .ZN(n9515) );
  AND2_X1 U10751 ( .A1(n9502), .A2(n9515), .ZN(n8420) );
  INV_X1 U10752 ( .A(n9513), .ZN(n8419) );
  OAI22_X1 U10753 ( .A1(n9517), .A2(n8420), .B1(n8419), .B2(n9514), .ZN(n8421)
         );
  INV_X1 U10754 ( .A(n8423), .ZN(n12275) );
  INV_X1 U10755 ( .A(P3_REG0_REG_29__SCAN_IN), .ZN(n8424) );
  INV_X1 U10756 ( .A(n8426), .ZN(n8427) );
  INV_X1 U10757 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n8428) );
  NAND2_X1 U10758 ( .A1(n8973), .A2(n8428), .ZN(n8905) );
  INV_X1 U10759 ( .A(n8905), .ZN(n8432) );
  NOR2_X1 U10760 ( .A1(P2_IR_REG_14__SCAN_IN), .A2(P2_IR_REG_18__SCAN_IN), 
        .ZN(n8431) );
  NOR2_X1 U10761 ( .A1(P2_IR_REG_17__SCAN_IN), .A2(P2_IR_REG_19__SCAN_IN), 
        .ZN(n8430) );
  AND4_X2 U10762 ( .A1(n8432), .A2(n8431), .A3(n8430), .A4(n8429), .ZN(n8436)
         );
  NOR2_X1 U10763 ( .A1(P2_IR_REG_6__SCAN_IN), .A2(P2_IR_REG_10__SCAN_IN), .ZN(
        n8435) );
  NOR2_X1 U10764 ( .A1(P2_IR_REG_8__SCAN_IN), .A2(P2_IR_REG_7__SCAN_IN), .ZN(
        n8434) );
  NOR2_X1 U10765 ( .A1(P2_IR_REG_9__SCAN_IN), .A2(P2_IR_REG_11__SCAN_IN), .ZN(
        n8433) );
  NOR2_X1 U10766 ( .A1(P2_IR_REG_22__SCAN_IN), .A2(P2_IR_REG_23__SCAN_IN), 
        .ZN(n8440) );
  NOR2_X1 U10767 ( .A1(P2_IR_REG_21__SCAN_IN), .A2(P2_IR_REG_20__SCAN_IN), 
        .ZN(n8439) );
  NOR2_X1 U10768 ( .A1(P2_IR_REG_24__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), 
        .ZN(n8438) );
  NAND2_X1 U10769 ( .A1(n8664), .A2(n8665), .ZN(n8668) );
  NAND2_X1 U10770 ( .A1(n8447), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8444) );
  MUX2_X1 U10771 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8444), .S(
        P2_IR_REG_26__SCAN_IN), .Z(n8445) );
  INV_X1 U10772 ( .A(n13435), .ZN(n8455) );
  NAND2_X1 U10773 ( .A1(n8452), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8446) );
  MUX2_X1 U10774 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8446), .S(
        P2_IR_REG_25__SCAN_IN), .Z(n8448) );
  NAND2_X1 U10775 ( .A1(n8448), .A2(n8447), .ZN(n13437) );
  INV_X1 U10776 ( .A(n8449), .ZN(n8450) );
  NAND2_X1 U10777 ( .A1(n8450), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8451) );
  MUX2_X1 U10778 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8451), .S(
        P2_IR_REG_24__SCAN_IN), .Z(n8453) );
  NAND2_X1 U10779 ( .A1(n8453), .A2(n8452), .ZN(n11087) );
  NOR2_X1 U10780 ( .A1(n13437), .A2(n11087), .ZN(n8454) );
  NAND2_X1 U10781 ( .A1(n8455), .A2(n8454), .ZN(n9319) );
  NAND2_X1 U10782 ( .A1(n8668), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8457) );
  XNOR2_X1 U10783 ( .A(n8457), .B(n8456), .ZN(n9318) );
  INV_X1 U10784 ( .A(n8940), .ZN(n8458) );
  NOR2_X1 U10785 ( .A1(n9319), .A2(n8458), .ZN(P2_U3947) );
  NAND4_X1 U10786 ( .A1(n8781), .A2(n8460), .A3(n8582), .A4(n8459), .ZN(n8463)
         );
  NAND4_X1 U10787 ( .A1(n8967), .A2(n8784), .A3(n8970), .A4(n8461), .ZN(n8462)
         );
  INV_X1 U10788 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n8471) );
  NOR2_X1 U10789 ( .A1(P1_IR_REG_23__SCAN_IN), .A2(P1_IR_REG_25__SCAN_IN), 
        .ZN(n8473) );
  NAND2_X1 U10790 ( .A1(n11195), .A2(n8473), .ZN(n8475) );
  NAND3_X1 U10791 ( .A1(n9269), .A2(n9273), .A3(n7012), .ZN(n8474) );
  NAND2_X1 U10792 ( .A1(n8479), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8478) );
  MUX2_X1 U10793 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8478), .S(
        P1_IR_REG_26__SCAN_IN), .Z(n8480) );
  NAND2_X1 U10794 ( .A1(n8480), .A2(n8725), .ZN(n14127) );
  NAND2_X2 U10795 ( .A1(n8483), .A2(n9253), .ZN(n9284) );
  NAND2_X1 U10796 ( .A1(n8484), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8485) );
  INV_X1 U10797 ( .A(n8738), .ZN(n8486) );
  OR2_X2 U10798 ( .A1(n9284), .A2(n8486), .ZN(n13667) );
  NAND2_X1 U10799 ( .A1(n8495), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8487) );
  OAI21_X2 U10800 ( .B1(n8495), .B2(n8488), .A(n8487), .ZN(n8491) );
  INV_X1 U10801 ( .A(n8491), .ZN(n8489) );
  INV_X1 U10802 ( .A(SI_2_), .ZN(n8618) );
  NOR2_X1 U10803 ( .A1(n8532), .A2(n8618), .ZN(n8492) );
  NAND2_X1 U10804 ( .A1(n8496), .A2(n8492), .ZN(n8493) );
  MUX2_X1 U10805 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(P1_DATAO_REG_2__SCAN_IN), 
        .S(n8495), .Z(n8526) );
  INV_X1 U10806 ( .A(n8526), .ZN(n8500) );
  NAND2_X1 U10807 ( .A1(n8496), .A2(n8497), .ZN(n8533) );
  OAI21_X1 U10808 ( .B1(n8533), .B2(n8532), .A(n8497), .ZN(n8498) );
  NAND2_X1 U10809 ( .A1(n8498), .A2(SI_2_), .ZN(n8499) );
  NAND2_X1 U10810 ( .A1(n8503), .A2(SI_3_), .ZN(n8505) );
  OAI21_X1 U10811 ( .B1(SI_3_), .B2(n8503), .A(n8505), .ZN(n8539) );
  INV_X1 U10812 ( .A(n8539), .ZN(n8504) );
  NAND2_X1 U10813 ( .A1(n8538), .A2(n8504), .ZN(n8506) );
  MUX2_X1 U10814 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n8495), .Z(n8507) );
  NAND2_X1 U10815 ( .A1(n8507), .A2(SI_4_), .ZN(n8509) );
  OAI21_X1 U10816 ( .B1(SI_4_), .B2(n8507), .A(n8509), .ZN(n8508) );
  INV_X1 U10817 ( .A(n8508), .ZN(n8519) );
  MUX2_X1 U10818 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n8495), .Z(n8510) );
  NAND2_X1 U10819 ( .A1(n8510), .A2(SI_5_), .ZN(n8558) );
  OAI21_X1 U10820 ( .B1(SI_5_), .B2(n8510), .A(n8558), .ZN(n8555) );
  XNOR2_X1 U10821 ( .A(n8557), .B(n8555), .ZN(n9841) );
  INV_X1 U10822 ( .A(n9841), .ZN(n8616) );
  AND2_X1 U10823 ( .A1(n11543), .A2(P2_U3088), .ZN(n11064) );
  INV_X2 U10824 ( .A(n11064), .ZN(n13438) );
  AND2_X1 U10825 ( .A1(n8511), .A2(n8429), .ZN(n8512) );
  INV_X1 U10826 ( .A(n8516), .ZN(n8513) );
  NAND2_X1 U10827 ( .A1(n8513), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8514) );
  MUX2_X1 U10828 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8514), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n8517) );
  INV_X1 U10829 ( .A(n8886), .ZN(n8553) );
  NOR2_X1 U10830 ( .A1(n11543), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13428) );
  AOI22_X1 U10831 ( .A1(n14652), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_5__SCAN_IN), .B2(n13428), .ZN(n8518) );
  OAI21_X1 U10832 ( .B1(n8616), .B2(n13438), .A(n8518), .ZN(P2_U3322) );
  OR2_X1 U10833 ( .A1(n8520), .A2(n8519), .ZN(n8521) );
  AND2_X1 U10834 ( .A1(n8522), .A2(n8521), .ZN(n9621) );
  INV_X1 U10835 ( .A(n9621), .ZN(n8589) );
  NAND2_X1 U10836 ( .A1(n8523), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8524) );
  XNOR2_X1 U10837 ( .A(n8524), .B(P2_IR_REG_4__SCAN_IN), .ZN(n14638) );
  AOI22_X1 U10838 ( .A1(n14638), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_4__SCAN_IN), .B2(n13428), .ZN(n8525) );
  OAI21_X1 U10839 ( .B1(n8589), .B2(n13438), .A(n8525), .ZN(P2_U3323) );
  INV_X2 U10840 ( .A(n13428), .ZN(n13440) );
  XNOR2_X1 U10841 ( .A(n8527), .B(n8526), .ZN(n9017) );
  INV_X1 U10842 ( .A(n9017), .ZN(n9570) );
  NAND2_X1 U10843 ( .A1(n8535), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8528) );
  MUX2_X1 U10844 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8528), .S(
        P2_IR_REG_2__SCAN_IN), .Z(n8530) );
  NAND2_X1 U10845 ( .A1(n8530), .A2(n8529), .ZN(n9019) );
  OAI222_X1 U10846 ( .A1(n13440), .A2(n8531), .B1(n13438), .B2(n9570), .C1(
        n9019), .C2(P2_U3088), .ZN(P2_U3325) );
  XNOR2_X1 U10847 ( .A(n8533), .B(n8532), .ZN(n9576) );
  NAND2_X1 U10848 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), 
        .ZN(n8534) );
  MUX2_X1 U10849 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8534), .S(
        P2_IR_REG_1__SCAN_IN), .Z(n8536) );
  OAI222_X1 U10850 ( .A1(n13440), .A2(n8537), .B1(n13438), .B2(n9576), .C1(
        n13069), .C2(P2_U3088), .ZN(P2_U3326) );
  XNOR2_X1 U10851 ( .A(n8538), .B(n8539), .ZN(n9600) );
  INV_X1 U10852 ( .A(n9600), .ZN(n8609) );
  NAND2_X1 U10853 ( .A1(n8529), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8540) );
  MUX2_X1 U10854 ( .A(P2_IR_REG_31__SCAN_IN), .B(n8540), .S(
        P2_IR_REG_3__SCAN_IN), .Z(n8541) );
  AND2_X1 U10855 ( .A1(n8541), .A2(n8523), .ZN(n9098) );
  INV_X1 U10856 ( .A(n9098), .ZN(n8749) );
  OAI222_X1 U10857 ( .A1(n13440), .A2(n8542), .B1(n13438), .B2(n8609), .C1(
        P2_U3088), .C2(n8749), .ZN(P2_U3324) );
  OR2_X1 U10858 ( .A1(n8543), .A2(n14111), .ZN(n8544) );
  XNOR2_X1 U10859 ( .A(n8544), .B(P1_IR_REG_2__SCAN_IN), .ZN(n13689) );
  INV_X1 U10860 ( .A(n13689), .ZN(n8546) );
  INV_X1 U10861 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n8545) );
  NAND2_X1 U10862 ( .A1(n11361), .A2(P1_U3086), .ZN(n14130) );
  OAI222_X1 U10863 ( .A1(P1_U3086), .A2(n8546), .B1(n14124), .B2(n8545), .C1(
        n14130), .C2(n9570), .ZN(P1_U3353) );
  INV_X1 U10864 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n13671) );
  NAND2_X1 U10865 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), 
        .ZN(n8547) );
  MUX2_X1 U10866 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8547), .S(
        P1_IR_REG_1__SCAN_IN), .Z(n8549) );
  INV_X1 U10867 ( .A(n8543), .ZN(n8548) );
  NAND2_X1 U10868 ( .A1(n8549), .A2(n8548), .ZN(n13669) );
  OAI222_X1 U10869 ( .A1(P1_U3086), .A2(n13669), .B1(n14124), .B2(n8488), .C1(
        n14130), .C2(n9576), .ZN(P1_U3354) );
  NAND2_X1 U10870 ( .A1(n11543), .A2(P3_U3151), .ZN(n12608) );
  NOR2_X1 U10871 ( .A1(n11543), .A2(P3_STATE_REG_SCAN_IN), .ZN(n12596) );
  INV_X1 U10872 ( .A(n12596), .ZN(n12607) );
  INV_X1 U10873 ( .A(n8550), .ZN(n8552) );
  OAI222_X1 U10874 ( .A1(n12608), .A2(n9280), .B1(n12607), .B2(n8552), .C1(
        P3_U3151), .C2(n8551), .ZN(P3_U3295) );
  NAND2_X1 U10875 ( .A1(n8553), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8554) );
  XNOR2_X1 U10876 ( .A(n8554), .B(P2_IR_REG_6__SCAN_IN), .ZN(n9191) );
  INV_X1 U10877 ( .A(n9191), .ZN(n13087) );
  INV_X1 U10878 ( .A(n8555), .ZN(n8556) );
  MUX2_X1 U10879 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n11543), .Z(n8559) );
  NAND2_X1 U10880 ( .A1(n8559), .A2(SI_6_), .ZN(n8573) );
  OAI21_X1 U10881 ( .B1(SI_6_), .B2(n8559), .A(n8573), .ZN(n8560) );
  INV_X1 U10882 ( .A(n8560), .ZN(n8561) );
  OR2_X1 U10883 ( .A1(n8562), .A2(n8561), .ZN(n8563) );
  NAND2_X1 U10884 ( .A1(n8563), .A2(n8574), .ZN(n9845) );
  OAI222_X1 U10885 ( .A1(P2_U3088), .A2(n13087), .B1(n13440), .B2(n8564), .C1(
        n13438), .C2(n9845), .ZN(P2_U3321) );
  INV_X1 U10886 ( .A(SI_10_), .ZN(n8565) );
  OAI222_X1 U10887 ( .A1(n12607), .A2(n8566), .B1(n14866), .B2(P3_U3151), .C1(
        n8565), .C2(n12608), .ZN(P3_U3285) );
  INV_X1 U10888 ( .A(SI_9_), .ZN(n8567) );
  OAI222_X1 U10889 ( .A1(n12607), .A2(n8568), .B1(n10341), .B2(P3_U3151), .C1(
        n8567), .C2(n12608), .ZN(P3_U3286) );
  INV_X1 U10890 ( .A(SI_7_), .ZN(n8569) );
  OAI222_X1 U10891 ( .A1(n12607), .A2(n8570), .B1(n9901), .B2(P3_U3151), .C1(
        n8569), .C2(n12608), .ZN(P3_U3288) );
  INV_X1 U10892 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n8571) );
  NAND2_X1 U10893 ( .A1(n8886), .A2(n8571), .ZN(n8637) );
  NAND2_X1 U10894 ( .A1(n8637), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8572) );
  XNOR2_X1 U10895 ( .A(n8572), .B(P2_IR_REG_7__SCAN_IN), .ZN(n13105) );
  INV_X1 U10896 ( .A(n13105), .ZN(n13103) );
  INV_X1 U10897 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n8580) );
  MUX2_X1 U10898 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(P1_DATAO_REG_7__SCAN_IN), 
        .S(n11543), .Z(n8575) );
  NAND2_X1 U10899 ( .A1(n8575), .A2(SI_7_), .ZN(n8593) );
  OAI21_X1 U10900 ( .B1(SI_7_), .B2(n8575), .A(n8593), .ZN(n8576) );
  INV_X1 U10901 ( .A(n8576), .ZN(n8577) );
  NAND2_X1 U10902 ( .A1(n8578), .A2(n8577), .ZN(n8594) );
  OR2_X1 U10903 ( .A1(n8578), .A2(n8577), .ZN(n8579) );
  NAND2_X1 U10904 ( .A1(n8594), .A2(n8579), .ZN(n10172) );
  OAI222_X1 U10905 ( .A1(P2_U3088), .A2(n13103), .B1(n13440), .B2(n8580), .C1(
        n13438), .C2(n10172), .ZN(P2_U3320) );
  NAND2_X1 U10906 ( .A1(n8581), .A2(n8582), .ZN(n8612) );
  NAND2_X1 U10907 ( .A1(n8600), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8583) );
  XNOR2_X1 U10908 ( .A(n8583), .B(P1_IR_REG_7__SCAN_IN), .ZN(n13747) );
  INV_X1 U10909 ( .A(n13747), .ZN(n8836) );
  OAI222_X1 U10910 ( .A1(n14124), .A2(n8584), .B1(n14130), .B2(n10172), .C1(
        n8836), .C2(P1_U3086), .ZN(P1_U3348) );
  INV_X1 U10911 ( .A(n8585), .ZN(n8586) );
  OAI222_X1 U10912 ( .A1(n12607), .A2(n8586), .B1(n12158), .B2(P3_U3151), .C1(
        n15174), .C2(n12608), .ZN(P3_U3283) );
  OR2_X1 U10913 ( .A1(n8587), .A2(P1_IR_REG_3__SCAN_IN), .ZN(n8607) );
  NAND2_X1 U10914 ( .A1(n8607), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8588) );
  XNOR2_X1 U10915 ( .A(n8588), .B(P1_IR_REG_4__SCAN_IN), .ZN(n13721) );
  INV_X1 U10916 ( .A(n13721), .ZN(n8590) );
  INV_X1 U10917 ( .A(P2_DATAO_REG_4__SCAN_IN), .ZN(n9624) );
  OAI222_X1 U10918 ( .A1(P1_U3086), .A2(n8590), .B1(n14124), .B2(n9624), .C1(
        n14130), .C2(n8589), .ZN(P1_U3351) );
  NAND2_X1 U10919 ( .A1(n8612), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8591) );
  XNOR2_X1 U10920 ( .A(n8591), .B(P1_IR_REG_6__SCAN_IN), .ZN(n9847) );
  INV_X1 U10921 ( .A(n9847), .ZN(n8985) );
  OAI222_X1 U10922 ( .A1(P1_U3086), .A2(n8985), .B1(n14124), .B2(n8592), .C1(
        n14130), .C2(n9845), .ZN(P1_U3349) );
  INV_X1 U10923 ( .A(n14130), .ZN(n11068) );
  INV_X1 U10924 ( .A(n11068), .ZN(n14119) );
  NAND2_X1 U10925 ( .A1(n8594), .A2(n8593), .ZN(n8598) );
  MUX2_X1 U10926 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n11543), .Z(n8595) );
  NAND2_X1 U10927 ( .A1(n8595), .A2(SI_8_), .ZN(n8640) );
  OAI21_X1 U10928 ( .B1(SI_8_), .B2(n8595), .A(n8640), .ZN(n8596) );
  INV_X1 U10929 ( .A(n8596), .ZN(n8597) );
  NAND2_X1 U10930 ( .A1(n8598), .A2(n8597), .ZN(n8641) );
  OR2_X1 U10931 ( .A1(n8598), .A2(n8597), .ZN(n8599) );
  NAND2_X1 U10932 ( .A1(n8641), .A2(n8599), .ZN(n10199) );
  OR2_X1 U10933 ( .A1(n8603), .A2(n14111), .ZN(n8601) );
  MUX2_X1 U10934 ( .A(n8601), .B(P1_IR_REG_31__SCAN_IN), .S(n8602), .Z(n8604)
         );
  NAND2_X1 U10935 ( .A1(n8603), .A2(n8602), .ZN(n8647) );
  NAND2_X1 U10936 ( .A1(n8604), .A2(n8647), .ZN(n8858) );
  OAI222_X1 U10937 ( .A1(n14124), .A2(n8605), .B1(n14119), .B2(n10199), .C1(
        n8858), .C2(P1_U3086), .ZN(P1_U3347) );
  NAND2_X1 U10938 ( .A1(n8587), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8606) );
  MUX2_X1 U10939 ( .A(P1_IR_REG_31__SCAN_IN), .B(n8606), .S(
        P1_IR_REG_3__SCAN_IN), .Z(n8608) );
  AND2_X1 U10940 ( .A1(n8608), .A2(n8607), .ZN(n13703) );
  INV_X1 U10941 ( .A(n13703), .ZN(n8610) );
  OAI222_X1 U10942 ( .A1(n8610), .A2(P1_U3086), .B1(n14119), .B2(n8609), .C1(
        n8502), .C2(n14124), .ZN(P1_U3352) );
  NOR2_X1 U10943 ( .A1(n8581), .A2(n14111), .ZN(n8611) );
  MUX2_X1 U10944 ( .A(n14111), .B(n8611), .S(P1_IR_REG_5__SCAN_IN), .Z(n8614)
         );
  INV_X1 U10945 ( .A(n8612), .ZN(n8613) );
  OR2_X1 U10946 ( .A1(n8614), .A2(n8613), .ZN(n13736) );
  INV_X1 U10947 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n8615) );
  OAI222_X1 U10948 ( .A1(n13736), .A2(P1_U3086), .B1(n14119), .B2(n8616), .C1(
        n8615), .C2(n14124), .ZN(P1_U3350) );
  INV_X1 U10949 ( .A(n12608), .ZN(n12594) );
  INV_X1 U10950 ( .A(n12594), .ZN(n12589) );
  OAI222_X1 U10951 ( .A1(n12589), .A2(n8618), .B1(n12607), .B2(n8617), .C1(
        P3_U3151), .C2(n9058), .ZN(P3_U3293) );
  INV_X1 U10952 ( .A(n8619), .ZN(n8621) );
  OAI222_X1 U10953 ( .A1(n12589), .A2(n15225), .B1(n12607), .B2(n8621), .C1(
        P3_U3151), .C2(n8620), .ZN(P3_U3289) );
  INV_X1 U10954 ( .A(n8622), .ZN(n8623) );
  OAI222_X1 U10955 ( .A1(n12589), .A2(n8625), .B1(n8624), .B2(P3_U3151), .C1(
        n12607), .C2(n8623), .ZN(P3_U3287) );
  INV_X1 U10956 ( .A(SI_5_), .ZN(n8628) );
  OAI222_X1 U10957 ( .A1(n12589), .A2(n8628), .B1(n12607), .B2(n8627), .C1(
        P3_U3151), .C2(n8626), .ZN(P3_U3290) );
  INV_X1 U10958 ( .A(n8629), .ZN(n8630) );
  OAI222_X1 U10959 ( .A1(n12589), .A2(n8631), .B1(n9226), .B2(P3_U3151), .C1(
        n12607), .C2(n8630), .ZN(P3_U3294) );
  INV_X1 U10960 ( .A(SI_3_), .ZN(n8634) );
  OAI222_X1 U10961 ( .A1(n12589), .A2(n8634), .B1(n12607), .B2(n8633), .C1(
        P3_U3151), .C2(n8632), .ZN(P3_U3292) );
  INV_X1 U10962 ( .A(SI_4_), .ZN(n8636) );
  OAI222_X1 U10963 ( .A1(n12589), .A2(n8636), .B1(n12607), .B2(n8635), .C1(
        P3_U3151), .C2(n9185), .ZN(P3_U3291) );
  NAND2_X1 U10964 ( .A1(n8652), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8638) );
  XNOR2_X1 U10965 ( .A(n8638), .B(P2_IR_REG_8__SCAN_IN), .ZN(n9731) );
  INV_X1 U10966 ( .A(n9731), .ZN(n8871) );
  INV_X1 U10967 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n8639) );
  OAI222_X1 U10968 ( .A1(P2_U3088), .A2(n8871), .B1(n13440), .B2(n8639), .C1(
        n13438), .C2(n10199), .ZN(P2_U3319) );
  MUX2_X1 U10969 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n11543), .Z(n8642) );
  NAND2_X1 U10970 ( .A1(n8642), .A2(SI_9_), .ZN(n8657) );
  OAI21_X1 U10971 ( .B1(SI_9_), .B2(n8642), .A(n8657), .ZN(n8643) );
  INV_X1 U10972 ( .A(n8643), .ZN(n8644) );
  OR2_X1 U10973 ( .A1(n8645), .A2(n8644), .ZN(n8646) );
  NAND2_X1 U10974 ( .A1(n8658), .A2(n8646), .ZN(n10205) );
  NAND2_X1 U10975 ( .A1(n8647), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8783) );
  INV_X1 U10976 ( .A(P1_IR_REG_9__SCAN_IN), .ZN(n8648) );
  NAND2_X1 U10977 ( .A1(n8783), .A2(n8648), .ZN(n8660) );
  OR2_X1 U10978 ( .A1(n8783), .A2(n8648), .ZN(n8649) );
  INV_X1 U10979 ( .A(n14124), .ZN(n14114) );
  AOI22_X1 U10980 ( .A1(n13769), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n14114), .ZN(n8650) );
  OAI21_X1 U10981 ( .B1(n10205), .B2(n14119), .A(n8650), .ZN(P1_U3346) );
  OAI222_X1 U10982 ( .A1(n12607), .A2(n8651), .B1(n14877), .B2(P3_U3151), .C1(
        n12589), .C2(n15209), .ZN(P3_U3284) );
  NAND2_X1 U10983 ( .A1(n8694), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8653) );
  XNOR2_X1 U10984 ( .A(n8653), .B(P2_IR_REG_9__SCAN_IN), .ZN(n9786) );
  INV_X1 U10985 ( .A(n9786), .ZN(n9080) );
  INV_X1 U10986 ( .A(P1_DATAO_REG_9__SCAN_IN), .ZN(n8654) );
  OAI222_X1 U10987 ( .A1(P2_U3088), .A2(n9080), .B1(n13440), .B2(n8654), .C1(
        n13438), .C2(n10205), .ZN(P2_U3318) );
  INV_X1 U10988 ( .A(SI_13_), .ZN(n15203) );
  OAI222_X1 U10989 ( .A1(n12608), .A2(n15203), .B1(n12607), .B2(n8656), .C1(
        P3_U3151), .C2(n8655), .ZN(P3_U3282) );
  MUX2_X1 U10990 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n11543), .Z(n8659) );
  NAND2_X1 U10991 ( .A1(n8659), .A2(SI_10_), .ZN(n8768) );
  OAI21_X1 U10992 ( .B1(SI_10_), .B2(n8659), .A(n8768), .ZN(n8765) );
  XNOR2_X1 U10993 ( .A(n8767), .B(n7416), .ZN(n10456) );
  INV_X1 U10994 ( .A(n10456), .ZN(n8699) );
  NAND2_X1 U10995 ( .A1(n8660), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8661) );
  XNOR2_X1 U10996 ( .A(n8661), .B(P1_IR_REG_10__SCAN_IN), .ZN(n10457) );
  AOI22_X1 U10997 ( .A1(n10457), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n14114), .ZN(n8662) );
  OAI21_X1 U10998 ( .B1(n8699), .B2(n14119), .A(n8662), .ZN(P1_U3345) );
  INV_X1 U10999 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n8663) );
  XNOR2_X1 U11000 ( .A(n13069), .B(P2_REG1_REG_1__SCAN_IN), .ZN(n13078) );
  NAND3_X1 U11001 ( .A1(n13078), .A2(P2_IR_REG_0__SCAN_IN), .A3(
        P2_REG1_REG_0__SCAN_IN), .ZN(n13076) );
  OAI21_X1 U11002 ( .B1(n13069), .B2(n8663), .A(n13076), .ZN(n8751) );
  XNOR2_X1 U11003 ( .A(n9019), .B(P2_REG1_REG_2__SCAN_IN), .ZN(n8750) );
  XNOR2_X1 U11004 ( .A(n8751), .B(n8750), .ZN(n8691) );
  INV_X1 U11005 ( .A(n9318), .ZN(n11065) );
  INV_X1 U11006 ( .A(n8931), .ZN(n14742) );
  NOR2_X1 U11007 ( .A1(n12720), .A2(n14742), .ZN(n9324) );
  NAND2_X1 U11008 ( .A1(n9324), .A2(n9318), .ZN(n8675) );
  INV_X1 U11009 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n8671) );
  NAND2_X1 U11010 ( .A1(n8675), .A2(n8899), .ZN(n8676) );
  OAI21_X1 U11011 ( .B1(n9319), .B2(n11065), .A(n8676), .ZN(n8679) );
  NOR2_X1 U11012 ( .A1(n8677), .A2(P2_U3088), .ZN(n13427) );
  NAND2_X1 U11013 ( .A1(n8679), .A2(n13427), .ZN(n8683) );
  INV_X1 U11014 ( .A(n13432), .ZN(n11867) );
  OR2_X1 U11015 ( .A1(n8679), .A2(P2_U3088), .ZN(n14671) );
  INV_X1 U11016 ( .A(n14671), .ZN(n14685) );
  AND2_X1 U11017 ( .A1(n8677), .A2(P2_STATE_REG_SCAN_IN), .ZN(n8678) );
  NAND2_X1 U11018 ( .A1(n8679), .A2(n8678), .ZN(n14667) );
  INV_X1 U11019 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n8680) );
  OAI22_X1 U11020 ( .A1(n14667), .A2(n9019), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8680), .ZN(n8681) );
  AOI21_X1 U11021 ( .B1(n14685), .B2(P2_ADDR_REG_2__SCAN_IN), .A(n8681), .ZN(
        n8690) );
  INV_X1 U11022 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n8682) );
  MUX2_X1 U11023 ( .A(n8682), .B(P2_REG2_REG_2__SCAN_IN), .S(n9019), .Z(n8688)
         );
  INV_X1 U11024 ( .A(n13069), .ZN(n8890) );
  INV_X1 U11025 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n9378) );
  MUX2_X1 U11026 ( .A(P2_REG2_REG_1__SCAN_IN), .B(n9378), .S(n13069), .Z(
        n13072) );
  INV_X1 U11027 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n14631) );
  NOR3_X1 U11028 ( .A1(n13072), .A2(n14631), .A3(n13075), .ZN(n13071) );
  AOI21_X1 U11029 ( .B1(n8890), .B2(P2_REG2_REG_1__SCAN_IN), .A(n13071), .ZN(
        n8686) );
  INV_X1 U11030 ( .A(n8686), .ZN(n8687) );
  INV_X1 U11031 ( .A(n8683), .ZN(n8684) );
  MUX2_X1 U11032 ( .A(P2_REG2_REG_2__SCAN_IN), .B(n8682), .S(n9019), .Z(n8685)
         );
  OAI211_X1 U11033 ( .C1(n8688), .C2(n8687), .A(n14692), .B(n8758), .ZN(n8689)
         );
  OAI211_X1 U11034 ( .C1(n8691), .C2(n14639), .A(n8690), .B(n8689), .ZN(
        P2_U3216) );
  OAI222_X1 U11035 ( .A1(n12607), .A2(n8693), .B1(n8692), .B2(P3_U3151), .C1(
        n15089), .C2(n12608), .ZN(P3_U3281) );
  INV_X1 U11036 ( .A(n8694), .ZN(n8696) );
  INV_X1 U11037 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n8695) );
  NAND2_X1 U11038 ( .A1(n8696), .A2(n8695), .ZN(n8763) );
  NAND2_X1 U11039 ( .A1(n8763), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8697) );
  XNOR2_X1 U11040 ( .A(n8697), .B(P2_IR_REG_10__SCAN_IN), .ZN(n9959) );
  INV_X1 U11041 ( .A(n9959), .ZN(n14666) );
  INV_X1 U11042 ( .A(P1_DATAO_REG_10__SCAN_IN), .ZN(n8698) );
  OAI222_X1 U11043 ( .A1(n14666), .A2(P2_U3088), .B1(n13438), .B2(n8699), .C1(
        n8698), .C2(n13440), .ZN(P2_U3317) );
  XNOR2_X2 U11044 ( .A(n8701), .B(n8700), .ZN(n11991) );
  AOI21_X1 U11045 ( .B1(n8702), .B2(n8672), .A(n8671), .ZN(n8703) );
  XNOR2_X2 U11046 ( .A(n8704), .B(P2_IR_REG_29__SCAN_IN), .ZN(n8710) );
  AND2_X2 U11047 ( .A1(n11991), .A2(n8710), .ZN(n9113) );
  INV_X1 U11048 ( .A(n9113), .ZN(n11872) );
  INV_X1 U11049 ( .A(P2_REG1_REG_31__SCAN_IN), .ZN(n8707) );
  INV_X1 U11050 ( .A(n8710), .ZN(n11188) );
  AND2_X2 U11051 ( .A1(n8711), .A2(n11188), .ZN(n9115) );
  NAND2_X1 U11052 ( .A1(n11688), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n8706) );
  AND2_X2 U11053 ( .A1(n11991), .A2(n11188), .ZN(n9030) );
  NAND2_X1 U11054 ( .A1(n11123), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n8705) );
  OAI211_X1 U11055 ( .C1(n11872), .C2(n8707), .A(n8706), .B(n8705), .ZN(n13164) );
  NAND2_X1 U11056 ( .A1(n6471), .A2(n13164), .ZN(n8708) );
  OAI21_X1 U11057 ( .B1(n6471), .B2(n8709), .A(n8708), .ZN(P2_U3562) );
  NAND2_X1 U11058 ( .A1(n6485), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n8715) );
  NAND2_X1 U11059 ( .A1(n9030), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n8714) );
  NAND2_X1 U11060 ( .A1(n9113), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n8713) );
  NAND2_X1 U11061 ( .A1(n9115), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n8712) );
  NAND2_X1 U11062 ( .A1(n6471), .A2(n9437), .ZN(n8716) );
  OAI21_X1 U11063 ( .B1(n6471), .B2(n6732), .A(n8716), .ZN(P2_U3531) );
  INV_X1 U11064 ( .A(n9277), .ZN(n8717) );
  NAND2_X1 U11065 ( .A1(n8717), .A2(P1_STATE_REG_SCAN_IN), .ZN(n11616) );
  NAND2_X1 U11066 ( .A1(n9301), .A2(n11616), .ZN(n8742) );
  INV_X1 U11067 ( .A(n8720), .ZN(n8721) );
  NAND2_X1 U11068 ( .A1(n8721), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8722) );
  NAND2_X1 U11069 ( .A1(n14544), .A2(n14545), .ZN(n11538) );
  INV_X1 U11070 ( .A(n11538), .ZN(n9275) );
  NAND2_X1 U11071 ( .A1(n9275), .A2(n9277), .ZN(n8729) );
  NAND2_X1 U11072 ( .A1(n8729), .A2(n11364), .ZN(n8740) );
  AND2_X1 U11073 ( .A1(n8742), .A2(n8740), .ZN(n14497) );
  NOR2_X1 U11074 ( .A1(n14497), .A2(P1_U4016), .ZN(P1_U3085) );
  INV_X1 U11075 ( .A(P1_B_REG_SCAN_IN), .ZN(n8732) );
  NOR2_X1 U11076 ( .A1(n9253), .A2(n8732), .ZN(n8731) );
  INV_X1 U11077 ( .A(n8730), .ZN(n11085) );
  MUX2_X1 U11078 ( .A(n8732), .B(n8731), .S(n11085), .Z(n8733) );
  INV_X1 U11079 ( .A(n9301), .ZN(n8735) );
  NAND2_X1 U11080 ( .A1(n9663), .A2(n8735), .ZN(n14539) );
  INV_X1 U11081 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n8737) );
  AND2_X1 U11082 ( .A1(n8738), .A2(n14127), .ZN(n8736) );
  INV_X1 U11083 ( .A(n9253), .ZN(n14128) );
  AOI22_X1 U11084 ( .A1(n14539), .A2(n8737), .B1(n8736), .B2(n14128), .ZN(
        P1_U3446) );
  INV_X1 U11085 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n8739) );
  NOR2_X1 U11086 ( .A1(n8730), .A2(n9252), .ZN(n9660) );
  AOI22_X1 U11087 ( .A1(n14539), .A2(n8739), .B1(n8738), .B2(n9660), .ZN(
        P1_U3445) );
  INV_X1 U11088 ( .A(n14497), .ZN(n14495) );
  INV_X1 U11089 ( .A(n8740), .ZN(n8741) );
  NAND2_X1 U11090 ( .A1(n8742), .A2(n8741), .ZN(n8839) );
  INV_X1 U11091 ( .A(n8839), .ZN(n8842) );
  INV_X1 U11092 ( .A(n14121), .ZN(n12002) );
  INV_X1 U11093 ( .A(n8743), .ZN(n13680) );
  INV_X1 U11094 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n8843) );
  NAND2_X1 U11095 ( .A1(n12002), .A2(n8843), .ZN(n8744) );
  AND2_X1 U11096 ( .A1(n13680), .A2(n8744), .ZN(n13683) );
  OAI21_X1 U11097 ( .B1(n12002), .B2(P1_REG1_REG_0__SCAN_IN), .A(n13683), .ZN(
        n8745) );
  XNOR2_X1 U11098 ( .A(n8745), .B(P1_IR_REG_0__SCAN_IN), .ZN(n8746) );
  AOI22_X1 U11099 ( .A1(n8842), .A2(n8746), .B1(P1_REG3_REG_0__SCAN_IN), .B2(
        P1_U3086), .ZN(n8747) );
  OAI21_X1 U11100 ( .B1(n14495), .B2(n6676), .A(n8747), .ZN(P1_U3243) );
  NAND2_X1 U11101 ( .A1(n14685), .A2(P2_ADDR_REG_3__SCAN_IN), .ZN(n8748) );
  NAND2_X1 U11102 ( .A1(P2_U3088), .A2(P2_REG3_REG_3__SCAN_IN), .ZN(n9453) );
  OAI211_X1 U11103 ( .C1(n14667), .C2(n8749), .A(n8748), .B(n9453), .ZN(n8762)
         );
  INV_X1 U11104 ( .A(n9019), .ZN(n8754) );
  AOI22_X1 U11105 ( .A1(n8751), .A2(n8750), .B1(P2_REG1_REG_2__SCAN_IN), .B2(
        n8754), .ZN(n8753) );
  INV_X1 U11106 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n14800) );
  MUX2_X1 U11107 ( .A(n14800), .B(P2_REG1_REG_3__SCAN_IN), .S(n9098), .Z(n8752) );
  NOR2_X1 U11108 ( .A1(n8753), .A2(n8752), .ZN(n8865) );
  AOI211_X1 U11109 ( .C1(n8753), .C2(n8752), .A(n8865), .B(n14639), .ZN(n8761)
         );
  INV_X1 U11110 ( .A(n14692), .ZN(n14677) );
  NAND2_X1 U11111 ( .A1(n8754), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8757) );
  INV_X1 U11112 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n8755) );
  MUX2_X1 U11113 ( .A(n8755), .B(P2_REG2_REG_3__SCAN_IN), .S(n9098), .Z(n8756)
         );
  AOI21_X1 U11114 ( .B1(n8758), .B2(n8757), .A(n8756), .ZN(n8872) );
  AND3_X1 U11115 ( .A1(n8758), .A2(n8757), .A3(n8756), .ZN(n8759) );
  NOR3_X1 U11116 ( .A1(n14677), .A2(n8872), .A3(n8759), .ZN(n8760) );
  OR3_X1 U11117 ( .A1(n8762), .A2(n8761), .A3(n8760), .ZN(P2_U3217) );
  OAI21_X1 U11118 ( .B1(n8763), .B2(P2_IR_REG_10__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n8764) );
  XNOR2_X1 U11119 ( .A(n8764), .B(P2_IR_REG_11__SCAN_IN), .ZN(n10059) );
  INV_X1 U11120 ( .A(n10059), .ZN(n10008) );
  INV_X1 U11121 ( .A(n8765), .ZN(n8766) );
  MUX2_X1 U11122 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n11543), .Z(n8822) );
  XNOR2_X1 U11123 ( .A(n8822), .B(SI_11_), .ZN(n8825) );
  XNOR2_X1 U11124 ( .A(n8826), .B(n8825), .ZN(n10615) );
  INV_X1 U11125 ( .A(n10615), .ZN(n8785) );
  INV_X1 U11126 ( .A(P1_DATAO_REG_11__SCAN_IN), .ZN(n8769) );
  OAI222_X1 U11127 ( .A1(n10008), .A2(P2_U3088), .B1(n13438), .B2(n8785), .C1(
        n8769), .C2(n13440), .ZN(P2_U3316) );
  NAND2_X1 U11128 ( .A1(n9633), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n9851) );
  NAND2_X1 U11129 ( .A1(n9869), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n10181) );
  INV_X1 U11130 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n10684) );
  INV_X1 U11131 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n10774) );
  NAND2_X1 U11132 ( .A1(n10981), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10989) );
  INV_X1 U11133 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n10988) );
  INV_X1 U11134 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n11099) );
  NOR2_X1 U11135 ( .A1(n11101), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n8770) );
  OR2_X1 U11136 ( .A1(n11312), .A2(n8770), .ZN(n13984) );
  NAND2_X1 U11137 ( .A1(n8773), .A2(n8774), .ZN(n14112) );
  INV_X1 U11138 ( .A(n11185), .ZN(n8776) );
  NAND2_X2 U11139 ( .A1(n14120), .A2(n8776), .ZN(n9593) );
  AOI22_X1 U11140 ( .A1(n6473), .A2(P1_REG1_REG_18__SCAN_IN), .B1(n6482), .B2(
        P1_REG2_REG_18__SCAN_IN), .ZN(n8779) );
  NAND2_X1 U11141 ( .A1(n11503), .A2(P1_REG0_REG_18__SCAN_IN), .ZN(n8778) );
  OAI211_X1 U11142 ( .C1(n13984), .C2(n11470), .A(n8779), .B(n8778), .ZN(
        n13530) );
  NAND2_X1 U11143 ( .A1(n13530), .A2(P1_U4016), .ZN(n8780) );
  OAI21_X1 U11144 ( .B1(P1_U4016), .B2(n9829), .A(n8780), .ZN(P1_U3578) );
  OR2_X1 U11145 ( .A1(n8781), .A2(n14111), .ZN(n8782) );
  NAND2_X1 U11146 ( .A1(n8783), .A2(n8782), .ZN(n8827) );
  XNOR2_X1 U11147 ( .A(n8827), .B(n8784), .ZN(n13783) );
  INV_X1 U11148 ( .A(n13783), .ZN(n9526) );
  OAI222_X1 U11149 ( .A1(n8786), .A2(n14124), .B1(P1_U3086), .B2(n9526), .C1(
        n14119), .C2(n8785), .ZN(P1_U3344) );
  NOR2_X1 U11150 ( .A1(n12586), .A2(n8787), .ZN(n8790) );
  CLKBUF_X1 U11151 ( .A(n8790), .Z(n8813) );
  INV_X1 U11152 ( .A(P3_D_REG_11__SCAN_IN), .ZN(n8788) );
  NOR2_X1 U11153 ( .A1(n8813), .A2(n8788), .ZN(P3_U3254) );
  INV_X1 U11154 ( .A(P3_D_REG_2__SCAN_IN), .ZN(n8789) );
  NOR2_X1 U11155 ( .A1(n8813), .A2(n8789), .ZN(P3_U3263) );
  INV_X1 U11156 ( .A(P3_D_REG_5__SCAN_IN), .ZN(n8791) );
  NOR2_X1 U11157 ( .A1(n8813), .A2(n8791), .ZN(P3_U3260) );
  INV_X1 U11158 ( .A(P3_D_REG_10__SCAN_IN), .ZN(n8792) );
  NOR2_X1 U11159 ( .A1(n8813), .A2(n8792), .ZN(P3_U3255) );
  INV_X1 U11160 ( .A(P3_D_REG_6__SCAN_IN), .ZN(n8793) );
  NOR2_X1 U11161 ( .A1(n8813), .A2(n8793), .ZN(P3_U3259) );
  INV_X1 U11162 ( .A(P3_D_REG_9__SCAN_IN), .ZN(n8794) );
  NOR2_X1 U11163 ( .A1(n8813), .A2(n8794), .ZN(P3_U3256) );
  INV_X1 U11164 ( .A(P3_D_REG_4__SCAN_IN), .ZN(n8795) );
  NOR2_X1 U11165 ( .A1(n8813), .A2(n8795), .ZN(P3_U3261) );
  INV_X1 U11166 ( .A(P3_D_REG_12__SCAN_IN), .ZN(n8796) );
  NOR2_X1 U11167 ( .A1(n8813), .A2(n8796), .ZN(P3_U3253) );
  INV_X1 U11168 ( .A(P3_D_REG_13__SCAN_IN), .ZN(n8797) );
  NOR2_X1 U11169 ( .A1(n8813), .A2(n8797), .ZN(P3_U3252) );
  INV_X1 U11170 ( .A(P3_D_REG_14__SCAN_IN), .ZN(n8798) );
  NOR2_X1 U11171 ( .A1(n8813), .A2(n8798), .ZN(P3_U3251) );
  INV_X1 U11172 ( .A(P3_D_REG_15__SCAN_IN), .ZN(n8799) );
  NOR2_X1 U11173 ( .A1(n8813), .A2(n8799), .ZN(P3_U3250) );
  INV_X1 U11174 ( .A(P3_D_REG_16__SCAN_IN), .ZN(n8800) );
  NOR2_X1 U11175 ( .A1(n8813), .A2(n8800), .ZN(P3_U3249) );
  INV_X1 U11176 ( .A(P3_D_REG_3__SCAN_IN), .ZN(n8801) );
  NOR2_X1 U11177 ( .A1(n8813), .A2(n8801), .ZN(P3_U3262) );
  INV_X1 U11178 ( .A(P3_D_REG_17__SCAN_IN), .ZN(n8802) );
  NOR2_X1 U11179 ( .A1(n8813), .A2(n8802), .ZN(P3_U3248) );
  INV_X1 U11180 ( .A(P3_D_REG_18__SCAN_IN), .ZN(n8803) );
  NOR2_X1 U11181 ( .A1(n8813), .A2(n8803), .ZN(P3_U3247) );
  INV_X1 U11182 ( .A(P3_D_REG_19__SCAN_IN), .ZN(n8804) );
  NOR2_X1 U11183 ( .A1(n8813), .A2(n8804), .ZN(P3_U3246) );
  INV_X1 U11184 ( .A(P3_D_REG_7__SCAN_IN), .ZN(n8805) );
  NOR2_X1 U11185 ( .A1(n8813), .A2(n8805), .ZN(P3_U3258) );
  INV_X1 U11186 ( .A(P3_D_REG_20__SCAN_IN), .ZN(n8806) );
  NOR2_X1 U11187 ( .A1(n8790), .A2(n8806), .ZN(P3_U3245) );
  INV_X1 U11188 ( .A(P3_D_REG_21__SCAN_IN), .ZN(n8807) );
  NOR2_X1 U11189 ( .A1(n8790), .A2(n8807), .ZN(P3_U3244) );
  INV_X1 U11190 ( .A(P3_D_REG_22__SCAN_IN), .ZN(n8808) );
  NOR2_X1 U11191 ( .A1(n8790), .A2(n8808), .ZN(P3_U3243) );
  INV_X1 U11192 ( .A(P3_D_REG_23__SCAN_IN), .ZN(n8809) );
  NOR2_X1 U11193 ( .A1(n8790), .A2(n8809), .ZN(P3_U3242) );
  INV_X1 U11194 ( .A(P3_D_REG_24__SCAN_IN), .ZN(n8810) );
  NOR2_X1 U11195 ( .A1(n8790), .A2(n8810), .ZN(P3_U3241) );
  INV_X1 U11196 ( .A(P3_D_REG_25__SCAN_IN), .ZN(n8811) );
  NOR2_X1 U11197 ( .A1(n8790), .A2(n8811), .ZN(P3_U3240) );
  INV_X1 U11198 ( .A(P3_D_REG_8__SCAN_IN), .ZN(n8812) );
  NOR2_X1 U11199 ( .A1(n8813), .A2(n8812), .ZN(P3_U3257) );
  INV_X1 U11200 ( .A(P3_D_REG_26__SCAN_IN), .ZN(n8814) );
  NOR2_X1 U11201 ( .A1(n8790), .A2(n8814), .ZN(P3_U3239) );
  INV_X1 U11202 ( .A(P3_D_REG_27__SCAN_IN), .ZN(n8815) );
  NOR2_X1 U11203 ( .A1(n8790), .A2(n8815), .ZN(P3_U3238) );
  INV_X1 U11204 ( .A(P3_D_REG_28__SCAN_IN), .ZN(n8816) );
  NOR2_X1 U11205 ( .A1(n8790), .A2(n8816), .ZN(P3_U3237) );
  INV_X1 U11206 ( .A(P3_D_REG_29__SCAN_IN), .ZN(n8817) );
  NOR2_X1 U11207 ( .A1(n8790), .A2(n8817), .ZN(P3_U3236) );
  INV_X1 U11208 ( .A(P3_D_REG_30__SCAN_IN), .ZN(n8818) );
  NOR2_X1 U11209 ( .A1(n8790), .A2(n8818), .ZN(P3_U3235) );
  INV_X1 U11210 ( .A(P3_D_REG_31__SCAN_IN), .ZN(n8819) );
  NOR2_X1 U11211 ( .A1(n8813), .A2(n8819), .ZN(P3_U3234) );
  INV_X1 U11212 ( .A(n8820), .ZN(n8821) );
  OAI222_X1 U11213 ( .A1(n12607), .A2(n8821), .B1(n12205), .B2(P3_U3151), .C1(
        n15194), .C2(n12608), .ZN(P3_U3280) );
  INV_X1 U11214 ( .A(n8822), .ZN(n8823) );
  NAND2_X1 U11215 ( .A1(n8823), .A2(n15209), .ZN(n8824) );
  MUX2_X1 U11216 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(P1_DATAO_REG_12__SCAN_IN), 
        .S(n11543), .Z(n8962) );
  XNOR2_X1 U11217 ( .A(n8961), .B(n8960), .ZN(n10678) );
  INV_X1 U11218 ( .A(n10678), .ZN(n8888) );
  NAND2_X1 U11219 ( .A1(n8828), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8968) );
  XNOR2_X1 U11220 ( .A(n8968), .B(P1_IR_REG_12__SCAN_IN), .ZN(n14491) );
  AOI22_X1 U11221 ( .A1(n14491), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n14114), .ZN(n8829) );
  OAI21_X1 U11222 ( .B1(n8888), .B2(n14119), .A(n8829), .ZN(P1_U3343) );
  INV_X1 U11223 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n10178) );
  MUX2_X1 U11224 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n10178), .S(n8858), .Z(n8838) );
  INV_X1 U11225 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n9871) );
  INV_X1 U11226 ( .A(n13736), .ZN(n13731) );
  INV_X1 U11227 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n9303) );
  MUX2_X1 U11228 ( .A(n9303), .B(P1_REG1_REG_1__SCAN_IN), .S(n13669), .Z(n8831) );
  AND2_X1 U11229 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n8830) );
  NAND2_X1 U11230 ( .A1(n8831), .A2(n8830), .ZN(n13686) );
  INV_X1 U11231 ( .A(n13669), .ZN(n13673) );
  NAND2_X1 U11232 ( .A1(n13673), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n13685) );
  NAND2_X1 U11233 ( .A1(n13686), .A2(n13685), .ZN(n8833) );
  INV_X1 U11234 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n9564) );
  MUX2_X1 U11235 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n9564), .S(n13689), .Z(n8832) );
  NAND2_X1 U11236 ( .A1(n8833), .A2(n8832), .ZN(n13705) );
  NAND2_X1 U11237 ( .A1(n13689), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n13704) );
  NAND2_X1 U11238 ( .A1(n13705), .A2(n13704), .ZN(n8835) );
  INV_X1 U11239 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n9592) );
  MUX2_X1 U11240 ( .A(P1_REG1_REG_3__SCAN_IN), .B(n9592), .S(n13703), .Z(n8834) );
  NAND2_X1 U11241 ( .A1(n8835), .A2(n8834), .ZN(n13718) );
  NAND2_X1 U11242 ( .A1(n13703), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n13717) );
  INV_X1 U11243 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n14617) );
  MUX2_X1 U11244 ( .A(n14617), .B(P1_REG1_REG_4__SCAN_IN), .S(n13721), .Z(
        n13716) );
  AOI21_X1 U11245 ( .B1(n13718), .B2(n13717), .A(n13716), .ZN(n13715) );
  AOI21_X1 U11246 ( .B1(n13721), .B2(P1_REG1_REG_4__SCAN_IN), .A(n13715), .ZN(
        n13733) );
  INV_X1 U11247 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n14619) );
  MUX2_X1 U11248 ( .A(n14619), .B(P1_REG1_REG_5__SCAN_IN), .S(n13736), .Z(
        n13734) );
  NAND2_X1 U11249 ( .A1(n13733), .A2(n13734), .ZN(n13732) );
  OAI21_X1 U11250 ( .B1(P1_REG1_REG_5__SCAN_IN), .B2(n13731), .A(n13732), .ZN(
        n8981) );
  INV_X1 U11251 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n14621) );
  MUX2_X1 U11252 ( .A(n14621), .B(P1_REG1_REG_6__SCAN_IN), .S(n9847), .Z(n8980) );
  NOR2_X1 U11253 ( .A1(n8981), .A2(n8980), .ZN(n13755) );
  NOR2_X1 U11254 ( .A1(n8985), .A2(n14621), .ZN(n13754) );
  MUX2_X1 U11255 ( .A(P1_REG1_REG_7__SCAN_IN), .B(n9871), .S(n13747), .Z(
        n13753) );
  OAI21_X1 U11256 ( .B1(n13755), .B2(n13754), .A(n13753), .ZN(n13757) );
  OAI21_X1 U11257 ( .B1(n8836), .B2(n9871), .A(n13757), .ZN(n8837) );
  NOR2_X1 U11258 ( .A1(n8837), .A2(n8838), .ZN(n13764) );
  AOI21_X1 U11259 ( .B1(n8838), .B2(n8837), .A(n13764), .ZN(n8864) );
  INV_X1 U11260 ( .A(n8858), .ZN(n10200) );
  INV_X1 U11261 ( .A(n14501), .ZN(n14490) );
  INV_X1 U11262 ( .A(P1_ADDR_REG_8__SCAN_IN), .ZN(n14137) );
  NAND2_X1 U11263 ( .A1(P1_REG3_REG_8__SCAN_IN), .A2(P1_U3086), .ZN(n10428) );
  OAI21_X1 U11264 ( .B1(n14495), .B2(n14137), .A(n10428), .ZN(n8840) );
  AOI21_X1 U11265 ( .B1(n10200), .B2(n14490), .A(n8840), .ZN(n8863) );
  NOR2_X1 U11266 ( .A1(n8743), .A2(n14121), .ZN(n8841) );
  INV_X1 U11267 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n10303) );
  MUX2_X1 U11268 ( .A(n10303), .B(P1_REG2_REG_5__SCAN_IN), .S(n13736), .Z(
        n8852) );
  INV_X1 U11269 ( .A(P1_REG2_REG_1__SCAN_IN), .ZN(n9305) );
  MUX2_X1 U11270 ( .A(n9305), .B(P1_REG2_REG_1__SCAN_IN), .S(n13669), .Z(
        n13668) );
  NOR2_X1 U11271 ( .A1(n13671), .A2(n8843), .ZN(n13679) );
  NAND2_X1 U11272 ( .A1(n13668), .A2(n13679), .ZN(n13692) );
  NAND2_X1 U11273 ( .A1(n13673), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n13691) );
  NAND2_X1 U11274 ( .A1(n13692), .A2(n13691), .ZN(n8846) );
  INV_X1 U11275 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n8844) );
  MUX2_X1 U11276 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n8844), .S(n13689), .Z(n8845) );
  NAND2_X1 U11277 ( .A1(n8846), .A2(n8845), .ZN(n13700) );
  NAND2_X1 U11278 ( .A1(n13689), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n13699) );
  NAND2_X1 U11279 ( .A1(n13700), .A2(n13699), .ZN(n8848) );
  INV_X1 U11280 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n9591) );
  MUX2_X1 U11281 ( .A(P1_REG2_REG_3__SCAN_IN), .B(n9591), .S(n13703), .Z(n8847) );
  NAND2_X1 U11282 ( .A1(n8848), .A2(n8847), .ZN(n13713) );
  NAND2_X1 U11283 ( .A1(n13703), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n13712) );
  NAND2_X1 U11284 ( .A1(n13713), .A2(n13712), .ZN(n8850) );
  INV_X1 U11285 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n9610) );
  MUX2_X1 U11286 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n9610), .S(n13721), .Z(n8849) );
  NAND2_X1 U11287 ( .A1(n8850), .A2(n8849), .ZN(n13738) );
  NAND2_X1 U11288 ( .A1(n13721), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n13737) );
  NAND2_X1 U11289 ( .A1(n13738), .A2(n13737), .ZN(n8851) );
  NAND2_X1 U11290 ( .A1(n8852), .A2(n8851), .ZN(n13741) );
  NAND2_X1 U11291 ( .A1(n13731), .A2(P1_REG2_REG_5__SCAN_IN), .ZN(n8853) );
  NAND2_X1 U11292 ( .A1(n13741), .A2(n8853), .ZN(n8978) );
  INV_X1 U11293 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n10289) );
  MUX2_X1 U11294 ( .A(P1_REG2_REG_6__SCAN_IN), .B(n10289), .S(n9847), .Z(n8977) );
  NAND2_X1 U11295 ( .A1(n8978), .A2(n8977), .ZN(n13750) );
  NAND2_X1 U11296 ( .A1(n9847), .A2(P1_REG2_REG_6__SCAN_IN), .ZN(n13749) );
  NAND2_X1 U11297 ( .A1(n13750), .A2(n13749), .ZN(n8855) );
  INV_X1 U11298 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n10319) );
  MUX2_X1 U11299 ( .A(P1_REG2_REG_7__SCAN_IN), .B(n10319), .S(n13747), .Z(
        n8854) );
  NAND2_X1 U11300 ( .A1(n8855), .A2(n8854), .ZN(n13752) );
  NAND2_X1 U11301 ( .A1(n13747), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n8860) );
  NAND2_X1 U11302 ( .A1(n13752), .A2(n8860), .ZN(n8857) );
  INV_X1 U11303 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n10179) );
  MUX2_X1 U11304 ( .A(n10179), .B(P1_REG2_REG_8__SCAN_IN), .S(n8858), .Z(n8856) );
  NAND2_X1 U11305 ( .A1(n8857), .A2(n8856), .ZN(n13772) );
  MUX2_X1 U11306 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n10179), .S(n8858), .Z(n8859) );
  NAND3_X1 U11307 ( .A1(n13752), .A2(n8860), .A3(n8859), .ZN(n8861) );
  NAND3_X1 U11308 ( .A1(n14508), .A2(n13772), .A3(n8861), .ZN(n8862) );
  OAI211_X1 U11309 ( .C1(n8864), .C2(n13801), .A(n8863), .B(n8862), .ZN(
        P1_U3251) );
  AOI21_X1 U11310 ( .B1(n9098), .B2(P2_REG1_REG_3__SCAN_IN), .A(n8865), .ZN(
        n14642) );
  INV_X1 U11311 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n14802) );
  MUX2_X1 U11312 ( .A(n14802), .B(P2_REG1_REG_4__SCAN_IN), .S(n14638), .Z(
        n14641) );
  NOR2_X1 U11313 ( .A1(n14642), .A2(n14641), .ZN(n14640) );
  AOI21_X1 U11314 ( .B1(n14638), .B2(P2_REG1_REG_4__SCAN_IN), .A(n14640), .ZN(
        n14654) );
  INV_X1 U11315 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n14804) );
  MUX2_X1 U11316 ( .A(n14804), .B(P2_REG1_REG_5__SCAN_IN), .S(n14652), .Z(
        n14653) );
  OR2_X1 U11317 ( .A1(n14654), .A2(n14653), .ZN(n14656) );
  NAND2_X1 U11318 ( .A1(n14652), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n13090) );
  INV_X1 U11319 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n9207) );
  MUX2_X1 U11320 ( .A(n9207), .B(P2_REG1_REG_6__SCAN_IN), .S(n9191), .Z(n13089) );
  AOI21_X1 U11321 ( .B1(n14656), .B2(n13090), .A(n13089), .ZN(n13111) );
  NOR2_X1 U11322 ( .A1(n13087), .A2(n9207), .ZN(n13106) );
  INV_X1 U11323 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n8866) );
  MUX2_X1 U11324 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n8866), .S(n13105), .Z(n8867) );
  OAI21_X1 U11325 ( .B1(n13111), .B2(n13106), .A(n8867), .ZN(n13109) );
  NAND2_X1 U11326 ( .A1(n13105), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n8869) );
  INV_X1 U11327 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n14806) );
  MUX2_X1 U11328 ( .A(n14806), .B(P2_REG1_REG_8__SCAN_IN), .S(n9731), .Z(n8868) );
  AOI21_X1 U11329 ( .B1(n13109), .B2(n8869), .A(n8868), .ZN(n8987) );
  NAND3_X1 U11330 ( .A1(n13109), .A2(n8869), .A3(n8868), .ZN(n8870) );
  NAND2_X1 U11331 ( .A1(n8870), .A2(n14686), .ZN(n8884) );
  NAND2_X1 U11332 ( .A1(P2_REG3_REG_8__SCAN_IN), .A2(P2_U3088), .ZN(n9752) );
  OAI21_X1 U11333 ( .B1(n14667), .B2(n8871), .A(n9752), .ZN(n8882) );
  AOI21_X1 U11334 ( .B1(n9098), .B2(P2_REG2_REG_3__SCAN_IN), .A(n8872), .ZN(
        n14646) );
  INV_X1 U11335 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n8873) );
  MUX2_X1 U11336 ( .A(n8873), .B(P2_REG2_REG_4__SCAN_IN), .S(n14638), .Z(
        n14645) );
  AOI21_X1 U11337 ( .B1(n14638), .B2(P2_REG2_REG_4__SCAN_IN), .A(n14644), .ZN(
        n14658) );
  MUX2_X1 U11338 ( .A(n9165), .B(P2_REG2_REG_5__SCAN_IN), .S(n14652), .Z(
        n14657) );
  OR2_X1 U11339 ( .A1(n14658), .A2(n14657), .ZN(n14660) );
  NAND2_X1 U11340 ( .A1(n14652), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n13083) );
  INV_X1 U11341 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n8874) );
  MUX2_X1 U11342 ( .A(n8874), .B(P2_REG2_REG_6__SCAN_IN), .S(n9191), .Z(n13082) );
  NOR2_X1 U11343 ( .A1(n13087), .A2(n8874), .ZN(n13096) );
  INV_X1 U11344 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n8875) );
  MUX2_X1 U11345 ( .A(P2_REG2_REG_7__SCAN_IN), .B(n8875), .S(n13105), .Z(n8876) );
  OAI21_X1 U11346 ( .B1(n13101), .B2(n13096), .A(n8876), .ZN(n13099) );
  NAND2_X1 U11347 ( .A1(n13105), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n8879) );
  INV_X1 U11348 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n8877) );
  MUX2_X1 U11349 ( .A(n8877), .B(P2_REG2_REG_8__SCAN_IN), .S(n9731), .Z(n8878)
         );
  AOI21_X1 U11350 ( .B1(n13099), .B2(n8879), .A(n8878), .ZN(n8986) );
  AND3_X1 U11351 ( .A1(n13099), .A2(n8879), .A3(n8878), .ZN(n8880) );
  NOR3_X1 U11352 ( .A1(n8986), .A2(n8880), .A3(n14677), .ZN(n8881) );
  AOI211_X1 U11353 ( .C1(n14685), .C2(P2_ADDR_REG_8__SCAN_IN), .A(n8882), .B(
        n8881), .ZN(n8883) );
  OAI21_X1 U11354 ( .B1(n8987), .B2(n8884), .A(n8883), .ZN(P2_U3222) );
  NAND2_X1 U11355 ( .A1(n8974), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8887) );
  XNOR2_X1 U11356 ( .A(n8887), .B(P2_IR_REG_12__SCAN_IN), .ZN(n10129) );
  INV_X1 U11357 ( .A(n10129), .ZN(n13120) );
  OAI222_X1 U11358 ( .A1(n13440), .A2(n8889), .B1(n13438), .B2(n8888), .C1(
        n13120), .C2(P2_U3088), .ZN(P2_U3315) );
  NAND2_X4 U11359 ( .A1(n8899), .A2(n11543), .ZN(n12931) );
  NAND2_X1 U11360 ( .A1(n9097), .A2(P1_DATAO_REG_1__SCAN_IN), .ZN(n8892) );
  NAND2_X1 U11361 ( .A1(n9142), .A2(n8890), .ZN(n8891) );
  NAND2_X1 U11362 ( .A1(n9113), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8896) );
  NAND2_X1 U11363 ( .A1(n6484), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n8895) );
  NAND2_X1 U11364 ( .A1(n9030), .A2(P2_REG0_REG_1__SCAN_IN), .ZN(n8893) );
  NAND4_X4 U11365 ( .A1(n8896), .A2(n8895), .A3(n8894), .A4(n8893), .ZN(n13067) );
  INV_X1 U11366 ( .A(n12995), .ZN(n8901) );
  NAND2_X1 U11367 ( .A1(n11543), .A2(SI_0_), .ZN(n8897) );
  XNOR2_X1 U11368 ( .A(n8897), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n13441) );
  OR2_X1 U11369 ( .A1(n9437), .A2(n9441), .ZN(n9438) );
  INV_X1 U11370 ( .A(n9438), .ZN(n8900) );
  NAND2_X1 U11371 ( .A1(n12995), .A2(n9438), .ZN(n8902) );
  NAND2_X1 U11372 ( .A1(n9028), .A2(n8902), .ZN(n8926) );
  INV_X1 U11373 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n8904) );
  NAND2_X1 U11374 ( .A1(n8904), .A2(n8903), .ZN(n8906) );
  NAND2_X1 U11375 ( .A1(n9243), .A2(n8907), .ZN(n9371) );
  AND2_X1 U11376 ( .A1(P2_IR_REG_19__SCAN_IN), .A2(P2_IR_REG_31__SCAN_IN), 
        .ZN(n8908) );
  XNOR2_X1 U11377 ( .A(P2_IR_REG_19__SCAN_IN), .B(P2_IR_REG_31__SCAN_IN), .ZN(
        n8912) );
  INV_X1 U11378 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n9825) );
  INV_X1 U11379 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n8910) );
  NAND3_X1 U11380 ( .A1(n9825), .A2(n8910), .A3(P2_IR_REG_19__SCAN_IN), .ZN(
        n8911) );
  AND2_X1 U11381 ( .A1(n8912), .A2(n8911), .ZN(n8913) );
  INV_X1 U11382 ( .A(n12720), .ZN(n13031) );
  NAND2_X1 U11383 ( .A1(n12988), .A2(n13031), .ZN(n12935) );
  INV_X1 U11384 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n8916) );
  NAND2_X1 U11385 ( .A1(n8931), .A2(n13026), .ZN(n8918) );
  INV_X1 U11386 ( .A(n9437), .ZN(n12725) );
  INV_X1 U11387 ( .A(n8677), .ZN(n8919) );
  NAND2_X1 U11388 ( .A1(n9324), .A2(n8919), .ZN(n14322) );
  OR2_X1 U11389 ( .A1(n12725), .A2(n14322), .ZN(n8925) );
  NAND2_X1 U11390 ( .A1(n9145), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n8923) );
  NAND2_X1 U11391 ( .A1(n9030), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n8922) );
  NAND2_X1 U11392 ( .A1(n9115), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n8921) );
  NAND2_X1 U11393 ( .A1(n9113), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n8920) );
  NAND4_X2 U11394 ( .A1(n8923), .A2(n8922), .A3(n8921), .A4(n8920), .ZN(n13066) );
  NAND2_X1 U11395 ( .A1(n13066), .A2(n12711), .ZN(n8924) );
  NAND2_X1 U11396 ( .A1(n8925), .A2(n8924), .ZN(n11983) );
  AOI21_X1 U11397 ( .B1(n8926), .B2(n14740), .A(n11983), .ZN(n9384) );
  NAND2_X1 U11398 ( .A1(n8928), .A2(n14714), .ZN(n8929) );
  OR2_X1 U11399 ( .A1(n8929), .A2(n9026), .ZN(n9379) );
  NAND2_X1 U11400 ( .A1(n12988), .A2(n12720), .ZN(n12723) );
  NAND2_X1 U11401 ( .A1(n12720), .A2(n7478), .ZN(n9313) );
  OAI21_X2 U11402 ( .B1(n12723), .B2(n8931), .A(n9313), .ZN(n14788) );
  AND2_X1 U11403 ( .A1(n9379), .A2(n8930), .ZN(n8935) );
  OR2_X1 U11404 ( .A1(n12725), .A2(n9441), .ZN(n9020) );
  XNOR2_X1 U11405 ( .A(n12995), .B(n9020), .ZN(n9377) );
  INV_X1 U11406 ( .A(n9327), .ZN(n12722) );
  XNOR2_X1 U11407 ( .A(n12722), .B(n12720), .ZN(n8932) );
  INV_X1 U11408 ( .A(n9328), .ZN(n14741) );
  NAND2_X1 U11409 ( .A1(n9377), .A2(n14741), .ZN(n8934) );
  INV_X1 U11410 ( .A(n14793), .ZN(n14761) );
  NAND2_X1 U11411 ( .A1(n9377), .A2(n14761), .ZN(n8933) );
  AND4_X1 U11412 ( .A1(n9384), .A2(n8935), .A3(n8934), .A4(n8933), .ZN(n14751)
         );
  XNOR2_X1 U11413 ( .A(n11087), .B(P2_B_REG_SCAN_IN), .ZN(n8936) );
  AND2_X1 U11414 ( .A1(n8936), .A2(n13437), .ZN(n8937) );
  INV_X1 U11415 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n14739) );
  NAND2_X1 U11416 ( .A1(n14732), .A2(n14739), .ZN(n8939) );
  NAND2_X1 U11417 ( .A1(n13435), .A2(n13437), .ZN(n8938) );
  NAND2_X1 U11418 ( .A1(n8939), .A2(n8938), .ZN(n9094) );
  AND2_X1 U11419 ( .A1(n9094), .A2(n14736), .ZN(n14737) );
  NOR2_X1 U11420 ( .A1(P2_D_REG_2__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .ZN(
        n8944) );
  NOR4_X1 U11421 ( .A1(P2_D_REG_29__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_4__SCAN_IN), .A4(P2_D_REG_5__SCAN_IN), .ZN(n8943) );
  NOR4_X1 U11422 ( .A1(P2_D_REG_10__SCAN_IN), .A2(P2_D_REG_11__SCAN_IN), .A3(
        P2_D_REG_12__SCAN_IN), .A4(P2_D_REG_13__SCAN_IN), .ZN(n8942) );
  NOR4_X1 U11423 ( .A1(P2_D_REG_6__SCAN_IN), .A2(P2_D_REG_7__SCAN_IN), .A3(
        P2_D_REG_8__SCAN_IN), .A4(P2_D_REG_9__SCAN_IN), .ZN(n8941) );
  AND4_X1 U11424 ( .A1(n8944), .A2(n8943), .A3(n8942), .A4(n8941), .ZN(n8950)
         );
  NOR4_X1 U11425 ( .A1(P2_D_REG_18__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_20__SCAN_IN), .A4(P2_D_REG_21__SCAN_IN), .ZN(n8948) );
  NOR4_X1 U11426 ( .A1(P2_D_REG_16__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_15__SCAN_IN), .A4(P2_D_REG_17__SCAN_IN), .ZN(n8947) );
  NOR4_X1 U11427 ( .A1(P2_D_REG_26__SCAN_IN), .A2(P2_D_REG_27__SCAN_IN), .A3(
        P2_D_REG_28__SCAN_IN), .A4(P2_D_REG_31__SCAN_IN), .ZN(n8946) );
  NOR4_X1 U11428 ( .A1(P2_D_REG_22__SCAN_IN), .A2(P2_D_REG_23__SCAN_IN), .A3(
        P2_D_REG_24__SCAN_IN), .A4(P2_D_REG_25__SCAN_IN), .ZN(n8945) );
  AND4_X1 U11429 ( .A1(n8948), .A2(n8947), .A3(n8946), .A4(n8945), .ZN(n8949)
         );
  NAND2_X1 U11430 ( .A1(n8950), .A2(n8949), .ZN(n8951) );
  NAND2_X1 U11431 ( .A1(n14732), .A2(n8951), .ZN(n9310) );
  NAND2_X1 U11432 ( .A1(n13253), .A2(n8952), .ZN(n9314) );
  AND2_X1 U11433 ( .A1(n9314), .A2(n8931), .ZN(n12934) );
  INV_X1 U11434 ( .A(n12934), .ZN(n8953) );
  NAND2_X1 U11435 ( .A1(n9310), .A2(n13027), .ZN(n9093) );
  NOR2_X1 U11436 ( .A1(n9093), .A2(n9315), .ZN(n8954) );
  INV_X1 U11437 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n14734) );
  NAND2_X1 U11438 ( .A1(n14732), .A2(n14734), .ZN(n8956) );
  NAND2_X1 U11439 ( .A1(n13435), .A2(n11087), .ZN(n8955) );
  NAND2_X1 U11440 ( .A1(n14808), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n8957) );
  OAI21_X1 U11441 ( .B1(n14751), .B2(n14808), .A(n8957), .ZN(P2_U3500) );
  INV_X1 U11442 ( .A(n8958), .ZN(n8959) );
  OAI222_X1 U11443 ( .A1(n12607), .A2(n8959), .B1(n12222), .B2(P3_U3151), .C1(
        n15144), .C2(n12589), .ZN(P3_U3279) );
  INV_X1 U11444 ( .A(n8962), .ZN(n8963) );
  NAND2_X1 U11445 ( .A1(n8963), .A2(n15174), .ZN(n8964) );
  MUX2_X1 U11446 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(P1_DATAO_REG_13__SCAN_IN), 
        .S(n11543), .Z(n9124) );
  XNOR2_X1 U11447 ( .A(n9124), .B(n15203), .ZN(n8966) );
  XNOR2_X1 U11448 ( .A(n9127), .B(n8966), .ZN(n10765) );
  INV_X1 U11449 ( .A(n10765), .ZN(n8976) );
  NAND2_X1 U11450 ( .A1(n8968), .A2(n8967), .ZN(n8969) );
  NAND2_X1 U11451 ( .A1(n8969), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n8971) );
  NAND2_X1 U11452 ( .A1(n8971), .A2(n8970), .ZN(n9130) );
  OR2_X1 U11453 ( .A1(n8971), .A2(n8970), .ZN(n8972) );
  INV_X1 U11454 ( .A(n10766), .ZN(n14500) );
  OAI222_X1 U11455 ( .A1(n14124), .A2(n7292), .B1(n14119), .B2(n8976), .C1(
        n14500), .C2(P1_U3086), .ZN(P1_U3342) );
  OR2_X1 U11456 ( .A1(n8974), .A2(P2_IR_REG_12__SCAN_IN), .ZN(n9212) );
  NAND2_X1 U11457 ( .A1(n9212), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n8975) );
  XNOR2_X1 U11458 ( .A(n8973), .B(n8975), .ZN(n10247) );
  OAI222_X1 U11459 ( .A1(P2_U3088), .A2(n10247), .B1(n13440), .B2(n7289), .C1(
        n13438), .C2(n8976), .ZN(P2_U3314) );
  NAND2_X1 U11460 ( .A1(P1_REG3_REG_6__SCAN_IN), .A2(P1_U3086), .ZN(n9877) );
  OAI211_X1 U11461 ( .C1(n8978), .C2(n8977), .A(n14508), .B(n13750), .ZN(n8979) );
  NAND2_X1 U11462 ( .A1(n9877), .A2(n8979), .ZN(n8983) );
  AOI211_X1 U11463 ( .C1(n8981), .C2(n8980), .A(n13755), .B(n13801), .ZN(n8982) );
  AOI211_X1 U11464 ( .C1(n14497), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n8983), .B(
        n8982), .ZN(n8984) );
  OAI21_X1 U11465 ( .B1(n8985), .B2(n14501), .A(n8984), .ZN(P1_U3249) );
  AOI21_X1 U11466 ( .B1(n9731), .B2(P2_REG2_REG_8__SCAN_IN), .A(n8986), .ZN(
        n8992) );
  INV_X1 U11467 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n8990) );
  NOR3_X1 U11468 ( .A1(n8992), .A2(n8990), .A3(n14677), .ZN(n8989) );
  INV_X1 U11469 ( .A(n14667), .ZN(n14691) );
  AOI21_X1 U11470 ( .B1(n9731), .B2(P2_REG1_REG_8__SCAN_IN), .A(n8987), .ZN(
        n8997) );
  INV_X1 U11471 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10023) );
  NOR3_X1 U11472 ( .A1(n8997), .A2(n10023), .A3(n14639), .ZN(n8988) );
  NOR3_X1 U11473 ( .A1(n8989), .A2(n14691), .A3(n8988), .ZN(n9001) );
  AND2_X1 U11474 ( .A1(P2_U3088), .A2(P2_REG3_REG_9__SCAN_IN), .ZN(n8995) );
  MUX2_X1 U11475 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n8990), .S(n9786), .Z(n8991)
         );
  NAND2_X1 U11476 ( .A1(n8992), .A2(n8991), .ZN(n9085) );
  OR3_X1 U11477 ( .A1(n8992), .A2(P2_REG2_REG_9__SCAN_IN), .A3(n9786), .ZN(
        n8993) );
  AOI21_X1 U11478 ( .B1(n9085), .B2(n8993), .A(n14677), .ZN(n8994) );
  AOI211_X1 U11479 ( .C1(n14685), .C2(P2_ADDR_REG_9__SCAN_IN), .A(n8995), .B(
        n8994), .ZN(n9000) );
  NOR3_X1 U11480 ( .A1(n8997), .A2(P2_REG1_REG_9__SCAN_IN), .A3(n9786), .ZN(
        n8998) );
  MUX2_X1 U11481 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10023), .S(n9786), .Z(n8996) );
  OAI21_X1 U11482 ( .B1(n8998), .B2(n9079), .A(n14686), .ZN(n8999) );
  OAI211_X1 U11483 ( .C1(n9001), .C2(n9080), .A(n9000), .B(n8999), .ZN(
        P2_U3223) );
  INV_X1 U11484 ( .A(n10457), .ZN(n9016) );
  NAND2_X1 U11485 ( .A1(n10200), .A2(P1_REG2_REG_8__SCAN_IN), .ZN(n13771) );
  NAND2_X1 U11486 ( .A1(n13772), .A2(n13771), .ZN(n9003) );
  INV_X1 U11487 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n10238) );
  MUX2_X1 U11488 ( .A(P1_REG2_REG_9__SCAN_IN), .B(n10238), .S(n13769), .Z(
        n9002) );
  NAND2_X1 U11489 ( .A1(n9003), .A2(n9002), .ZN(n13774) );
  NAND2_X1 U11490 ( .A1(n13769), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n9007) );
  NAND2_X1 U11491 ( .A1(n13774), .A2(n9007), .ZN(n9005) );
  INV_X1 U11492 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n10227) );
  MUX2_X1 U11493 ( .A(P1_REG2_REG_10__SCAN_IN), .B(n10227), .S(n10457), .Z(
        n9004) );
  NAND2_X1 U11494 ( .A1(n9005), .A2(n9004), .ZN(n13786) );
  MUX2_X1 U11495 ( .A(n10227), .B(P1_REG2_REG_10__SCAN_IN), .S(n10457), .Z(
        n9006) );
  NAND3_X1 U11496 ( .A1(n13774), .A2(n9007), .A3(n9006), .ZN(n9008) );
  NAND3_X1 U11497 ( .A1(n14508), .A2(n13786), .A3(n9008), .ZN(n9015) );
  NAND2_X1 U11498 ( .A1(P1_REG3_REG_10__SCAN_IN), .A2(P1_U3086), .ZN(n10850)
         );
  INV_X1 U11499 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n14628) );
  MUX2_X1 U11500 ( .A(n14628), .B(P1_REG1_REG_10__SCAN_IN), .S(n10457), .Z(
        n9010) );
  NOR2_X1 U11501 ( .A1(n10200), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n13762) );
  INV_X1 U11502 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n14625) );
  MUX2_X1 U11503 ( .A(P1_REG1_REG_9__SCAN_IN), .B(n14625), .S(n13769), .Z(
        n13763) );
  OAI21_X1 U11504 ( .B1(n13764), .B2(n13762), .A(n13763), .ZN(n13761) );
  OAI21_X1 U11505 ( .B1(n13769), .B2(P1_REG1_REG_9__SCAN_IN), .A(n13761), .ZN(
        n9009) );
  NOR2_X1 U11506 ( .A1(n9009), .A2(n9010), .ZN(n9525) );
  AOI211_X1 U11507 ( .C1(n9010), .C2(n9009), .A(n9525), .B(n13801), .ZN(n9011)
         );
  INV_X1 U11508 ( .A(n9011), .ZN(n9012) );
  NAND2_X1 U11509 ( .A1(n10850), .A2(n9012), .ZN(n9013) );
  AOI21_X1 U11510 ( .B1(n14497), .B2(P1_ADDR_REG_10__SCAN_IN), .A(n9013), .ZN(
        n9014) );
  OAI211_X1 U11511 ( .C1(n14501), .C2(n9016), .A(n9015), .B(n9014), .ZN(
        P1_U3253) );
  INV_X1 U11512 ( .A(n12931), .ZN(n9018) );
  INV_X1 U11513 ( .A(n13067), .ZN(n9035) );
  NAND2_X1 U11514 ( .A1(n9035), .A2(n9021), .ZN(n9022) );
  NAND2_X1 U11515 ( .A1(n9023), .A2(n9022), .ZN(n9102) );
  XNOR2_X1 U11516 ( .A(n9101), .B(n9102), .ZN(n14726) );
  AND2_X1 U11517 ( .A1(n9026), .A2(n9024), .ZN(n9107) );
  INV_X1 U11518 ( .A(n9107), .ZN(n9025) );
  OAI211_X1 U11519 ( .C1(n9024), .C2(n9026), .A(n9025), .B(n14714), .ZN(n14723) );
  OAI21_X1 U11520 ( .B1(n9024), .B2(n14774), .A(n14723), .ZN(n9038) );
  NAND2_X1 U11521 ( .A1(n9028), .A2(n9027), .ZN(n9110) );
  INV_X1 U11522 ( .A(n9101), .ZN(n9109) );
  XNOR2_X1 U11523 ( .A(n9110), .B(n9109), .ZN(n9036) );
  INV_X1 U11524 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n9029) );
  NAND2_X1 U11525 ( .A1(n9145), .A2(n9029), .ZN(n9034) );
  NAND2_X1 U11526 ( .A1(n11701), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n9033) );
  NAND2_X1 U11527 ( .A1(n9115), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n9032) );
  NAND2_X1 U11528 ( .A1(n11123), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n9031) );
  NAND4_X2 U11529 ( .A1(n9034), .A2(n9033), .A3(n9032), .A4(n9031), .ZN(n13065) );
  INV_X1 U11530 ( .A(n13065), .ZN(n9153) );
  INV_X1 U11531 ( .A(n12711), .ZN(n14324) );
  OAI22_X1 U11532 ( .A1(n9035), .A2(n14322), .B1(n9153), .B2(n14324), .ZN(
        n9322) );
  AOI21_X1 U11533 ( .B1(n9036), .B2(n14740), .A(n9322), .ZN(n14730) );
  INV_X1 U11534 ( .A(n14730), .ZN(n9037) );
  AOI211_X1 U11535 ( .C1(n14726), .C2(n14768), .A(n9038), .B(n9037), .ZN(
        n14753) );
  NAND2_X1 U11536 ( .A1(n14808), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n9039) );
  OAI21_X1 U11537 ( .B1(n14753), .B2(n14808), .A(n9039), .ZN(P2_U3501) );
  OAI21_X1 U11538 ( .B1(n9042), .B2(n9041), .A(n9040), .ZN(n9043) );
  NAND2_X1 U11539 ( .A1(n9043), .A2(n14843), .ZN(n9057) );
  AOI21_X1 U11540 ( .B1(n9046), .B2(n9045), .A(n9044), .ZN(n9049) );
  NAND2_X1 U11541 ( .A1(P3_U3151), .A2(P3_REG3_REG_2__SCAN_IN), .ZN(n9048) );
  NAND2_X1 U11542 ( .A1(n14869), .A2(P3_ADDR_REG_2__SCAN_IN), .ZN(n9047) );
  OAI211_X1 U11543 ( .C1(n14887), .C2(n9049), .A(n9048), .B(n9047), .ZN(n9055)
         );
  AOI21_X1 U11544 ( .B1(n9052), .B2(n9051), .A(n9050), .ZN(n9053) );
  NOR2_X1 U11545 ( .A1(n14893), .A2(n9053), .ZN(n9054) );
  NOR2_X1 U11546 ( .A1(n9055), .A2(n9054), .ZN(n9056) );
  OAI211_X1 U11547 ( .C1(n14878), .C2(n9058), .A(n9057), .B(n9056), .ZN(
        P3_U3184) );
  INV_X1 U11548 ( .A(n9059), .ZN(n9061) );
  OAI222_X1 U11549 ( .A1(n12607), .A2(n9061), .B1(n9060), .B2(P3_U3151), .C1(
        n15072), .C2(n12589), .ZN(P3_U3278) );
  AOI21_X1 U11550 ( .B1(n9064), .B2(n9063), .A(n9062), .ZN(n9065) );
  NOR2_X1 U11551 ( .A1(n14893), .A2(n9065), .ZN(n9071) );
  AOI21_X1 U11552 ( .B1(n15026), .B2(n9067), .A(n9066), .ZN(n9069) );
  NAND2_X1 U11553 ( .A1(P3_U3151), .A2(P3_REG3_REG_3__SCAN_IN), .ZN(n9987) );
  NAND2_X1 U11554 ( .A1(n14869), .A2(P3_ADDR_REG_3__SCAN_IN), .ZN(n9068) );
  OAI211_X1 U11555 ( .C1(n14887), .C2(n9069), .A(n9987), .B(n9068), .ZN(n9070)
         );
  AOI211_X1 U11556 ( .C1(n14846), .C2(n9072), .A(n9071), .B(n9070), .ZN(n9078)
         );
  OAI21_X1 U11557 ( .B1(n9075), .B2(n9074), .A(n9073), .ZN(n9076) );
  NAND2_X1 U11558 ( .A1(n9076), .A2(n14843), .ZN(n9077) );
  NAND2_X1 U11559 ( .A1(n9078), .A2(n9077), .ZN(P3_U3185) );
  AOI21_X1 U11560 ( .B1(n10023), .B2(n9080), .A(n9079), .ZN(n14675) );
  INV_X1 U11561 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n9081) );
  MUX2_X1 U11562 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n9081), .S(n9959), .Z(
        n14674) );
  NAND2_X1 U11563 ( .A1(n14675), .A2(n14674), .ZN(n14673) );
  NAND2_X1 U11564 ( .A1(n9959), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9083) );
  INV_X1 U11565 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n10451) );
  MUX2_X1 U11566 ( .A(n10451), .B(P2_REG1_REG_11__SCAN_IN), .S(n10059), .Z(
        n9082) );
  AOI21_X1 U11567 ( .B1(n14673), .B2(n9083), .A(n9082), .ZN(n10001) );
  NAND3_X1 U11568 ( .A1(n14673), .A2(n9083), .A3(n9082), .ZN(n9084) );
  NAND2_X1 U11569 ( .A1(n9084), .A2(n14686), .ZN(n9092) );
  OAI21_X1 U11570 ( .B1(n9786), .B2(P2_REG2_REG_9__SCAN_IN), .A(n9085), .ZN(
        n14678) );
  MUX2_X1 U11571 ( .A(n10050), .B(P2_REG2_REG_10__SCAN_IN), .S(n9959), .Z(
        n14679) );
  AOI21_X1 U11572 ( .B1(P2_REG2_REG_10__SCAN_IN), .B2(n9959), .A(n14676), .ZN(
        n9087) );
  INV_X1 U11573 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n10007) );
  MUX2_X1 U11574 ( .A(P2_REG2_REG_11__SCAN_IN), .B(n10007), .S(n10059), .Z(
        n9086) );
  NAND2_X1 U11575 ( .A1(n9087), .A2(n9086), .ZN(n13117) );
  OAI21_X1 U11576 ( .B1(n9087), .B2(n9086), .A(n13117), .ZN(n9088) );
  NAND2_X1 U11577 ( .A1(n9088), .A2(n14692), .ZN(n9091) );
  NAND2_X1 U11578 ( .A1(P2_U3088), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n10405)
         );
  OAI21_X1 U11579 ( .B1(n14667), .B2(n10008), .A(n10405), .ZN(n9089) );
  AOI21_X1 U11580 ( .B1(n14685), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n9089), .ZN(
        n9090) );
  OAI211_X1 U11581 ( .C1(n10001), .C2(n9092), .A(n9091), .B(n9090), .ZN(
        P2_U3225) );
  INV_X1 U11582 ( .A(n9093), .ZN(n9095) );
  INV_X1 U11583 ( .A(n9094), .ZN(n9311) );
  NAND4_X1 U11584 ( .A1(n9095), .A2(n9311), .A3(n14736), .A4(n14735), .ZN(
        n9105) );
  INV_X2 U11585 ( .A(n13316), .ZN(n14731) );
  NOR2_X1 U11586 ( .A1(n12721), .A2(n14741), .ZN(n9096) );
  INV_X2 U11587 ( .A(n12931), .ZN(n11860) );
  NAND2_X1 U11588 ( .A1(n9600), .A2(n11860), .ZN(n9100) );
  AOI22_X1 U11589 ( .A1(n9097), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n9142), .B2(
        n9098), .ZN(n9099) );
  XNOR2_X2 U11590 ( .A(n12759), .B(n13065), .ZN(n12998) );
  NAND2_X1 U11591 ( .A1(n9102), .A2(n9101), .ZN(n9104) );
  INV_X1 U11592 ( .A(n13066), .ZN(n9120) );
  NAND2_X1 U11593 ( .A1(n9120), .A2(n9024), .ZN(n9103) );
  NAND2_X1 U11594 ( .A1(n9104), .A2(n9103), .ZN(n9137) );
  XNOR2_X1 U11595 ( .A(n12998), .B(n9137), .ZN(n14757) );
  INV_X1 U11596 ( .A(n12759), .ZN(n14755) );
  INV_X1 U11597 ( .A(n14715), .ZN(n9106) );
  OAI211_X1 U11598 ( .C1(n14755), .C2(n9107), .A(n9106), .B(n14714), .ZN(
        n14754) );
  OAI22_X1 U11599 ( .A1(n13282), .A2(n14754), .B1(P2_REG3_REG_3__SCAN_IN), 
        .B2(n14706), .ZN(n9108) );
  AOI21_X1 U11600 ( .B1(n14341), .B2(n12759), .A(n9108), .ZN(n9123) );
  NAND2_X1 U11601 ( .A1(n9110), .A2(n9109), .ZN(n9112) );
  NAND2_X1 U11602 ( .A1(n9120), .A2(n12740), .ZN(n9111) );
  NAND2_X1 U11603 ( .A1(n9112), .A2(n9111), .ZN(n9152) );
  XNOR2_X1 U11604 ( .A(n9152), .B(n12998), .ZN(n9121) );
  NAND2_X1 U11605 ( .A1(n11123), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n9119) );
  NAND2_X1 U11606 ( .A1(n11701), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n9118) );
  NOR2_X1 U11607 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_REG3_REG_3__SCAN_IN), 
        .ZN(n9114) );
  NOR2_X1 U11608 ( .A1(n9146), .A2(n9114), .ZN(n9690) );
  NAND2_X1 U11609 ( .A1(n9145), .A2(n9690), .ZN(n9117) );
  NAND2_X1 U11610 ( .A1(n9115), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n9116) );
  INV_X1 U11611 ( .A(n13064), .ZN(n9156) );
  OAI22_X1 U11612 ( .A1(n9120), .A2(n14322), .B1(n9156), .B2(n14324), .ZN(
        n9452) );
  AOI21_X1 U11613 ( .B1(n9121), .B2(n14740), .A(n9452), .ZN(n14756) );
  MUX2_X1 U11614 ( .A(n8755), .B(n14756), .S(n13316), .Z(n9122) );
  OAI211_X1 U11615 ( .C1(n13304), .C2(n14757), .A(n9123), .B(n9122), .ZN(
        P2_U3262) );
  NOR2_X1 U11616 ( .A1(n9124), .A2(SI_13_), .ZN(n9126) );
  NAND2_X1 U11617 ( .A1(n9124), .A2(SI_13_), .ZN(n9125) );
  NAND2_X1 U11618 ( .A1(n9232), .A2(SI_14_), .ZN(n9129) );
  MUX2_X1 U11619 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(P1_DATAO_REG_14__SCAN_IN), 
        .S(n11543), .Z(n9348) );
  INV_X1 U11620 ( .A(n10970), .ZN(n9214) );
  NAND2_X1 U11621 ( .A1(n9130), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9131) );
  XNOR2_X1 U11622 ( .A(n9131), .B(P1_IR_REG_14__SCAN_IN), .ZN(n10971) );
  AOI22_X1 U11623 ( .A1(n10971), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(n14114), .ZN(n9132) );
  OAI21_X1 U11624 ( .B1(n9214), .B2(n14119), .A(n9132), .ZN(P1_U3341) );
  INV_X1 U11625 ( .A(n9133), .ZN(n9135) );
  OAI222_X1 U11626 ( .A1(n12607), .A2(n9135), .B1(n9134), .B2(P3_U3151), .C1(
        n9821), .C2(n12608), .ZN(P3_U3277) );
  INV_X1 U11627 ( .A(n12998), .ZN(n9136) );
  OR2_X1 U11628 ( .A1(n13065), .A2(n12759), .ZN(n9138) );
  INV_X2 U11629 ( .A(n12931), .ZN(n12943) );
  NAND2_X1 U11630 ( .A1(n9621), .A2(n12943), .ZN(n9140) );
  AOI22_X1 U11631 ( .A1(n9097), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n9142), .B2(
        n14638), .ZN(n9139) );
  NAND2_X1 U11632 ( .A1(n9140), .A2(n9139), .ZN(n12754) );
  INV_X1 U11633 ( .A(n14701), .ZN(n14712) );
  OR2_X1 U11634 ( .A1(n12754), .A2(n13064), .ZN(n9141) );
  NAND2_X1 U11635 ( .A1(n9841), .A2(n12943), .ZN(n9144) );
  AOI22_X1 U11636 ( .A1(n9097), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n9142), .B2(
        n14652), .ZN(n9143) );
  NAND2_X1 U11637 ( .A1(n9144), .A2(n9143), .ZN(n12773) );
  NAND2_X1 U11638 ( .A1(n11701), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n9151) );
  NAND2_X1 U11639 ( .A1(n11688), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n9150) );
  NOR2_X1 U11640 ( .A1(n9146), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n9147) );
  NOR2_X1 U11641 ( .A1(n9157), .A2(n9147), .ZN(n9166) );
  NAND2_X1 U11642 ( .A1(n9145), .A2(n9166), .ZN(n9149) );
  NAND2_X1 U11643 ( .A1(n11123), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n9148) );
  XNOR2_X1 U11644 ( .A(n12773), .B(n9188), .ZN(n13000) );
  INV_X1 U11645 ( .A(n13000), .ZN(n9186) );
  XNOR2_X1 U11646 ( .A(n9196), .B(n9186), .ZN(n14776) );
  INV_X1 U11647 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n9165) );
  NAND2_X1 U11648 ( .A1(n9152), .A2(n12998), .ZN(n9155) );
  NAND2_X1 U11649 ( .A1(n9153), .A2(n12759), .ZN(n9154) );
  XNOR2_X1 U11650 ( .A(n9187), .B(n9186), .ZN(n9164) );
  NAND2_X1 U11651 ( .A1(n11123), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n9162) );
  NAND2_X1 U11652 ( .A1(n11701), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n9161) );
  NOR2_X1 U11653 ( .A1(n9157), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n9158) );
  NOR2_X1 U11654 ( .A1(n9198), .A2(n9158), .ZN(n9712) );
  NAND2_X1 U11655 ( .A1(n9145), .A2(n9712), .ZN(n9160) );
  NAND2_X1 U11656 ( .A1(n11688), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n9159) );
  NAND4_X1 U11657 ( .A1(n9162), .A2(n9161), .A3(n9160), .A4(n9159), .ZN(n13062) );
  AOI22_X1 U11658 ( .A1(n12710), .A2(n13064), .B1(n13062), .B2(n12711), .ZN(
        n9702) );
  INV_X1 U11659 ( .A(n9702), .ZN(n9163) );
  AOI21_X1 U11660 ( .B1(n9164), .B2(n14740), .A(n9163), .ZN(n14773) );
  MUX2_X1 U11661 ( .A(n9165), .B(n14773), .S(n13316), .Z(n9169) );
  INV_X1 U11662 ( .A(n12754), .ZN(n14764) );
  NAND2_X1 U11663 ( .A1(n14715), .A2(n14764), .ZN(n14713) );
  AOI211_X1 U11664 ( .C1(n12773), .C2(n14713), .A(n9329), .B(n9197), .ZN(
        n14771) );
  INV_X1 U11665 ( .A(n12773), .ZN(n14775) );
  INV_X1 U11666 ( .A(n9166), .ZN(n9706) );
  OAI22_X1 U11667 ( .A1(n14721), .A2(n14775), .B1(n9706), .B2(n14706), .ZN(
        n9167) );
  AOI21_X1 U11668 ( .B1(n14771), .B2(n14725), .A(n9167), .ZN(n9168) );
  OAI211_X1 U11669 ( .C1(n13304), .C2(n14776), .A(n9169), .B(n9168), .ZN(
        P2_U3260) );
  OAI21_X1 U11670 ( .B1(n9172), .B2(n9171), .A(n9170), .ZN(n9173) );
  NAND2_X1 U11671 ( .A1(n9173), .A2(n14843), .ZN(n9184) );
  AOI21_X1 U11672 ( .B1(n6612), .B2(n9175), .A(n9174), .ZN(n9177) );
  NAND2_X1 U11673 ( .A1(P3_U3151), .A2(P3_REG3_REG_4__SCAN_IN), .ZN(n10097) );
  NAND2_X1 U11674 ( .A1(n14869), .A2(P3_ADDR_REG_4__SCAN_IN), .ZN(n9176) );
  OAI211_X1 U11675 ( .C1(n14887), .C2(n9177), .A(n10097), .B(n9176), .ZN(n9182) );
  AOI21_X1 U11676 ( .B1(n6613), .B2(n9179), .A(n9178), .ZN(n9180) );
  NOR2_X1 U11677 ( .A1(n14893), .A2(n9180), .ZN(n9181) );
  NOR2_X1 U11678 ( .A1(n9182), .A2(n9181), .ZN(n9183) );
  OAI211_X1 U11679 ( .C1(n14878), .C2(n9185), .A(n9184), .B(n9183), .ZN(
        P3_U3186) );
  NAND2_X1 U11680 ( .A1(n12773), .A2(n9188), .ZN(n9189) );
  NAND2_X1 U11681 ( .A1(n9190), .A2(n9189), .ZN(n9402) );
  OR2_X1 U11682 ( .A1(n9845), .A2(n12931), .ZN(n9193) );
  AOI22_X1 U11683 ( .A1(n9097), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n9142), .B2(
        n9191), .ZN(n9192) );
  XNOR2_X1 U11684 ( .A(n12776), .B(n13062), .ZN(n12996) );
  INV_X1 U11685 ( .A(n12996), .ZN(n9415) );
  XNOR2_X1 U11686 ( .A(n9402), .B(n9415), .ZN(n9448) );
  NOR2_X1 U11687 ( .A1(n12773), .A2(n13063), .ZN(n9195) );
  NAND2_X1 U11688 ( .A1(n12773), .A2(n13063), .ZN(n9194) );
  OAI21_X2 U11689 ( .B1(n9196), .B2(n9195), .A(n9194), .ZN(n9416) );
  XNOR2_X1 U11690 ( .A(n9416), .B(n12996), .ZN(n9446) );
  INV_X1 U11691 ( .A(n12776), .ZN(n9203) );
  OAI211_X1 U11692 ( .C1(n9197), .C2(n9203), .A(n14714), .B(n9414), .ZN(n9444)
         );
  NAND2_X1 U11693 ( .A1(n11701), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n9202) );
  NAND2_X1 U11694 ( .A1(n11123), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n9201) );
  OAI21_X1 U11695 ( .B1(n9198), .B2(P2_REG3_REG_7__SCAN_IN), .A(n9744), .ZN(
        n9484) );
  INV_X1 U11696 ( .A(n9484), .ZN(n9426) );
  NAND2_X1 U11697 ( .A1(n9145), .A2(n9426), .ZN(n9200) );
  NAND2_X1 U11698 ( .A1(n11688), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n9199) );
  NAND4_X1 U11699 ( .A1(n9202), .A2(n9201), .A3(n9200), .A4(n9199), .ZN(n13061) );
  AOI22_X1 U11700 ( .A1(n12711), .A2(n13061), .B1(n13063), .B2(n12710), .ZN(
        n9710) );
  OAI211_X1 U11701 ( .C1(n9203), .C2(n14774), .A(n9444), .B(n9710), .ZN(n9204)
         );
  AOI21_X1 U11702 ( .B1(n9446), .B2(n14768), .A(n9204), .ZN(n9205) );
  OAI21_X1 U11703 ( .B1(n9448), .B2(n14352), .A(n9205), .ZN(n9209) );
  NAND2_X1 U11704 ( .A1(n9209), .A2(n6470), .ZN(n9206) );
  OAI21_X1 U11705 ( .B1(n6470), .B2(n9207), .A(n9206), .ZN(P2_U3505) );
  INV_X2 U11706 ( .A(n14795), .ZN(n14797) );
  INV_X1 U11707 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n9211) );
  NAND2_X1 U11708 ( .A1(n9209), .A2(n14797), .ZN(n9210) );
  OAI21_X1 U11709 ( .B1(n14797), .B2(n9211), .A(n9210), .ZN(P2_U3448) );
  NAND2_X1 U11710 ( .A1(n9354), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9213) );
  XNOR2_X1 U11711 ( .A(n9213), .B(P2_IR_REG_14__SCAN_IN), .ZN(n10725) );
  INV_X1 U11712 ( .A(n10725), .ZN(n10479) );
  OAI222_X1 U11713 ( .A1(n13440), .A2(n9215), .B1(n13438), .B2(n9214), .C1(
        n10479), .C2(P2_U3088), .ZN(P2_U3313) );
  OAI21_X1 U11714 ( .B1(n9217), .B2(n14813), .A(n9216), .ZN(n9229) );
  AOI21_X1 U11715 ( .B1(n15022), .B2(n9219), .A(n9218), .ZN(n9225) );
  AOI21_X1 U11716 ( .B1(n14976), .B2(n9221), .A(n9220), .ZN(n9222) );
  OR2_X1 U11717 ( .A1(n14893), .A2(n9222), .ZN(n9224) );
  AOI22_X1 U11718 ( .A1(n14869), .A2(P3_ADDR_REG_1__SCAN_IN), .B1(
        P3_REG3_REG_1__SCAN_IN), .B2(P3_U3151), .ZN(n9223) );
  OAI211_X1 U11719 ( .C1(n9225), .C2(n14887), .A(n9224), .B(n9223), .ZN(n9228)
         );
  NOR2_X1 U11720 ( .A1(n14878), .A2(n9226), .ZN(n9227) );
  AOI211_X1 U11721 ( .C1(n14843), .C2(n9229), .A(n9228), .B(n9227), .ZN(n9230)
         );
  INV_X1 U11722 ( .A(n9230), .ZN(P3_U3183) );
  NAND2_X1 U11723 ( .A1(n9236), .A2(n15089), .ZN(n9231) );
  MUX2_X1 U11724 ( .A(n7296), .B(n9358), .S(n11543), .Z(n9233) );
  INV_X1 U11725 ( .A(n9233), .ZN(n9234) );
  NAND2_X1 U11726 ( .A1(n9234), .A2(SI_15_), .ZN(n9235) );
  NAND2_X1 U11727 ( .A1(n9238), .A2(n9235), .ZN(n9350) );
  NOR2_X1 U11728 ( .A1(n9236), .A2(n15089), .ZN(n9237) );
  NAND2_X1 U11729 ( .A1(n9239), .A2(n9238), .ZN(n9363) );
  MUX2_X1 U11730 ( .A(n9251), .B(n9246), .S(n11543), .Z(n9240) );
  INV_X1 U11731 ( .A(n9240), .ZN(n9241) );
  NAND2_X1 U11732 ( .A1(n9241), .A2(SI_16_), .ZN(n9242) );
  XNOR2_X1 U11733 ( .A(n9363), .B(n9362), .ZN(n11088) );
  INV_X1 U11734 ( .A(n11088), .ZN(n9250) );
  INV_X1 U11735 ( .A(n9243), .ZN(n9244) );
  NAND2_X1 U11736 ( .A1(n9244), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9245) );
  XNOR2_X1 U11737 ( .A(n9245), .B(P2_IR_REG_16__SCAN_IN), .ZN(n10928) );
  INV_X1 U11738 ( .A(n10928), .ZN(n10822) );
  OAI222_X1 U11739 ( .A1(n13440), .A2(n9246), .B1(n13438), .B2(n9250), .C1(
        n10822), .C2(P2_U3088), .ZN(P2_U3311) );
  INV_X1 U11740 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n9248) );
  NAND2_X1 U11741 ( .A1(n9247), .A2(n9248), .ZN(n9367) );
  NAND2_X1 U11742 ( .A1(n9367), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9249) );
  XNOR2_X1 U11743 ( .A(n9249), .B(P1_IR_REG_16__SCAN_IN), .ZN(n11089) );
  OAI222_X1 U11744 ( .A1(n14124), .A2(n9251), .B1(n14130), .B2(n9250), .C1(
        n10714), .C2(P1_U3086), .ZN(P1_U3339) );
  OR2_X1 U11745 ( .A1(n9253), .A2(n9252), .ZN(n9254) );
  INV_X1 U11746 ( .A(n9937), .ZN(n9268) );
  INV_X1 U11747 ( .A(n9663), .ZN(n9267) );
  NOR4_X1 U11748 ( .A1(P1_D_REG_18__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_20__SCAN_IN), .A4(P1_D_REG_21__SCAN_IN), .ZN(n9259) );
  NOR4_X1 U11749 ( .A1(P1_D_REG_16__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_15__SCAN_IN), .A4(P1_D_REG_17__SCAN_IN), .ZN(n9258) );
  NOR4_X1 U11750 ( .A1(P1_D_REG_26__SCAN_IN), .A2(P1_D_REG_27__SCAN_IN), .A3(
        P1_D_REG_28__SCAN_IN), .A4(P1_D_REG_31__SCAN_IN), .ZN(n9257) );
  NOR4_X1 U11751 ( .A1(P1_D_REG_22__SCAN_IN), .A2(P1_D_REG_23__SCAN_IN), .A3(
        P1_D_REG_24__SCAN_IN), .A4(P1_D_REG_25__SCAN_IN), .ZN(n9256) );
  NAND4_X1 U11752 ( .A1(n9259), .A2(n9258), .A3(n9257), .A4(n9256), .ZN(n9265)
         );
  NOR2_X1 U11753 ( .A1(P1_D_REG_2__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .ZN(
        n9263) );
  NOR4_X1 U11754 ( .A1(P1_D_REG_29__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_4__SCAN_IN), .A4(P1_D_REG_5__SCAN_IN), .ZN(n9262) );
  NOR4_X1 U11755 ( .A1(P1_D_REG_10__SCAN_IN), .A2(P1_D_REG_11__SCAN_IN), .A3(
        P1_D_REG_12__SCAN_IN), .A4(P1_D_REG_13__SCAN_IN), .ZN(n9261) );
  NOR4_X1 U11756 ( .A1(P1_D_REG_6__SCAN_IN), .A2(P1_D_REG_7__SCAN_IN), .A3(
        P1_D_REG_8__SCAN_IN), .A4(P1_D_REG_9__SCAN_IN), .ZN(n9260) );
  NAND4_X1 U11757 ( .A1(n9263), .A2(n9262), .A3(n9261), .A4(n9260), .ZN(n9264)
         );
  NOR2_X1 U11758 ( .A1(n9265), .A2(n9264), .ZN(n9662) );
  NAND2_X1 U11759 ( .A1(n9662), .A2(P1_D_REG_0__SCAN_IN), .ZN(n9266) );
  AOI21_X1 U11760 ( .B1(n9267), .B2(n9266), .A(n9660), .ZN(n9686) );
  NAND2_X1 U11761 ( .A1(n9268), .A2(n9686), .ZN(n9302) );
  NAND2_X1 U11762 ( .A1(n11199), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9270) );
  NAND2_X1 U11763 ( .A1(n9274), .A2(n11199), .ZN(n13806) );
  NAND2_X1 U11764 ( .A1(n11206), .A2(n13806), .ZN(n9296) );
  AND2_X1 U11765 ( .A1(n9275), .A2(n9296), .ZN(n9300) );
  INV_X1 U11766 ( .A(n14544), .ZN(n9276) );
  NAND2_X1 U11767 ( .A1(n9276), .A2(n11206), .ZN(n9666) );
  NOR2_X1 U11768 ( .A1(n14596), .A2(n13806), .ZN(n9658) );
  INV_X1 U11769 ( .A(n9658), .ZN(n9282) );
  OAI21_X1 U11770 ( .B1(n9302), .B2(n9300), .A(n9282), .ZN(n9279) );
  AND2_X1 U11771 ( .A1(n9284), .A2(n9277), .ZN(n9278) );
  NAND2_X1 U11772 ( .A1(n9279), .A2(n9278), .ZN(n9632) );
  OR2_X1 U11773 ( .A1(n9632), .A2(P1_U3086), .ZN(n9655) );
  INV_X1 U11774 ( .A(n9655), .ZN(n9309) );
  INV_X1 U11775 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n9981) );
  NOR2_X1 U11776 ( .A1(n11543), .A2(n9280), .ZN(n9281) );
  XNOR2_X1 U11777 ( .A(n9281), .B(P2_DATAO_REG_0__SCAN_IN), .ZN(n14133) );
  MUX2_X1 U11778 ( .A(n13671), .B(n14133), .S(n11364), .Z(n14546) );
  INV_X1 U11779 ( .A(n14546), .ZN(n9668) );
  NOR2_X1 U11780 ( .A1(n9302), .A2(n9301), .ZN(n9295) );
  NAND2_X1 U11781 ( .A1(n7146), .A2(n7147), .ZN(n11605) );
  NOR2_X1 U11782 ( .A1(n14544), .A2(n11605), .ZN(n9944) );
  NAND2_X1 U11783 ( .A1(n9295), .A2(n9944), .ZN(n9283) );
  OR2_X2 U11784 ( .A1(n9301), .A2(n9282), .ZN(n14532) );
  NAND2_X2 U11785 ( .A1(n9284), .A2(n9940), .ZN(n13535) );
  INV_X1 U11786 ( .A(n9284), .ZN(n9285) );
  NAND2_X1 U11787 ( .A1(n11502), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n9291) );
  OR2_X1 U11788 ( .A1(n6476), .A2(n9981), .ZN(n9290) );
  INV_X1 U11789 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n9286) );
  OR2_X1 U11790 ( .A1(n9853), .A2(n9286), .ZN(n9289) );
  INV_X1 U11791 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n9287) );
  OR2_X1 U11792 ( .A1(n9593), .A2(n9287), .ZN(n9288) );
  NAND4_X2 U11793 ( .A1(n9291), .A2(n9290), .A3(n9289), .A4(n9288), .ZN(n14526) );
  NAND2_X1 U11794 ( .A1(n14526), .A2(n9619), .ZN(n9292) );
  AOI21_X1 U11795 ( .B1(n9575), .B2(n9294), .A(n9574), .ZN(n13678) );
  INV_X1 U11796 ( .A(n9295), .ZN(n9299) );
  NAND2_X1 U11797 ( .A1(n7146), .A2(n9296), .ZN(n9297) );
  NAND2_X1 U11798 ( .A1(n14606), .A2(n11538), .ZN(n9298) );
  OR2_X1 U11799 ( .A1(n9302), .A2(n11613), .ZN(n13513) );
  NOR2_X2 U11800 ( .A1(n13513), .A2(n14008), .ZN(n13639) );
  INV_X1 U11801 ( .A(P1_REG3_REG_1__SCAN_IN), .ZN(n14533) );
  OAI22_X1 U11802 ( .A1(n13678), .A2(n13650), .B1(n13617), .B2(n6669), .ZN(
        n9307) );
  AOI21_X1 U11803 ( .B1(n9668), .B2(n13647), .A(n9307), .ZN(n9308) );
  OAI21_X1 U11804 ( .B1(n9309), .B2(n9981), .A(n9308), .ZN(P1_U3232) );
  NAND3_X1 U11805 ( .A1(n9312), .A2(n9311), .A3(n9310), .ZN(n9317) );
  OR2_X1 U11806 ( .A1(n9317), .A2(n14738), .ZN(n9323) );
  INV_X1 U11807 ( .A(n12703), .ZN(n12719) );
  NOR2_X2 U11808 ( .A1(n9323), .A2(n9314), .ZN(n14330) );
  INV_X1 U11809 ( .A(n9315), .ZN(n9316) );
  NAND2_X1 U11810 ( .A1(n9317), .A2(n9316), .ZN(n9321) );
  AND3_X1 U11811 ( .A1(n9319), .A2(n9318), .A3(n13027), .ZN(n9320) );
  NAND2_X1 U11812 ( .A1(n9321), .A2(n9320), .ZN(n9451) );
  OR2_X1 U11813 ( .A1(n9451), .A2(P2_U3088), .ZN(n11982) );
  AOI22_X1 U11814 ( .A1(n14330), .A2(n9322), .B1(n11982), .B2(
        P2_REG3_REG_2__SCAN_IN), .ZN(n9346) );
  INV_X1 U11815 ( .A(n9323), .ZN(n9326) );
  NOR2_X1 U11816 ( .A1(n14788), .A2(n9324), .ZN(n9325) );
  XNOR2_X1 U11817 ( .A(n12740), .B(n11628), .ZN(n9333) );
  INV_X1 U11818 ( .A(n9333), .ZN(n9331) );
  NOR2_X2 U11819 ( .A1(n9329), .A2(n12988), .ZN(n9335) );
  NAND2_X1 U11820 ( .A1(n13066), .A2(n11749), .ZN(n9332) );
  INV_X1 U11821 ( .A(n9332), .ZN(n9330) );
  NAND2_X1 U11822 ( .A1(n9331), .A2(n9330), .ZN(n9334) );
  NAND2_X1 U11823 ( .A1(n9333), .A2(n9332), .ZN(n9449) );
  AND2_X1 U11824 ( .A1(n9334), .A2(n9449), .ZN(n9343) );
  XNOR2_X1 U11825 ( .A(n9339), .B(n9338), .ZN(n11986) );
  NAND2_X1 U11826 ( .A1(n9335), .A2(n14743), .ZN(n9434) );
  AND2_X1 U11827 ( .A1(n9438), .A2(n9434), .ZN(n9488) );
  NAND2_X1 U11828 ( .A1(n9441), .A2(n11750), .ZN(n9337) );
  NAND2_X1 U11829 ( .A1(n9488), .A2(n9337), .ZN(n11985) );
  INV_X1 U11830 ( .A(n9338), .ZN(n9340) );
  NAND2_X1 U11831 ( .A1(n9340), .A2(n9339), .ZN(n9341) );
  NAND2_X1 U11832 ( .A1(n11984), .A2(n9341), .ZN(n9342) );
  NAND2_X1 U11833 ( .A1(n9342), .A2(n9343), .ZN(n9450) );
  OAI21_X1 U11834 ( .B1(n9343), .B2(n9342), .A(n9450), .ZN(n9344) );
  NAND2_X1 U11835 ( .A1(n14328), .A2(n9344), .ZN(n9345) );
  OAI211_X1 U11836 ( .C1(n12719), .C2(n9024), .A(n9346), .B(n9345), .ZN(
        P2_U3209) );
  OAI21_X1 U11837 ( .B1(n9349), .B2(n9348), .A(n9347), .ZN(n9352) );
  INV_X1 U11838 ( .A(n9350), .ZN(n9351) );
  XNOR2_X1 U11839 ( .A(n9352), .B(n9351), .ZN(n10976) );
  INV_X1 U11840 ( .A(n10976), .ZN(n9357) );
  OR2_X1 U11841 ( .A1(n9247), .A2(n14111), .ZN(n9353) );
  XNOR2_X1 U11842 ( .A(n9353), .B(P1_IR_REG_15__SCAN_IN), .ZN(n10977) );
  INV_X1 U11843 ( .A(n10977), .ZN(n10090) );
  OAI222_X1 U11844 ( .A1(n14124), .A2(n7296), .B1(n14119), .B2(n9357), .C1(
        n10090), .C2(P1_U3086), .ZN(P1_U3340) );
  OAI21_X1 U11845 ( .B1(n9354), .B2(P2_IR_REG_14__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n9355) );
  XNOR2_X1 U11846 ( .A(n9355), .B(P2_IR_REG_15__SCAN_IN), .ZN(n10730) );
  INV_X1 U11847 ( .A(n10730), .ZN(n9356) );
  OAI222_X1 U11848 ( .A1(n13440), .A2(n9358), .B1(n13438), .B2(n9357), .C1(
        n9356), .C2(P2_U3088), .ZN(P2_U3312) );
  INV_X1 U11849 ( .A(n9359), .ZN(n9361) );
  OAI222_X1 U11850 ( .A1(n12607), .A2(n9361), .B1(n9360), .B2(P3_U3151), .C1(
        n15045), .C2(n12608), .ZN(P3_U3276) );
  NAND2_X1 U11851 ( .A1(n9363), .A2(n9362), .ZN(n9365) );
  NAND2_X1 U11852 ( .A1(n9365), .A2(n9364), .ZN(n9817) );
  MUX2_X1 U11853 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(P1_DATAO_REG_17__SCAN_IN), 
        .S(n11543), .Z(n9815) );
  XNOR2_X1 U11854 ( .A(n9815), .B(n15072), .ZN(n9366) );
  XNOR2_X1 U11855 ( .A(n9817), .B(n9366), .ZN(n11305) );
  INV_X1 U11856 ( .A(n11305), .ZN(n9373) );
  OR2_X1 U11857 ( .A1(n9367), .A2(P1_IR_REG_16__SCAN_IN), .ZN(n9822) );
  NAND2_X1 U11858 ( .A1(n9822), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n9369) );
  INV_X1 U11859 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n9368) );
  XNOR2_X1 U11860 ( .A(n9369), .B(n9368), .ZN(n10953) );
  OAI222_X1 U11861 ( .A1(n14124), .A2(n9370), .B1(n14119), .B2(n9373), .C1(
        n10953), .C2(P1_U3086), .ZN(P1_U3338) );
  INV_X1 U11862 ( .A(n9371), .ZN(n9826) );
  NAND2_X1 U11863 ( .A1(n9371), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9372) );
  XNOR2_X1 U11864 ( .A(n9372), .B(P2_IR_REG_17__SCAN_IN), .ZN(n11027) );
  INV_X1 U11865 ( .A(n11027), .ZN(n13136) );
  OAI222_X1 U11866 ( .A1(n13440), .A2(n9374), .B1(n13438), .B2(n9373), .C1(
        n13136), .C2(P2_U3088), .ZN(P2_U3310) );
  NAND2_X1 U11867 ( .A1(n12143), .A2(P3_DATAO_REG_29__SCAN_IN), .ZN(n9375) );
  OAI21_X1 U11868 ( .B1(n9376), .B2(n12143), .A(n9375), .ZN(P3_U3520) );
  NAND2_X1 U11869 ( .A1(n14727), .A2(n9377), .ZN(n9383) );
  INV_X1 U11870 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n13068) );
  OAI22_X1 U11871 ( .A1(n13282), .A2(n9379), .B1(n13068), .B2(n14706), .ZN(
        n9381) );
  NOR2_X1 U11872 ( .A1(n14721), .A2(n9021), .ZN(n9380) );
  AOI211_X1 U11873 ( .C1(n14731), .C2(P2_REG2_REG_1__SCAN_IN), .A(n9381), .B(
        n9380), .ZN(n9382) );
  OAI211_X1 U11874 ( .C1(n14731), .C2(n9384), .A(n9383), .B(n9382), .ZN(
        P2_U3264) );
  AOI21_X1 U11875 ( .B1(n9387), .B2(n9386), .A(n9385), .ZN(n9401) );
  OAI21_X1 U11876 ( .B1(n9390), .B2(n9389), .A(n9388), .ZN(n9396) );
  AOI21_X1 U11877 ( .B1(n9393), .B2(n9392), .A(n9391), .ZN(n9394) );
  NOR2_X1 U11878 ( .A1(n9394), .A2(n14893), .ZN(n9395) );
  AOI21_X1 U11879 ( .B1(n14843), .B2(n9396), .A(n9395), .ZN(n9400) );
  NAND2_X1 U11880 ( .A1(P3_U3151), .A2(P3_REG3_REG_5__SCAN_IN), .ZN(n10034) );
  OAI21_X1 U11881 ( .B1(n14875), .B2(n6688), .A(n10034), .ZN(n9397) );
  AOI21_X1 U11882 ( .B1(n9398), .B2(n14846), .A(n9397), .ZN(n9399) );
  OAI211_X1 U11883 ( .C1(n9401), .C2(n14887), .A(n9400), .B(n9399), .ZN(
        P3_U3187) );
  INV_X1 U11884 ( .A(n13062), .ZN(n9403) );
  NAND2_X1 U11885 ( .A1(n12776), .A2(n9403), .ZN(n9404) );
  OR2_X1 U11886 ( .A1(n10172), .A2(n12931), .ZN(n9406) );
  AOI22_X1 U11887 ( .A1(n9097), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n9142), .B2(
        n13105), .ZN(n9405) );
  NAND2_X1 U11888 ( .A1(n9406), .A2(n9405), .ZN(n12791) );
  INV_X1 U11889 ( .A(n13061), .ZN(n9773) );
  XNOR2_X1 U11890 ( .A(n9769), .B(n13001), .ZN(n9433) );
  NAND2_X1 U11891 ( .A1(n13062), .A2(n12710), .ZN(n9412) );
  NAND2_X1 U11892 ( .A1(n11701), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n9410) );
  NAND2_X1 U11893 ( .A1(n11123), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n9409) );
  XNOR2_X1 U11894 ( .A(n9744), .B(P2_REG3_REG_8__SCAN_IN), .ZN(n9741) );
  NAND2_X1 U11895 ( .A1(n9145), .A2(n9741), .ZN(n9408) );
  NAND2_X1 U11896 ( .A1(n11688), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n9407) );
  NAND4_X1 U11897 ( .A1(n9410), .A2(n9409), .A3(n9408), .A4(n9407), .ZN(n13060) );
  NAND2_X1 U11898 ( .A1(n13060), .A2(n12711), .ZN(n9411) );
  NAND2_X1 U11899 ( .A1(n9412), .A2(n9411), .ZN(n9482) );
  INV_X1 U11900 ( .A(n9780), .ZN(n9413) );
  AOI211_X1 U11901 ( .C1(n12791), .C2(n9414), .A(n9329), .B(n9413), .ZN(n9424)
         );
  AOI211_X1 U11902 ( .C1(n12791), .C2(n14788), .A(n9482), .B(n9424), .ZN(n9419) );
  NAND2_X1 U11903 ( .A1(n12776), .A2(n13062), .ZN(n9417) );
  XOR2_X1 U11904 ( .A(n9765), .B(n13001), .Z(n9431) );
  NAND2_X1 U11905 ( .A1(n9431), .A2(n14768), .ZN(n9418) );
  OAI211_X1 U11906 ( .C1(n14352), .C2(n9433), .A(n9419), .B(n9418), .ZN(n9421)
         );
  NAND2_X1 U11907 ( .A1(n9421), .A2(n6470), .ZN(n9420) );
  OAI21_X1 U11908 ( .B1(n6470), .B2(n8866), .A(n9420), .ZN(P2_U3506) );
  INV_X1 U11909 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n9423) );
  NAND2_X1 U11910 ( .A1(n9421), .A2(n14797), .ZN(n9422) );
  OAI21_X1 U11911 ( .B1(n14797), .B2(n9423), .A(n9422), .ZN(P2_U3451) );
  OR2_X1 U11912 ( .A1(n14731), .A2(n14352), .ZN(n13198) );
  INV_X1 U11913 ( .A(n12791), .ZN(n9429) );
  NAND2_X1 U11914 ( .A1(n9424), .A2(n14725), .ZN(n9428) );
  INV_X1 U11915 ( .A(n14706), .ZN(n14719) );
  MUX2_X1 U11916 ( .A(n9482), .B(P2_REG2_REG_7__SCAN_IN), .S(n14731), .Z(n9425) );
  AOI21_X1 U11917 ( .B1(n14719), .B2(n9426), .A(n9425), .ZN(n9427) );
  OAI211_X1 U11918 ( .C1(n9429), .C2(n14721), .A(n9428), .B(n9427), .ZN(n9430)
         );
  AOI21_X1 U11919 ( .B1(n14727), .B2(n9431), .A(n9430), .ZN(n9432) );
  OAI21_X1 U11920 ( .B1(n9433), .B2(n13198), .A(n9432), .ZN(P2_U3258) );
  INV_X1 U11921 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n14635) );
  NAND2_X1 U11922 ( .A1(n13067), .A2(n12711), .ZN(n14745) );
  OAI211_X1 U11923 ( .C1(n14706), .C2(n14635), .A(n9434), .B(n14745), .ZN(
        n9436) );
  NOR2_X1 U11924 ( .A1(n13316), .A2(n14631), .ZN(n9435) );
  AOI21_X1 U11925 ( .B1(n13316), .B2(n9436), .A(n9435), .ZN(n9440) );
  INV_X1 U11926 ( .A(n13198), .ZN(n13284) );
  NAND2_X1 U11927 ( .A1(n9438), .A2(n12731), .ZN(n14748) );
  OAI21_X1 U11928 ( .B1(n14727), .B2(n13284), .A(n14748), .ZN(n9439) );
  OAI211_X1 U11929 ( .C1(n14721), .C2(n9441), .A(n9440), .B(n9439), .ZN(
        P2_U3265) );
  AOI22_X1 U11930 ( .A1(n14341), .A2(n12776), .B1(n9712), .B2(n14719), .ZN(
        n9443) );
  MUX2_X1 U11931 ( .A(n9710), .B(n8874), .S(n14731), .Z(n9442) );
  OAI211_X1 U11932 ( .C1(n9444), .C2(n13282), .A(n9443), .B(n9442), .ZN(n9445)
         );
  AOI21_X1 U11933 ( .B1(n9446), .B2(n14727), .A(n9445), .ZN(n9447) );
  OAI21_X1 U11934 ( .B1(n9448), .B2(n13198), .A(n9447), .ZN(P2_U3259) );
  NAND2_X1 U11935 ( .A1(n9450), .A2(n9449), .ZN(n9458) );
  XNOR2_X1 U11936 ( .A(n12759), .B(n11628), .ZN(n9460) );
  NAND2_X1 U11937 ( .A1(n13065), .A2(n11749), .ZN(n9461) );
  XNOR2_X1 U11938 ( .A(n9460), .B(n9461), .ZN(n9459) );
  XNOR2_X1 U11939 ( .A(n9458), .B(n9459), .ZN(n9457) );
  INV_X1 U11940 ( .A(n14334), .ZN(n12717) );
  NAND2_X1 U11941 ( .A1(n14330), .A2(n9452), .ZN(n9454) );
  OAI211_X1 U11942 ( .C1(n12719), .C2(n14755), .A(n9454), .B(n9453), .ZN(n9455) );
  AOI21_X1 U11943 ( .B1(n12717), .B2(n9029), .A(n9455), .ZN(n9456) );
  OAI21_X1 U11944 ( .B1(n9457), .B2(n12705), .A(n9456), .ZN(P2_U3190) );
  INV_X1 U11945 ( .A(n9460), .ZN(n9463) );
  INV_X1 U11946 ( .A(n9461), .ZN(n9462) );
  XNOR2_X1 U11947 ( .A(n12754), .B(n11628), .ZN(n9465) );
  NAND2_X1 U11948 ( .A1(n13064), .A2(n11749), .ZN(n9466) );
  NAND2_X1 U11949 ( .A1(n9465), .A2(n9466), .ZN(n9470) );
  INV_X1 U11950 ( .A(n9465), .ZN(n9468) );
  INV_X1 U11951 ( .A(n9466), .ZN(n9467) );
  NAND2_X1 U11952 ( .A1(n9468), .A2(n9467), .ZN(n9469) );
  AND2_X1 U11953 ( .A1(n9470), .A2(n9469), .ZN(n9693) );
  XNOR2_X1 U11954 ( .A(n12773), .B(n11628), .ZN(n9471) );
  NAND2_X1 U11955 ( .A1(n13063), .A2(n11749), .ZN(n9472) );
  NAND2_X1 U11956 ( .A1(n9471), .A2(n9472), .ZN(n9476) );
  INV_X1 U11957 ( .A(n9471), .ZN(n9474) );
  INV_X1 U11958 ( .A(n9472), .ZN(n9473) );
  NAND2_X1 U11959 ( .A1(n9474), .A2(n9473), .ZN(n9475) );
  AND2_X1 U11960 ( .A1(n9476), .A2(n9475), .ZN(n9700) );
  NAND2_X1 U11961 ( .A1(n9699), .A2(n9700), .ZN(n9698) );
  XNOR2_X1 U11962 ( .A(n12776), .B(n11628), .ZN(n9477) );
  NAND2_X1 U11963 ( .A1(n13062), .A2(n11749), .ZN(n9478) );
  XNOR2_X1 U11964 ( .A(n9477), .B(n9478), .ZN(n9707) );
  INV_X1 U11965 ( .A(n9477), .ZN(n9480) );
  INV_X1 U11966 ( .A(n9478), .ZN(n9479) );
  NAND2_X1 U11967 ( .A1(n9480), .A2(n9479), .ZN(n9481) );
  XNOR2_X1 U11968 ( .A(n12791), .B(n11750), .ZN(n9730) );
  NAND2_X1 U11969 ( .A1(n13061), .A2(n11749), .ZN(n9728) );
  XNOR2_X1 U11970 ( .A(n9730), .B(n9728), .ZN(n9726) );
  XNOR2_X1 U11971 ( .A(n9727), .B(n9726), .ZN(n9487) );
  NAND2_X1 U11972 ( .A1(n14330), .A2(n9482), .ZN(n9483) );
  NAND2_X1 U11973 ( .A1(P2_U3088), .A2(P2_REG3_REG_7__SCAN_IN), .ZN(n13102) );
  OAI211_X1 U11974 ( .C1(n14334), .C2(n9484), .A(n9483), .B(n13102), .ZN(n9485) );
  AOI21_X1 U11975 ( .B1(n12791), .B2(n12703), .A(n9485), .ZN(n9486) );
  OAI21_X1 U11976 ( .B1(n9487), .B2(n12705), .A(n9486), .ZN(P2_U3185) );
  INV_X1 U11977 ( .A(n14330), .ZN(n12715) );
  AOI22_X1 U11978 ( .A1(n14331), .A2(n14743), .B1(n11982), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n9491) );
  OAI21_X1 U11979 ( .B1(n9335), .B2(n12731), .A(n9488), .ZN(n9489) );
  NAND2_X1 U11980 ( .A1(n14328), .A2(n9489), .ZN(n9490) );
  OAI211_X1 U11981 ( .C1(n12715), .C2(n14745), .A(n9491), .B(n9490), .ZN(
        P2_U3204) );
  NAND2_X1 U11982 ( .A1(n9502), .A2(n14298), .ZN(n9492) );
  NAND2_X1 U11983 ( .A1(n12142), .A2(n12437), .ZN(n9512) );
  OAI21_X1 U11984 ( .B1(n9519), .B2(n9492), .A(n9512), .ZN(n10110) );
  INV_X1 U11985 ( .A(n10110), .ZN(n9494) );
  AOI22_X1 U11986 ( .A1(n10361), .A2(n9522), .B1(n15036), .B2(
        P3_REG1_REG_0__SCAN_IN), .ZN(n9493) );
  OAI21_X1 U11987 ( .B1(n9494), .B2(n15036), .A(n9493), .ZN(P3_U3459) );
  NAND2_X1 U11988 ( .A1(n9517), .A2(n9513), .ZN(n9500) );
  NOR2_X1 U11989 ( .A1(n9496), .A2(n9495), .ZN(n9499) );
  INV_X1 U11990 ( .A(n9515), .ZN(n9497) );
  NAND2_X1 U11991 ( .A1(n9514), .A2(n9497), .ZN(n9498) );
  NAND4_X1 U11992 ( .A1(n9500), .A2(n9499), .A3(n9886), .A4(n9498), .ZN(n9501)
         );
  NAND2_X1 U11993 ( .A1(n9501), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9505) );
  NOR2_X1 U11994 ( .A1(n9509), .A2(n9502), .ZN(n9503) );
  NAND2_X1 U11995 ( .A1(n9514), .A2(n9503), .ZN(n9504) );
  NOR2_X1 U11996 ( .A1(n12112), .A2(P3_U3151), .ZN(n9725) );
  INV_X1 U11997 ( .A(P3_REG3_REG_0__SCAN_IN), .ZN(n9524) );
  NAND2_X1 U11998 ( .A1(n9517), .A2(n14969), .ZN(n9507) );
  NOR2_X1 U11999 ( .A1(n9509), .A2(n14298), .ZN(n9506) );
  INV_X1 U12000 ( .A(n9514), .ZN(n9511) );
  NOR2_X1 U12001 ( .A1(n9509), .A2(n9508), .ZN(n9510) );
  NOR2_X1 U12002 ( .A1(n9512), .A2(n14281), .ZN(n9521) );
  NAND2_X1 U12003 ( .A1(n9513), .A2(n14298), .ZN(n9516) );
  OAI22_X1 U12004 ( .A1(n9517), .A2(n9516), .B1(n9515), .B2(n9514), .ZN(n9518)
         );
  NOR2_X1 U12005 ( .A1(n9519), .A2(n12115), .ZN(n9520) );
  AOI211_X1 U12006 ( .C1(n14274), .C2(n9522), .A(n9521), .B(n9520), .ZN(n9523)
         );
  OAI21_X1 U12007 ( .B1(n9725), .B2(n9524), .A(n9523), .ZN(P3_U3172) );
  INV_X1 U12008 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n14440) );
  INV_X1 U12009 ( .A(n14491), .ZN(n9527) );
  AOI21_X1 U12010 ( .B1(n10457), .B2(P1_REG1_REG_10__SCAN_IN), .A(n9525), .ZN(
        n13778) );
  INV_X1 U12011 ( .A(P1_REG1_REG_11__SCAN_IN), .ZN(n14446) );
  MUX2_X1 U12012 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n14446), .S(n13783), .Z(
        n13779) );
  NAND2_X1 U12013 ( .A1(n13778), .A2(n13779), .ZN(n14483) );
  NAND2_X1 U12014 ( .A1(n9526), .A2(n14446), .ZN(n14481) );
  INV_X1 U12015 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n10608) );
  MUX2_X1 U12016 ( .A(n10608), .B(P1_REG1_REG_12__SCAN_IN), .S(n14491), .Z(
        n14482) );
  AOI21_X1 U12017 ( .B1(n14483), .B2(n14481), .A(n14482), .ZN(n14480) );
  AOI21_X1 U12018 ( .B1(n10608), .B2(n9527), .A(n14480), .ZN(n14506) );
  MUX2_X1 U12019 ( .A(P1_REG1_REG_13__SCAN_IN), .B(n14440), .S(n10766), .Z(
        n14505) );
  NAND2_X1 U12020 ( .A1(n14506), .A2(n14505), .ZN(n14503) );
  OAI21_X1 U12021 ( .B1(n14500), .B2(n14440), .A(n14503), .ZN(n9529) );
  INV_X1 U12022 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n10773) );
  MUX2_X1 U12023 ( .A(n10773), .B(P1_REG1_REG_14__SCAN_IN), .S(n10971), .Z(
        n9528) );
  NOR2_X1 U12024 ( .A1(n9528), .A2(n9529), .ZN(n10084) );
  AOI21_X1 U12025 ( .B1(n9529), .B2(n9528), .A(n10084), .ZN(n9545) );
  NAND2_X1 U12026 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n10766), .ZN(n9538) );
  INV_X1 U12027 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n9530) );
  MUX2_X1 U12028 ( .A(n9530), .B(P1_REG2_REG_13__SCAN_IN), .S(n10766), .Z(
        n9531) );
  INV_X1 U12029 ( .A(n9531), .ZN(n14509) );
  NAND2_X1 U12030 ( .A1(n10457), .A2(P1_REG2_REG_10__SCAN_IN), .ZN(n13785) );
  NAND2_X1 U12031 ( .A1(n13786), .A2(n13785), .ZN(n9533) );
  INV_X1 U12032 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n10625) );
  MUX2_X1 U12033 ( .A(P1_REG2_REG_11__SCAN_IN), .B(n10625), .S(n13783), .Z(
        n9532) );
  NAND2_X1 U12034 ( .A1(n9533), .A2(n9532), .ZN(n13788) );
  NAND2_X1 U12035 ( .A1(n13783), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n9534) );
  AND2_X1 U12036 ( .A1(n13788), .A2(n9534), .ZN(n14487) );
  INV_X1 U12037 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n9535) );
  MUX2_X1 U12038 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n9535), .S(n14491), .Z(
        n14488) );
  NAND2_X1 U12039 ( .A1(n14487), .A2(n14488), .ZN(n14486) );
  INV_X1 U12040 ( .A(n14486), .ZN(n9537) );
  NOR2_X1 U12041 ( .A1(n14491), .A2(P1_REG2_REG_12__SCAN_IN), .ZN(n9536) );
  NOR2_X1 U12042 ( .A1(n9537), .A2(n9536), .ZN(n14510) );
  NAND2_X1 U12043 ( .A1(n14509), .A2(n14510), .ZN(n14507) );
  NAND2_X1 U12044 ( .A1(n9538), .A2(n14507), .ZN(n9541) );
  INV_X1 U12045 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n9539) );
  MUX2_X1 U12046 ( .A(P1_REG2_REG_14__SCAN_IN), .B(n9539), .S(n10971), .Z(
        n9540) );
  NAND2_X1 U12047 ( .A1(n9541), .A2(n9540), .ZN(n10082) );
  OAI211_X1 U12048 ( .C1(n9541), .C2(n9540), .A(n10082), .B(n14508), .ZN(n9544) );
  INV_X1 U12049 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n14225) );
  NAND2_X1 U12050 ( .A1(P1_REG3_REG_14__SCAN_IN), .A2(P1_U3086), .ZN(n13503)
         );
  OAI21_X1 U12051 ( .B1(n14495), .B2(n14225), .A(n13503), .ZN(n9542) );
  AOI21_X1 U12052 ( .B1(n10971), .B2(n14490), .A(n9542), .ZN(n9543) );
  OAI211_X1 U12053 ( .C1(n9545), .C2(n13801), .A(n9544), .B(n9543), .ZN(
        P1_U3257) );
  INV_X1 U12054 ( .A(P3_REG3_REG_1__SCAN_IN), .ZN(n9562) );
  AOI21_X1 U12055 ( .B1(n10112), .B2(n9758), .A(n9547), .ZN(n9548) );
  NAND3_X1 U12056 ( .A1(n12142), .A2(n6508), .A3(n9552), .ZN(n9553) );
  NAND2_X1 U12057 ( .A1(n14960), .A2(n6508), .ZN(n9554) );
  NAND2_X1 U12058 ( .A1(n9555), .A2(n9554), .ZN(n9556) );
  NAND2_X1 U12059 ( .A1(n6539), .A2(n9556), .ZN(n9717) );
  NAND3_X1 U12060 ( .A1(n14966), .A2(n14967), .A3(n11971), .ZN(n9557) );
  OAI211_X1 U12061 ( .C1(n6539), .C2(n14960), .A(n9717), .B(n9557), .ZN(n9558)
         );
  NAND2_X1 U12062 ( .A1(n9558), .A2(n14276), .ZN(n9561) );
  NAND2_X1 U12063 ( .A1(n12144), .A2(n12440), .ZN(n9559) );
  OAI21_X1 U12064 ( .B1(n9992), .B2(n12100), .A(n9559), .ZN(n14963) );
  AOI22_X1 U12065 ( .A1(n14963), .A2(n12104), .B1(n14274), .B2(n9552), .ZN(
        n9560) );
  OAI211_X1 U12066 ( .C1(n9725), .C2(n9562), .A(n9561), .B(n9560), .ZN(
        P3_U3162) );
  NAND2_X1 U12067 ( .A1(n11502), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n9568) );
  INV_X1 U12068 ( .A(P1_REG3_REG_2__SCAN_IN), .ZN(n10161) );
  OR2_X1 U12069 ( .A1(n6475), .A2(n10161), .ZN(n9567) );
  INV_X1 U12070 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n9563) );
  OR2_X1 U12071 ( .A1(n9853), .A2(n9563), .ZN(n9566) );
  OR2_X1 U12072 ( .A1(n9593), .A2(n9564), .ZN(n9565) );
  AND2_X2 U12073 ( .A1(n11364), .A2(n11543), .ZN(n9620) );
  NAND2_X1 U12074 ( .A1(n9620), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n9569) );
  INV_X4 U12075 ( .A(n11364), .ZN(n11317) );
  AOI22_X1 U12076 ( .A1(n13485), .A2(n14525), .B1(n9619), .B2(n10164), .ZN(
        n9590) );
  NAND2_X1 U12077 ( .A1(n14525), .A2(n9619), .ZN(n9572) );
  OR2_X1 U12078 ( .A1(n13535), .A2(n14555), .ZN(n9571) );
  NAND2_X1 U12079 ( .A1(n9572), .A2(n9571), .ZN(n9573) );
  NAND2_X1 U12080 ( .A1(n14544), .A2(n13806), .ZN(n9941) );
  NAND2_X4 U12081 ( .A1(n9941), .A2(n9940), .ZN(n13536) );
  XNOR2_X1 U12082 ( .A(n9573), .B(n13536), .ZN(n9588) );
  INV_X1 U12083 ( .A(n9588), .ZN(n9589) );
  NAND2_X1 U12084 ( .A1(n6479), .A2(n9619), .ZN(n9582) );
  NAND2_X1 U12085 ( .A1(n9620), .A2(P2_DATAO_REG_1__SCAN_IN), .ZN(n9580) );
  INV_X1 U12086 ( .A(n9576), .ZN(n9577) );
  NAND2_X1 U12087 ( .A1(n9599), .A2(n9577), .ZN(n9579) );
  NAND2_X1 U12088 ( .A1(n11317), .A2(n13673), .ZN(n9578) );
  OR2_X1 U12089 ( .A1(n13535), .A2(n14550), .ZN(n9581) );
  NAND2_X1 U12090 ( .A1(n9582), .A2(n9581), .ZN(n9583) );
  XNOR2_X1 U12091 ( .A(n9583), .B(n13471), .ZN(n9585) );
  NAND2_X1 U12092 ( .A1(n9585), .A2(n9584), .ZN(n9586) );
  OAI21_X1 U12093 ( .B1(n9585), .B2(n9584), .A(n9586), .ZN(n9644) );
  INV_X1 U12094 ( .A(n9586), .ZN(n9587) );
  XOR2_X1 U12095 ( .A(n9590), .B(n9588), .Z(n9651) );
  NAND2_X1 U12096 ( .A1(n11503), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n9598) );
  OR2_X1 U12097 ( .A1(n6487), .A2(n9591), .ZN(n9597) );
  OR2_X1 U12098 ( .A1(n9593), .A2(n9592), .ZN(n9596) );
  OR2_X1 U12099 ( .A1(n6475), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n9595) );
  NAND4_X2 U12100 ( .A1(n9598), .A2(n9597), .A3(n9596), .A4(n9595), .ZN(n13666) );
  NAND2_X1 U12101 ( .A1(n13666), .A2(n9619), .ZN(n9605) );
  NAND2_X1 U12102 ( .A1(n9599), .A2(n9600), .ZN(n9603) );
  NAND2_X1 U12103 ( .A1(n9620), .A2(P2_DATAO_REG_3__SCAN_IN), .ZN(n9602) );
  NAND2_X1 U12104 ( .A1(n11317), .A2(n13703), .ZN(n9601) );
  OR2_X1 U12105 ( .A1(n13535), .A2(n11160), .ZN(n9604) );
  NAND2_X1 U12106 ( .A1(n9605), .A2(n9604), .ZN(n9606) );
  XNOR2_X1 U12107 ( .A(n9606), .B(n13536), .ZN(n9609) );
  INV_X1 U12108 ( .A(n11160), .ZN(n13519) );
  AOI22_X1 U12109 ( .A1(n13485), .A2(n13666), .B1(n9619), .B2(n13519), .ZN(
        n9607) );
  XNOR2_X1 U12110 ( .A(n9609), .B(n9607), .ZN(n13517) );
  NAND2_X1 U12111 ( .A1(n13518), .A2(n13517), .ZN(n9835) );
  INV_X1 U12112 ( .A(n9607), .ZN(n9608) );
  NAND2_X1 U12113 ( .A1(n9609), .A2(n9608), .ZN(n9831) );
  NAND2_X1 U12114 ( .A1(n9835), .A2(n9831), .ZN(n9631) );
  NAND2_X1 U12115 ( .A1(n11503), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n9618) );
  OR2_X1 U12116 ( .A1(n6487), .A2(n9610), .ZN(n9617) );
  INV_X1 U12117 ( .A(n9633), .ZN(n9614) );
  INV_X1 U12118 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n9612) );
  INV_X1 U12119 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n9611) );
  NAND2_X1 U12120 ( .A1(n9612), .A2(n9611), .ZN(n9613) );
  NAND2_X1 U12121 ( .A1(n9614), .A2(n9613), .ZN(n9947) );
  OR2_X1 U12122 ( .A1(n6476), .A2(n9947), .ZN(n9616) );
  NAND2_X1 U12123 ( .A1(n13485), .A2(n13665), .ZN(n9626) );
  NAND2_X1 U12124 ( .A1(n11547), .A2(n9621), .ZN(n9623) );
  NAND2_X1 U12125 ( .A1(n11317), .A2(n13721), .ZN(n9622) );
  NAND2_X1 U12126 ( .A1(n13442), .A2(n11228), .ZN(n9625) );
  AND2_X1 U12127 ( .A1(n9626), .A2(n9625), .ZN(n9832) );
  INV_X1 U12128 ( .A(n9832), .ZN(n9838) );
  NAND2_X1 U12129 ( .A1(n13665), .A2(n13442), .ZN(n9628) );
  NAND2_X1 U12130 ( .A1(n13481), .A2(n11228), .ZN(n9627) );
  NAND2_X1 U12131 ( .A1(n9628), .A2(n9627), .ZN(n9629) );
  XNOR2_X1 U12132 ( .A(n9629), .B(n13471), .ZN(n9836) );
  XNOR2_X1 U12133 ( .A(n9838), .B(n9836), .ZN(n9630) );
  XNOR2_X1 U12134 ( .A(n9631), .B(n9630), .ZN(n9642) );
  OR2_X1 U12135 ( .A1(n11538), .A2(n8743), .ZN(n14006) );
  NOR2_X2 U12136 ( .A1(n13513), .A2(n14006), .ZN(n13620) );
  NAND2_X1 U12137 ( .A1(P1_REG3_REG_4__SCAN_IN), .A2(P1_U3086), .ZN(n13722) );
  NAND2_X1 U12138 ( .A1(n11503), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n9637) );
  OR2_X1 U12139 ( .A1(n9593), .A2(n14619), .ZN(n9636) );
  OR2_X1 U12140 ( .A1(n6487), .A2(n10303), .ZN(n9635) );
  OAI21_X1 U12141 ( .B1(n9633), .B2(P1_REG3_REG_5__SCAN_IN), .A(n9851), .ZN(
        n10307) );
  OR2_X1 U12142 ( .A1(n6468), .A2(n10307), .ZN(n9634) );
  NAND2_X1 U12143 ( .A1(n13639), .A2(n13664), .ZN(n9638) );
  OAI211_X1 U12144 ( .C1(n13644), .C2(n9947), .A(n13722), .B(n9638), .ZN(n9640) );
  NOR2_X1 U12145 ( .A1(n13636), .A2(n14561), .ZN(n9639) );
  AOI211_X1 U12146 ( .C1(n13620), .C2(n13666), .A(n9640), .B(n9639), .ZN(n9641) );
  OAI21_X1 U12147 ( .B1(n9642), .B2(n13650), .A(n9641), .ZN(P1_U3230) );
  AOI21_X1 U12148 ( .B1(n9645), .B2(n9644), .A(n9643), .ZN(n9649) );
  AOI22_X1 U12149 ( .A1(n13620), .A2(n14526), .B1(n13639), .B2(n14525), .ZN(
        n9646) );
  OAI21_X1 U12150 ( .B1(n14550), .B2(n13636), .A(n9646), .ZN(n9647) );
  AOI21_X1 U12151 ( .B1(P1_REG3_REG_1__SCAN_IN), .B2(n9655), .A(n9647), .ZN(
        n9648) );
  OAI21_X1 U12152 ( .B1(n9649), .B2(n13650), .A(n9648), .ZN(P1_U3222) );
  AOI21_X1 U12153 ( .B1(n9652), .B2(n9651), .A(n9650), .ZN(n9657) );
  AOI22_X1 U12154 ( .A1(n13620), .A2(n6480), .B1(n13639), .B2(n13666), .ZN(
        n9653) );
  OAI21_X1 U12155 ( .B1(n14555), .B2(n13636), .A(n9653), .ZN(n9654) );
  AOI21_X1 U12156 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(n9655), .A(n9654), .ZN(
        n9656) );
  OAI21_X1 U12157 ( .B1(n9657), .B2(n13650), .A(n9656), .ZN(P1_U3237) );
  NOR2_X1 U12158 ( .A1(n11613), .A2(n9658), .ZN(n9659) );
  AND2_X1 U12159 ( .A1(n9937), .A2(n9659), .ZN(n9687) );
  INV_X1 U12160 ( .A(n9660), .ZN(n9661) );
  OAI21_X1 U12161 ( .B1(n9663), .B2(P1_D_REG_0__SCAN_IN), .A(n9661), .ZN(n9665) );
  OR2_X1 U12162 ( .A1(n9663), .A2(n9662), .ZN(n9664) );
  INV_X1 U12163 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n9685) );
  OR2_X1 U12164 ( .A1(n9666), .A2(n13806), .ZN(n14585) );
  NAND2_X1 U12165 ( .A1(n14526), .A2(n9668), .ZN(n14515) );
  OR2_X1 U12166 ( .A1(n6480), .A2(n9667), .ZN(n9670) );
  OR2_X1 U12167 ( .A1(n14525), .A2(n10164), .ZN(n9671) );
  OR2_X1 U12168 ( .A1(n13666), .A2(n11160), .ZN(n11221) );
  NAND2_X1 U12169 ( .A1(n13666), .A2(n11160), .ZN(n11222) );
  OR2_X1 U12170 ( .A1(n9672), .A2(n11219), .ZN(n9673) );
  NAND2_X1 U12171 ( .A1(n9936), .A2(n9673), .ZN(n11155) );
  NAND2_X1 U12172 ( .A1(n14550), .A2(n14546), .ZN(n14517) );
  INV_X1 U12173 ( .A(n9946), .ZN(n9675) );
  NAND2_X1 U12174 ( .A1(n10160), .A2(n13519), .ZN(n9674) );
  NAND2_X1 U12175 ( .A1(n9675), .A2(n9674), .ZN(n11156) );
  OAI22_X1 U12176 ( .A1(n11156), .A2(n14596), .B1(n11160), .B2(n14606), .ZN(
        n9683) );
  NAND2_X1 U12177 ( .A1(n14544), .A2(n11204), .ZN(n9676) );
  NAND2_X1 U12178 ( .A1(n14545), .A2(n7147), .ZN(n11509) );
  NAND2_X1 U12179 ( .A1(n9676), .A2(n11509), .ZN(n14392) );
  OR2_X1 U12180 ( .A1(n14526), .A2(n14546), .ZN(n11212) );
  NAND2_X1 U12181 ( .A1(n11209), .A2(n11212), .ZN(n9677) );
  AND2_X1 U12182 ( .A1(n9677), .A2(n11213), .ZN(n10154) );
  NAND2_X1 U12183 ( .A1(n10154), .A2(n11576), .ZN(n10153) );
  NOR2_X1 U12184 ( .A1(n14525), .A2(n14555), .ZN(n11216) );
  INV_X1 U12185 ( .A(n11216), .ZN(n9678) );
  XNOR2_X1 U12186 ( .A(n11219), .B(n9949), .ZN(n9682) );
  AOI21_X1 U12187 ( .B1(n14544), .B2(n11190), .A(n11204), .ZN(n9679) );
  NAND2_X1 U12188 ( .A1(n13536), .A2(n9679), .ZN(n14023) );
  NAND2_X1 U12189 ( .A1(n11155), .A2(n14523), .ZN(n9681) );
  AOI22_X1 U12190 ( .A1(n14527), .A2(n14525), .B1(n13665), .B2(n14524), .ZN(
        n9680) );
  OAI211_X1 U12191 ( .C1(n14542), .C2(n9682), .A(n9681), .B(n9680), .ZN(n11154) );
  AOI211_X1 U12192 ( .C1(n14599), .C2(n11155), .A(n9683), .B(n11154), .ZN(
        n9688) );
  OR2_X1 U12193 ( .A1(n9688), .A2(n14611), .ZN(n9684) );
  OAI21_X1 U12194 ( .B1(n14613), .B2(n9685), .A(n9684), .ZN(P1_U3468) );
  OR2_X1 U12195 ( .A1(n9688), .A2(n14627), .ZN(n9689) );
  OAI21_X1 U12196 ( .B1(n14630), .B2(n9592), .A(n9689), .ZN(P1_U3531) );
  INV_X1 U12197 ( .A(n9690), .ZN(n14705) );
  AOI22_X1 U12198 ( .A1(n12710), .A2(n13065), .B1(n13063), .B2(n12711), .ZN(
        n14702) );
  NAND2_X1 U12199 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3088), .ZN(n14650) );
  OAI21_X1 U12200 ( .B1(n12715), .B2(n14702), .A(n14650), .ZN(n9691) );
  AOI21_X1 U12201 ( .B1(n12754), .B2(n14331), .A(n9691), .ZN(n9697) );
  OAI21_X1 U12202 ( .B1(n9694), .B2(n9693), .A(n9692), .ZN(n9695) );
  NAND2_X1 U12203 ( .A1(n9695), .A2(n14328), .ZN(n9696) );
  OAI211_X1 U12204 ( .C1(n14334), .C2(n14705), .A(n9697), .B(n9696), .ZN(
        P2_U3202) );
  OAI21_X1 U12205 ( .B1(n9700), .B2(n9699), .A(n9698), .ZN(n9701) );
  NAND2_X1 U12206 ( .A1(n9701), .A2(n14328), .ZN(n9705) );
  NAND2_X1 U12207 ( .A1(P2_REG3_REG_5__SCAN_IN), .A2(P2_U3088), .ZN(n14663) );
  OAI21_X1 U12208 ( .B1(n12715), .B2(n9702), .A(n14663), .ZN(n9703) );
  AOI21_X1 U12209 ( .B1(n12773), .B2(n14331), .A(n9703), .ZN(n9704) );
  OAI211_X1 U12210 ( .C1(n14334), .C2(n9706), .A(n9705), .B(n9704), .ZN(
        P2_U3199) );
  XNOR2_X1 U12211 ( .A(n9708), .B(n9707), .ZN(n9714) );
  NAND2_X1 U12212 ( .A1(P2_U3088), .A2(P2_REG3_REG_6__SCAN_IN), .ZN(n13086) );
  NAND2_X1 U12213 ( .A1(n14331), .A2(n12776), .ZN(n9709) );
  OAI211_X1 U12214 ( .C1(n12715), .C2(n9710), .A(n13086), .B(n9709), .ZN(n9711) );
  AOI21_X1 U12215 ( .B1(n9712), .B2(n12717), .A(n9711), .ZN(n9713) );
  OAI21_X1 U12216 ( .B1(n9714), .B2(n12705), .A(n9713), .ZN(P2_U3211) );
  INV_X1 U12217 ( .A(P3_REG3_REG_2__SCAN_IN), .ZN(n9724) );
  XNOR2_X1 U12218 ( .A(n9715), .B(n11971), .ZN(n9990) );
  XNOR2_X1 U12219 ( .A(n9992), .B(n9990), .ZN(n9719) );
  NAND2_X1 U12220 ( .A1(n9717), .A2(n9716), .ZN(n9718) );
  NAND2_X1 U12221 ( .A1(n9718), .A2(n9719), .ZN(n9994) );
  OAI21_X1 U12222 ( .B1(n9719), .B2(n9718), .A(n9994), .ZN(n9720) );
  NAND2_X1 U12223 ( .A1(n9720), .A2(n14276), .ZN(n9723) );
  AOI22_X1 U12224 ( .A1(n12440), .A2(n12142), .B1(n12140), .B2(n12437), .ZN(
        n10121) );
  INV_X1 U12225 ( .A(n10121), .ZN(n9721) );
  AOI22_X1 U12226 ( .A1(n9721), .A2(n12104), .B1(n10117), .B2(n14274), .ZN(
        n9722) );
  OAI211_X1 U12227 ( .C1(n9725), .C2(n9724), .A(n9723), .B(n9722), .ZN(
        P3_U3177) );
  INV_X1 U12228 ( .A(n9728), .ZN(n9729) );
  OR2_X1 U12229 ( .A1(n10199), .A2(n12931), .ZN(n9733) );
  AOI22_X1 U12230 ( .A1(n9097), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n9142), .B2(
        n9731), .ZN(n9732) );
  NAND2_X2 U12231 ( .A1(n9733), .A2(n9732), .ZN(n14781) );
  XNOR2_X1 U12232 ( .A(n14781), .B(n11628), .ZN(n9734) );
  NAND2_X1 U12233 ( .A1(n13060), .A2(n11749), .ZN(n9735) );
  NAND2_X1 U12234 ( .A1(n9734), .A2(n9735), .ZN(n9922) );
  INV_X1 U12235 ( .A(n9734), .ZN(n9737) );
  INV_X1 U12236 ( .A(n9735), .ZN(n9736) );
  NAND2_X1 U12237 ( .A1(n9737), .A2(n9736), .ZN(n9738) );
  NAND2_X1 U12238 ( .A1(n9922), .A2(n9738), .ZN(n9739) );
  AOI21_X1 U12239 ( .B1(n9740), .B2(n9739), .A(n7251), .ZN(n9756) );
  INV_X1 U12240 ( .A(n9741), .ZN(n9781) );
  NAND2_X1 U12241 ( .A1(n13061), .A2(n12710), .ZN(n9751) );
  NAND2_X1 U12242 ( .A1(n11123), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n9749) );
  NAND2_X1 U12243 ( .A1(n11701), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n9748) );
  INV_X1 U12244 ( .A(n9744), .ZN(n9742) );
  AOI21_X1 U12245 ( .B1(n9742), .B2(P2_REG3_REG_8__SCAN_IN), .A(
        P2_REG3_REG_9__SCAN_IN), .ZN(n9745) );
  NAND2_X1 U12246 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_REG3_REG_8__SCAN_IN), 
        .ZN(n9743) );
  OR2_X1 U12247 ( .A1(n9745), .A2(n9794), .ZN(n9929) );
  INV_X1 U12248 ( .A(n9929), .ZN(n9809) );
  NAND2_X1 U12249 ( .A1(n9145), .A2(n9809), .ZN(n9747) );
  NAND2_X1 U12250 ( .A1(n11688), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n9746) );
  NAND4_X1 U12251 ( .A1(n9749), .A2(n9748), .A3(n9747), .A4(n9746), .ZN(n13059) );
  NAND2_X1 U12252 ( .A1(n13059), .A2(n12711), .ZN(n9750) );
  NAND2_X1 U12253 ( .A1(n9751), .A2(n9750), .ZN(n9778) );
  NAND2_X1 U12254 ( .A1(n14330), .A2(n9778), .ZN(n9753) );
  OAI211_X1 U12255 ( .C1(n14334), .C2(n9781), .A(n9753), .B(n9752), .ZN(n9754)
         );
  AOI21_X1 U12256 ( .B1(n14781), .B2(n12703), .A(n9754), .ZN(n9755) );
  OAI21_X1 U12257 ( .B1(n9756), .B2(n12705), .A(n9755), .ZN(P2_U3193) );
  INV_X1 U12258 ( .A(SI_20_), .ZN(n10533) );
  INV_X1 U12259 ( .A(n9757), .ZN(n9759) );
  OAI222_X1 U12260 ( .A1(n12608), .A2(n10533), .B1(n12607), .B2(n9759), .C1(
        P3_U3151), .C2(n9758), .ZN(P3_U3275) );
  NAND2_X1 U12261 ( .A1(n10112), .A2(P3_STATE_REG_SCAN_IN), .ZN(n9760) );
  OAI21_X1 U12262 ( .B1(n12608), .B2(n9761), .A(n9760), .ZN(n9762) );
  AOI21_X1 U12263 ( .B1(n9763), .B2(n12596), .A(n9762), .ZN(n9764) );
  INV_X1 U12264 ( .A(n9764), .ZN(P3_U3274) );
  INV_X1 U12265 ( .A(n13060), .ZN(n9766) );
  NAND2_X1 U12266 ( .A1(n14781), .A2(n9766), .ZN(n9791) );
  OR2_X1 U12267 ( .A1(n14781), .A2(n9766), .ZN(n9767) );
  XOR2_X1 U12268 ( .A(n9802), .B(n13002), .Z(n9779) );
  INV_X1 U12269 ( .A(n9779), .ZN(n14784) );
  INV_X1 U12270 ( .A(n12721), .ZN(n9768) );
  OR2_X1 U12271 ( .A1(n14731), .A2(n9768), .ZN(n13320) );
  INV_X1 U12272 ( .A(n9769), .ZN(n9772) );
  AND2_X1 U12273 ( .A1(n12791), .A2(n9773), .ZN(n9770) );
  INV_X1 U12274 ( .A(n9770), .ZN(n9771) );
  OR2_X1 U12275 ( .A1(n12791), .A2(n9773), .ZN(n9774) );
  NAND2_X1 U12276 ( .A1(n9775), .A2(n13002), .ZN(n9776) );
  AOI21_X1 U12277 ( .B1(n9792), .B2(n9776), .A(n14352), .ZN(n9777) );
  AOI211_X1 U12278 ( .C1(n9779), .C2(n14741), .A(n9778), .B(n9777), .ZN(n14783) );
  MUX2_X1 U12279 ( .A(n8877), .B(n14783), .S(n13316), .Z(n9785) );
  AOI211_X1 U12280 ( .C1(n14781), .C2(n9780), .A(n9329), .B(n9807), .ZN(n14780) );
  INV_X1 U12281 ( .A(n14781), .ZN(n9782) );
  OAI22_X1 U12282 ( .A1(n9782), .A2(n14721), .B1(n9781), .B2(n14706), .ZN(
        n9783) );
  AOI21_X1 U12283 ( .B1(n14780), .B2(n14725), .A(n9783), .ZN(n9784) );
  OAI211_X1 U12284 ( .C1(n14784), .C2(n13320), .A(n9785), .B(n9784), .ZN(
        P2_U3257) );
  OR2_X1 U12285 ( .A1(n10205), .A2(n12931), .ZN(n9788) );
  AOI22_X1 U12286 ( .A1(n9142), .A2(n9786), .B1(n11862), .B2(
        P1_DATAO_REG_9__SCAN_IN), .ZN(n9787) );
  INV_X1 U12287 ( .A(n13059), .ZN(n9789) );
  NAND2_X1 U12288 ( .A1(n12801), .A2(n9789), .ZN(n10044) );
  OR2_X1 U12289 ( .A1(n12801), .A2(n9789), .ZN(n9790) );
  OAI21_X1 U12290 ( .B1(n13004), .B2(n9793), .A(n10045), .ZN(n9806) );
  NAND2_X1 U12291 ( .A1(n13060), .A2(n12710), .ZN(n9801) );
  NAND2_X1 U12292 ( .A1(n11123), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n9799) );
  NAND2_X1 U12293 ( .A1(n11701), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n9798) );
  NAND2_X1 U12294 ( .A1(n9794), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9964) );
  OR2_X1 U12295 ( .A1(n9794), .A2(P2_REG3_REG_10__SCAN_IN), .ZN(n9795) );
  AND2_X1 U12296 ( .A1(n9964), .A2(n9795), .ZN(n9962) );
  NAND2_X1 U12297 ( .A1(n9145), .A2(n9962), .ZN(n9797) );
  NAND2_X1 U12298 ( .A1(n11688), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n9796) );
  NAND4_X1 U12299 ( .A1(n9799), .A2(n9798), .A3(n9797), .A4(n9796), .ZN(n13058) );
  NAND2_X1 U12300 ( .A1(n13058), .A2(n12711), .ZN(n9800) );
  NAND2_X1 U12301 ( .A1(n9801), .A2(n9800), .ZN(n9926) );
  NAND2_X1 U12302 ( .A1(n9802), .A2(n13002), .ZN(n9804) );
  NAND2_X1 U12303 ( .A1(n14781), .A2(n13060), .ZN(n9803) );
  INV_X1 U12304 ( .A(n13004), .ZN(n10039) );
  XNOR2_X1 U12305 ( .A(n10040), .B(n10039), .ZN(n10018) );
  NOR2_X1 U12306 ( .A1(n10018), .A2(n9328), .ZN(n9805) );
  AOI211_X1 U12307 ( .C1(n14740), .C2(n9806), .A(n9926), .B(n9805), .ZN(n10017) );
  INV_X1 U12308 ( .A(n9807), .ZN(n9808) );
  INV_X1 U12309 ( .A(n12801), .ZN(n9811) );
  NAND2_X1 U12310 ( .A1(n9811), .A2(n9807), .ZN(n10052) );
  AOI211_X1 U12311 ( .C1(n12801), .C2(n9808), .A(n9329), .B(n6850), .ZN(n10015) );
  AOI22_X1 U12312 ( .A1(n14731), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n9809), .B2(
        n14719), .ZN(n9810) );
  OAI21_X1 U12313 ( .B1(n9811), .B2(n14721), .A(n9810), .ZN(n9813) );
  NOR2_X1 U12314 ( .A1(n10018), .A2(n13320), .ZN(n9812) );
  AOI211_X1 U12315 ( .C1(n10015), .C2(n14725), .A(n9813), .B(n9812), .ZN(n9814) );
  OAI21_X1 U12316 ( .B1(n10017), .B2(n14708), .A(n9814), .ZN(P2_U3256) );
  OAI21_X1 U12317 ( .B1(n9817), .B2(n15072), .A(n9816), .ZN(n9819) );
  NAND2_X1 U12318 ( .A1(n9817), .A2(n15072), .ZN(n9818) );
  MUX2_X1 U12319 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(P1_DATAO_REG_18__SCAN_IN), 
        .S(n11543), .Z(n9933) );
  INV_X1 U12320 ( .A(n11316), .ZN(n9830) );
  OAI21_X1 U12321 ( .B1(n9822), .B2(P1_IR_REG_17__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .ZN(n9823) );
  XNOR2_X1 U12322 ( .A(n9823), .B(P1_IR_REG_18__SCAN_IN), .ZN(n13797) );
  INV_X1 U12323 ( .A(n13797), .ZN(n10959) );
  OAI222_X1 U12324 ( .A1(n14124), .A2(n9824), .B1(n14119), .B2(n9830), .C1(
        n10959), .C2(P1_U3086), .ZN(P1_U3337) );
  NAND2_X1 U12325 ( .A1(n9826), .A2(n9825), .ZN(n9827) );
  NAND2_X1 U12326 ( .A1(n9827), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n9828) );
  XNOR2_X1 U12327 ( .A(n9828), .B(P2_IR_REG_18__SCAN_IN), .ZN(n13149) );
  INV_X1 U12328 ( .A(n13149), .ZN(n13134) );
  INV_X1 U12329 ( .A(P1_DATAO_REG_18__SCAN_IN), .ZN(n9829) );
  OAI222_X1 U12330 ( .A1(P2_U3088), .A2(n13134), .B1(n13438), .B2(n9830), .C1(
        n9829), .C2(n13440), .ZN(P2_U3309) );
  NAND2_X1 U12331 ( .A1(n9835), .A2(n9834), .ZN(n9840) );
  INV_X1 U12332 ( .A(n9836), .ZN(n9837) );
  NAND2_X1 U12333 ( .A1(n9840), .A2(n9839), .ZN(n9910) );
  NAND2_X1 U12334 ( .A1(n9841), .A2(n9599), .ZN(n9843) );
  INV_X2 U12335 ( .A(n9846), .ZN(n11548) );
  AOI22_X1 U12336 ( .A1(n11548), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n11317), 
        .B2(n13731), .ZN(n9842) );
  NAND2_X1 U12337 ( .A1(n9843), .A2(n9842), .ZN(n11233) );
  AOI22_X1 U12338 ( .A1(n13485), .A2(n13664), .B1(n13442), .B2(n11233), .ZN(
        n9864) );
  AOI22_X1 U12339 ( .A1(n13664), .A2(n13442), .B1(n13481), .B2(n11233), .ZN(
        n9844) );
  XNOR2_X1 U12340 ( .A(n9844), .B(n13536), .ZN(n9865) );
  XOR2_X1 U12341 ( .A(n9864), .B(n9865), .Z(n9911) );
  NAND2_X1 U12342 ( .A1(n9910), .A2(n9911), .ZN(n9866) );
  OR2_X1 U12343 ( .A1(n9845), .A2(n11490), .ZN(n9849) );
  AOI22_X1 U12344 ( .A1(n11548), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n11317), 
        .B2(n9847), .ZN(n9848) );
  NAND2_X1 U12345 ( .A1(n9849), .A2(n9848), .ZN(n11238) );
  NAND2_X1 U12346 ( .A1(n11238), .A2(n13481), .ZN(n9860) );
  NAND2_X1 U12347 ( .A1(n6473), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n9858) );
  OR2_X1 U12348 ( .A1(n6487), .A2(n10289), .ZN(n9857) );
  AND2_X1 U12349 ( .A1(n9851), .A2(n9850), .ZN(n9852) );
  OR2_X1 U12350 ( .A1(n9852), .A2(n9869), .ZN(n10292) );
  OR2_X1 U12351 ( .A1(n11470), .A2(n10292), .ZN(n9856) );
  INV_X1 U12352 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n9854) );
  OR2_X1 U12353 ( .A1(n11516), .A2(n9854), .ZN(n9855) );
  NAND4_X1 U12354 ( .A1(n9858), .A2(n9857), .A3(n9856), .A4(n9855), .ZN(n13663) );
  NAND2_X1 U12355 ( .A1(n13663), .A2(n13442), .ZN(n9859) );
  NAND2_X1 U12356 ( .A1(n9860), .A2(n9859), .ZN(n9861) );
  XNOR2_X1 U12357 ( .A(n9861), .B(n13471), .ZN(n10169) );
  NAND2_X1 U12358 ( .A1(n13485), .A2(n13663), .ZN(n9863) );
  NAND2_X1 U12359 ( .A1(n11238), .A2(n13442), .ZN(n9862) );
  NAND2_X1 U12360 ( .A1(n9863), .A2(n9862), .ZN(n10167) );
  XNOR2_X1 U12361 ( .A(n10169), .B(n10167), .ZN(n9867) );
  NAND2_X1 U12362 ( .A1(n9865), .A2(n9864), .ZN(n9868) );
  NAND2_X1 U12363 ( .A1(n10171), .A2(n13626), .ZN(n9882) );
  AOI21_X1 U12364 ( .B1(n9866), .B2(n9868), .A(n9867), .ZN(n9881) );
  NAND2_X1 U12365 ( .A1(n11503), .A2(P1_REG0_REG_7__SCAN_IN), .ZN(n9875) );
  OR2_X1 U12366 ( .A1(n6487), .A2(n10319), .ZN(n9874) );
  OR2_X1 U12367 ( .A1(n9869), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n9870) );
  NAND2_X1 U12368 ( .A1(n10181), .A2(n9870), .ZN(n10321) );
  OR2_X1 U12369 ( .A1(n11470), .A2(n10321), .ZN(n9873) );
  OR2_X1 U12370 ( .A1(n6483), .A2(n9871), .ZN(n9872) );
  NAND4_X1 U12371 ( .A1(n9875), .A2(n9874), .A3(n9873), .A4(n9872), .ZN(n13662) );
  NAND2_X1 U12372 ( .A1(n13639), .A2(n13662), .ZN(n9876) );
  OAI211_X1 U12373 ( .C1(n13644), .C2(n10292), .A(n9877), .B(n9876), .ZN(n9879) );
  INV_X1 U12374 ( .A(n11238), .ZN(n14573) );
  NOR2_X1 U12375 ( .A1(n13636), .A2(n14573), .ZN(n9878) );
  AOI211_X1 U12376 ( .C1(n13620), .C2(n13664), .A(n9879), .B(n9878), .ZN(n9880) );
  OAI21_X1 U12377 ( .B1(n9882), .B2(n9881), .A(n9880), .ZN(P1_U3239) );
  INV_X1 U12378 ( .A(n9883), .ZN(n9884) );
  XNOR2_X1 U12379 ( .A(n12585), .B(n9884), .ZN(n9885) );
  NAND3_X1 U12380 ( .A1(n9887), .A2(n9886), .A3(n9885), .ZN(n9890) );
  INV_X1 U12381 ( .A(n14969), .ZN(n10118) );
  OR2_X1 U12382 ( .A1(n9890), .A2(n10118), .ZN(n12458) );
  NOR2_X1 U12383 ( .A1(n14298), .A2(n14969), .ZN(n9888) );
  NAND2_X1 U12384 ( .A1(n10110), .A2(n14977), .ZN(n9893) );
  AOI22_X1 U12385 ( .A1(n14979), .A2(P3_REG2_REG_0__SCAN_IN), .B1(
        P3_REG3_REG_0__SCAN_IN), .B2(n14973), .ZN(n9892) );
  OAI211_X1 U12386 ( .C1(n10108), .C2(n14906), .A(n9893), .B(n9892), .ZN(
        P3_U3233) );
  AOI21_X1 U12387 ( .B1(n9896), .B2(n9895), .A(n9894), .ZN(n9909) );
  OAI21_X1 U12388 ( .B1(n9899), .B2(n9898), .A(n9897), .ZN(n9907) );
  AOI22_X1 U12389 ( .A1(n14869), .A2(P3_ADDR_REG_7__SCAN_IN), .B1(
        P3_REG3_REG_7__SCAN_IN), .B2(P3_U3151), .ZN(n9900) );
  OAI21_X1 U12390 ( .B1(n14878), .B2(n9901), .A(n9900), .ZN(n9906) );
  AOI21_X1 U12391 ( .B1(n15030), .B2(n9903), .A(n9902), .ZN(n9904) );
  NOR2_X1 U12392 ( .A1(n9904), .A2(n14887), .ZN(n9905) );
  AOI211_X1 U12393 ( .C1(n14843), .C2(n9907), .A(n9906), .B(n9905), .ZN(n9908)
         );
  OAI21_X1 U12394 ( .B1(n9909), .B2(n14893), .A(n9908), .ZN(P3_U3189) );
  OAI21_X1 U12395 ( .B1(n9911), .B2(n9910), .A(n9866), .ZN(n9915) );
  INV_X1 U12396 ( .A(n13620), .ZN(n13629) );
  OAI22_X1 U12397 ( .A1(n13636), .A2(n6874), .B1(n13629), .B2(n10192), .ZN(
        n9914) );
  NAND2_X1 U12398 ( .A1(P1_REG3_REG_5__SCAN_IN), .A2(P1_U3086), .ZN(n13729) );
  NAND2_X1 U12399 ( .A1(n13639), .A2(n13663), .ZN(n9912) );
  OAI211_X1 U12400 ( .C1(n13644), .C2(n10307), .A(n13729), .B(n9912), .ZN(
        n9913) );
  AOI211_X1 U12401 ( .C1(n9915), .C2(n13626), .A(n9914), .B(n9913), .ZN(n9916)
         );
  INV_X1 U12402 ( .A(n9916), .ZN(P1_U3227) );
  XNOR2_X1 U12403 ( .A(n12801), .B(n11628), .ZN(n9917) );
  NAND2_X1 U12404 ( .A1(n13059), .A2(n11749), .ZN(n9918) );
  NAND2_X1 U12405 ( .A1(n9917), .A2(n9918), .ZN(n9957) );
  INV_X1 U12406 ( .A(n9917), .ZN(n9920) );
  INV_X1 U12407 ( .A(n9918), .ZN(n9919) );
  NAND2_X1 U12408 ( .A1(n9920), .A2(n9919), .ZN(n9921) );
  AND2_X1 U12409 ( .A1(n9957), .A2(n9921), .ZN(n9925) );
  OAI21_X1 U12410 ( .B1(n9925), .B2(n9924), .A(n9958), .ZN(n9931) );
  NAND2_X1 U12411 ( .A1(n12801), .A2(n14331), .ZN(n9928) );
  AOI22_X1 U12412 ( .A1(n14330), .A2(n9926), .B1(P2_REG3_REG_9__SCAN_IN), .B2(
        P2_U3088), .ZN(n9927) );
  OAI211_X1 U12413 ( .C1(n14334), .C2(n9929), .A(n9928), .B(n9927), .ZN(n9930)
         );
  AOI21_X1 U12414 ( .B1(n9931), .B2(n14328), .A(n9930), .ZN(n9932) );
  INV_X1 U12415 ( .A(n9932), .ZN(P2_U3203) );
  MUX2_X1 U12416 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(P1_DATAO_REG_19__SCAN_IN), 
        .S(n11543), .Z(n10529) );
  XNOR2_X1 U12417 ( .A(n10529), .B(SI_19_), .ZN(n10531) );
  XNOR2_X1 U12418 ( .A(n10532), .B(n10531), .ZN(n11309) );
  INV_X1 U12419 ( .A(n11309), .ZN(n12012) );
  OAI222_X1 U12420 ( .A1(n14124), .A2(n7510), .B1(n14119), .B2(n12012), .C1(
        P1_U3086), .C2(n13806), .ZN(P1_U3336) );
  XNOR2_X1 U12421 ( .A(n13665), .B(n14561), .ZN(n11578) );
  OR2_X1 U12422 ( .A1(n13666), .A2(n13519), .ZN(n9935) );
  XOR2_X1 U12423 ( .A(n11578), .B(n10193), .Z(n14560) );
  NOR2_X1 U12424 ( .A1(n9937), .A2(n11613), .ZN(n9939) );
  INV_X2 U12425 ( .A(n14388), .ZN(n13893) );
  OAI21_X1 U12426 ( .B1(n9941), .B2(n9940), .A(n13536), .ZN(n9942) );
  INV_X1 U12427 ( .A(n9942), .ZN(n9943) );
  NAND2_X1 U12428 ( .A1(n9946), .A2(n14561), .ZN(n10304) );
  OAI21_X1 U12429 ( .B1(n9946), .B2(n14561), .A(n10304), .ZN(n14562) );
  OAI22_X1 U12430 ( .A1(n13989), .A2(n14562), .B1(n9947), .B2(n14532), .ZN(
        n9948) );
  AOI21_X1 U12431 ( .B1(n14398), .B2(n11228), .A(n9948), .ZN(n9956) );
  INV_X1 U12432 ( .A(n11219), .ZN(n11577) );
  INV_X1 U12433 ( .A(n11578), .ZN(n9950) );
  XNOR2_X1 U12434 ( .A(n10216), .B(n9950), .ZN(n9951) );
  NAND2_X1 U12435 ( .A1(n9951), .A2(n14392), .ZN(n9953) );
  AOI22_X1 U12436 ( .A1(n14527), .A2(n13666), .B1(n13664), .B2(n14524), .ZN(
        n9952) );
  NAND2_X1 U12437 ( .A1(n9953), .A2(n9952), .ZN(n14564) );
  MUX2_X1 U12438 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n14564), .S(n13893), .Z(
        n9954) );
  INV_X1 U12439 ( .A(n9954), .ZN(n9955) );
  OAI211_X1 U12440 ( .C1(n14560), .C2(n14015), .A(n9956), .B(n9955), .ZN(
        P1_U3289) );
  NAND2_X1 U12441 ( .A1(n10456), .A2(n11860), .ZN(n9961) );
  AOI22_X1 U12442 ( .A1(n9959), .A2(n9142), .B1(P1_DATAO_REG_10__SCAN_IN), 
        .B2(n9097), .ZN(n9960) );
  XNOR2_X1 U12443 ( .A(n14789), .B(n11628), .ZN(n10391) );
  NAND2_X1 U12444 ( .A1(n13058), .A2(n11749), .ZN(n10390) );
  XNOR2_X1 U12445 ( .A(n10391), .B(n10390), .ZN(n10392) );
  XNOR2_X1 U12446 ( .A(n10393), .B(n10392), .ZN(n9976) );
  INV_X1 U12447 ( .A(n9962), .ZN(n10053) );
  NAND2_X1 U12448 ( .A1(n13059), .A2(n12710), .ZN(n9971) );
  NAND2_X1 U12449 ( .A1(n11123), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n9969) );
  NAND2_X1 U12450 ( .A1(n11701), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n9968) );
  NAND2_X1 U12451 ( .A1(n9964), .A2(n9963), .ZN(n9965) );
  AND2_X1 U12452 ( .A1(n10064), .A2(n9965), .ZN(n10404) );
  NAND2_X1 U12453 ( .A1(n9145), .A2(n10404), .ZN(n9967) );
  NAND2_X1 U12454 ( .A1(n11688), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n9966) );
  NAND4_X1 U12455 ( .A1(n9969), .A2(n9968), .A3(n9967), .A4(n9966), .ZN(n13057) );
  NAND2_X1 U12456 ( .A1(n13057), .A2(n12711), .ZN(n9970) );
  NAND2_X1 U12457 ( .A1(n9971), .A2(n9970), .ZN(n10048) );
  INV_X1 U12458 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n9972) );
  NOR2_X1 U12459 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n9972), .ZN(n14665) );
  AOI21_X1 U12460 ( .B1(n14330), .B2(n10048), .A(n14665), .ZN(n9973) );
  OAI21_X1 U12461 ( .B1(n10053), .B2(n14334), .A(n9973), .ZN(n9974) );
  AOI21_X1 U12462 ( .B1(n14789), .B2(n12703), .A(n9974), .ZN(n9975) );
  OAI21_X1 U12463 ( .B1(n9976), .B2(n12705), .A(n9975), .ZN(P2_U3189) );
  INV_X1 U12464 ( .A(n9977), .ZN(n9980) );
  OAI22_X1 U12465 ( .A1(n9978), .A2(P3_U3151), .B1(SI_22_), .B2(n12589), .ZN(
        n9979) );
  AOI21_X1 U12466 ( .B1(n9980), .B2(n12596), .A(n9979), .ZN(P3_U3273) );
  NAND2_X1 U12467 ( .A1(n14526), .A2(n14546), .ZN(n11191) );
  AND2_X1 U12468 ( .A1(n11212), .A2(n11191), .ZN(n14540) );
  AND2_X1 U12469 ( .A1(n13893), .A2(n14392), .ZN(n12010) );
  NOR2_X1 U12470 ( .A1(n14383), .A2(n12010), .ZN(n9985) );
  NAND2_X1 U12471 ( .A1(n6479), .A2(n14524), .ZN(n14543) );
  OAI22_X1 U12472 ( .A1(n14388), .A2(n14543), .B1(n9981), .B2(n14532), .ZN(
        n9983) );
  AOI21_X1 U12473 ( .B1(n14534), .B2(n13989), .A(n14546), .ZN(n9982) );
  AOI211_X1 U12474 ( .C1(n14388), .C2(P1_REG2_REG_0__SCAN_IN), .A(n9983), .B(
        n9982), .ZN(n9984) );
  OAI21_X1 U12475 ( .B1(n14540), .B2(n9985), .A(n9984), .ZN(P1_U3293) );
  INV_X1 U12476 ( .A(P3_REG3_REG_3__SCAN_IN), .ZN(n15067) );
  OR2_X1 U12477 ( .A1(n10033), .A2(n12100), .ZN(n9986) );
  OAI21_X1 U12478 ( .B1(n9992), .B2(n12103), .A(n9986), .ZN(n14952) );
  NAND2_X1 U12479 ( .A1(n14952), .A2(n12104), .ZN(n9988) );
  OAI211_X1 U12480 ( .C1(n12095), .C2(n9989), .A(n9988), .B(n9987), .ZN(n9999)
         );
  XNOR2_X1 U12481 ( .A(n9989), .B(n6508), .ZN(n10025) );
  XNOR2_X1 U12482 ( .A(n10025), .B(n12140), .ZN(n9995) );
  INV_X1 U12483 ( .A(n9990), .ZN(n9991) );
  NAND2_X1 U12484 ( .A1(n9992), .A2(n9991), .ZN(n9996) );
  AND2_X1 U12485 ( .A1(n9996), .A2(n9995), .ZN(n9993) );
  NAND2_X1 U12486 ( .A1(n9994), .A2(n9993), .ZN(n10028) );
  INV_X1 U12487 ( .A(n10028), .ZN(n10101) );
  AOI21_X1 U12488 ( .B1(n9994), .B2(n9996), .A(n9995), .ZN(n9997) );
  NOR3_X1 U12489 ( .A1(n10101), .A2(n9997), .A3(n12115), .ZN(n9998) );
  AOI211_X1 U12490 ( .C1(n15067), .C2(n12112), .A(n9999), .B(n9998), .ZN(
        n10000) );
  INV_X1 U12491 ( .A(n10000), .ZN(P3_U3158) );
  INV_X1 U12492 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10564) );
  INV_X1 U12493 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n14373) );
  AOI21_X1 U12494 ( .B1(n10059), .B2(P2_REG1_REG_11__SCAN_IN), .A(n10001), 
        .ZN(n13124) );
  MUX2_X1 U12495 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n14373), .S(n10129), .Z(
        n13123) );
  AOI21_X1 U12496 ( .B1(n14373), .B2(n13120), .A(n13125), .ZN(n14689) );
  MUX2_X1 U12497 ( .A(n10564), .B(P2_REG1_REG_13__SCAN_IN), .S(n10247), .Z(
        n14688) );
  NAND2_X1 U12498 ( .A1(n14689), .A2(n14688), .ZN(n14687) );
  OAI21_X1 U12499 ( .B1(n10564), .B2(n10247), .A(n14687), .ZN(n10004) );
  INV_X1 U12500 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10002) );
  MUX2_X1 U12501 ( .A(P2_REG1_REG_14__SCAN_IN), .B(n10002), .S(n10725), .Z(
        n10003) );
  NAND2_X1 U12502 ( .A1(n10003), .A2(n10004), .ZN(n10478) );
  OAI211_X1 U12503 ( .C1(n10004), .C2(n10003), .A(n14686), .B(n10478), .ZN(
        n10006) );
  NAND2_X1 U12504 ( .A1(n14685), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n10005) );
  OAI211_X1 U12505 ( .C1(n14667), .C2(n10479), .A(n10006), .B(n10005), .ZN(
        n10014) );
  NAND2_X1 U12506 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(P2_U3088), .ZN(n14332)
         );
  INV_X1 U12507 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n10010) );
  INV_X1 U12508 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n10009) );
  NAND2_X1 U12509 ( .A1(n10008), .A2(n10007), .ZN(n13115) );
  MUX2_X1 U12510 ( .A(n10009), .B(P2_REG2_REG_12__SCAN_IN), .S(n10129), .Z(
        n13116) );
  AOI21_X1 U12511 ( .B1(n13117), .B2(n13115), .A(n13116), .ZN(n13119) );
  MUX2_X1 U12512 ( .A(n10010), .B(P2_REG2_REG_13__SCAN_IN), .S(n10247), .Z(
        n14694) );
  NAND2_X1 U12513 ( .A1(n14695), .A2(n14694), .ZN(n14693) );
  OAI21_X1 U12514 ( .B1(n10010), .B2(n10247), .A(n14693), .ZN(n10481) );
  XNOR2_X1 U12515 ( .A(n10479), .B(n10481), .ZN(n10011) );
  NAND2_X1 U12516 ( .A1(P2_REG2_REG_14__SCAN_IN), .A2(n10011), .ZN(n10482) );
  OAI211_X1 U12517 ( .C1(P2_REG2_REG_14__SCAN_IN), .C2(n10011), .A(n14692), 
        .B(n10482), .ZN(n10012) );
  NAND2_X1 U12518 ( .A1(n14332), .A2(n10012), .ZN(n10013) );
  OR2_X1 U12519 ( .A1(n10014), .A2(n10013), .ZN(P2_U3228) );
  INV_X1 U12520 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10020) );
  AOI21_X1 U12521 ( .B1(n12801), .B2(n14788), .A(n10015), .ZN(n10016) );
  OAI211_X1 U12522 ( .C1(n14793), .C2(n10018), .A(n10017), .B(n10016), .ZN(
        n10021) );
  NAND2_X1 U12523 ( .A1(n10021), .A2(n14797), .ZN(n10019) );
  OAI21_X1 U12524 ( .B1(n14797), .B2(n10020), .A(n10019), .ZN(P2_U3457) );
  NAND2_X1 U12525 ( .A1(n10021), .A2(n6470), .ZN(n10022) );
  OAI21_X1 U12526 ( .B1(n6470), .B2(n10023), .A(n10022), .ZN(P2_U3508) );
  INV_X1 U12527 ( .A(n14939), .ZN(n10038) );
  XNOR2_X1 U12528 ( .A(n10364), .B(n11971), .ZN(n10434) );
  XNOR2_X1 U12529 ( .A(n7638), .B(n10434), .ZN(n10031) );
  XNOR2_X1 U12530 ( .A(n10327), .B(n6508), .ZN(n10024) );
  NAND2_X1 U12531 ( .A1(n10033), .A2(n10024), .ZN(n10029) );
  OAI21_X1 U12532 ( .B1(n10033), .B2(n10024), .A(n10029), .ZN(n10099) );
  INV_X1 U12533 ( .A(n10025), .ZN(n10026) );
  AND2_X1 U12534 ( .A1(n12140), .A2(n10026), .ZN(n10100) );
  NOR2_X1 U12535 ( .A1(n10099), .A2(n10100), .ZN(n10027) );
  NAND2_X1 U12536 ( .A1(n10028), .A2(n10027), .ZN(n10102) );
  NAND2_X1 U12537 ( .A1(n10102), .A2(n10029), .ZN(n10030) );
  NAND2_X1 U12538 ( .A1(n10030), .A2(n10031), .ZN(n10511) );
  OAI21_X1 U12539 ( .B1(n10031), .B2(n10030), .A(n10511), .ZN(n10032) );
  NAND2_X1 U12540 ( .A1(n10032), .A2(n14276), .ZN(n10037) );
  INV_X1 U12541 ( .A(n12137), .ZN(n10507) );
  OAI22_X1 U12542 ( .A1(n10507), .A2(n12100), .B1(n10033), .B2(n12103), .ZN(
        n10358) );
  OAI21_X1 U12543 ( .B1(n12095), .B2(n10364), .A(n10034), .ZN(n10035) );
  AOI21_X1 U12544 ( .B1(n10358), .B2(n12104), .A(n10035), .ZN(n10036) );
  OAI211_X1 U12545 ( .C1(n10038), .C2(n14286), .A(n10037), .B(n10036), .ZN(
        P3_U3167) );
  NAND2_X1 U12546 ( .A1(n12801), .A2(n13059), .ZN(n10041) );
  INV_X1 U12547 ( .A(n13058), .ZN(n10042) );
  NAND2_X1 U12548 ( .A1(n14789), .A2(n10042), .ZN(n10057) );
  OR2_X1 U12549 ( .A1(n14789), .A2(n10042), .ZN(n10043) );
  INV_X1 U12550 ( .A(n13005), .ZN(n10072) );
  XNOR2_X1 U12551 ( .A(n10073), .B(n10072), .ZN(n14792) );
  INV_X1 U12552 ( .A(P2_REG2_REG_10__SCAN_IN), .ZN(n10050) );
  NAND2_X1 U12553 ( .A1(n10045), .A2(n10044), .ZN(n10046) );
  NAND2_X1 U12554 ( .A1(n10046), .A2(n13005), .ZN(n10058) );
  OAI21_X1 U12555 ( .B1(n13005), .B2(n10046), .A(n10058), .ZN(n10049) );
  NOR2_X1 U12556 ( .A1(n14792), .A2(n9328), .ZN(n10047) );
  AOI211_X1 U12557 ( .C1(n14740), .C2(n10049), .A(n10048), .B(n10047), .ZN(
        n14791) );
  MUX2_X1 U12558 ( .A(n10050), .B(n14791), .S(n13316), .Z(n10056) );
  INV_X1 U12559 ( .A(n10077), .ZN(n10051) );
  AOI211_X1 U12560 ( .C1(n14789), .C2(n10052), .A(n9329), .B(n10051), .ZN(
        n14787) );
  OAI22_X1 U12561 ( .A1(n6849), .A2(n14721), .B1(n14706), .B2(n10053), .ZN(
        n10054) );
  AOI21_X1 U12562 ( .B1(n14787), .B2(n14725), .A(n10054), .ZN(n10055) );
  OAI211_X1 U12563 ( .C1(n14792), .C2(n13320), .A(n10056), .B(n10055), .ZN(
        P2_U3255) );
  NAND2_X1 U12564 ( .A1(n10058), .A2(n10057), .ZN(n10063) );
  NAND2_X1 U12565 ( .A1(n10615), .A2(n12943), .ZN(n10061) );
  AOI22_X1 U12566 ( .A1(n10059), .A2(n9142), .B1(P1_DATAO_REG_11__SCAN_IN), 
        .B2(n9097), .ZN(n10060) );
  INV_X1 U12567 ( .A(n13057), .ZN(n12812) );
  XNOR2_X1 U12568 ( .A(n12810), .B(n12812), .ZN(n13008) );
  INV_X1 U12569 ( .A(n13008), .ZN(n10062) );
  OAI21_X1 U12570 ( .B1(n10063), .B2(n10062), .A(n10128), .ZN(n10075) );
  NAND2_X1 U12571 ( .A1(n13058), .A2(n12710), .ZN(n10071) );
  NAND2_X1 U12572 ( .A1(n11123), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n10069) );
  NAND2_X1 U12573 ( .A1(n11701), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n10068) );
  NAND2_X1 U12574 ( .A1(n10064), .A2(n10500), .ZN(n10065) );
  NAND2_X1 U12575 ( .A1(n10257), .A2(n10065), .ZN(n10501) );
  INV_X1 U12576 ( .A(n10501), .ZN(n10145) );
  NAND2_X1 U12577 ( .A1(n9145), .A2(n10145), .ZN(n10067) );
  NAND2_X1 U12578 ( .A1(n11688), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n10066) );
  NAND4_X1 U12579 ( .A1(n10069), .A2(n10068), .A3(n10067), .A4(n10066), .ZN(
        n13056) );
  NAND2_X1 U12580 ( .A1(n13056), .A2(n12711), .ZN(n10070) );
  NAND2_X1 U12581 ( .A1(n10071), .A2(n10070), .ZN(n10407) );
  XNOR2_X1 U12582 ( .A(n10140), .B(n13008), .ZN(n10446) );
  NOR2_X1 U12583 ( .A1(n10446), .A2(n9328), .ZN(n10074) );
  AOI211_X1 U12584 ( .C1(n14740), .C2(n10075), .A(n10407), .B(n10074), .ZN(
        n10445) );
  INV_X1 U12585 ( .A(n10142), .ZN(n10076) );
  AOI211_X1 U12586 ( .C1(n12810), .C2(n10077), .A(n9329), .B(n10076), .ZN(
        n10443) );
  AOI22_X1 U12587 ( .A1(n14708), .A2(P2_REG2_REG_11__SCAN_IN), .B1(n10404), 
        .B2(n14719), .ZN(n10078) );
  OAI21_X1 U12588 ( .B1(n6847), .B2(n14721), .A(n10078), .ZN(n10080) );
  NOR2_X1 U12589 ( .A1(n10446), .A2(n13320), .ZN(n10079) );
  AOI211_X1 U12590 ( .C1(n10443), .C2(n14725), .A(n10080), .B(n10079), .ZN(
        n10081) );
  OAI21_X1 U12591 ( .B1(n10445), .B2(n14731), .A(n10081), .ZN(P2_U3254) );
  INV_X1 U12592 ( .A(n10971), .ZN(n10085) );
  OAI21_X1 U12593 ( .B1(n9539), .B2(n10085), .A(n10082), .ZN(n10540) );
  XOR2_X1 U12594 ( .A(n10540), .B(n10090), .Z(n10083) );
  NOR2_X1 U12595 ( .A1(P1_REG2_REG_15__SCAN_IN), .A2(n10083), .ZN(n10541) );
  AOI21_X1 U12596 ( .B1(P1_REG2_REG_15__SCAN_IN), .B2(n10083), .A(n10541), 
        .ZN(n10095) );
  INV_X1 U12597 ( .A(n14508), .ZN(n10094) );
  AOI21_X1 U12598 ( .B1(n10773), .B2(n10085), .A(n10084), .ZN(n10546) );
  XNOR2_X1 U12599 ( .A(n10546), .B(n10977), .ZN(n10086) );
  NOR2_X1 U12600 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n10086), .ZN(n10547) );
  AOI21_X1 U12601 ( .B1(P1_REG1_REG_15__SCAN_IN), .B2(n10086), .A(n10547), 
        .ZN(n10087) );
  NOR2_X1 U12602 ( .A1(n10087), .A2(n13801), .ZN(n10092) );
  INV_X1 U12603 ( .A(P1_REG3_REG_15__SCAN_IN), .ZN(n13641) );
  NOR2_X1 U12604 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n13641), .ZN(n10088) );
  AOI21_X1 U12605 ( .B1(n14497), .B2(P1_ADDR_REG_15__SCAN_IN), .A(n10088), 
        .ZN(n10089) );
  OAI21_X1 U12606 ( .B1(n10090), .B2(n14501), .A(n10089), .ZN(n10091) );
  NOR2_X1 U12607 ( .A1(n10092), .A2(n10091), .ZN(n10093) );
  OAI21_X1 U12608 ( .B1(n10095), .B2(n10094), .A(n10093), .ZN(P1_U3258) );
  NAND2_X1 U12609 ( .A1(n12140), .A2(n12440), .ZN(n10096) );
  OAI21_X1 U12610 ( .B1(n7638), .B2(n12100), .A(n10096), .ZN(n10279) );
  NAND2_X1 U12611 ( .A1(n10279), .A2(n12104), .ZN(n10098) );
  OAI211_X1 U12612 ( .C1(n12095), .C2(n10327), .A(n10098), .B(n10097), .ZN(
        n10105) );
  OAI21_X1 U12613 ( .B1(n10101), .B2(n10100), .A(n10099), .ZN(n10103) );
  AOI21_X1 U12614 ( .B1(n10103), .B2(n10102), .A(n12115), .ZN(n10104) );
  AOI211_X1 U12615 ( .C1(n10382), .C2(n12112), .A(n10105), .B(n10104), .ZN(
        n10106) );
  INV_X1 U12616 ( .A(n10106), .ZN(P3_U3170) );
  INV_X1 U12617 ( .A(P3_REG0_REG_0__SCAN_IN), .ZN(n10107) );
  OAI22_X1 U12618 ( .A1(n12583), .A2(n10108), .B1(n15015), .B2(n10107), .ZN(
        n10109) );
  AOI21_X1 U12619 ( .B1(n10110), .B2(n15015), .A(n10109), .ZN(n10111) );
  INV_X1 U12620 ( .A(n10111), .ZN(P3_U3390) );
  AND2_X1 U12621 ( .A1(n10118), .A2(n10112), .ZN(n14895) );
  NAND2_X1 U12622 ( .A1(n14977), .A2(n14895), .ZN(n10640) );
  NAND2_X1 U12623 ( .A1(n14977), .A2(n14968), .ZN(n10113) );
  OAI21_X1 U12624 ( .B1(n10115), .B2(n10120), .A(n10114), .ZN(n10116) );
  INV_X1 U12625 ( .A(n10116), .ZN(n14988) );
  INV_X1 U12626 ( .A(P3_REG2_REG_2__SCAN_IN), .ZN(n10125) );
  NAND2_X1 U12627 ( .A1(n10117), .A2(n15016), .ZN(n14986) );
  NOR2_X1 U12628 ( .A1(n14986), .A2(n10118), .ZN(n10123) );
  XNOR2_X1 U12629 ( .A(n10119), .B(n10120), .ZN(n10122) );
  OAI21_X1 U12630 ( .B1(n10122), .B2(n14949), .A(n10121), .ZN(n14985) );
  AOI211_X1 U12631 ( .C1(n14973), .C2(P3_REG3_REG_2__SCAN_IN), .A(n10123), .B(
        n14985), .ZN(n10124) );
  MUX2_X1 U12632 ( .A(n10125), .B(n10124), .S(n14977), .Z(n10126) );
  OAI21_X1 U12633 ( .B1(n12486), .B2(n14988), .A(n10126), .ZN(P3_U3231) );
  NAND2_X1 U12634 ( .A1(n12810), .A2(n12812), .ZN(n10127) );
  NAND2_X1 U12635 ( .A1(n10128), .A2(n10127), .ZN(n10244) );
  NAND2_X1 U12636 ( .A1(n10678), .A2(n11860), .ZN(n10131) );
  AOI22_X1 U12637 ( .A1(n9097), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n9142), 
        .B2(n10129), .ZN(n10130) );
  OR2_X1 U12638 ( .A1(n12823), .A2(n13056), .ZN(n10250) );
  NAND2_X1 U12639 ( .A1(n12823), .A2(n13056), .ZN(n10252) );
  NAND2_X1 U12640 ( .A1(n10250), .A2(n10252), .ZN(n13006) );
  XNOR2_X1 U12641 ( .A(n10244), .B(n13006), .ZN(n10138) );
  NAND2_X1 U12642 ( .A1(n13057), .A2(n12710), .ZN(n10137) );
  NAND2_X1 U12643 ( .A1(n11701), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n10135) );
  XNOR2_X1 U12644 ( .A(n10257), .B(P2_REG3_REG_13__SCAN_IN), .ZN(n10574) );
  NAND2_X1 U12645 ( .A1(n9145), .A2(n10574), .ZN(n10134) );
  NAND2_X1 U12646 ( .A1(n11688), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10133) );
  NAND2_X1 U12647 ( .A1(n11123), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n10132) );
  NAND4_X1 U12648 ( .A1(n10135), .A2(n10134), .A3(n10133), .A4(n10132), .ZN(
        n13055) );
  NAND2_X1 U12649 ( .A1(n13055), .A2(n12711), .ZN(n10136) );
  NAND2_X1 U12650 ( .A1(n10137), .A2(n10136), .ZN(n10503) );
  AOI21_X1 U12651 ( .B1(n10138), .B2(n14740), .A(n10503), .ZN(n14372) );
  INV_X1 U12652 ( .A(n13006), .ZN(n10141) );
  XNOR2_X1 U12653 ( .A(n10253), .B(n10141), .ZN(n14370) );
  NAND2_X1 U12654 ( .A1(n12823), .A2(n10142), .ZN(n10143) );
  NAND2_X1 U12655 ( .A1(n10143), .A2(n14714), .ZN(n10144) );
  OR2_X1 U12656 ( .A1(n10254), .A2(n10144), .ZN(n14367) );
  AOI22_X1 U12657 ( .A1(n14731), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n10145), 
        .B2(n14719), .ZN(n10147) );
  NAND2_X1 U12658 ( .A1(n12823), .A2(n14341), .ZN(n10146) );
  OAI211_X1 U12659 ( .C1(n14367), .C2(n13282), .A(n10147), .B(n10146), .ZN(
        n10148) );
  AOI21_X1 U12660 ( .B1(n14370), .B2(n14727), .A(n10148), .ZN(n10149) );
  OAI21_X1 U12661 ( .B1(n14372), .B2(n14731), .A(n10149), .ZN(P2_U3253) );
  OAI21_X1 U12662 ( .B1(n10152), .B2(n10151), .A(n10150), .ZN(n14559) );
  INV_X1 U12663 ( .A(n14559), .ZN(n10158) );
  AOI22_X1 U12664 ( .A1(n14527), .A2(n6480), .B1(n13666), .B2(n14524), .ZN(
        n10157) );
  OAI21_X1 U12665 ( .B1(n10154), .B2(n11576), .A(n10153), .ZN(n10155) );
  NAND2_X1 U12666 ( .A1(n10155), .A2(n14392), .ZN(n10156) );
  OAI211_X1 U12667 ( .C1(n10158), .C2(n14023), .A(n10157), .B(n10156), .ZN(
        n14557) );
  AND2_X1 U12668 ( .A1(n14531), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n10163) );
  NAND2_X1 U12669 ( .A1(n14517), .A2(n10164), .ZN(n10159) );
  NAND2_X1 U12670 ( .A1(n10160), .A2(n10159), .ZN(n14556) );
  OAI22_X1 U12671 ( .A1(n13989), .A2(n14556), .B1(n10161), .B2(n14532), .ZN(
        n10162) );
  AOI211_X1 U12672 ( .C1(n14557), .C2(n13893), .A(n10163), .B(n10162), .ZN(
        n10166) );
  NAND2_X1 U12673 ( .A1(n11190), .A2(n11204), .ZN(n11539) );
  AOI22_X1 U12674 ( .A1(n14520), .A2(n14559), .B1(n14398), .B2(n10164), .ZN(
        n10165) );
  NAND2_X1 U12675 ( .A1(n10166), .A2(n10165), .ZN(P1_U3291) );
  INV_X1 U12676 ( .A(n10167), .ZN(n10168) );
  OR2_X1 U12677 ( .A1(n10172), .A2(n11490), .ZN(n10174) );
  AOI22_X1 U12678 ( .A1(n11548), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n11317), 
        .B2(n13747), .ZN(n10173) );
  NAND2_X1 U12679 ( .A1(n10174), .A2(n10173), .ZN(n14579) );
  INV_X1 U12680 ( .A(n14579), .ZN(n10322) );
  OAI22_X1 U12681 ( .A1(n10322), .A2(n13539), .B1(n10376), .B2(n13538), .ZN(
        n10413) );
  NAND2_X1 U12682 ( .A1(n14579), .A2(n13481), .ZN(n10176) );
  NAND2_X1 U12683 ( .A1(n13662), .A2(n13442), .ZN(n10175) );
  NAND2_X1 U12684 ( .A1(n10176), .A2(n10175), .ZN(n10177) );
  XNOR2_X1 U12685 ( .A(n10177), .B(n13536), .ZN(n10414) );
  XOR2_X1 U12686 ( .A(n10413), .B(n10414), .Z(n10416) );
  XOR2_X1 U12687 ( .A(n10417), .B(n10416), .Z(n10190) );
  INV_X1 U12688 ( .A(n13663), .ZN(n10221) );
  OAI22_X1 U12689 ( .A1(n13636), .A2(n10322), .B1(n13629), .B2(n10221), .ZN(
        n10189) );
  NAND2_X1 U12690 ( .A1(P1_U3086), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n13745) );
  NAND2_X1 U12691 ( .A1(n11503), .A2(P1_REG0_REG_8__SCAN_IN), .ZN(n10186) );
  OR2_X1 U12692 ( .A1(n6483), .A2(n10178), .ZN(n10185) );
  OR2_X1 U12693 ( .A1(n6487), .A2(n10179), .ZN(n10184) );
  NAND2_X1 U12694 ( .A1(n10181), .A2(n10180), .ZN(n10182) );
  NAND2_X1 U12695 ( .A1(n10209), .A2(n10182), .ZN(n10429) );
  OR2_X1 U12696 ( .A1(n11470), .A2(n10429), .ZN(n10183) );
  NAND4_X1 U12697 ( .A1(n10186), .A2(n10185), .A3(n10184), .A4(n10183), .ZN(
        n13661) );
  NAND2_X1 U12698 ( .A1(n13639), .A2(n13661), .ZN(n10187) );
  OAI211_X1 U12699 ( .C1(n13644), .C2(n10321), .A(n13745), .B(n10187), .ZN(
        n10188) );
  AOI211_X1 U12700 ( .C1(n10190), .C2(n13626), .A(n10189), .B(n10188), .ZN(
        n10191) );
  INV_X1 U12701 ( .A(n10191), .ZN(P1_U3213) );
  XNOR2_X1 U12702 ( .A(n13664), .B(n11233), .ZN(n11580) );
  OR2_X1 U12703 ( .A1(n13664), .A2(n11233), .ZN(n10194) );
  XNOR2_X1 U12704 ( .A(n11238), .B(n13663), .ZN(n11581) );
  NAND2_X1 U12705 ( .A1(n10284), .A2(n7037), .ZN(n10196) );
  OR2_X1 U12706 ( .A1(n11238), .A2(n13663), .ZN(n10195) );
  NAND2_X1 U12707 ( .A1(n10196), .A2(n10195), .ZN(n10312) );
  XNOR2_X1 U12708 ( .A(n14579), .B(n13662), .ZN(n11582) );
  NAND2_X1 U12709 ( .A1(n10312), .A2(n10313), .ZN(n10198) );
  OR2_X1 U12710 ( .A1(n14579), .A2(n13662), .ZN(n10197) );
  NAND2_X1 U12711 ( .A1(n10198), .A2(n10197), .ZN(n10368) );
  OR2_X1 U12712 ( .A1(n10199), .A2(n11490), .ZN(n10202) );
  AOI22_X1 U12713 ( .A1(n11548), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n11317), 
        .B2(n10200), .ZN(n10201) );
  NAND2_X1 U12714 ( .A1(n10202), .A2(n10201), .ZN(n11250) );
  INV_X1 U12715 ( .A(n13661), .ZN(n10224) );
  XNOR2_X1 U12716 ( .A(n11250), .B(n10224), .ZN(n11585) );
  NAND2_X1 U12717 ( .A1(n10368), .A2(n11585), .ZN(n10204) );
  OR2_X1 U12718 ( .A1(n11250), .A2(n13661), .ZN(n10203) );
  NAND2_X1 U12719 ( .A1(n10204), .A2(n10203), .ZN(n10453) );
  OR2_X1 U12720 ( .A1(n10205), .A2(n11490), .ZN(n10207) );
  AOI22_X1 U12721 ( .A1(n11548), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n11317), 
        .B2(n13769), .ZN(n10206) );
  NAND2_X1 U12722 ( .A1(n11503), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n10214) );
  OR2_X1 U12723 ( .A1(n6487), .A2(n10238), .ZN(n10213) );
  OR2_X1 U12724 ( .A1(n6483), .A2(n14625), .ZN(n10212) );
  AND2_X1 U12725 ( .A1(n10209), .A2(n10208), .ZN(n10210) );
  OR2_X1 U12726 ( .A1(n10210), .A2(n10228), .ZN(n10799) );
  OR2_X1 U12727 ( .A1(n11470), .A2(n10799), .ZN(n10211) );
  NAND4_X1 U12728 ( .A1(n10214), .A2(n10213), .A3(n10212), .A4(n10211), .ZN(
        n13660) );
  XNOR2_X1 U12729 ( .A(n11259), .B(n13660), .ZN(n11586) );
  INV_X1 U12730 ( .A(n11586), .ZN(n10452) );
  XNOR2_X1 U12731 ( .A(n10453), .B(n10452), .ZN(n14600) );
  NAND2_X1 U12732 ( .A1(n13665), .A2(n14561), .ZN(n10215) );
  OR2_X1 U12733 ( .A1(n13665), .A2(n14561), .ZN(n10217) );
  NAND2_X1 U12734 ( .A1(n10218), .A2(n10217), .ZN(n10299) );
  NAND2_X1 U12735 ( .A1(n10299), .A2(n11580), .ZN(n10220) );
  OR2_X1 U12736 ( .A1(n13664), .A2(n6874), .ZN(n10219) );
  NAND2_X1 U12737 ( .A1(n10220), .A2(n10219), .ZN(n10285) );
  NAND2_X1 U12738 ( .A1(n10221), .A2(n11238), .ZN(n10222) );
  AND2_X1 U12739 ( .A1(n14579), .A2(n10376), .ZN(n10223) );
  INV_X1 U12740 ( .A(n11585), .ZN(n10373) );
  NAND2_X1 U12741 ( .A1(n10225), .A2(n11586), .ZN(n10470) );
  OAI21_X1 U12742 ( .B1(n10225), .B2(n11586), .A(n10470), .ZN(n10226) );
  NAND2_X1 U12743 ( .A1(n10226), .A2(n14392), .ZN(n10235) );
  NAND2_X1 U12744 ( .A1(n11503), .A2(P1_REG0_REG_10__SCAN_IN), .ZN(n10233) );
  OR2_X1 U12745 ( .A1(n6487), .A2(n10227), .ZN(n10232) );
  NOR2_X1 U12746 ( .A1(n10228), .A2(P1_REG3_REG_10__SCAN_IN), .ZN(n10229) );
  OR2_X1 U12747 ( .A1(n10461), .A2(n10229), .ZN(n10849) );
  OR2_X1 U12748 ( .A1(n11470), .A2(n10849), .ZN(n10231) );
  OR2_X1 U12749 ( .A1(n6483), .A2(n14628), .ZN(n10230) );
  NAND4_X1 U12750 ( .A1(n10233), .A2(n10232), .A3(n10231), .A4(n10230), .ZN(
        n13659) );
  AOI22_X1 U12751 ( .A1(n14527), .A2(n13661), .B1(n13659), .B2(n14524), .ZN(
        n10234) );
  NAND2_X1 U12752 ( .A1(n10235), .A2(n10234), .ZN(n10236) );
  AOI21_X1 U12753 ( .B1(n14600), .B2(n14523), .A(n10236), .ZN(n14602) );
  INV_X1 U12754 ( .A(n11250), .ZN(n14589) );
  NAND2_X1 U12755 ( .A1(n10369), .A2(n11259), .ZN(n10237) );
  NAND2_X1 U12756 ( .A1(n10460), .A2(n10237), .ZN(n14597) );
  OAI22_X1 U12757 ( .A1(n13893), .A2(n10238), .B1(n10799), .B2(n14532), .ZN(
        n10239) );
  AOI21_X1 U12758 ( .B1(n14398), .B2(n11259), .A(n10239), .ZN(n10240) );
  OAI21_X1 U12759 ( .B1(n14597), .B2(n13989), .A(n10240), .ZN(n10241) );
  AOI21_X1 U12760 ( .B1(n14600), .B2(n14520), .A(n10241), .ZN(n10242) );
  OAI21_X1 U12761 ( .B1(n14602), .B2(n14388), .A(n10242), .ZN(P1_U3284) );
  INV_X1 U12762 ( .A(n13056), .ZN(n10245) );
  OR2_X1 U12763 ( .A1(n12823), .A2(n10245), .ZN(n10243) );
  NAND2_X1 U12764 ( .A1(n12823), .A2(n10245), .ZN(n10246) );
  NAND2_X1 U12765 ( .A1(n10765), .A2(n11860), .ZN(n10249) );
  INV_X1 U12766 ( .A(n10247), .ZN(n14690) );
  AOI22_X1 U12767 ( .A1(n9142), .A2(n14690), .B1(n11862), .B2(
        P1_DATAO_REG_13__SCAN_IN), .ZN(n10248) );
  XNOR2_X1 U12768 ( .A(n12830), .B(n14323), .ZN(n13009) );
  XNOR2_X1 U12769 ( .A(n10721), .B(n13009), .ZN(n10562) );
  INV_X1 U12770 ( .A(n10250), .ZN(n10251) );
  XOR2_X1 U12771 ( .A(n13009), .B(n10743), .Z(n10560) );
  OAI211_X1 U12772 ( .C1(n10741), .C2(n10254), .A(n14714), .B(n14346), .ZN(
        n10558) );
  NAND2_X1 U12773 ( .A1(P2_REG3_REG_13__SCAN_IN), .A2(P2_REG3_REG_14__SCAN_IN), 
        .ZN(n10255) );
  INV_X1 U12774 ( .A(n10733), .ZN(n10259) );
  INV_X1 U12775 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n10570) );
  INV_X1 U12776 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n10256) );
  OAI21_X1 U12777 ( .B1(n10257), .B2(n10570), .A(n10256), .ZN(n10258) );
  NAND2_X1 U12778 ( .A1(n10259), .A2(n10258), .ZN(n14339) );
  OR2_X1 U12779 ( .A1(n11663), .A2(n14339), .ZN(n10263) );
  NAND2_X1 U12780 ( .A1(n11701), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n10262) );
  NAND2_X1 U12781 ( .A1(n11688), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n10261) );
  NAND2_X1 U12782 ( .A1(n11123), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n10260) );
  NAND4_X1 U12783 ( .A1(n10263), .A2(n10262), .A3(n10261), .A4(n10260), .ZN(
        n13054) );
  NAND2_X1 U12784 ( .A1(n13054), .A2(n12711), .ZN(n10265) );
  NAND2_X1 U12785 ( .A1(n13056), .A2(n12710), .ZN(n10264) );
  AND2_X1 U12786 ( .A1(n10265), .A2(n10264), .ZN(n10571) );
  NAND2_X1 U12787 ( .A1(n14708), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n10267) );
  NAND2_X1 U12788 ( .A1(n14719), .A2(n10574), .ZN(n10266) );
  OAI211_X1 U12789 ( .C1(n14708), .C2(n10571), .A(n10267), .B(n10266), .ZN(
        n10268) );
  AOI21_X1 U12790 ( .B1(n12830), .B2(n14341), .A(n10268), .ZN(n10269) );
  OAI21_X1 U12791 ( .B1(n10558), .B2(n13282), .A(n10269), .ZN(n10270) );
  AOI21_X1 U12792 ( .B1(n10560), .B2(n14727), .A(n10270), .ZN(n10271) );
  OAI21_X1 U12793 ( .B1(n10562), .B2(n13198), .A(n10271), .ZN(P2_U3252) );
  INV_X1 U12794 ( .A(n14983), .ZN(n14989) );
  OAI21_X1 U12795 ( .B1(n10273), .B2(n10278), .A(n10272), .ZN(n10274) );
  INV_X1 U12796 ( .A(n10274), .ZN(n10386) );
  NOR2_X1 U12797 ( .A1(n10275), .A2(n14950), .ZN(n14948) );
  NOR2_X1 U12798 ( .A1(n14948), .A2(n10276), .ZN(n10277) );
  NOR2_X1 U12799 ( .A1(n10277), .A2(n10278), .ZN(n10355) );
  AOI211_X1 U12800 ( .C1(n10278), .C2(n10277), .A(n14949), .B(n10355), .ZN(
        n10280) );
  NOR2_X1 U12801 ( .A1(n10280), .A2(n10279), .ZN(n10380) );
  OAI21_X1 U12802 ( .B1(n14989), .B2(n10386), .A(n10380), .ZN(n10329) );
  INV_X1 U12803 ( .A(P3_REG1_REG_4__SCAN_IN), .ZN(n10281) );
  OAI22_X1 U12804 ( .A1(n12537), .A2(n10327), .B1(n15038), .B2(n10281), .ZN(
        n10282) );
  AOI21_X1 U12805 ( .B1(n10329), .B2(n15038), .A(n10282), .ZN(n10283) );
  INV_X1 U12806 ( .A(n10283), .ZN(P3_U3463) );
  XNOR2_X1 U12807 ( .A(n10284), .B(n7037), .ZN(n14578) );
  INV_X1 U12808 ( .A(n14578), .ZN(n10296) );
  INV_X1 U12809 ( .A(n14520), .ZN(n13901) );
  XNOR2_X1 U12810 ( .A(n10285), .B(n7037), .ZN(n10287) );
  AOI22_X1 U12811 ( .A1(n14527), .A2(n13664), .B1(n13662), .B2(n14524), .ZN(
        n10286) );
  OAI21_X1 U12812 ( .B1(n10287), .B2(n14542), .A(n10286), .ZN(n10288) );
  AOI21_X1 U12813 ( .B1(n14578), .B2(n14523), .A(n10288), .ZN(n14575) );
  MUX2_X1 U12814 ( .A(n10289), .B(n14575), .S(n13893), .Z(n10295) );
  INV_X1 U12815 ( .A(n10306), .ZN(n10291) );
  INV_X1 U12816 ( .A(n10290), .ZN(n10320) );
  OAI21_X1 U12817 ( .B1(n14573), .B2(n10291), .A(n10320), .ZN(n14574) );
  OAI22_X1 U12818 ( .A1(n14574), .A2(n13989), .B1(n10292), .B2(n14532), .ZN(
        n10293) );
  AOI21_X1 U12819 ( .B1(n14398), .B2(n11238), .A(n10293), .ZN(n10294) );
  OAI211_X1 U12820 ( .C1(n10296), .C2(n13901), .A(n10295), .B(n10294), .ZN(
        P1_U3287) );
  XNOR2_X1 U12821 ( .A(n10297), .B(n10298), .ZN(n14569) );
  INV_X1 U12822 ( .A(n14569), .ZN(n10311) );
  XNOR2_X1 U12823 ( .A(n10298), .B(n10299), .ZN(n10301) );
  AOI22_X1 U12824 ( .A1(n14527), .A2(n13665), .B1(n13663), .B2(n14524), .ZN(
        n10300) );
  OAI21_X1 U12825 ( .B1(n10301), .B2(n14542), .A(n10300), .ZN(n10302) );
  AOI21_X1 U12826 ( .B1(n14569), .B2(n14523), .A(n10302), .ZN(n14571) );
  MUX2_X1 U12827 ( .A(n10303), .B(n14571), .S(n13893), .Z(n10310) );
  NAND2_X1 U12828 ( .A1(n10304), .A2(n11233), .ZN(n10305) );
  NAND2_X1 U12829 ( .A1(n10306), .A2(n10305), .ZN(n14567) );
  OAI22_X1 U12830 ( .A1(n13989), .A2(n14567), .B1(n10307), .B2(n14532), .ZN(
        n10308) );
  AOI21_X1 U12831 ( .B1(n14398), .B2(n11233), .A(n10308), .ZN(n10309) );
  OAI211_X1 U12832 ( .C1(n10311), .C2(n13901), .A(n10310), .B(n10309), .ZN(
        P1_U3288) );
  XNOR2_X1 U12833 ( .A(n10312), .B(n10313), .ZN(n10318) );
  INV_X1 U12834 ( .A(n10318), .ZN(n14586) );
  XNOR2_X1 U12835 ( .A(n10314), .B(n10313), .ZN(n10316) );
  AOI22_X1 U12836 ( .A1(n14527), .A2(n13663), .B1(n13661), .B2(n14524), .ZN(
        n10315) );
  OAI21_X1 U12837 ( .B1(n10316), .B2(n14542), .A(n10315), .ZN(n10317) );
  AOI21_X1 U12838 ( .B1(n10318), .B2(n14523), .A(n10317), .ZN(n14584) );
  MUX2_X1 U12839 ( .A(n10319), .B(n14584), .S(n13893), .Z(n10325) );
  AOI21_X1 U12840 ( .B1(n14579), .B2(n10320), .A(n10370), .ZN(n14582) );
  OAI22_X1 U12841 ( .A1(n14534), .A2(n10322), .B1(n10321), .B2(n14532), .ZN(
        n10323) );
  AOI21_X1 U12842 ( .B1(n14582), .B2(n14519), .A(n10323), .ZN(n10324) );
  OAI211_X1 U12843 ( .C1(n14586), .C2(n13901), .A(n10325), .B(n10324), .ZN(
        P1_U3286) );
  INV_X1 U12844 ( .A(P3_REG0_REG_4__SCAN_IN), .ZN(n10326) );
  OAI22_X1 U12845 ( .A1(n12583), .A2(n10327), .B1(n15015), .B2(n10326), .ZN(
        n10328) );
  AOI21_X1 U12846 ( .B1(n10329), .B2(n15015), .A(n10328), .ZN(n10330) );
  INV_X1 U12847 ( .A(n10330), .ZN(P3_U3402) );
  AOI21_X1 U12848 ( .B1(n10333), .B2(n10332), .A(n10331), .ZN(n10349) );
  INV_X1 U12849 ( .A(n10334), .ZN(n10336) );
  AND2_X1 U12850 ( .A1(n10336), .A2(n10335), .ZN(n10337) );
  XNOR2_X1 U12851 ( .A(n10338), .B(n10337), .ZN(n10347) );
  NOR2_X1 U12852 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n7686), .ZN(n10339) );
  AOI21_X1 U12853 ( .B1(n14869), .B2(P3_ADDR_REG_9__SCAN_IN), .A(n10339), .ZN(
        n10340) );
  OAI21_X1 U12854 ( .B1(n14878), .B2(n10341), .A(n10340), .ZN(n10346) );
  AOI21_X1 U12855 ( .B1(n15034), .B2(n10343), .A(n10342), .ZN(n10344) );
  NOR2_X1 U12856 ( .A1(n10344), .A2(n14887), .ZN(n10345) );
  AOI211_X1 U12857 ( .C1(n14843), .C2(n10347), .A(n10346), .B(n10345), .ZN(
        n10348) );
  OAI21_X1 U12858 ( .B1(n10349), .B2(n14893), .A(n10348), .ZN(P3_U3191) );
  OAI21_X1 U12859 ( .B1(n10351), .B2(n10353), .A(n10350), .ZN(n14942) );
  INV_X1 U12860 ( .A(n10352), .ZN(n10354) );
  OAI21_X1 U12861 ( .B1(n10355), .B2(n10354), .A(n10353), .ZN(n10357) );
  AOI21_X1 U12862 ( .B1(n10357), .B2(n10356), .A(n14949), .ZN(n10359) );
  NOR2_X1 U12863 ( .A1(n10359), .A2(n10358), .ZN(n14945) );
  INV_X1 U12864 ( .A(n14945), .ZN(n10360) );
  AOI21_X1 U12865 ( .B1(n14983), .B2(n14942), .A(n10360), .ZN(n10367) );
  AOI22_X1 U12866 ( .A1(n10361), .A2(n14940), .B1(n15036), .B2(
        P3_REG1_REG_5__SCAN_IN), .ZN(n10362) );
  OAI21_X1 U12867 ( .B1(n10367), .B2(n15036), .A(n10362), .ZN(P3_U3464) );
  INV_X1 U12868 ( .A(P3_REG0_REG_5__SCAN_IN), .ZN(n10363) );
  OAI22_X1 U12869 ( .A1(n12583), .A2(n10364), .B1(n15015), .B2(n10363), .ZN(
        n10365) );
  INV_X1 U12870 ( .A(n10365), .ZN(n10366) );
  OAI21_X1 U12871 ( .B1(n10367), .B2(n8422), .A(n10366), .ZN(P3_U3405) );
  XNOR2_X1 U12872 ( .A(n10368), .B(n11585), .ZN(n14593) );
  OAI21_X1 U12873 ( .B1(n10370), .B2(n14589), .A(n10369), .ZN(n14590) );
  INV_X1 U12874 ( .A(n10429), .ZN(n10371) );
  INV_X1 U12875 ( .A(n14532), .ZN(n13996) );
  AOI22_X1 U12876 ( .A1(n14398), .A2(n11250), .B1(n10371), .B2(n13996), .ZN(
        n10372) );
  OAI21_X1 U12877 ( .B1(n14590), .B2(n13989), .A(n10372), .ZN(n10378) );
  INV_X1 U12878 ( .A(n13660), .ZN(n10792) );
  XNOR2_X1 U12879 ( .A(n10374), .B(n10373), .ZN(n10375) );
  OAI222_X1 U12880 ( .A1(n14008), .A2(n10792), .B1(n14006), .B2(n10376), .C1(
        n10375), .C2(n14542), .ZN(n14591) );
  MUX2_X1 U12881 ( .A(P1_REG2_REG_8__SCAN_IN), .B(n14591), .S(n13893), .Z(
        n10377) );
  AOI211_X1 U12882 ( .C1(n14383), .C2(n14593), .A(n10378), .B(n10377), .ZN(
        n10379) );
  INV_X1 U12883 ( .A(n10379), .ZN(P1_U3285) );
  INV_X1 U12884 ( .A(P3_REG2_REG_4__SCAN_IN), .ZN(n10381) );
  MUX2_X1 U12885 ( .A(n10381), .B(n10380), .S(n14977), .Z(n10385) );
  AOI22_X1 U12886 ( .A1(n14957), .A2(n10383), .B1(n14973), .B2(n10382), .ZN(
        n10384) );
  OAI211_X1 U12887 ( .C1(n12486), .C2(n10386), .A(n10385), .B(n10384), .ZN(
        P3_U3229) );
  INV_X1 U12888 ( .A(SI_23_), .ZN(n11075) );
  NAND2_X1 U12889 ( .A1(n10387), .A2(n12596), .ZN(n10389) );
  OAI211_X1 U12890 ( .C1(n11075), .C2(n12589), .A(n10389), .B(n10388), .ZN(
        P3_U3272) );
  XNOR2_X1 U12891 ( .A(n12810), .B(n11628), .ZN(n10394) );
  NAND2_X1 U12892 ( .A1(n13057), .A2(n11749), .ZN(n10395) );
  NAND2_X1 U12893 ( .A1(n10394), .A2(n10395), .ZN(n10495) );
  INV_X1 U12894 ( .A(n10394), .ZN(n10397) );
  INV_X1 U12895 ( .A(n10395), .ZN(n10396) );
  NAND2_X1 U12896 ( .A1(n10397), .A2(n10396), .ZN(n10398) );
  NAND2_X1 U12897 ( .A1(n10495), .A2(n10398), .ZN(n10402) );
  INV_X1 U12898 ( .A(n10403), .ZN(n10400) );
  INV_X1 U12899 ( .A(n10496), .ZN(n10401) );
  AOI21_X1 U12900 ( .B1(n10403), .B2(n10402), .A(n10401), .ZN(n10412) );
  INV_X1 U12901 ( .A(n10404), .ZN(n10409) );
  INV_X1 U12902 ( .A(n10405), .ZN(n10406) );
  AOI21_X1 U12903 ( .B1(n14330), .B2(n10407), .A(n10406), .ZN(n10408) );
  OAI21_X1 U12904 ( .B1(n10409), .B2(n14334), .A(n10408), .ZN(n10410) );
  AOI21_X1 U12905 ( .B1(n12810), .B2(n12703), .A(n10410), .ZN(n10411) );
  OAI21_X1 U12906 ( .B1(n10412), .B2(n12705), .A(n10411), .ZN(P2_U3208) );
  NAND2_X1 U12907 ( .A1(n11250), .A2(n13481), .ZN(n10419) );
  NAND2_X1 U12908 ( .A1(n13661), .A2(n13442), .ZN(n10418) );
  NAND2_X1 U12909 ( .A1(n10419), .A2(n10418), .ZN(n10420) );
  XNOR2_X1 U12910 ( .A(n10420), .B(n13536), .ZN(n10424) );
  NAND2_X1 U12911 ( .A1(n11250), .A2(n13442), .ZN(n10422) );
  NAND2_X1 U12912 ( .A1(n13485), .A2(n13661), .ZN(n10421) );
  NAND2_X1 U12913 ( .A1(n10422), .A2(n10421), .ZN(n10423) );
  NOR2_X1 U12914 ( .A1(n10424), .A2(n10423), .ZN(n10789) );
  AOI21_X1 U12915 ( .B1(n10424), .B2(n10423), .A(n10789), .ZN(n10425) );
  OAI21_X1 U12916 ( .B1(n10426), .B2(n10425), .A(n10791), .ZN(n10432) );
  NAND2_X1 U12917 ( .A1(n13620), .A2(n13662), .ZN(n10427) );
  OAI211_X1 U12918 ( .C1(n13617), .C2(n10792), .A(n10428), .B(n10427), .ZN(
        n10431) );
  OAI22_X1 U12919 ( .A1(n13636), .A2(n14589), .B1(n10429), .B2(n13644), .ZN(
        n10430) );
  AOI211_X1 U12920 ( .C1(n10432), .C2(n13626), .A(n10431), .B(n10430), .ZN(
        n10433) );
  INV_X1 U12921 ( .A(n10433), .ZN(P1_U3221) );
  INV_X1 U12922 ( .A(n10434), .ZN(n10435) );
  NAND2_X1 U12923 ( .A1(n7638), .A2(n10435), .ZN(n10509) );
  AND2_X1 U12924 ( .A1(n10511), .A2(n10509), .ZN(n12098) );
  XNOR2_X1 U12925 ( .A(n14996), .B(n11971), .ZN(n10506) );
  XNOR2_X1 U12926 ( .A(n12137), .B(n10506), .ZN(n12097) );
  NAND2_X1 U12927 ( .A1(n12098), .A2(n12097), .ZN(n12096) );
  INV_X1 U12928 ( .A(n10506), .ZN(n10436) );
  NAND2_X1 U12929 ( .A1(n10436), .A2(n12137), .ZN(n10512) );
  NAND2_X1 U12930 ( .A1(n12096), .A2(n10512), .ZN(n10646) );
  XNOR2_X1 U12931 ( .A(n14912), .B(n11971), .ZN(n10645) );
  XNOR2_X1 U12932 ( .A(n10646), .B(n10645), .ZN(n10442) );
  NAND2_X1 U12933 ( .A1(n12137), .A2(n12440), .ZN(n10437) );
  OAI21_X1 U12934 ( .B1(n10521), .B2(n12100), .A(n10437), .ZN(n14919) );
  INV_X1 U12935 ( .A(P3_REG3_REG_7__SCAN_IN), .ZN(n15176) );
  OAI22_X1 U12936 ( .A1(n12095), .A2(n10438), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15176), .ZN(n10440) );
  NOR2_X1 U12937 ( .A1(n14286), .A2(n14924), .ZN(n10439) );
  AOI211_X1 U12938 ( .C1(n12104), .C2(n14919), .A(n10440), .B(n10439), .ZN(
        n10441) );
  OAI21_X1 U12939 ( .B1(n10442), .B2(n12115), .A(n10441), .ZN(P3_U3153) );
  INV_X1 U12940 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10448) );
  AOI21_X1 U12941 ( .B1(n12810), .B2(n14788), .A(n10443), .ZN(n10444) );
  OAI211_X1 U12942 ( .C1(n10446), .C2(n14793), .A(n10445), .B(n10444), .ZN(
        n10449) );
  NAND2_X1 U12943 ( .A1(n10449), .A2(n14797), .ZN(n10447) );
  OAI21_X1 U12944 ( .B1(n14797), .B2(n10448), .A(n10447), .ZN(P2_U3463) );
  NAND2_X1 U12945 ( .A1(n10449), .A2(n6470), .ZN(n10450) );
  OAI21_X1 U12946 ( .B1(n6470), .B2(n10451), .A(n10450), .ZN(P2_U3510) );
  NAND2_X1 U12947 ( .A1(n10453), .A2(n10452), .ZN(n10455) );
  OR2_X1 U12948 ( .A1(n11259), .A2(n13660), .ZN(n10454) );
  NAND2_X1 U12949 ( .A1(n10456), .A2(n11547), .ZN(n10459) );
  AOI22_X1 U12950 ( .A1(n11548), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n11317), 
        .B2(n10457), .ZN(n10458) );
  XNOR2_X1 U12951 ( .A(n11268), .B(n13659), .ZN(n11587) );
  XNOR2_X1 U12952 ( .A(n10620), .B(n10619), .ZN(n14610) );
  INV_X1 U12953 ( .A(n14610), .ZN(n10477) );
  AOI21_X1 U12954 ( .B1(n10460), .B2(n11268), .A(n14596), .ZN(n10468) );
  NAND2_X1 U12955 ( .A1(n6482), .A2(P1_REG2_REG_11__SCAN_IN), .ZN(n10467) );
  OR2_X1 U12956 ( .A1(n6483), .A2(n14446), .ZN(n10466) );
  OR2_X1 U12957 ( .A1(n10461), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n10462) );
  NAND2_X1 U12958 ( .A1(n10606), .A2(n10462), .ZN(n10893) );
  OR2_X1 U12959 ( .A1(n11470), .A2(n10893), .ZN(n10465) );
  INV_X1 U12960 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n10463) );
  OR2_X1 U12961 ( .A1(n11516), .A2(n10463), .ZN(n10464) );
  NAND4_X1 U12962 ( .A1(n10467), .A2(n10466), .A3(n10465), .A4(n10464), .ZN(
        n13658) );
  AOI22_X1 U12963 ( .A1(n10468), .A2(n10623), .B1(n14524), .B2(n13658), .ZN(
        n14604) );
  NAND2_X1 U12964 ( .A1(n11259), .A2(n10792), .ZN(n10469) );
  AOI21_X1 U12965 ( .B1(n10471), .B2(n10619), .A(n14542), .ZN(n10472) );
  AOI22_X1 U12966 ( .A1(n10472), .A2(n10614), .B1(n14527), .B2(n13660), .ZN(
        n14605) );
  OAI21_X1 U12967 ( .B1(n11204), .B2(n14604), .A(n14605), .ZN(n10475) );
  INV_X1 U12968 ( .A(n11268), .ZN(n14607) );
  NOR2_X1 U12969 ( .A1(n14607), .A2(n14534), .ZN(n10474) );
  OAI22_X1 U12970 ( .A1(n13893), .A2(n10227), .B1(n10849), .B2(n14532), .ZN(
        n10473) );
  AOI211_X1 U12971 ( .C1(n10475), .C2(n13893), .A(n10474), .B(n10473), .ZN(
        n10476) );
  OAI21_X1 U12972 ( .B1(n14015), .B2(n10477), .A(n10476), .ZN(P1_U3283) );
  OAI21_X1 U12973 ( .B1(n10002), .B2(n10479), .A(n10478), .ZN(n10595) );
  XOR2_X1 U12974 ( .A(n10730), .B(n10595), .Z(n10480) );
  NAND2_X1 U12975 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n10480), .ZN(n10596) );
  OAI21_X1 U12976 ( .B1(P2_REG1_REG_15__SCAN_IN), .B2(n10480), .A(n10596), 
        .ZN(n10489) );
  NAND2_X1 U12977 ( .A1(n10725), .A2(n10481), .ZN(n10483) );
  NAND2_X1 U12978 ( .A1(P2_REG2_REG_15__SCAN_IN), .A2(n10484), .ZN(n10591) );
  OAI211_X1 U12979 ( .C1(n10484), .C2(P2_REG2_REG_15__SCAN_IN), .A(n14692), 
        .B(n10591), .ZN(n10488) );
  INV_X1 U12980 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n10485) );
  INV_X1 U12981 ( .A(P2_ADDR_REG_15__SCAN_IN), .ZN(n14228) );
  OAI22_X1 U12982 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10485), .B1(n14671), .B2(
        n14228), .ZN(n10486) );
  AOI21_X1 U12983 ( .B1(n14691), .B2(n10730), .A(n10486), .ZN(n10487) );
  OAI211_X1 U12984 ( .C1(n10489), .C2(n14639), .A(n10488), .B(n10487), .ZN(
        P2_U3229) );
  INV_X1 U12985 ( .A(n12823), .ZN(n14368) );
  XNOR2_X1 U12986 ( .A(n12823), .B(n11628), .ZN(n10490) );
  NAND2_X1 U12987 ( .A1(n13056), .A2(n11749), .ZN(n10491) );
  NAND2_X1 U12988 ( .A1(n10490), .A2(n10491), .ZN(n10568) );
  INV_X1 U12989 ( .A(n10490), .ZN(n10493) );
  INV_X1 U12990 ( .A(n10491), .ZN(n10492) );
  NAND2_X1 U12991 ( .A1(n10493), .A2(n10492), .ZN(n10494) );
  AND2_X1 U12992 ( .A1(n10568), .A2(n10494), .ZN(n10498) );
  OAI21_X1 U12993 ( .B1(n10498), .B2(n10497), .A(n10569), .ZN(n10499) );
  NAND2_X1 U12994 ( .A1(n10499), .A2(n14328), .ZN(n10505) );
  NOR2_X1 U12995 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10500), .ZN(n13122) );
  NOR2_X1 U12996 ( .A1(n14334), .A2(n10501), .ZN(n10502) );
  AOI211_X1 U12997 ( .C1(n14330), .C2(n10503), .A(n13122), .B(n10502), .ZN(
        n10504) );
  OAI211_X1 U12998 ( .C1(n14368), .C2(n12719), .A(n10505), .B(n10504), .ZN(
        P2_U3196) );
  XNOR2_X1 U12999 ( .A(n10811), .B(n11971), .ZN(n10577) );
  XNOR2_X1 U13000 ( .A(n10577), .B(n12134), .ZN(n10658) );
  XNOR2_X1 U13001 ( .A(n10649), .B(n6508), .ZN(n10515) );
  XNOR2_X1 U13002 ( .A(n10521), .B(n10515), .ZN(n10647) );
  NAND2_X1 U13003 ( .A1(n10507), .A2(n10506), .ZN(n10508) );
  AND4_X1 U13004 ( .A1(n10645), .A2(n10647), .A3(n10509), .A4(n10508), .ZN(
        n10510) );
  NAND2_X1 U13005 ( .A1(n10511), .A2(n10510), .ZN(n10519) );
  INV_X1 U13006 ( .A(n10647), .ZN(n10514) );
  OAI21_X1 U13007 ( .B1(n10514), .B2(n10512), .A(n10645), .ZN(n10517) );
  INV_X1 U13008 ( .A(n10645), .ZN(n10513) );
  OAI21_X1 U13009 ( .B1(n12101), .B2(n10514), .A(n10513), .ZN(n10516) );
  AOI22_X1 U13010 ( .A1(n10517), .A2(n10516), .B1(n10515), .B2(n12135), .ZN(
        n10518) );
  OR2_X1 U13011 ( .A1(n10662), .A2(n10658), .ZN(n10582) );
  INV_X1 U13012 ( .A(n10582), .ZN(n10520) );
  AOI21_X1 U13013 ( .B1(n10658), .B2(n10662), .A(n10520), .ZN(n10528) );
  OR2_X1 U13014 ( .A1(n10580), .A2(n12100), .ZN(n10523) );
  OR2_X1 U13015 ( .A1(n10521), .A2(n12103), .ZN(n10522) );
  AND2_X1 U13016 ( .A1(n10523), .A2(n10522), .ZN(n10809) );
  AOI22_X1 U13017 ( .A1(n14274), .A2(n10524), .B1(P3_REG3_REG_9__SCAN_IN), 
        .B2(P3_U3151), .ZN(n10525) );
  OAI21_X1 U13018 ( .B1(n10809), .B2(n14281), .A(n10525), .ZN(n10526) );
  AOI21_X1 U13019 ( .B1(n10812), .B2(n12112), .A(n10526), .ZN(n10527) );
  OAI21_X1 U13020 ( .B1(n10528), .B2(n12115), .A(n10527), .ZN(P3_U3171) );
  INV_X1 U13021 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n10539) );
  INV_X1 U13022 ( .A(n10529), .ZN(n10530) );
  NAND2_X1 U13023 ( .A1(n10534), .A2(n10533), .ZN(n10535) );
  INV_X1 U13024 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n10557) );
  MUX2_X1 U13025 ( .A(n10539), .B(n10557), .S(n11543), .Z(n10536) );
  NAND2_X1 U13026 ( .A1(n10537), .A2(n10536), .ZN(n10538) );
  AND2_X1 U13027 ( .A1(n10701), .A2(n10538), .ZN(n11639) );
  INV_X1 U13028 ( .A(n11639), .ZN(n10556) );
  OAI222_X1 U13029 ( .A1(n14124), .A2(n10539), .B1(n14119), .B2(n10556), .C1(
        n11206), .C2(P1_U3086), .ZN(P1_U3335) );
  NOR2_X1 U13030 ( .A1(n10977), .A2(n10540), .ZN(n10542) );
  NOR2_X1 U13031 ( .A1(n10542), .A2(n10541), .ZN(n10545) );
  INV_X1 U13032 ( .A(P1_REG2_REG_16__SCAN_IN), .ZN(n11110) );
  NOR2_X1 U13033 ( .A1(n10714), .A2(n11110), .ZN(n10543) );
  AOI21_X1 U13034 ( .B1(n11110), .B2(n10714), .A(n10543), .ZN(n10544) );
  NAND2_X1 U13035 ( .A1(n10544), .A2(n10545), .ZN(n10710) );
  OAI211_X1 U13036 ( .C1(n10545), .C2(n10544), .A(n14508), .B(n10710), .ZN(
        n10555) );
  NAND2_X1 U13037 ( .A1(P1_U3086), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n13572)
         );
  NOR2_X1 U13038 ( .A1(n10977), .A2(n10546), .ZN(n10548) );
  NOR2_X1 U13039 ( .A1(n10548), .A2(n10547), .ZN(n10551) );
  INV_X1 U13040 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n14417) );
  NOR2_X1 U13041 ( .A1(n14417), .A2(n10714), .ZN(n10549) );
  AOI21_X1 U13042 ( .B1(n14417), .B2(n10714), .A(n10549), .ZN(n10550) );
  NAND2_X1 U13043 ( .A1(n10550), .A2(n10551), .ZN(n10713) );
  OAI211_X1 U13044 ( .C1(n10551), .C2(n10550), .A(n14504), .B(n10713), .ZN(
        n10552) );
  NAND2_X1 U13045 ( .A1(n13572), .A2(n10552), .ZN(n10553) );
  AOI21_X1 U13046 ( .B1(n14497), .B2(P1_ADDR_REG_16__SCAN_IN), .A(n10553), 
        .ZN(n10554) );
  OAI211_X1 U13047 ( .C1(n14501), .C2(n10714), .A(n10555), .B(n10554), .ZN(
        P1_U3259) );
  OAI222_X1 U13048 ( .A1(n13440), .A2(n10557), .B1(P2_U3088), .B2(n8952), .C1(
        n13438), .C2(n10556), .ZN(P2_U3307) );
  OAI211_X1 U13049 ( .C1(n10741), .C2(n14774), .A(n10558), .B(n10571), .ZN(
        n10559) );
  AOI21_X1 U13050 ( .B1(n10560), .B2(n14768), .A(n10559), .ZN(n10561) );
  OAI21_X1 U13051 ( .B1(n14352), .B2(n10562), .A(n10561), .ZN(n10565) );
  NAND2_X1 U13052 ( .A1(n10565), .A2(n6470), .ZN(n10563) );
  OAI21_X1 U13053 ( .B1(n6470), .B2(n10564), .A(n10563), .ZN(P2_U3512) );
  INV_X1 U13054 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10567) );
  NAND2_X1 U13055 ( .A1(n10565), .A2(n14797), .ZN(n10566) );
  OAI21_X1 U13056 ( .B1(n14797), .B2(n10567), .A(n10566), .ZN(P2_U3469) );
  XNOR2_X1 U13057 ( .A(n12830), .B(n11628), .ZN(n11007) );
  NAND2_X1 U13058 ( .A1(n13055), .A2(n11749), .ZN(n11008) );
  XNOR2_X1 U13059 ( .A(n11007), .B(n11008), .ZN(n11006) );
  XNOR2_X1 U13060 ( .A(n11012), .B(n11006), .ZN(n10576) );
  OAI22_X1 U13061 ( .A1(n12715), .A2(n10571), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10570), .ZN(n10573) );
  NOR2_X1 U13062 ( .A1(n10741), .A2(n12719), .ZN(n10572) );
  AOI211_X1 U13063 ( .C1(n12717), .C2(n10574), .A(n10573), .B(n10572), .ZN(
        n10575) );
  OAI21_X1 U13064 ( .B1(n10576), .B2(n12705), .A(n10575), .ZN(P2_U3206) );
  INV_X1 U13065 ( .A(n10577), .ZN(n10578) );
  NAND2_X1 U13066 ( .A1(n10579), .A2(n10578), .ZN(n10581) );
  AND2_X1 U13067 ( .A1(n10582), .A2(n10581), .ZN(n10585) );
  XNOR2_X1 U13068 ( .A(n14905), .B(n11971), .ZN(n10657) );
  XNOR2_X1 U13069 ( .A(n10580), .B(n10657), .ZN(n10584) );
  AND2_X1 U13070 ( .A1(n10584), .A2(n10581), .ZN(n10659) );
  NAND2_X1 U13071 ( .A1(n10582), .A2(n10659), .ZN(n10583) );
  OAI211_X1 U13072 ( .C1(n10585), .C2(n10584), .A(n14276), .B(n10583), .ZN(
        n10589) );
  NAND2_X1 U13073 ( .A1(n12134), .A2(n12440), .ZN(n10586) );
  OAI21_X1 U13074 ( .B1(n10861), .B2(n12100), .A(n10586), .ZN(n14901) );
  NAND2_X1 U13075 ( .A1(P3_U3151), .A2(P3_REG3_REG_10__SCAN_IN), .ZN(n14860)
         );
  OAI21_X1 U13076 ( .B1(n12095), .B2(n14905), .A(n14860), .ZN(n10587) );
  AOI21_X1 U13077 ( .B1(n12104), .B2(n14901), .A(n10587), .ZN(n10588) );
  OAI211_X1 U13078 ( .C1(n14910), .C2(n14286), .A(n10589), .B(n10588), .ZN(
        P3_U3157) );
  INV_X1 U13079 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n10818) );
  AOI22_X1 U13080 ( .A1(n10928), .A2(P2_REG2_REG_16__SCAN_IN), .B1(n10818), 
        .B2(n10822), .ZN(n10594) );
  NAND2_X1 U13081 ( .A1(n10730), .A2(n10590), .ZN(n10592) );
  NAND2_X1 U13082 ( .A1(n10592), .A2(n10591), .ZN(n10593) );
  OAI21_X1 U13083 ( .B1(n10594), .B2(n10593), .A(n10817), .ZN(n10604) );
  NAND2_X1 U13084 ( .A1(P2_U3088), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n12656)
         );
  OAI21_X1 U13085 ( .B1(n14667), .B2(n10822), .A(n12656), .ZN(n10602) );
  INV_X1 U13086 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n10823) );
  AOI22_X1 U13087 ( .A1(n10928), .A2(P2_REG1_REG_16__SCAN_IN), .B1(n10823), 
        .B2(n10822), .ZN(n10599) );
  NAND2_X1 U13088 ( .A1(n10730), .A2(n10595), .ZN(n10597) );
  NAND2_X1 U13089 ( .A1(n10597), .A2(n10596), .ZN(n10598) );
  NAND2_X1 U13090 ( .A1(n10599), .A2(n10598), .ZN(n10821) );
  OAI21_X1 U13091 ( .B1(n10599), .B2(n10598), .A(n10821), .ZN(n10600) );
  NOR2_X1 U13092 ( .A1(n10600), .A2(n14639), .ZN(n10601) );
  AOI211_X1 U13093 ( .C1(n14685), .C2(P2_ADDR_REG_16__SCAN_IN), .A(n10602), 
        .B(n10601), .ZN(n10603) );
  OAI21_X1 U13094 ( .B1(n10604), .B2(n14677), .A(n10603), .ZN(P2_U3230) );
  NAND2_X1 U13095 ( .A1(n11503), .A2(P1_REG0_REG_12__SCAN_IN), .ZN(n10612) );
  NAND2_X1 U13096 ( .A1(n10606), .A2(n10605), .ZN(n10607) );
  NAND2_X1 U13097 ( .A1(n10685), .A2(n10607), .ZN(n10911) );
  OR2_X1 U13098 ( .A1(n11470), .A2(n10911), .ZN(n10611) );
  OR2_X1 U13099 ( .A1(n6487), .A2(n9535), .ZN(n10610) );
  OR2_X1 U13100 ( .A1(n6483), .A2(n10608), .ZN(n10609) );
  NAND4_X1 U13101 ( .A1(n10612), .A2(n10611), .A3(n10610), .A4(n10609), .ZN(
        n13657) );
  INV_X1 U13102 ( .A(n13659), .ZN(n10842) );
  OR2_X1 U13103 ( .A1(n11268), .A2(n10842), .ZN(n10613) );
  NAND2_X1 U13104 ( .A1(n10615), .A2(n11547), .ZN(n10617) );
  AOI22_X1 U13105 ( .A1(n11548), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n11317), 
        .B2(n13783), .ZN(n10616) );
  XNOR2_X1 U13106 ( .A(n11273), .B(n13658), .ZN(n11589) );
  XNOR2_X1 U13107 ( .A(n10681), .B(n11589), .ZN(n10618) );
  OAI222_X1 U13108 ( .A1(n14008), .A2(n11285), .B1(n14006), .B2(n10842), .C1(
        n10618), .C2(n14542), .ZN(n14443) );
  INV_X1 U13109 ( .A(n14443), .ZN(n10630) );
  NAND2_X1 U13110 ( .A1(n10620), .A2(n10619), .ZN(n10622) );
  OR2_X1 U13111 ( .A1(n11268), .A2(n13659), .ZN(n10621) );
  NAND2_X1 U13112 ( .A1(n10622), .A2(n10621), .ZN(n10675) );
  INV_X1 U13113 ( .A(n11589), .ZN(n10674) );
  XNOR2_X1 U13114 ( .A(n10675), .B(n10674), .ZN(n14445) );
  AND2_X1 U13115 ( .A1(n10623), .A2(n11273), .ZN(n10624) );
  OR2_X1 U13116 ( .A1(n10624), .A2(n10694), .ZN(n14442) );
  OAI22_X1 U13117 ( .A1(n13893), .A2(n10625), .B1(n10893), .B2(n14532), .ZN(
        n10626) );
  AOI21_X1 U13118 ( .B1(n11273), .B2(n14398), .A(n10626), .ZN(n10627) );
  OAI21_X1 U13119 ( .B1(n14442), .B2(n13989), .A(n10627), .ZN(n10628) );
  AOI21_X1 U13120 ( .B1(n14445), .B2(n14383), .A(n10628), .ZN(n10629) );
  OAI21_X1 U13121 ( .B1(n10630), .B2(n14388), .A(n10629), .ZN(P1_U3282) );
  XNOR2_X1 U13122 ( .A(n10631), .B(n10632), .ZN(n15007) );
  NAND2_X1 U13123 ( .A1(n15007), .A2(n14968), .ZN(n10639) );
  NAND2_X1 U13124 ( .A1(n10633), .A2(n10632), .ZN(n10634) );
  NAND2_X1 U13125 ( .A1(n10635), .A2(n10634), .ZN(n10637) );
  NAND2_X1 U13126 ( .A1(n12134), .A2(n12437), .ZN(n10636) );
  OAI21_X1 U13127 ( .B1(n12101), .B2(n12103), .A(n10636), .ZN(n10652) );
  AOI21_X1 U13128 ( .B1(n10637), .B2(n14961), .A(n10652), .ZN(n10638) );
  INV_X1 U13129 ( .A(n10640), .ZN(n14974) );
  INV_X1 U13130 ( .A(P3_REG2_REG_8__SCAN_IN), .ZN(n10642) );
  AND2_X1 U13131 ( .A1(n10649), .A2(n15016), .ZN(n15006) );
  AOI22_X1 U13132 ( .A1(n12479), .A2(n15006), .B1(n14973), .B2(n10653), .ZN(
        n10641) );
  OAI21_X1 U13133 ( .B1(n10642), .B2(n14977), .A(n10641), .ZN(n10643) );
  AOI21_X1 U13134 ( .B1(n15007), .B2(n14974), .A(n10643), .ZN(n10644) );
  OAI21_X1 U13135 ( .B1(n15009), .B2(n14979), .A(n10644), .ZN(P3_U3225) );
  MUX2_X1 U13136 ( .A(n12136), .B(n10646), .S(n10645), .Z(n10648) );
  XNOR2_X1 U13137 ( .A(n10648), .B(n10647), .ZN(n10656) );
  NAND2_X1 U13138 ( .A1(n14274), .A2(n10649), .ZN(n10650) );
  OAI21_X1 U13139 ( .B1(P3_STATE_REG_SCAN_IN), .B2(n15058), .A(n10650), .ZN(
        n10651) );
  AOI21_X1 U13140 ( .B1(n10652), .B2(n12104), .A(n10651), .ZN(n10655) );
  NAND2_X1 U13141 ( .A1(n12112), .A2(n10653), .ZN(n10654) );
  OAI211_X1 U13142 ( .C1(n10656), .C2(n12115), .A(n10655), .B(n10654), .ZN(
        P3_U3161) );
  AND2_X1 U13143 ( .A1(n12133), .A2(n10657), .ZN(n10660) );
  XNOR2_X1 U13144 ( .A(n10918), .B(n6508), .ZN(n10859) );
  INV_X1 U13145 ( .A(n10859), .ZN(n10664) );
  XNOR2_X1 U13146 ( .A(n10663), .B(n6508), .ZN(n10863) );
  OAI22_X1 U13147 ( .A1(n12132), .A2(n10664), .B1(n10863), .B2(n12131), .ZN(
        n10668) );
  NOR2_X1 U13148 ( .A1(n10861), .A2(n10859), .ZN(n10665) );
  NAND2_X1 U13149 ( .A1(n10665), .A2(n12131), .ZN(n10667) );
  OAI21_X1 U13150 ( .B1(n10665), .B2(n12131), .A(n10863), .ZN(n10666) );
  XNOR2_X1 U13151 ( .A(n14299), .B(n11971), .ZN(n10871) );
  XNOR2_X1 U13152 ( .A(n10871), .B(n10873), .ZN(n10669) );
  XNOR2_X1 U13153 ( .A(n10870), .B(n10669), .ZN(n10673) );
  AOI22_X1 U13154 ( .A1(n12440), .A2(n12131), .B1(n12439), .B2(n12437), .ZN(
        n12466) );
  NAND2_X1 U13155 ( .A1(P3_U3151), .A2(P3_REG3_REG_13__SCAN_IN), .ZN(n12171)
         );
  OAI21_X1 U13156 ( .B1(n12466), .B2(n14281), .A(n12171), .ZN(n10671) );
  NOR2_X1 U13157 ( .A1(n14299), .A2(n12095), .ZN(n10670) );
  AOI211_X1 U13158 ( .C1(n12468), .C2(n12112), .A(n10671), .B(n10670), .ZN(
        n10672) );
  OAI21_X1 U13159 ( .B1(n10673), .B2(n12115), .A(n10672), .ZN(P3_U3174) );
  NAND2_X1 U13160 ( .A1(n10675), .A2(n10674), .ZN(n10677) );
  OR2_X1 U13161 ( .A1(n11273), .A2(n13658), .ZN(n10676) );
  NAND2_X1 U13162 ( .A1(n10678), .A2(n11547), .ZN(n10680) );
  AOI22_X1 U13163 ( .A1(n11548), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n14491), 
        .B2(n11317), .ZN(n10679) );
  NAND2_X1 U13164 ( .A1(n10680), .A2(n10679), .ZN(n11281) );
  XNOR2_X1 U13165 ( .A(n11281), .B(n11285), .ZN(n11592) );
  XNOR2_X1 U13166 ( .A(n10769), .B(n11592), .ZN(n14263) );
  INV_X1 U13167 ( .A(n13658), .ZN(n10882) );
  OR2_X1 U13168 ( .A1(n11273), .A2(n10882), .ZN(n10682) );
  INV_X1 U13169 ( .A(n11592), .ZN(n10762) );
  XNOR2_X1 U13170 ( .A(n10763), .B(n10762), .ZN(n10692) );
  NAND2_X1 U13171 ( .A1(n11503), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n10690) );
  OR2_X1 U13172 ( .A1(n6483), .A2(n14440), .ZN(n10689) );
  OR2_X1 U13173 ( .A1(n6487), .A2(n9530), .ZN(n10688) );
  NAND2_X1 U13174 ( .A1(n10685), .A2(n10684), .ZN(n10686) );
  NAND2_X1 U13175 ( .A1(n10775), .A2(n10686), .ZN(n11055) );
  OR2_X1 U13176 ( .A1(n11470), .A2(n11055), .ZN(n10687) );
  NAND4_X1 U13177 ( .A1(n10690), .A2(n10689), .A3(n10688), .A4(n10687), .ZN(
        n14394) );
  AOI22_X1 U13178 ( .A1(n14527), .A2(n13658), .B1(n14394), .B2(n14524), .ZN(
        n10691) );
  OAI21_X1 U13179 ( .B1(n10692), .B2(n14542), .A(n10691), .ZN(n10693) );
  AOI21_X1 U13180 ( .B1(n14263), .B2(n14523), .A(n10693), .ZN(n14265) );
  INV_X1 U13181 ( .A(n11281), .ZN(n14260) );
  NAND2_X1 U13182 ( .A1(n10694), .A2(n14260), .ZN(n10771) );
  OR2_X1 U13183 ( .A1(n10694), .A2(n14260), .ZN(n10695) );
  NAND2_X1 U13184 ( .A1(n10771), .A2(n10695), .ZN(n14261) );
  OAI22_X1 U13185 ( .A1(n13893), .A2(n9535), .B1(n10911), .B2(n14532), .ZN(
        n10696) );
  AOI21_X1 U13186 ( .B1(n11281), .B2(n14398), .A(n10696), .ZN(n10697) );
  OAI21_X1 U13187 ( .B1(n14261), .B2(n13989), .A(n10697), .ZN(n10698) );
  AOI21_X1 U13188 ( .B1(n14263), .B2(n14520), .A(n10698), .ZN(n10699) );
  OAI21_X1 U13189 ( .B1(n14265), .B2(n14388), .A(n10699), .ZN(P1_U3281) );
  MUX2_X1 U13190 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(P1_DATAO_REG_21__SCAN_IN), 
        .S(n11543), .Z(n10702) );
  NAND2_X1 U13191 ( .A1(n10702), .A2(SI_21_), .ZN(n10960) );
  OAI21_X1 U13192 ( .B1(SI_21_), .B2(n10702), .A(n10960), .ZN(n10705) );
  INV_X1 U13193 ( .A(n10705), .ZN(n10703) );
  INV_X1 U13194 ( .A(n10704), .ZN(n10706) );
  NAND2_X1 U13195 ( .A1(n10706), .A2(n10705), .ZN(n10707) );
  AND2_X1 U13196 ( .A1(n10961), .A2(n10707), .ZN(n11646) );
  INV_X1 U13197 ( .A(n11646), .ZN(n10760) );
  OAI222_X1 U13198 ( .A1(n14124), .A2(n10708), .B1(n14130), .B2(n10760), .C1(
        n7146), .C2(P1_U3086), .ZN(P1_U3334) );
  INV_X1 U13199 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n10950) );
  NOR2_X1 U13200 ( .A1(n10953), .A2(n10950), .ZN(n10709) );
  AOI21_X1 U13201 ( .B1(n10950), .B2(n10953), .A(n10709), .ZN(n10712) );
  OAI21_X1 U13202 ( .B1(n10714), .B2(n11110), .A(n10710), .ZN(n10711) );
  NAND2_X1 U13203 ( .A1(n10712), .A2(n10711), .ZN(n10949) );
  OAI211_X1 U13204 ( .C1(n10712), .C2(n10711), .A(n14508), .B(n10949), .ZN(
        n10720) );
  NAND2_X1 U13205 ( .A1(P1_U3086), .A2(P1_REG3_REG_17__SCAN_IN), .ZN(n13585)
         );
  INV_X1 U13206 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n11103) );
  INV_X1 U13207 ( .A(n10953), .ZN(n11306) );
  MUX2_X1 U13208 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n11103), .S(n11306), .Z(
        n10716) );
  OAI21_X1 U13209 ( .B1(n14417), .B2(n10714), .A(n10713), .ZN(n10715) );
  NAND2_X1 U13210 ( .A1(n10716), .A2(n10715), .ZN(n10952) );
  OAI211_X1 U13211 ( .C1(n10716), .C2(n10715), .A(n10952), .B(n14504), .ZN(
        n10717) );
  NAND2_X1 U13212 ( .A1(n13585), .A2(n10717), .ZN(n10718) );
  AOI21_X1 U13213 ( .B1(n14497), .B2(P1_ADDR_REG_17__SCAN_IN), .A(n10718), 
        .ZN(n10719) );
  OAI211_X1 U13214 ( .C1(n14501), .C2(n10953), .A(n10720), .B(n10719), .ZN(
        P1_U3260) );
  AND2_X1 U13215 ( .A1(n12830), .A2(n14323), .ZN(n10722) );
  OR2_X1 U13216 ( .A1(n12830), .A2(n14323), .ZN(n10723) );
  NAND2_X1 U13217 ( .A1(n10970), .A2(n12943), .ZN(n10727) );
  AOI22_X1 U13218 ( .A1(n10725), .A2(n9142), .B1(n11862), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n10726) );
  NAND2_X2 U13219 ( .A1(n10727), .A2(n10726), .ZN(n14342) );
  INV_X1 U13220 ( .A(n13054), .ZN(n10728) );
  NOR2_X1 U13221 ( .A1(n14342), .A2(n10728), .ZN(n10729) );
  INV_X1 U13222 ( .A(n14342), .ZN(n14362) );
  NAND2_X1 U13223 ( .A1(n10976), .A2(n12943), .ZN(n10732) );
  AOI22_X1 U13224 ( .A1(n10730), .A2(n9142), .B1(n11862), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n10731) );
  NAND2_X1 U13225 ( .A1(n10733), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n10747) );
  OR2_X1 U13226 ( .A1(n10733), .A2(P2_REG3_REG_15__SCAN_IN), .ZN(n10734) );
  NAND2_X1 U13227 ( .A1(n10747), .A2(n10734), .ZN(n11022) );
  NAND2_X1 U13228 ( .A1(n11688), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n10735) );
  OAI21_X1 U13229 ( .B1(n11022), .B2(n11663), .A(n10735), .ZN(n10739) );
  NAND2_X1 U13230 ( .A1(n11123), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n10737) );
  NAND2_X1 U13231 ( .A1(n11701), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n10736) );
  NAND2_X1 U13232 ( .A1(n10737), .A2(n10736), .ZN(n10738) );
  XNOR2_X1 U13233 ( .A(n10934), .B(n13010), .ZN(n14353) );
  NOR2_X1 U13234 ( .A1(n10741), .A2(n14323), .ZN(n10742) );
  OAI21_X1 U13235 ( .B1(n10744), .B2(n13010), .A(n10942), .ZN(n14359) );
  INV_X1 U13236 ( .A(n12842), .ZN(n14356) );
  OAI211_X1 U13237 ( .C1(n14356), .C2(n10745), .A(n14714), .B(n10931), .ZN(
        n14355) );
  INV_X1 U13238 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10746) );
  NAND2_X1 U13239 ( .A1(n10747), .A2(n10746), .ZN(n10748) );
  NAND2_X1 U13240 ( .A1(n10936), .A2(n10748), .ZN(n12655) );
  NAND2_X1 U13241 ( .A1(n11123), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n10750) );
  NAND2_X1 U13242 ( .A1(n11701), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n10749) );
  AND2_X1 U13243 ( .A1(n10750), .A2(n10749), .ZN(n10752) );
  NAND2_X1 U13244 ( .A1(n11688), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n10751) );
  OAI211_X1 U13245 ( .C1(n12655), .C2(n11663), .A(n10752), .B(n10751), .ZN(
        n13052) );
  NAND2_X1 U13246 ( .A1(n13052), .A2(n12711), .ZN(n10754) );
  NAND2_X1 U13247 ( .A1(n13054), .A2(n12710), .ZN(n10753) );
  NAND2_X1 U13248 ( .A1(n10754), .A2(n10753), .ZN(n11020) );
  INV_X1 U13249 ( .A(n11020), .ZN(n14354) );
  OAI22_X1 U13250 ( .A1(n14708), .A2(n14354), .B1(n11022), .B2(n14706), .ZN(
        n10756) );
  NOR2_X1 U13251 ( .A1(n14356), .A2(n14721), .ZN(n10755) );
  AOI211_X1 U13252 ( .C1(n14708), .C2(P2_REG2_REG_15__SCAN_IN), .A(n10756), 
        .B(n10755), .ZN(n10757) );
  OAI21_X1 U13253 ( .B1(n13282), .B2(n14355), .A(n10757), .ZN(n10758) );
  AOI21_X1 U13254 ( .B1(n14359), .B2(n14727), .A(n10758), .ZN(n10759) );
  OAI21_X1 U13255 ( .B1(n14353), .B2(n13198), .A(n10759), .ZN(P2_U3250) );
  OAI222_X1 U13256 ( .A1(n13440), .A2(n10761), .B1(P2_U3088), .B2(n14742), 
        .C1(n13438), .C2(n10760), .ZN(P2_U3306) );
  OR2_X1 U13257 ( .A1(n11281), .A2(n11285), .ZN(n10764) );
  NAND2_X1 U13258 ( .A1(n10765), .A2(n9599), .ZN(n10768) );
  AOI22_X1 U13259 ( .A1(n10766), .A2(n11317), .B1(n11548), .B2(
        P2_DATAO_REG_13__SCAN_IN), .ZN(n10767) );
  XNOR2_X1 U13260 ( .A(n14432), .B(n11283), .ZN(n11591) );
  INV_X1 U13261 ( .A(n11591), .ZN(n10968) );
  XNOR2_X1 U13262 ( .A(n10969), .B(n10968), .ZN(n14436) );
  INV_X1 U13263 ( .A(n12010), .ZN(n13877) );
  OR2_X1 U13264 ( .A1(n11281), .A2(n13657), .ZN(n10770) );
  XNOR2_X1 U13265 ( .A(n10997), .B(n11591), .ZN(n14439) );
  NAND2_X1 U13266 ( .A1(n14439), .A2(n14383), .ZN(n10788) );
  NAND2_X1 U13267 ( .A1(n10771), .A2(n14432), .ZN(n10772) );
  NAND2_X1 U13268 ( .A1(n14381), .A2(n10772), .ZN(n14435) );
  INV_X1 U13269 ( .A(n14435), .ZN(n10786) );
  INV_X1 U13270 ( .A(n14432), .ZN(n10784) );
  NAND2_X1 U13271 ( .A1(n6482), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n10781) );
  OR2_X1 U13272 ( .A1(n6483), .A2(n10773), .ZN(n10780) );
  AND2_X1 U13273 ( .A1(n10775), .A2(n10774), .ZN(n10776) );
  OR2_X1 U13274 ( .A1(n10776), .A2(n10981), .ZN(n14386) );
  OR2_X1 U13275 ( .A1(n11470), .A2(n14386), .ZN(n10779) );
  INV_X1 U13276 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n10777) );
  OR2_X1 U13277 ( .A1(n11516), .A2(n10777), .ZN(n10778) );
  NAND4_X1 U13278 ( .A1(n10781), .A2(n10780), .A3(n10779), .A4(n10778), .ZN(
        n13656) );
  AOI22_X1 U13279 ( .A1(n14527), .A2(n13657), .B1(n13656), .B2(n14524), .ZN(
        n14434) );
  OAI22_X1 U13280 ( .A1(n14388), .A2(n14434), .B1(n11055), .B2(n14532), .ZN(
        n10782) );
  AOI21_X1 U13281 ( .B1(P1_REG2_REG_13__SCAN_IN), .B2(n14531), .A(n10782), 
        .ZN(n10783) );
  OAI21_X1 U13282 ( .B1(n10784), .B2(n14534), .A(n10783), .ZN(n10785) );
  AOI21_X1 U13283 ( .B1(n10786), .B2(n14519), .A(n10785), .ZN(n10787) );
  OAI211_X1 U13284 ( .C1(n14436), .C2(n13877), .A(n10788), .B(n10787), .ZN(
        P1_U3280) );
  INV_X1 U13285 ( .A(n11259), .ZN(n14595) );
  INV_X1 U13286 ( .A(n10789), .ZN(n10790) );
  NAND2_X1 U13287 ( .A1(n10791), .A2(n10790), .ZN(n10838) );
  NOR2_X1 U13288 ( .A1(n10792), .A2(n13538), .ZN(n10793) );
  AOI21_X1 U13289 ( .B1(n11259), .B2(n13442), .A(n10793), .ZN(n10837) );
  INV_X1 U13290 ( .A(n10837), .ZN(n10794) );
  AOI22_X1 U13291 ( .A1(n11259), .A2(n13481), .B1(n13442), .B2(n13660), .ZN(
        n10795) );
  XNOR2_X1 U13292 ( .A(n10795), .B(n13536), .ZN(n10796) );
  OAI21_X1 U13293 ( .B1(n10797), .B2(n10796), .A(n10846), .ZN(n10798) );
  NAND2_X1 U13294 ( .A1(n10798), .A2(n13626), .ZN(n10803) );
  NOR2_X1 U13295 ( .A1(n13644), .A2(n10799), .ZN(n10801) );
  NAND2_X1 U13296 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3086), .ZN(n13767) );
  OAI21_X1 U13297 ( .B1(n13617), .B2(n10842), .A(n13767), .ZN(n10800) );
  AOI211_X1 U13298 ( .C1(n13620), .C2(n13661), .A(n10801), .B(n10800), .ZN(
        n10802) );
  OAI211_X1 U13299 ( .C1(n14595), .C2(n13636), .A(n10803), .B(n10802), .ZN(
        P1_U3231) );
  XNOR2_X1 U13300 ( .A(n10804), .B(n10806), .ZN(n10810) );
  INV_X1 U13301 ( .A(n14968), .ZN(n12340) );
  OAI211_X1 U13302 ( .C1(n10807), .C2(n10806), .A(n10805), .B(n14961), .ZN(
        n10808) );
  OAI211_X1 U13303 ( .C1(n10810), .C2(n12340), .A(n10809), .B(n10808), .ZN(
        n15011) );
  INV_X1 U13304 ( .A(n15011), .ZN(n10816) );
  INV_X1 U13305 ( .A(n10810), .ZN(n15013) );
  NOR2_X1 U13306 ( .A1(n10811), .A2(n14298), .ZN(n15012) );
  AOI22_X1 U13307 ( .A1(n12479), .A2(n15012), .B1(n14973), .B2(n10812), .ZN(
        n10813) );
  OAI21_X1 U13308 ( .B1(n10333), .B2(n14977), .A(n10813), .ZN(n10814) );
  AOI21_X1 U13309 ( .B1(n15013), .B2(n14974), .A(n10814), .ZN(n10815) );
  OAI21_X1 U13310 ( .B1(n10816), .B2(n14979), .A(n10815), .ZN(P3_U3224) );
  INV_X1 U13311 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n13131) );
  AOI22_X1 U13312 ( .A1(n11027), .A2(P2_REG2_REG_17__SCAN_IN), .B1(n13131), 
        .B2(n13136), .ZN(n10820) );
  NAND2_X1 U13313 ( .A1(n10820), .A2(n10819), .ZN(n13130) );
  OAI21_X1 U13314 ( .B1(n10820), .B2(n10819), .A(n13130), .ZN(n10830) );
  NAND2_X1 U13315 ( .A1(P2_U3088), .A2(P2_REG3_REG_17__SCAN_IN), .ZN(n12666)
         );
  OAI21_X1 U13316 ( .B1(n14667), .B2(n13136), .A(n12666), .ZN(n10828) );
  INV_X1 U13317 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n13137) );
  AOI22_X1 U13318 ( .A1(n11027), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n13137), 
        .B2(n13136), .ZN(n10825) );
  OAI21_X1 U13319 ( .B1(n10823), .B2(n10822), .A(n10821), .ZN(n10824) );
  NAND2_X1 U13320 ( .A1(n10825), .A2(n10824), .ZN(n13135) );
  OAI21_X1 U13321 ( .B1(n10825), .B2(n10824), .A(n13135), .ZN(n10826) );
  NOR2_X1 U13322 ( .A1(n10826), .A2(n14639), .ZN(n10827) );
  AOI211_X1 U13323 ( .C1(n14685), .C2(P2_ADDR_REG_17__SCAN_IN), .A(n10828), 
        .B(n10827), .ZN(n10829) );
  OAI21_X1 U13324 ( .B1(n10830), .B2(n14677), .A(n10829), .ZN(P2_U3231) );
  INV_X1 U13325 ( .A(n10831), .ZN(n10919) );
  XNOR2_X1 U13326 ( .A(n10860), .B(n10859), .ZN(n10862) );
  XNOR2_X1 U13327 ( .A(n10862), .B(n12132), .ZN(n10832) );
  NAND2_X1 U13328 ( .A1(n10832), .A2(n14276), .ZN(n10836) );
  INV_X1 U13329 ( .A(P3_REG3_REG_11__SCAN_IN), .ZN(n15073) );
  NOR2_X1 U13330 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n15073), .ZN(n14891) );
  AOI22_X1 U13331 ( .A1(n12133), .A2(n12440), .B1(n12437), .B2(n12131), .ZN(
        n10923) );
  NOR2_X1 U13332 ( .A1(n10923), .A2(n14281), .ZN(n10833) );
  AOI211_X1 U13333 ( .C1(n14274), .C2(n10834), .A(n14891), .B(n10833), .ZN(
        n10835) );
  OAI211_X1 U13334 ( .C1(n10919), .C2(n14286), .A(n10836), .B(n10835), .ZN(
        P3_U3176) );
  NAND2_X1 U13335 ( .A1(n10838), .A2(n10837), .ZN(n10844) );
  AND2_X1 U13336 ( .A1(n10844), .A2(n10846), .ZN(n10848) );
  NAND2_X1 U13337 ( .A1(n11268), .A2(n13481), .ZN(n10840) );
  NAND2_X1 U13338 ( .A1(n13659), .A2(n13442), .ZN(n10839) );
  NAND2_X1 U13339 ( .A1(n10840), .A2(n10839), .ZN(n10841) );
  XNOR2_X1 U13340 ( .A(n10841), .B(n13536), .ZN(n10886) );
  NOR2_X1 U13341 ( .A1(n10842), .A2(n13538), .ZN(n10843) );
  AOI21_X1 U13342 ( .B1(n11268), .B2(n13442), .A(n10843), .ZN(n10884) );
  XNOR2_X1 U13343 ( .A(n10886), .B(n10884), .ZN(n10847) );
  OAI211_X1 U13344 ( .C1(n10848), .C2(n10847), .A(n13626), .B(n10890), .ZN(
        n10854) );
  NOR2_X1 U13345 ( .A1(n13644), .A2(n10849), .ZN(n10852) );
  OAI21_X1 U13346 ( .B1(n13617), .B2(n10882), .A(n10850), .ZN(n10851) );
  AOI211_X1 U13347 ( .C1(n13620), .C2(n13660), .A(n10852), .B(n10851), .ZN(
        n10853) );
  OAI211_X1 U13348 ( .C1(n14607), .C2(n13636), .A(n10854), .B(n10853), .ZN(
        P1_U3217) );
  OAI22_X1 U13349 ( .A1(n10855), .A2(P3_U3151), .B1(n15171), .B2(n12589), .ZN(
        n10856) );
  AOI21_X1 U13350 ( .B1(n10857), .B2(n12596), .A(n10856), .ZN(n10858) );
  INV_X1 U13351 ( .A(n10858), .ZN(P3_U3271) );
  OAI22_X1 U13352 ( .A1(n10862), .A2(n10861), .B1(n10860), .B2(n10859), .ZN(
        n10865) );
  XNOR2_X1 U13353 ( .A(n10863), .B(n12131), .ZN(n10864) );
  XNOR2_X1 U13354 ( .A(n10865), .B(n10864), .ZN(n10866) );
  NAND2_X1 U13355 ( .A1(n10866), .A2(n14276), .ZN(n10869) );
  AND2_X1 U13356 ( .A1(P3_U3151), .A2(P3_REG3_REG_12__SCAN_IN), .ZN(n12152) );
  AOI22_X1 U13357 ( .A1(n12132), .A2(n12440), .B1(n12437), .B2(n12130), .ZN(
        n12482) );
  NOR2_X1 U13358 ( .A1(n12482), .A2(n14281), .ZN(n10867) );
  AOI211_X1 U13359 ( .C1(n12476), .C2(n12112), .A(n12152), .B(n10867), .ZN(
        n10868) );
  OAI211_X1 U13360 ( .C1(n12475), .C2(n12095), .A(n10869), .B(n10868), .ZN(
        P3_U3164) );
  INV_X1 U13361 ( .A(n10871), .ZN(n10872) );
  XNOR2_X1 U13362 ( .A(n12455), .B(n11971), .ZN(n11927) );
  XNOR2_X1 U13363 ( .A(n11927), .B(n11930), .ZN(n10874) );
  NAND2_X1 U13364 ( .A1(n10875), .A2(n10874), .ZN(n11928) );
  OAI211_X1 U13365 ( .C1(n10875), .C2(n10874), .A(n11928), .B(n14276), .ZN(
        n10878) );
  AOI22_X1 U13366 ( .A1(n12440), .A2(n12130), .B1(n12129), .B2(n12437), .ZN(
        n12453) );
  NAND2_X1 U13367 ( .A1(P3_U3151), .A2(P3_REG3_REG_14__SCAN_IN), .ZN(n12190)
         );
  OAI21_X1 U13368 ( .B1(n12453), .B2(n14281), .A(n12190), .ZN(n10876) );
  AOI21_X1 U13369 ( .B1(n12456), .B2(n12112), .A(n10876), .ZN(n10877) );
  OAI211_X1 U13370 ( .C1(n12095), .C2(n12455), .A(n10878), .B(n10877), .ZN(
        P3_U3155) );
  INV_X1 U13371 ( .A(n11273), .ZN(n14441) );
  NAND2_X1 U13372 ( .A1(n11273), .A2(n13481), .ZN(n10880) );
  NAND2_X1 U13373 ( .A1(n13658), .A2(n13442), .ZN(n10879) );
  NAND2_X1 U13374 ( .A1(n10880), .A2(n10879), .ZN(n10881) );
  XNOR2_X1 U13375 ( .A(n10881), .B(n13536), .ZN(n10901) );
  NOR2_X1 U13376 ( .A1(n10882), .A2(n13538), .ZN(n10883) );
  AOI21_X1 U13377 ( .B1(n11273), .B2(n13442), .A(n10883), .ZN(n10902) );
  XNOR2_X1 U13378 ( .A(n10901), .B(n10902), .ZN(n10888) );
  INV_X1 U13379 ( .A(n10884), .ZN(n10885) );
  NAND2_X1 U13380 ( .A1(n10886), .A2(n10885), .ZN(n10889) );
  INV_X1 U13381 ( .A(n10908), .ZN(n10892) );
  AOI21_X1 U13382 ( .B1(n10890), .B2(n10889), .A(n10888), .ZN(n10891) );
  OAI21_X1 U13383 ( .B1(n10892), .B2(n10891), .A(n13626), .ZN(n10897) );
  NOR2_X1 U13384 ( .A1(n13644), .A2(n10893), .ZN(n10895) );
  NAND2_X1 U13385 ( .A1(P1_REG3_REG_11__SCAN_IN), .A2(P1_U3086), .ZN(n13781)
         );
  OAI21_X1 U13386 ( .B1(n13617), .B2(n11285), .A(n13781), .ZN(n10894) );
  AOI211_X1 U13387 ( .C1(n13620), .C2(n13659), .A(n10895), .B(n10894), .ZN(
        n10896) );
  OAI211_X1 U13388 ( .C1(n14441), .C2(n13636), .A(n10897), .B(n10896), .ZN(
        P1_U3236) );
  INV_X1 U13389 ( .A(SI_25_), .ZN(n15088) );
  INV_X1 U13390 ( .A(n10898), .ZN(n10900) );
  OAI222_X1 U13391 ( .A1(n12589), .A2(n15088), .B1(n12607), .B2(n10900), .C1(
        n10899), .C2(P3_U3151), .ZN(P3_U3270) );
  INV_X1 U13392 ( .A(n10901), .ZN(n10903) );
  NAND2_X1 U13393 ( .A1(n10903), .A2(n10902), .ZN(n10906) );
  AND2_X1 U13394 ( .A1(n10908), .A2(n10906), .ZN(n10910) );
  OAI22_X1 U13395 ( .A1(n14260), .A2(n13535), .B1(n11285), .B2(n13539), .ZN(
        n10904) );
  XNOR2_X1 U13396 ( .A(n10904), .B(n13536), .ZN(n11048) );
  NOR2_X1 U13397 ( .A1(n11285), .A2(n13538), .ZN(n10905) );
  AOI21_X1 U13398 ( .B1(n11281), .B2(n13442), .A(n10905), .ZN(n11049) );
  XNOR2_X1 U13399 ( .A(n11048), .B(n11049), .ZN(n10909) );
  OAI211_X1 U13400 ( .C1(n10910), .C2(n10909), .A(n13626), .B(n11052), .ZN(
        n10915) );
  NOR2_X1 U13401 ( .A1(n13644), .A2(n10911), .ZN(n10913) );
  NAND2_X1 U13402 ( .A1(P1_REG3_REG_12__SCAN_IN), .A2(P1_U3086), .ZN(n14493)
         );
  OAI21_X1 U13403 ( .B1(n13617), .B2(n11283), .A(n14493), .ZN(n10912) );
  AOI211_X1 U13404 ( .C1(n13620), .C2(n13658), .A(n10913), .B(n10912), .ZN(
        n10914) );
  OAI211_X1 U13405 ( .C1(n14260), .C2(n13636), .A(n10915), .B(n10914), .ZN(
        P1_U3224) );
  OAI21_X1 U13406 ( .B1(n6607), .B2(n10917), .A(n10916), .ZN(n14310) );
  INV_X1 U13407 ( .A(n14310), .ZN(n10927) );
  NOR2_X1 U13408 ( .A1(n10918), .A2(n14298), .ZN(n14309) );
  OAI22_X1 U13409 ( .A1(n14977), .A2(n14874), .B1(n10919), .B2(n14959), .ZN(
        n10920) );
  AOI21_X1 U13410 ( .B1(n12479), .B2(n14309), .A(n10920), .ZN(n10926) );
  XNOR2_X1 U13411 ( .A(n10921), .B(n10922), .ZN(n10924) );
  OAI21_X1 U13412 ( .B1(n10924), .B2(n14949), .A(n10923), .ZN(n14308) );
  NAND2_X1 U13413 ( .A1(n14308), .A2(n14977), .ZN(n10925) );
  OAI211_X1 U13414 ( .C1(n10927), .C2(n12486), .A(n10926), .B(n10925), .ZN(
        P3_U3222) );
  NAND2_X1 U13415 ( .A1(n11088), .A2(n11860), .ZN(n10930) );
  AOI22_X1 U13416 ( .A1(n9097), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n10928), 
        .B2(n9142), .ZN(n10929) );
  AOI211_X1 U13417 ( .C1(n13404), .C2(n10931), .A(n9329), .B(n11036), .ZN(
        n13403) );
  AND2_X1 U13418 ( .A1(n12842), .A2(n10740), .ZN(n10933) );
  OR2_X1 U13419 ( .A1(n12842), .A2(n10740), .ZN(n10932) );
  XNOR2_X1 U13420 ( .A(n13404), .B(n13052), .ZN(n13011) );
  XNOR2_X1 U13421 ( .A(n11032), .B(n13011), .ZN(n10940) );
  INV_X1 U13422 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n10935) );
  AND2_X1 U13423 ( .A1(n10936), .A2(n10935), .ZN(n10937) );
  OR2_X1 U13424 ( .A1(n10937), .A2(n11037), .ZN(n12665) );
  AOI22_X1 U13425 ( .A1(n11701), .A2(P2_REG1_REG_17__SCAN_IN), .B1(n11123), 
        .B2(P2_REG0_REG_17__SCAN_IN), .ZN(n10939) );
  NAND2_X1 U13426 ( .A1(n11688), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n10938) );
  OAI211_X1 U13427 ( .C1(n12665), .C2(n11663), .A(n10939), .B(n10938), .ZN(
        n13051) );
  AOI22_X1 U13428 ( .A1(n13051), .A2(n12711), .B1(n12710), .B2(n13053), .ZN(
        n12657) );
  OAI21_X1 U13429 ( .B1(n10940), .B2(n14352), .A(n12657), .ZN(n13402) );
  AOI21_X1 U13430 ( .B1(n13403), .B2(n13253), .A(n13402), .ZN(n10948) );
  OAI22_X1 U13431 ( .A1(n13316), .A2(n10818), .B1(n12655), .B2(n14706), .ZN(
        n10946) );
  NAND2_X1 U13432 ( .A1(n10942), .A2(n10941), .ZN(n10943) );
  NOR2_X1 U13433 ( .A1(n10943), .A2(n13011), .ZN(n11026) );
  AOI21_X1 U13434 ( .B1(n13011), .B2(n10943), .A(n11026), .ZN(n10944) );
  INV_X1 U13435 ( .A(n10944), .ZN(n13407) );
  NOR2_X1 U13436 ( .A1(n13407), .A2(n13304), .ZN(n10945) );
  AOI211_X1 U13437 ( .C1(n14341), .C2(n13404), .A(n10946), .B(n10945), .ZN(
        n10947) );
  OAI21_X1 U13438 ( .B1(n14731), .B2(n10948), .A(n10947), .ZN(P2_U3249) );
  OAI21_X1 U13439 ( .B1(n10950), .B2(n10953), .A(n10949), .ZN(n13792) );
  XNOR2_X1 U13440 ( .A(n10959), .B(n13792), .ZN(n10951) );
  NAND2_X1 U13441 ( .A1(P1_REG2_REG_18__SCAN_IN), .A2(n10951), .ZN(n13794) );
  OAI211_X1 U13442 ( .C1(P1_REG2_REG_18__SCAN_IN), .C2(n10951), .A(n14508), 
        .B(n13794), .ZN(n10958) );
  NAND2_X1 U13443 ( .A1(P1_U3086), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n13615)
         );
  OAI21_X1 U13444 ( .B1(n11103), .B2(n10953), .A(n10952), .ZN(n13796) );
  XNOR2_X1 U13445 ( .A(n13796), .B(n10959), .ZN(n10954) );
  NAND2_X1 U13446 ( .A1(P1_REG1_REG_18__SCAN_IN), .A2(n10954), .ZN(n13799) );
  OAI211_X1 U13447 ( .C1(P1_REG1_REG_18__SCAN_IN), .C2(n10954), .A(n14504), 
        .B(n13799), .ZN(n10955) );
  NAND2_X1 U13448 ( .A1(n13615), .A2(n10955), .ZN(n10956) );
  AOI21_X1 U13449 ( .B1(n14497), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n10956), 
        .ZN(n10957) );
  OAI211_X1 U13450 ( .C1(n14501), .C2(n10959), .A(n10958), .B(n10957), .ZN(
        P1_U3261) );
  NAND2_X1 U13451 ( .A1(n11071), .A2(SI_22_), .ZN(n11060) );
  MUX2_X1 U13452 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(P1_DATAO_REG_22__SCAN_IN), 
        .S(n11543), .Z(n11072) );
  NAND2_X1 U13453 ( .A1(n11362), .A2(n11072), .ZN(n11061) );
  INV_X1 U13454 ( .A(n11362), .ZN(n10964) );
  INV_X1 U13455 ( .A(n11072), .ZN(n10963) );
  NAND2_X1 U13456 ( .A1(n10964), .A2(n10963), .ZN(n10965) );
  INV_X1 U13457 ( .A(n11659), .ZN(n10966) );
  OAI222_X1 U13458 ( .A1(n13440), .A2(n10967), .B1(P2_U3088), .B2(n12720), 
        .C1(n13438), .C2(n10966), .ZN(P2_U3305) );
  AOI22_X1 U13459 ( .A1(n10971), .A2(n11317), .B1(n11548), .B2(
        P2_DATAO_REG_14__SCAN_IN), .ZN(n10972) );
  NAND2_X2 U13460 ( .A1(n10973), .A2(n10972), .ZN(n14397) );
  NAND2_X1 U13461 ( .A1(n14390), .A2(n14391), .ZN(n10975) );
  INV_X1 U13462 ( .A(n13656), .ZN(n10974) );
  OR2_X1 U13463 ( .A1(n14397), .A2(n10974), .ZN(n11295) );
  NAND2_X1 U13464 ( .A1(n10975), .A2(n11295), .ZN(n11093) );
  NAND2_X1 U13465 ( .A1(n10976), .A2(n9599), .ZN(n10979) );
  AOI22_X1 U13466 ( .A1(n11548), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n11317), 
        .B2(n10977), .ZN(n10978) );
  NAND2_X1 U13467 ( .A1(n11503), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n10986) );
  INV_X1 U13468 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n10980) );
  OR2_X1 U13469 ( .A1(n6483), .A2(n10980), .ZN(n10985) );
  INV_X1 U13470 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n11000) );
  OR2_X1 U13471 ( .A1(n6487), .A2(n11000), .ZN(n10984) );
  OR2_X1 U13472 ( .A1(n10981), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n10982) );
  NAND2_X1 U13473 ( .A1(n10989), .A2(n10982), .ZN(n13645) );
  OR2_X1 U13474 ( .A1(n6468), .A2(n13645), .ZN(n10983) );
  NAND2_X1 U13475 ( .A1(n13648), .A2(n13504), .ZN(n11298) );
  NAND2_X1 U13476 ( .A1(n11297), .A2(n11298), .ZN(n11593) );
  XNOR2_X1 U13477 ( .A(n11093), .B(n11593), .ZN(n10987) );
  NAND2_X1 U13478 ( .A1(n10987), .A2(n14392), .ZN(n10996) );
  NAND2_X1 U13479 ( .A1(n10989), .A2(n10988), .ZN(n10990) );
  NAND2_X1 U13480 ( .A1(n11100), .A2(n10990), .ZN(n13576) );
  OR2_X1 U13481 ( .A1(n11470), .A2(n13576), .ZN(n10994) );
  NAND2_X1 U13482 ( .A1(n11503), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n10993) );
  OR2_X1 U13483 ( .A1(n6483), .A2(n14417), .ZN(n10992) );
  OR2_X1 U13484 ( .A1(n6487), .A2(n11110), .ZN(n10991) );
  NAND4_X1 U13485 ( .A1(n10994), .A2(n10993), .A3(n10992), .A4(n10991), .ZN(
        n13655) );
  AOI22_X1 U13486 ( .A1(n14524), .A2(n13655), .B1(n13656), .B2(n14527), .ZN(
        n10995) );
  NAND2_X1 U13487 ( .A1(n10996), .A2(n10995), .ZN(n14421) );
  INV_X1 U13488 ( .A(n14421), .ZN(n11005) );
  NAND2_X1 U13489 ( .A1(n14397), .A2(n13656), .ZN(n10998) );
  INV_X1 U13490 ( .A(n11593), .ZN(n11092) );
  OAI21_X1 U13491 ( .B1(n6507), .B2(n11593), .A(n11098), .ZN(n14422) );
  INV_X1 U13492 ( .A(n13648), .ZN(n14418) );
  INV_X1 U13493 ( .A(n10999), .ZN(n14380) );
  INV_X1 U13494 ( .A(n11113), .ZN(n11111) );
  OAI21_X1 U13495 ( .B1(n14418), .B2(n14380), .A(n11111), .ZN(n14419) );
  OAI22_X1 U13496 ( .A1(n13893), .A2(n11000), .B1(n13645), .B2(n14532), .ZN(
        n11001) );
  AOI21_X1 U13497 ( .B1(n13648), .B2(n14398), .A(n11001), .ZN(n11002) );
  OAI21_X1 U13498 ( .B1(n14419), .B2(n13989), .A(n11002), .ZN(n11003) );
  AOI21_X1 U13499 ( .B1(n14422), .B2(n14383), .A(n11003), .ZN(n11004) );
  OAI21_X1 U13500 ( .B1(n14531), .B2(n11005), .A(n11004), .ZN(P1_U3278) );
  INV_X1 U13501 ( .A(n11007), .ZN(n11010) );
  INV_X1 U13502 ( .A(n11008), .ZN(n11009) );
  NAND2_X1 U13503 ( .A1(n11010), .A2(n11009), .ZN(n11011) );
  INV_X1 U13504 ( .A(n11013), .ZN(n14326) );
  XNOR2_X1 U13505 ( .A(n14342), .B(n11628), .ZN(n11014) );
  NAND2_X1 U13506 ( .A1(n13054), .A2(n11749), .ZN(n11015) );
  NAND2_X1 U13507 ( .A1(n11014), .A2(n11015), .ZN(n11019) );
  INV_X1 U13508 ( .A(n11014), .ZN(n11017) );
  INV_X1 U13509 ( .A(n11015), .ZN(n11016) );
  NAND2_X1 U13510 ( .A1(n11017), .A2(n11016), .ZN(n11018) );
  AND2_X1 U13511 ( .A1(n11019), .A2(n11018), .ZN(n14327) );
  NAND2_X1 U13512 ( .A1(n14326), .A2(n14327), .ZN(n14325) );
  NAND2_X1 U13513 ( .A1(n13053), .A2(n11749), .ZN(n11622) );
  XNOR2_X1 U13514 ( .A(n11623), .B(n11622), .ZN(n11025) );
  AOI22_X1 U13515 ( .A1(n14330), .A2(n11020), .B1(P2_REG3_REG_15__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11021) );
  OAI21_X1 U13516 ( .B1(n11022), .B2(n14334), .A(n11021), .ZN(n11023) );
  AOI21_X1 U13517 ( .B1(n12842), .B2(n12703), .A(n11023), .ZN(n11024) );
  OAI21_X1 U13518 ( .B1(n11025), .B2(n12705), .A(n11024), .ZN(P2_U3213) );
  NAND2_X1 U13519 ( .A1(n11305), .A2(n12943), .ZN(n11029) );
  AOI22_X1 U13520 ( .A1(n11027), .A2(n9142), .B1(n11862), .B2(
        P1_DATAO_REG_17__SCAN_IN), .ZN(n11028) );
  XNOR2_X1 U13521 ( .A(n12851), .B(n13051), .ZN(n13013) );
  NOR2_X1 U13522 ( .A1(n11030), .A2(n13013), .ZN(n11133) );
  AOI21_X1 U13523 ( .B1(n11030), .B2(n13013), .A(n11133), .ZN(n11031) );
  INV_X1 U13524 ( .A(n11031), .ZN(n13401) );
  NAND2_X1 U13525 ( .A1(n11032), .A2(n13011), .ZN(n11035) );
  INV_X1 U13526 ( .A(n13052), .ZN(n11033) );
  OR2_X1 U13527 ( .A1(n13404), .A2(n11033), .ZN(n11034) );
  XOR2_X1 U13528 ( .A(n13013), .B(n11136), .Z(n13399) );
  INV_X1 U13529 ( .A(n12851), .ZN(n13397) );
  OAI211_X1 U13530 ( .C1(n11036), .C2(n13397), .A(n13313), .B(n14714), .ZN(
        n13396) );
  NOR2_X1 U13531 ( .A1(n13396), .A2(n13282), .ZN(n11046) );
  NAND2_X1 U13532 ( .A1(n12851), .A2(n14341), .ZN(n11044) );
  NAND2_X1 U13533 ( .A1(n11037), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n11121) );
  OR2_X1 U13534 ( .A1(n11037), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n11038) );
  NAND2_X1 U13535 ( .A1(n11121), .A2(n11038), .ZN(n13315) );
  AOI22_X1 U13536 ( .A1(n9113), .A2(P2_REG1_REG_18__SCAN_IN), .B1(n11688), 
        .B2(P2_REG2_REG_18__SCAN_IN), .ZN(n11040) );
  NAND2_X1 U13537 ( .A1(n11123), .A2(P2_REG0_REG_18__SCAN_IN), .ZN(n11039) );
  OAI211_X1 U13538 ( .C1(n13315), .C2(n11663), .A(n11040), .B(n11039), .ZN(
        n13050) );
  AND2_X1 U13539 ( .A1(n13052), .A2(n12710), .ZN(n11041) );
  AOI21_X1 U13540 ( .B1(n13050), .B2(n12711), .A(n11041), .ZN(n13395) );
  OAI22_X1 U13541 ( .A1(n14708), .A2(n13395), .B1(n12665), .B2(n14706), .ZN(
        n11042) );
  INV_X1 U13542 ( .A(n11042), .ZN(n11043) );
  OAI211_X1 U13543 ( .C1(n13316), .C2(n13131), .A(n11044), .B(n11043), .ZN(
        n11045) );
  AOI211_X1 U13544 ( .C1(n13399), .C2(n13284), .A(n11046), .B(n11045), .ZN(
        n11047) );
  OAI21_X1 U13545 ( .B1(n13401), .B2(n13304), .A(n11047), .ZN(P2_U3248) );
  INV_X1 U13546 ( .A(n11049), .ZN(n11050) );
  NOR2_X1 U13547 ( .A1(n11283), .A2(n13538), .ZN(n11053) );
  AOI21_X1 U13548 ( .B1(n14432), .B2(n13442), .A(n11053), .ZN(n11767) );
  AOI22_X1 U13549 ( .A1(n14432), .A2(n13481), .B1(n13442), .B2(n14394), .ZN(
        n11054) );
  XNOR2_X1 U13550 ( .A(n11054), .B(n13536), .ZN(n11766) );
  XOR2_X1 U13551 ( .A(n11767), .B(n11766), .Z(n11771) );
  XNOR2_X1 U13552 ( .A(n11772), .B(n11771), .ZN(n11059) );
  NOR2_X1 U13553 ( .A1(n13644), .A2(n11055), .ZN(n11057) );
  NAND2_X1 U13554 ( .A1(P1_U3086), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n14499)
         );
  OAI21_X1 U13555 ( .B1(n13513), .B2(n14434), .A(n14499), .ZN(n11056) );
  AOI211_X1 U13556 ( .C1(n14432), .C2(n13647), .A(n11057), .B(n11056), .ZN(
        n11058) );
  OAI21_X1 U13557 ( .B1(n11059), .B2(n13650), .A(n11058), .ZN(P1_U3234) );
  NAND2_X1 U13558 ( .A1(n11061), .A2(n11060), .ZN(n11063) );
  MUX2_X1 U13559 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(P1_DATAO_REG_23__SCAN_IN), 
        .S(n11543), .Z(n11074) );
  XNOR2_X1 U13560 ( .A(n11074), .B(SI_23_), .ZN(n11062) );
  XNOR2_X1 U13561 ( .A(n11063), .B(n11062), .ZN(n11387) );
  NAND2_X1 U13562 ( .A1(n11387), .A2(n11064), .ZN(n11066) );
  AND2_X1 U13563 ( .A1(n11065), .A2(P2_STATE_REG_SCAN_IN), .ZN(n13032) );
  INV_X1 U13564 ( .A(n13032), .ZN(n13030) );
  OAI211_X1 U13565 ( .C1(n11067), .C2(n13440), .A(n11066), .B(n13030), .ZN(
        P2_U3304) );
  NAND2_X1 U13566 ( .A1(n11387), .A2(n11068), .ZN(n11069) );
  OAI211_X1 U13567 ( .C1(n11070), .C2(n14124), .A(n11069), .B(n11616), .ZN(
        P1_U3332) );
  AOI22_X1 U13568 ( .A1(SI_22_), .A2(n11072), .B1(n11074), .B2(SI_23_), .ZN(
        n11073) );
  INV_X1 U13569 ( .A(n11074), .ZN(n11076) );
  NAND2_X1 U13570 ( .A1(n11076), .A2(n11075), .ZN(n11077) );
  MUX2_X1 U13571 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(P1_DATAO_REG_24__SCAN_IN), 
        .S(n11543), .Z(n11080) );
  INV_X1 U13572 ( .A(n11080), .ZN(n11081) );
  NAND2_X1 U13573 ( .A1(n11082), .A2(n11081), .ZN(n11083) );
  NAND2_X1 U13574 ( .A1(n11167), .A2(n11083), .ZN(n11685) );
  OAI222_X1 U13575 ( .A1(P1_U3086), .A2(n11085), .B1(n14119), .B2(n11685), 
        .C1(n11084), .C2(n14124), .ZN(P1_U3331) );
  OAI222_X1 U13576 ( .A1(n11087), .A2(P2_U3088), .B1(n13438), .B2(n11685), 
        .C1(n11086), .C2(n13440), .ZN(P2_U3303) );
  NAND2_X1 U13577 ( .A1(n11088), .A2(n11547), .ZN(n11091) );
  AOI22_X1 U13578 ( .A1(n11548), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(n11317), 
        .B2(n11089), .ZN(n11090) );
  INV_X1 U13579 ( .A(n13655), .ZN(n14007) );
  XNOR2_X1 U13580 ( .A(n14409), .B(n14007), .ZN(n11905) );
  NAND2_X1 U13581 ( .A1(n11093), .A2(n11092), .ZN(n11094) );
  NAND2_X1 U13582 ( .A1(n11094), .A2(n11297), .ZN(n11096) );
  INV_X1 U13583 ( .A(n14003), .ZN(n11095) );
  AOI21_X1 U13584 ( .B1(n11905), .B2(n11096), .A(n11095), .ZN(n14414) );
  INV_X1 U13585 ( .A(n13504), .ZN(n14385) );
  OR2_X1 U13586 ( .A1(n13648), .A2(n14385), .ZN(n11097) );
  XNOR2_X1 U13587 ( .A(n11906), .B(n11905), .ZN(n14416) );
  NAND2_X1 U13588 ( .A1(n14416), .A2(n14383), .ZN(n11117) );
  AND2_X1 U13589 ( .A1(n11100), .A2(n11099), .ZN(n11102) );
  OR2_X1 U13590 ( .A1(n11102), .A2(n11101), .ZN(n13995) );
  OR2_X1 U13591 ( .A1(n6483), .A2(n11103), .ZN(n11105) );
  OR2_X1 U13592 ( .A1(n6487), .A2(n10950), .ZN(n11104) );
  AND2_X1 U13593 ( .A1(n11105), .A2(n11104), .ZN(n11107) );
  NAND2_X1 U13594 ( .A1(n11503), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n11106) );
  OAI211_X1 U13595 ( .C1(n13995), .C2(n6468), .A(n11107), .B(n11106), .ZN(
        n13977) );
  INV_X1 U13596 ( .A(n13977), .ZN(n13573) );
  OAI22_X1 U13597 ( .A1(n13573), .A2(n14008), .B1(n13504), .B2(n14006), .ZN(
        n14408) );
  INV_X1 U13598 ( .A(n13576), .ZN(n11108) );
  AOI22_X1 U13599 ( .A1(n13893), .A2(n14408), .B1(n11108), .B2(n13996), .ZN(
        n11109) );
  OAI21_X1 U13600 ( .B1(n11110), .B2(n13893), .A(n11109), .ZN(n11115) );
  NAND2_X1 U13601 ( .A1(n11111), .A2(n14409), .ZN(n14411) );
  INV_X1 U13602 ( .A(n14409), .ZN(n11112) );
  AND3_X1 U13603 ( .A1(n14411), .A2(n14519), .A3(n14410), .ZN(n11114) );
  AOI211_X1 U13604 ( .C1(n14398), .C2(n14409), .A(n11115), .B(n11114), .ZN(
        n11116) );
  OAI211_X1 U13605 ( .C1(n14414), .C2(n13877), .A(n11117), .B(n11116), .ZN(
        P1_U3277) );
  NAND2_X1 U13606 ( .A1(n11309), .A2(n12943), .ZN(n11119) );
  AOI22_X1 U13607 ( .A1(n12988), .A2(n9142), .B1(n11862), .B2(
        P1_DATAO_REG_19__SCAN_IN), .ZN(n11118) );
  INV_X1 U13608 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n11120) );
  NAND2_X1 U13609 ( .A1(n11121), .A2(n11120), .ZN(n11122) );
  AND2_X1 U13610 ( .A1(n11141), .A2(n11122), .ZN(n12633) );
  NAND2_X1 U13611 ( .A1(n12633), .A2(n9145), .ZN(n11129) );
  INV_X1 U13612 ( .A(P2_REG1_REG_19__SCAN_IN), .ZN(n11126) );
  NAND2_X1 U13613 ( .A1(n11123), .A2(P2_REG0_REG_19__SCAN_IN), .ZN(n11125) );
  NAND2_X1 U13614 ( .A1(n11688), .A2(P2_REG2_REG_19__SCAN_IN), .ZN(n11124) );
  OAI211_X1 U13615 ( .C1(n11872), .C2(n11126), .A(n11125), .B(n11124), .ZN(
        n11127) );
  INV_X1 U13616 ( .A(n11127), .ZN(n11128) );
  NAND2_X1 U13617 ( .A1(n11129), .A2(n11128), .ZN(n13049) );
  INV_X1 U13618 ( .A(n13049), .ZN(n12700) );
  NAND2_X1 U13619 ( .A1(n12873), .A2(n12700), .ZN(n11848) );
  OR2_X1 U13620 ( .A1(n12873), .A2(n12700), .ZN(n11130) );
  NAND2_X1 U13621 ( .A1(n11848), .A2(n11130), .ZN(n13016) );
  NAND2_X1 U13622 ( .A1(n11316), .A2(n11860), .ZN(n11132) );
  AOI22_X1 U13623 ( .A1(n13149), .A2(n9142), .B1(n11862), .B2(
        P1_DATAO_REG_18__SCAN_IN), .ZN(n11131) );
  INV_X1 U13624 ( .A(n13050), .ZN(n11137) );
  XNOR2_X1 U13625 ( .A(n13390), .B(n11137), .ZN(n13307) );
  XOR2_X1 U13626 ( .A(n13016), .B(n11876), .Z(n13389) );
  INV_X1 U13627 ( .A(n13051), .ZN(n12853) );
  NOR2_X1 U13628 ( .A1(n12851), .A2(n12853), .ZN(n11135) );
  NAND2_X1 U13629 ( .A1(n12851), .A2(n12853), .ZN(n11134) );
  OAI21_X2 U13630 ( .B1(n11136), .B2(n11135), .A(n11134), .ZN(n13308) );
  AND2_X1 U13631 ( .A1(n13390), .A2(n11137), .ZN(n11139) );
  OR2_X1 U13632 ( .A1(n13390), .A2(n11137), .ZN(n11138) );
  INV_X1 U13633 ( .A(n13016), .ZN(n11140) );
  OAI21_X1 U13634 ( .B1(n6597), .B2(n11140), .A(n11849), .ZN(n13387) );
  OAI211_X1 U13635 ( .C1(n6859), .C2(n6860), .A(n14714), .B(n13296), .ZN(
        n13385) );
  INV_X1 U13636 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n12683) );
  AND2_X1 U13637 ( .A1(n11141), .A2(n12683), .ZN(n11142) );
  OR2_X1 U13638 ( .A1(n11142), .A2(n11649), .ZN(n13294) );
  INV_X1 U13639 ( .A(P2_REG1_REG_20__SCAN_IN), .ZN(n11145) );
  NAND2_X1 U13640 ( .A1(n11123), .A2(P2_REG0_REG_20__SCAN_IN), .ZN(n11144) );
  NAND2_X1 U13641 ( .A1(n11688), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n11143) );
  OAI211_X1 U13642 ( .C1(n11872), .C2(n11145), .A(n11144), .B(n11143), .ZN(
        n11146) );
  INV_X1 U13643 ( .A(n11146), .ZN(n11147) );
  OAI21_X1 U13644 ( .B1(n13294), .B2(n11663), .A(n11147), .ZN(n13048) );
  AOI22_X1 U13645 ( .A1(n13048), .A2(n12711), .B1(n12710), .B2(n13050), .ZN(
        n13384) );
  INV_X1 U13646 ( .A(n12633), .ZN(n11148) );
  OAI22_X1 U13647 ( .A1(n13384), .A2(n14708), .B1(n11148), .B2(n14706), .ZN(
        n11150) );
  NOR2_X1 U13648 ( .A1(n6859), .A2(n14721), .ZN(n11149) );
  AOI211_X1 U13649 ( .C1(n14708), .C2(P2_REG2_REG_19__SCAN_IN), .A(n11150), 
        .B(n11149), .ZN(n11151) );
  OAI21_X1 U13650 ( .B1(n13282), .B2(n13385), .A(n11151), .ZN(n11152) );
  AOI21_X1 U13651 ( .B1(n13387), .B2(n13284), .A(n11152), .ZN(n11153) );
  OAI21_X1 U13652 ( .B1(n13389), .B2(n13304), .A(n11153), .ZN(P2_U3246) );
  MUX2_X1 U13653 ( .A(n11154), .B(P1_REG2_REG_3__SCAN_IN), .S(n14531), .Z(
        n11162) );
  NAND2_X1 U13654 ( .A1(n11155), .A2(n14520), .ZN(n11159) );
  OAI22_X1 U13655 ( .A1(n13989), .A2(n11156), .B1(P1_REG3_REG_3__SCAN_IN), 
        .B2(n14532), .ZN(n11157) );
  INV_X1 U13656 ( .A(n11157), .ZN(n11158) );
  OAI211_X1 U13657 ( .C1(n11160), .C2(n14534), .A(n11159), .B(n11158), .ZN(
        n11161) );
  OR2_X1 U13658 ( .A1(n11162), .A2(n11161), .ZN(P1_U3290) );
  INV_X1 U13659 ( .A(n12583), .ZN(n11164) );
  INV_X1 U13660 ( .A(n11165), .ZN(P3_U3455) );
  MUX2_X1 U13661 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(P1_DATAO_REG_25__SCAN_IN), 
        .S(n11543), .Z(n11168) );
  XNOR2_X1 U13662 ( .A(n11168), .B(SI_25_), .ZN(n11420) );
  INV_X1 U13663 ( .A(n11168), .ZN(n11169) );
  NAND2_X1 U13664 ( .A1(n11169), .A2(n15088), .ZN(n11170) );
  MUX2_X1 U13665 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(P1_DATAO_REG_26__SCAN_IN), 
        .S(n11543), .Z(n11173) );
  NAND2_X1 U13666 ( .A1(n11173), .A2(SI_26_), .ZN(n11175) );
  OAI21_X1 U13667 ( .B1(SI_26_), .B2(n11173), .A(n11175), .ZN(n11428) );
  INV_X1 U13668 ( .A(n11428), .ZN(n11174) );
  MUX2_X1 U13669 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(P1_DATAO_REG_27__SCAN_IN), 
        .S(n11543), .Z(n11458) );
  INV_X1 U13670 ( .A(n11458), .ZN(n11176) );
  INV_X1 U13671 ( .A(SI_27_), .ZN(n15169) );
  NAND2_X1 U13672 ( .A1(n11176), .A2(n15169), .ZN(n11177) );
  NAND2_X1 U13673 ( .A1(n11458), .A2(SI_27_), .ZN(n11178) );
  MUX2_X1 U13674 ( .A(n11618), .B(n11180), .S(n11543), .Z(n11181) );
  INV_X1 U13675 ( .A(SI_28_), .ZN(n15047) );
  NAND2_X1 U13676 ( .A1(n11181), .A2(n15047), .ZN(n11184) );
  INV_X1 U13677 ( .A(n11181), .ZN(n11182) );
  NAND2_X1 U13678 ( .A1(n11182), .A2(SI_28_), .ZN(n11183) );
  NAND2_X1 U13679 ( .A1(n11184), .A2(n11183), .ZN(n11477) );
  MUX2_X1 U13680 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(P1_DATAO_REG_29__SCAN_IN), 
        .S(n11543), .Z(n11482) );
  INV_X1 U13681 ( .A(SI_29_), .ZN(n11483) );
  XNOR2_X1 U13682 ( .A(n11482), .B(n11483), .ZN(n11480) );
  XNOR2_X1 U13683 ( .A(n11481), .B(n11480), .ZN(n11861) );
  INV_X1 U13684 ( .A(n11861), .ZN(n11187) );
  OAI222_X1 U13685 ( .A1(n14124), .A2(n11186), .B1(n14130), .B2(n11187), .C1(
        n11185), .C2(P1_U3086), .ZN(P1_U3326) );
  OAI222_X1 U13686 ( .A1(n13440), .A2(n11189), .B1(P2_U3088), .B2(n11188), 
        .C1(n13438), .C2(n11187), .ZN(P2_U3298) );
  NAND2_X1 U13687 ( .A1(n11191), .A2(n11190), .ZN(n11207) );
  NAND2_X1 U13688 ( .A1(n11192), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n11194) );
  NAND2_X1 U13689 ( .A1(n14111), .A2(P1_IR_REG_22__SCAN_IN), .ZN(n11193) );
  NAND2_X1 U13690 ( .A1(n11194), .A2(n11193), .ZN(n11202) );
  INV_X1 U13691 ( .A(n11195), .ZN(n11197) );
  NAND2_X1 U13692 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), 
        .ZN(n11196) );
  OAI211_X1 U13693 ( .C1(n11197), .C2(P1_IR_REG_20__SCAN_IN), .A(
        P1_IR_REG_31__SCAN_IN), .B(n11196), .ZN(n11198) );
  NOR2_X1 U13694 ( .A1(n11199), .A2(n11198), .ZN(n11200) );
  AOI21_X1 U13695 ( .B1(n11201), .B2(n11202), .A(n11200), .ZN(n11205) );
  INV_X1 U13696 ( .A(n11202), .ZN(n11203) );
  NAND3_X1 U13697 ( .A1(n11207), .A2(n11212), .A3(n11554), .ZN(n11208) );
  NAND2_X1 U13698 ( .A1(n11208), .A2(n11209), .ZN(n11211) );
  INV_X1 U13699 ( .A(n11209), .ZN(n11210) );
  INV_X1 U13700 ( .A(n11212), .ZN(n11214) );
  NAND2_X1 U13701 ( .A1(n11216), .A2(n11551), .ZN(n11218) );
  NAND3_X1 U13702 ( .A1(n11554), .A2(n14525), .A3(n14555), .ZN(n11217) );
  NAND3_X1 U13703 ( .A1(n11220), .A2(n7472), .A3(n11577), .ZN(n11227) );
  INV_X1 U13704 ( .A(n11221), .ZN(n11224) );
  INV_X1 U13705 ( .A(n11222), .ZN(n11223) );
  MUX2_X1 U13706 ( .A(n11224), .B(n11223), .S(n11551), .Z(n11225) );
  INV_X1 U13707 ( .A(n11225), .ZN(n11226) );
  MUX2_X1 U13708 ( .A(n13665), .B(n11228), .S(n11551), .Z(n11231) );
  MUX2_X1 U13709 ( .A(n13665), .B(n11228), .S(n11554), .Z(n11229) );
  OAI21_X1 U13710 ( .B1(n11232), .B2(n11231), .A(n11230), .ZN(n11235) );
  MUX2_X1 U13711 ( .A(n13664), .B(n11233), .S(n11554), .Z(n11236) );
  MUX2_X1 U13712 ( .A(n13664), .B(n11233), .S(n11551), .Z(n11234) );
  INV_X1 U13713 ( .A(n11236), .ZN(n11237) );
  MUX2_X1 U13714 ( .A(n11238), .B(n13663), .S(n11554), .Z(n11242) );
  NAND2_X1 U13715 ( .A1(n11241), .A2(n11242), .ZN(n11240) );
  MUX2_X1 U13716 ( .A(n11238), .B(n13663), .S(n11551), .Z(n11239) );
  NAND2_X1 U13717 ( .A1(n11240), .A2(n11239), .ZN(n11246) );
  INV_X1 U13718 ( .A(n11242), .ZN(n11243) );
  NAND2_X1 U13719 ( .A1(n11244), .A2(n11243), .ZN(n11245) );
  MUX2_X1 U13720 ( .A(n13662), .B(n14579), .S(n11554), .Z(n11248) );
  MUX2_X1 U13721 ( .A(n13662), .B(n14579), .S(n11551), .Z(n11247) );
  INV_X1 U13722 ( .A(n11248), .ZN(n11249) );
  MUX2_X1 U13723 ( .A(n13661), .B(n11250), .S(n11551), .Z(n11254) );
  NAND2_X1 U13724 ( .A1(n11253), .A2(n11254), .ZN(n11252) );
  MUX2_X1 U13725 ( .A(n13661), .B(n11250), .S(n11554), .Z(n11251) );
  NAND2_X1 U13726 ( .A1(n11252), .A2(n11251), .ZN(n11258) );
  INV_X1 U13727 ( .A(n11253), .ZN(n11256) );
  INV_X1 U13728 ( .A(n11254), .ZN(n11255) );
  NAND2_X1 U13729 ( .A1(n11256), .A2(n11255), .ZN(n11257) );
  NAND2_X1 U13730 ( .A1(n11258), .A2(n11257), .ZN(n11262) );
  MUX2_X1 U13731 ( .A(n13660), .B(n11259), .S(n11554), .Z(n11263) );
  NAND2_X1 U13732 ( .A1(n11262), .A2(n11263), .ZN(n11261) );
  MUX2_X1 U13733 ( .A(n13660), .B(n11259), .S(n11551), .Z(n11260) );
  NAND2_X1 U13734 ( .A1(n11261), .A2(n11260), .ZN(n11267) );
  INV_X1 U13735 ( .A(n11262), .ZN(n11265) );
  INV_X1 U13736 ( .A(n11263), .ZN(n11264) );
  NAND2_X1 U13737 ( .A1(n11265), .A2(n11264), .ZN(n11266) );
  NAND2_X1 U13738 ( .A1(n11267), .A2(n11266), .ZN(n11270) );
  MUX2_X1 U13739 ( .A(n13659), .B(n11268), .S(n11551), .Z(n11271) );
  MUX2_X1 U13740 ( .A(n13659), .B(n11268), .S(n11554), .Z(n11269) );
  INV_X1 U13741 ( .A(n11271), .ZN(n11272) );
  MUX2_X1 U13742 ( .A(n13658), .B(n11273), .S(n11554), .Z(n11277) );
  MUX2_X1 U13743 ( .A(n13658), .B(n11273), .S(n11551), .Z(n11274) );
  NAND2_X1 U13744 ( .A1(n11275), .A2(n11274), .ZN(n11280) );
  INV_X1 U13745 ( .A(n11276), .ZN(n11278) );
  NAND2_X1 U13746 ( .A1(n11278), .A2(n7130), .ZN(n11279) );
  NAND2_X1 U13747 ( .A1(n11280), .A2(n11279), .ZN(n11288) );
  MUX2_X1 U13748 ( .A(n13657), .B(n11281), .S(n11551), .Z(n11287) );
  MUX2_X1 U13749 ( .A(n14394), .B(n14432), .S(n11554), .Z(n11291) );
  NAND2_X1 U13750 ( .A1(n14432), .A2(n11551), .ZN(n11282) );
  OAI211_X1 U13751 ( .C1(n11283), .C2(n11551), .A(n11291), .B(n11282), .ZN(
        n11284) );
  MUX2_X1 U13752 ( .A(n11285), .B(n14260), .S(n11554), .Z(n11286) );
  INV_X1 U13753 ( .A(n14397), .ZN(n14426) );
  OAI21_X1 U13754 ( .B1(n14426), .B2(n13656), .A(n11298), .ZN(n11293) );
  OR2_X1 U13755 ( .A1(n14394), .A2(n11551), .ZN(n11289) );
  OAI21_X1 U13756 ( .B1(n14432), .B2(n11554), .A(n11289), .ZN(n11290) );
  NOR2_X1 U13757 ( .A1(n11291), .A2(n11290), .ZN(n11292) );
  AOI22_X1 U13758 ( .A1(n11293), .A2(n11551), .B1(n11292), .B2(n14391), .ZN(
        n11294) );
  AOI21_X1 U13759 ( .B1(n11297), .B2(n11295), .A(n11551), .ZN(n11296) );
  MUX2_X1 U13760 ( .A(n13655), .B(n14409), .S(n11554), .Z(n11299) );
  OR2_X1 U13761 ( .A1(n11300), .A2(n11299), .ZN(n11304) );
  NAND2_X1 U13762 ( .A1(n11300), .A2(n11299), .ZN(n11302) );
  MUX2_X1 U13763 ( .A(n13655), .B(n14409), .S(n11551), .Z(n11301) );
  NAND2_X1 U13764 ( .A1(n11302), .A2(n11301), .ZN(n11303) );
  NAND2_X1 U13765 ( .A1(n11304), .A2(n11303), .ZN(n11321) );
  NAND2_X1 U13766 ( .A1(n11305), .A2(n11547), .ZN(n11308) );
  AOI22_X1 U13767 ( .A1(n11548), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(n11317), 
        .B2(n11306), .ZN(n11307) );
  NAND2_X1 U13768 ( .A1(n14090), .A2(n13977), .ZN(n11909) );
  NAND2_X1 U13769 ( .A1(n11309), .A2(n11547), .ZN(n11311) );
  AOI22_X1 U13770 ( .A1(n11548), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n11204), 
        .B2(n11317), .ZN(n11310) );
  OR2_X1 U13771 ( .A1(n11312), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n11313) );
  NAND2_X1 U13772 ( .A1(n11332), .A2(n11313), .ZN(n13966) );
  AOI22_X1 U13773 ( .A1(n6473), .A2(P1_REG1_REG_19__SCAN_IN), .B1(n6482), .B2(
        P1_REG2_REG_19__SCAN_IN), .ZN(n11315) );
  NAND2_X1 U13774 ( .A1(n11503), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n11314) );
  OAI211_X1 U13775 ( .C1(n13966), .C2(n6468), .A(n11315), .B(n11314), .ZN(
        n13978) );
  XNOR2_X1 U13776 ( .A(n13969), .B(n13978), .ZN(n11574) );
  NAND2_X1 U13777 ( .A1(n11316), .A2(n9599), .ZN(n11319) );
  AOI22_X1 U13778 ( .A1(n11548), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(n11317), 
        .B2(n13797), .ZN(n11318) );
  XNOR2_X1 U13779 ( .A(n13987), .B(n13530), .ZN(n13975) );
  NOR2_X1 U13780 ( .A1(n14090), .A2(n13977), .ZN(n11910) );
  MUX2_X1 U13781 ( .A(n13977), .B(n14090), .S(n11551), .Z(n11320) );
  INV_X1 U13782 ( .A(n13530), .ZN(n14009) );
  NAND3_X1 U13783 ( .A1(n13987), .A2(n14009), .A3(n11551), .ZN(n11323) );
  OR3_X1 U13784 ( .A1(n13987), .A2(n14009), .A3(n11551), .ZN(n11322) );
  NAND2_X1 U13785 ( .A1(n11323), .A2(n11322), .ZN(n11324) );
  NAND2_X1 U13786 ( .A1(n11574), .A2(n11324), .ZN(n11328) );
  NAND2_X1 U13787 ( .A1(n13969), .A2(n11551), .ZN(n11326) );
  OR2_X1 U13788 ( .A1(n13969), .A2(n11551), .ZN(n11325) );
  MUX2_X1 U13789 ( .A(n11326), .B(n11325), .S(n13978), .Z(n11327) );
  NAND2_X1 U13790 ( .A1(n11639), .A2(n9599), .ZN(n11330) );
  NAND2_X1 U13791 ( .A1(n11548), .A2(P2_DATAO_REG_20__SCAN_IN), .ZN(n11329) );
  INV_X1 U13792 ( .A(P1_REG3_REG_20__SCAN_IN), .ZN(n11331) );
  NAND2_X1 U13793 ( .A1(n11332), .A2(n11331), .ZN(n11333) );
  AND2_X1 U13794 ( .A1(n11344), .A2(n11333), .ZN(n13953) );
  INV_X1 U13795 ( .A(n6476), .ZN(n11380) );
  NAND2_X1 U13796 ( .A1(n13953), .A2(n11380), .ZN(n11339) );
  INV_X1 U13797 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n11336) );
  NAND2_X1 U13798 ( .A1(n6482), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n11335) );
  NAND2_X1 U13799 ( .A1(n11503), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n11334) );
  OAI211_X1 U13800 ( .C1(n6483), .C2(n11336), .A(n11335), .B(n11334), .ZN(
        n11337) );
  INV_X1 U13801 ( .A(n11337), .ZN(n11338) );
  NAND2_X1 U13802 ( .A1(n11339), .A2(n11338), .ZN(n13935) );
  MUX2_X1 U13803 ( .A(n14078), .B(n13935), .S(n11551), .Z(n11340) );
  INV_X1 U13804 ( .A(n11340), .ZN(n11342) );
  MUX2_X1 U13805 ( .A(n13935), .B(n14078), .S(n11551), .Z(n11341) );
  INV_X1 U13806 ( .A(P1_REG3_REG_21__SCAN_IN), .ZN(n11343) );
  AND2_X1 U13807 ( .A1(n11344), .A2(n11343), .ZN(n11345) );
  OR2_X1 U13808 ( .A1(n11345), .A2(n11365), .ZN(n13930) );
  INV_X1 U13809 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n11348) );
  NAND2_X1 U13810 ( .A1(n11503), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n11347) );
  NAND2_X1 U13811 ( .A1(n6482), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n11346) );
  OAI211_X1 U13812 ( .C1(n6483), .C2(n11348), .A(n11347), .B(n11346), .ZN(
        n11349) );
  INV_X1 U13813 ( .A(n11349), .ZN(n11350) );
  OAI21_X1 U13814 ( .B1(n13930), .B2(n6468), .A(n11350), .ZN(n13945) );
  NAND2_X1 U13815 ( .A1(n11646), .A2(n9599), .ZN(n11352) );
  NAND2_X1 U13816 ( .A1(n11548), .A2(P2_DATAO_REG_21__SCAN_IN), .ZN(n11351) );
  MUX2_X1 U13817 ( .A(n13945), .B(n14072), .S(n11551), .Z(n11356) );
  NAND2_X1 U13818 ( .A1(n11355), .A2(n11356), .ZN(n11354) );
  MUX2_X1 U13819 ( .A(n14072), .B(n13945), .S(n11551), .Z(n11353) );
  NAND2_X1 U13820 ( .A1(n11354), .A2(n11353), .ZN(n11360) );
  INV_X1 U13821 ( .A(n11355), .ZN(n11358) );
  INV_X1 U13822 ( .A(n11356), .ZN(n11357) );
  NAND2_X1 U13823 ( .A1(n11358), .A2(n11357), .ZN(n11359) );
  NAND2_X1 U13824 ( .A1(n11360), .A2(n11359), .ZN(n11376) );
  NAND2_X1 U13825 ( .A1(n11362), .A2(n11361), .ZN(n11363) );
  NOR2_X1 U13826 ( .A1(n11365), .A2(P1_REG3_REG_22__SCAN_IN), .ZN(n11366) );
  NOR2_X1 U13827 ( .A1(n11378), .A2(n11366), .ZN(n13923) );
  NAND2_X1 U13828 ( .A1(n13923), .A2(n11380), .ZN(n11372) );
  INV_X1 U13829 ( .A(P1_REG1_REG_22__SCAN_IN), .ZN(n11369) );
  NAND2_X1 U13830 ( .A1(n11503), .A2(P1_REG0_REG_22__SCAN_IN), .ZN(n11368) );
  NAND2_X1 U13831 ( .A1(n6482), .A2(P1_REG2_REG_22__SCAN_IN), .ZN(n11367) );
  OAI211_X1 U13832 ( .C1(n6483), .C2(n11369), .A(n11368), .B(n11367), .ZN(
        n11370) );
  INV_X1 U13833 ( .A(n11370), .ZN(n11371) );
  MUX2_X1 U13834 ( .A(n11572), .B(n11917), .S(n11551), .Z(n11373) );
  INV_X1 U13835 ( .A(n11373), .ZN(n11375) );
  MUX2_X1 U13836 ( .A(n11917), .B(n11572), .S(n11551), .Z(n11374) );
  NOR2_X1 U13837 ( .A1(n11376), .A2(n11375), .ZN(n11377) );
  OR2_X1 U13838 ( .A1(n11378), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n11379) );
  AND2_X1 U13839 ( .A1(n11379), .A2(n11395), .ZN(n13906) );
  NAND2_X1 U13840 ( .A1(n13906), .A2(n11380), .ZN(n11386) );
  INV_X1 U13841 ( .A(P1_REG1_REG_23__SCAN_IN), .ZN(n11383) );
  NAND2_X1 U13842 ( .A1(n11503), .A2(P1_REG0_REG_23__SCAN_IN), .ZN(n11382) );
  NAND2_X1 U13843 ( .A1(n6482), .A2(P1_REG2_REG_23__SCAN_IN), .ZN(n11381) );
  OAI211_X1 U13844 ( .C1(n6483), .C2(n11383), .A(n11382), .B(n11381), .ZN(
        n11384) );
  INV_X1 U13845 ( .A(n11384), .ZN(n11385) );
  NAND2_X1 U13846 ( .A1(n11386), .A2(n11385), .ZN(n13888) );
  NAND2_X1 U13847 ( .A1(n11387), .A2(n11547), .ZN(n11389) );
  NAND2_X1 U13848 ( .A1(n11548), .A2(P2_DATAO_REG_23__SCAN_IN), .ZN(n11388) );
  MUX2_X1 U13849 ( .A(n13888), .B(n14062), .S(n11551), .Z(n11391) );
  MUX2_X1 U13850 ( .A(n14062), .B(n13888), .S(n11551), .Z(n11390) );
  NAND2_X1 U13851 ( .A1(n11548), .A2(P2_DATAO_REG_24__SCAN_IN), .ZN(n11392) );
  NAND2_X1 U13852 ( .A1(n6482), .A2(P1_REG2_REG_24__SCAN_IN), .ZN(n11401) );
  INV_X1 U13853 ( .A(P1_REG1_REG_24__SCAN_IN), .ZN(n11394) );
  OR2_X1 U13854 ( .A1(n9593), .A2(n11394), .ZN(n11400) );
  OAI21_X1 U13855 ( .B1(P1_REG3_REG_24__SCAN_IN), .B2(n11396), .A(n11413), 
        .ZN(n13895) );
  OR2_X1 U13856 ( .A1(n6468), .A2(n13895), .ZN(n11399) );
  INV_X1 U13857 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n11397) );
  OR2_X1 U13858 ( .A1(n11516), .A2(n11397), .ZN(n11398) );
  NAND4_X1 U13859 ( .A1(n11401), .A2(n11400), .A3(n11399), .A4(n11398), .ZN(
        n13865) );
  MUX2_X1 U13860 ( .A(n13898), .B(n13865), .S(n11551), .Z(n11405) );
  NAND2_X1 U13861 ( .A1(n11404), .A2(n11405), .ZN(n11403) );
  MUX2_X1 U13862 ( .A(n13865), .B(n13898), .S(n11551), .Z(n11402) );
  NAND2_X1 U13863 ( .A1(n11403), .A2(n11402), .ZN(n11409) );
  INV_X1 U13864 ( .A(n11405), .ZN(n11406) );
  NAND2_X1 U13865 ( .A1(n11407), .A2(n11406), .ZN(n11408) );
  NAND2_X1 U13866 ( .A1(n6482), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n11419) );
  INV_X1 U13867 ( .A(P1_REG1_REG_25__SCAN_IN), .ZN(n11410) );
  OR2_X1 U13868 ( .A1(n6483), .A2(n11410), .ZN(n11418) );
  INV_X1 U13869 ( .A(n11413), .ZN(n11411) );
  NAND2_X1 U13870 ( .A1(n11411), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n11435) );
  INV_X1 U13871 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n11412) );
  NAND2_X1 U13872 ( .A1(n11413), .A2(n11412), .ZN(n11414) );
  NAND2_X1 U13873 ( .A1(n11435), .A2(n11414), .ZN(n13869) );
  OR2_X1 U13874 ( .A1(n11470), .A2(n13869), .ZN(n11417) );
  INV_X1 U13875 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n11415) );
  OR2_X1 U13876 ( .A1(n11516), .A2(n11415), .ZN(n11416) );
  NAND4_X1 U13877 ( .A1(n11419), .A2(n11418), .A3(n11417), .A4(n11416), .ZN(
        n13887) );
  XNOR2_X1 U13878 ( .A(n11421), .B(n11420), .ZN(n13436) );
  NAND2_X1 U13879 ( .A1(n13436), .A2(n11547), .ZN(n11423) );
  NAND2_X1 U13880 ( .A1(n11548), .A2(P2_DATAO_REG_25__SCAN_IN), .ZN(n11422) );
  MUX2_X1 U13881 ( .A(n13887), .B(n14049), .S(n11551), .Z(n11426) );
  MUX2_X1 U13882 ( .A(n13887), .B(n14049), .S(n11554), .Z(n11424) );
  INV_X1 U13883 ( .A(n11426), .ZN(n11427) );
  NAND2_X1 U13884 ( .A1(n11172), .A2(n11428), .ZN(n11429) );
  NAND2_X1 U13885 ( .A1(n13434), .A2(n9599), .ZN(n11432) );
  NAND2_X1 U13886 ( .A1(n11548), .A2(P2_DATAO_REG_26__SCAN_IN), .ZN(n11431) );
  NAND2_X1 U13887 ( .A1(n6473), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n11441) );
  INV_X1 U13888 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n13853) );
  OR2_X1 U13889 ( .A1(n6487), .A2(n13853), .ZN(n11440) );
  INV_X1 U13890 ( .A(n11435), .ZN(n11433) );
  NAND2_X1 U13891 ( .A1(n11433), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n11450) );
  INV_X1 U13892 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n11434) );
  NAND2_X1 U13893 ( .A1(n11435), .A2(n11434), .ZN(n11436) );
  NAND2_X1 U13894 ( .A1(n11450), .A2(n11436), .ZN(n13849) );
  OR2_X1 U13895 ( .A1(n11470), .A2(n13849), .ZN(n11439) );
  INV_X1 U13896 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n11437) );
  OR2_X1 U13897 ( .A1(n11516), .A2(n11437), .ZN(n11438) );
  NAND4_X1 U13898 ( .A1(n11441), .A2(n11440), .A3(n11439), .A4(n11438), .ZN(
        n13866) );
  MUX2_X1 U13899 ( .A(n14043), .B(n13866), .S(n11551), .Z(n11444) );
  MUX2_X1 U13900 ( .A(n13866), .B(n14043), .S(n11551), .Z(n11442) );
  NAND2_X1 U13901 ( .A1(n11443), .A2(n11442), .ZN(n11446) );
  NAND2_X1 U13902 ( .A1(n6473), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n11456) );
  INV_X1 U13903 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n13837) );
  OR2_X1 U13904 ( .A1(n6487), .A2(n13837), .ZN(n11455) );
  INV_X1 U13905 ( .A(n11450), .ZN(n11448) );
  NAND2_X1 U13906 ( .A1(n11448), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n11513) );
  INV_X1 U13907 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n11449) );
  NAND2_X1 U13908 ( .A1(n11450), .A2(n11449), .ZN(n11451) );
  NAND2_X1 U13909 ( .A1(n11513), .A2(n11451), .ZN(n13836) );
  OR2_X1 U13910 ( .A1(n6468), .A2(n13836), .ZN(n11454) );
  INV_X1 U13911 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n11452) );
  OR2_X1 U13912 ( .A1(n11516), .A2(n11452), .ZN(n11453) );
  XNOR2_X1 U13913 ( .A(n11458), .B(SI_27_), .ZN(n11459) );
  NAND2_X1 U13914 ( .A1(n13431), .A2(n9599), .ZN(n11461) );
  NAND2_X1 U13915 ( .A1(n11548), .A2(P2_DATAO_REG_27__SCAN_IN), .ZN(n11460) );
  MUX2_X1 U13916 ( .A(n13847), .B(n14038), .S(n11551), .Z(n11465) );
  NAND2_X1 U13917 ( .A1(n11464), .A2(n11465), .ZN(n11463) );
  MUX2_X1 U13918 ( .A(n14038), .B(n13847), .S(n11551), .Z(n11462) );
  INV_X1 U13919 ( .A(n11464), .ZN(n11467) );
  INV_X1 U13920 ( .A(n11465), .ZN(n11466) );
  NAND2_X1 U13921 ( .A1(n6473), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n11475) );
  INV_X1 U13922 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n11468) );
  OR2_X1 U13923 ( .A1(n6487), .A2(n11468), .ZN(n11474) );
  INV_X1 U13924 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n11469) );
  XNOR2_X1 U13925 ( .A(n11513), .B(n11469), .ZN(n13546) );
  INV_X1 U13926 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n11471) );
  OR2_X1 U13927 ( .A1(n11516), .A2(n11471), .ZN(n11472) );
  NAND4_X1 U13928 ( .A1(n11475), .A2(n11474), .A3(n11473), .A4(n11472), .ZN(
        n13654) );
  NAND2_X1 U13929 ( .A1(n11737), .A2(n11547), .ZN(n11479) );
  NAND2_X1 U13930 ( .A1(n11548), .A2(P2_DATAO_REG_28__SCAN_IN), .ZN(n11478) );
  MUX2_X1 U13931 ( .A(n13654), .B(n14032), .S(n11554), .Z(n11525) );
  INV_X1 U13932 ( .A(n11482), .ZN(n11484) );
  NAND2_X1 U13933 ( .A1(n11484), .A2(n11483), .ZN(n11485) );
  MUX2_X1 U13934 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(P1_DATAO_REG_30__SCAN_IN), 
        .S(n11543), .Z(n11486) );
  NAND2_X1 U13935 ( .A1(n11486), .A2(SI_30_), .ZN(n11541) );
  OAI21_X1 U13936 ( .B1(SI_30_), .B2(n11486), .A(n11541), .ZN(n11488) );
  NAND2_X1 U13937 ( .A1(n11487), .A2(n11488), .ZN(n11489) );
  NAND2_X1 U13938 ( .A1(n11548), .A2(P2_DATAO_REG_30__SCAN_IN), .ZN(n11491) );
  INV_X1 U13939 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n11493) );
  NOR2_X1 U13940 ( .A1(n9593), .A2(n11493), .ZN(n11498) );
  INV_X1 U13941 ( .A(P1_REG2_REG_31__SCAN_IN), .ZN(n11494) );
  NOR2_X1 U13942 ( .A1(n6487), .A2(n11494), .ZN(n11497) );
  INV_X1 U13943 ( .A(P1_REG0_REG_31__SCAN_IN), .ZN(n11495) );
  NOR2_X1 U13944 ( .A1(n11516), .A2(n11495), .ZN(n11496) );
  NAND2_X1 U13945 ( .A1(n13814), .A2(n11551), .ZN(n11501) );
  NAND2_X1 U13946 ( .A1(n11499), .A2(n7146), .ZN(n11500) );
  NAND2_X1 U13947 ( .A1(n11501), .A2(n11500), .ZN(n11507) );
  INV_X1 U13948 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n11506) );
  NAND2_X1 U13949 ( .A1(n6482), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n11505) );
  NAND2_X1 U13950 ( .A1(n11503), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n11504) );
  OAI211_X1 U13951 ( .C1(n9593), .C2(n11506), .A(n11505), .B(n11504), .ZN(
        n13652) );
  AND2_X1 U13952 ( .A1(n11507), .A2(n13652), .ZN(n11508) );
  AOI21_X1 U13953 ( .B1(n13818), .B2(n11554), .A(n11508), .ZN(n11532) );
  OAI21_X1 U13954 ( .B1(n13814), .B2(n11509), .A(n13652), .ZN(n11510) );
  INV_X1 U13955 ( .A(n11510), .ZN(n11511) );
  MUX2_X1 U13956 ( .A(n11511), .B(n13818), .S(n11551), .Z(n11526) );
  NAND2_X1 U13957 ( .A1(n6473), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n11520) );
  INV_X1 U13958 ( .A(P1_REG2_REG_29__SCAN_IN), .ZN(n11512) );
  OR2_X1 U13959 ( .A1(n6487), .A2(n11512), .ZN(n11519) );
  INV_X1 U13960 ( .A(n11513), .ZN(n11514) );
  NAND2_X1 U13961 ( .A1(n11514), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n12003) );
  OR2_X1 U13962 ( .A1(n6468), .A2(n12003), .ZN(n11518) );
  INV_X1 U13963 ( .A(P1_REG0_REG_29__SCAN_IN), .ZN(n11515) );
  OR2_X1 U13964 ( .A1(n11516), .A2(n11515), .ZN(n11517) );
  NAND2_X1 U13965 ( .A1(n11861), .A2(n9599), .ZN(n11522) );
  NAND2_X1 U13966 ( .A1(n11548), .A2(P2_DATAO_REG_29__SCAN_IN), .ZN(n11521) );
  MUX2_X1 U13967 ( .A(n11569), .B(n14027), .S(n11554), .Z(n11528) );
  MUX2_X1 U13968 ( .A(n13653), .B(n11570), .S(n11551), .Z(n11527) );
  AOI22_X1 U13969 ( .A1(n11532), .A2(n11526), .B1(n11528), .B2(n11527), .ZN(
        n11523) );
  INV_X1 U13970 ( .A(n13654), .ZN(n13829) );
  INV_X1 U13971 ( .A(n14032), .ZN(n13540) );
  MUX2_X1 U13972 ( .A(n13829), .B(n13540), .S(n11551), .Z(n11524) );
  INV_X1 U13973 ( .A(n11526), .ZN(n11536) );
  INV_X1 U13974 ( .A(n11527), .ZN(n11530) );
  INV_X1 U13975 ( .A(n11528), .ZN(n11529) );
  NAND2_X1 U13976 ( .A1(n11530), .A2(n11529), .ZN(n11531) );
  NAND2_X1 U13977 ( .A1(n11532), .A2(n11531), .ZN(n11535) );
  INV_X1 U13978 ( .A(n11531), .ZN(n11534) );
  INV_X1 U13979 ( .A(n11532), .ZN(n11533) );
  AOI22_X1 U13980 ( .A1(n11536), .A2(n11535), .B1(n11534), .B2(n11533), .ZN(
        n11537) );
  NAND2_X1 U13981 ( .A1(n11538), .A2(n9666), .ZN(n11540) );
  NAND2_X1 U13982 ( .A1(n11540), .A2(n11539), .ZN(n11556) );
  INV_X1 U13983 ( .A(n11556), .ZN(n11555) );
  MUX2_X1 U13984 ( .A(P2_DATAO_REG_31__SCAN_IN), .B(P1_DATAO_REG_31__SCAN_IN), 
        .S(n11543), .Z(n11544) );
  XNOR2_X1 U13985 ( .A(n11544), .B(SI_31_), .ZN(n11545) );
  NAND2_X1 U13986 ( .A1(n12944), .A2(n11547), .ZN(n11550) );
  NAND2_X1 U13987 ( .A1(n11548), .A2(P2_DATAO_REG_31__SCAN_IN), .ZN(n11549) );
  XNOR2_X1 U13988 ( .A(n13812), .B(n13814), .ZN(n11568) );
  OR2_X1 U13989 ( .A1(n13812), .A2(n11551), .ZN(n11562) );
  INV_X1 U13990 ( .A(n11562), .ZN(n11552) );
  XOR2_X1 U13991 ( .A(n11556), .B(n11552), .Z(n11553) );
  NAND4_X1 U13992 ( .A1(n11553), .A2(n14018), .A3(n11605), .A4(n13814), .ZN(
        n11560) );
  NOR2_X1 U13993 ( .A1(n14018), .A2(n11554), .ZN(n11565) );
  INV_X1 U13994 ( .A(n13814), .ZN(n11564) );
  NAND3_X1 U13995 ( .A1(n11565), .A2(n11564), .A3(n11555), .ZN(n11559) );
  INV_X1 U13996 ( .A(n11565), .ZN(n11557) );
  AND2_X1 U13997 ( .A1(n11556), .A2(n11605), .ZN(n11561) );
  NAND4_X1 U13998 ( .A1(n11557), .A2(n11564), .A3(n11561), .A4(n13812), .ZN(
        n11558) );
  OAI21_X1 U13999 ( .B1(n11562), .B2(n11564), .A(n11561), .ZN(n11563) );
  INV_X1 U14000 ( .A(n11568), .ZN(n11603) );
  XNOR2_X1 U14001 ( .A(n13818), .B(n13652), .ZN(n11601) );
  INV_X1 U14002 ( .A(n14043), .ZN(n13854) );
  NAND2_X1 U14003 ( .A1(n13854), .A2(n13866), .ZN(n11571) );
  INV_X1 U14004 ( .A(n13866), .ZN(n13830) );
  NAND2_X1 U14005 ( .A1(n14043), .A2(n13830), .ZN(n13825) );
  INV_X1 U14006 ( .A(n13888), .ZN(n13918) );
  XNOR2_X1 U14007 ( .A(n13898), .B(n13865), .ZN(n13885) );
  INV_X1 U14008 ( .A(n14078), .ZN(n11816) );
  NAND2_X1 U14009 ( .A1(n11816), .A2(n13935), .ZN(n11897) );
  INV_X1 U14010 ( .A(n13935), .ZN(n13964) );
  NAND2_X1 U14011 ( .A1(n14078), .A2(n13964), .ZN(n11573) );
  NAND2_X1 U14012 ( .A1(n11897), .A2(n11573), .ZN(n13949) );
  INV_X1 U14013 ( .A(n13975), .ZN(n11596) );
  NAND4_X1 U14014 ( .A1(n11577), .A2(n14521), .A3(n14540), .A4(n11576), .ZN(
        n11579) );
  NOR2_X1 U14015 ( .A1(n11579), .A2(n11578), .ZN(n11583) );
  NAND4_X1 U14016 ( .A1(n11583), .A2(n11582), .A3(n11581), .A4(n11580), .ZN(
        n11584) );
  NOR2_X1 U14017 ( .A1(n11585), .A2(n11584), .ZN(n11588) );
  NAND4_X1 U14018 ( .A1(n11589), .A2(n11588), .A3(n11587), .A4(n11586), .ZN(
        n11590) );
  OR4_X1 U14019 ( .A1(n11593), .A2(n11592), .A3(n11591), .A4(n11590), .ZN(
        n11595) );
  NAND2_X1 U14020 ( .A1(n7120), .A2(n11909), .ZN(n14001) );
  NAND2_X1 U14021 ( .A1(n14001), .A2(n14391), .ZN(n11594) );
  OR4_X1 U14022 ( .A1(n11596), .A2(n11905), .A3(n11595), .A4(n11594), .ZN(
        n11597) );
  NOR3_X1 U14023 ( .A1(n13949), .A2(n13962), .A3(n11597), .ZN(n11598) );
  XNOR2_X1 U14024 ( .A(n14072), .B(n13945), .ZN(n13934) );
  NAND4_X1 U14025 ( .A1(n13885), .A2(n11916), .A3(n11598), .A4(n13934), .ZN(
        n11599) );
  NOR4_X1 U14026 ( .A1(n13842), .A2(n13860), .A3(n13903), .A4(n11599), .ZN(
        n11600) );
  NAND4_X1 U14027 ( .A1(n11601), .A2(n11600), .A3(n11923), .A4(n11921), .ZN(
        n11602) );
  XNOR2_X1 U14028 ( .A(n11604), .B(n13806), .ZN(n11607) );
  INV_X1 U14029 ( .A(n11605), .ZN(n11606) );
  NAND2_X1 U14030 ( .A1(n11607), .A2(n11606), .ZN(n11608) );
  OAI21_X1 U14031 ( .B1(n11610), .B2(n11609), .A(n11608), .ZN(n11611) );
  NOR2_X1 U14032 ( .A1(n11612), .A2(n11611), .ZN(n11617) );
  NOR3_X1 U14033 ( .A1(n11613), .A2(n14121), .A3(n14006), .ZN(n11615) );
  OAI21_X1 U14034 ( .B1(n11616), .B2(n14544), .A(P1_B_REG_SCAN_IN), .ZN(n11614) );
  INV_X1 U14035 ( .A(n11737), .ZN(n13430) );
  OAI222_X1 U14036 ( .A1(n14124), .A2(n11618), .B1(n14130), .B2(n13430), .C1(
        P1_U3086), .C2(n8743), .ZN(P1_U3327) );
  NAND2_X1 U14037 ( .A1(n11387), .A2(n12943), .ZN(n11620) );
  NAND2_X1 U14038 ( .A1(n11862), .A2(P1_DATAO_REG_23__SCAN_IN), .ZN(n11619) );
  INV_X1 U14039 ( .A(n13363), .ZN(n11879) );
  XNOR2_X1 U14040 ( .A(n11879), .B(n11750), .ZN(n12619) );
  INV_X1 U14041 ( .A(n12619), .ZN(n11684) );
  XNOR2_X1 U14042 ( .A(n13404), .B(n11628), .ZN(n11625) );
  NAND2_X1 U14043 ( .A1(n13052), .A2(n11749), .ZN(n11624) );
  NAND2_X1 U14044 ( .A1(n11625), .A2(n11624), .ZN(n11626) );
  OAI21_X1 U14045 ( .B1(n11625), .B2(n11624), .A(n11626), .ZN(n12654) );
  INV_X1 U14046 ( .A(n11626), .ZN(n11627) );
  NOR2_X1 U14047 ( .A1(n12652), .A2(n11627), .ZN(n12664) );
  XNOR2_X1 U14048 ( .A(n12851), .B(n11628), .ZN(n11630) );
  NAND2_X1 U14049 ( .A1(n13051), .A2(n11749), .ZN(n11629) );
  NAND2_X1 U14050 ( .A1(n11630), .A2(n11629), .ZN(n11631) );
  OAI21_X1 U14051 ( .B1(n11630), .B2(n11629), .A(n11631), .ZN(n12663) );
  NOR2_X2 U14052 ( .A1(n12664), .A2(n12663), .ZN(n12662) );
  INV_X1 U14053 ( .A(n11631), .ZN(n11632) );
  XNOR2_X1 U14054 ( .A(n13390), .B(n11750), .ZN(n11634) );
  NAND2_X1 U14055 ( .A1(n13050), .A2(n11749), .ZN(n11633) );
  XNOR2_X1 U14056 ( .A(n11634), .B(n11633), .ZN(n12698) );
  INV_X1 U14057 ( .A(n11633), .ZN(n11635) );
  AND2_X1 U14058 ( .A1(n13049), .A2(n11749), .ZN(n11637) );
  XNOR2_X1 U14059 ( .A(n12873), .B(n11750), .ZN(n11636) );
  NOR2_X1 U14060 ( .A1(n11636), .A2(n11637), .ZN(n11638) );
  AOI21_X1 U14061 ( .B1(n11637), .B2(n11636), .A(n11638), .ZN(n12629) );
  AND2_X1 U14062 ( .A1(n13048), .A2(n11749), .ZN(n11643) );
  NAND2_X1 U14063 ( .A1(n11639), .A2(n11860), .ZN(n11641) );
  NAND2_X1 U14064 ( .A1(n11862), .A2(P1_DATAO_REG_20__SCAN_IN), .ZN(n11640) );
  XNOR2_X1 U14065 ( .A(n13380), .B(n11750), .ZN(n11642) );
  NOR2_X1 U14066 ( .A1(n11642), .A2(n11643), .ZN(n11644) );
  AOI21_X1 U14067 ( .B1(n11643), .B2(n11642), .A(n11644), .ZN(n12681) );
  NAND2_X1 U14068 ( .A1(n12680), .A2(n12681), .ZN(n12679) );
  INV_X1 U14069 ( .A(n11644), .ZN(n11645) );
  NAND2_X1 U14070 ( .A1(n11646), .A2(n12943), .ZN(n11648) );
  NAND2_X1 U14071 ( .A1(n11862), .A2(P1_DATAO_REG_21__SCAN_IN), .ZN(n11647) );
  XNOR2_X1 U14072 ( .A(n13374), .B(n11750), .ZN(n11658) );
  OR2_X1 U14073 ( .A1(n11649), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n11650) );
  NAND2_X1 U14074 ( .A1(n11649), .A2(P2_REG3_REG_21__SCAN_IN), .ZN(n11665) );
  AND2_X1 U14075 ( .A1(n11650), .A2(n11665), .ZN(n12638) );
  NAND2_X1 U14076 ( .A1(n12638), .A2(n6485), .ZN(n11656) );
  INV_X1 U14077 ( .A(P2_REG1_REG_21__SCAN_IN), .ZN(n11653) );
  NAND2_X1 U14078 ( .A1(n11123), .A2(P2_REG0_REG_21__SCAN_IN), .ZN(n11652) );
  NAND2_X1 U14079 ( .A1(n11688), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n11651) );
  OAI211_X1 U14080 ( .C1(n11872), .C2(n11653), .A(n11652), .B(n11651), .ZN(
        n11654) );
  INV_X1 U14081 ( .A(n11654), .ZN(n11655) );
  NAND2_X1 U14082 ( .A1(n11656), .A2(n11655), .ZN(n13047) );
  NAND2_X1 U14083 ( .A1(n13047), .A2(n11749), .ZN(n11657) );
  XNOR2_X1 U14084 ( .A(n11658), .B(n11657), .ZN(n12636) );
  NAND2_X1 U14085 ( .A1(n11659), .A2(n11860), .ZN(n11661) );
  NAND2_X1 U14086 ( .A1(n11862), .A2(P1_DATAO_REG_22__SCAN_IN), .ZN(n11660) );
  XNOR2_X1 U14087 ( .A(n13368), .B(n11750), .ZN(n11672) );
  NAND2_X1 U14088 ( .A1(n11123), .A2(P2_REG0_REG_22__SCAN_IN), .ZN(n11671) );
  NAND2_X1 U14089 ( .A1(n11701), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n11670) );
  INV_X1 U14090 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n11664) );
  NAND2_X1 U14091 ( .A1(n11664), .A2(n11665), .ZN(n11667) );
  INV_X1 U14092 ( .A(n11665), .ZN(n11666) );
  NAND2_X1 U14093 ( .A1(P2_REG3_REG_22__SCAN_IN), .A2(n11666), .ZN(n11676) );
  AND2_X1 U14094 ( .A1(n11667), .A2(n11676), .ZN(n13265) );
  NAND2_X1 U14095 ( .A1(n9145), .A2(n13265), .ZN(n11669) );
  NAND2_X1 U14096 ( .A1(n11688), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n11668) );
  NAND4_X1 U14097 ( .A1(n11671), .A2(n11670), .A3(n11669), .A4(n11668), .ZN(
        n13046) );
  INV_X1 U14098 ( .A(n13046), .ZN(n12898) );
  NOR2_X1 U14099 ( .A1(n12898), .A2(n9335), .ZN(n12689) );
  INV_X1 U14100 ( .A(n12621), .ZN(n11683) );
  NAND2_X1 U14101 ( .A1(n11123), .A2(P2_REG0_REG_23__SCAN_IN), .ZN(n11681) );
  NAND2_X1 U14102 ( .A1(n9113), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n11680) );
  INV_X1 U14103 ( .A(n11676), .ZN(n11674) );
  NAND2_X1 U14104 ( .A1(n11674), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n11691) );
  INV_X1 U14105 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n11675) );
  NAND2_X1 U14106 ( .A1(n11676), .A2(n11675), .ZN(n11677) );
  AND2_X1 U14107 ( .A1(n11691), .A2(n11677), .ZN(n12622) );
  NAND2_X1 U14108 ( .A1(n9145), .A2(n12622), .ZN(n11679) );
  NAND2_X1 U14109 ( .A1(n11688), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n11678) );
  NAND4_X1 U14110 ( .A1(n11681), .A2(n11680), .A3(n11679), .A4(n11678), .ZN(
        n13045) );
  NAND2_X1 U14111 ( .A1(n13045), .A2(n11749), .ZN(n12618) );
  AOI21_X1 U14112 ( .B1(n12621), .B2(n12619), .A(n12618), .ZN(n11682) );
  NAND2_X1 U14113 ( .A1(n11862), .A2(P1_DATAO_REG_24__SCAN_IN), .ZN(n11686) );
  XNOR2_X1 U14114 ( .A(n13236), .B(n11750), .ZN(n11698) );
  NAND2_X1 U14115 ( .A1(n11701), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n11696) );
  NAND2_X1 U14116 ( .A1(n11688), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n11695) );
  INV_X1 U14117 ( .A(n11691), .ZN(n11689) );
  NAND2_X1 U14118 ( .A1(n11689), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n11704) );
  INV_X1 U14119 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n11690) );
  NAND2_X1 U14120 ( .A1(n11691), .A2(n11690), .ZN(n11692) );
  AND2_X1 U14121 ( .A1(n11704), .A2(n11692), .ZN(n12673) );
  NAND2_X1 U14122 ( .A1(n9145), .A2(n12673), .ZN(n11694) );
  NAND2_X1 U14123 ( .A1(n11123), .A2(P2_REG0_REG_24__SCAN_IN), .ZN(n11693) );
  NAND4_X1 U14124 ( .A1(n11696), .A2(n11695), .A3(n11694), .A4(n11693), .ZN(
        n13044) );
  NAND2_X1 U14125 ( .A1(n13044), .A2(n11749), .ZN(n11697) );
  XNOR2_X1 U14126 ( .A(n11698), .B(n11697), .ZN(n12671) );
  OAI22_X2 U14127 ( .A1(n12672), .A2(n12671), .B1(n11698), .B2(n11697), .ZN(
        n12644) );
  NAND2_X1 U14128 ( .A1(n13436), .A2(n11860), .ZN(n11700) );
  NAND2_X1 U14129 ( .A1(n11862), .A2(P1_DATAO_REG_25__SCAN_IN), .ZN(n11699) );
  XNOR2_X1 U14130 ( .A(n13352), .B(n11750), .ZN(n11712) );
  NAND2_X1 U14131 ( .A1(n11701), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n11709) );
  NAND2_X1 U14132 ( .A1(n11688), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n11708) );
  INV_X1 U14133 ( .A(n11704), .ZN(n11702) );
  NAND2_X1 U14134 ( .A1(n11702), .A2(P2_REG3_REG_25__SCAN_IN), .ZN(n11714) );
  INV_X1 U14135 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n11703) );
  NAND2_X1 U14136 ( .A1(n11704), .A2(n11703), .ZN(n11705) );
  AND2_X1 U14137 ( .A1(n11714), .A2(n11705), .ZN(n13216) );
  NAND2_X1 U14138 ( .A1(n9145), .A2(n13216), .ZN(n11707) );
  NAND2_X1 U14139 ( .A1(n11123), .A2(P2_REG0_REG_25__SCAN_IN), .ZN(n11706) );
  NAND4_X1 U14140 ( .A1(n11709), .A2(n11708), .A3(n11707), .A4(n11706), .ZN(
        n13043) );
  NAND2_X1 U14141 ( .A1(n13043), .A2(n11749), .ZN(n11710) );
  XNOR2_X1 U14142 ( .A(n11712), .B(n11710), .ZN(n12643) );
  INV_X1 U14143 ( .A(n11710), .ZN(n11711) );
  NAND2_X1 U14144 ( .A1(n11123), .A2(P2_REG0_REG_26__SCAN_IN), .ZN(n11719) );
  NAND2_X1 U14145 ( .A1(n11701), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n11718) );
  INV_X1 U14146 ( .A(n11714), .ZN(n11713) );
  NAND2_X1 U14147 ( .A1(n11713), .A2(P2_REG3_REG_26__SCAN_IN), .ZN(n11727) );
  INV_X1 U14148 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n12714) );
  NAND2_X1 U14149 ( .A1(n11714), .A2(n12714), .ZN(n11715) );
  AND2_X1 U14150 ( .A1(n11727), .A2(n11715), .ZN(n13204) );
  NAND2_X1 U14151 ( .A1(n9145), .A2(n13204), .ZN(n11717) );
  NAND2_X1 U14152 ( .A1(n11688), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n11716) );
  NAND4_X1 U14153 ( .A1(n11719), .A2(n11718), .A3(n11717), .A4(n11716), .ZN(
        n13042) );
  AND2_X1 U14154 ( .A1(n13042), .A2(n11749), .ZN(n11723) );
  NAND2_X1 U14155 ( .A1(n13434), .A2(n12943), .ZN(n11721) );
  NAND2_X1 U14156 ( .A1(n11862), .A2(P1_DATAO_REG_26__SCAN_IN), .ZN(n11720) );
  XNOR2_X1 U14157 ( .A(n12922), .B(n11750), .ZN(n11722) );
  NOR2_X1 U14158 ( .A1(n11722), .A2(n11723), .ZN(n11724) );
  AOI21_X1 U14159 ( .B1(n11723), .B2(n11722), .A(n11724), .ZN(n12708) );
  NAND2_X1 U14160 ( .A1(n11123), .A2(P2_REG0_REG_27__SCAN_IN), .ZN(n11732) );
  NAND2_X1 U14161 ( .A1(n9113), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n11731) );
  INV_X1 U14162 ( .A(n11727), .ZN(n11725) );
  NAND2_X1 U14163 ( .A1(n11725), .A2(P2_REG3_REG_27__SCAN_IN), .ZN(n11742) );
  INV_X1 U14164 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n11726) );
  NAND2_X1 U14165 ( .A1(n11727), .A2(n11726), .ZN(n11728) );
  NAND2_X1 U14166 ( .A1(n9145), .A2(n13191), .ZN(n11730) );
  NAND2_X1 U14167 ( .A1(n11688), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n11729) );
  NAND4_X1 U14168 ( .A1(n11732), .A2(n11731), .A3(n11730), .A4(n11729), .ZN(
        n13041) );
  NAND2_X1 U14169 ( .A1(n13041), .A2(n11749), .ZN(n11736) );
  NAND2_X1 U14170 ( .A1(n13431), .A2(n11860), .ZN(n11734) );
  NAND2_X1 U14171 ( .A1(n11862), .A2(P1_DATAO_REG_27__SCAN_IN), .ZN(n11733) );
  XNOR2_X1 U14172 ( .A(n13339), .B(n11750), .ZN(n11735) );
  XOR2_X1 U14173 ( .A(n11736), .B(n11735), .Z(n12609) );
  NAND2_X1 U14174 ( .A1(n11737), .A2(n12943), .ZN(n11739) );
  NAND2_X1 U14175 ( .A1(n9097), .A2(P1_DATAO_REG_28__SCAN_IN), .ZN(n11738) );
  NAND2_X1 U14176 ( .A1(n11123), .A2(P2_REG0_REG_28__SCAN_IN), .ZN(n11748) );
  NAND2_X1 U14177 ( .A1(n11701), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n11747) );
  INV_X1 U14178 ( .A(n11742), .ZN(n11740) );
  INV_X1 U14179 ( .A(n11887), .ZN(n11744) );
  INV_X1 U14180 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n11741) );
  NAND2_X1 U14181 ( .A1(n11742), .A2(n11741), .ZN(n11743) );
  NAND2_X1 U14182 ( .A1(n6485), .A2(n13181), .ZN(n11746) );
  NAND2_X1 U14183 ( .A1(n11688), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n11745) );
  NAND4_X1 U14184 ( .A1(n11748), .A2(n11747), .A3(n11746), .A4(n11745), .ZN(
        n13040) );
  NAND2_X1 U14185 ( .A1(n13040), .A2(n11749), .ZN(n11751) );
  XNOR2_X1 U14186 ( .A(n11751), .B(n11750), .ZN(n11752) );
  XNOR2_X1 U14187 ( .A(n13331), .B(n11752), .ZN(n11753) );
  XNOR2_X1 U14188 ( .A(n11754), .B(n11753), .ZN(n11765) );
  INV_X1 U14189 ( .A(n13181), .ZN(n11762) );
  NAND2_X1 U14190 ( .A1(n9113), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n11758) );
  NAND2_X1 U14191 ( .A1(n11688), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n11757) );
  NAND2_X1 U14192 ( .A1(n6485), .A2(n11887), .ZN(n11756) );
  NAND2_X1 U14193 ( .A1(n11123), .A2(P2_REG0_REG_29__SCAN_IN), .ZN(n11755) );
  NAND4_X1 U14194 ( .A1(n11758), .A2(n11757), .A3(n11756), .A4(n11755), .ZN(
        n13039) );
  NAND2_X1 U14195 ( .A1(n13039), .A2(n12711), .ZN(n11760) );
  NAND2_X1 U14196 ( .A1(n13041), .A2(n12710), .ZN(n11759) );
  NAND2_X1 U14197 ( .A1(n11760), .A2(n11759), .ZN(n13175) );
  AOI22_X1 U14198 ( .A1(n14330), .A2(n13175), .B1(P2_REG3_REG_28__SCAN_IN), 
        .B2(P2_U3088), .ZN(n11761) );
  OAI21_X1 U14199 ( .B1(n11762), .B2(n14334), .A(n11761), .ZN(n11763) );
  AOI21_X1 U14200 ( .B1(n13331), .B2(n12703), .A(n11763), .ZN(n11764) );
  OAI21_X1 U14201 ( .B1(n11765), .B2(n12705), .A(n11764), .ZN(P2_U3192) );
  INV_X1 U14202 ( .A(n11766), .ZN(n11769) );
  INV_X1 U14203 ( .A(n11767), .ZN(n11768) );
  AOI21_X2 U14204 ( .B1(n11772), .B2(n11771), .A(n11770), .ZN(n13500) );
  NAND2_X1 U14205 ( .A1(n14397), .A2(n13481), .ZN(n11774) );
  NAND2_X1 U14206 ( .A1(n13656), .A2(n13442), .ZN(n11773) );
  NAND2_X1 U14207 ( .A1(n11774), .A2(n11773), .ZN(n11775) );
  XNOR2_X1 U14208 ( .A(n11775), .B(n13536), .ZN(n11779) );
  NAND2_X1 U14209 ( .A1(n14397), .A2(n13442), .ZN(n11777) );
  NAND2_X1 U14210 ( .A1(n13485), .A2(n13656), .ZN(n11776) );
  NAND2_X1 U14211 ( .A1(n11777), .A2(n11776), .ZN(n11778) );
  NOR2_X1 U14212 ( .A1(n11779), .A2(n11778), .ZN(n11780) );
  AOI21_X1 U14213 ( .B1(n11779), .B2(n11778), .A(n11780), .ZN(n13501) );
  INV_X1 U14214 ( .A(n11780), .ZN(n11781) );
  NAND2_X1 U14215 ( .A1(n13648), .A2(n13481), .ZN(n11783) );
  OR2_X1 U14216 ( .A1(n13504), .A2(n13539), .ZN(n11782) );
  NAND2_X1 U14217 ( .A1(n11783), .A2(n11782), .ZN(n11784) );
  XNOR2_X1 U14218 ( .A(n11784), .B(n13471), .ZN(n11785) );
  AOI22_X1 U14219 ( .A1(n13648), .A2(n13442), .B1(n13485), .B2(n14385), .ZN(
        n13637) );
  NAND2_X1 U14220 ( .A1(n14409), .A2(n13481), .ZN(n11787) );
  NAND2_X1 U14221 ( .A1(n13655), .A2(n13442), .ZN(n11786) );
  NAND2_X1 U14222 ( .A1(n11787), .A2(n11786), .ZN(n11788) );
  XNOR2_X1 U14223 ( .A(n11788), .B(n13471), .ZN(n11791) );
  AND2_X1 U14224 ( .A1(n13485), .A2(n13655), .ZN(n11789) );
  AOI21_X1 U14225 ( .B1(n14409), .B2(n13442), .A(n11789), .ZN(n11790) );
  NAND2_X1 U14226 ( .A1(n11791), .A2(n11790), .ZN(n11792) );
  OAI21_X1 U14227 ( .B1(n11791), .B2(n11790), .A(n11792), .ZN(n13571) );
  INV_X1 U14228 ( .A(n11792), .ZN(n13582) );
  NAND2_X1 U14229 ( .A1(n14090), .A2(n13481), .ZN(n11794) );
  NAND2_X1 U14230 ( .A1(n13977), .A2(n13442), .ZN(n11793) );
  NAND2_X1 U14231 ( .A1(n11794), .A2(n11793), .ZN(n11795) );
  XNOR2_X1 U14232 ( .A(n11795), .B(n13471), .ZN(n11797) );
  AND2_X1 U14233 ( .A1(n13485), .A2(n13977), .ZN(n11796) );
  AOI21_X1 U14234 ( .B1(n14090), .B2(n13442), .A(n11796), .ZN(n11798) );
  NAND2_X1 U14235 ( .A1(n11797), .A2(n11798), .ZN(n11802) );
  INV_X1 U14236 ( .A(n11797), .ZN(n11800) );
  INV_X1 U14237 ( .A(n11798), .ZN(n11799) );
  NAND2_X1 U14238 ( .A1(n11800), .A2(n11799), .ZN(n11801) );
  AND2_X1 U14239 ( .A1(n11802), .A2(n11801), .ZN(n13581) );
  NAND2_X1 U14240 ( .A1(n13580), .A2(n11802), .ZN(n13612) );
  NAND2_X1 U14241 ( .A1(n13987), .A2(n13481), .ZN(n11804) );
  NAND2_X1 U14242 ( .A1(n13530), .A2(n13442), .ZN(n11803) );
  NAND2_X1 U14243 ( .A1(n11804), .A2(n11803), .ZN(n11805) );
  XNOR2_X1 U14244 ( .A(n11805), .B(n13536), .ZN(n11808) );
  AOI22_X1 U14245 ( .A1(n13987), .A2(n13442), .B1(n13485), .B2(n13530), .ZN(
        n11809) );
  XNOR2_X1 U14246 ( .A(n11808), .B(n11809), .ZN(n13613) );
  INV_X1 U14247 ( .A(n13978), .ZN(n13616) );
  OAI22_X1 U14248 ( .A1(n14083), .A2(n13535), .B1(n13616), .B2(n13539), .ZN(
        n11806) );
  XNOR2_X1 U14249 ( .A(n11806), .B(n13536), .ZN(n11812) );
  AND2_X1 U14250 ( .A1(n13978), .A2(n13485), .ZN(n11807) );
  AOI21_X1 U14251 ( .B1(n13969), .B2(n13442), .A(n11807), .ZN(n11813) );
  XNOR2_X1 U14252 ( .A(n11812), .B(n11813), .ZN(n13526) );
  INV_X1 U14253 ( .A(n11808), .ZN(n11810) );
  NAND2_X1 U14254 ( .A1(n11810), .A2(n11809), .ZN(n13524) );
  NAND2_X1 U14255 ( .A1(n13611), .A2(n11811), .ZN(n13525) );
  INV_X1 U14256 ( .A(n11813), .ZN(n11814) );
  NAND2_X1 U14257 ( .A1(n13525), .A2(n11815), .ZN(n13602) );
  OAI22_X1 U14258 ( .A1(n11816), .A2(n13539), .B1(n13964), .B2(n13538), .ZN(
        n11820) );
  NAND2_X1 U14259 ( .A1(n14078), .A2(n13481), .ZN(n11818) );
  NAND2_X1 U14260 ( .A1(n13935), .A2(n13442), .ZN(n11817) );
  NAND2_X1 U14261 ( .A1(n11818), .A2(n11817), .ZN(n11819) );
  XNOR2_X1 U14262 ( .A(n11819), .B(n13536), .ZN(n11821) );
  XOR2_X1 U14263 ( .A(n11820), .B(n11821), .Z(n13601) );
  NAND2_X1 U14264 ( .A1(n11821), .A2(n11820), .ZN(n11822) );
  NAND2_X1 U14265 ( .A1(n14072), .A2(n13481), .ZN(n11824) );
  NAND2_X1 U14266 ( .A1(n13945), .A2(n13442), .ZN(n11823) );
  NAND2_X1 U14267 ( .A1(n11824), .A2(n11823), .ZN(n11825) );
  XNOR2_X1 U14268 ( .A(n11825), .B(n13471), .ZN(n11828) );
  AND2_X1 U14269 ( .A1(n13945), .A2(n13485), .ZN(n11826) );
  AOI21_X1 U14270 ( .B1(n14072), .B2(n13442), .A(n11826), .ZN(n11827) );
  NAND2_X1 U14271 ( .A1(n11828), .A2(n11827), .ZN(n11838) );
  OAI21_X1 U14272 ( .B1(n11828), .B2(n11827), .A(n11838), .ZN(n13551) );
  INV_X1 U14273 ( .A(n11839), .ZN(n13550) );
  INV_X1 U14274 ( .A(n11838), .ZN(n11837) );
  OAI22_X1 U14275 ( .A1(n11572), .A2(n13535), .B1(n11917), .B2(n13539), .ZN(
        n11830) );
  XNOR2_X1 U14276 ( .A(n11830), .B(n13471), .ZN(n11832) );
  NOR2_X1 U14277 ( .A1(n11917), .A2(n13538), .ZN(n11831) );
  AOI21_X1 U14278 ( .B1(n6886), .B2(n13442), .A(n11831), .ZN(n11833) );
  NAND2_X1 U14279 ( .A1(n11832), .A2(n11833), .ZN(n13450) );
  INV_X1 U14280 ( .A(n11832), .ZN(n11835) );
  INV_X1 U14281 ( .A(n11833), .ZN(n11834) );
  NAND2_X1 U14282 ( .A1(n11835), .A2(n11834), .ZN(n11836) );
  AND2_X1 U14283 ( .A1(n13450), .A2(n11836), .ZN(n11840) );
  NOR3_X1 U14284 ( .A1(n13550), .A2(n11837), .A3(n11840), .ZN(n11843) );
  NAND2_X1 U14285 ( .A1(n11839), .A2(n11838), .ZN(n11841) );
  INV_X1 U14286 ( .A(n13451), .ZN(n11842) );
  OAI21_X1 U14287 ( .B1(n11843), .B2(n11842), .A(n13626), .ZN(n11847) );
  INV_X1 U14288 ( .A(n13644), .ZN(n13632) );
  INV_X1 U14289 ( .A(n13945), .ZN(n13917) );
  AOI22_X1 U14290 ( .A1(n13888), .A2(n13639), .B1(P1_REG3_REG_22__SCAN_IN), 
        .B2(P1_U3086), .ZN(n11844) );
  OAI21_X1 U14291 ( .B1(n13917), .B2(n13629), .A(n11844), .ZN(n11845) );
  AOI21_X1 U14292 ( .B1(n13923), .B2(n13632), .A(n11845), .ZN(n11846) );
  OAI211_X1 U14293 ( .C1(n13636), .C2(n11572), .A(n11847), .B(n11846), .ZN(
        P1_U3235) );
  XNOR2_X1 U14294 ( .A(n13368), .B(n13046), .ZN(n13260) );
  INV_X1 U14295 ( .A(n13260), .ZN(n13268) );
  INV_X1 U14296 ( .A(n13048), .ZN(n12879) );
  XNOR2_X1 U14297 ( .A(n13380), .B(n12879), .ZN(n13017) );
  NAND2_X1 U14298 ( .A1(n13380), .A2(n12879), .ZN(n11850) );
  INV_X1 U14299 ( .A(n13047), .ZN(n12692) );
  OR2_X1 U14300 ( .A1(n12885), .A2(n12692), .ZN(n11851) );
  NAND2_X1 U14301 ( .A1(n13275), .A2(n11851), .ZN(n11853) );
  NAND2_X1 U14302 ( .A1(n12885), .A2(n12692), .ZN(n11852) );
  NAND2_X1 U14303 ( .A1(n13363), .A2(n12691), .ZN(n11855) );
  INV_X1 U14304 ( .A(n13043), .ZN(n12674) );
  INV_X1 U14305 ( .A(n13042), .ZN(n11856) );
  INV_X1 U14306 ( .A(n13041), .ZN(n11857) );
  AOI22_X1 U14307 ( .A1(n13187), .A2(n13189), .B1(n11857), .B2(n13339), .ZN(
        n13172) );
  INV_X1 U14308 ( .A(n13040), .ZN(n11884) );
  NAND2_X1 U14309 ( .A1(n13331), .A2(n11884), .ZN(n11858) );
  NAND2_X1 U14310 ( .A1(n13172), .A2(n13173), .ZN(n13176) );
  NAND2_X1 U14311 ( .A1(n13176), .A2(n11859), .ZN(n11866) );
  NAND2_X1 U14312 ( .A1(n11861), .A2(n11860), .ZN(n11864) );
  NAND2_X1 U14313 ( .A1(n11862), .A2(P1_DATAO_REG_29__SCAN_IN), .ZN(n11863) );
  INV_X1 U14314 ( .A(n13039), .ZN(n11865) );
  XNOR2_X1 U14315 ( .A(n11866), .B(n13022), .ZN(n11875) );
  NAND2_X1 U14316 ( .A1(n11867), .A2(P2_B_REG_SCAN_IN), .ZN(n11868) );
  AND2_X1 U14317 ( .A1(n12711), .A2(n11868), .ZN(n13163) );
  INV_X1 U14318 ( .A(P2_REG1_REG_30__SCAN_IN), .ZN(n11871) );
  NAND2_X1 U14319 ( .A1(n11688), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n11870) );
  NAND2_X1 U14320 ( .A1(n9030), .A2(P2_REG0_REG_30__SCAN_IN), .ZN(n11869) );
  OAI211_X1 U14321 ( .C1(n11872), .C2(n11871), .A(n11870), .B(n11869), .ZN(
        n13038) );
  INV_X1 U14322 ( .A(n11873), .ZN(n11874) );
  AOI21_X2 U14323 ( .B1(n11875), .B2(n14740), .A(n11874), .ZN(n13328) );
  INV_X1 U14324 ( .A(n13380), .ZN(n12688) );
  OAI21_X1 U14325 ( .B1(n12688), .B2(n12879), .A(n13286), .ZN(n11877) );
  XNOR2_X1 U14326 ( .A(n12885), .B(n13047), .ZN(n13274) );
  INV_X1 U14327 ( .A(n13274), .ZN(n11878) );
  INV_X1 U14328 ( .A(n13247), .ZN(n13245) );
  OAI21_X1 U14329 ( .B1(n13236), .B2(n12623), .A(n13230), .ZN(n13214) );
  INV_X1 U14330 ( .A(n13214), .ZN(n11881) );
  NAND2_X1 U14331 ( .A1(n11881), .A2(n11880), .ZN(n13212) );
  NAND2_X1 U14332 ( .A1(n13212), .A2(n11882), .ZN(n13199) );
  NAND2_X1 U14333 ( .A1(n12922), .A2(n13042), .ZN(n11883) );
  INV_X1 U14334 ( .A(n13331), .ZN(n11886) );
  INV_X1 U14335 ( .A(n13022), .ZN(n11885) );
  INV_X1 U14336 ( .A(n13327), .ZN(n11890) );
  NOR2_X4 U14337 ( .A1(n13380), .A2(n13296), .ZN(n13299) );
  OR2_X1 U14338 ( .A1(n13238), .A2(n13352), .ZN(n13221) );
  INV_X1 U14339 ( .A(n13221), .ZN(n13203) );
  AOI211_X1 U14340 ( .C1(n13327), .C2(n13178), .A(n9329), .B(n13168), .ZN(
        n13326) );
  NAND2_X1 U14341 ( .A1(n13326), .A2(n14725), .ZN(n11889) );
  AOI22_X1 U14342 ( .A1(n14708), .A2(P2_REG2_REG_29__SCAN_IN), .B1(n11887), 
        .B2(n14719), .ZN(n11888) );
  OAI211_X1 U14343 ( .C1(n11890), .C2(n14721), .A(n11889), .B(n11888), .ZN(
        n11891) );
  AOI21_X1 U14344 ( .B1(n13325), .B2(n14727), .A(n11891), .ZN(n11892) );
  OAI21_X1 U14345 ( .B1(n13328), .B2(n14731), .A(n11892), .ZN(P2_U3236) );
  AND2_X1 U14346 ( .A1(n13969), .A2(n13616), .ZN(n13942) );
  NOR2_X1 U14347 ( .A1(n13949), .A2(n13942), .ZN(n11896) );
  NAND2_X1 U14348 ( .A1(n14409), .A2(n14007), .ZN(n14002) );
  AND2_X1 U14349 ( .A1(n14001), .A2(n14002), .ZN(n11893) );
  OR2_X1 U14350 ( .A1(n14090), .A2(n13573), .ZN(n11894) );
  OR2_X1 U14351 ( .A1(n13987), .A2(n14009), .ZN(n11895) );
  NOR2_X1 U14352 ( .A1(n11572), .A2(n13936), .ZN(n11898) );
  NAND2_X1 U14353 ( .A1(n14056), .A2(n13865), .ZN(n11899) );
  INV_X1 U14354 ( .A(n14049), .ZN(n13873) );
  INV_X1 U14355 ( .A(n13842), .ZN(n13846) );
  NAND2_X1 U14356 ( .A1(n11900), .A2(n11921), .ZN(n13828) );
  INV_X1 U14357 ( .A(n13847), .ZN(n11901) );
  NAND2_X1 U14358 ( .A1(n14038), .A2(n11901), .ZN(n11902) );
  INV_X1 U14359 ( .A(n14038), .ZN(n13835) );
  OR2_X1 U14360 ( .A1(n14410), .A2(n14090), .ZN(n13993) );
  NOR2_X2 U14361 ( .A1(n13987), .A2(n13993), .ZN(n13983) );
  NOR2_X2 U14362 ( .A1(n13833), .A2(n14032), .ZN(n12000) );
  AOI21_X1 U14363 ( .B1(n14032), .B2(n13833), .A(n12000), .ZN(n14033) );
  NOR2_X1 U14364 ( .A1(n14532), .A2(n13546), .ZN(n11903) );
  AOI21_X1 U14365 ( .B1(n14388), .B2(P1_REG2_REG_28__SCAN_IN), .A(n11903), 
        .ZN(n11904) );
  OAI21_X1 U14366 ( .B1(n13540), .B2(n14534), .A(n11904), .ZN(n11925) );
  INV_X1 U14367 ( .A(n13865), .ZN(n13462) );
  OR2_X1 U14368 ( .A1(n14409), .A2(n13655), .ZN(n11907) );
  AND2_X1 U14369 ( .A1(n13987), .A2(n13530), .ZN(n11912) );
  OR2_X1 U14370 ( .A1(n13987), .A2(n13530), .ZN(n11911) );
  NAND2_X1 U14371 ( .A1(n14078), .A2(n13935), .ZN(n11913) );
  OR2_X1 U14372 ( .A1(n14072), .A2(n13945), .ZN(n11914) );
  NAND2_X1 U14373 ( .A1(n11572), .A2(n11917), .ZN(n11918) );
  NAND2_X1 U14374 ( .A1(n14062), .A2(n13888), .ZN(n11919) );
  NAND2_X1 U14375 ( .A1(n13824), .A2(n13826), .ZN(n13823) );
  OAI21_X1 U14376 ( .B1(n14038), .B2(n13847), .A(n13823), .ZN(n11922) );
  NOR2_X1 U14377 ( .A1(n14031), .A2(n14015), .ZN(n11924) );
  OAI21_X1 U14378 ( .B1(n14035), .B2(n14388), .A(n11926), .ZN(P1_U3265) );
  XNOR2_X1 U14379 ( .A(n12562), .B(n11971), .ZN(n11951) );
  INV_X1 U14380 ( .A(n11951), .ZN(n11952) );
  XNOR2_X1 U14381 ( .A(n12575), .B(n11971), .ZN(n11938) );
  INV_X1 U14382 ( .A(n11938), .ZN(n11939) );
  INV_X1 U14383 ( .A(n11927), .ZN(n11929) );
  OAI21_X1 U14384 ( .B1(n11930), .B2(n11929), .A(n11928), .ZN(n14279) );
  XNOR2_X1 U14385 ( .A(n14275), .B(n11971), .ZN(n11931) );
  XNOR2_X1 U14386 ( .A(n11931), .B(n12129), .ZN(n14278) );
  NAND2_X1 U14387 ( .A1(n14279), .A2(n14278), .ZN(n14277) );
  INV_X1 U14388 ( .A(n11931), .ZN(n11933) );
  NAND2_X1 U14389 ( .A1(n11933), .A2(n12129), .ZN(n11934) );
  XNOR2_X1 U14390 ( .A(n12579), .B(n11971), .ZN(n11935) );
  XNOR2_X1 U14391 ( .A(n11935), .B(n12438), .ZN(n12054) );
  INV_X1 U14392 ( .A(n11935), .ZN(n11937) );
  XNOR2_X1 U14393 ( .A(n11938), .B(n11940), .ZN(n12061) );
  OAI21_X1 U14394 ( .B1(n11940), .B2(n11939), .A(n12060), .ZN(n12091) );
  XNOR2_X1 U14395 ( .A(n12088), .B(n11971), .ZN(n11942) );
  XNOR2_X1 U14396 ( .A(n11942), .B(n12127), .ZN(n12090) );
  NAND2_X1 U14397 ( .A1(n12091), .A2(n12090), .ZN(n12089) );
  NAND2_X1 U14398 ( .A1(n12089), .A2(n11943), .ZN(n12036) );
  XNOR2_X1 U14399 ( .A(n12518), .B(n11971), .ZN(n11945) );
  XNOR2_X1 U14400 ( .A(n11945), .B(n12126), .ZN(n12035) );
  NAND2_X1 U14401 ( .A1(n12036), .A2(n12035), .ZN(n12034) );
  NAND2_X1 U14402 ( .A1(n12034), .A2(n11946), .ZN(n12078) );
  XNOR2_X1 U14403 ( .A(n11947), .B(n11971), .ZN(n11949) );
  XNOR2_X1 U14404 ( .A(n11949), .B(n12125), .ZN(n12077) );
  XNOR2_X1 U14405 ( .A(n11951), .B(n12124), .ZN(n12041) );
  XNOR2_X1 U14406 ( .A(n12355), .B(n11971), .ZN(n11955) );
  XNOR2_X1 U14407 ( .A(n11954), .B(n11955), .ZN(n12083) );
  XNOR2_X1 U14408 ( .A(n12031), .B(n11971), .ZN(n11957) );
  XNOR2_X1 U14409 ( .A(n11956), .B(n11957), .ZN(n12025) );
  NAND2_X1 U14410 ( .A1(n12025), .A2(n12070), .ZN(n11960) );
  INV_X1 U14411 ( .A(n11956), .ZN(n11958) );
  NAND2_X1 U14412 ( .A1(n11960), .A2(n11959), .ZN(n12067) );
  XNOR2_X1 U14413 ( .A(n12499), .B(n11971), .ZN(n11961) );
  XNOR2_X1 U14414 ( .A(n11961), .B(n12027), .ZN(n12068) );
  NAND2_X1 U14415 ( .A1(n12067), .A2(n12068), .ZN(n11964) );
  INV_X1 U14416 ( .A(n11961), .ZN(n11962) );
  XNOR2_X1 U14417 ( .A(n12317), .B(n11971), .ZN(n11965) );
  XNOR2_X1 U14418 ( .A(n11965), .B(n12120), .ZN(n12047) );
  XNOR2_X1 U14419 ( .A(n12304), .B(n11971), .ZN(n11969) );
  XNOR2_X1 U14420 ( .A(n11969), .B(n12119), .ZN(n12110) );
  NAND2_X1 U14421 ( .A1(n11969), .A2(n11968), .ZN(n11970) );
  XNOR2_X1 U14422 ( .A(n12022), .B(n11971), .ZN(n11972) );
  XNOR2_X1 U14423 ( .A(n11972), .B(n7281), .ZN(n12018) );
  XNOR2_X1 U14424 ( .A(n11974), .B(n11971), .ZN(n11975) );
  INV_X1 U14425 ( .A(n11976), .ZN(n12280) );
  NOR2_X1 U14426 ( .A1(n12280), .A2(n14286), .ZN(n11979) );
  OAI22_X1 U14427 ( .A1(n11977), .A2(n14281), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15066), .ZN(n11978) );
  AOI211_X1 U14428 ( .C1(n12282), .C2(n14274), .A(n11979), .B(n11978), .ZN(
        n11980) );
  OAI21_X1 U14429 ( .B1(n11981), .B2(n12115), .A(n11980), .ZN(P3_U3160) );
  AOI22_X1 U14430 ( .A1(n14330), .A2(n11983), .B1(n11982), .B2(
        P2_REG3_REG_1__SCAN_IN), .ZN(n11989) );
  OAI21_X1 U14431 ( .B1(n11986), .B2(n11985), .A(n11984), .ZN(n11987) );
  NAND2_X1 U14432 ( .A1(n14328), .A2(n11987), .ZN(n11988) );
  OAI211_X1 U14433 ( .C1(n12719), .C2(n9021), .A(n11989), .B(n11988), .ZN(
        P2_U3194) );
  OAI222_X1 U14434 ( .A1(P2_U3088), .A2(n11991), .B1(n13438), .B2(n14118), 
        .C1(n11990), .C2(n13440), .ZN(P2_U3297) );
  OR2_X1 U14435 ( .A1(n12275), .A2(n12537), .ZN(n11994) );
  OR2_X1 U14436 ( .A1(n14032), .A2(n13829), .ZN(n11996) );
  AND2_X1 U14437 ( .A1(n14032), .A2(n13829), .ZN(n11995) );
  AOI21_X1 U14438 ( .B1(n11997), .B2(n11996), .A(n11995), .ZN(n11999) );
  XNOR2_X1 U14439 ( .A(n11999), .B(n11998), .ZN(n14029) );
  NAND2_X1 U14440 ( .A1(n14027), .A2(n12000), .ZN(n13819) );
  OR2_X1 U14441 ( .A1(n14027), .A2(n12000), .ZN(n12001) );
  NOR2_X1 U14442 ( .A1(n14024), .A2(n13989), .ZN(n12009) );
  AOI21_X1 U14443 ( .B1(n12002), .B2(P1_B_REG_SCAN_IN), .A(n14008), .ZN(n13813) );
  NAND2_X1 U14444 ( .A1(n13652), .A2(n13813), .ZN(n14025) );
  OAI22_X1 U14445 ( .A1(n12004), .A2(n14025), .B1(n12003), .B2(n14532), .ZN(
        n12006) );
  NAND2_X1 U14446 ( .A1(n13654), .A2(n14527), .ZN(n14026) );
  NOR2_X1 U14447 ( .A1(n14531), .A2(n14026), .ZN(n12005) );
  AOI211_X1 U14448 ( .C1(n14388), .C2(P1_REG2_REG_29__SCAN_IN), .A(n12006), 
        .B(n12005), .ZN(n12007) );
  OAI21_X1 U14449 ( .B1(n14027), .B2(n14534), .A(n12007), .ZN(n12008) );
  AOI211_X1 U14450 ( .C1(n14029), .C2(n12010), .A(n12009), .B(n12008), .ZN(
        n12011) );
  OAI21_X1 U14451 ( .B1(n14030), .B2(n14015), .A(n12011), .ZN(P1_U3356) );
  OAI222_X1 U14452 ( .A1(n13440), .A2(n12013), .B1(n13438), .B2(n12012), .C1(
        n13253), .C2(P2_U3088), .ZN(P2_U3308) );
  INV_X1 U14453 ( .A(n12014), .ZN(n12016) );
  INV_X1 U14454 ( .A(SI_30_), .ZN(n15056) );
  OAI222_X1 U14455 ( .A1(n12607), .A2(n12016), .B1(n12015), .B2(P3_U3151), 
        .C1(n15056), .C2(n12608), .ZN(P3_U3265) );
  XOR2_X1 U14456 ( .A(n12018), .B(n12017), .Z(n12024) );
  AOI22_X1 U14457 ( .A1(n12112), .A2(n12288), .B1(P3_REG3_REG_27__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12019) );
  OAI21_X1 U14458 ( .B1(n12020), .B2(n14281), .A(n12019), .ZN(n12021) );
  AOI21_X1 U14459 ( .B1(n12022), .B2(n14274), .A(n12021), .ZN(n12023) );
  OAI21_X1 U14460 ( .B1(n12024), .B2(n12115), .A(n12023), .ZN(P3_U3154) );
  XNOR2_X1 U14461 ( .A(n12025), .B(n12122), .ZN(n12033) );
  INV_X1 U14462 ( .A(n12342), .ZN(n12029) );
  OAI22_X1 U14463 ( .A1(n12027), .A2(n12100), .B1(n12026), .B2(n12103), .ZN(
        n12337) );
  AOI22_X1 U14464 ( .A1(n12337), .A2(n12104), .B1(P3_REG3_REG_23__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12028) );
  OAI21_X1 U14465 ( .B1(n12029), .B2(n14286), .A(n12028), .ZN(n12030) );
  AOI21_X1 U14466 ( .B1(n12031), .B2(n14274), .A(n12030), .ZN(n12032) );
  OAI21_X1 U14467 ( .B1(n12033), .B2(n12115), .A(n12032), .ZN(P3_U3156) );
  OAI211_X1 U14468 ( .C1(n12036), .C2(n12035), .A(n12034), .B(n14276), .ZN(
        n12039) );
  AOI22_X1 U14469 ( .A1(n12440), .A2(n12127), .B1(n12125), .B2(n12437), .ZN(
        n12388) );
  INV_X1 U14470 ( .A(P3_REG3_REG_19__SCAN_IN), .ZN(n15204) );
  OAI22_X1 U14471 ( .A1(n12388), .A2(n14281), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15204), .ZN(n12037) );
  AOI21_X1 U14472 ( .B1(n12390), .B2(n12112), .A(n12037), .ZN(n12038) );
  OAI211_X1 U14473 ( .C1(n12392), .C2(n12095), .A(n12039), .B(n12038), .ZN(
        P3_U3159) );
  AOI21_X1 U14474 ( .B1(n12041), .B2(n12040), .A(n6598), .ZN(n12045) );
  AOI22_X1 U14475 ( .A1(n12440), .A2(n12125), .B1(n12123), .B2(n12437), .ZN(
        n12364) );
  OAI22_X1 U14476 ( .A1(n12364), .A2(n14281), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15192), .ZN(n12043) );
  NOR2_X1 U14477 ( .A1(n12562), .A2(n12095), .ZN(n12042) );
  AOI211_X1 U14478 ( .C1(n12366), .C2(n12112), .A(n12043), .B(n12042), .ZN(
        n12044) );
  OAI21_X1 U14479 ( .B1(n12045), .B2(n12115), .A(n12044), .ZN(P3_U3163) );
  XOR2_X1 U14480 ( .A(n12047), .B(n12046), .Z(n12051) );
  AOI22_X1 U14481 ( .A1(n12119), .A2(n12437), .B1(n12440), .B2(n12121), .ZN(
        n12315) );
  AOI22_X1 U14482 ( .A1(n12112), .A2(n12318), .B1(P3_REG3_REG_25__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12048) );
  OAI21_X1 U14483 ( .B1(n12315), .B2(n14281), .A(n12048), .ZN(n12049) );
  AOI21_X1 U14484 ( .B1(n12317), .B2(n14274), .A(n12049), .ZN(n12050) );
  OAI21_X1 U14485 ( .B1(n12051), .B2(n12115), .A(n12050), .ZN(P3_U3165) );
  AOI21_X1 U14486 ( .B1(n12054), .B2(n12053), .A(n12052), .ZN(n12059) );
  AOI22_X1 U14487 ( .A1(n12440), .A2(n12129), .B1(n12128), .B2(n12437), .ZN(
        n12426) );
  NAND2_X1 U14488 ( .A1(n12112), .A2(n12431), .ZN(n12055) );
  NAND2_X1 U14489 ( .A1(P3_U3151), .A2(P3_REG3_REG_16__SCAN_IN), .ZN(n12221)
         );
  OAI211_X1 U14490 ( .C1(n12426), .C2(n14281), .A(n12055), .B(n12221), .ZN(
        n12056) );
  AOI21_X1 U14491 ( .B1(n12057), .B2(n14274), .A(n12056), .ZN(n12058) );
  OAI21_X1 U14492 ( .B1(n12059), .B2(n12115), .A(n12058), .ZN(P3_U3166) );
  OAI211_X1 U14493 ( .C1(n12062), .C2(n12061), .A(n12060), .B(n14276), .ZN(
        n12066) );
  AOI22_X1 U14494 ( .A1(n12127), .A2(n12437), .B1(n12440), .B2(n12438), .ZN(
        n12418) );
  OAI22_X1 U14495 ( .A1(n12418), .A2(n14281), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12063), .ZN(n12064) );
  AOI21_X1 U14496 ( .B1(n12420), .B2(n12112), .A(n12064), .ZN(n12065) );
  OAI211_X1 U14497 ( .C1(n12575), .C2(n12095), .A(n12066), .B(n12065), .ZN(
        P3_U3168) );
  XOR2_X1 U14498 ( .A(n12068), .B(n12067), .Z(n12075) );
  INV_X1 U14499 ( .A(n12069), .ZN(n12327) );
  OAI22_X1 U14500 ( .A1(n12071), .A2(n12100), .B1(n12070), .B2(n12103), .ZN(
        n12324) );
  AOI22_X1 U14501 ( .A1(n12324), .A2(n12104), .B1(P3_REG3_REG_24__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12072) );
  OAI21_X1 U14502 ( .B1(n12327), .B2(n14286), .A(n12072), .ZN(n12073) );
  AOI21_X1 U14503 ( .B1(n12330), .B2(n14274), .A(n12073), .ZN(n12074) );
  OAI21_X1 U14504 ( .B1(n12075), .B2(n12115), .A(n12074), .ZN(P3_U3169) );
  OAI211_X1 U14505 ( .C1(n12078), .C2(n12077), .A(n12076), .B(n14276), .ZN(
        n12082) );
  AOI22_X1 U14506 ( .A1(n12440), .A2(n12126), .B1(n12124), .B2(n12437), .ZN(
        n12372) );
  OAI22_X1 U14507 ( .A1(n12372), .A2(n14281), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12079), .ZN(n12080) );
  AOI21_X1 U14508 ( .B1(n12374), .B2(n12112), .A(n12080), .ZN(n12081) );
  OAI211_X1 U14509 ( .C1(n12566), .C2(n12095), .A(n12082), .B(n12081), .ZN(
        P3_U3173) );
  XNOR2_X1 U14510 ( .A(n12083), .B(n12123), .ZN(n12087) );
  AOI22_X1 U14511 ( .A1(n12437), .A2(n12122), .B1(n12124), .B2(n12440), .ZN(
        n12353) );
  INV_X1 U14512 ( .A(P3_REG3_REG_22__SCAN_IN), .ZN(n15082) );
  OAI22_X1 U14513 ( .A1(n12353), .A2(n14281), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15082), .ZN(n12084) );
  AOI21_X1 U14514 ( .B1(n12356), .B2(n12112), .A(n12084), .ZN(n12086) );
  NAND2_X1 U14515 ( .A1(n12355), .A2(n14274), .ZN(n12085) );
  OAI211_X1 U14516 ( .C1(n12087), .C2(n12115), .A(n12086), .B(n12085), .ZN(
        P3_U3175) );
  INV_X1 U14517 ( .A(n12088), .ZN(n12571) );
  OAI211_X1 U14518 ( .C1(n12091), .C2(n12090), .A(n12089), .B(n14276), .ZN(
        n12094) );
  AOI22_X1 U14519 ( .A1(n12126), .A2(n12437), .B1(n12440), .B2(n12128), .ZN(
        n12403) );
  NAND2_X1 U14520 ( .A1(P3_U3151), .A2(P3_REG3_REG_18__SCAN_IN), .ZN(n12258)
         );
  OAI21_X1 U14521 ( .B1(n12403), .B2(n14281), .A(n12258), .ZN(n12092) );
  AOI21_X1 U14522 ( .B1(n12405), .B2(n12112), .A(n12092), .ZN(n12093) );
  OAI211_X1 U14523 ( .C1(n12571), .C2(n12095), .A(n12094), .B(n12093), .ZN(
        P3_U3178) );
  OAI211_X1 U14524 ( .C1(n12098), .C2(n12097), .A(n12096), .B(n14276), .ZN(
        n12108) );
  AOI22_X1 U14525 ( .A1(n14274), .A2(n14996), .B1(P3_REG3_REG_6__SCAN_IN), 
        .B2(P3_U3151), .ZN(n12107) );
  NAND2_X1 U14526 ( .A1(n12112), .A2(n12099), .ZN(n12106) );
  OR2_X1 U14527 ( .A1(n12101), .A2(n12100), .ZN(n12102) );
  OAI21_X1 U14528 ( .B1(n7638), .B2(n12103), .A(n12102), .ZN(n14933) );
  NAND2_X1 U14529 ( .A1(n14933), .A2(n12104), .ZN(n12105) );
  NAND4_X1 U14530 ( .A1(n12108), .A2(n12107), .A3(n12106), .A4(n12105), .ZN(
        P3_U3179) );
  XOR2_X1 U14531 ( .A(n12110), .B(n12109), .Z(n12116) );
  AOI22_X1 U14532 ( .A1(n7281), .A2(n12437), .B1(n12440), .B2(n12120), .ZN(
        n12302) );
  OAI22_X1 U14533 ( .A1(n12302), .A2(n14281), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n15206), .ZN(n12111) );
  AOI21_X1 U14534 ( .B1(n12305), .B2(n12112), .A(n12111), .ZN(n12114) );
  NAND2_X1 U14535 ( .A1(n12304), .A2(n14274), .ZN(n12113) );
  OAI211_X1 U14536 ( .C1(n12116), .C2(n12115), .A(n12114), .B(n12113), .ZN(
        P3_U3180) );
  MUX2_X1 U14537 ( .A(n12267), .B(P3_DATAO_REG_31__SCAN_IN), .S(n12143), .Z(
        P3_U3522) );
  MUX2_X1 U14538 ( .A(n12117), .B(P3_DATAO_REG_30__SCAN_IN), .S(n12143), .Z(
        P3_U3521) );
  MUX2_X1 U14539 ( .A(P3_DATAO_REG_28__SCAN_IN), .B(n12118), .S(P3_U3897), .Z(
        P3_U3519) );
  MUX2_X1 U14540 ( .A(n7281), .B(P3_DATAO_REG_27__SCAN_IN), .S(n12143), .Z(
        P3_U3518) );
  MUX2_X1 U14541 ( .A(P3_DATAO_REG_26__SCAN_IN), .B(n12119), .S(P3_U3897), .Z(
        P3_U3517) );
  MUX2_X1 U14542 ( .A(n12120), .B(P3_DATAO_REG_25__SCAN_IN), .S(n12143), .Z(
        P3_U3516) );
  MUX2_X1 U14543 ( .A(n12121), .B(P3_DATAO_REG_24__SCAN_IN), .S(n12143), .Z(
        P3_U3515) );
  MUX2_X1 U14544 ( .A(P3_DATAO_REG_23__SCAN_IN), .B(n12122), .S(P3_U3897), .Z(
        P3_U3514) );
  MUX2_X1 U14545 ( .A(P3_DATAO_REG_22__SCAN_IN), .B(n12123), .S(P3_U3897), .Z(
        P3_U3513) );
  MUX2_X1 U14546 ( .A(P3_DATAO_REG_21__SCAN_IN), .B(n12124), .S(P3_U3897), .Z(
        P3_U3512) );
  MUX2_X1 U14547 ( .A(P3_DATAO_REG_20__SCAN_IN), .B(n12125), .S(P3_U3897), .Z(
        P3_U3511) );
  MUX2_X1 U14548 ( .A(P3_DATAO_REG_19__SCAN_IN), .B(n12126), .S(P3_U3897), .Z(
        P3_U3510) );
  MUX2_X1 U14549 ( .A(P3_DATAO_REG_18__SCAN_IN), .B(n12127), .S(P3_U3897), .Z(
        P3_U3509) );
  MUX2_X1 U14550 ( .A(n12128), .B(P3_DATAO_REG_17__SCAN_IN), .S(n12143), .Z(
        P3_U3508) );
  MUX2_X1 U14551 ( .A(n12438), .B(P3_DATAO_REG_16__SCAN_IN), .S(n12143), .Z(
        P3_U3507) );
  MUX2_X1 U14552 ( .A(n12129), .B(P3_DATAO_REG_15__SCAN_IN), .S(n12143), .Z(
        P3_U3506) );
  MUX2_X1 U14553 ( .A(n12439), .B(P3_DATAO_REG_14__SCAN_IN), .S(n12143), .Z(
        P3_U3505) );
  MUX2_X1 U14554 ( .A(n12130), .B(P3_DATAO_REG_13__SCAN_IN), .S(n12143), .Z(
        P3_U3504) );
  MUX2_X1 U14555 ( .A(n12131), .B(P3_DATAO_REG_12__SCAN_IN), .S(n12143), .Z(
        P3_U3503) );
  MUX2_X1 U14556 ( .A(P3_DATAO_REG_11__SCAN_IN), .B(n12132), .S(P3_U3897), .Z(
        P3_U3502) );
  MUX2_X1 U14557 ( .A(P3_DATAO_REG_10__SCAN_IN), .B(n12133), .S(P3_U3897), .Z(
        P3_U3501) );
  MUX2_X1 U14558 ( .A(n12134), .B(P3_DATAO_REG_9__SCAN_IN), .S(n12143), .Z(
        P3_U3500) );
  MUX2_X1 U14559 ( .A(P3_DATAO_REG_8__SCAN_IN), .B(n12135), .S(P3_U3897), .Z(
        P3_U3499) );
  MUX2_X1 U14560 ( .A(P3_DATAO_REG_7__SCAN_IN), .B(n12136), .S(P3_U3897), .Z(
        P3_U3498) );
  MUX2_X1 U14561 ( .A(n12137), .B(P3_DATAO_REG_6__SCAN_IN), .S(n12143), .Z(
        P3_U3497) );
  MUX2_X1 U14562 ( .A(P3_DATAO_REG_5__SCAN_IN), .B(n12138), .S(P3_U3897), .Z(
        P3_U3496) );
  MUX2_X1 U14563 ( .A(P3_DATAO_REG_4__SCAN_IN), .B(n12139), .S(P3_U3897), .Z(
        P3_U3495) );
  MUX2_X1 U14564 ( .A(n12140), .B(P3_DATAO_REG_3__SCAN_IN), .S(n12143), .Z(
        P3_U3494) );
  MUX2_X1 U14565 ( .A(P3_DATAO_REG_2__SCAN_IN), .B(n12141), .S(P3_U3897), .Z(
        P3_U3493) );
  MUX2_X1 U14566 ( .A(n12142), .B(P3_DATAO_REG_1__SCAN_IN), .S(n12143), .Z(
        P3_U3492) );
  MUX2_X1 U14567 ( .A(n12144), .B(P3_DATAO_REG_0__SCAN_IN), .S(n12143), .Z(
        P3_U3491) );
  AOI21_X1 U14568 ( .B1(n12147), .B2(n12146), .A(n12145), .ZN(n12148) );
  NOR2_X1 U14569 ( .A1(n12148), .A2(n14893), .ZN(n12161) );
  AOI21_X1 U14570 ( .B1(n6595), .B2(n12150), .A(n12149), .ZN(n12151) );
  NOR2_X1 U14571 ( .A1(n12151), .A2(n14887), .ZN(n12160) );
  AOI21_X1 U14572 ( .B1(n14869), .B2(P3_ADDR_REG_12__SCAN_IN), .A(n12152), 
        .ZN(n12157) );
  XNOR2_X1 U14573 ( .A(n12153), .B(n12154), .ZN(n12155) );
  NAND2_X1 U14574 ( .A1(n12155), .A2(n14843), .ZN(n12156) );
  OAI211_X1 U14575 ( .C1(n14878), .C2(n12158), .A(n12157), .B(n12156), .ZN(
        n12159) );
  OR3_X1 U14576 ( .A1(n12161), .A2(n12160), .A3(n12159), .ZN(P3_U3194) );
  AOI21_X1 U14577 ( .B1(n14303), .B2(n12163), .A(n12162), .ZN(n12177) );
  AOI21_X1 U14578 ( .B1(n12166), .B2(n12165), .A(n12164), .ZN(n12167) );
  OR2_X1 U14579 ( .A1(n12167), .A2(n14893), .ZN(n12176) );
  AOI21_X1 U14580 ( .B1(n12169), .B2(n12168), .A(n12185), .ZN(n12170) );
  INV_X1 U14581 ( .A(n14843), .ZN(n14885) );
  NOR2_X1 U14582 ( .A1(n12170), .A2(n14885), .ZN(n12174) );
  INV_X1 U14583 ( .A(P3_ADDR_REG_13__SCAN_IN), .ZN(n12172) );
  OAI21_X1 U14584 ( .B1(n14875), .B2(n12172), .A(n12171), .ZN(n12173) );
  AOI211_X1 U14585 ( .C1(n14846), .C2(n8266), .A(n12174), .B(n12173), .ZN(
        n12175) );
  OAI211_X1 U14586 ( .C1(n12177), .C2(n14887), .A(n12176), .B(n12175), .ZN(
        P3_U3195) );
  AOI21_X1 U14587 ( .B1(n6596), .B2(n12179), .A(n12178), .ZN(n12196) );
  AOI21_X1 U14588 ( .B1(n12182), .B2(n12181), .A(n12180), .ZN(n12183) );
  OR2_X1 U14589 ( .A1(n12183), .A2(n14893), .ZN(n12195) );
  INV_X1 U14590 ( .A(P3_ADDR_REG_14__SCAN_IN), .ZN(n12191) );
  OAI21_X1 U14591 ( .B1(n12186), .B2(n12185), .A(n12184), .ZN(n12188) );
  NAND3_X1 U14592 ( .A1(n12188), .A2(n14843), .A3(n12187), .ZN(n12189) );
  OAI211_X1 U14593 ( .C1(n14875), .C2(n12191), .A(n12190), .B(n12189), .ZN(
        n12192) );
  AOI21_X1 U14594 ( .B1(n12193), .B2(n14846), .A(n12192), .ZN(n12194) );
  OAI211_X1 U14595 ( .C1(n12196), .C2(n14887), .A(n12195), .B(n12194), .ZN(
        P3_U3196) );
  AOI21_X1 U14596 ( .B1(n12199), .B2(n12198), .A(n12197), .ZN(n12213) );
  AOI21_X1 U14597 ( .B1(n12202), .B2(n12201), .A(n12200), .ZN(n12203) );
  INV_X1 U14598 ( .A(n12203), .ZN(n12211) );
  NAND2_X1 U14599 ( .A1(P3_U3151), .A2(P3_REG3_REG_15__SCAN_IN), .ZN(n14272)
         );
  NAND2_X1 U14600 ( .A1(n14869), .A2(P3_ADDR_REG_15__SCAN_IN), .ZN(n12204) );
  OAI211_X1 U14601 ( .C1(n14878), .C2(n12205), .A(n14272), .B(n12204), .ZN(
        n12210) );
  AOI21_X1 U14602 ( .B1(n12535), .B2(n12207), .A(n12206), .ZN(n12208) );
  NOR2_X1 U14603 ( .A1(n12208), .A2(n14887), .ZN(n12209) );
  AOI211_X1 U14604 ( .C1(n14843), .C2(n12211), .A(n12210), .B(n12209), .ZN(
        n12212) );
  OAI21_X1 U14605 ( .B1(n12213), .B2(n14893), .A(n12212), .ZN(P3_U3197) );
  AOI21_X1 U14606 ( .B1(n6535), .B2(n12215), .A(n12214), .ZN(n12231) );
  NOR2_X1 U14607 ( .A1(n12217), .A2(n12216), .ZN(n12219) );
  XOR2_X1 U14608 ( .A(n12219), .B(n12218), .Z(n12229) );
  NAND2_X1 U14609 ( .A1(n14869), .A2(P3_ADDR_REG_16__SCAN_IN), .ZN(n12220) );
  OAI211_X1 U14610 ( .C1(n14878), .C2(n12222), .A(n12221), .B(n12220), .ZN(
        n12228) );
  AOI21_X1 U14611 ( .B1(n12225), .B2(n12224), .A(n12223), .ZN(n12226) );
  NOR2_X1 U14612 ( .A1(n12226), .A2(n14887), .ZN(n12227) );
  AOI211_X1 U14613 ( .C1(n14843), .C2(n12229), .A(n12228), .B(n12227), .ZN(
        n12230) );
  OAI21_X1 U14614 ( .B1(n12231), .B2(n14893), .A(n12230), .ZN(P3_U3198) );
  AOI21_X1 U14615 ( .B1(n12234), .B2(n12233), .A(n12232), .ZN(n12249) );
  NAND2_X1 U14616 ( .A1(n12236), .A2(n12235), .ZN(n12237) );
  NAND2_X1 U14617 ( .A1(n12237), .A2(n14843), .ZN(n12240) );
  NOR2_X1 U14618 ( .A1(P3_STATE_REG_SCAN_IN), .A2(n12063), .ZN(n12238) );
  AOI21_X1 U14619 ( .B1(n14869), .B2(P3_ADDR_REG_17__SCAN_IN), .A(n12238), 
        .ZN(n12239) );
  OAI21_X1 U14620 ( .B1(n12241), .B2(n12240), .A(n12239), .ZN(n12246) );
  AOI21_X1 U14621 ( .B1(n12527), .B2(n12243), .A(n12242), .ZN(n12244) );
  NOR2_X1 U14622 ( .A1(n12244), .A2(n14887), .ZN(n12245) );
  AOI211_X1 U14623 ( .C1(n14846), .C2(n12247), .A(n12246), .B(n12245), .ZN(
        n12248) );
  OAI21_X1 U14624 ( .B1(n12249), .B2(n14893), .A(n12248), .ZN(P3_U3199) );
  AOI21_X1 U14625 ( .B1(n12252), .B2(n12251), .A(n12250), .ZN(n12264) );
  INV_X1 U14626 ( .A(P3_ADDR_REG_18__SCAN_IN), .ZN(n12259) );
  OAI21_X1 U14627 ( .B1(n12255), .B2(n12254), .A(n12253), .ZN(n12256) );
  NAND2_X1 U14628 ( .A1(n14843), .A2(n12256), .ZN(n12257) );
  NAND2_X1 U14629 ( .A1(n12273), .A2(n14973), .ZN(n12268) );
  INV_X1 U14630 ( .A(n12265), .ZN(n12266) );
  NAND2_X1 U14631 ( .A1(n12267), .A2(n12266), .ZN(n14291) );
  AOI21_X1 U14632 ( .B1(n12268), .B2(n14291), .A(n14979), .ZN(n12270) );
  AOI21_X1 U14633 ( .B1(n14979), .B2(P3_REG2_REG_31__SCAN_IN), .A(n12270), 
        .ZN(n12269) );
  OAI21_X1 U14634 ( .B1(n14288), .B2(n14906), .A(n12269), .ZN(P3_U3202) );
  AOI21_X1 U14635 ( .B1(n14979), .B2(P3_REG2_REG_30__SCAN_IN), .A(n12270), 
        .ZN(n12271) );
  OAI21_X1 U14636 ( .B1(n14292), .B2(n14906), .A(n12271), .ZN(P3_U3203) );
  AOI22_X1 U14637 ( .A1(n12273), .A2(n14973), .B1(P3_REG2_REG_29__SCAN_IN), 
        .B2(n14979), .ZN(n12274) );
  OAI21_X1 U14638 ( .B1(n12275), .B2(n14906), .A(n12274), .ZN(n12276) );
  AOI21_X1 U14639 ( .B1(n12277), .B2(n14941), .A(n12276), .ZN(n12278) );
  OAI21_X1 U14640 ( .B1(n7173), .B2(n14979), .A(n12278), .ZN(P3_U3204) );
  INV_X1 U14641 ( .A(P3_REG2_REG_28__SCAN_IN), .ZN(n12279) );
  OAI22_X1 U14642 ( .A1(n12280), .A2(n14959), .B1(n14977), .B2(n12279), .ZN(
        n12281) );
  AOI21_X1 U14643 ( .B1(n12282), .B2(n14957), .A(n12281), .ZN(n12285) );
  NAND2_X1 U14644 ( .A1(n12283), .A2(n14941), .ZN(n12284) );
  OAI211_X1 U14645 ( .C1(n12286), .C2(n14979), .A(n12285), .B(n12284), .ZN(
        P3_U3205) );
  INV_X1 U14646 ( .A(n12287), .ZN(n12293) );
  AOI22_X1 U14647 ( .A1(n12288), .A2(n14973), .B1(n14979), .B2(
        P3_REG2_REG_27__SCAN_IN), .ZN(n12289) );
  OAI21_X1 U14648 ( .B1(n12541), .B2(n14906), .A(n12289), .ZN(n12290) );
  AOI21_X1 U14649 ( .B1(n12291), .B2(n14977), .A(n12290), .ZN(n12292) );
  OAI21_X1 U14650 ( .B1(n12486), .B2(n12293), .A(n12292), .ZN(P3_U3206) );
  NAND2_X1 U14651 ( .A1(n12294), .A2(n12295), .ZN(n12310) );
  NAND2_X1 U14652 ( .A1(n12310), .A2(n12312), .ZN(n12297) );
  NAND2_X1 U14653 ( .A1(n12297), .A2(n12296), .ZN(n12298) );
  XOR2_X1 U14654 ( .A(n12300), .B(n12298), .Z(n12489) );
  INV_X1 U14655 ( .A(n12489), .ZN(n12309) );
  NAND2_X1 U14656 ( .A1(n12313), .A2(n12299), .ZN(n12301) );
  XNOR2_X1 U14657 ( .A(n12301), .B(n12300), .ZN(n12303) );
  OAI21_X1 U14658 ( .B1(n12303), .B2(n14949), .A(n12302), .ZN(n12488) );
  INV_X1 U14659 ( .A(n12304), .ZN(n12545) );
  AOI22_X1 U14660 ( .A1(n12305), .A2(n14973), .B1(n14979), .B2(
        P3_REG2_REG_26__SCAN_IN), .ZN(n12306) );
  OAI21_X1 U14661 ( .B1(n12545), .B2(n14906), .A(n12306), .ZN(n12307) );
  AOI21_X1 U14662 ( .B1(n12488), .B2(n14977), .A(n12307), .ZN(n12308) );
  OAI21_X1 U14663 ( .B1(n12309), .B2(n12486), .A(n12308), .ZN(P3_U3207) );
  XNOR2_X1 U14664 ( .A(n12310), .B(n12312), .ZN(n12493) );
  INV_X1 U14665 ( .A(n12493), .ZN(n12322) );
  INV_X1 U14666 ( .A(n12312), .ZN(n12314) );
  OAI211_X1 U14667 ( .C1(n7380), .C2(n12314), .A(n14961), .B(n12313), .ZN(
        n12316) );
  NAND2_X1 U14668 ( .A1(n12316), .A2(n12315), .ZN(n12492) );
  INV_X1 U14669 ( .A(n12317), .ZN(n12549) );
  AOI22_X1 U14670 ( .A1(n14979), .A2(P3_REG2_REG_25__SCAN_IN), .B1(n12318), 
        .B2(n14973), .ZN(n12319) );
  OAI21_X1 U14671 ( .B1(n12549), .B2(n14906), .A(n12319), .ZN(n12320) );
  AOI21_X1 U14672 ( .B1(n12492), .B2(n14977), .A(n12320), .ZN(n12321) );
  OAI21_X1 U14673 ( .B1(n12322), .B2(n12486), .A(n12321), .ZN(P3_U3208) );
  XNOR2_X1 U14674 ( .A(n12323), .B(n12326), .ZN(n12325) );
  AOI21_X1 U14675 ( .B1(n12325), .B2(n14961), .A(n12324), .ZN(n12497) );
  OAI21_X1 U14676 ( .B1(n6541), .B2(n12326), .A(n12294), .ZN(n12496) );
  NAND2_X1 U14677 ( .A1(n12496), .A2(n14941), .ZN(n12332) );
  INV_X1 U14678 ( .A(P3_REG2_REG_24__SCAN_IN), .ZN(n12328) );
  OAI22_X1 U14679 ( .A1(n14977), .A2(n12328), .B1(n12327), .B2(n14959), .ZN(
        n12329) );
  AOI21_X1 U14680 ( .B1(n12330), .B2(n14957), .A(n12329), .ZN(n12331) );
  OAI211_X1 U14681 ( .C1(n14979), .C2(n12497), .A(n12332), .B(n12331), .ZN(
        P3_U3209) );
  OAI21_X1 U14682 ( .B1(n12334), .B2(n12335), .A(n12333), .ZN(n12341) );
  XNOR2_X1 U14683 ( .A(n12336), .B(n12335), .ZN(n12338) );
  AOI21_X1 U14684 ( .B1(n12338), .B2(n14961), .A(n12337), .ZN(n12339) );
  OAI21_X1 U14685 ( .B1(n12341), .B2(n12340), .A(n12339), .ZN(n12500) );
  INV_X1 U14686 ( .A(n12500), .ZN(n12346) );
  INV_X1 U14687 ( .A(n12341), .ZN(n12501) );
  AOI22_X1 U14688 ( .A1(n14979), .A2(P3_REG2_REG_23__SCAN_IN), .B1(n14973), 
        .B2(n12342), .ZN(n12343) );
  OAI21_X1 U14689 ( .B1(n12554), .B2(n14906), .A(n12343), .ZN(n12344) );
  AOI21_X1 U14690 ( .B1(n12501), .B2(n14974), .A(n12344), .ZN(n12345) );
  OAI21_X1 U14691 ( .B1(n12346), .B2(n14979), .A(n12345), .ZN(P3_U3210) );
  NAND2_X1 U14692 ( .A1(n12361), .A2(n12347), .ZN(n12349) );
  NAND2_X1 U14693 ( .A1(n12349), .A2(n12348), .ZN(n12350) );
  XNOR2_X1 U14694 ( .A(n12350), .B(n12352), .ZN(n12505) );
  INV_X1 U14695 ( .A(n12505), .ZN(n12360) );
  XOR2_X1 U14696 ( .A(n12352), .B(n12351), .Z(n12354) );
  OAI21_X1 U14697 ( .B1(n12354), .B2(n14949), .A(n12353), .ZN(n12504) );
  INV_X1 U14698 ( .A(n12355), .ZN(n12558) );
  AOI22_X1 U14699 ( .A1(n14979), .A2(P3_REG2_REG_22__SCAN_IN), .B1(n14973), 
        .B2(n12356), .ZN(n12357) );
  OAI21_X1 U14700 ( .B1(n12558), .B2(n14906), .A(n12357), .ZN(n12358) );
  AOI21_X1 U14701 ( .B1(n12504), .B2(n14977), .A(n12358), .ZN(n12359) );
  OAI21_X1 U14702 ( .B1(n12486), .B2(n12360), .A(n12359), .ZN(P3_U3211) );
  XOR2_X1 U14703 ( .A(n12363), .B(n12361), .Z(n12509) );
  INV_X1 U14704 ( .A(n12509), .ZN(n12370) );
  XOR2_X1 U14705 ( .A(n12363), .B(n12362), .Z(n12365) );
  OAI21_X1 U14706 ( .B1(n12365), .B2(n14949), .A(n12364), .ZN(n12508) );
  AOI22_X1 U14707 ( .A1(n14979), .A2(P3_REG2_REG_21__SCAN_IN), .B1(n12366), 
        .B2(n14973), .ZN(n12367) );
  OAI21_X1 U14708 ( .B1(n12562), .B2(n14906), .A(n12367), .ZN(n12368) );
  AOI21_X1 U14709 ( .B1(n12508), .B2(n14977), .A(n12368), .ZN(n12369) );
  OAI21_X1 U14710 ( .B1(n12370), .B2(n12486), .A(n12369), .ZN(P3_U3212) );
  XNOR2_X1 U14711 ( .A(n12371), .B(n12379), .ZN(n12373) );
  OAI21_X1 U14712 ( .B1(n12373), .B2(n14949), .A(n12372), .ZN(n12513) );
  AOI22_X1 U14713 ( .A1(n14979), .A2(P3_REG2_REG_20__SCAN_IN), .B1(n14973), 
        .B2(n12374), .ZN(n12375) );
  OAI21_X1 U14714 ( .B1(n12566), .B2(n14906), .A(n12375), .ZN(n12383) );
  INV_X1 U14715 ( .A(n12376), .ZN(n12381) );
  NAND2_X1 U14716 ( .A1(n12378), .A2(n12377), .ZN(n12380) );
  AND2_X1 U14717 ( .A1(n12380), .A2(n12379), .ZN(n12512) );
  NOR3_X1 U14718 ( .A1(n12381), .A2(n12512), .A3(n12486), .ZN(n12382) );
  AOI211_X1 U14719 ( .C1(n14977), .C2(n12513), .A(n12383), .B(n12382), .ZN(
        n12384) );
  INV_X1 U14720 ( .A(n12384), .ZN(P3_U3213) );
  XNOR2_X1 U14721 ( .A(n12385), .B(n12387), .ZN(n12520) );
  XNOR2_X1 U14722 ( .A(n12386), .B(n12387), .ZN(n12389) );
  OAI21_X1 U14723 ( .B1(n12389), .B2(n14949), .A(n12388), .ZN(n12517) );
  AOI22_X1 U14724 ( .A1(n14979), .A2(P3_REG2_REG_19__SCAN_IN), .B1(n14973), 
        .B2(n12390), .ZN(n12391) );
  OAI21_X1 U14725 ( .B1(n12392), .B2(n14906), .A(n12391), .ZN(n12393) );
  AOI21_X1 U14726 ( .B1(n12517), .B2(n14977), .A(n12393), .ZN(n12394) );
  OAI21_X1 U14727 ( .B1(n12486), .B2(n12520), .A(n12394), .ZN(P3_U3214) );
  INV_X1 U14728 ( .A(n12395), .ZN(n12396) );
  AOI21_X1 U14729 ( .B1(n12398), .B2(n12397), .A(n12396), .ZN(n12522) );
  INV_X1 U14730 ( .A(n12522), .ZN(n12409) );
  INV_X1 U14731 ( .A(n12399), .ZN(n12400) );
  AOI21_X1 U14732 ( .B1(n12402), .B2(n12401), .A(n12400), .ZN(n12404) );
  OAI21_X1 U14733 ( .B1(n12404), .B2(n14949), .A(n12403), .ZN(n12521) );
  AOI22_X1 U14734 ( .A1(n14979), .A2(P3_REG2_REG_18__SCAN_IN), .B1(n14973), 
        .B2(n12405), .ZN(n12406) );
  OAI21_X1 U14735 ( .B1(n12571), .B2(n14906), .A(n12406), .ZN(n12407) );
  AOI21_X1 U14736 ( .B1(n12521), .B2(n14977), .A(n12407), .ZN(n12408) );
  OAI21_X1 U14737 ( .B1(n12409), .B2(n12486), .A(n12408), .ZN(P3_U3215) );
  OAI21_X1 U14738 ( .B1(n12412), .B2(n12411), .A(n12410), .ZN(n12526) );
  INV_X1 U14739 ( .A(n12526), .ZN(n12424) );
  AND2_X1 U14740 ( .A1(n12414), .A2(n12413), .ZN(n12417) );
  OAI211_X1 U14741 ( .C1(n12417), .C2(n12416), .A(n14961), .B(n12415), .ZN(
        n12419) );
  NAND2_X1 U14742 ( .A1(n12419), .A2(n12418), .ZN(n12525) );
  AOI22_X1 U14743 ( .A1(n14979), .A2(P3_REG2_REG_17__SCAN_IN), .B1(n14973), 
        .B2(n12420), .ZN(n12421) );
  OAI21_X1 U14744 ( .B1(n12575), .B2(n14906), .A(n12421), .ZN(n12422) );
  AOI21_X1 U14745 ( .B1(n12525), .B2(n14977), .A(n12422), .ZN(n12423) );
  OAI21_X1 U14746 ( .B1(n12424), .B2(n12486), .A(n12423), .ZN(P3_U3216) );
  XOR2_X1 U14747 ( .A(n12429), .B(n12425), .Z(n12427) );
  OAI21_X1 U14748 ( .B1(n12427), .B2(n14949), .A(n12426), .ZN(n12529) );
  INV_X1 U14749 ( .A(n12529), .ZN(n12435) );
  OAI21_X1 U14750 ( .B1(n12430), .B2(n12429), .A(n12428), .ZN(n12530) );
  AOI22_X1 U14751 ( .A1(n14979), .A2(P3_REG2_REG_16__SCAN_IN), .B1(n14973), 
        .B2(n12431), .ZN(n12432) );
  OAI21_X1 U14752 ( .B1(n12579), .B2(n14906), .A(n12432), .ZN(n12433) );
  AOI21_X1 U14753 ( .B1(n12530), .B2(n14941), .A(n12433), .ZN(n12434) );
  OAI21_X1 U14754 ( .B1(n12435), .B2(n14979), .A(n12434), .ZN(P3_U3217) );
  XNOR2_X1 U14755 ( .A(n12436), .B(n7149), .ZN(n12441) );
  AOI22_X1 U14756 ( .A1(n12440), .A2(n12439), .B1(n12438), .B2(n12437), .ZN(
        n14282) );
  OAI21_X1 U14757 ( .B1(n12441), .B2(n14949), .A(n14282), .ZN(n12533) );
  INV_X1 U14758 ( .A(n12533), .ZN(n12449) );
  OAI21_X1 U14759 ( .B1(n12444), .B2(n12443), .A(n12442), .ZN(n12534) );
  AOI22_X1 U14760 ( .A1(n14979), .A2(P3_REG2_REG_15__SCAN_IN), .B1(n14973), 
        .B2(n12445), .ZN(n12446) );
  OAI21_X1 U14761 ( .B1(n12584), .B2(n14906), .A(n12446), .ZN(n12447) );
  AOI21_X1 U14762 ( .B1(n12534), .B2(n14941), .A(n12447), .ZN(n12448) );
  OAI21_X1 U14763 ( .B1(n12449), .B2(n14979), .A(n12448), .ZN(P3_U3218) );
  XNOR2_X1 U14764 ( .A(n12450), .B(n12451), .ZN(n14296) );
  INV_X1 U14765 ( .A(n14296), .ZN(n12462) );
  XNOR2_X1 U14766 ( .A(n12452), .B(n12451), .ZN(n12454) );
  OAI21_X1 U14767 ( .B1(n12454), .B2(n14949), .A(n12453), .ZN(n14294) );
  NOR2_X1 U14768 ( .A1(n12455), .A2(n14298), .ZN(n14295) );
  INV_X1 U14769 ( .A(n14295), .ZN(n12459) );
  AOI22_X1 U14770 ( .A1(n14979), .A2(P3_REG2_REG_14__SCAN_IN), .B1(n14973), 
        .B2(n12456), .ZN(n12457) );
  OAI21_X1 U14771 ( .B1(n12459), .B2(n12458), .A(n12457), .ZN(n12460) );
  AOI21_X1 U14772 ( .B1(n14294), .B2(n14977), .A(n12460), .ZN(n12461) );
  OAI21_X1 U14773 ( .B1(n12486), .B2(n12462), .A(n12461), .ZN(P3_U3219) );
  XOR2_X1 U14774 ( .A(n12464), .B(n12463), .Z(n14302) );
  INV_X1 U14775 ( .A(n14302), .ZN(n12472) );
  XNOR2_X1 U14776 ( .A(n12465), .B(n12464), .ZN(n12467) );
  OAI21_X1 U14777 ( .B1(n12467), .B2(n14949), .A(n12466), .ZN(n14300) );
  AOI22_X1 U14778 ( .A1(n14979), .A2(P3_REG2_REG_13__SCAN_IN), .B1(n12468), 
        .B2(n14973), .ZN(n12469) );
  OAI21_X1 U14779 ( .B1(n14299), .B2(n14906), .A(n12469), .ZN(n12470) );
  AOI21_X1 U14780 ( .B1(n14300), .B2(n14977), .A(n12470), .ZN(n12471) );
  OAI21_X1 U14781 ( .B1(n12472), .B2(n12486), .A(n12471), .ZN(P3_U3220) );
  XNOR2_X1 U14782 ( .A(n12474), .B(n12473), .ZN(n14306) );
  INV_X1 U14783 ( .A(n14306), .ZN(n12487) );
  NOR2_X1 U14784 ( .A1(n12475), .A2(n14298), .ZN(n14305) );
  INV_X1 U14785 ( .A(n12476), .ZN(n12477) );
  OAI22_X1 U14786 ( .A1(n14977), .A2(n8264), .B1(n12477), .B2(n14959), .ZN(
        n12478) );
  AOI21_X1 U14787 ( .B1(n12479), .B2(n14305), .A(n12478), .ZN(n12485) );
  XNOR2_X1 U14788 ( .A(n12481), .B(n12480), .ZN(n12483) );
  OAI21_X1 U14789 ( .B1(n12483), .B2(n14949), .A(n12482), .ZN(n14304) );
  NAND2_X1 U14790 ( .A1(n14304), .A2(n14977), .ZN(n12484) );
  OAI211_X1 U14791 ( .C1(n12487), .C2(n12486), .A(n12485), .B(n12484), .ZN(
        P3_U3221) );
  INV_X1 U14792 ( .A(P3_REG1_REG_26__SCAN_IN), .ZN(n12490) );
  AOI21_X1 U14793 ( .B1(n12489), .B2(n14983), .A(n12488), .ZN(n12542) );
  MUX2_X1 U14794 ( .A(n12490), .B(n12542), .S(n15038), .Z(n12491) );
  OAI21_X1 U14795 ( .B1(n12545), .B2(n12537), .A(n12491), .ZN(P3_U3485) );
  INV_X1 U14796 ( .A(P3_REG1_REG_25__SCAN_IN), .ZN(n12494) );
  AOI21_X1 U14797 ( .B1(n12493), .B2(n14983), .A(n12492), .ZN(n12546) );
  MUX2_X1 U14798 ( .A(n12494), .B(n12546), .S(n15038), .Z(n12495) );
  OAI21_X1 U14799 ( .B1(n12549), .B2(n12537), .A(n12495), .ZN(P3_U3484) );
  NAND2_X1 U14800 ( .A1(n12496), .A2(n14983), .ZN(n12498) );
  OAI211_X1 U14801 ( .C1(n12499), .C2(n14298), .A(n12498), .B(n12497), .ZN(
        n12550) );
  MUX2_X1 U14802 ( .A(P3_REG1_REG_24__SCAN_IN), .B(n12550), .S(n15038), .Z(
        P3_U3483) );
  INV_X1 U14803 ( .A(P3_REG1_REG_23__SCAN_IN), .ZN(n12502) );
  AOI21_X1 U14804 ( .B1(n6604), .B2(n12501), .A(n12500), .ZN(n12551) );
  MUX2_X1 U14805 ( .A(n12502), .B(n12551), .S(n15038), .Z(n12503) );
  OAI21_X1 U14806 ( .B1(n12554), .B2(n12537), .A(n12503), .ZN(P3_U3482) );
  INV_X1 U14807 ( .A(P3_REG1_REG_22__SCAN_IN), .ZN(n12506) );
  AOI21_X1 U14808 ( .B1(n14983), .B2(n12505), .A(n12504), .ZN(n12555) );
  MUX2_X1 U14809 ( .A(n12506), .B(n12555), .S(n15038), .Z(n12507) );
  OAI21_X1 U14810 ( .B1(n12558), .B2(n12537), .A(n12507), .ZN(P3_U3481) );
  INV_X1 U14811 ( .A(P3_REG1_REG_21__SCAN_IN), .ZN(n12510) );
  AOI21_X1 U14812 ( .B1(n12509), .B2(n14983), .A(n12508), .ZN(n12559) );
  MUX2_X1 U14813 ( .A(n12510), .B(n12559), .S(n15038), .Z(n12511) );
  OAI21_X1 U14814 ( .B1(n12562), .B2(n12537), .A(n12511), .ZN(P3_U3480) );
  INV_X1 U14815 ( .A(P3_REG1_REG_20__SCAN_IN), .ZN(n12515) );
  NOR2_X1 U14816 ( .A1(n12512), .A2(n14989), .ZN(n12514) );
  AOI21_X1 U14817 ( .B1(n12514), .B2(n12376), .A(n12513), .ZN(n12563) );
  MUX2_X1 U14818 ( .A(n12515), .B(n12563), .S(n15038), .Z(n12516) );
  OAI21_X1 U14819 ( .B1(n12566), .B2(n12537), .A(n12516), .ZN(P3_U3479) );
  AOI21_X1 U14820 ( .B1(n15016), .B2(n12518), .A(n12517), .ZN(n12519) );
  OAI21_X1 U14821 ( .B1(n14989), .B2(n12520), .A(n12519), .ZN(n12567) );
  MUX2_X1 U14822 ( .A(P3_REG1_REG_19__SCAN_IN), .B(n12567), .S(n15038), .Z(
        P3_U3478) );
  AOI21_X1 U14823 ( .B1(n12522), .B2(n14983), .A(n12521), .ZN(n12568) );
  MUX2_X1 U14824 ( .A(n12523), .B(n12568), .S(n15038), .Z(n12524) );
  OAI21_X1 U14825 ( .B1(n12571), .B2(n12537), .A(n12524), .ZN(P3_U3477) );
  AOI21_X1 U14826 ( .B1(n12526), .B2(n14983), .A(n12525), .ZN(n12572) );
  MUX2_X1 U14827 ( .A(n12527), .B(n12572), .S(n15038), .Z(n12528) );
  OAI21_X1 U14828 ( .B1(n12575), .B2(n12537), .A(n12528), .ZN(P3_U3476) );
  AOI21_X1 U14829 ( .B1(n14983), .B2(n12530), .A(n12529), .ZN(n12576) );
  MUX2_X1 U14830 ( .A(n12531), .B(n12576), .S(n15038), .Z(n12532) );
  OAI21_X1 U14831 ( .B1(n12579), .B2(n12537), .A(n12532), .ZN(P3_U3475) );
  AOI21_X1 U14832 ( .B1(n14983), .B2(n12534), .A(n12533), .ZN(n12580) );
  MUX2_X1 U14833 ( .A(n12535), .B(n12580), .S(n15038), .Z(n12536) );
  OAI21_X1 U14834 ( .B1(n12584), .B2(n12537), .A(n12536), .ZN(P3_U3474) );
  INV_X1 U14835 ( .A(P3_REG0_REG_27__SCAN_IN), .ZN(n12539) );
  OAI21_X1 U14836 ( .B1(n12541), .B2(n12583), .A(n12540), .ZN(P3_U3454) );
  INV_X1 U14837 ( .A(P3_REG0_REG_26__SCAN_IN), .ZN(n12543) );
  MUX2_X1 U14838 ( .A(n12543), .B(n12542), .S(n15015), .Z(n12544) );
  OAI21_X1 U14839 ( .B1(n12545), .B2(n12583), .A(n12544), .ZN(P3_U3453) );
  INV_X1 U14840 ( .A(P3_REG0_REG_25__SCAN_IN), .ZN(n12547) );
  MUX2_X1 U14841 ( .A(n12547), .B(n12546), .S(n15015), .Z(n12548) );
  OAI21_X1 U14842 ( .B1(n12549), .B2(n12583), .A(n12548), .ZN(P3_U3452) );
  MUX2_X1 U14843 ( .A(P3_REG0_REG_24__SCAN_IN), .B(n12550), .S(n15015), .Z(
        P3_U3451) );
  INV_X1 U14844 ( .A(P3_REG0_REG_23__SCAN_IN), .ZN(n12552) );
  MUX2_X1 U14845 ( .A(n12552), .B(n12551), .S(n15015), .Z(n12553) );
  OAI21_X1 U14846 ( .B1(n12554), .B2(n12583), .A(n12553), .ZN(P3_U3450) );
  INV_X1 U14847 ( .A(P3_REG0_REG_22__SCAN_IN), .ZN(n12556) );
  MUX2_X1 U14848 ( .A(n12556), .B(n12555), .S(n15015), .Z(n12557) );
  OAI21_X1 U14849 ( .B1(n12558), .B2(n12583), .A(n12557), .ZN(P3_U3449) );
  INV_X1 U14850 ( .A(P3_REG0_REG_21__SCAN_IN), .ZN(n12560) );
  MUX2_X1 U14851 ( .A(n12560), .B(n12559), .S(n15015), .Z(n12561) );
  OAI21_X1 U14852 ( .B1(n12562), .B2(n12583), .A(n12561), .ZN(P3_U3448) );
  INV_X1 U14853 ( .A(P3_REG0_REG_20__SCAN_IN), .ZN(n12564) );
  MUX2_X1 U14854 ( .A(n12564), .B(n12563), .S(n15015), .Z(n12565) );
  OAI21_X1 U14855 ( .B1(n12566), .B2(n12583), .A(n12565), .ZN(P3_U3447) );
  MUX2_X1 U14856 ( .A(P3_REG0_REG_19__SCAN_IN), .B(n12567), .S(n15015), .Z(
        P3_U3446) );
  INV_X1 U14857 ( .A(P3_REG0_REG_18__SCAN_IN), .ZN(n12569) );
  MUX2_X1 U14858 ( .A(n12569), .B(n12568), .S(n15015), .Z(n12570) );
  OAI21_X1 U14859 ( .B1(n12571), .B2(n12583), .A(n12570), .ZN(P3_U3444) );
  INV_X1 U14860 ( .A(P3_REG0_REG_17__SCAN_IN), .ZN(n12573) );
  MUX2_X1 U14861 ( .A(n12573), .B(n12572), .S(n15015), .Z(n12574) );
  OAI21_X1 U14862 ( .B1(n12575), .B2(n12583), .A(n12574), .ZN(P3_U3441) );
  INV_X1 U14863 ( .A(P3_REG0_REG_16__SCAN_IN), .ZN(n12577) );
  MUX2_X1 U14864 ( .A(n12577), .B(n12576), .S(n15015), .Z(n12578) );
  OAI21_X1 U14865 ( .B1(n12579), .B2(n12583), .A(n12578), .ZN(P3_U3438) );
  INV_X1 U14866 ( .A(P3_REG0_REG_15__SCAN_IN), .ZN(n12581) );
  MUX2_X1 U14867 ( .A(n12581), .B(n12580), .S(n15015), .Z(n12582) );
  OAI21_X1 U14868 ( .B1(n12584), .B2(n12583), .A(n12582), .ZN(P3_U3435) );
  MUX2_X1 U14869 ( .A(n12585), .B(P3_D_REG_1__SCAN_IN), .S(n12586), .Z(
        P3_U3377) );
  MUX2_X1 U14870 ( .A(n12587), .B(P3_D_REG_0__SCAN_IN), .S(n12586), .Z(
        P3_U3376) );
  NAND3_X1 U14871 ( .A1(n12588), .A2(P3_STATE_REG_SCAN_IN), .A3(
        P3_IR_REG_31__SCAN_IN), .ZN(n12590) );
  OAI22_X1 U14872 ( .A1(n7554), .A2(n12590), .B1(n15074), .B2(n12589), .ZN(
        n12591) );
  AOI21_X1 U14873 ( .B1(n12592), .B2(n12596), .A(n12591), .ZN(n12593) );
  INV_X1 U14874 ( .A(n12593), .ZN(P3_U3264) );
  AOI222_X1 U14875 ( .A1(n12597), .A2(n12596), .B1(P3_STATE_REG_SCAN_IN), .B2(
        n12595), .C1(SI_29_), .C2(n12594), .ZN(n12598) );
  INV_X1 U14876 ( .A(n12598), .ZN(P3_U3266) );
  INV_X1 U14877 ( .A(n12599), .ZN(n12600) );
  OAI222_X1 U14878 ( .A1(n12607), .A2(n12600), .B1(P3_U3151), .B2(n7945), .C1(
        n15047), .C2(n12608), .ZN(P3_U3267) );
  INV_X1 U14879 ( .A(n12601), .ZN(n12603) );
  OAI222_X1 U14880 ( .A1(n12607), .A2(n12603), .B1(P3_U3151), .B2(n12602), 
        .C1(n15169), .C2(n12608), .ZN(P3_U3268) );
  INV_X1 U14881 ( .A(SI_26_), .ZN(n15084) );
  INV_X1 U14882 ( .A(n12604), .ZN(n12606) );
  OAI222_X1 U14883 ( .A1(n12608), .A2(n15084), .B1(n12607), .B2(n12606), .C1(
        n12605), .C2(P3_U3151), .ZN(P3_U3269) );
  XNOR2_X1 U14884 ( .A(n12610), .B(n12609), .ZN(n12617) );
  INV_X1 U14885 ( .A(n13191), .ZN(n12614) );
  NAND2_X1 U14886 ( .A1(n13040), .A2(n12711), .ZN(n12612) );
  NAND2_X1 U14887 ( .A1(n13042), .A2(n12710), .ZN(n12611) );
  NAND2_X1 U14888 ( .A1(n12612), .A2(n12611), .ZN(n13338) );
  AOI22_X1 U14889 ( .A1(n14330), .A2(n13338), .B1(P2_REG3_REG_27__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12613) );
  OAI21_X1 U14890 ( .B1(n12614), .B2(n14334), .A(n12613), .ZN(n12615) );
  AOI21_X1 U14891 ( .B1(n13339), .B2(n12703), .A(n12615), .ZN(n12616) );
  OAI21_X1 U14892 ( .B1(n12617), .B2(n12705), .A(n12616), .ZN(P2_U3186) );
  XNOR2_X1 U14893 ( .A(n12619), .B(n12618), .ZN(n12620) );
  XNOR2_X1 U14894 ( .A(n12621), .B(n12620), .ZN(n12627) );
  INV_X1 U14895 ( .A(n12622), .ZN(n13255) );
  OAI22_X1 U14896 ( .A1(n12623), .A2(n14324), .B1(n12898), .B2(n14322), .ZN(
        n13249) );
  AOI22_X1 U14897 ( .A1(n14330), .A2(n13249), .B1(P2_REG3_REG_23__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12624) );
  OAI21_X1 U14898 ( .B1(n13255), .B2(n14334), .A(n12624), .ZN(n12625) );
  AOI21_X1 U14899 ( .B1(n13363), .B2(n14331), .A(n12625), .ZN(n12626) );
  OAI21_X1 U14900 ( .B1(n12627), .B2(n12705), .A(n12626), .ZN(P2_U3188) );
  OAI21_X1 U14901 ( .B1(n12630), .B2(n12629), .A(n12628), .ZN(n12631) );
  NAND2_X1 U14902 ( .A1(n12631), .A2(n14328), .ZN(n12635) );
  NAND2_X1 U14903 ( .A1(P2_U3088), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n13159)
         );
  OAI21_X1 U14904 ( .B1(n13384), .B2(n12715), .A(n13159), .ZN(n12632) );
  AOI21_X1 U14905 ( .B1(n12633), .B2(n12717), .A(n12632), .ZN(n12634) );
  OAI211_X1 U14906 ( .C1(n6859), .C2(n12719), .A(n12635), .B(n12634), .ZN(
        P2_U3191) );
  XNOR2_X1 U14907 ( .A(n12637), .B(n12636), .ZN(n12642) );
  INV_X1 U14908 ( .A(n12638), .ZN(n13278) );
  OAI22_X1 U14909 ( .A1(n12879), .A2(n14322), .B1(n12898), .B2(n14324), .ZN(
        n13277) );
  AOI22_X1 U14910 ( .A1(n13277), .A2(n14330), .B1(P2_REG3_REG_21__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12639) );
  OAI21_X1 U14911 ( .B1(n13278), .B2(n14334), .A(n12639), .ZN(n12640) );
  AOI21_X1 U14912 ( .B1(n12885), .B2(n12703), .A(n12640), .ZN(n12641) );
  OAI21_X1 U14913 ( .B1(n12642), .B2(n12705), .A(n12641), .ZN(P2_U3195) );
  XNOR2_X1 U14914 ( .A(n12644), .B(n12643), .ZN(n12651) );
  INV_X1 U14915 ( .A(n13216), .ZN(n12648) );
  NAND2_X1 U14916 ( .A1(n13044), .A2(n12710), .ZN(n12646) );
  NAND2_X1 U14917 ( .A1(n13042), .A2(n12711), .ZN(n12645) );
  NAND2_X1 U14918 ( .A1(n12646), .A2(n12645), .ZN(n13351) );
  AOI22_X1 U14919 ( .A1(n14330), .A2(n13351), .B1(P2_REG3_REG_25__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12647) );
  OAI21_X1 U14920 ( .B1(n12648), .B2(n14334), .A(n12647), .ZN(n12649) );
  AOI21_X1 U14921 ( .B1(n13352), .B2(n14331), .A(n12649), .ZN(n12650) );
  OAI21_X1 U14922 ( .B1(n12651), .B2(n12705), .A(n12650), .ZN(P2_U3197) );
  AOI21_X1 U14923 ( .B1(n12654), .B2(n12653), .A(n12652), .ZN(n12661) );
  NOR2_X1 U14924 ( .A1(n14334), .A2(n12655), .ZN(n12659) );
  OAI21_X1 U14925 ( .B1(n12715), .B2(n12657), .A(n12656), .ZN(n12658) );
  AOI211_X1 U14926 ( .C1(n13404), .C2(n14331), .A(n12659), .B(n12658), .ZN(
        n12660) );
  OAI21_X1 U14927 ( .B1(n12661), .B2(n12705), .A(n12660), .ZN(P2_U3198) );
  AOI21_X1 U14928 ( .B1(n12664), .B2(n12663), .A(n12662), .ZN(n12670) );
  NOR2_X1 U14929 ( .A1(n14334), .A2(n12665), .ZN(n12668) );
  OAI21_X1 U14930 ( .B1(n12715), .B2(n13395), .A(n12666), .ZN(n12667) );
  AOI211_X1 U14931 ( .C1(n12851), .C2(n14331), .A(n12668), .B(n12667), .ZN(
        n12669) );
  OAI21_X1 U14932 ( .B1(n12670), .B2(n12705), .A(n12669), .ZN(P2_U3200) );
  XNOR2_X1 U14933 ( .A(n12672), .B(n12671), .ZN(n12678) );
  INV_X1 U14934 ( .A(n12673), .ZN(n13234) );
  OAI22_X1 U14935 ( .A1(n12674), .A2(n14324), .B1(n12691), .B2(n14322), .ZN(
        n13228) );
  AOI22_X1 U14936 ( .A1(n14330), .A2(n13228), .B1(P2_REG3_REG_24__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12675) );
  OAI21_X1 U14937 ( .B1(n13234), .B2(n14334), .A(n12675), .ZN(n12676) );
  AOI21_X1 U14938 ( .B1(n13358), .B2(n14331), .A(n12676), .ZN(n12677) );
  OAI21_X1 U14939 ( .B1(n12678), .B2(n12705), .A(n12677), .ZN(P2_U3201) );
  OAI21_X1 U14940 ( .B1(n12681), .B2(n12680), .A(n12679), .ZN(n12682) );
  NAND2_X1 U14941 ( .A1(n12682), .A2(n14328), .ZN(n12687) );
  INV_X1 U14942 ( .A(n13294), .ZN(n12685) );
  AOI22_X1 U14943 ( .A1(n13047), .A2(n12711), .B1(n12710), .B2(n13049), .ZN(
        n13290) );
  OAI22_X1 U14944 ( .A1(n13290), .A2(n12715), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12683), .ZN(n12684) );
  AOI21_X1 U14945 ( .B1(n12685), .B2(n12717), .A(n12684), .ZN(n12686) );
  OAI211_X1 U14946 ( .C1(n12688), .C2(n12719), .A(n12687), .B(n12686), .ZN(
        P2_U3205) );
  XNOR2_X1 U14947 ( .A(n12690), .B(n12689), .ZN(n12697) );
  INV_X1 U14948 ( .A(n13265), .ZN(n12694) );
  OAI22_X1 U14949 ( .A1(n12692), .A2(n14322), .B1(n12691), .B2(n14324), .ZN(
        n13261) );
  AOI22_X1 U14950 ( .A1(n13261), .A2(n14330), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3088), .ZN(n12693) );
  OAI21_X1 U14951 ( .B1(n12694), .B2(n14334), .A(n12693), .ZN(n12695) );
  AOI21_X1 U14952 ( .B1(n13368), .B2(n14331), .A(n12695), .ZN(n12696) );
  OAI21_X1 U14953 ( .B1(n12697), .B2(n12705), .A(n12696), .ZN(P2_U3207) );
  XNOR2_X1 U14954 ( .A(n12699), .B(n12698), .ZN(n12706) );
  OAI22_X1 U14955 ( .A1(n12700), .A2(n14324), .B1(n12853), .B2(n14322), .ZN(
        n13310) );
  NAND2_X1 U14956 ( .A1(n14330), .A2(n13310), .ZN(n12701) );
  NAND2_X1 U14957 ( .A1(P2_U3088), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n13133)
         );
  OAI211_X1 U14958 ( .C1(n14334), .C2(n13315), .A(n12701), .B(n13133), .ZN(
        n12702) );
  AOI21_X1 U14959 ( .B1(n13390), .B2(n12703), .A(n12702), .ZN(n12704) );
  OAI21_X1 U14960 ( .B1(n12706), .B2(n12705), .A(n12704), .ZN(P2_U3210) );
  OAI21_X1 U14961 ( .B1(n6536), .B2(n12708), .A(n12707), .ZN(n12709) );
  NAND2_X1 U14962 ( .A1(n13043), .A2(n12710), .ZN(n12713) );
  NAND2_X1 U14963 ( .A1(n13041), .A2(n12711), .ZN(n12712) );
  AND2_X1 U14964 ( .A1(n12713), .A2(n12712), .ZN(n13343) );
  OAI22_X1 U14965 ( .A1(n12715), .A2(n13343), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n12714), .ZN(n12716) );
  AOI21_X1 U14966 ( .B1(n13204), .B2(n12717), .A(n12716), .ZN(n12718) );
  NAND2_X1 U14967 ( .A1(n6477), .A2(n14743), .ZN(n12724) );
  NAND2_X1 U14968 ( .A1(n12723), .A2(n12722), .ZN(n12727) );
  NAND2_X1 U14969 ( .A1(n12724), .A2(n12727), .ZN(n12726) );
  NAND2_X1 U14970 ( .A1(n12726), .A2(n12725), .ZN(n12730) );
  INV_X1 U14971 ( .A(n12727), .ZN(n12728) );
  NAND2_X1 U14972 ( .A1(n12728), .A2(n14743), .ZN(n12729) );
  AOI22_X1 U14973 ( .A1(n6477), .A2(n13067), .B1(n12932), .B2(n12732), .ZN(
        n12737) );
  NAND2_X1 U14974 ( .A1(n6477), .A2(n12732), .ZN(n12733) );
  NAND2_X1 U14975 ( .A1(n12734), .A2(n12733), .ZN(n12735) );
  NAND2_X1 U14976 ( .A1(n12737), .A2(n12736), .ZN(n12744) );
  NAND2_X1 U14977 ( .A1(n6477), .A2(n12740), .ZN(n12739) );
  NAND2_X1 U14978 ( .A1(n13066), .A2(n12932), .ZN(n12738) );
  NAND2_X1 U14979 ( .A1(n12739), .A2(n12738), .ZN(n12746) );
  AND2_X1 U14980 ( .A1(n12742), .A2(n12741), .ZN(n12747) );
  NAND2_X1 U14981 ( .A1(n12746), .A2(n12747), .ZN(n12743) );
  NAND3_X1 U14982 ( .A1(n12745), .A2(n12744), .A3(n12743), .ZN(n12751) );
  INV_X1 U14983 ( .A(n12746), .ZN(n12749) );
  INV_X1 U14984 ( .A(n12747), .ZN(n12748) );
  NAND2_X1 U14985 ( .A1(n12749), .A2(n12748), .ZN(n12750) );
  NAND2_X1 U14986 ( .A1(n6477), .A2(n13065), .ZN(n12753) );
  NAND2_X1 U14987 ( .A1(n12759), .A2(n12772), .ZN(n12752) );
  NAND2_X1 U14988 ( .A1(n12753), .A2(n12752), .ZN(n12758) );
  AOI22_X1 U14989 ( .A1(n12754), .A2(n12772), .B1(n6477), .B2(n13064), .ZN(
        n12765) );
  INV_X2 U14990 ( .A(n12976), .ZN(n12949) );
  NAND2_X1 U14991 ( .A1(n12949), .A2(n13064), .ZN(n12756) );
  NAND2_X1 U14992 ( .A1(n12754), .A2(n6477), .ZN(n12755) );
  NAND2_X1 U14993 ( .A1(n12756), .A2(n12755), .ZN(n12764) );
  NAND2_X1 U14994 ( .A1(n12765), .A2(n12764), .ZN(n12757) );
  AOI22_X1 U14995 ( .A1(n6477), .A2(n12759), .B1(n12949), .B2(n13065), .ZN(
        n12760) );
  INV_X1 U14996 ( .A(n12760), .ZN(n12761) );
  NAND2_X1 U14997 ( .A1(n12762), .A2(n12761), .ZN(n12763) );
  NAND2_X1 U14998 ( .A1(n6560), .A2(n12763), .ZN(n12769) );
  INV_X1 U14999 ( .A(n12764), .ZN(n12767) );
  INV_X1 U15000 ( .A(n12765), .ZN(n12766) );
  NAND2_X1 U15001 ( .A1(n12767), .A2(n12766), .ZN(n12768) );
  NAND2_X1 U15002 ( .A1(n12769), .A2(n12768), .ZN(n12780) );
  NAND2_X1 U15003 ( .A1(n12773), .A2(n12949), .ZN(n12771) );
  NAND2_X1 U15004 ( .A1(n6477), .A2(n13063), .ZN(n12770) );
  NAND2_X1 U15005 ( .A1(n12771), .A2(n12770), .ZN(n12779) );
  AOI22_X1 U15006 ( .A1(n12773), .A2(n12959), .B1(n12949), .B2(n13063), .ZN(
        n12774) );
  AOI21_X1 U15007 ( .B1(n12780), .B2(n12779), .A(n12774), .ZN(n12785) );
  AND2_X1 U15008 ( .A1(n12932), .A2(n13062), .ZN(n12775) );
  NAND2_X1 U15009 ( .A1(n12776), .A2(n12949), .ZN(n12778) );
  NAND2_X1 U15010 ( .A1(n6477), .A2(n13062), .ZN(n12777) );
  NAND2_X1 U15011 ( .A1(n12778), .A2(n12777), .ZN(n12781) );
  OAI22_X1 U15012 ( .A1(n12780), .A2(n12779), .B1(n12782), .B2(n12781), .ZN(
        n12784) );
  NAND2_X1 U15013 ( .A1(n12782), .A2(n12781), .ZN(n12783) );
  NAND2_X1 U15014 ( .A1(n12791), .A2(n12949), .ZN(n12787) );
  NAND2_X1 U15015 ( .A1(n12959), .A2(n13061), .ZN(n12786) );
  NAND2_X1 U15016 ( .A1(n12787), .A2(n12786), .ZN(n12793) );
  AND2_X1 U15017 ( .A1(n12932), .A2(n13060), .ZN(n12788) );
  AOI21_X1 U15018 ( .B1(n14781), .B2(n12959), .A(n12788), .ZN(n12796) );
  NAND2_X1 U15019 ( .A1(n14781), .A2(n12949), .ZN(n12790) );
  NAND2_X1 U15020 ( .A1(n6477), .A2(n13060), .ZN(n12789) );
  NAND2_X1 U15021 ( .A1(n12790), .A2(n12789), .ZN(n12795) );
  OAI22_X1 U15022 ( .A1(n12794), .A2(n12793), .B1(n12796), .B2(n12795), .ZN(
        n12798) );
  AOI22_X1 U15023 ( .A1(n12791), .A2(n12959), .B1(n12949), .B2(n13061), .ZN(
        n12792) );
  AOI21_X1 U15024 ( .B1(n12794), .B2(n12793), .A(n12792), .ZN(n12797) );
  NAND2_X1 U15025 ( .A1(n12801), .A2(n12949), .ZN(n12800) );
  NAND2_X1 U15026 ( .A1(n12959), .A2(n13059), .ZN(n12799) );
  NAND2_X1 U15027 ( .A1(n12800), .A2(n12799), .ZN(n12803) );
  AOI22_X1 U15028 ( .A1(n12801), .A2(n12959), .B1(n12772), .B2(n13059), .ZN(
        n12802) );
  NAND2_X1 U15029 ( .A1(n14789), .A2(n12959), .ZN(n12805) );
  NAND2_X1 U15030 ( .A1(n12949), .A2(n13058), .ZN(n12804) );
  NAND2_X1 U15031 ( .A1(n12805), .A2(n12804), .ZN(n12807) );
  AOI22_X1 U15032 ( .A1(n14789), .A2(n12772), .B1(n12959), .B2(n13058), .ZN(
        n12806) );
  NAND2_X1 U15033 ( .A1(n12810), .A2(n12772), .ZN(n12809) );
  NAND2_X1 U15034 ( .A1(n12959), .A2(n13057), .ZN(n12808) );
  NAND2_X1 U15035 ( .A1(n12809), .A2(n12808), .ZN(n12816) );
  NAND2_X1 U15036 ( .A1(n12815), .A2(n12816), .ZN(n12814) );
  NAND2_X1 U15037 ( .A1(n12810), .A2(n6477), .ZN(n12811) );
  NAND2_X1 U15038 ( .A1(n12814), .A2(n12813), .ZN(n12820) );
  INV_X1 U15039 ( .A(n12815), .ZN(n12818) );
  NAND2_X1 U15040 ( .A1(n12818), .A2(n12817), .ZN(n12819) );
  NAND2_X1 U15041 ( .A1(n12820), .A2(n12819), .ZN(n12827) );
  NAND2_X1 U15042 ( .A1(n12823), .A2(n12959), .ZN(n12822) );
  NAND2_X1 U15043 ( .A1(n12949), .A2(n13056), .ZN(n12821) );
  NAND2_X1 U15044 ( .A1(n12822), .A2(n12821), .ZN(n12826) );
  AOI22_X1 U15045 ( .A1(n12823), .A2(n12949), .B1(n6477), .B2(n13056), .ZN(
        n12824) );
  NAND2_X1 U15046 ( .A1(n12830), .A2(n12772), .ZN(n12829) );
  NAND2_X1 U15047 ( .A1(n6477), .A2(n13055), .ZN(n12828) );
  NAND2_X1 U15048 ( .A1(n12830), .A2(n6477), .ZN(n12831) );
  OAI21_X1 U15049 ( .B1(n14323), .B2(n6477), .A(n12831), .ZN(n12832) );
  NAND2_X1 U15050 ( .A1(n14342), .A2(n12959), .ZN(n12834) );
  NAND2_X1 U15051 ( .A1(n12949), .A2(n13054), .ZN(n12833) );
  NAND2_X1 U15052 ( .A1(n12834), .A2(n12833), .ZN(n12836) );
  AOI22_X1 U15053 ( .A1(n14342), .A2(n12949), .B1(n12959), .B2(n13054), .ZN(
        n12835) );
  AOI21_X1 U15054 ( .B1(n12837), .B2(n12836), .A(n12835), .ZN(n12839) );
  NOR2_X1 U15055 ( .A1(n12837), .A2(n12836), .ZN(n12838) );
  OR2_X1 U15056 ( .A1(n12839), .A2(n12838), .ZN(n12845) );
  NAND2_X1 U15057 ( .A1(n12842), .A2(n12772), .ZN(n12841) );
  NAND2_X1 U15058 ( .A1(n12959), .A2(n13053), .ZN(n12840) );
  NAND2_X1 U15059 ( .A1(n12841), .A2(n12840), .ZN(n12844) );
  AOI22_X1 U15060 ( .A1(n12842), .A2(n12959), .B1(n12772), .B2(n13053), .ZN(
        n12843) );
  NAND2_X1 U15061 ( .A1(n13404), .A2(n12959), .ZN(n12847) );
  NAND2_X1 U15062 ( .A1(n13052), .A2(n12772), .ZN(n12846) );
  AOI22_X1 U15063 ( .A1(n13404), .A2(n12772), .B1(n12959), .B2(n13052), .ZN(
        n12848) );
  AND2_X1 U15064 ( .A1(n13051), .A2(n12959), .ZN(n12849) );
  AOI21_X1 U15065 ( .B1(n12851), .B2(n12949), .A(n12849), .ZN(n12857) );
  INV_X1 U15066 ( .A(n12857), .ZN(n12850) );
  NAND2_X1 U15067 ( .A1(n12856), .A2(n12850), .ZN(n12855) );
  NAND2_X1 U15068 ( .A1(n12851), .A2(n12959), .ZN(n12852) );
  NAND2_X1 U15069 ( .A1(n12855), .A2(n12854), .ZN(n12860) );
  INV_X1 U15070 ( .A(n12856), .ZN(n12858) );
  NAND2_X1 U15071 ( .A1(n12858), .A2(n12857), .ZN(n12859) );
  NAND2_X1 U15072 ( .A1(n12860), .A2(n12859), .ZN(n12867) );
  AND2_X1 U15073 ( .A1(n13050), .A2(n12932), .ZN(n12861) );
  AOI21_X1 U15074 ( .B1(n13390), .B2(n12959), .A(n12861), .ZN(n12868) );
  INV_X1 U15075 ( .A(n12868), .ZN(n12862) );
  NAND2_X1 U15076 ( .A1(n12867), .A2(n12862), .ZN(n12866) );
  NAND2_X1 U15077 ( .A1(n13390), .A2(n12949), .ZN(n12864) );
  NAND2_X1 U15078 ( .A1(n13050), .A2(n12959), .ZN(n12863) );
  NAND2_X1 U15079 ( .A1(n12864), .A2(n12863), .ZN(n12865) );
  INV_X1 U15080 ( .A(n12867), .ZN(n12869) );
  NAND2_X1 U15081 ( .A1(n12869), .A2(n12868), .ZN(n12870) );
  NAND2_X1 U15082 ( .A1(n12873), .A2(n12949), .ZN(n12872) );
  NAND2_X1 U15083 ( .A1(n13049), .A2(n6477), .ZN(n12871) );
  NAND2_X1 U15084 ( .A1(n12872), .A2(n12871), .ZN(n12875) );
  AOI22_X1 U15085 ( .A1(n12873), .A2(n12959), .B1(n12772), .B2(n13049), .ZN(
        n12874) );
  NAND2_X1 U15086 ( .A1(n13380), .A2(n12959), .ZN(n12877) );
  NAND2_X1 U15087 ( .A1(n13048), .A2(n12772), .ZN(n12876) );
  NAND2_X1 U15088 ( .A1(n12877), .A2(n12876), .ZN(n12882) );
  NAND2_X1 U15089 ( .A1(n13380), .A2(n12772), .ZN(n12878) );
  OAI21_X1 U15090 ( .B1(n12772), .B2(n12879), .A(n12878), .ZN(n12880) );
  NAND2_X1 U15091 ( .A1(n12885), .A2(n12949), .ZN(n12884) );
  NAND2_X1 U15092 ( .A1(n13047), .A2(n12959), .ZN(n12883) );
  NAND2_X1 U15093 ( .A1(n12884), .A2(n12883), .ZN(n12890) );
  AOI22_X1 U15094 ( .A1(n12885), .A2(n12959), .B1(n12949), .B2(n13047), .ZN(
        n12886) );
  INV_X1 U15095 ( .A(n12886), .ZN(n12887) );
  NAND2_X1 U15096 ( .A1(n12888), .A2(n12887), .ZN(n12894) );
  NAND2_X1 U15097 ( .A1(n12892), .A2(n12891), .ZN(n12893) );
  NAND2_X1 U15098 ( .A1(n13368), .A2(n12959), .ZN(n12896) );
  NAND2_X1 U15099 ( .A1(n12949), .A2(n13046), .ZN(n12895) );
  NAND2_X1 U15100 ( .A1(n13368), .A2(n12772), .ZN(n12897) );
  OAI21_X1 U15101 ( .B1(n12772), .B2(n12898), .A(n12897), .ZN(n12899) );
  NAND2_X1 U15102 ( .A1(n13363), .A2(n12949), .ZN(n12901) );
  NAND2_X1 U15103 ( .A1(n12959), .A2(n13045), .ZN(n12900) );
  NAND2_X1 U15104 ( .A1(n12901), .A2(n12900), .ZN(n12903) );
  AOI22_X1 U15105 ( .A1(n13363), .A2(n12959), .B1(n12772), .B2(n13045), .ZN(
        n12902) );
  NAND2_X1 U15106 ( .A1(n13358), .A2(n12959), .ZN(n12905) );
  NAND2_X1 U15107 ( .A1(n12949), .A2(n13044), .ZN(n12904) );
  NAND2_X1 U15108 ( .A1(n12905), .A2(n12904), .ZN(n12907) );
  AOI22_X1 U15109 ( .A1(n13358), .A2(n12772), .B1(n12959), .B2(n13044), .ZN(
        n12906) );
  AOI21_X1 U15110 ( .B1(n12908), .B2(n12907), .A(n12906), .ZN(n12910) );
  NOR2_X1 U15111 ( .A1(n12908), .A2(n12907), .ZN(n12909) );
  NAND2_X1 U15112 ( .A1(n13352), .A2(n12949), .ZN(n12912) );
  NAND2_X1 U15113 ( .A1(n12959), .A2(n13043), .ZN(n12911) );
  NAND2_X1 U15114 ( .A1(n12912), .A2(n12911), .ZN(n12914) );
  AOI22_X1 U15115 ( .A1(n13352), .A2(n12959), .B1(n12932), .B2(n13043), .ZN(
        n12913) );
  AND2_X1 U15116 ( .A1(n12932), .A2(n13042), .ZN(n12916) );
  AOI21_X1 U15117 ( .B1(n12922), .B2(n12959), .A(n12916), .ZN(n12920) );
  NAND2_X1 U15118 ( .A1(n12919), .A2(n12920), .ZN(n12954) );
  NAND2_X1 U15119 ( .A1(n13339), .A2(n12959), .ZN(n12918) );
  NAND2_X1 U15120 ( .A1(n12949), .A2(n13041), .ZN(n12917) );
  NAND2_X1 U15121 ( .A1(n12918), .A2(n12917), .ZN(n12947) );
  AND2_X1 U15122 ( .A1(n12954), .A2(n12947), .ZN(n12952) );
  INV_X1 U15123 ( .A(n12920), .ZN(n12921) );
  NAND2_X1 U15124 ( .A1(n12922), .A2(n12772), .ZN(n12924) );
  NAND2_X1 U15125 ( .A1(n12959), .A2(n13042), .ZN(n12923) );
  NAND2_X1 U15126 ( .A1(n12924), .A2(n12923), .ZN(n12925) );
  NAND2_X1 U15127 ( .A1(n12926), .A2(n12925), .ZN(n12956) );
  AND2_X1 U15128 ( .A1(n12932), .A2(n13040), .ZN(n12927) );
  AOI21_X1 U15129 ( .B1(n13331), .B2(n12959), .A(n12927), .ZN(n12969) );
  NAND2_X1 U15130 ( .A1(n13331), .A2(n12772), .ZN(n12929) );
  NAND2_X1 U15131 ( .A1(n12959), .A2(n13040), .ZN(n12928) );
  NAND2_X1 U15132 ( .A1(n12929), .A2(n12928), .ZN(n12968) );
  NAND2_X1 U15133 ( .A1(n9097), .A2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12930) );
  AND2_X1 U15134 ( .A1(n12932), .A2(n13038), .ZN(n12933) );
  AOI21_X1 U15135 ( .B1(n13161), .B2(n12959), .A(n12933), .ZN(n12963) );
  INV_X1 U15136 ( .A(n13038), .ZN(n12939) );
  OAI21_X1 U15137 ( .B1(n12935), .B2(n13026), .A(n12934), .ZN(n12936) );
  AOI21_X1 U15138 ( .B1(n12959), .B2(n13164), .A(n12936), .ZN(n12938) );
  NAND2_X1 U15139 ( .A1(n13161), .A2(n12772), .ZN(n12937) );
  OAI21_X1 U15140 ( .B1(n12939), .B2(n12938), .A(n12937), .ZN(n12962) );
  AND2_X1 U15141 ( .A1(n12959), .A2(n13039), .ZN(n12940) );
  AOI21_X1 U15142 ( .B1(n13327), .B2(n12949), .A(n12940), .ZN(n12965) );
  NAND2_X1 U15143 ( .A1(n13327), .A2(n12959), .ZN(n12942) );
  NAND2_X1 U15144 ( .A1(n12772), .A2(n13039), .ZN(n12941) );
  NAND2_X1 U15145 ( .A1(n12942), .A2(n12941), .ZN(n12964) );
  NAND2_X1 U15146 ( .A1(n12965), .A2(n12964), .ZN(n12970) );
  NAND2_X1 U15147 ( .A1(n12944), .A2(n12943), .ZN(n12946) );
  NAND2_X1 U15148 ( .A1(n9097), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(n12945) );
  INV_X1 U15149 ( .A(n12947), .ZN(n12951) );
  AND2_X1 U15150 ( .A1(n12959), .A2(n13041), .ZN(n12948) );
  AOI21_X1 U15151 ( .B1(n13339), .B2(n12949), .A(n12948), .ZN(n12953) );
  INV_X1 U15152 ( .A(n12953), .ZN(n12950) );
  NAND2_X1 U15153 ( .A1(n12956), .A2(n12955), .ZN(n12957) );
  NAND2_X1 U15154 ( .A1(n12958), .A2(n12957), .ZN(n12985) );
  MUX2_X1 U15155 ( .A(n13164), .B(n12949), .S(n12975), .Z(n12961) );
  NAND2_X1 U15156 ( .A1(n12949), .A2(n13164), .ZN(n12960) );
  NAND2_X1 U15157 ( .A1(n12961), .A2(n12960), .ZN(n12973) );
  INV_X1 U15158 ( .A(n12962), .ZN(n12967) );
  INV_X1 U15159 ( .A(n12963), .ZN(n12966) );
  OAI22_X1 U15160 ( .A1(n12967), .A2(n12966), .B1(n12965), .B2(n12964), .ZN(
        n12972) );
  AND3_X1 U15161 ( .A1(n12970), .A2(n12969), .A3(n12968), .ZN(n12971) );
  AOI22_X1 U15162 ( .A1(n12973), .A2(n12972), .B1(n12971), .B2(n12994), .ZN(
        n12982) );
  INV_X1 U15163 ( .A(n12974), .ZN(n12981) );
  INV_X1 U15164 ( .A(n13164), .ZN(n12977) );
  OR3_X1 U15165 ( .A1(n12975), .A2(n12977), .A3(n12959), .ZN(n12979) );
  NAND3_X1 U15166 ( .A1(n12975), .A2(n12977), .A3(n6477), .ZN(n12978) );
  AND2_X1 U15167 ( .A1(n12979), .A2(n12978), .ZN(n12980) );
  OAI21_X1 U15168 ( .B1(n12982), .B2(n12981), .A(n12980), .ZN(n12983) );
  AOI21_X1 U15169 ( .B1(n12720), .B2(n8952), .A(n13253), .ZN(n12986) );
  INV_X1 U15170 ( .A(n12986), .ZN(n12987) );
  NOR2_X1 U15171 ( .A1(n13030), .A2(n7478), .ZN(n12991) );
  OAI21_X1 U15172 ( .B1(n13031), .B2(n9327), .A(n12988), .ZN(n12989) );
  NAND3_X1 U15173 ( .A1(n12992), .A2(n12991), .A3(n12990), .ZN(n13037) );
  INV_X1 U15174 ( .A(n12994), .ZN(n13024) );
  XOR2_X1 U15175 ( .A(n13038), .B(n13161), .Z(n13023) );
  NOR4_X1 U15176 ( .A1(n14748), .A2(n12995), .A3(n9101), .A4(n8952), .ZN(
        n12997) );
  NAND4_X1 U15177 ( .A1(n12998), .A2(n12997), .A3(n12996), .A4(n14701), .ZN(
        n12999) );
  NOR4_X1 U15178 ( .A1(n13002), .A2(n13001), .A3(n13000), .A4(n12999), .ZN(
        n13003) );
  NAND4_X1 U15179 ( .A1(n13006), .A2(n13005), .A3(n13004), .A4(n13003), .ZN(
        n13007) );
  NOR4_X1 U15180 ( .A1(n14336), .A2(n13009), .A3(n13008), .A4(n13007), .ZN(
        n13014) );
  NAND4_X1 U15181 ( .A1(n13014), .A2(n13013), .A3(n13012), .A4(n13011), .ZN(
        n13015) );
  NOR4_X1 U15182 ( .A1(n13017), .A2(n13307), .A3(n13016), .A4(n13015), .ZN(
        n13018) );
  NAND3_X1 U15183 ( .A1(n13260), .A2(n13018), .A3(n13274), .ZN(n13019) );
  NOR4_X1 U15184 ( .A1(n13200), .A2(n13231), .A3(n13247), .A4(n13019), .ZN(
        n13020) );
  NAND4_X1 U15185 ( .A1(n13173), .A2(n13020), .A3(n13189), .A4(n13215), .ZN(
        n13021) );
  NOR4_X1 U15186 ( .A1(n13024), .A2(n13023), .A3(n13022), .A4(n13021), .ZN(
        n13033) );
  NOR4_X1 U15187 ( .A1(n13033), .A2(n8931), .A3(n13253), .A4(n13030), .ZN(
        n13025) );
  OAI21_X1 U15188 ( .B1(n12993), .B2(n13026), .A(n13025), .ZN(n13036) );
  NOR2_X1 U15189 ( .A1(n14322), .A2(n13432), .ZN(n13028) );
  NAND3_X1 U15190 ( .A1(n14736), .A2(n13028), .A3(n13027), .ZN(n13029) );
  OAI211_X1 U15191 ( .C1(n13031), .C2(n13030), .A(n13029), .B(P2_B_REG_SCAN_IN), .ZN(n13035) );
  NAND4_X1 U15192 ( .A1(n13033), .A2(n13032), .A3(n13253), .A4(n14742), .ZN(
        n13034) );
  NAND4_X1 U15193 ( .A1(n13037), .A2(n13036), .A3(n13035), .A4(n13034), .ZN(
        P2_U3328) );
  MUX2_X1 U15194 ( .A(P2_DATAO_REG_30__SCAN_IN), .B(n13038), .S(n6471), .Z(
        P2_U3561) );
  MUX2_X1 U15195 ( .A(P2_DATAO_REG_29__SCAN_IN), .B(n13039), .S(n6471), .Z(
        P2_U3560) );
  MUX2_X1 U15196 ( .A(P2_DATAO_REG_28__SCAN_IN), .B(n13040), .S(n6471), .Z(
        P2_U3559) );
  MUX2_X1 U15197 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n13041), .S(n6471), .Z(
        P2_U3558) );
  MUX2_X1 U15198 ( .A(P2_DATAO_REG_26__SCAN_IN), .B(n13042), .S(n6471), .Z(
        P2_U3557) );
  MUX2_X1 U15199 ( .A(P2_DATAO_REG_25__SCAN_IN), .B(n13043), .S(n6471), .Z(
        P2_U3556) );
  MUX2_X1 U15200 ( .A(P2_DATAO_REG_24__SCAN_IN), .B(n13044), .S(n6471), .Z(
        P2_U3555) );
  MUX2_X1 U15201 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n13045), .S(n6471), .Z(
        P2_U3554) );
  MUX2_X1 U15202 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n13046), .S(n6471), .Z(
        P2_U3553) );
  MUX2_X1 U15203 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n13047), .S(n6471), .Z(
        P2_U3552) );
  MUX2_X1 U15204 ( .A(P2_DATAO_REG_20__SCAN_IN), .B(n13048), .S(n6471), .Z(
        P2_U3551) );
  MUX2_X1 U15205 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n13049), .S(n6471), .Z(
        P2_U3550) );
  MUX2_X1 U15206 ( .A(P2_DATAO_REG_18__SCAN_IN), .B(n13050), .S(n6471), .Z(
        P2_U3549) );
  MUX2_X1 U15207 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n13051), .S(n6471), .Z(
        P2_U3548) );
  MUX2_X1 U15208 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n13052), .S(n6471), .Z(
        P2_U3547) );
  MUX2_X1 U15209 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n13053), .S(n6471), .Z(
        P2_U3546) );
  MUX2_X1 U15210 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n13054), .S(n6471), .Z(
        P2_U3545) );
  MUX2_X1 U15211 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n13055), .S(n6471), .Z(
        P2_U3544) );
  MUX2_X1 U15212 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n13056), .S(n6471), .Z(
        P2_U3543) );
  MUX2_X1 U15213 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n13057), .S(n6471), .Z(
        P2_U3542) );
  MUX2_X1 U15214 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n13058), .S(n6471), .Z(
        P2_U3541) );
  MUX2_X1 U15215 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n13059), .S(n6471), .Z(
        P2_U3540) );
  MUX2_X1 U15216 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n13060), .S(n6471), .Z(
        P2_U3539) );
  MUX2_X1 U15217 ( .A(P2_DATAO_REG_7__SCAN_IN), .B(n13061), .S(n6471), .Z(
        P2_U3538) );
  MUX2_X1 U15218 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(n13062), .S(n6471), .Z(
        P2_U3537) );
  MUX2_X1 U15219 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(n13063), .S(n6471), .Z(
        P2_U3536) );
  MUX2_X1 U15220 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n13064), .S(n6471), .Z(
        P2_U3535) );
  MUX2_X1 U15221 ( .A(P2_DATAO_REG_3__SCAN_IN), .B(n13065), .S(n6471), .Z(
        P2_U3534) );
  MUX2_X1 U15222 ( .A(P2_DATAO_REG_2__SCAN_IN), .B(n13066), .S(n6471), .Z(
        P2_U3533) );
  MUX2_X1 U15223 ( .A(P2_DATAO_REG_1__SCAN_IN), .B(n13067), .S(n6471), .Z(
        P2_U3532) );
  OAI22_X1 U15224 ( .A1(n14667), .A2(n13069), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n13068), .ZN(n13070) );
  AOI21_X1 U15225 ( .B1(n14685), .B2(P2_ADDR_REG_1__SCAN_IN), .A(n13070), .ZN(
        n13081) );
  INV_X1 U15226 ( .A(n13071), .ZN(n13074) );
  OAI21_X1 U15227 ( .B1(n14631), .B2(n13075), .A(n13072), .ZN(n13073) );
  NAND3_X1 U15228 ( .A1(n14692), .A2(n13074), .A3(n13073), .ZN(n13080) );
  INV_X1 U15229 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n14798) );
  NOR2_X1 U15230 ( .A1(n13075), .A2(n14798), .ZN(n13077) );
  OAI211_X1 U15231 ( .C1(n13078), .C2(n13077), .A(n14686), .B(n13076), .ZN(
        n13079) );
  NAND3_X1 U15232 ( .A1(n13081), .A2(n13080), .A3(n13079), .ZN(P2_U3215) );
  INV_X1 U15233 ( .A(n13101), .ZN(n13085) );
  NAND3_X1 U15234 ( .A1(n14660), .A2(n13083), .A3(n13082), .ZN(n13084) );
  NAND3_X1 U15235 ( .A1(n13085), .A2(n14692), .A3(n13084), .ZN(n13095) );
  OAI21_X1 U15236 ( .B1(n14667), .B2(n13087), .A(n13086), .ZN(n13088) );
  AOI21_X1 U15237 ( .B1(n14685), .B2(P2_ADDR_REG_6__SCAN_IN), .A(n13088), .ZN(
        n13094) );
  INV_X1 U15238 ( .A(n13111), .ZN(n13092) );
  NAND3_X1 U15239 ( .A1(n14656), .A2(n13090), .A3(n13089), .ZN(n13091) );
  NAND3_X1 U15240 ( .A1(n13092), .A2(n14686), .A3(n13091), .ZN(n13093) );
  NAND3_X1 U15241 ( .A1(n13095), .A2(n13094), .A3(n13093), .ZN(P2_U3220) );
  MUX2_X1 U15242 ( .A(n8875), .B(P2_REG2_REG_7__SCAN_IN), .S(n13105), .Z(
        n13098) );
  INV_X1 U15243 ( .A(n13096), .ZN(n13097) );
  NAND2_X1 U15244 ( .A1(n13098), .A2(n13097), .ZN(n13100) );
  OAI211_X1 U15245 ( .C1(n13101), .C2(n13100), .A(n13099), .B(n14692), .ZN(
        n13114) );
  OAI21_X1 U15246 ( .B1(n14667), .B2(n13103), .A(n13102), .ZN(n13104) );
  AOI21_X1 U15247 ( .B1(n14685), .B2(P2_ADDR_REG_7__SCAN_IN), .A(n13104), .ZN(
        n13113) );
  MUX2_X1 U15248 ( .A(n8866), .B(P2_REG1_REG_7__SCAN_IN), .S(n13105), .Z(
        n13108) );
  INV_X1 U15249 ( .A(n13106), .ZN(n13107) );
  NAND2_X1 U15250 ( .A1(n13108), .A2(n13107), .ZN(n13110) );
  OAI211_X1 U15251 ( .C1(n13111), .C2(n13110), .A(n13109), .B(n14686), .ZN(
        n13112) );
  NAND3_X1 U15252 ( .A1(n13114), .A2(n13113), .A3(n13112), .ZN(P2_U3221) );
  AND3_X1 U15253 ( .A1(n13117), .A2(n13116), .A3(n13115), .ZN(n13118) );
  OAI21_X1 U15254 ( .B1(n13119), .B2(n13118), .A(n14692), .ZN(n13129) );
  NOR2_X1 U15255 ( .A1(n14667), .A2(n13120), .ZN(n13121) );
  AOI211_X1 U15256 ( .C1(n14685), .C2(P2_ADDR_REG_12__SCAN_IN), .A(n13122), 
        .B(n13121), .ZN(n13128) );
  NOR2_X1 U15257 ( .A1(n13124), .A2(n13123), .ZN(n13126) );
  OAI21_X1 U15258 ( .B1(n13126), .B2(n13125), .A(n14686), .ZN(n13127) );
  NAND3_X1 U15259 ( .A1(n13129), .A2(n13128), .A3(n13127), .ZN(P2_U3226) );
  XNOR2_X1 U15260 ( .A(n13149), .B(n13144), .ZN(n13132) );
  NOR2_X1 U15261 ( .A1(P2_REG2_REG_18__SCAN_IN), .A2(n13132), .ZN(n13146) );
  AOI21_X1 U15262 ( .B1(P2_REG2_REG_18__SCAN_IN), .B2(n13132), .A(n13146), 
        .ZN(n13143) );
  OAI21_X1 U15263 ( .B1(n14667), .B2(n13134), .A(n13133), .ZN(n13141) );
  OAI21_X1 U15264 ( .B1(n13137), .B2(n13136), .A(n13135), .ZN(n13148) );
  XOR2_X1 U15265 ( .A(n13149), .B(n13148), .Z(n13138) );
  NAND2_X1 U15266 ( .A1(P2_REG1_REG_18__SCAN_IN), .A2(n13138), .ZN(n13151) );
  OAI21_X1 U15267 ( .B1(P2_REG1_REG_18__SCAN_IN), .B2(n13138), .A(n13151), 
        .ZN(n13139) );
  NOR2_X1 U15268 ( .A1(n13139), .A2(n14639), .ZN(n13140) );
  AOI211_X1 U15269 ( .C1(n14685), .C2(P2_ADDR_REG_18__SCAN_IN), .A(n13141), 
        .B(n13140), .ZN(n13142) );
  OAI21_X1 U15270 ( .B1(n13143), .B2(n14677), .A(n13142), .ZN(P2_U3232) );
  NOR2_X1 U15271 ( .A1(n13149), .A2(n13144), .ZN(n13145) );
  NOR2_X1 U15272 ( .A1(n13146), .A2(n13145), .ZN(n13147) );
  INV_X1 U15273 ( .A(n13156), .ZN(n13154) );
  NAND2_X1 U15274 ( .A1(n13149), .A2(n13148), .ZN(n13150) );
  NAND2_X1 U15275 ( .A1(n13151), .A2(n13150), .ZN(n13152) );
  XOR2_X1 U15276 ( .A(n13152), .B(P2_REG1_REG_19__SCAN_IN), .Z(n13155) );
  OAI21_X1 U15277 ( .B1(n13155), .B2(n14639), .A(n14667), .ZN(n13153) );
  AOI21_X1 U15278 ( .B1(n13154), .B2(n14692), .A(n13153), .ZN(n13158) );
  MUX2_X1 U15279 ( .A(n13158), .B(n13157), .S(n13253), .Z(n13160) );
  OAI211_X1 U15280 ( .C1(n7543), .C2(n14671), .A(n13160), .B(n13159), .ZN(
        P2_U3233) );
  NAND2_X1 U15281 ( .A1(n13162), .A2(n14714), .ZN(n13321) );
  NAND2_X1 U15282 ( .A1(n13164), .A2(n13163), .ZN(n13322) );
  NOR2_X1 U15283 ( .A1(n14731), .A2(n13322), .ZN(n13170) );
  NOR2_X1 U15284 ( .A1(n6858), .A2(n14721), .ZN(n13165) );
  AOI211_X1 U15285 ( .C1(n14708), .C2(P2_REG2_REG_31__SCAN_IN), .A(n13170), 
        .B(n13165), .ZN(n13166) );
  OAI21_X1 U15286 ( .B1(n13321), .B2(n13282), .A(n13166), .ZN(P2_U3234) );
  OAI211_X1 U15287 ( .C1(n13324), .C2(n13168), .A(n13167), .B(n14714), .ZN(
        n13323) );
  NOR2_X1 U15288 ( .A1(n13324), .A2(n14721), .ZN(n13169) );
  AOI211_X1 U15289 ( .C1(n14708), .C2(P2_REG2_REG_30__SCAN_IN), .A(n13170), 
        .B(n13169), .ZN(n13171) );
  OAI21_X1 U15290 ( .B1(n13282), .B2(n13323), .A(n13171), .ZN(P2_U3235) );
  AOI22_X1 U15291 ( .A1(n13331), .A2(n14341), .B1(n14708), .B2(
        P2_REG2_REG_28__SCAN_IN), .ZN(n13185) );
  INV_X1 U15292 ( .A(n13172), .ZN(n13174) );
  AOI21_X1 U15293 ( .B1(n13174), .B2(n7215), .A(n14352), .ZN(n13177) );
  AOI21_X1 U15294 ( .B1(n13177), .B2(n13176), .A(n13175), .ZN(n13334) );
  INV_X1 U15295 ( .A(n13190), .ZN(n13180) );
  INV_X1 U15296 ( .A(n13178), .ZN(n13179) );
  AOI21_X1 U15297 ( .B1(n13331), .B2(n13180), .A(n13179), .ZN(n13332) );
  AOI22_X1 U15298 ( .A1(n13332), .A2(n9335), .B1(n13181), .B2(n14719), .ZN(
        n13182) );
  AOI21_X1 U15299 ( .B1(n13334), .B2(n13182), .A(n14708), .ZN(n13183) );
  INV_X1 U15300 ( .A(n13183), .ZN(n13184) );
  OAI211_X1 U15301 ( .C1(n13335), .C2(n13304), .A(n13185), .B(n13184), .ZN(
        P2_U3237) );
  XNOR2_X1 U15302 ( .A(n13187), .B(n13186), .ZN(n13342) );
  XNOR2_X1 U15303 ( .A(n13188), .B(n13189), .ZN(n13336) );
  NAND2_X1 U15304 ( .A1(n13336), .A2(n14727), .ZN(n13197) );
  AOI211_X1 U15305 ( .C1(n13339), .C2(n13202), .A(n9329), .B(n13190), .ZN(
        n13337) );
  INV_X1 U15306 ( .A(n13339), .ZN(n13194) );
  AOI22_X1 U15307 ( .A1(n13316), .A2(n13338), .B1(n13191), .B2(n14719), .ZN(
        n13193) );
  NAND2_X1 U15308 ( .A1(n14731), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n13192) );
  OAI211_X1 U15309 ( .C1(n13194), .C2(n14721), .A(n13193), .B(n13192), .ZN(
        n13195) );
  AOI21_X1 U15310 ( .B1(n13337), .B2(n14725), .A(n13195), .ZN(n13196) );
  OAI211_X1 U15311 ( .C1(n13342), .C2(n13198), .A(n13197), .B(n13196), .ZN(
        P2_U3238) );
  XOR2_X1 U15312 ( .A(n13199), .B(n13200), .Z(n13349) );
  XNOR2_X1 U15313 ( .A(n13201), .B(n13200), .ZN(n13347) );
  OAI211_X1 U15314 ( .C1(n13345), .C2(n13203), .A(n14714), .B(n13202), .ZN(
        n13344) );
  INV_X1 U15315 ( .A(n13204), .ZN(n13205) );
  OAI22_X1 U15316 ( .A1(n14708), .A2(n13343), .B1(n13205), .B2(n14706), .ZN(
        n13207) );
  NOR2_X1 U15317 ( .A1(n13345), .A2(n14721), .ZN(n13206) );
  AOI211_X1 U15318 ( .C1(n14731), .C2(P2_REG2_REG_26__SCAN_IN), .A(n13207), 
        .B(n13206), .ZN(n13208) );
  OAI21_X1 U15319 ( .B1(n13282), .B2(n13344), .A(n13208), .ZN(n13209) );
  AOI21_X1 U15320 ( .B1(n13347), .B2(n13284), .A(n13209), .ZN(n13210) );
  OAI21_X1 U15321 ( .B1(n13349), .B2(n13304), .A(n13210), .ZN(P2_U3239) );
  XNOR2_X1 U15322 ( .A(n13211), .B(n13215), .ZN(n13353) );
  INV_X1 U15323 ( .A(n13212), .ZN(n13213) );
  AOI21_X1 U15324 ( .B1(n13215), .B2(n13214), .A(n13213), .ZN(n13356) );
  INV_X1 U15325 ( .A(n13351), .ZN(n13219) );
  NAND2_X1 U15326 ( .A1(n14708), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n13218) );
  NAND2_X1 U15327 ( .A1(n14719), .A2(n13216), .ZN(n13217) );
  OAI211_X1 U15328 ( .C1(n14731), .C2(n13219), .A(n13218), .B(n13217), .ZN(
        n13220) );
  AOI21_X1 U15329 ( .B1(n13352), .B2(n14341), .A(n13220), .ZN(n13224) );
  AOI21_X1 U15330 ( .B1(n13238), .B2(n13352), .A(n9329), .ZN(n13222) );
  AND2_X1 U15331 ( .A1(n13222), .A2(n13221), .ZN(n13350) );
  NAND2_X1 U15332 ( .A1(n13350), .A2(n14725), .ZN(n13223) );
  OAI211_X1 U15333 ( .C1(n13356), .C2(n13304), .A(n13224), .B(n13223), .ZN(
        n13225) );
  AOI21_X1 U15334 ( .B1(n13284), .B2(n13353), .A(n13225), .ZN(n13226) );
  INV_X1 U15335 ( .A(n13226), .ZN(P2_U3240) );
  XNOR2_X1 U15336 ( .A(n13227), .B(n13231), .ZN(n13229) );
  AOI21_X1 U15337 ( .B1(n13229), .B2(n14740), .A(n13228), .ZN(n13360) );
  OAI21_X1 U15338 ( .B1(n13232), .B2(n13231), .A(n13230), .ZN(n13361) );
  NAND2_X1 U15339 ( .A1(n14708), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n13233) );
  OAI21_X1 U15340 ( .B1(n14706), .B2(n13234), .A(n13233), .ZN(n13235) );
  AOI21_X1 U15341 ( .B1(n13358), .B2(n14341), .A(n13235), .ZN(n13240) );
  OR2_X1 U15342 ( .A1(n13236), .A2(n6519), .ZN(n13237) );
  AND3_X1 U15343 ( .A1(n13238), .A2(n13237), .A3(n14714), .ZN(n13357) );
  NAND2_X1 U15344 ( .A1(n13357), .A2(n14725), .ZN(n13239) );
  OAI211_X1 U15345 ( .C1(n13361), .C2(n13304), .A(n13240), .B(n13239), .ZN(
        n13241) );
  INV_X1 U15346 ( .A(n13241), .ZN(n13242) );
  OAI21_X1 U15347 ( .B1(n14731), .B2(n13360), .A(n13242), .ZN(P2_U3241) );
  AOI21_X1 U15348 ( .B1(n13245), .B2(n13244), .A(n13243), .ZN(n13366) );
  AOI22_X1 U15349 ( .A1(n13363), .A2(n14341), .B1(P2_REG2_REG_23__SCAN_IN), 
        .B2(n14731), .ZN(n13258) );
  AOI21_X1 U15350 ( .B1(n13247), .B2(n13246), .A(n6549), .ZN(n13248) );
  NOR2_X1 U15351 ( .A1(n13248), .A2(n14352), .ZN(n13250) );
  NOR2_X1 U15352 ( .A1(n13250), .A2(n13249), .ZN(n13365) );
  NAND2_X1 U15353 ( .A1(n13363), .A2(n13263), .ZN(n13251) );
  NAND2_X1 U15354 ( .A1(n13251), .A2(n14714), .ZN(n13252) );
  NOR2_X1 U15355 ( .A1(n6519), .A2(n13252), .ZN(n13362) );
  NAND2_X1 U15356 ( .A1(n13362), .A2(n13253), .ZN(n13254) );
  OAI211_X1 U15357 ( .C1(n14706), .C2(n13255), .A(n13365), .B(n13254), .ZN(
        n13256) );
  NAND2_X1 U15358 ( .A1(n13256), .A2(n13316), .ZN(n13257) );
  OAI211_X1 U15359 ( .C1(n13366), .C2(n13304), .A(n13258), .B(n13257), .ZN(
        P2_U3242) );
  XNOR2_X1 U15360 ( .A(n13259), .B(n13260), .ZN(n13262) );
  AOI21_X1 U15361 ( .B1(n13262), .B2(n14740), .A(n13261), .ZN(n13370) );
  INV_X1 U15362 ( .A(n13263), .ZN(n13264) );
  AOI211_X1 U15363 ( .C1(n13368), .C2(n13276), .A(n9329), .B(n13264), .ZN(
        n13367) );
  AOI22_X1 U15364 ( .A1(n14731), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n13265), 
        .B2(n14719), .ZN(n13266) );
  OAI21_X1 U15365 ( .B1(n6939), .B2(n14721), .A(n13266), .ZN(n13271) );
  OAI21_X1 U15366 ( .B1(n13269), .B2(n13268), .A(n13267), .ZN(n13371) );
  NOR2_X1 U15367 ( .A1(n13371), .A2(n13304), .ZN(n13270) );
  AOI211_X1 U15368 ( .C1(n13367), .C2(n14725), .A(n13271), .B(n13270), .ZN(
        n13272) );
  OAI21_X1 U15369 ( .B1(n14708), .B2(n13370), .A(n13272), .ZN(P2_U3243) );
  XNOR2_X1 U15370 ( .A(n13273), .B(n13274), .ZN(n13378) );
  XNOR2_X1 U15371 ( .A(n13275), .B(n13274), .ZN(n13376) );
  OAI211_X1 U15372 ( .C1(n13374), .C2(n13299), .A(n14714), .B(n13276), .ZN(
        n13373) );
  INV_X1 U15373 ( .A(n13277), .ZN(n13372) );
  OAI22_X1 U15374 ( .A1(n13372), .A2(n14708), .B1(n13278), .B2(n14706), .ZN(
        n13280) );
  NOR2_X1 U15375 ( .A1(n13374), .A2(n14721), .ZN(n13279) );
  AOI211_X1 U15376 ( .C1(n14708), .C2(P2_REG2_REG_21__SCAN_IN), .A(n13280), 
        .B(n13279), .ZN(n13281) );
  OAI21_X1 U15377 ( .B1(n13282), .B2(n13373), .A(n13281), .ZN(n13283) );
  AOI21_X1 U15378 ( .B1(n13284), .B2(n13376), .A(n13283), .ZN(n13285) );
  OAI21_X1 U15379 ( .B1(n13378), .B2(n13304), .A(n13285), .ZN(P2_U3244) );
  XNOR2_X1 U15380 ( .A(n13286), .B(n13288), .ZN(n13383) );
  OAI21_X1 U15381 ( .B1(n13289), .B2(n13288), .A(n13287), .ZN(n13292) );
  INV_X1 U15382 ( .A(n13290), .ZN(n13291) );
  AOI21_X1 U15383 ( .B1(n13292), .B2(n14740), .A(n13291), .ZN(n13382) );
  NAND2_X1 U15384 ( .A1(n14708), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n13293) );
  OAI21_X1 U15385 ( .B1(n14706), .B2(n13294), .A(n13293), .ZN(n13295) );
  AOI21_X1 U15386 ( .B1(n13380), .B2(n14341), .A(n13295), .ZN(n13301) );
  NAND2_X1 U15387 ( .A1(n13380), .A2(n13296), .ZN(n13297) );
  NAND2_X1 U15388 ( .A1(n13297), .A2(n14714), .ZN(n13298) );
  NOR2_X1 U15389 ( .A1(n13299), .A2(n13298), .ZN(n13379) );
  NAND2_X1 U15390 ( .A1(n13379), .A2(n14725), .ZN(n13300) );
  OAI211_X1 U15391 ( .C1(n13382), .C2(n14731), .A(n13301), .B(n13300), .ZN(
        n13302) );
  INV_X1 U15392 ( .A(n13302), .ZN(n13303) );
  OAI21_X1 U15393 ( .B1(n13383), .B2(n13304), .A(n13303), .ZN(P2_U3245) );
  OAI21_X1 U15394 ( .B1(n13306), .B2(n13307), .A(n13305), .ZN(n13312) );
  INV_X1 U15395 ( .A(n13312), .ZN(n13394) );
  XNOR2_X1 U15396 ( .A(n13308), .B(n13307), .ZN(n13309) );
  NOR2_X1 U15397 ( .A1(n13309), .A2(n14352), .ZN(n13311) );
  AOI211_X1 U15398 ( .C1(n13312), .C2(n14741), .A(n13311), .B(n13310), .ZN(
        n13393) );
  AOI21_X1 U15399 ( .B1(n13390), .B2(n13313), .A(n6860), .ZN(n13391) );
  NAND2_X1 U15400 ( .A1(n13391), .A2(n9335), .ZN(n13314) );
  OAI211_X1 U15401 ( .C1(n14706), .C2(n13315), .A(n13393), .B(n13314), .ZN(
        n13317) );
  NAND2_X1 U15402 ( .A1(n13317), .A2(n13316), .ZN(n13319) );
  AOI22_X1 U15403 ( .A1(n13390), .A2(n14341), .B1(n14708), .B2(
        P2_REG2_REG_18__SCAN_IN), .ZN(n13318) );
  OAI211_X1 U15404 ( .C1(n13394), .C2(n13320), .A(n13319), .B(n13318), .ZN(
        P2_U3247) );
  OAI211_X1 U15405 ( .C1(n6858), .C2(n14774), .A(n13321), .B(n13322), .ZN(
        n13408) );
  MUX2_X1 U15406 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n13408), .S(n6470), .Z(
        P2_U3530) );
  OAI211_X1 U15407 ( .C1(n13324), .C2(n14774), .A(n13323), .B(n13322), .ZN(
        n13409) );
  MUX2_X1 U15408 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n13409), .S(n6470), .Z(
        P2_U3529) );
  NAND2_X1 U15409 ( .A1(n13325), .A2(n14768), .ZN(n13330) );
  AOI21_X1 U15410 ( .B1(n13327), .B2(n14788), .A(n13326), .ZN(n13329) );
  MUX2_X1 U15411 ( .A(P2_REG1_REG_29__SCAN_IN), .B(n13410), .S(n6470), .Z(
        P2_U3528) );
  AOI22_X1 U15412 ( .A1(n13332), .A2(n14714), .B1(n13331), .B2(n14788), .ZN(
        n13333) );
  MUX2_X1 U15413 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n13411), .S(n6470), .Z(
        P2_U3527) );
  NAND2_X1 U15414 ( .A1(n13336), .A2(n14768), .ZN(n13341) );
  AOI211_X1 U15415 ( .C1(n13339), .C2(n14788), .A(n13338), .B(n13337), .ZN(
        n13340) );
  OAI211_X1 U15416 ( .C1(n14352), .C2(n13342), .A(n13341), .B(n13340), .ZN(
        n13412) );
  MUX2_X1 U15417 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n13412), .S(n6470), .Z(
        P2_U3526) );
  OAI211_X1 U15418 ( .C1(n13345), .C2(n14774), .A(n13344), .B(n13343), .ZN(
        n13346) );
  AOI21_X1 U15419 ( .B1(n13347), .B2(n14740), .A(n13346), .ZN(n13348) );
  OAI21_X1 U15420 ( .B1(n13349), .B2(n13406), .A(n13348), .ZN(n13413) );
  MUX2_X1 U15421 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n13413), .S(n6470), .Z(
        P2_U3525) );
  AOI211_X1 U15422 ( .C1(n13352), .C2(n14788), .A(n13351), .B(n13350), .ZN(
        n13355) );
  NAND2_X1 U15423 ( .A1(n13353), .A2(n14740), .ZN(n13354) );
  OAI211_X1 U15424 ( .C1(n13356), .C2(n13406), .A(n13355), .B(n13354), .ZN(
        n13414) );
  MUX2_X1 U15425 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n13414), .S(n6470), .Z(
        P2_U3524) );
  AOI21_X1 U15426 ( .B1(n13358), .B2(n14788), .A(n13357), .ZN(n13359) );
  OAI211_X1 U15427 ( .C1(n13361), .C2(n13406), .A(n13360), .B(n13359), .ZN(
        n13415) );
  MUX2_X1 U15428 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n13415), .S(n6470), .Z(
        P2_U3523) );
  AOI21_X1 U15429 ( .B1(n13363), .B2(n14788), .A(n13362), .ZN(n13364) );
  OAI211_X1 U15430 ( .C1(n13366), .C2(n13406), .A(n13365), .B(n13364), .ZN(
        n13416) );
  MUX2_X1 U15431 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n13416), .S(n6470), .Z(
        P2_U3522) );
  AOI21_X1 U15432 ( .B1(n13368), .B2(n14788), .A(n13367), .ZN(n13369) );
  OAI211_X1 U15433 ( .C1(n13371), .C2(n13406), .A(n13370), .B(n13369), .ZN(
        n13417) );
  MUX2_X1 U15434 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n13417), .S(n6470), .Z(
        P2_U3521) );
  OAI211_X1 U15435 ( .C1(n13374), .C2(n14774), .A(n13373), .B(n13372), .ZN(
        n13375) );
  AOI21_X1 U15436 ( .B1(n13376), .B2(n14740), .A(n13375), .ZN(n13377) );
  OAI21_X1 U15437 ( .B1(n13378), .B2(n13406), .A(n13377), .ZN(n13418) );
  MUX2_X1 U15438 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n13418), .S(n6470), .Z(
        P2_U3520) );
  AOI21_X1 U15439 ( .B1(n13380), .B2(n14788), .A(n13379), .ZN(n13381) );
  OAI211_X1 U15440 ( .C1(n13383), .C2(n13406), .A(n13382), .B(n13381), .ZN(
        n13419) );
  MUX2_X1 U15441 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n13419), .S(n6470), .Z(
        P2_U3519) );
  OAI211_X1 U15442 ( .C1(n6859), .C2(n14774), .A(n13385), .B(n13384), .ZN(
        n13386) );
  AOI21_X1 U15443 ( .B1(n13387), .B2(n14740), .A(n13386), .ZN(n13388) );
  OAI21_X1 U15444 ( .B1(n13389), .B2(n13406), .A(n13388), .ZN(n13420) );
  MUX2_X1 U15445 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n13420), .S(n6470), .Z(
        P2_U3518) );
  AOI22_X1 U15446 ( .A1(n13391), .A2(n14714), .B1(n13390), .B2(n14788), .ZN(
        n13392) );
  OAI211_X1 U15447 ( .C1(n13394), .C2(n14793), .A(n13393), .B(n13392), .ZN(
        n13421) );
  MUX2_X1 U15448 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n13421), .S(n6470), .Z(
        P2_U3517) );
  OAI211_X1 U15449 ( .C1(n13397), .C2(n14774), .A(n13396), .B(n13395), .ZN(
        n13398) );
  AOI21_X1 U15450 ( .B1(n13399), .B2(n14740), .A(n13398), .ZN(n13400) );
  OAI21_X1 U15451 ( .B1(n13401), .B2(n13406), .A(n13400), .ZN(n13422) );
  MUX2_X1 U15452 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n13422), .S(n6470), .Z(
        P2_U3516) );
  AOI211_X1 U15453 ( .C1(n13404), .C2(n14788), .A(n13403), .B(n13402), .ZN(
        n13405) );
  OAI21_X1 U15454 ( .B1(n13407), .B2(n13406), .A(n13405), .ZN(n13423) );
  MUX2_X1 U15455 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n13423), .S(n6470), .Z(
        P2_U3515) );
  MUX2_X1 U15456 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n13408), .S(n14797), .Z(
        P2_U3498) );
  MUX2_X1 U15457 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n13409), .S(n14797), .Z(
        P2_U3497) );
  MUX2_X1 U15458 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n13410), .S(n14797), .Z(
        P2_U3496) );
  MUX2_X1 U15459 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n13412), .S(n14797), .Z(
        P2_U3494) );
  MUX2_X1 U15460 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n13413), .S(n14797), .Z(
        P2_U3493) );
  MUX2_X1 U15461 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n13414), .S(n14797), .Z(
        P2_U3492) );
  MUX2_X1 U15462 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n13415), .S(n14797), .Z(
        P2_U3491) );
  MUX2_X1 U15463 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n13416), .S(n14797), .Z(
        P2_U3490) );
  MUX2_X1 U15464 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n13417), .S(n14797), .Z(
        P2_U3489) );
  MUX2_X1 U15465 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n13418), .S(n14797), .Z(
        P2_U3488) );
  MUX2_X1 U15466 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n13419), .S(n14797), .Z(
        P2_U3487) );
  MUX2_X1 U15467 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n13420), .S(n14797), .Z(
        P2_U3486) );
  MUX2_X1 U15468 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n13421), .S(n14797), .Z(
        P2_U3484) );
  MUX2_X1 U15469 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n13422), .S(n14797), .Z(
        P2_U3481) );
  MUX2_X1 U15470 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n13423), .S(n14797), .Z(
        P2_U3478) );
  INV_X1 U15471 ( .A(n12944), .ZN(n14116) );
  NOR4_X1 U15472 ( .A1(n13424), .A2(P2_IR_REG_30__SCAN_IN), .A3(n8671), .A4(
        P2_U3088), .ZN(n13425) );
  AOI21_X1 U15473 ( .B1(n13428), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n13425), 
        .ZN(n13426) );
  OAI21_X1 U15474 ( .B1(n14116), .B2(n13438), .A(n13426), .ZN(P2_U3296) );
  AOI21_X1 U15475 ( .B1(n13428), .B2(P1_DATAO_REG_28__SCAN_IN), .A(n13427), 
        .ZN(n13429) );
  OAI21_X1 U15476 ( .B1(n13430), .B2(n13438), .A(n13429), .ZN(P2_U3299) );
  INV_X1 U15477 ( .A(n13431), .ZN(n14122) );
  OAI222_X1 U15478 ( .A1(n13440), .A2(n13433), .B1(n13438), .B2(n14122), .C1(
        n13432), .C2(P2_U3088), .ZN(P2_U3300) );
  INV_X1 U15479 ( .A(n13434), .ZN(n14126) );
  OAI222_X1 U15480 ( .A1(n13435), .A2(P2_U3088), .B1(n13438), .B2(n14126), 
        .C1(n6834), .C2(n13440), .ZN(P2_U3301) );
  INV_X1 U15481 ( .A(n13436), .ZN(n14129) );
  OAI222_X1 U15482 ( .A1(n13440), .A2(n13439), .B1(n13438), .B2(n14129), .C1(
        n13437), .C2(P2_U3088), .ZN(P2_U3302) );
  MUX2_X1 U15483 ( .A(n13441), .B(P2_IR_REG_0__SCAN_IN), .S(
        P2_STATE_REG_SCAN_IN), .Z(P2_U3327) );
  NAND2_X1 U15484 ( .A1(n14038), .A2(n13481), .ZN(n13444) );
  NAND2_X1 U15485 ( .A1(n13847), .A2(n13442), .ZN(n13443) );
  NAND2_X1 U15486 ( .A1(n13444), .A2(n13443), .ZN(n13445) );
  XNOR2_X1 U15487 ( .A(n13445), .B(n13536), .ZN(n13449) );
  NAND2_X1 U15488 ( .A1(n14038), .A2(n13442), .ZN(n13447) );
  NAND2_X1 U15489 ( .A1(n13485), .A2(n13847), .ZN(n13446) );
  NAND2_X1 U15490 ( .A1(n13447), .A2(n13446), .ZN(n13448) );
  NOR2_X1 U15491 ( .A1(n13449), .A2(n13448), .ZN(n13533) );
  AOI21_X1 U15492 ( .B1(n13449), .B2(n13448), .A(n13533), .ZN(n13493) );
  NAND2_X1 U15493 ( .A1(n14062), .A2(n13481), .ZN(n13453) );
  NAND2_X1 U15494 ( .A1(n13888), .A2(n13442), .ZN(n13452) );
  NAND2_X1 U15495 ( .A1(n13453), .A2(n13452), .ZN(n13454) );
  XNOR2_X1 U15496 ( .A(n13454), .B(n13536), .ZN(n13458) );
  NAND2_X1 U15497 ( .A1(n14062), .A2(n13442), .ZN(n13456) );
  NAND2_X1 U15498 ( .A1(n13888), .A2(n13485), .ZN(n13455) );
  NAND2_X1 U15499 ( .A1(n13456), .A2(n13455), .ZN(n13457) );
  NOR2_X1 U15500 ( .A1(n13458), .A2(n13457), .ZN(n13592) );
  AOI21_X1 U15501 ( .B1(n13458), .B2(n13457), .A(n13592), .ZN(n13510) );
  NAND2_X1 U15502 ( .A1(n13898), .A2(n13481), .ZN(n13460) );
  NAND2_X1 U15503 ( .A1(n13865), .A2(n13442), .ZN(n13459) );
  NAND2_X1 U15504 ( .A1(n13460), .A2(n13459), .ZN(n13461) );
  XNOR2_X1 U15505 ( .A(n13461), .B(n13471), .ZN(n13464) );
  NOR2_X1 U15506 ( .A1(n13462), .A2(n13538), .ZN(n13463) );
  AOI21_X1 U15507 ( .B1(n13898), .B2(n13442), .A(n13463), .ZN(n13465) );
  NAND2_X1 U15508 ( .A1(n13464), .A2(n13465), .ZN(n13563) );
  INV_X1 U15509 ( .A(n13464), .ZN(n13467) );
  INV_X1 U15510 ( .A(n13465), .ZN(n13466) );
  NAND2_X1 U15511 ( .A1(n13467), .A2(n13466), .ZN(n13468) );
  NAND2_X1 U15512 ( .A1(n14049), .A2(n13481), .ZN(n13470) );
  NAND2_X1 U15513 ( .A1(n13887), .A2(n9619), .ZN(n13469) );
  NAND2_X1 U15514 ( .A1(n13470), .A2(n13469), .ZN(n13472) );
  XNOR2_X1 U15515 ( .A(n13472), .B(n13471), .ZN(n13474) );
  NOR2_X1 U15516 ( .A1(n13630), .A2(n13538), .ZN(n13473) );
  AOI21_X1 U15517 ( .B1(n14049), .B2(n13442), .A(n13473), .ZN(n13475) );
  NAND2_X1 U15518 ( .A1(n13474), .A2(n13475), .ZN(n13480) );
  INV_X1 U15519 ( .A(n13474), .ZN(n13477) );
  INV_X1 U15520 ( .A(n13475), .ZN(n13476) );
  NAND2_X1 U15521 ( .A1(n13477), .A2(n13476), .ZN(n13478) );
  NAND2_X1 U15522 ( .A1(n13479), .A2(n13561), .ZN(n13565) );
  NAND2_X1 U15523 ( .A1(n14043), .A2(n13481), .ZN(n13483) );
  NAND2_X1 U15524 ( .A1(n13866), .A2(n9619), .ZN(n13482) );
  NAND2_X1 U15525 ( .A1(n13483), .A2(n13482), .ZN(n13484) );
  XNOR2_X1 U15526 ( .A(n13484), .B(n13536), .ZN(n13489) );
  NAND2_X1 U15527 ( .A1(n14043), .A2(n9619), .ZN(n13487) );
  NAND2_X1 U15528 ( .A1(n13485), .A2(n13866), .ZN(n13486) );
  NAND2_X1 U15529 ( .A1(n13487), .A2(n13486), .ZN(n13488) );
  NOR2_X1 U15530 ( .A1(n13489), .A2(n13488), .ZN(n13490) );
  AOI21_X1 U15531 ( .B1(n13489), .B2(n13488), .A(n13490), .ZN(n13625) );
  INV_X1 U15532 ( .A(n13490), .ZN(n13491) );
  OAI21_X1 U15533 ( .B1(n13493), .B2(n13492), .A(n13534), .ZN(n13494) );
  INV_X1 U15534 ( .A(n13836), .ZN(n13497) );
  AOI22_X1 U15535 ( .A1(n13639), .A2(n13654), .B1(P1_REG3_REG_27__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13495) );
  OAI21_X1 U15536 ( .B1(n13830), .B2(n13629), .A(n13495), .ZN(n13496) );
  AOI21_X1 U15537 ( .B1(n13497), .B2(n13632), .A(n13496), .ZN(n13498) );
  OAI21_X1 U15538 ( .B1(n13501), .B2(n13500), .A(n13499), .ZN(n13502) );
  NAND2_X1 U15539 ( .A1(n13502), .A2(n13626), .ZN(n13508) );
  NOR2_X1 U15540 ( .A1(n13644), .A2(n14386), .ZN(n13506) );
  OAI21_X1 U15541 ( .B1(n13617), .B2(n13504), .A(n13503), .ZN(n13505) );
  AOI211_X1 U15542 ( .C1(n13620), .C2(n14394), .A(n13506), .B(n13505), .ZN(
        n13507) );
  OAI211_X1 U15543 ( .C1(n14426), .C2(n13636), .A(n13508), .B(n13507), .ZN(
        P1_U3215) );
  INV_X1 U15544 ( .A(n14062), .ZN(n13908) );
  OAI21_X1 U15545 ( .B1(n13510), .B2(n13509), .A(n13590), .ZN(n13511) );
  NAND2_X1 U15546 ( .A1(n13511), .A2(n13626), .ZN(n13516) );
  AOI22_X1 U15547 ( .A1(n13936), .A2(n14527), .B1(n14524), .B2(n13865), .ZN(
        n13910) );
  INV_X1 U15548 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n13512) );
  OAI22_X1 U15549 ( .A1(n13910), .A2(n13513), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n13512), .ZN(n13514) );
  AOI21_X1 U15550 ( .B1(n13906), .B2(n13632), .A(n13514), .ZN(n13515) );
  OAI211_X1 U15551 ( .C1(n13908), .C2(n13636), .A(n13516), .B(n13515), .ZN(
        P1_U3216) );
  OAI211_X1 U15552 ( .C1(n13518), .C2(n13517), .A(n9835), .B(n13626), .ZN(
        n13523) );
  AOI22_X1 U15553 ( .A1(n13647), .A2(n13519), .B1(n13620), .B2(n14525), .ZN(
        n13522) );
  NOR2_X1 U15554 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9612), .ZN(n13698) );
  NOR2_X1 U15555 ( .A1(n13644), .A2(P1_REG3_REG_3__SCAN_IN), .ZN(n13520) );
  AOI211_X1 U15556 ( .C1(n13639), .C2(n13665), .A(n13698), .B(n13520), .ZN(
        n13521) );
  NAND3_X1 U15557 ( .A1(n13523), .A2(n13522), .A3(n13521), .ZN(P1_U3218) );
  AND2_X1 U15558 ( .A1(n13611), .A2(n13524), .ZN(n13527) );
  OAI211_X1 U15559 ( .C1(n13527), .C2(n13526), .A(n13626), .B(n13525), .ZN(
        n13532) );
  NOR2_X1 U15560 ( .A1(n13644), .A2(n13966), .ZN(n13529) );
  NAND2_X1 U15561 ( .A1(P1_U3086), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n13809)
         );
  OAI21_X1 U15562 ( .B1(n13617), .B2(n13964), .A(n13809), .ZN(n13528) );
  AOI211_X1 U15563 ( .C1(n13620), .C2(n13530), .A(n13529), .B(n13528), .ZN(
        n13531) );
  OAI211_X1 U15564 ( .C1(n14083), .C2(n13636), .A(n13532), .B(n13531), .ZN(
        P1_U3219) );
  OAI22_X1 U15565 ( .A1(n13540), .A2(n13535), .B1(n13829), .B2(n13539), .ZN(
        n13537) );
  XNOR2_X1 U15566 ( .A(n13537), .B(n13536), .ZN(n13542) );
  OAI22_X1 U15567 ( .A1(n13540), .A2(n13539), .B1(n13829), .B2(n13538), .ZN(
        n13541) );
  XNOR2_X1 U15568 ( .A(n13542), .B(n13541), .ZN(n13543) );
  AOI22_X1 U15569 ( .A1(n13620), .A2(n13847), .B1(P1_REG3_REG_28__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13545) );
  NAND2_X1 U15570 ( .A1(n13639), .A2(n13653), .ZN(n13544) );
  OAI211_X1 U15571 ( .C1(n13644), .C2(n13546), .A(n13545), .B(n13544), .ZN(
        n13547) );
  AOI21_X1 U15572 ( .B1(n14032), .B2(n13647), .A(n13547), .ZN(n13548) );
  OAI21_X1 U15573 ( .B1(n13549), .B2(n13650), .A(n13548), .ZN(P1_U3220) );
  AOI21_X1 U15574 ( .B1(n13552), .B2(n13551), .A(n13550), .ZN(n13557) );
  AOI22_X1 U15575 ( .A1(n13936), .A2(n13639), .B1(P1_REG3_REG_21__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13554) );
  NAND2_X1 U15576 ( .A1(n13620), .A2(n13935), .ZN(n13553) );
  OAI211_X1 U15577 ( .C1(n13644), .C2(n13930), .A(n13554), .B(n13553), .ZN(
        n13555) );
  AOI21_X1 U15578 ( .B1(n14072), .B2(n13647), .A(n13555), .ZN(n13556) );
  OAI21_X1 U15579 ( .B1(n13557), .B2(n13650), .A(n13556), .ZN(P1_U3223) );
  AOI22_X1 U15580 ( .A1(n13639), .A2(n13866), .B1(P1_REG3_REG_25__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13559) );
  NAND2_X1 U15581 ( .A1(n13620), .A2(n13865), .ZN(n13558) );
  OAI211_X1 U15582 ( .C1(n13644), .C2(n13869), .A(n13559), .B(n13558), .ZN(
        n13567) );
  INV_X1 U15583 ( .A(n13561), .ZN(n13562) );
  NAND3_X1 U15584 ( .A1(n13560), .A2(n13563), .A3(n13562), .ZN(n13564) );
  AOI21_X1 U15585 ( .B1(n13565), .B2(n13564), .A(n13650), .ZN(n13566) );
  AOI211_X1 U15586 ( .C1(n14049), .C2(n13647), .A(n13567), .B(n13566), .ZN(
        n13568) );
  INV_X1 U15587 ( .A(n13568), .ZN(P1_U3225) );
  AOI21_X1 U15588 ( .B1(n13571), .B2(n13570), .A(n13569), .ZN(n13579) );
  OAI21_X1 U15589 ( .B1(n13617), .B2(n13573), .A(n13572), .ZN(n13574) );
  AOI21_X1 U15590 ( .B1(n13620), .B2(n14385), .A(n13574), .ZN(n13575) );
  OAI21_X1 U15591 ( .B1(n13576), .B2(n13644), .A(n13575), .ZN(n13577) );
  AOI21_X1 U15592 ( .B1(n14409), .B2(n13647), .A(n13577), .ZN(n13578) );
  OAI21_X1 U15593 ( .B1(n13579), .B2(n13650), .A(n13578), .ZN(P1_U3226) );
  INV_X1 U15594 ( .A(n14090), .ZN(n13999) );
  INV_X1 U15595 ( .A(n13580), .ZN(n13584) );
  NOR3_X1 U15596 ( .A1(n13569), .A2(n13582), .A3(n13581), .ZN(n13583) );
  OAI21_X1 U15597 ( .B1(n13584), .B2(n13583), .A(n13626), .ZN(n13589) );
  NOR2_X1 U15598 ( .A1(n13644), .A2(n13995), .ZN(n13587) );
  OAI21_X1 U15599 ( .B1(n13617), .B2(n14009), .A(n13585), .ZN(n13586) );
  AOI211_X1 U15600 ( .C1(n13620), .C2(n13655), .A(n13587), .B(n13586), .ZN(
        n13588) );
  OAI211_X1 U15601 ( .C1(n13999), .C2(n13636), .A(n13589), .B(n13588), .ZN(
        P1_U3228) );
  INV_X1 U15602 ( .A(n13590), .ZN(n13593) );
  NOR3_X1 U15603 ( .A1(n13593), .A2(n13592), .A3(n13591), .ZN(n13595) );
  INV_X1 U15604 ( .A(n13560), .ZN(n13594) );
  OAI21_X1 U15605 ( .B1(n13595), .B2(n13594), .A(n13626), .ZN(n13600) );
  INV_X1 U15606 ( .A(n13895), .ZN(n13598) );
  AOI22_X1 U15607 ( .A1(n13639), .A2(n13887), .B1(P1_REG3_REG_24__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13596) );
  OAI21_X1 U15608 ( .B1(n13918), .B2(n13629), .A(n13596), .ZN(n13597) );
  AOI21_X1 U15609 ( .B1(n13598), .B2(n13632), .A(n13597), .ZN(n13599) );
  OAI211_X1 U15610 ( .C1(n14056), .C2(n13636), .A(n13600), .B(n13599), .ZN(
        P1_U3229) );
  XNOR2_X1 U15611 ( .A(n13602), .B(n13601), .ZN(n13610) );
  INV_X1 U15612 ( .A(n13953), .ZN(n13603) );
  OR2_X1 U15613 ( .A1(n13644), .A2(n13603), .ZN(n13607) );
  NAND2_X1 U15614 ( .A1(n13620), .A2(n13978), .ZN(n13606) );
  NAND2_X1 U15615 ( .A1(P1_U3086), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n13605)
         );
  NAND2_X1 U15616 ( .A1(n13639), .A2(n13945), .ZN(n13604) );
  NAND4_X1 U15617 ( .A1(n13607), .A2(n13606), .A3(n13605), .A4(n13604), .ZN(
        n13608) );
  AOI21_X1 U15618 ( .B1(n14078), .B2(n13647), .A(n13608), .ZN(n13609) );
  OAI21_X1 U15619 ( .B1(n13610), .B2(n13650), .A(n13609), .ZN(P1_U3233) );
  INV_X1 U15620 ( .A(n13987), .ZN(n14401) );
  OAI21_X1 U15621 ( .B1(n13613), .B2(n13612), .A(n13611), .ZN(n13614) );
  NAND2_X1 U15622 ( .A1(n13614), .A2(n13626), .ZN(n13622) );
  NOR2_X1 U15623 ( .A1(n13644), .A2(n13984), .ZN(n13619) );
  OAI21_X1 U15624 ( .B1(n13617), .B2(n13616), .A(n13615), .ZN(n13618) );
  AOI211_X1 U15625 ( .C1(n13620), .C2(n13977), .A(n13619), .B(n13618), .ZN(
        n13621) );
  OAI211_X1 U15626 ( .C1(n14401), .C2(n13636), .A(n13622), .B(n13621), .ZN(
        P1_U3238) );
  OAI21_X1 U15627 ( .B1(n13625), .B2(n13624), .A(n13623), .ZN(n13627) );
  NAND2_X1 U15628 ( .A1(n13627), .A2(n13626), .ZN(n13635) );
  INV_X1 U15629 ( .A(n13849), .ZN(n13633) );
  AOI22_X1 U15630 ( .A1(n13639), .A2(n13847), .B1(P1_REG3_REG_26__SCAN_IN), 
        .B2(P1_U3086), .ZN(n13628) );
  OAI21_X1 U15631 ( .B1(n13630), .B2(n13629), .A(n13628), .ZN(n13631) );
  AOI21_X1 U15632 ( .B1(n13633), .B2(n13632), .A(n13631), .ZN(n13634) );
  OAI211_X1 U15633 ( .C1(n13854), .C2(n13636), .A(n13635), .B(n13634), .ZN(
        P1_U3240) );
  XNOR2_X1 U15634 ( .A(n13638), .B(n13637), .ZN(n13651) );
  NAND2_X1 U15635 ( .A1(n13639), .A2(n13655), .ZN(n13640) );
  OAI21_X1 U15636 ( .B1(P1_STATE_REG_SCAN_IN), .B2(n13641), .A(n13640), .ZN(
        n13642) );
  AOI21_X1 U15637 ( .B1(n13620), .B2(n13656), .A(n13642), .ZN(n13643) );
  OAI21_X1 U15638 ( .B1(n13645), .B2(n13644), .A(n13643), .ZN(n13646) );
  AOI21_X1 U15639 ( .B1(n13648), .B2(n13647), .A(n13646), .ZN(n13649) );
  OAI21_X1 U15640 ( .B1(n13651), .B2(n13650), .A(n13649), .ZN(P1_U3241) );
  MUX2_X1 U15641 ( .A(n13814), .B(P1_DATAO_REG_31__SCAN_IN), .S(n13667), .Z(
        P1_U3591) );
  MUX2_X1 U15642 ( .A(n13652), .B(P1_DATAO_REG_30__SCAN_IN), .S(n13667), .Z(
        P1_U3590) );
  MUX2_X1 U15643 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n13653), .S(P1_U4016), .Z(
        P1_U3589) );
  MUX2_X1 U15644 ( .A(n13654), .B(P1_DATAO_REG_28__SCAN_IN), .S(n13667), .Z(
        P1_U3588) );
  MUX2_X1 U15645 ( .A(n13847), .B(P1_DATAO_REG_27__SCAN_IN), .S(n13667), .Z(
        P1_U3587) );
  MUX2_X1 U15646 ( .A(n13866), .B(P1_DATAO_REG_26__SCAN_IN), .S(n13667), .Z(
        P1_U3586) );
  MUX2_X1 U15647 ( .A(n13887), .B(P1_DATAO_REG_25__SCAN_IN), .S(n13667), .Z(
        P1_U3585) );
  MUX2_X1 U15648 ( .A(n13865), .B(P1_DATAO_REG_24__SCAN_IN), .S(n13667), .Z(
        P1_U3584) );
  MUX2_X1 U15649 ( .A(n13888), .B(P1_DATAO_REG_23__SCAN_IN), .S(n13667), .Z(
        P1_U3583) );
  MUX2_X1 U15650 ( .A(n13936), .B(P1_DATAO_REG_22__SCAN_IN), .S(n13667), .Z(
        P1_U3582) );
  MUX2_X1 U15651 ( .A(n13945), .B(P1_DATAO_REG_21__SCAN_IN), .S(n13667), .Z(
        P1_U3581) );
  MUX2_X1 U15652 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n13935), .S(P1_U4016), .Z(
        P1_U3580) );
  MUX2_X1 U15653 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n13978), .S(P1_U4016), .Z(
        P1_U3579) );
  MUX2_X1 U15654 ( .A(n13977), .B(P1_DATAO_REG_17__SCAN_IN), .S(n13667), .Z(
        P1_U3577) );
  MUX2_X1 U15655 ( .A(n13655), .B(P1_DATAO_REG_16__SCAN_IN), .S(n13667), .Z(
        P1_U3576) );
  MUX2_X1 U15656 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n14385), .S(P1_U4016), .Z(
        P1_U3575) );
  MUX2_X1 U15657 ( .A(n13656), .B(P1_DATAO_REG_14__SCAN_IN), .S(n13667), .Z(
        P1_U3574) );
  MUX2_X1 U15658 ( .A(n14394), .B(P1_DATAO_REG_13__SCAN_IN), .S(n13667), .Z(
        P1_U3573) );
  MUX2_X1 U15659 ( .A(n13657), .B(P1_DATAO_REG_12__SCAN_IN), .S(n13667), .Z(
        P1_U3572) );
  MUX2_X1 U15660 ( .A(n13658), .B(P1_DATAO_REG_11__SCAN_IN), .S(n13667), .Z(
        P1_U3571) );
  MUX2_X1 U15661 ( .A(n13659), .B(P1_DATAO_REG_10__SCAN_IN), .S(n13667), .Z(
        P1_U3570) );
  MUX2_X1 U15662 ( .A(n13660), .B(P1_DATAO_REG_9__SCAN_IN), .S(n13667), .Z(
        P1_U3569) );
  MUX2_X1 U15663 ( .A(n13661), .B(P1_DATAO_REG_8__SCAN_IN), .S(n13667), .Z(
        P1_U3568) );
  MUX2_X1 U15664 ( .A(n13662), .B(P1_DATAO_REG_7__SCAN_IN), .S(n13667), .Z(
        P1_U3567) );
  MUX2_X1 U15665 ( .A(n13663), .B(P1_DATAO_REG_6__SCAN_IN), .S(n13667), .Z(
        P1_U3566) );
  MUX2_X1 U15666 ( .A(n13664), .B(P1_DATAO_REG_5__SCAN_IN), .S(n13667), .Z(
        P1_U3565) );
  MUX2_X1 U15667 ( .A(n13665), .B(P1_DATAO_REG_4__SCAN_IN), .S(n13667), .Z(
        P1_U3564) );
  MUX2_X1 U15668 ( .A(n13666), .B(P1_DATAO_REG_3__SCAN_IN), .S(n13667), .Z(
        P1_U3563) );
  MUX2_X1 U15669 ( .A(n14525), .B(P1_DATAO_REG_2__SCAN_IN), .S(n13667), .Z(
        P1_U3562) );
  MUX2_X1 U15670 ( .A(n6479), .B(P1_DATAO_REG_1__SCAN_IN), .S(n13667), .Z(
        P1_U3561) );
  MUX2_X1 U15671 ( .A(n14526), .B(P1_DATAO_REG_0__SCAN_IN), .S(n13667), .Z(
        P1_U3560) );
  OAI211_X1 U15672 ( .C1(n13679), .C2(n13668), .A(n14508), .B(n13692), .ZN(
        n13677) );
  MUX2_X1 U15673 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n9303), .S(n13669), .Z(
        n13670) );
  OAI21_X1 U15674 ( .B1(n9287), .B2(n13671), .A(n13670), .ZN(n13672) );
  NAND3_X1 U15675 ( .A1(n14504), .A2(n13686), .A3(n13672), .ZN(n13676) );
  NAND2_X1 U15676 ( .A1(n14490), .A2(n13673), .ZN(n13675) );
  AOI22_X1 U15677 ( .A1(n14497), .A2(P1_ADDR_REG_1__SCAN_IN), .B1(
        P1_REG3_REG_1__SCAN_IN), .B2(P1_U3086), .ZN(n13674) );
  NAND4_X1 U15678 ( .A1(n13677), .A2(n13676), .A3(n13675), .A4(n13674), .ZN(
        P1_U3244) );
  MUX2_X1 U15679 ( .A(n13679), .B(n13678), .S(n14121), .Z(n13681) );
  NAND2_X1 U15680 ( .A1(n13681), .A2(n13680), .ZN(n13682) );
  OAI211_X1 U15681 ( .C1(P1_IR_REG_0__SCAN_IN), .C2(n13683), .A(n13682), .B(
        P1_U4016), .ZN(n13728) );
  AOI22_X1 U15682 ( .A1(n14497), .A2(P1_ADDR_REG_2__SCAN_IN), .B1(
        P1_REG3_REG_2__SCAN_IN), .B2(P1_U3086), .ZN(n13696) );
  MUX2_X1 U15683 ( .A(n9564), .B(P1_REG1_REG_2__SCAN_IN), .S(n13689), .Z(
        n13684) );
  NAND3_X1 U15684 ( .A1(n13686), .A2(n13685), .A3(n13684), .ZN(n13687) );
  AND3_X1 U15685 ( .A1(n14504), .A2(n13705), .A3(n13687), .ZN(n13688) );
  AOI21_X1 U15686 ( .B1(n14490), .B2(n13689), .A(n13688), .ZN(n13695) );
  MUX2_X1 U15687 ( .A(n8844), .B(P1_REG2_REG_2__SCAN_IN), .S(n13689), .Z(
        n13690) );
  NAND3_X1 U15688 ( .A1(n13692), .A2(n13691), .A3(n13690), .ZN(n13693) );
  NAND3_X1 U15689 ( .A1(n14508), .A2(n13700), .A3(n13693), .ZN(n13694) );
  NAND4_X1 U15690 ( .A1(n13728), .A2(n13696), .A3(n13695), .A4(n13694), .ZN(
        P1_U3245) );
  NOR2_X1 U15691 ( .A1(n14495), .A2(n14142), .ZN(n13697) );
  AOI211_X1 U15692 ( .C1(n14490), .C2(n13703), .A(n13698), .B(n13697), .ZN(
        n13710) );
  MUX2_X1 U15693 ( .A(n9591), .B(P1_REG2_REG_3__SCAN_IN), .S(n13703), .Z(
        n13701) );
  NAND3_X1 U15694 ( .A1(n13701), .A2(n13700), .A3(n13699), .ZN(n13702) );
  NAND3_X1 U15695 ( .A1(n14508), .A2(n13713), .A3(n13702), .ZN(n13709) );
  MUX2_X1 U15696 ( .A(n9592), .B(P1_REG1_REG_3__SCAN_IN), .S(n13703), .Z(
        n13706) );
  NAND3_X1 U15697 ( .A1(n13706), .A2(n13705), .A3(n13704), .ZN(n13707) );
  NAND3_X1 U15698 ( .A1(n14504), .A2(n13718), .A3(n13707), .ZN(n13708) );
  NAND3_X1 U15699 ( .A1(n13710), .A2(n13709), .A3(n13708), .ZN(P1_U3246) );
  NAND2_X1 U15700 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(n14497), .ZN(n13727) );
  MUX2_X1 U15701 ( .A(n9610), .B(P1_REG2_REG_4__SCAN_IN), .S(n13721), .Z(
        n13711) );
  NAND3_X1 U15702 ( .A1(n13713), .A2(n13712), .A3(n13711), .ZN(n13714) );
  NAND3_X1 U15703 ( .A1(n14508), .A2(n13738), .A3(n13714), .ZN(n13725) );
  INV_X1 U15704 ( .A(n13715), .ZN(n13720) );
  NAND3_X1 U15705 ( .A1(n13718), .A2(n13717), .A3(n13716), .ZN(n13719) );
  NAND3_X1 U15706 ( .A1(n14504), .A2(n13720), .A3(n13719), .ZN(n13724) );
  NAND2_X1 U15707 ( .A1(n14490), .A2(n13721), .ZN(n13723) );
  AND4_X1 U15708 ( .A1(n13725), .A2(n13724), .A3(n13723), .A4(n13722), .ZN(
        n13726) );
  NAND3_X1 U15709 ( .A1(n13728), .A2(n13727), .A3(n13726), .ZN(P1_U3247) );
  INV_X1 U15710 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n14149) );
  OAI21_X1 U15711 ( .B1(n14495), .B2(n14149), .A(n13729), .ZN(n13730) );
  AOI21_X1 U15712 ( .B1(n13731), .B2(n14490), .A(n13730), .ZN(n13744) );
  OAI21_X1 U15713 ( .B1(n13734), .B2(n13733), .A(n13732), .ZN(n13735) );
  NAND2_X1 U15714 ( .A1(n14504), .A2(n13735), .ZN(n13743) );
  MUX2_X1 U15715 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n10303), .S(n13736), .Z(
        n13739) );
  NAND3_X1 U15716 ( .A1(n13739), .A2(n13738), .A3(n13737), .ZN(n13740) );
  NAND3_X1 U15717 ( .A1(n14508), .A2(n13741), .A3(n13740), .ZN(n13742) );
  NAND3_X1 U15718 ( .A1(n13744), .A2(n13743), .A3(n13742), .ZN(P1_U3248) );
  INV_X1 U15719 ( .A(P1_ADDR_REG_7__SCAN_IN), .ZN(n14154) );
  OAI21_X1 U15720 ( .B1(n14495), .B2(n14154), .A(n13745), .ZN(n13746) );
  AOI21_X1 U15721 ( .B1(n13747), .B2(n14490), .A(n13746), .ZN(n13760) );
  MUX2_X1 U15722 ( .A(n10319), .B(P1_REG2_REG_7__SCAN_IN), .S(n13747), .Z(
        n13748) );
  NAND3_X1 U15723 ( .A1(n13750), .A2(n13749), .A3(n13748), .ZN(n13751) );
  NAND3_X1 U15724 ( .A1(n14508), .A2(n13752), .A3(n13751), .ZN(n13759) );
  OR3_X1 U15725 ( .A1(n13755), .A2(n13754), .A3(n13753), .ZN(n13756) );
  NAND3_X1 U15726 ( .A1(n14504), .A2(n13757), .A3(n13756), .ZN(n13758) );
  NAND3_X1 U15727 ( .A1(n13760), .A2(n13759), .A3(n13758), .ZN(P1_U3250) );
  INV_X1 U15728 ( .A(n13761), .ZN(n13766) );
  NOR3_X1 U15729 ( .A1(n13764), .A2(n13763), .A3(n13762), .ZN(n13765) );
  OAI21_X1 U15730 ( .B1(n13766), .B2(n13765), .A(n14504), .ZN(n13777) );
  INV_X1 U15731 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n14136) );
  OAI21_X1 U15732 ( .B1(n14495), .B2(n14136), .A(n13767), .ZN(n13768) );
  AOI21_X1 U15733 ( .B1(n13769), .B2(n14490), .A(n13768), .ZN(n13776) );
  MUX2_X1 U15734 ( .A(n10238), .B(P1_REG2_REG_9__SCAN_IN), .S(n13769), .Z(
        n13770) );
  NAND3_X1 U15735 ( .A1(n13772), .A2(n13771), .A3(n13770), .ZN(n13773) );
  NAND3_X1 U15736 ( .A1(n14508), .A2(n13774), .A3(n13773), .ZN(n13775) );
  NAND3_X1 U15737 ( .A1(n13777), .A2(n13776), .A3(n13775), .ZN(P1_U3252) );
  OAI21_X1 U15738 ( .B1(n13779), .B2(n13778), .A(n14483), .ZN(n13780) );
  NAND2_X1 U15739 ( .A1(n13780), .A2(n14504), .ZN(n13791) );
  INV_X1 U15740 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n14135) );
  OAI21_X1 U15741 ( .B1(n14495), .B2(n14135), .A(n13781), .ZN(n13782) );
  AOI21_X1 U15742 ( .B1(n14490), .B2(n13783), .A(n13782), .ZN(n13790) );
  MUX2_X1 U15743 ( .A(n10625), .B(P1_REG2_REG_11__SCAN_IN), .S(n13783), .Z(
        n13784) );
  NAND3_X1 U15744 ( .A1(n13786), .A2(n13785), .A3(n13784), .ZN(n13787) );
  NAND3_X1 U15745 ( .A1(n14508), .A2(n13788), .A3(n13787), .ZN(n13789) );
  NAND3_X1 U15746 ( .A1(n13791), .A2(n13790), .A3(n13789), .ZN(P1_U3254) );
  NAND2_X1 U15747 ( .A1(n13797), .A2(n13792), .ZN(n13793) );
  NAND2_X1 U15748 ( .A1(n13794), .A2(n13793), .ZN(n13795) );
  XOR2_X1 U15749 ( .A(n13795), .B(P1_REG2_REG_19__SCAN_IN), .Z(n13805) );
  INV_X1 U15750 ( .A(n13805), .ZN(n13803) );
  NAND2_X1 U15751 ( .A1(n13797), .A2(n13796), .ZN(n13798) );
  NAND2_X1 U15752 ( .A1(n13799), .A2(n13798), .ZN(n13800) );
  XOR2_X1 U15753 ( .A(n13800), .B(P1_REG1_REG_19__SCAN_IN), .Z(n13804) );
  OAI21_X1 U15754 ( .B1(n13804), .B2(n13801), .A(n14501), .ZN(n13802) );
  AOI21_X1 U15755 ( .B1(n14508), .B2(n13803), .A(n13802), .ZN(n13808) );
  AOI22_X1 U15756 ( .A1(n13805), .A2(n14508), .B1(n13804), .B2(n14504), .ZN(
        n13807) );
  MUX2_X1 U15757 ( .A(n13808), .B(n13807), .S(n13806), .Z(n13810) );
  OAI211_X1 U15758 ( .C1(n13811), .C2(n14495), .A(n13810), .B(n13809), .ZN(
        P1_U3262) );
  NOR2_X1 U15759 ( .A1(n13818), .A2(n13819), .ZN(n13817) );
  XNOR2_X1 U15760 ( .A(n13817), .B(n13812), .ZN(n14016) );
  NAND2_X1 U15761 ( .A1(n14016), .A2(n14519), .ZN(n13816) );
  NAND2_X1 U15762 ( .A1(n13814), .A2(n13813), .ZN(n14020) );
  NOR2_X1 U15763 ( .A1(n14531), .A2(n14020), .ZN(n13820) );
  AOI21_X1 U15764 ( .B1(n14388), .B2(P1_REG2_REG_31__SCAN_IN), .A(n13820), 
        .ZN(n13815) );
  OAI211_X1 U15765 ( .C1(n14018), .C2(n14534), .A(n13816), .B(n13815), .ZN(
        P1_U3263) );
  INV_X1 U15766 ( .A(n13818), .ZN(n14022) );
  AOI21_X1 U15767 ( .B1(n13819), .B2(n13818), .A(n13817), .ZN(n14019) );
  NAND2_X1 U15768 ( .A1(n14019), .A2(n14519), .ZN(n13822) );
  AOI21_X1 U15769 ( .B1(n14388), .B2(P1_REG2_REG_30__SCAN_IN), .A(n13820), 
        .ZN(n13821) );
  OAI211_X1 U15770 ( .C1(n14022), .C2(n14534), .A(n13822), .B(n13821), .ZN(
        P1_U3264) );
  OAI21_X1 U15771 ( .B1(n13824), .B2(n13826), .A(n13823), .ZN(n14037) );
  NAND3_X1 U15772 ( .A1(n13826), .A2(n13844), .A3(n13825), .ZN(n13827) );
  AOI21_X1 U15773 ( .B1(n13828), .B2(n13827), .A(n14542), .ZN(n13832) );
  OAI22_X1 U15774 ( .A1(n13830), .A2(n14006), .B1(n13829), .B2(n14008), .ZN(
        n13831) );
  INV_X1 U15775 ( .A(n13833), .ZN(n13834) );
  AOI21_X1 U15776 ( .B1(n14038), .B2(n6880), .A(n13834), .ZN(n14039) );
  NOR2_X1 U15777 ( .A1(n13835), .A2(n14534), .ZN(n13839) );
  OAI22_X1 U15778 ( .A1(n13893), .A2(n13837), .B1(n13836), .B2(n14532), .ZN(
        n13838) );
  AOI211_X1 U15779 ( .C1(n14039), .C2(n14519), .A(n13839), .B(n13838), .ZN(
        n13841) );
  NAND2_X1 U15780 ( .A1(n14037), .A2(n14520), .ZN(n13840) );
  OAI211_X1 U15781 ( .C1(n14041), .C2(n14531), .A(n13841), .B(n13840), .ZN(
        P1_U3266) );
  XNOR2_X1 U15782 ( .A(n6472), .B(n13842), .ZN(n14047) );
  OAI21_X1 U15783 ( .B1(n13846), .B2(n13845), .A(n13844), .ZN(n13848) );
  AOI222_X1 U15784 ( .A1(n14392), .A2(n13848), .B1(n13847), .B2(n14524), .C1(
        n13887), .C2(n14527), .ZN(n14046) );
  OAI21_X1 U15785 ( .B1(n13849), .B2(n14532), .A(n14046), .ZN(n13850) );
  NAND2_X1 U15786 ( .A1(n13850), .A2(n13893), .ZN(n13857) );
  AND2_X1 U15787 ( .A1(n14043), .A2(n13864), .ZN(n13851) );
  NOR2_X1 U15788 ( .A1(n13852), .A2(n13851), .ZN(n14044) );
  OAI22_X1 U15789 ( .A1(n13854), .A2(n14534), .B1(n13853), .B2(n13893), .ZN(
        n13855) );
  AOI21_X1 U15790 ( .B1(n14044), .B2(n14519), .A(n13855), .ZN(n13856) );
  OAI211_X1 U15791 ( .C1(n14047), .C2(n14015), .A(n13857), .B(n13856), .ZN(
        P1_U3267) );
  XOR2_X1 U15792 ( .A(n13860), .B(n13858), .Z(n14055) );
  OAI21_X1 U15793 ( .B1(n13861), .B2(n13860), .A(n13859), .ZN(n13862) );
  INV_X1 U15794 ( .A(n13862), .ZN(n14053) );
  NAND2_X1 U15795 ( .A1(n13883), .A2(n14049), .ZN(n13863) );
  NAND2_X1 U15796 ( .A1(n13864), .A2(n13863), .ZN(n14051) );
  NOR2_X1 U15797 ( .A1(n14051), .A2(n13989), .ZN(n13875) );
  NAND2_X1 U15798 ( .A1(n13865), .A2(n14527), .ZN(n13868) );
  NAND2_X1 U15799 ( .A1(n13866), .A2(n14524), .ZN(n13867) );
  NAND2_X1 U15800 ( .A1(n13868), .A2(n13867), .ZN(n14048) );
  INV_X1 U15801 ( .A(n13869), .ZN(n13870) );
  AOI22_X1 U15802 ( .A1(n13893), .A2(n14048), .B1(n13870), .B2(n13996), .ZN(
        n13872) );
  NAND2_X1 U15803 ( .A1(n14388), .A2(P1_REG2_REG_25__SCAN_IN), .ZN(n13871) );
  OAI211_X1 U15804 ( .C1(n13873), .C2(n14534), .A(n13872), .B(n13871), .ZN(
        n13874) );
  AOI211_X1 U15805 ( .C1(n14053), .C2(n14383), .A(n13875), .B(n13874), .ZN(
        n13876) );
  OAI21_X1 U15806 ( .B1(n13877), .B2(n14055), .A(n13876), .ZN(P1_U3268) );
  AND2_X1 U15807 ( .A1(n13878), .A2(n13885), .ZN(n13879) );
  INV_X1 U15808 ( .A(n14059), .ZN(n13902) );
  INV_X1 U15809 ( .A(n13881), .ZN(n13892) );
  OR2_X1 U15810 ( .A1(n14056), .A2(n13905), .ZN(n13882) );
  NAND2_X1 U15811 ( .A1(n13883), .A2(n13882), .ZN(n14057) );
  OAI211_X1 U15812 ( .C1(n13886), .C2(n13885), .A(n13884), .B(n14392), .ZN(
        n13890) );
  AOI22_X1 U15813 ( .A1(n13888), .A2(n14527), .B1(n14524), .B2(n13887), .ZN(
        n13889) );
  NAND2_X1 U15814 ( .A1(n13890), .A2(n13889), .ZN(n13891) );
  AOI21_X1 U15815 ( .B1(n14059), .B2(n14523), .A(n13891), .ZN(n14061) );
  OAI21_X1 U15816 ( .B1(n13892), .B2(n14057), .A(n14061), .ZN(n13894) );
  NAND2_X1 U15817 ( .A1(n13894), .A2(n13893), .ZN(n13900) );
  INV_X1 U15818 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n13896) );
  OAI22_X1 U15819 ( .A1(n13893), .A2(n13896), .B1(n13895), .B2(n14532), .ZN(
        n13897) );
  AOI21_X1 U15820 ( .B1(n13898), .B2(n14398), .A(n13897), .ZN(n13899) );
  OAI211_X1 U15821 ( .C1(n13902), .C2(n13901), .A(n13900), .B(n13899), .ZN(
        P1_U3269) );
  XNOR2_X1 U15822 ( .A(n13904), .B(n7063), .ZN(n14066) );
  AOI21_X1 U15823 ( .B1(n14062), .B2(n13922), .A(n13905), .ZN(n14063) );
  AOI22_X1 U15824 ( .A1(n14531), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n13906), 
        .B2(n13996), .ZN(n13907) );
  OAI21_X1 U15825 ( .B1(n13908), .B2(n14534), .A(n13907), .ZN(n13914) );
  OAI21_X1 U15826 ( .B1(n6544), .B2(n7063), .A(n13909), .ZN(n13912) );
  INV_X1 U15827 ( .A(n13910), .ZN(n13911) );
  AOI21_X1 U15828 ( .B1(n13912), .B2(n14392), .A(n13911), .ZN(n14065) );
  NOR2_X1 U15829 ( .A1(n14065), .A2(n14388), .ZN(n13913) );
  AOI211_X1 U15830 ( .C1(n14063), .C2(n14519), .A(n13914), .B(n13913), .ZN(
        n13915) );
  OAI21_X1 U15831 ( .B1(n14015), .B2(n14066), .A(n13915), .ZN(P1_U3270) );
  XNOR2_X1 U15832 ( .A(n13920), .B(n6574), .ZN(n13916) );
  OAI222_X1 U15833 ( .A1(n14008), .A2(n13918), .B1(n14006), .B2(n13917), .C1(
        n14542), .C2(n13916), .ZN(n14068) );
  INV_X1 U15834 ( .A(n14068), .ZN(n13928) );
  OAI21_X1 U15835 ( .B1(n13921), .B2(n13920), .A(n13919), .ZN(n14070) );
  OAI21_X1 U15836 ( .B1(n11572), .B2(n6591), .A(n13922), .ZN(n14067) );
  AOI22_X1 U15837 ( .A1(n14531), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n13923), 
        .B2(n13996), .ZN(n13925) );
  NAND2_X1 U15838 ( .A1(n6886), .A2(n14398), .ZN(n13924) );
  OAI211_X1 U15839 ( .C1(n14067), .C2(n13989), .A(n13925), .B(n13924), .ZN(
        n13926) );
  AOI21_X1 U15840 ( .B1(n14070), .B2(n14383), .A(n13926), .ZN(n13927) );
  OAI21_X1 U15841 ( .B1(n13928), .B2(n14388), .A(n13927), .ZN(P1_U3271) );
  XOR2_X1 U15842 ( .A(n13929), .B(n13934), .Z(n14076) );
  AOI21_X1 U15843 ( .B1(n14072), .B2(n13952), .A(n6591), .ZN(n14073) );
  INV_X1 U15844 ( .A(n13930), .ZN(n13931) );
  AOI22_X1 U15845 ( .A1(n14531), .A2(P1_REG2_REG_21__SCAN_IN), .B1(n13931), 
        .B2(n13996), .ZN(n13932) );
  OAI21_X1 U15846 ( .B1(n6884), .B2(n14534), .A(n13932), .ZN(n13939) );
  XOR2_X1 U15847 ( .A(n13934), .B(n13933), .Z(n13937) );
  AOI222_X1 U15848 ( .A1(n14392), .A2(n13937), .B1(n13936), .B2(n14524), .C1(
        n13935), .C2(n14527), .ZN(n14075) );
  NOR2_X1 U15849 ( .A1(n14075), .A2(n14388), .ZN(n13938) );
  AOI211_X1 U15850 ( .C1(n14073), .C2(n14519), .A(n13939), .B(n13938), .ZN(
        n13940) );
  OAI21_X1 U15851 ( .B1(n14076), .B2(n14015), .A(n13940), .ZN(P1_U3272) );
  INV_X1 U15852 ( .A(n13941), .ZN(n13960) );
  OAI21_X1 U15853 ( .B1(n13960), .B2(n13942), .A(n13949), .ZN(n13944) );
  NAND3_X1 U15854 ( .A1(n13944), .A2(n14392), .A3(n13943), .ZN(n13947) );
  AOI22_X1 U15855 ( .A1(n13945), .A2(n14524), .B1(n14527), .B2(n13978), .ZN(
        n13946) );
  AND2_X1 U15856 ( .A1(n13947), .A2(n13946), .ZN(n14081) );
  OAI21_X1 U15857 ( .B1(n13950), .B2(n13949), .A(n13948), .ZN(n14082) );
  INV_X1 U15858 ( .A(n14082), .ZN(n13957) );
  NAND2_X1 U15859 ( .A1(n14078), .A2(n13965), .ZN(n13951) );
  NAND2_X1 U15860 ( .A1(n13952), .A2(n13951), .ZN(n14077) );
  AOI22_X1 U15861 ( .A1(n14388), .A2(P1_REG2_REG_20__SCAN_IN), .B1(n13953), 
        .B2(n13996), .ZN(n13955) );
  NAND2_X1 U15862 ( .A1(n14078), .A2(n14398), .ZN(n13954) );
  OAI211_X1 U15863 ( .C1(n14077), .C2(n13989), .A(n13955), .B(n13954), .ZN(
        n13956) );
  AOI21_X1 U15864 ( .B1(n13957), .B2(n14383), .A(n13956), .ZN(n13958) );
  OAI21_X1 U15865 ( .B1(n14531), .B2(n14081), .A(n13958), .ZN(P1_U3273) );
  XNOR2_X1 U15866 ( .A(n13959), .B(n13962), .ZN(n14087) );
  INV_X1 U15867 ( .A(n14087), .ZN(n13973) );
  AOI21_X1 U15868 ( .B1(n13962), .B2(n13961), .A(n13960), .ZN(n13963) );
  OAI222_X1 U15869 ( .A1(n14008), .A2(n13964), .B1(n14006), .B2(n14009), .C1(
        n14542), .C2(n13963), .ZN(n14085) );
  OAI21_X1 U15870 ( .B1(n14083), .B2(n13983), .A(n13965), .ZN(n14084) );
  INV_X1 U15871 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n13967) );
  OAI22_X1 U15872 ( .A1(n13893), .A2(n13967), .B1(n13966), .B2(n14532), .ZN(
        n13968) );
  AOI21_X1 U15873 ( .B1(n13969), .B2(n14398), .A(n13968), .ZN(n13970) );
  OAI21_X1 U15874 ( .B1(n14084), .B2(n13989), .A(n13970), .ZN(n13971) );
  AOI21_X1 U15875 ( .B1(n14085), .B2(n13893), .A(n13971), .ZN(n13972) );
  OAI21_X1 U15876 ( .B1(n14015), .B2(n13973), .A(n13972), .ZN(P1_U3274) );
  XNOR2_X1 U15877 ( .A(n13974), .B(n13975), .ZN(n14404) );
  XNOR2_X1 U15878 ( .A(n13976), .B(n13975), .ZN(n13980) );
  AOI22_X1 U15879 ( .A1(n13978), .A2(n14524), .B1(n14527), .B2(n13977), .ZN(
        n13979) );
  OAI21_X1 U15880 ( .B1(n13980), .B2(n14542), .A(n13979), .ZN(n13981) );
  AOI21_X1 U15881 ( .B1(n14404), .B2(n14523), .A(n13981), .ZN(n14406) );
  AND2_X1 U15882 ( .A1(n13987), .A2(n13993), .ZN(n13982) );
  OR2_X1 U15883 ( .A1(n13983), .A2(n13982), .ZN(n14402) );
  INV_X1 U15884 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n13985) );
  OAI22_X1 U15885 ( .A1(n13893), .A2(n13985), .B1(n13984), .B2(n14532), .ZN(
        n13986) );
  AOI21_X1 U15886 ( .B1(n13987), .B2(n14398), .A(n13986), .ZN(n13988) );
  OAI21_X1 U15887 ( .B1(n14402), .B2(n13989), .A(n13988), .ZN(n13990) );
  AOI21_X1 U15888 ( .B1(n14404), .B2(n14520), .A(n13990), .ZN(n13991) );
  OAI21_X1 U15889 ( .B1(n14406), .B2(n14388), .A(n13991), .ZN(P1_U3275) );
  XNOR2_X1 U15890 ( .A(n13992), .B(n14001), .ZN(n14094) );
  INV_X1 U15891 ( .A(n13993), .ZN(n13994) );
  AOI21_X1 U15892 ( .B1(n14090), .B2(n14410), .A(n13994), .ZN(n14091) );
  INV_X1 U15893 ( .A(n13995), .ZN(n13997) );
  AOI22_X1 U15894 ( .A1(n14531), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n13997), 
        .B2(n13996), .ZN(n13998) );
  OAI21_X1 U15895 ( .B1(n13999), .B2(n14534), .A(n13998), .ZN(n14013) );
  INV_X1 U15896 ( .A(n14000), .ZN(n14005) );
  AOI21_X1 U15897 ( .B1(n14003), .B2(n14002), .A(n14001), .ZN(n14004) );
  NOR3_X1 U15898 ( .A1(n14005), .A2(n14004), .A3(n14542), .ZN(n14011) );
  OAI22_X1 U15899 ( .A1(n14009), .A2(n14008), .B1(n14007), .B2(n14006), .ZN(
        n14010) );
  NOR2_X1 U15900 ( .A1(n14011), .A2(n14010), .ZN(n14093) );
  NOR2_X1 U15901 ( .A1(n14093), .A2(n14388), .ZN(n14012) );
  AOI211_X1 U15902 ( .C1(n14091), .C2(n14519), .A(n14013), .B(n14012), .ZN(
        n14014) );
  OAI21_X1 U15903 ( .B1(n14015), .B2(n14094), .A(n14014), .ZN(P1_U3276) );
  INV_X1 U15904 ( .A(n14596), .ZN(n14581) );
  NAND2_X1 U15905 ( .A1(n14016), .A2(n14581), .ZN(n14017) );
  OAI211_X1 U15906 ( .C1(n14018), .C2(n14606), .A(n14017), .B(n14020), .ZN(
        n14095) );
  MUX2_X1 U15907 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n14095), .S(n14630), .Z(
        P1_U3559) );
  NAND2_X1 U15908 ( .A1(n14019), .A2(n14581), .ZN(n14021) );
  OAI211_X1 U15909 ( .C1(n14022), .C2(n14606), .A(n14021), .B(n14020), .ZN(
        n14096) );
  MUX2_X1 U15910 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n14096), .S(n14630), .Z(
        P1_U3558) );
  OAI211_X1 U15911 ( .C1(n14027), .C2(n14606), .A(n14026), .B(n14025), .ZN(
        n14028) );
  AOI22_X1 U15912 ( .A1(n14033), .A2(n14581), .B1(n14580), .B2(n14032), .ZN(
        n14034) );
  MUX2_X1 U15913 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n14098), .S(n14630), .Z(
        P1_U3556) );
  INV_X1 U15914 ( .A(n14037), .ZN(n14042) );
  AOI22_X1 U15915 ( .A1(n14039), .A2(n14581), .B1(n14580), .B2(n14038), .ZN(
        n14040) );
  OAI211_X1 U15916 ( .C1(n14042), .C2(n14585), .A(n14041), .B(n14040), .ZN(
        n14099) );
  MUX2_X1 U15917 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n14099), .S(n14630), .Z(
        P1_U3555) );
  AOI22_X1 U15918 ( .A1(n14044), .A2(n14581), .B1(n14580), .B2(n14043), .ZN(
        n14045) );
  OAI211_X1 U15919 ( .C1(n14047), .C2(n14541), .A(n14046), .B(n14045), .ZN(
        n14100) );
  MUX2_X1 U15920 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n14100), .S(n14630), .Z(
        P1_U3554) );
  AOI21_X1 U15921 ( .B1(n14049), .B2(n14580), .A(n14048), .ZN(n14050) );
  OAI21_X1 U15922 ( .B1(n14051), .B2(n14596), .A(n14050), .ZN(n14052) );
  AOI21_X1 U15923 ( .B1(n14053), .B2(n14609), .A(n14052), .ZN(n14054) );
  OAI21_X1 U15924 ( .B1(n14542), .B2(n14055), .A(n14054), .ZN(n14101) );
  MUX2_X1 U15925 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n14101), .S(n14630), .Z(
        P1_U3553) );
  OAI22_X1 U15926 ( .A1(n14057), .A2(n14596), .B1(n14056), .B2(n14606), .ZN(
        n14058) );
  AOI21_X1 U15927 ( .B1(n14059), .B2(n14599), .A(n14058), .ZN(n14060) );
  NAND2_X1 U15928 ( .A1(n14061), .A2(n14060), .ZN(n14102) );
  MUX2_X1 U15929 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n14102), .S(n14630), .Z(
        P1_U3552) );
  AOI22_X1 U15930 ( .A1(n14063), .A2(n14581), .B1(n14580), .B2(n14062), .ZN(
        n14064) );
  OAI211_X1 U15931 ( .C1(n14066), .C2(n14541), .A(n14065), .B(n14064), .ZN(
        n14103) );
  MUX2_X1 U15932 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n14103), .S(n14630), .Z(
        P1_U3551) );
  OAI22_X1 U15933 ( .A1(n14067), .A2(n14596), .B1(n11572), .B2(n14606), .ZN(
        n14069) );
  AOI211_X1 U15934 ( .C1(n14609), .C2(n14070), .A(n14069), .B(n14068), .ZN(
        n14071) );
  INV_X1 U15935 ( .A(n14071), .ZN(n14104) );
  MUX2_X1 U15936 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n14104), .S(n14630), .Z(
        P1_U3550) );
  AOI22_X1 U15937 ( .A1(n14073), .A2(n14581), .B1(n14580), .B2(n14072), .ZN(
        n14074) );
  OAI211_X1 U15938 ( .C1(n14076), .C2(n14541), .A(n14075), .B(n14074), .ZN(
        n14105) );
  MUX2_X1 U15939 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n14105), .S(n14630), .Z(
        P1_U3549) );
  INV_X1 U15940 ( .A(n14077), .ZN(n14079) );
  AOI22_X1 U15941 ( .A1(n14079), .A2(n14581), .B1(n14580), .B2(n14078), .ZN(
        n14080) );
  OAI211_X1 U15942 ( .C1(n14082), .C2(n14541), .A(n14081), .B(n14080), .ZN(
        n14106) );
  MUX2_X1 U15943 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n14106), .S(n14630), .Z(
        P1_U3548) );
  INV_X1 U15944 ( .A(P1_REG1_REG_19__SCAN_IN), .ZN(n14088) );
  OAI22_X1 U15945 ( .A1(n14084), .A2(n14596), .B1(n14083), .B2(n14606), .ZN(
        n14086) );
  AOI211_X1 U15946 ( .C1(n14087), .C2(n14609), .A(n14086), .B(n14085), .ZN(
        n14107) );
  MUX2_X1 U15947 ( .A(n14088), .B(n14107), .S(n14630), .Z(n14089) );
  INV_X1 U15948 ( .A(n14089), .ZN(P1_U3547) );
  AOI22_X1 U15949 ( .A1(n14091), .A2(n14581), .B1(n14580), .B2(n14090), .ZN(
        n14092) );
  OAI211_X1 U15950 ( .C1(n14094), .C2(n14541), .A(n14093), .B(n14092), .ZN(
        n14110) );
  MUX2_X1 U15951 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n14110), .S(n14630), .Z(
        P1_U3545) );
  MUX2_X1 U15952 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n14095), .S(n14613), .Z(
        P1_U3527) );
  MUX2_X1 U15953 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n14096), .S(n14613), .Z(
        P1_U3526) );
  MUX2_X1 U15954 ( .A(P1_REG0_REG_28__SCAN_IN), .B(n14098), .S(n14613), .Z(
        P1_U3524) );
  MUX2_X1 U15955 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n14099), .S(n14613), .Z(
        P1_U3523) );
  MUX2_X1 U15956 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n14100), .S(n14613), .Z(
        P1_U3522) );
  MUX2_X1 U15957 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n14101), .S(n14613), .Z(
        P1_U3521) );
  MUX2_X1 U15958 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n14102), .S(n14613), .Z(
        P1_U3520) );
  MUX2_X1 U15959 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n14103), .S(n14613), .Z(
        P1_U3519) );
  MUX2_X1 U15960 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n14104), .S(n14613), .Z(
        P1_U3518) );
  MUX2_X1 U15961 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n14105), .S(n14613), .Z(
        P1_U3517) );
  MUX2_X1 U15962 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n14106), .S(n14613), .Z(
        P1_U3516) );
  INV_X1 U15963 ( .A(P1_REG0_REG_19__SCAN_IN), .ZN(n14108) );
  MUX2_X1 U15964 ( .A(n14108), .B(n14107), .S(n14613), .Z(n14109) );
  INV_X1 U15965 ( .A(n14109), .ZN(P1_U3515) );
  MUX2_X1 U15966 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n14110), .S(n14613), .Z(
        P1_U3510) );
  NOR4_X1 U15967 ( .A1(n14112), .A2(P1_IR_REG_30__SCAN_IN), .A3(n14111), .A4(
        P1_U3086), .ZN(n14113) );
  AOI21_X1 U15968 ( .B1(n14114), .B2(P2_DATAO_REG_31__SCAN_IN), .A(n14113), 
        .ZN(n14115) );
  OAI21_X1 U15969 ( .B1(n14116), .B2(n14119), .A(n14115), .ZN(P1_U3324) );
  OAI222_X1 U15970 ( .A1(n14124), .A2(n14123), .B1(n14130), .B2(n14122), .C1(
        P1_U3086), .C2(n14121), .ZN(P1_U3328) );
  OAI222_X1 U15971 ( .A1(P1_U3086), .A2(n14127), .B1(n14130), .B2(n14126), 
        .C1(n14125), .C2(n14124), .ZN(P1_U3329) );
  OAI222_X1 U15972 ( .A1(n14124), .A2(n14131), .B1(n14130), .B2(n14129), .C1(
        P1_U3086), .C2(n14128), .ZN(P1_U3330) );
  MUX2_X1 U15973 ( .A(n14132), .B(n14544), .S(P1_STATE_REG_SCAN_IN), .Z(
        P1_U3333) );
  INV_X1 U15974 ( .A(n14133), .ZN(n14134) );
  MUX2_X1 U15975 ( .A(n14134), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3355) );
  INV_X1 U15976 ( .A(P2_ADDR_REG_17__SCAN_IN), .ZN(n14238) );
  INV_X1 U15977 ( .A(P2_ADDR_REG_16__SCAN_IN), .ZN(n14478) );
  INV_X1 U15978 ( .A(P2_ADDR_REG_14__SCAN_IN), .ZN(n14221) );
  XOR2_X1 U15979 ( .A(P3_ADDR_REG_14__SCAN_IN), .B(n14225), .Z(n14223) );
  INV_X1 U15980 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n14217) );
  INV_X1 U15981 ( .A(P3_ADDR_REG_12__SCAN_IN), .ZN(n14166) );
  INV_X1 U15982 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n14496) );
  XNOR2_X1 U15983 ( .A(n14496), .B(n14166), .ZN(n14213) );
  INV_X1 U15984 ( .A(P3_ADDR_REG_11__SCAN_IN), .ZN(n14876) );
  XNOR2_X1 U15985 ( .A(n14135), .B(n14876), .ZN(n14211) );
  INV_X1 U15986 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n14161) );
  INV_X1 U15987 ( .A(P3_ADDR_REG_9__SCAN_IN), .ZN(n14159) );
  XNOR2_X1 U15988 ( .A(n14136), .B(n14159), .ZN(n14168) );
  XNOR2_X1 U15989 ( .A(n14137), .B(n14853), .ZN(n14202) );
  XOR2_X1 U15990 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n14833), .Z(n14195) );
  NAND2_X1 U15991 ( .A1(P3_ADDR_REG_3__SCAN_IN), .A2(n14141), .ZN(n14144) );
  NAND2_X1 U15992 ( .A1(P3_ADDR_REG_4__SCAN_IN), .A2(n14145), .ZN(n14147) );
  NAND2_X1 U15993 ( .A1(n14170), .A2(n14171), .ZN(n14146) );
  NAND2_X1 U15994 ( .A1(P3_ADDR_REG_5__SCAN_IN), .A2(n14148), .ZN(n14151) );
  NAND2_X1 U15995 ( .A1(n14189), .A2(n14149), .ZN(n14150) );
  NAND2_X1 U15996 ( .A1(n14151), .A2(n14150), .ZN(n14196) );
  NAND2_X1 U15997 ( .A1(n14195), .A2(n14196), .ZN(n14152) );
  NAND2_X1 U15998 ( .A1(P3_ADDR_REG_7__SCAN_IN), .A2(n14153), .ZN(n14156) );
  XOR2_X1 U15999 ( .A(n14153), .B(P3_ADDR_REG_7__SCAN_IN), .Z(n14199) );
  NAND2_X1 U16000 ( .A1(n14199), .A2(n14154), .ZN(n14155) );
  NAND2_X1 U16001 ( .A1(n14156), .A2(n14155), .ZN(n14203) );
  NAND2_X1 U16002 ( .A1(n14202), .A2(n14203), .ZN(n14157) );
  NAND2_X1 U16003 ( .A1(n14168), .A2(n14169), .ZN(n14158) );
  NAND2_X1 U16004 ( .A1(n14161), .A2(n14160), .ZN(n14163) );
  XOR2_X1 U16005 ( .A(n14161), .B(n14160), .Z(n14208) );
  NAND2_X1 U16006 ( .A1(n14208), .A2(P3_ADDR_REG_10__SCAN_IN), .ZN(n14162) );
  NAND2_X1 U16007 ( .A1(n14163), .A2(n14162), .ZN(n14212) );
  NAND2_X1 U16008 ( .A1(n14211), .A2(n14212), .ZN(n14164) );
  NAND2_X1 U16009 ( .A1(n14213), .A2(n14214), .ZN(n14165) );
  OR2_X1 U16010 ( .A1(n14217), .A2(P3_ADDR_REG_13__SCAN_IN), .ZN(n14167) );
  XOR2_X1 U16011 ( .A(n14223), .B(n14222), .Z(n14469) );
  XNOR2_X1 U16012 ( .A(n14169), .B(n14168), .ZN(n14206) );
  NAND2_X1 U16013 ( .A1(P2_ADDR_REG_4__SCAN_IN), .A2(n14172), .ZN(n14188) );
  INV_X1 U16014 ( .A(P2_ADDR_REG_2__SCAN_IN), .ZN(n14182) );
  XNOR2_X1 U16015 ( .A(n14174), .B(n14173), .ZN(n14250) );
  XNOR2_X1 U16016 ( .A(n14175), .B(n14176), .ZN(n14178) );
  NAND2_X1 U16017 ( .A1(P2_ADDR_REG_1__SCAN_IN), .A2(n14178), .ZN(n14180) );
  AOI21_X1 U16018 ( .B1(P1_ADDR_REG_0__SCAN_IN), .B2(n14177), .A(n14176), .ZN(
        n15248) );
  INV_X1 U16019 ( .A(P2_ADDR_REG_0__SCAN_IN), .ZN(n15247) );
  NOR2_X1 U16020 ( .A1(n15248), .A2(n15247), .ZN(n15253) );
  NAND2_X1 U16021 ( .A1(n14180), .A2(n14179), .ZN(n14251) );
  NAND2_X1 U16022 ( .A1(n14250), .A2(n14251), .ZN(n14181) );
  NOR2_X1 U16023 ( .A1(n14250), .A2(n14251), .ZN(n14249) );
  XOR2_X1 U16024 ( .A(P1_ADDR_REG_3__SCAN_IN), .B(n14183), .Z(n14184) );
  NAND2_X1 U16025 ( .A1(n14185), .A2(n14184), .ZN(n14187) );
  NAND2_X1 U16026 ( .A1(n14187), .A2(n14186), .ZN(n15244) );
  XOR2_X1 U16027 ( .A(P1_ADDR_REG_5__SCAN_IN), .B(n14189), .Z(n14190) );
  NOR2_X1 U16028 ( .A1(n14191), .A2(n14190), .ZN(n14193) );
  XNOR2_X1 U16029 ( .A(n14190), .B(n14191), .ZN(n15246) );
  NOR2_X1 U16030 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n15246), .ZN(n14192) );
  NAND2_X1 U16031 ( .A1(n14194), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n14197) );
  XNOR2_X1 U16032 ( .A(n14196), .B(n14195), .ZN(n14253) );
  NOR2_X1 U16033 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n14198), .ZN(n14201) );
  XOR2_X1 U16034 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n14199), .Z(n15249) );
  NOR2_X1 U16035 ( .A1(n15250), .A2(n15249), .ZN(n14200) );
  XNOR2_X1 U16036 ( .A(n14203), .B(n14202), .ZN(n14204) );
  XOR2_X1 U16037 ( .A(n14208), .B(P3_ADDR_REG_10__SCAN_IN), .Z(n14209) );
  XNOR2_X1 U16038 ( .A(n14212), .B(n14211), .ZN(n14458) );
  XNOR2_X1 U16039 ( .A(n14214), .B(n14213), .ZN(n14216) );
  XNOR2_X1 U16040 ( .A(n14216), .B(n14215), .ZN(n14461) );
  XOR2_X1 U16041 ( .A(n14217), .B(P3_ADDR_REG_13__SCAN_IN), .Z(n14219) );
  XNOR2_X1 U16042 ( .A(n14219), .B(n14218), .ZN(n14463) );
  INV_X1 U16043 ( .A(P2_ADDR_REG_13__SCAN_IN), .ZN(n14465) );
  NAND2_X1 U16044 ( .A1(n14469), .A2(n14468), .ZN(n14220) );
  INV_X1 U16045 ( .A(P3_ADDR_REG_15__SCAN_IN), .ZN(n14229) );
  XOR2_X1 U16046 ( .A(P1_ADDR_REG_15__SCAN_IN), .B(n14229), .Z(n14226) );
  NAND2_X1 U16047 ( .A1(n14223), .A2(n14222), .ZN(n14224) );
  XOR2_X1 U16048 ( .A(n14226), .B(n14230), .Z(n14472) );
  XOR2_X1 U16049 ( .A(P3_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .Z(n14234) );
  AND2_X1 U16050 ( .A1(n14229), .A2(P1_ADDR_REG_15__SCAN_IN), .ZN(n14231) );
  OAI22_X1 U16051 ( .A1(n14231), .A2(n14230), .B1(P1_ADDR_REG_15__SCAN_IN), 
        .B2(n14229), .ZN(n14233) );
  XOR2_X1 U16052 ( .A(n14234), .B(n14233), .Z(n14476) );
  NAND2_X1 U16053 ( .A1(n14477), .A2(n14476), .ZN(n14475) );
  INV_X1 U16054 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n14239) );
  INV_X1 U16055 ( .A(P3_ADDR_REG_16__SCAN_IN), .ZN(n14236) );
  NOR2_X1 U16056 ( .A1(n14234), .A2(n14233), .ZN(n14235) );
  AOI21_X1 U16057 ( .B1(P1_ADDR_REG_16__SCAN_IN), .B2(n14236), .A(n14235), 
        .ZN(n14240) );
  XOR2_X1 U16058 ( .A(n14239), .B(n14240), .Z(n14241) );
  XNOR2_X1 U16059 ( .A(P3_ADDR_REG_17__SCAN_IN), .B(n14241), .ZN(n14269) );
  NAND2_X1 U16060 ( .A1(n14270), .A2(n14269), .ZN(n14237) );
  NAND2_X1 U16061 ( .A1(n14240), .A2(n14239), .ZN(n14243) );
  NAND2_X1 U16062 ( .A1(P3_ADDR_REG_17__SCAN_IN), .A2(n14241), .ZN(n14242) );
  NAND2_X1 U16063 ( .A1(n14243), .A2(n14242), .ZN(n15234) );
  XOR2_X1 U16064 ( .A(n12259), .B(P1_ADDR_REG_18__SCAN_IN), .Z(n15235) );
  XNOR2_X1 U16065 ( .A(n15234), .B(n15235), .ZN(n14245) );
  NOR2_X1 U16066 ( .A1(n14244), .A2(n14245), .ZN(n15040) );
  NOR2_X1 U16067 ( .A1(n15040), .A2(n15039), .ZN(n14246) );
  XOR2_X1 U16068 ( .A(P2_ADDR_REG_18__SCAN_IN), .B(n14246), .Z(SUB_1596_U62)
         );
  AOI21_X1 U16069 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(
        P3_WR_REG_SCAN_IN), .ZN(n14247) );
  OAI21_X1 U16070 ( .B1(P2_WR_REG_SCAN_IN), .B2(P1_WR_REG_SCAN_IN), .A(n14247), 
        .ZN(U28) );
  INV_X1 U16071 ( .A(P1_RD_REG_SCAN_IN), .ZN(n14248) );
  INV_X1 U16072 ( .A(P3_RD_REG_SCAN_IN), .ZN(n15168) );
  OAI221_X1 U16073 ( .B1(P2_RD_REG_SCAN_IN), .B2(P1_RD_REG_SCAN_IN), .C1(n6729), .C2(n14248), .A(n15168), .ZN(U29) );
  AOI21_X1 U16074 ( .B1(n14251), .B2(n14250), .A(n14249), .ZN(n14252) );
  XOR2_X1 U16075 ( .A(n14252), .B(P2_ADDR_REG_2__SCAN_IN), .Z(SUB_1596_U61) );
  XOR2_X1 U16076 ( .A(n14254), .B(n14253), .Z(SUB_1596_U57) );
  XNOR2_X1 U16077 ( .A(n14255), .B(P2_ADDR_REG_8__SCAN_IN), .ZN(SUB_1596_U55)
         );
  XOR2_X1 U16078 ( .A(n14256), .B(P2_ADDR_REG_9__SCAN_IN), .Z(SUB_1596_U54) );
  NOR2_X1 U16079 ( .A1(n14258), .A2(n14257), .ZN(n14259) );
  XOR2_X1 U16080 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(n14259), .Z(SUB_1596_U70)
         );
  OAI22_X1 U16081 ( .A1(n14261), .A2(n14596), .B1(n14260), .B2(n14606), .ZN(
        n14262) );
  AOI21_X1 U16082 ( .B1(n14263), .B2(n14599), .A(n14262), .ZN(n14264) );
  AND2_X1 U16083 ( .A1(n14265), .A2(n14264), .ZN(n14267) );
  INV_X1 U16084 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n14266) );
  AOI22_X1 U16085 ( .A1(n14613), .A2(n14267), .B1(n14266), .B2(n14611), .ZN(
        P1_U3495) );
  AOI22_X1 U16086 ( .A1(n14630), .A2(n14267), .B1(n10608), .B2(n14627), .ZN(
        P1_U3540) );
  AOI21_X1 U16087 ( .B1(n14270), .B2(n14269), .A(n14268), .ZN(n14271) );
  XOR2_X1 U16088 ( .A(n14271), .B(P2_ADDR_REG_17__SCAN_IN), .Z(SUB_1596_U63)
         );
  INV_X1 U16089 ( .A(n14272), .ZN(n14273) );
  AOI21_X1 U16090 ( .B1(n14275), .B2(n14274), .A(n14273), .ZN(n14285) );
  OAI211_X1 U16091 ( .C1(n14279), .C2(n14278), .A(n14277), .B(n14276), .ZN(
        n14280) );
  OAI21_X1 U16092 ( .B1(n14282), .B2(n14281), .A(n14280), .ZN(n14283) );
  INV_X1 U16093 ( .A(n14283), .ZN(n14284) );
  OAI211_X1 U16094 ( .C1(n14287), .C2(n14286), .A(n14285), .B(n14284), .ZN(
        P3_U3181) );
  OR2_X1 U16095 ( .A1(n14288), .A2(n14298), .ZN(n14289) );
  AOI22_X1 U16096 ( .A1(n15038), .A2(n6509), .B1(n14290), .B2(n15036), .ZN(
        P3_U3490) );
  OAI21_X1 U16097 ( .B1(n14292), .B2(n14298), .A(n14291), .ZN(n14312) );
  OAI22_X1 U16098 ( .A1(n15036), .A2(n14312), .B1(P3_REG1_REG_30__SCAN_IN), 
        .B2(n15038), .ZN(n14293) );
  INV_X1 U16099 ( .A(n14293), .ZN(P3_U3489) );
  AOI211_X1 U16100 ( .C1(n14983), .C2(n14296), .A(n14295), .B(n14294), .ZN(
        n14315) );
  INV_X1 U16101 ( .A(P3_REG1_REG_14__SCAN_IN), .ZN(n14297) );
  AOI22_X1 U16102 ( .A1(n15038), .A2(n14315), .B1(n14297), .B2(n15036), .ZN(
        P3_U3473) );
  NOR2_X1 U16103 ( .A1(n14299), .A2(n14298), .ZN(n14301) );
  AOI211_X1 U16104 ( .C1(n14302), .C2(n14983), .A(n14301), .B(n14300), .ZN(
        n14317) );
  AOI22_X1 U16105 ( .A1(n15038), .A2(n14317), .B1(n14303), .B2(n15036), .ZN(
        P3_U3472) );
  AOI211_X1 U16106 ( .C1(n14306), .C2(n14983), .A(n14305), .B(n14304), .ZN(
        n14319) );
  AOI22_X1 U16107 ( .A1(n15038), .A2(n14319), .B1(n14307), .B2(n15036), .ZN(
        P3_U3471) );
  AOI211_X1 U16108 ( .C1(n14983), .C2(n14310), .A(n14309), .B(n14308), .ZN(
        n14321) );
  AOI22_X1 U16109 ( .A1(n15038), .A2(n14321), .B1(n14881), .B2(n15036), .ZN(
        P3_U3470) );
  INV_X1 U16110 ( .A(P3_REG0_REG_31__SCAN_IN), .ZN(n14311) );
  AOI22_X1 U16111 ( .A1(n15015), .A2(n6509), .B1(n14311), .B2(n8422), .ZN(
        P3_U3458) );
  OAI22_X1 U16112 ( .A1(n8422), .A2(n14312), .B1(P3_REG0_REG_30__SCAN_IN), 
        .B2(n15015), .ZN(n14313) );
  INV_X1 U16113 ( .A(n14313), .ZN(P3_U3457) );
  INV_X1 U16114 ( .A(P3_REG0_REG_14__SCAN_IN), .ZN(n14314) );
  AOI22_X1 U16115 ( .A1(n15015), .A2(n14315), .B1(n14314), .B2(n8422), .ZN(
        P3_U3432) );
  INV_X1 U16116 ( .A(P3_REG0_REG_13__SCAN_IN), .ZN(n14316) );
  AOI22_X1 U16117 ( .A1(n15015), .A2(n14317), .B1(n14316), .B2(n8422), .ZN(
        P3_U3429) );
  INV_X1 U16118 ( .A(P3_REG0_REG_12__SCAN_IN), .ZN(n14318) );
  AOI22_X1 U16119 ( .A1(n15015), .A2(n14319), .B1(n14318), .B2(n8422), .ZN(
        P3_U3426) );
  INV_X1 U16120 ( .A(P3_REG0_REG_11__SCAN_IN), .ZN(n14320) );
  AOI22_X1 U16121 ( .A1(n15015), .A2(n14321), .B1(n14320), .B2(n8422), .ZN(
        P3_U3423) );
  OAI22_X1 U16122 ( .A1(n10740), .A2(n14324), .B1(n14323), .B2(n14322), .ZN(
        n14337) );
  OAI21_X1 U16123 ( .B1(n14327), .B2(n14326), .A(n14325), .ZN(n14329) );
  AOI222_X1 U16124 ( .A1(n14331), .A2(n14342), .B1(n14337), .B2(n14330), .C1(
        n14329), .C2(n14328), .ZN(n14333) );
  OAI211_X1 U16125 ( .C1(n14334), .C2(n14339), .A(n14333), .B(n14332), .ZN(
        P2_U3187) );
  XNOR2_X1 U16126 ( .A(n14336), .B(n14335), .ZN(n14338) );
  AOI21_X1 U16127 ( .B1(n14338), .B2(n14740), .A(n14337), .ZN(n14363) );
  INV_X1 U16128 ( .A(n14339), .ZN(n14340) );
  AOI222_X1 U16129 ( .A1(n14342), .A2(n14341), .B1(P2_REG2_REG_14__SCAN_IN), 
        .B2(n14731), .C1(n14719), .C2(n14340), .ZN(n14351) );
  AOI21_X1 U16130 ( .B1(n14345), .B2(n14344), .A(n14343), .ZN(n14366) );
  INV_X1 U16131 ( .A(n14346), .ZN(n14348) );
  OAI211_X1 U16132 ( .C1(n14362), .C2(n14348), .A(n14714), .B(n14347), .ZN(
        n14361) );
  INV_X1 U16133 ( .A(n14361), .ZN(n14349) );
  AOI22_X1 U16134 ( .A1(n14366), .A2(n14727), .B1(n14725), .B2(n14349), .ZN(
        n14350) );
  OAI211_X1 U16135 ( .C1(n14731), .C2(n14363), .A(n14351), .B(n14350), .ZN(
        P2_U3251) );
  NOR2_X1 U16136 ( .A1(n14353), .A2(n14352), .ZN(n14358) );
  OAI211_X1 U16137 ( .C1(n14356), .C2(n14774), .A(n14355), .B(n14354), .ZN(
        n14357) );
  AOI211_X1 U16138 ( .C1(n14359), .C2(n14768), .A(n14358), .B(n14357), .ZN(
        n14375) );
  INV_X1 U16139 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n14360) );
  AOI22_X1 U16140 ( .A1(n6470), .A2(n14375), .B1(n14360), .B2(n14808), .ZN(
        P2_U3514) );
  OAI21_X1 U16141 ( .B1(n14362), .B2(n14774), .A(n14361), .ZN(n14365) );
  INV_X1 U16142 ( .A(n14363), .ZN(n14364) );
  AOI211_X1 U16143 ( .C1(n14366), .C2(n14768), .A(n14365), .B(n14364), .ZN(
        n14377) );
  AOI22_X1 U16144 ( .A1(n6470), .A2(n14377), .B1(n10002), .B2(n14808), .ZN(
        P2_U3513) );
  OAI21_X1 U16145 ( .B1(n14368), .B2(n14774), .A(n14367), .ZN(n14369) );
  AOI21_X1 U16146 ( .B1(n14370), .B2(n14768), .A(n14369), .ZN(n14371) );
  AND2_X1 U16147 ( .A1(n14372), .A2(n14371), .ZN(n14379) );
  AOI22_X1 U16148 ( .A1(n6470), .A2(n14379), .B1(n14373), .B2(n14808), .ZN(
        P2_U3511) );
  INV_X1 U16149 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n14374) );
  AOI22_X1 U16150 ( .A1(n14797), .A2(n14375), .B1(n14374), .B2(n14795), .ZN(
        P2_U3475) );
  INV_X1 U16151 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n14376) );
  AOI22_X1 U16152 ( .A1(n14797), .A2(n14377), .B1(n14376), .B2(n14795), .ZN(
        P2_U3472) );
  INV_X1 U16153 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n14378) );
  AOI22_X1 U16154 ( .A1(n14797), .A2(n14379), .B1(n14378), .B2(n14795), .ZN(
        P2_U3466) );
  AOI21_X1 U16155 ( .B1(n14397), .B2(n14381), .A(n14380), .ZN(n14428) );
  NAND2_X1 U16156 ( .A1(n14382), .A2(n14391), .ZN(n14423) );
  AND3_X1 U16157 ( .A1(n7474), .A2(n14383), .A3(n14423), .ZN(n14384) );
  AOI21_X1 U16158 ( .B1(n14428), .B2(n14519), .A(n14384), .ZN(n14400) );
  NAND2_X1 U16159 ( .A1(n14385), .A2(n14524), .ZN(n14425) );
  NOR2_X1 U16160 ( .A1(n14532), .A2(n14386), .ZN(n14387) );
  AOI21_X1 U16161 ( .B1(n14388), .B2(P1_REG2_REG_14__SCAN_IN), .A(n14387), 
        .ZN(n14389) );
  OAI21_X1 U16162 ( .B1(n14531), .B2(n14425), .A(n14389), .ZN(n14396) );
  XOR2_X1 U16163 ( .A(n14391), .B(n14390), .Z(n14393) );
  NAND2_X1 U16164 ( .A1(n14393), .A2(n14392), .ZN(n14430) );
  NAND2_X1 U16165 ( .A1(n14394), .A2(n14527), .ZN(n14424) );
  AOI21_X1 U16166 ( .B1(n14430), .B2(n14424), .A(n14531), .ZN(n14395) );
  AOI211_X1 U16167 ( .C1(n14398), .C2(n14397), .A(n14396), .B(n14395), .ZN(
        n14399) );
  NAND2_X1 U16168 ( .A1(n14400), .A2(n14399), .ZN(P1_U3279) );
  OAI22_X1 U16169 ( .A1(n14402), .A2(n14596), .B1(n14401), .B2(n14606), .ZN(
        n14403) );
  AOI21_X1 U16170 ( .B1(n14404), .B2(n14599), .A(n14403), .ZN(n14405) );
  AND2_X1 U16171 ( .A1(n14406), .A2(n14405), .ZN(n14448) );
  INV_X1 U16172 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n14407) );
  AOI22_X1 U16173 ( .A1(n14630), .A2(n14448), .B1(n14407), .B2(n14627), .ZN(
        P1_U3546) );
  AOI21_X1 U16174 ( .B1(n14409), .B2(n14580), .A(n14408), .ZN(n14413) );
  NAND3_X1 U16175 ( .A1(n14411), .A2(n14581), .A3(n14410), .ZN(n14412) );
  OAI211_X1 U16176 ( .C1(n14414), .C2(n14542), .A(n14413), .B(n14412), .ZN(
        n14415) );
  AOI21_X1 U16177 ( .B1(n14416), .B2(n14609), .A(n14415), .ZN(n14450) );
  AOI22_X1 U16178 ( .A1(n14630), .A2(n14450), .B1(n14417), .B2(n14627), .ZN(
        P1_U3544) );
  OAI22_X1 U16179 ( .A1(n14419), .A2(n14596), .B1(n14418), .B2(n14606), .ZN(
        n14420) );
  AOI211_X1 U16180 ( .C1(n14422), .C2(n14609), .A(n14421), .B(n14420), .ZN(
        n14452) );
  AOI22_X1 U16181 ( .A1(n14630), .A2(n14452), .B1(n10980), .B2(n14627), .ZN(
        P1_U3543) );
  NAND3_X1 U16182 ( .A1(n7474), .A2(n14423), .A3(n14609), .ZN(n14431) );
  OAI211_X1 U16183 ( .C1(n14426), .C2(n14606), .A(n14425), .B(n14424), .ZN(
        n14427) );
  AOI21_X1 U16184 ( .B1(n14428), .B2(n14581), .A(n14427), .ZN(n14429) );
  AOI22_X1 U16185 ( .A1(n14630), .A2(n14453), .B1(n10773), .B2(n14627), .ZN(
        P1_U3542) );
  NAND2_X1 U16186 ( .A1(n14432), .A2(n14580), .ZN(n14433) );
  OAI211_X1 U16187 ( .C1(n14435), .C2(n14596), .A(n14434), .B(n14433), .ZN(
        n14438) );
  NOR2_X1 U16188 ( .A1(n14436), .A2(n14542), .ZN(n14437) );
  AOI211_X1 U16189 ( .C1(n14439), .C2(n14609), .A(n14438), .B(n14437), .ZN(
        n14455) );
  AOI22_X1 U16190 ( .A1(n14630), .A2(n14455), .B1(n14440), .B2(n14627), .ZN(
        P1_U3541) );
  OAI22_X1 U16191 ( .A1(n14442), .A2(n14596), .B1(n14441), .B2(n14606), .ZN(
        n14444) );
  AOI211_X1 U16192 ( .C1(n14445), .C2(n14609), .A(n14444), .B(n14443), .ZN(
        n14456) );
  AOI22_X1 U16193 ( .A1(n14630), .A2(n14456), .B1(n14446), .B2(n14627), .ZN(
        P1_U3539) );
  INV_X1 U16194 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n14447) );
  AOI22_X1 U16195 ( .A1(n14613), .A2(n14448), .B1(n14447), .B2(n14611), .ZN(
        P1_U3513) );
  INV_X1 U16196 ( .A(P1_REG0_REG_16__SCAN_IN), .ZN(n14449) );
  AOI22_X1 U16197 ( .A1(n14613), .A2(n14450), .B1(n14449), .B2(n14611), .ZN(
        P1_U3507) );
  INV_X1 U16198 ( .A(P1_REG0_REG_15__SCAN_IN), .ZN(n14451) );
  AOI22_X1 U16199 ( .A1(n14613), .A2(n14452), .B1(n14451), .B2(n14611), .ZN(
        P1_U3504) );
  AOI22_X1 U16200 ( .A1(n14613), .A2(n14453), .B1(n10777), .B2(n14611), .ZN(
        P1_U3501) );
  INV_X1 U16201 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n14454) );
  AOI22_X1 U16202 ( .A1(n14613), .A2(n14455), .B1(n14454), .B2(n14611), .ZN(
        P1_U3498) );
  AOI22_X1 U16203 ( .A1(n14613), .A2(n14456), .B1(n10463), .B2(n14611), .ZN(
        P1_U3492) );
  AOI21_X1 U16204 ( .B1(n14459), .B2(n14458), .A(n14457), .ZN(n14460) );
  XOR2_X1 U16205 ( .A(n14460), .B(P2_ADDR_REG_11__SCAN_IN), .Z(SUB_1596_U69)
         );
  XNOR2_X1 U16206 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(n14461), .ZN(SUB_1596_U68)
         );
  OAI21_X1 U16207 ( .B1(n14464), .B2(n14463), .A(n14462), .ZN(n14466) );
  XOR2_X1 U16208 ( .A(n14466), .B(n14465), .Z(SUB_1596_U67) );
  AOI21_X1 U16209 ( .B1(n14469), .B2(n14468), .A(n14467), .ZN(n14470) );
  XOR2_X1 U16210 ( .A(n14470), .B(P2_ADDR_REG_14__SCAN_IN), .Z(SUB_1596_U66)
         );
  AOI21_X1 U16211 ( .B1(n14473), .B2(n14472), .A(n14471), .ZN(n14474) );
  XOR2_X1 U16212 ( .A(n14474), .B(P2_ADDR_REG_15__SCAN_IN), .Z(SUB_1596_U65)
         );
  OAI21_X1 U16213 ( .B1(n14477), .B2(n14476), .A(n14475), .ZN(n14479) );
  XOR2_X1 U16214 ( .A(n14479), .B(n14478), .Z(SUB_1596_U64) );
  INV_X1 U16215 ( .A(n14480), .ZN(n14485) );
  NAND3_X1 U16216 ( .A1(n14483), .A2(n14482), .A3(n14481), .ZN(n14484) );
  NAND2_X1 U16217 ( .A1(n14485), .A2(n14484), .ZN(n14492) );
  OAI21_X1 U16218 ( .B1(n14488), .B2(n14487), .A(n14486), .ZN(n14489) );
  AOI222_X1 U16219 ( .A1(n14492), .A2(n14504), .B1(n14491), .B2(n14490), .C1(
        n14489), .C2(n14508), .ZN(n14494) );
  OAI211_X1 U16220 ( .C1(n14496), .C2(n14495), .A(n14494), .B(n14493), .ZN(
        P1_U3255) );
  NAND2_X1 U16221 ( .A1(n14497), .A2(P1_ADDR_REG_13__SCAN_IN), .ZN(n14498) );
  OAI211_X1 U16222 ( .C1(n14501), .C2(n14500), .A(n14499), .B(n14498), .ZN(
        n14502) );
  INV_X1 U16223 ( .A(n14502), .ZN(n14513) );
  OAI211_X1 U16224 ( .C1(n14506), .C2(n14505), .A(n14504), .B(n14503), .ZN(
        n14512) );
  OAI211_X1 U16225 ( .C1(n14510), .C2(n14509), .A(n14508), .B(n14507), .ZN(
        n14511) );
  NAND3_X1 U16226 ( .A1(n14513), .A2(n14512), .A3(n14511), .ZN(P1_U3256) );
  OAI21_X1 U16227 ( .B1(n11575), .B2(n14515), .A(n14514), .ZN(n14554) );
  OR2_X1 U16228 ( .A1(n14546), .A2(n14550), .ZN(n14516) );
  NAND2_X1 U16229 ( .A1(n14517), .A2(n14516), .ZN(n14551) );
  INV_X1 U16230 ( .A(n14551), .ZN(n14518) );
  AOI22_X1 U16231 ( .A1(n14520), .A2(n14554), .B1(n14519), .B2(n14518), .ZN(
        n14538) );
  XOR2_X1 U16232 ( .A(n14551), .B(n6479), .Z(n14522) );
  MUX2_X1 U16233 ( .A(n14522), .B(n14521), .S(n14526), .Z(n14530) );
  NAND2_X1 U16234 ( .A1(n14554), .A2(n14523), .ZN(n14529) );
  AOI22_X1 U16235 ( .A1(n14527), .A2(n14526), .B1(n14525), .B2(n14524), .ZN(
        n14528) );
  OAI211_X1 U16236 ( .C1(n14530), .C2(n14542), .A(n14529), .B(n14528), .ZN(
        n14552) );
  MUX2_X1 U16237 ( .A(n14552), .B(P1_REG2_REG_1__SCAN_IN), .S(n14531), .Z(
        n14536) );
  OAI22_X1 U16238 ( .A1(n14534), .A2(n14550), .B1(n14533), .B2(n14532), .ZN(
        n14535) );
  NOR2_X1 U16239 ( .A1(n14536), .A2(n14535), .ZN(n14537) );
  NAND2_X1 U16240 ( .A1(n14538), .A2(n14537), .ZN(P1_U3292) );
  AND2_X1 U16241 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n14539), .ZN(P1_U3294) );
  AND2_X1 U16242 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n14539), .ZN(P1_U3295) );
  AND2_X1 U16243 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n14539), .ZN(P1_U3296) );
  AND2_X1 U16244 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n14539), .ZN(P1_U3297) );
  AND2_X1 U16245 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n14539), .ZN(P1_U3298) );
  AND2_X1 U16246 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n14539), .ZN(P1_U3299) );
  AND2_X1 U16247 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n14539), .ZN(P1_U3300) );
  AND2_X1 U16248 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n14539), .ZN(P1_U3301) );
  AND2_X1 U16249 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n14539), .ZN(P1_U3302) );
  AND2_X1 U16250 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n14539), .ZN(P1_U3303) );
  AND2_X1 U16251 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n14539), .ZN(P1_U3304) );
  AND2_X1 U16252 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n14539), .ZN(P1_U3305) );
  AND2_X1 U16253 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n14539), .ZN(P1_U3306) );
  AND2_X1 U16254 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n14539), .ZN(P1_U3307) );
  AND2_X1 U16255 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n14539), .ZN(P1_U3308) );
  AND2_X1 U16256 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n14539), .ZN(P1_U3309) );
  AND2_X1 U16257 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n14539), .ZN(P1_U3310) );
  AND2_X1 U16258 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n14539), .ZN(P1_U3311) );
  AND2_X1 U16259 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n14539), .ZN(P1_U3312) );
  AND2_X1 U16260 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n14539), .ZN(P1_U3313) );
  AND2_X1 U16261 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n14539), .ZN(P1_U3314) );
  AND2_X1 U16262 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n14539), .ZN(P1_U3315) );
  AND2_X1 U16263 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n14539), .ZN(P1_U3316) );
  AND2_X1 U16264 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n14539), .ZN(P1_U3317) );
  AND2_X1 U16265 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n14539), .ZN(P1_U3318) );
  AND2_X1 U16266 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n14539), .ZN(P1_U3319) );
  AND2_X1 U16267 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n14539), .ZN(P1_U3320) );
  AND2_X1 U16268 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n14539), .ZN(P1_U3321) );
  AND2_X1 U16269 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n14539), .ZN(P1_U3322) );
  AND2_X1 U16270 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n14539), .ZN(P1_U3323) );
  AOI21_X1 U16271 ( .B1(n14542), .B2(n14541), .A(n14540), .ZN(n14549) );
  INV_X1 U16272 ( .A(n14543), .ZN(n14548) );
  NOR3_X1 U16273 ( .A1(n14546), .A2(n14545), .A3(n14544), .ZN(n14547) );
  NOR3_X1 U16274 ( .A1(n14549), .A2(n14548), .A3(n14547), .ZN(n14614) );
  AOI22_X1 U16275 ( .A1(n14613), .A2(n14614), .B1(n9286), .B2(n14611), .ZN(
        P1_U3459) );
  OAI22_X1 U16276 ( .A1(n14551), .A2(n14596), .B1(n14550), .B2(n14606), .ZN(
        n14553) );
  AOI211_X1 U16277 ( .C1(n14599), .C2(n14554), .A(n14553), .B(n14552), .ZN(
        n14615) );
  AOI22_X1 U16278 ( .A1(n14613), .A2(n14615), .B1(n7312), .B2(n14611), .ZN(
        P1_U3462) );
  OAI22_X1 U16279 ( .A1(n14556), .A2(n14596), .B1(n14555), .B2(n14606), .ZN(
        n14558) );
  AOI211_X1 U16280 ( .C1(n14599), .C2(n14559), .A(n14558), .B(n14557), .ZN(
        n14616) );
  AOI22_X1 U16281 ( .A1(n14613), .A2(n14616), .B1(n9563), .B2(n14611), .ZN(
        P1_U3465) );
  INV_X1 U16282 ( .A(n14560), .ZN(n14565) );
  OAI22_X1 U16283 ( .A1(n14562), .A2(n14596), .B1(n14561), .B2(n14606), .ZN(
        n14563) );
  AOI211_X1 U16284 ( .C1(n14565), .C2(n14609), .A(n14564), .B(n14563), .ZN(
        n14618) );
  INV_X1 U16285 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n14566) );
  AOI22_X1 U16286 ( .A1(n14613), .A2(n14618), .B1(n14566), .B2(n14611), .ZN(
        P1_U3471) );
  OAI22_X1 U16287 ( .A1(n14567), .A2(n14596), .B1(n6874), .B2(n14606), .ZN(
        n14568) );
  AOI21_X1 U16288 ( .B1(n14569), .B2(n14599), .A(n14568), .ZN(n14570) );
  AND2_X1 U16289 ( .A1(n14571), .A2(n14570), .ZN(n14620) );
  INV_X1 U16290 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n14572) );
  AOI22_X1 U16291 ( .A1(n14613), .A2(n14620), .B1(n14572), .B2(n14611), .ZN(
        P1_U3474) );
  OAI22_X1 U16292 ( .A1(n14574), .A2(n14596), .B1(n14573), .B2(n14606), .ZN(
        n14577) );
  INV_X1 U16293 ( .A(n14575), .ZN(n14576) );
  AOI211_X1 U16294 ( .C1(n14599), .C2(n14578), .A(n14577), .B(n14576), .ZN(
        n14622) );
  AOI22_X1 U16295 ( .A1(n14613), .A2(n14622), .B1(n9854), .B2(n14611), .ZN(
        P1_U3477) );
  AOI22_X1 U16296 ( .A1(n14582), .A2(n14581), .B1(n14580), .B2(n14579), .ZN(
        n14583) );
  OAI211_X1 U16297 ( .C1(n14586), .C2(n14585), .A(n14584), .B(n14583), .ZN(
        n14587) );
  INV_X1 U16298 ( .A(n14587), .ZN(n14623) );
  INV_X1 U16299 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n14588) );
  AOI22_X1 U16300 ( .A1(n14613), .A2(n14623), .B1(n14588), .B2(n14611), .ZN(
        P1_U3480) );
  OAI22_X1 U16301 ( .A1(n14590), .A2(n14596), .B1(n14589), .B2(n14606), .ZN(
        n14592) );
  AOI211_X1 U16302 ( .C1(n14593), .C2(n14609), .A(n14592), .B(n14591), .ZN(
        n14624) );
  INV_X1 U16303 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n14594) );
  AOI22_X1 U16304 ( .A1(n14613), .A2(n14624), .B1(n14594), .B2(n14611), .ZN(
        P1_U3483) );
  OAI22_X1 U16305 ( .A1(n14597), .A2(n14596), .B1(n14595), .B2(n14606), .ZN(
        n14598) );
  AOI21_X1 U16306 ( .B1(n14600), .B2(n14599), .A(n14598), .ZN(n14601) );
  AND2_X1 U16307 ( .A1(n14602), .A2(n14601), .ZN(n14626) );
  INV_X1 U16308 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n14603) );
  AOI22_X1 U16309 ( .A1(n14613), .A2(n14626), .B1(n14603), .B2(n14611), .ZN(
        P1_U3486) );
  OAI211_X1 U16310 ( .C1(n14607), .C2(n14606), .A(n14605), .B(n14604), .ZN(
        n14608) );
  AOI21_X1 U16311 ( .B1(n14610), .B2(n14609), .A(n14608), .ZN(n14629) );
  INV_X1 U16312 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n14612) );
  AOI22_X1 U16313 ( .A1(n14613), .A2(n14629), .B1(n14612), .B2(n14611), .ZN(
        P1_U3489) );
  AOI22_X1 U16314 ( .A1(n14630), .A2(n14614), .B1(n9287), .B2(n14627), .ZN(
        P1_U3528) );
  AOI22_X1 U16315 ( .A1(n14630), .A2(n14615), .B1(n9303), .B2(n14627), .ZN(
        P1_U3529) );
  AOI22_X1 U16316 ( .A1(n14630), .A2(n14616), .B1(n9564), .B2(n14627), .ZN(
        P1_U3530) );
  AOI22_X1 U16317 ( .A1(n14630), .A2(n14618), .B1(n14617), .B2(n14627), .ZN(
        P1_U3532) );
  AOI22_X1 U16318 ( .A1(n14630), .A2(n14620), .B1(n14619), .B2(n14627), .ZN(
        P1_U3533) );
  AOI22_X1 U16319 ( .A1(n14630), .A2(n14622), .B1(n14621), .B2(n14627), .ZN(
        P1_U3534) );
  AOI22_X1 U16320 ( .A1(n14630), .A2(n14623), .B1(n9871), .B2(n14627), .ZN(
        P1_U3535) );
  AOI22_X1 U16321 ( .A1(n14630), .A2(n14624), .B1(n10178), .B2(n14627), .ZN(
        P1_U3536) );
  AOI22_X1 U16322 ( .A1(n14630), .A2(n14626), .B1(n14625), .B2(n14627), .ZN(
        P1_U3537) );
  AOI22_X1 U16323 ( .A1(n14630), .A2(n14629), .B1(n14628), .B2(n14627), .ZN(
        P1_U3538) );
  NOR2_X1 U16324 ( .A1(n14685), .A2(n6471), .ZN(P2_U3087) );
  NAND2_X1 U16325 ( .A1(n14686), .A2(n14798), .ZN(n14633) );
  NAND2_X1 U16326 ( .A1(n14692), .A2(n14631), .ZN(n14632) );
  AND4_X1 U16327 ( .A1(n14633), .A2(n14632), .A3(P2_IR_REG_0__SCAN_IN), .A4(
        n14667), .ZN(n14637) );
  OAI22_X1 U16328 ( .A1(n14677), .A2(n14631), .B1(n14798), .B2(n14639), .ZN(
        n14634) );
  NOR2_X1 U16329 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(n14634), .ZN(n14636) );
  OAI222_X1 U16330 ( .A1(n15247), .A2(n14671), .B1(n14637), .B2(n14636), .C1(
        n14635), .C2(P2_STATE_REG_SCAN_IN), .ZN(P2_U3214) );
  AOI22_X1 U16331 ( .A1(n14685), .A2(P2_ADDR_REG_4__SCAN_IN), .B1(n14691), 
        .B2(n14638), .ZN(n14651) );
  AOI211_X1 U16332 ( .C1(n14642), .C2(n14641), .A(n14640), .B(n14639), .ZN(
        n14643) );
  INV_X1 U16333 ( .A(n14643), .ZN(n14649) );
  AOI211_X1 U16334 ( .C1(n14646), .C2(n14645), .A(n14644), .B(n14677), .ZN(
        n14647) );
  INV_X1 U16335 ( .A(n14647), .ZN(n14648) );
  NAND4_X1 U16336 ( .A1(n14651), .A2(n14650), .A3(n14649), .A4(n14648), .ZN(
        P2_U3218) );
  AOI22_X1 U16337 ( .A1(n14685), .A2(P2_ADDR_REG_5__SCAN_IN), .B1(n14691), 
        .B2(n14652), .ZN(n14664) );
  NAND2_X1 U16338 ( .A1(n14654), .A2(n14653), .ZN(n14655) );
  NAND3_X1 U16339 ( .A1(n14686), .A2(n14656), .A3(n14655), .ZN(n14662) );
  NAND2_X1 U16340 ( .A1(n14658), .A2(n14657), .ZN(n14659) );
  NAND3_X1 U16341 ( .A1(n14660), .A2(n14692), .A3(n14659), .ZN(n14661) );
  NAND4_X1 U16342 ( .A1(n14664), .A2(n14663), .A3(n14662), .A4(n14661), .ZN(
        P2_U3219) );
  INV_X1 U16343 ( .A(P2_ADDR_REG_10__SCAN_IN), .ZN(n14670) );
  INV_X1 U16344 ( .A(n14665), .ZN(n14669) );
  OR2_X1 U16345 ( .A1(n14667), .A2(n14666), .ZN(n14668) );
  OAI211_X1 U16346 ( .C1(n14671), .C2(n14670), .A(n14669), .B(n14668), .ZN(
        n14672) );
  INV_X1 U16347 ( .A(n14672), .ZN(n14683) );
  OAI211_X1 U16348 ( .C1(n14675), .C2(n14674), .A(n14673), .B(n14686), .ZN(
        n14682) );
  AOI211_X1 U16349 ( .C1(n14679), .C2(n14678), .A(n14677), .B(n14676), .ZN(
        n14680) );
  INV_X1 U16350 ( .A(n14680), .ZN(n14681) );
  NAND3_X1 U16351 ( .A1(n14683), .A2(n14682), .A3(n14681), .ZN(P2_U3224) );
  AOI22_X1 U16352 ( .A1(n14685), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3088), .ZN(n14699) );
  OAI211_X1 U16353 ( .C1(n14689), .C2(n14688), .A(n14687), .B(n14686), .ZN(
        n14698) );
  NAND2_X1 U16354 ( .A1(n14691), .A2(n14690), .ZN(n14697) );
  OAI211_X1 U16355 ( .C1(n14695), .C2(n14694), .A(n14693), .B(n14692), .ZN(
        n14696) );
  NAND4_X1 U16356 ( .A1(n14699), .A2(n14698), .A3(n14697), .A4(n14696), .ZN(
        P2_U3227) );
  XNOR2_X1 U16357 ( .A(n14701), .B(n14700), .ZN(n14704) );
  INV_X1 U16358 ( .A(n14702), .ZN(n14703) );
  AOI21_X1 U16359 ( .B1(n14704), .B2(n14740), .A(n14703), .ZN(n14765) );
  NOR2_X1 U16360 ( .A1(n14706), .A2(n14705), .ZN(n14707) );
  AOI21_X1 U16361 ( .B1(n14708), .B2(P2_REG2_REG_4__SCAN_IN), .A(n14707), .ZN(
        n14709) );
  OAI21_X1 U16362 ( .B1(n14721), .B2(n14764), .A(n14709), .ZN(n14710) );
  INV_X1 U16363 ( .A(n14710), .ZN(n14718) );
  XNOR2_X1 U16364 ( .A(n14712), .B(n14711), .ZN(n14769) );
  OAI211_X1 U16365 ( .C1(n14715), .C2(n14764), .A(n14714), .B(n14713), .ZN(
        n14763) );
  INV_X1 U16366 ( .A(n14763), .ZN(n14716) );
  AOI22_X1 U16367 ( .A1(n14769), .A2(n14727), .B1(n14725), .B2(n14716), .ZN(
        n14717) );
  OAI211_X1 U16368 ( .C1(n14731), .C2(n14765), .A(n14718), .B(n14717), .ZN(
        P2_U3261) );
  AOI22_X1 U16369 ( .A1(n14708), .A2(P2_REG2_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(n14719), .ZN(n14720) );
  OAI21_X1 U16370 ( .B1(n14721), .B2(n9024), .A(n14720), .ZN(n14722) );
  INV_X1 U16371 ( .A(n14722), .ZN(n14729) );
  INV_X1 U16372 ( .A(n14723), .ZN(n14724) );
  AOI22_X1 U16373 ( .A1(n14727), .A2(n14726), .B1(n14725), .B2(n14724), .ZN(
        n14728) );
  OAI211_X1 U16374 ( .C1(n14731), .C2(n14730), .A(n14729), .B(n14728), .ZN(
        P2_U3263) );
  AND2_X1 U16375 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n14733), .ZN(P2_U3266) );
  AND2_X1 U16376 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n14733), .ZN(P2_U3267) );
  AND2_X1 U16377 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n14733), .ZN(P2_U3268) );
  AND2_X1 U16378 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n14733), .ZN(P2_U3269) );
  AND2_X1 U16379 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n14733), .ZN(P2_U3270) );
  AND2_X1 U16380 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n14733), .ZN(P2_U3271) );
  AND2_X1 U16381 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n14733), .ZN(P2_U3272) );
  AND2_X1 U16382 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n14733), .ZN(P2_U3273) );
  AND2_X1 U16383 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n14733), .ZN(P2_U3274) );
  AND2_X1 U16384 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n14733), .ZN(P2_U3275) );
  AND2_X1 U16385 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n14733), .ZN(P2_U3276) );
  AND2_X1 U16386 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n14733), .ZN(P2_U3277) );
  AND2_X1 U16387 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n14733), .ZN(P2_U3278) );
  AND2_X1 U16388 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n14733), .ZN(P2_U3279) );
  AND2_X1 U16389 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n14733), .ZN(P2_U3280) );
  AND2_X1 U16390 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n14733), .ZN(P2_U3281) );
  AND2_X1 U16391 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n14733), .ZN(P2_U3282) );
  AND2_X1 U16392 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n14733), .ZN(P2_U3283) );
  AND2_X1 U16393 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n14733), .ZN(P2_U3284) );
  AND2_X1 U16394 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n14733), .ZN(P2_U3285) );
  AND2_X1 U16395 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n14733), .ZN(P2_U3286) );
  AND2_X1 U16396 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n14733), .ZN(P2_U3287) );
  AND2_X1 U16397 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n14733), .ZN(P2_U3288) );
  AND2_X1 U16398 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n14733), .ZN(P2_U3289) );
  AND2_X1 U16399 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n14733), .ZN(P2_U3290) );
  AND2_X1 U16400 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n14733), .ZN(P2_U3291) );
  AND2_X1 U16401 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n14733), .ZN(P2_U3292) );
  AND2_X1 U16402 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n14733), .ZN(P2_U3293) );
  AND2_X1 U16403 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n14733), .ZN(P2_U3294) );
  AND2_X1 U16404 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n14733), .ZN(P2_U3295) );
  AOI22_X1 U16405 ( .A1(n14736), .A2(n14735), .B1(n14734), .B2(n14738), .ZN(
        P2_U3416) );
  AOI21_X1 U16406 ( .B1(n14739), .B2(n14738), .A(n14737), .ZN(P2_U3417) );
  OAI21_X1 U16407 ( .B1(n14741), .B2(n14740), .A(n14748), .ZN(n14746) );
  NAND3_X1 U16408 ( .A1(n14743), .A2(n12720), .A3(n14742), .ZN(n14744) );
  NAND3_X1 U16409 ( .A1(n14746), .A2(n14745), .A3(n14744), .ZN(n14747) );
  AOI21_X1 U16410 ( .B1(n14761), .B2(n14748), .A(n14747), .ZN(n14799) );
  INV_X1 U16411 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n14749) );
  AOI22_X1 U16412 ( .A1(n14797), .A2(n14799), .B1(n14749), .B2(n14795), .ZN(
        P2_U3430) );
  INV_X1 U16413 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n14750) );
  AOI22_X1 U16414 ( .A1(n14797), .A2(n14751), .B1(n14750), .B2(n14795), .ZN(
        P2_U3433) );
  INV_X1 U16415 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n14752) );
  AOI22_X1 U16416 ( .A1(n14797), .A2(n14753), .B1(n14752), .B2(n14795), .ZN(
        P2_U3436) );
  INV_X1 U16417 ( .A(n14757), .ZN(n14760) );
  OAI21_X1 U16418 ( .B1(n14755), .B2(n14774), .A(n14754), .ZN(n14759) );
  OAI21_X1 U16419 ( .B1(n9328), .B2(n14757), .A(n14756), .ZN(n14758) );
  AOI211_X1 U16420 ( .C1(n14761), .C2(n14760), .A(n14759), .B(n14758), .ZN(
        n14801) );
  INV_X1 U16421 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n14762) );
  AOI22_X1 U16422 ( .A1(n14797), .A2(n14801), .B1(n14762), .B2(n14795), .ZN(
        P2_U3439) );
  OAI21_X1 U16423 ( .B1(n14764), .B2(n14774), .A(n14763), .ZN(n14767) );
  INV_X1 U16424 ( .A(n14765), .ZN(n14766) );
  AOI211_X1 U16425 ( .C1(n14769), .C2(n14768), .A(n14767), .B(n14766), .ZN(
        n14803) );
  INV_X1 U16426 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n14770) );
  AOI22_X1 U16427 ( .A1(n14797), .A2(n14803), .B1(n14770), .B2(n14795), .ZN(
        P2_U3442) );
  INV_X1 U16428 ( .A(n14771), .ZN(n14772) );
  OAI211_X1 U16429 ( .C1(n14775), .C2(n14774), .A(n14773), .B(n14772), .ZN(
        n14778) );
  AOI21_X1 U16430 ( .B1(n9328), .B2(n14793), .A(n14776), .ZN(n14777) );
  NOR2_X1 U16431 ( .A1(n14778), .A2(n14777), .ZN(n14805) );
  INV_X1 U16432 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n14779) );
  AOI22_X1 U16433 ( .A1(n14797), .A2(n14805), .B1(n14779), .B2(n14795), .ZN(
        P2_U3445) );
  AOI21_X1 U16434 ( .B1(n14781), .B2(n14788), .A(n14780), .ZN(n14782) );
  OAI211_X1 U16435 ( .C1(n14793), .C2(n14784), .A(n14783), .B(n14782), .ZN(
        n14785) );
  INV_X1 U16436 ( .A(n14785), .ZN(n14807) );
  INV_X1 U16437 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n14786) );
  AOI22_X1 U16438 ( .A1(n14797), .A2(n14807), .B1(n14786), .B2(n14795), .ZN(
        P2_U3454) );
  AOI21_X1 U16439 ( .B1(n14789), .B2(n14788), .A(n14787), .ZN(n14790) );
  OAI211_X1 U16440 ( .C1(n14793), .C2(n14792), .A(n14791), .B(n14790), .ZN(
        n14794) );
  INV_X1 U16441 ( .A(n14794), .ZN(n14809) );
  INV_X1 U16442 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n14796) );
  AOI22_X1 U16443 ( .A1(n14797), .A2(n14809), .B1(n14796), .B2(n14795), .ZN(
        P2_U3460) );
  AOI22_X1 U16444 ( .A1(n6470), .A2(n14799), .B1(n14798), .B2(n14808), .ZN(
        P2_U3499) );
  AOI22_X1 U16445 ( .A1(n6470), .A2(n14801), .B1(n14800), .B2(n14808), .ZN(
        P2_U3502) );
  AOI22_X1 U16446 ( .A1(n6470), .A2(n14803), .B1(n14802), .B2(n14808), .ZN(
        P2_U3503) );
  AOI22_X1 U16447 ( .A1(n6470), .A2(n14805), .B1(n14804), .B2(n14808), .ZN(
        P2_U3504) );
  AOI22_X1 U16448 ( .A1(n6470), .A2(n14807), .B1(n14806), .B2(n14808), .ZN(
        P2_U3507) );
  AOI22_X1 U16449 ( .A1(n6470), .A2(n14809), .B1(n9081), .B2(n14808), .ZN(
        P2_U3509) );
  NOR2_X1 U16450 ( .A1(P3_U3897), .A2(n14869), .ZN(P3_U3150) );
  AOI22_X1 U16451 ( .A1(n14846), .A2(P3_IR_REG_0__SCAN_IN), .B1(n14869), .B2(
        P3_ADDR_REG_0__SCAN_IN), .ZN(n14815) );
  NOR2_X1 U16452 ( .A1(n14810), .A2(P3_IR_REG_0__SCAN_IN), .ZN(n14812) );
  NAND3_X1 U16453 ( .A1(n14893), .A2(n14887), .A3(n14885), .ZN(n14811) );
  OAI21_X1 U16454 ( .B1(n14813), .B2(n14812), .A(n14811), .ZN(n14814) );
  OAI211_X1 U16455 ( .C1(P3_STATE_REG_SCAN_IN), .C2(n9524), .A(n14815), .B(
        n14814), .ZN(P3_U3182) );
  AOI21_X1 U16456 ( .B1(n6616), .B2(n14817), .A(n14816), .ZN(n14829) );
  AOI21_X1 U16457 ( .B1(n14820), .B2(n14819), .A(n14818), .ZN(n14821) );
  OR2_X1 U16458 ( .A1(n14821), .A2(n14893), .ZN(n14828) );
  OAI21_X1 U16459 ( .B1(n14824), .B2(n14823), .A(n14822), .ZN(n14825) );
  AOI22_X1 U16460 ( .A1(n14826), .A2(n14846), .B1(n14825), .B2(n14843), .ZN(
        n14827) );
  OAI211_X1 U16461 ( .C1(n14829), .C2(n14887), .A(n14828), .B(n14827), .ZN(
        n14830) );
  INV_X1 U16462 ( .A(n14830), .ZN(n14832) );
  NAND2_X1 U16463 ( .A1(P3_REG3_REG_6__SCAN_IN), .A2(P3_U3151), .ZN(n14831) );
  OAI211_X1 U16464 ( .C1(n14833), .C2(n14875), .A(n14832), .B(n14831), .ZN(
        P3_U3188) );
  AOI21_X1 U16465 ( .B1(n14836), .B2(n14835), .A(n14834), .ZN(n14849) );
  AOI21_X1 U16466 ( .B1(n14839), .B2(n14838), .A(n14837), .ZN(n14840) );
  OR2_X1 U16467 ( .A1(n14840), .A2(n14893), .ZN(n14848) );
  XNOR2_X1 U16468 ( .A(n14842), .B(n14841), .ZN(n14844) );
  AOI22_X1 U16469 ( .A1(n14846), .A2(n14845), .B1(n14844), .B2(n14843), .ZN(
        n14847) );
  OAI211_X1 U16470 ( .C1(n14849), .C2(n14887), .A(n14848), .B(n14847), .ZN(
        n14850) );
  INV_X1 U16471 ( .A(n14850), .ZN(n14852) );
  NAND2_X1 U16472 ( .A1(P3_REG3_REG_8__SCAN_IN), .A2(P3_U3151), .ZN(n14851) );
  OAI211_X1 U16473 ( .C1(n14853), .C2(n14875), .A(n14852), .B(n14851), .ZN(
        P3_U3190) );
  AOI21_X1 U16474 ( .B1(n14856), .B2(n14855), .A(n14854), .ZN(n14871) );
  AOI21_X1 U16475 ( .B1(n14859), .B2(n14858), .A(n14857), .ZN(n14861) );
  OAI21_X1 U16476 ( .B1(n14861), .B2(n14887), .A(n14860), .ZN(n14868) );
  AOI21_X1 U16477 ( .B1(n14864), .B2(n14863), .A(n14862), .ZN(n14865) );
  OAI22_X1 U16478 ( .A1(n14878), .A2(n14866), .B1(n14865), .B2(n14885), .ZN(
        n14867) );
  AOI211_X1 U16479 ( .C1(n14869), .C2(P3_ADDR_REG_10__SCAN_IN), .A(n14868), 
        .B(n14867), .ZN(n14870) );
  OAI21_X1 U16480 ( .B1(n14871), .B2(n14893), .A(n14870), .ZN(P3_U3192) );
  AOI21_X1 U16481 ( .B1(n14874), .B2(n14873), .A(n14872), .ZN(n14894) );
  OAI22_X1 U16482 ( .A1(n14878), .A2(n14877), .B1(n14876), .B2(n14875), .ZN(
        n14890) );
  AOI21_X1 U16483 ( .B1(n14881), .B2(n14880), .A(n14879), .ZN(n14888) );
  AOI21_X1 U16484 ( .B1(n14884), .B2(n14883), .A(n14882), .ZN(n14886) );
  OAI22_X1 U16485 ( .A1(n14888), .A2(n14887), .B1(n14886), .B2(n14885), .ZN(
        n14889) );
  NOR3_X1 U16486 ( .A1(n14891), .A2(n14890), .A3(n14889), .ZN(n14892) );
  OAI21_X1 U16487 ( .B1(n14894), .B2(n14893), .A(n14892), .ZN(P3_U3193) );
  INV_X1 U16488 ( .A(n14895), .ZN(n14953) );
  XOR2_X1 U16489 ( .A(n14896), .B(n14898), .Z(n15018) );
  INV_X1 U16490 ( .A(n15018), .ZN(n14903) );
  OAI211_X1 U16491 ( .C1(n14899), .C2(n14898), .A(n14897), .B(n14961), .ZN(
        n14900) );
  INV_X1 U16492 ( .A(n14900), .ZN(n14902) );
  AOI211_X1 U16493 ( .C1(n15018), .C2(n14968), .A(n14902), .B(n14901), .ZN(
        n15020) );
  OAI21_X1 U16494 ( .B1(n14953), .B2(n14903), .A(n15020), .ZN(n14908) );
  OAI22_X1 U16495 ( .A1(n14906), .A2(n14905), .B1(n14904), .B2(n14977), .ZN(
        n14907) );
  AOI21_X1 U16496 ( .B1(n14908), .B2(n14977), .A(n14907), .ZN(n14909) );
  OAI21_X1 U16497 ( .B1(n14910), .B2(n14959), .A(n14909), .ZN(P3_U3223) );
  OAI21_X1 U16498 ( .B1(n14913), .B2(n14912), .A(n14911), .ZN(n15002) );
  INV_X1 U16499 ( .A(n15002), .ZN(n14920) );
  OAI211_X1 U16500 ( .C1(n14916), .C2(n14915), .A(n14914), .B(n14961), .ZN(
        n14917) );
  INV_X1 U16501 ( .A(n14917), .ZN(n14918) );
  AOI211_X1 U16502 ( .C1(n15002), .C2(n14968), .A(n14919), .B(n14918), .ZN(
        n15004) );
  OAI21_X1 U16503 ( .B1(n14920), .B2(n14953), .A(n15004), .ZN(n14921) );
  MUX2_X1 U16504 ( .A(P3_REG2_REG_7__SCAN_IN), .B(n14921), .S(n14977), .Z(
        n14922) );
  AOI21_X1 U16505 ( .B1(n14957), .B2(n15001), .A(n14922), .ZN(n14923) );
  OAI21_X1 U16506 ( .B1(n14924), .B2(n14959), .A(n14923), .ZN(P3_U3226) );
  OAI21_X1 U16507 ( .B1(n14927), .B2(n14926), .A(n14925), .ZN(n14997) );
  INV_X1 U16508 ( .A(n14997), .ZN(n14934) );
  OAI211_X1 U16509 ( .C1(n14930), .C2(n14929), .A(n14928), .B(n14961), .ZN(
        n14931) );
  INV_X1 U16510 ( .A(n14931), .ZN(n14932) );
  AOI211_X1 U16511 ( .C1(n14997), .C2(n14968), .A(n14933), .B(n14932), .ZN(
        n14999) );
  OAI21_X1 U16512 ( .B1(n14934), .B2(n14953), .A(n14999), .ZN(n14935) );
  MUX2_X1 U16513 ( .A(P3_REG2_REG_6__SCAN_IN), .B(n14935), .S(n14977), .Z(
        n14936) );
  AOI21_X1 U16514 ( .B1(n14957), .B2(n14996), .A(n14936), .ZN(n14937) );
  OAI21_X1 U16515 ( .B1(n14938), .B2(n14959), .A(n14937), .ZN(P3_U3227) );
  AOI22_X1 U16516 ( .A1(n14979), .A2(P3_REG2_REG_5__SCAN_IN), .B1(n14973), 
        .B2(n14939), .ZN(n14944) );
  AOI22_X1 U16517 ( .A1(n14942), .A2(n14941), .B1(n14940), .B2(n14957), .ZN(
        n14943) );
  OAI211_X1 U16518 ( .C1(n14979), .C2(n14945), .A(n14944), .B(n14943), .ZN(
        P3_U3228) );
  OAI21_X1 U16519 ( .B1(n14947), .B2(n14950), .A(n14946), .ZN(n14992) );
  INV_X1 U16520 ( .A(n14992), .ZN(n14954) );
  AOI211_X1 U16521 ( .C1(n14950), .C2(n10275), .A(n14949), .B(n14948), .ZN(
        n14951) );
  AOI211_X1 U16522 ( .C1(n14968), .C2(n14992), .A(n14952), .B(n14951), .ZN(
        n14994) );
  OAI21_X1 U16523 ( .B1(n14954), .B2(n14953), .A(n14994), .ZN(n14955) );
  MUX2_X1 U16524 ( .A(P3_REG2_REG_3__SCAN_IN), .B(n14955), .S(n14977), .Z(
        n14956) );
  AOI21_X1 U16525 ( .B1(n14957), .B2(n14991), .A(n14956), .ZN(n14958) );
  OAI21_X1 U16526 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(n14959), .A(n14958), .ZN(
        P3_U3230) );
  XNOR2_X1 U16527 ( .A(n14966), .B(n14960), .ZN(n14962) );
  NAND2_X1 U16528 ( .A1(n14962), .A2(n14961), .ZN(n14965) );
  INV_X1 U16529 ( .A(n14963), .ZN(n14964) );
  NAND2_X1 U16530 ( .A1(n14965), .A2(n14964), .ZN(n14980) );
  INV_X1 U16531 ( .A(n14980), .ZN(n14972) );
  XNOR2_X1 U16532 ( .A(n14967), .B(n14966), .ZN(n14982) );
  NAND2_X1 U16533 ( .A1(n14982), .A2(n14968), .ZN(n14971) );
  AND2_X1 U16534 ( .A1(n9552), .A2(n15016), .ZN(n14981) );
  NAND2_X1 U16535 ( .A1(n14981), .A2(n14969), .ZN(n14970) );
  AND3_X1 U16536 ( .A1(n14972), .A2(n14971), .A3(n14970), .ZN(n14978) );
  AOI22_X1 U16537 ( .A1(n14982), .A2(n14974), .B1(P3_REG3_REG_1__SCAN_IN), 
        .B2(n14973), .ZN(n14975) );
  OAI221_X1 U16538 ( .B1(n14979), .B2(n14978), .C1(n14977), .C2(n14976), .A(
        n14975), .ZN(P3_U3232) );
  AOI211_X1 U16539 ( .C1(n14983), .C2(n14982), .A(n14981), .B(n14980), .ZN(
        n15023) );
  INV_X1 U16540 ( .A(P3_REG0_REG_1__SCAN_IN), .ZN(n14984) );
  AOI22_X1 U16541 ( .A1(n15015), .A2(n15023), .B1(n14984), .B2(n8422), .ZN(
        P3_U3393) );
  INV_X1 U16542 ( .A(n14985), .ZN(n14987) );
  OAI211_X1 U16543 ( .C1(n14989), .C2(n14988), .A(n14987), .B(n14986), .ZN(
        n15024) );
  OAI22_X1 U16544 ( .A1(n8422), .A2(n15024), .B1(P3_REG0_REG_2__SCAN_IN), .B2(
        n15015), .ZN(n14990) );
  INV_X1 U16545 ( .A(n14990), .ZN(P3_U3396) );
  AOI22_X1 U16546 ( .A1(n14992), .A2(n6604), .B1(n14991), .B2(n15016), .ZN(
        n14993) );
  AND2_X1 U16547 ( .A1(n14994), .A2(n14993), .ZN(n15027) );
  INV_X1 U16548 ( .A(P3_REG0_REG_3__SCAN_IN), .ZN(n14995) );
  AOI22_X1 U16549 ( .A1(n15015), .A2(n15027), .B1(n14995), .B2(n8422), .ZN(
        P3_U3399) );
  AOI22_X1 U16550 ( .A1(n14997), .A2(n6604), .B1(n15016), .B2(n14996), .ZN(
        n14998) );
  AND2_X1 U16551 ( .A1(n14999), .A2(n14998), .ZN(n15029) );
  INV_X1 U16552 ( .A(P3_REG0_REG_6__SCAN_IN), .ZN(n15000) );
  AOI22_X1 U16553 ( .A1(n15015), .A2(n15029), .B1(n15000), .B2(n8422), .ZN(
        P3_U3408) );
  AOI22_X1 U16554 ( .A1(n15002), .A2(n6604), .B1(n15001), .B2(n15016), .ZN(
        n15003) );
  AND2_X1 U16555 ( .A1(n15004), .A2(n15003), .ZN(n15031) );
  INV_X1 U16556 ( .A(P3_REG0_REG_7__SCAN_IN), .ZN(n15005) );
  AOI22_X1 U16557 ( .A1(n15015), .A2(n15031), .B1(n15005), .B2(n8422), .ZN(
        P3_U3411) );
  AOI21_X1 U16558 ( .B1(n15007), .B2(n6604), .A(n15006), .ZN(n15008) );
  INV_X1 U16559 ( .A(P3_REG0_REG_8__SCAN_IN), .ZN(n15010) );
  AOI22_X1 U16560 ( .A1(n15015), .A2(n15033), .B1(n15010), .B2(n8422), .ZN(
        P3_U3414) );
  AOI211_X1 U16561 ( .C1(n15013), .C2(n6604), .A(n15012), .B(n15011), .ZN(
        n15035) );
  INV_X1 U16562 ( .A(P3_REG0_REG_9__SCAN_IN), .ZN(n15014) );
  AOI22_X1 U16563 ( .A1(n15015), .A2(n15035), .B1(n15014), .B2(n8422), .ZN(
        P3_U3417) );
  AOI22_X1 U16564 ( .A1(n15018), .A2(n6604), .B1(n15017), .B2(n15016), .ZN(
        n15019) );
  AND2_X1 U16565 ( .A1(n15020), .A2(n15019), .ZN(n15037) );
  INV_X1 U16566 ( .A(P3_REG0_REG_10__SCAN_IN), .ZN(n15021) );
  AOI22_X1 U16567 ( .A1(n15015), .A2(n15037), .B1(n15021), .B2(n8422), .ZN(
        P3_U3420) );
  AOI22_X1 U16568 ( .A1(n15038), .A2(n15023), .B1(n15022), .B2(n15036), .ZN(
        P3_U3460) );
  OAI22_X1 U16569 ( .A1(n15036), .A2(n15024), .B1(P3_REG1_REG_2__SCAN_IN), 
        .B2(n15038), .ZN(n15025) );
  INV_X1 U16570 ( .A(n15025), .ZN(P3_U3461) );
  AOI22_X1 U16571 ( .A1(n15038), .A2(n15027), .B1(n15026), .B2(n15036), .ZN(
        P3_U3462) );
  INV_X1 U16572 ( .A(P3_REG1_REG_6__SCAN_IN), .ZN(n15028) );
  AOI22_X1 U16573 ( .A1(n15038), .A2(n15029), .B1(n15028), .B2(n15036), .ZN(
        P3_U3465) );
  AOI22_X1 U16574 ( .A1(n15038), .A2(n15031), .B1(n15030), .B2(n15036), .ZN(
        P3_U3466) );
  INV_X1 U16575 ( .A(P3_REG1_REG_8__SCAN_IN), .ZN(n15032) );
  AOI22_X1 U16576 ( .A1(n15038), .A2(n15033), .B1(n15032), .B2(n15036), .ZN(
        P3_U3467) );
  AOI22_X1 U16577 ( .A1(n15038), .A2(n15035), .B1(n15034), .B2(n15036), .ZN(
        P3_U3468) );
  AOI22_X1 U16578 ( .A1(n15038), .A2(n15037), .B1(n8319), .B2(n15036), .ZN(
        P3_U3469) );
  INV_X1 U16579 ( .A(P3_REG3_REG_24__SCAN_IN), .ZN(n15043) );
  AOI22_X1 U16580 ( .A1(n15043), .A2(keyinput_g51), .B1(keyinput_g16), .B2(
        n15144), .ZN(n15042) );
  OAI221_X1 U16581 ( .B1(n15043), .B2(keyinput_g51), .C1(n15144), .C2(
        keyinput_g16), .A(n15042), .ZN(n15053) );
  AOI22_X1 U16582 ( .A1(n15045), .A2(keyinput_g13), .B1(n7686), .B2(
        keyinput_g53), .ZN(n15044) );
  OAI221_X1 U16583 ( .B1(n15045), .B2(keyinput_g13), .C1(n7686), .C2(
        keyinput_g53), .A(n15044), .ZN(n15052) );
  AOI22_X1 U16584 ( .A1(n15048), .A2(keyinput_g36), .B1(keyinput_g4), .B2(
        n15047), .ZN(n15046) );
  OAI221_X1 U16585 ( .B1(n15048), .B2(keyinput_g36), .C1(n15047), .C2(
        keyinput_g4), .A(n15046), .ZN(n15051) );
  AOI22_X1 U16586 ( .A1(n9724), .A2(keyinput_g59), .B1(keyinput_g33), .B2(
        n15168), .ZN(n15049) );
  OAI221_X1 U16587 ( .B1(n9724), .B2(keyinput_g59), .C1(n15168), .C2(
        keyinput_g33), .A(n15049), .ZN(n15050) );
  NOR4_X1 U16588 ( .A1(n15053), .A2(n15052), .A3(n15051), .A4(n15050), .ZN(
        n15097) );
  AOI22_X1 U16589 ( .A1(SI_0_), .A2(keyinput_g32), .B1(SI_24_), .B2(
        keyinput_g8), .ZN(n15054) );
  OAI221_X1 U16590 ( .B1(SI_0_), .B2(keyinput_g32), .C1(SI_24_), .C2(
        keyinput_g8), .A(n15054), .ZN(n15064) );
  AOI22_X1 U16591 ( .A1(n15204), .A2(keyinput_g41), .B1(keyinput_g2), .B2(
        n15056), .ZN(n15055) );
  OAI221_X1 U16592 ( .B1(n15204), .B2(keyinput_g41), .C1(n15056), .C2(
        keyinput_g2), .A(n15055), .ZN(n15063) );
  AOI22_X1 U16593 ( .A1(P3_REG3_REG_1__SCAN_IN), .A2(keyinput_g44), .B1(
        P3_REG3_REG_4__SCAN_IN), .B2(keyinput_g52), .ZN(n15057) );
  OAI221_X1 U16594 ( .B1(P3_REG3_REG_1__SCAN_IN), .B2(keyinput_g44), .C1(
        P3_REG3_REG_4__SCAN_IN), .C2(keyinput_g52), .A(n15057), .ZN(n15062) );
  XNOR2_X1 U16595 ( .A(n15058), .B(keyinput_g43), .ZN(n15060) );
  XNOR2_X1 U16596 ( .A(SI_3_), .B(keyinput_g29), .ZN(n15059) );
  NAND2_X1 U16597 ( .A1(n15060), .A2(n15059), .ZN(n15061) );
  NOR4_X1 U16598 ( .A1(n15064), .A2(n15063), .A3(n15062), .A4(n15061), .ZN(
        n15096) );
  AOI22_X1 U16599 ( .A1(n15067), .A2(keyinput_g40), .B1(n15066), .B2(
        keyinput_g42), .ZN(n15065) );
  OAI221_X1 U16600 ( .B1(n15067), .B2(keyinput_g40), .C1(n15066), .C2(
        keyinput_g42), .A(n15065), .ZN(n15080) );
  INV_X1 U16601 ( .A(P3_REG3_REG_6__SCAN_IN), .ZN(n15070) );
  INV_X1 U16602 ( .A(P3_REG3_REG_23__SCAN_IN), .ZN(n15069) );
  AOI22_X1 U16603 ( .A1(n15070), .A2(keyinput_g61), .B1(n15069), .B2(
        keyinput_g38), .ZN(n15068) );
  OAI221_X1 U16604 ( .B1(n15070), .B2(keyinput_g61), .C1(n15069), .C2(
        keyinput_g38), .A(n15068), .ZN(n15079) );
  AOI22_X1 U16605 ( .A1(n15073), .A2(keyinput_g58), .B1(keyinput_g15), .B2(
        n15072), .ZN(n15071) );
  OAI221_X1 U16606 ( .B1(n15073), .B2(keyinput_g58), .C1(n15072), .C2(
        keyinput_g15), .A(n15071), .ZN(n15078) );
  INV_X1 U16607 ( .A(SI_31_), .ZN(n15074) );
  XOR2_X1 U16608 ( .A(n15074), .B(keyinput_g1), .Z(n15076) );
  XNOR2_X1 U16609 ( .A(SI_2_), .B(keyinput_g30), .ZN(n15075) );
  NAND2_X1 U16610 ( .A1(n15076), .A2(n15075), .ZN(n15077) );
  NOR4_X1 U16611 ( .A1(n15080), .A2(n15079), .A3(n15078), .A4(n15077), .ZN(
        n15095) );
  AOI22_X1 U16612 ( .A1(n15082), .A2(keyinput_g57), .B1(keyinput_g17), .B2(
        n15194), .ZN(n15081) );
  OAI221_X1 U16613 ( .B1(n15082), .B2(keyinput_g57), .C1(n15194), .C2(
        keyinput_g17), .A(n15081), .ZN(n15093) );
  AOI22_X1 U16614 ( .A1(n15206), .A2(keyinput_g62), .B1(keyinput_g6), .B2(
        n15084), .ZN(n15083) );
  OAI221_X1 U16615 ( .B1(n15206), .B2(keyinput_g62), .C1(n15084), .C2(
        keyinput_g6), .A(n15083), .ZN(n15092) );
  INV_X1 U16616 ( .A(P3_REG3_REG_10__SCAN_IN), .ZN(n15086) );
  AOI22_X1 U16617 ( .A1(n15176), .A2(keyinput_g35), .B1(n15086), .B2(
        keyinput_g39), .ZN(n15085) );
  OAI221_X1 U16618 ( .B1(n15176), .B2(keyinput_g35), .C1(n15086), .C2(
        keyinput_g39), .A(n15085), .ZN(n15091) );
  AOI22_X1 U16619 ( .A1(n15089), .A2(keyinput_g18), .B1(keyinput_g7), .B2(
        n15088), .ZN(n15087) );
  OAI221_X1 U16620 ( .B1(n15089), .B2(keyinput_g18), .C1(n15088), .C2(
        keyinput_g7), .A(n15087), .ZN(n15090) );
  NOR4_X1 U16621 ( .A1(n15093), .A2(n15092), .A3(n15091), .A4(n15090), .ZN(
        n15094) );
  NAND4_X1 U16622 ( .A1(n15097), .A2(n15096), .A3(n15095), .A4(n15094), .ZN(
        n15233) );
  AOI22_X1 U16623 ( .A1(SI_22_), .A2(keyinput_g10), .B1(P3_REG3_REG_5__SCAN_IN), .B2(keyinput_g49), .ZN(n15098) );
  OAI221_X1 U16624 ( .B1(SI_22_), .B2(keyinput_g10), .C1(
        P3_REG3_REG_5__SCAN_IN), .C2(keyinput_g49), .A(n15098), .ZN(n15105) );
  AOI22_X1 U16625 ( .A1(SI_9_), .A2(keyinput_g23), .B1(SI_21_), .B2(
        keyinput_g11), .ZN(n15099) );
  OAI221_X1 U16626 ( .B1(SI_9_), .B2(keyinput_g23), .C1(SI_21_), .C2(
        keyinput_g11), .A(n15099), .ZN(n15104) );
  AOI22_X1 U16627 ( .A1(SI_23_), .A2(keyinput_g9), .B1(P3_REG3_REG_21__SCAN_IN), .B2(keyinput_g45), .ZN(n15100) );
  OAI221_X1 U16628 ( .B1(SI_23_), .B2(keyinput_g9), .C1(
        P3_REG3_REG_21__SCAN_IN), .C2(keyinput_g45), .A(n15100), .ZN(n15103)
         );
  AOI22_X1 U16629 ( .A1(P3_REG3_REG_0__SCAN_IN), .A2(keyinput_g54), .B1(SI_5_), 
        .B2(keyinput_g27), .ZN(n15101) );
  OAI221_X1 U16630 ( .B1(P3_REG3_REG_0__SCAN_IN), .B2(keyinput_g54), .C1(SI_5_), .C2(keyinput_g27), .A(n15101), .ZN(n15102) );
  NOR4_X1 U16631 ( .A1(n15105), .A2(n15104), .A3(n15103), .A4(n15102), .ZN(
        n15132) );
  XNOR2_X1 U16632 ( .A(n15210), .B(keyinput_g48), .ZN(n15112) );
  AOI22_X1 U16633 ( .A1(SI_7_), .A2(keyinput_g25), .B1(SI_27_), .B2(
        keyinput_g5), .ZN(n15106) );
  OAI221_X1 U16634 ( .B1(SI_7_), .B2(keyinput_g25), .C1(SI_27_), .C2(
        keyinput_g5), .A(n15106), .ZN(n15111) );
  AOI22_X1 U16635 ( .A1(SI_18_), .A2(keyinput_g14), .B1(
        P3_REG3_REG_17__SCAN_IN), .B2(keyinput_g50), .ZN(n15107) );
  OAI221_X1 U16636 ( .B1(SI_18_), .B2(keyinput_g14), .C1(
        P3_REG3_REG_17__SCAN_IN), .C2(keyinput_g50), .A(n15107), .ZN(n15110)
         );
  AOI22_X1 U16637 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(keyinput_g46), .B1(
        P3_REG3_REG_14__SCAN_IN), .B2(keyinput_g37), .ZN(n15108) );
  OAI221_X1 U16638 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput_g46), .C1(
        P3_REG3_REG_14__SCAN_IN), .C2(keyinput_g37), .A(n15108), .ZN(n15109)
         );
  NOR4_X1 U16639 ( .A1(n15112), .A2(n15111), .A3(n15110), .A4(n15109), .ZN(
        n15131) );
  AOI22_X1 U16640 ( .A1(SI_1_), .A2(keyinput_g31), .B1(SI_11_), .B2(
        keyinput_g21), .ZN(n15113) );
  OAI221_X1 U16641 ( .B1(SI_1_), .B2(keyinput_g31), .C1(SI_11_), .C2(
        keyinput_g21), .A(n15113), .ZN(n15120) );
  AOI22_X1 U16642 ( .A1(SI_13_), .A2(keyinput_g19), .B1(
        P3_REG3_REG_13__SCAN_IN), .B2(keyinput_g56), .ZN(n15114) );
  OAI221_X1 U16643 ( .B1(SI_13_), .B2(keyinput_g19), .C1(
        P3_REG3_REG_13__SCAN_IN), .C2(keyinput_g56), .A(n15114), .ZN(n15119)
         );
  AOI22_X1 U16644 ( .A1(SI_10_), .A2(keyinput_g22), .B1(
        P3_REG3_REG_25__SCAN_IN), .B2(keyinput_g47), .ZN(n15115) );
  OAI221_X1 U16645 ( .B1(SI_10_), .B2(keyinput_g22), .C1(
        P3_REG3_REG_25__SCAN_IN), .C2(keyinput_g47), .A(n15115), .ZN(n15118)
         );
  AOI22_X1 U16646 ( .A1(P3_WR_REG_SCAN_IN), .A2(keyinput_g0), .B1(
        P3_REG3_REG_15__SCAN_IN), .B2(keyinput_g63), .ZN(n15116) );
  OAI221_X1 U16647 ( .B1(P3_WR_REG_SCAN_IN), .B2(keyinput_g0), .C1(
        P3_REG3_REG_15__SCAN_IN), .C2(keyinput_g63), .A(n15116), .ZN(n15117)
         );
  NOR4_X1 U16648 ( .A1(n15120), .A2(n15119), .A3(n15118), .A4(n15117), .ZN(
        n15130) );
  AOI22_X1 U16649 ( .A1(P3_REG3_REG_18__SCAN_IN), .A2(keyinput_g60), .B1(
        P3_STATE_REG_SCAN_IN), .B2(keyinput_g34), .ZN(n15121) );
  OAI221_X1 U16650 ( .B1(P3_REG3_REG_18__SCAN_IN), .B2(keyinput_g60), .C1(
        P3_STATE_REG_SCAN_IN), .C2(keyinput_g34), .A(n15121), .ZN(n15128) );
  AOI22_X1 U16651 ( .A1(SI_12_), .A2(keyinput_g20), .B1(SI_29_), .B2(
        keyinput_g3), .ZN(n15122) );
  OAI221_X1 U16652 ( .B1(SI_12_), .B2(keyinput_g20), .C1(SI_29_), .C2(
        keyinput_g3), .A(n15122), .ZN(n15127) );
  AOI22_X1 U16653 ( .A1(SI_20_), .A2(keyinput_g12), .B1(
        P3_REG3_REG_20__SCAN_IN), .B2(keyinput_g55), .ZN(n15123) );
  OAI221_X1 U16654 ( .B1(SI_20_), .B2(keyinput_g12), .C1(
        P3_REG3_REG_20__SCAN_IN), .C2(keyinput_g55), .A(n15123), .ZN(n15126)
         );
  AOI22_X1 U16655 ( .A1(SI_4_), .A2(keyinput_g28), .B1(SI_8_), .B2(
        keyinput_g24), .ZN(n15124) );
  OAI221_X1 U16656 ( .B1(SI_4_), .B2(keyinput_g28), .C1(SI_8_), .C2(
        keyinput_g24), .A(n15124), .ZN(n15125) );
  NOR4_X1 U16657 ( .A1(n15128), .A2(n15127), .A3(n15126), .A4(n15125), .ZN(
        n15129) );
  NAND4_X1 U16658 ( .A1(n15132), .A2(n15131), .A3(n15130), .A4(n15129), .ZN(
        n15232) );
  OAI22_X1 U16659 ( .A1(SI_31_), .A2(keyinput_f1), .B1(keyinput_f0), .B2(
        P3_WR_REG_SCAN_IN), .ZN(n15133) );
  AOI221_X1 U16660 ( .B1(SI_31_), .B2(keyinput_f1), .C1(P3_WR_REG_SCAN_IN), 
        .C2(keyinput_f0), .A(n15133), .ZN(n15150) );
  OAI22_X1 U16661 ( .A1(SI_21_), .A2(keyinput_f11), .B1(keyinput_f12), .B2(
        SI_20_), .ZN(n15134) );
  AOI221_X1 U16662 ( .B1(SI_21_), .B2(keyinput_f11), .C1(SI_20_), .C2(
        keyinput_f12), .A(n15134), .ZN(n15149) );
  AOI22_X1 U16663 ( .A1(SI_26_), .A2(keyinput_f6), .B1(P3_REG3_REG_18__SCAN_IN), .B2(keyinput_f60), .ZN(n15135) );
  OAI221_X1 U16664 ( .B1(SI_26_), .B2(keyinput_f6), .C1(
        P3_REG3_REG_18__SCAN_IN), .C2(keyinput_f60), .A(n15135), .ZN(n15142)
         );
  AOI22_X1 U16665 ( .A1(SI_7_), .A2(keyinput_f25), .B1(P3_REG3_REG_5__SCAN_IN), 
        .B2(keyinput_f49), .ZN(n15136) );
  OAI221_X1 U16666 ( .B1(SI_7_), .B2(keyinput_f25), .C1(P3_REG3_REG_5__SCAN_IN), .C2(keyinput_f49), .A(n15136), .ZN(n15141) );
  AOI22_X1 U16667 ( .A1(SI_28_), .A2(keyinput_f4), .B1(P3_REG3_REG_4__SCAN_IN), 
        .B2(keyinput_f52), .ZN(n15137) );
  OAI221_X1 U16668 ( .B1(SI_28_), .B2(keyinput_f4), .C1(P3_REG3_REG_4__SCAN_IN), .C2(keyinput_f52), .A(n15137), .ZN(n15140) );
  AOI22_X1 U16669 ( .A1(SI_17_), .A2(keyinput_f15), .B1(
        P3_REG3_REG_20__SCAN_IN), .B2(keyinput_f55), .ZN(n15138) );
  OAI221_X1 U16670 ( .B1(SI_17_), .B2(keyinput_f15), .C1(
        P3_REG3_REG_20__SCAN_IN), .C2(keyinput_f55), .A(n15138), .ZN(n15139)
         );
  NOR4_X1 U16671 ( .A1(n15142), .A2(n15141), .A3(n15140), .A4(n15139), .ZN(
        n15146) );
  OAI22_X1 U16672 ( .A1(n15144), .A2(keyinput_f16), .B1(keyinput_f30), .B2(
        SI_2_), .ZN(n15143) );
  AOI221_X1 U16673 ( .B1(n15144), .B2(keyinput_f16), .C1(SI_2_), .C2(
        keyinput_f30), .A(n15143), .ZN(n15145) );
  OAI211_X1 U16674 ( .C1(P3_REG3_REG_22__SCAN_IN), .C2(keyinput_f57), .A(
        n15146), .B(n15145), .ZN(n15147) );
  AOI21_X1 U16675 ( .B1(P3_REG3_REG_22__SCAN_IN), .B2(keyinput_f57), .A(n15147), .ZN(n15148) );
  NAND3_X1 U16676 ( .A1(n15150), .A2(n15149), .A3(n15148), .ZN(n15224) );
  OAI22_X1 U16677 ( .A1(P3_REG3_REG_12__SCAN_IN), .A2(keyinput_f46), .B1(
        keyinput_f18), .B2(SI_14_), .ZN(n15151) );
  AOI221_X1 U16678 ( .B1(P3_REG3_REG_12__SCAN_IN), .B2(keyinput_f46), .C1(
        SI_14_), .C2(keyinput_f18), .A(n15151), .ZN(n15158) );
  OAI22_X1 U16679 ( .A1(SI_10_), .A2(keyinput_f22), .B1(SI_23_), .B2(
        keyinput_f9), .ZN(n15152) );
  AOI221_X1 U16680 ( .B1(SI_10_), .B2(keyinput_f22), .C1(keyinput_f9), .C2(
        SI_23_), .A(n15152), .ZN(n15157) );
  OAI22_X1 U16681 ( .A1(P3_REG3_REG_3__SCAN_IN), .A2(keyinput_f40), .B1(
        keyinput_f32), .B2(SI_0_), .ZN(n15153) );
  AOI221_X1 U16682 ( .B1(P3_REG3_REG_3__SCAN_IN), .B2(keyinput_f40), .C1(SI_0_), .C2(keyinput_f32), .A(n15153), .ZN(n15156) );
  OAI22_X1 U16683 ( .A1(P3_REG3_REG_27__SCAN_IN), .A2(keyinput_f36), .B1(
        keyinput_f7), .B2(SI_25_), .ZN(n15154) );
  AOI221_X1 U16684 ( .B1(P3_REG3_REG_27__SCAN_IN), .B2(keyinput_f36), .C1(
        SI_25_), .C2(keyinput_f7), .A(n15154), .ZN(n15155) );
  NAND4_X1 U16685 ( .A1(n15158), .A2(n15157), .A3(n15156), .A4(n15155), .ZN(
        n15223) );
  OAI22_X1 U16686 ( .A1(P3_REG3_REG_10__SCAN_IN), .A2(keyinput_f39), .B1(
        P3_REG3_REG_9__SCAN_IN), .B2(keyinput_f53), .ZN(n15159) );
  AOI221_X1 U16687 ( .B1(P3_REG3_REG_10__SCAN_IN), .B2(keyinput_f39), .C1(
        keyinput_f53), .C2(P3_REG3_REG_9__SCAN_IN), .A(n15159), .ZN(n15166) );
  OAI22_X1 U16688 ( .A1(P3_REG3_REG_24__SCAN_IN), .A2(keyinput_f51), .B1(SI_8_), .B2(keyinput_f24), .ZN(n15160) );
  AOI221_X1 U16689 ( .B1(P3_REG3_REG_24__SCAN_IN), .B2(keyinput_f51), .C1(
        keyinput_f24), .C2(SI_8_), .A(n15160), .ZN(n15165) );
  OAI22_X1 U16690 ( .A1(SI_5_), .A2(keyinput_f27), .B1(keyinput_f44), .B2(
        P3_REG3_REG_1__SCAN_IN), .ZN(n15161) );
  AOI221_X1 U16691 ( .B1(SI_5_), .B2(keyinput_f27), .C1(P3_REG3_REG_1__SCAN_IN), .C2(keyinput_f44), .A(n15161), .ZN(n15164) );
  OAI22_X1 U16692 ( .A1(P3_REG3_REG_15__SCAN_IN), .A2(keyinput_f63), .B1(
        P3_REG3_REG_11__SCAN_IN), .B2(keyinput_f58), .ZN(n15162) );
  AOI221_X1 U16693 ( .B1(P3_REG3_REG_15__SCAN_IN), .B2(keyinput_f63), .C1(
        keyinput_f58), .C2(P3_REG3_REG_11__SCAN_IN), .A(n15162), .ZN(n15163)
         );
  NAND4_X1 U16694 ( .A1(n15166), .A2(n15165), .A3(n15164), .A4(n15163), .ZN(
        n15222) );
  AOI22_X1 U16695 ( .A1(n15169), .A2(keyinput_f5), .B1(keyinput_f33), .B2(
        n15168), .ZN(n15167) );
  OAI221_X1 U16696 ( .B1(n15169), .B2(keyinput_f5), .C1(n15168), .C2(
        keyinput_f33), .A(n15167), .ZN(n15180) );
  AOI22_X1 U16697 ( .A1(n9724), .A2(keyinput_f59), .B1(n15171), .B2(
        keyinput_f8), .ZN(n15170) );
  OAI221_X1 U16698 ( .B1(n9724), .B2(keyinput_f59), .C1(n15171), .C2(
        keyinput_f8), .A(n15170), .ZN(n15179) );
  INV_X1 U16699 ( .A(P3_REG3_REG_14__SCAN_IN), .ZN(n15173) );
  AOI22_X1 U16700 ( .A1(n15174), .A2(keyinput_f20), .B1(n15173), .B2(
        keyinput_f37), .ZN(n15172) );
  OAI221_X1 U16701 ( .B1(n15174), .B2(keyinput_f20), .C1(n15173), .C2(
        keyinput_f37), .A(n15172), .ZN(n15178) );
  AOI22_X1 U16702 ( .A1(n6673), .A2(keyinput_f10), .B1(n15176), .B2(
        keyinput_f35), .ZN(n15175) );
  OAI221_X1 U16703 ( .B1(n6673), .B2(keyinput_f10), .C1(n15176), .C2(
        keyinput_f35), .A(n15175), .ZN(n15177) );
  NOR4_X1 U16704 ( .A1(n15180), .A2(n15179), .A3(n15178), .A4(n15177), .ZN(
        n15220) );
  INV_X1 U16705 ( .A(P3_REG3_REG_13__SCAN_IN), .ZN(n15182) );
  AOI22_X1 U16706 ( .A1(n15182), .A2(keyinput_f56), .B1(n12063), .B2(
        keyinput_f50), .ZN(n15181) );
  OAI221_X1 U16707 ( .B1(n15182), .B2(keyinput_f56), .C1(n12063), .C2(
        keyinput_f50), .A(n15181), .ZN(n15190) );
  AOI22_X1 U16708 ( .A1(SI_19_), .A2(keyinput_f13), .B1(
        P3_REG3_REG_23__SCAN_IN), .B2(keyinput_f38), .ZN(n15183) );
  OAI221_X1 U16709 ( .B1(SI_19_), .B2(keyinput_f13), .C1(
        P3_REG3_REG_23__SCAN_IN), .C2(keyinput_f38), .A(n15183), .ZN(n15189)
         );
  AOI22_X1 U16710 ( .A1(SI_30_), .A2(keyinput_f2), .B1(SI_29_), .B2(
        keyinput_f3), .ZN(n15184) );
  OAI221_X1 U16711 ( .B1(SI_30_), .B2(keyinput_f2), .C1(SI_29_), .C2(
        keyinput_f3), .A(n15184), .ZN(n15188) );
  XNOR2_X1 U16712 ( .A(P3_REG3_REG_6__SCAN_IN), .B(keyinput_f61), .ZN(n15186)
         );
  XNOR2_X1 U16713 ( .A(SI_1_), .B(keyinput_f31), .ZN(n15185) );
  NAND2_X1 U16714 ( .A1(n15186), .A2(n15185), .ZN(n15187) );
  NOR4_X1 U16715 ( .A1(n15190), .A2(n15189), .A3(n15188), .A4(n15187), .ZN(
        n15219) );
  AOI22_X1 U16716 ( .A1(n9524), .A2(keyinput_f54), .B1(n15192), .B2(
        keyinput_f45), .ZN(n15191) );
  OAI221_X1 U16717 ( .B1(n9524), .B2(keyinput_f54), .C1(n15192), .C2(
        keyinput_f45), .A(n15191), .ZN(n15201) );
  AOI22_X1 U16718 ( .A1(P3_U3151), .A2(keyinput_f34), .B1(keyinput_f17), .B2(
        n15194), .ZN(n15193) );
  OAI221_X1 U16719 ( .B1(P3_U3151), .B2(keyinput_f34), .C1(n15194), .C2(
        keyinput_f17), .A(n15193), .ZN(n15200) );
  XNOR2_X1 U16720 ( .A(SI_9_), .B(keyinput_f23), .ZN(n15198) );
  XNOR2_X1 U16721 ( .A(P3_REG3_REG_8__SCAN_IN), .B(keyinput_f43), .ZN(n15197)
         );
  XNOR2_X1 U16722 ( .A(P3_REG3_REG_28__SCAN_IN), .B(keyinput_f42), .ZN(n15196)
         );
  XNOR2_X1 U16723 ( .A(SI_3_), .B(keyinput_f29), .ZN(n15195) );
  NAND4_X1 U16724 ( .A1(n15198), .A2(n15197), .A3(n15196), .A4(n15195), .ZN(
        n15199) );
  NOR3_X1 U16725 ( .A1(n15201), .A2(n15200), .A3(n15199), .ZN(n15218) );
  AOI22_X1 U16726 ( .A1(n15204), .A2(keyinput_f41), .B1(keyinput_f19), .B2(
        n15203), .ZN(n15202) );
  OAI221_X1 U16727 ( .B1(n15204), .B2(keyinput_f41), .C1(n15203), .C2(
        keyinput_f19), .A(n15202), .ZN(n15216) );
  INV_X1 U16728 ( .A(P3_REG3_REG_25__SCAN_IN), .ZN(n15207) );
  AOI22_X1 U16729 ( .A1(n15207), .A2(keyinput_f47), .B1(n15206), .B2(
        keyinput_f62), .ZN(n15205) );
  OAI221_X1 U16730 ( .B1(n15207), .B2(keyinput_f47), .C1(n15206), .C2(
        keyinput_f62), .A(n15205), .ZN(n15215) );
  AOI22_X1 U16731 ( .A1(n15210), .A2(keyinput_f48), .B1(keyinput_f21), .B2(
        n15209), .ZN(n15208) );
  OAI221_X1 U16732 ( .B1(n15210), .B2(keyinput_f48), .C1(n15209), .C2(
        keyinput_f21), .A(n15208), .ZN(n15214) );
  XNOR2_X1 U16733 ( .A(SI_4_), .B(keyinput_f28), .ZN(n15212) );
  XNOR2_X1 U16734 ( .A(SI_18_), .B(keyinput_f14), .ZN(n15211) );
  NAND2_X1 U16735 ( .A1(n15212), .A2(n15211), .ZN(n15213) );
  NOR4_X1 U16736 ( .A1(n15216), .A2(n15215), .A3(n15214), .A4(n15213), .ZN(
        n15217) );
  NAND4_X1 U16737 ( .A1(n15220), .A2(n15219), .A3(n15218), .A4(n15217), .ZN(
        n15221) );
  NOR4_X1 U16738 ( .A1(n15224), .A2(n15223), .A3(n15222), .A4(n15221), .ZN(
        n15227) );
  INV_X1 U16739 ( .A(keyinput_g26), .ZN(n15226) );
  OAI211_X1 U16740 ( .C1(n15227), .C2(keyinput_f26), .A(n15226), .B(n15225), 
        .ZN(n15230) );
  INV_X1 U16741 ( .A(keyinput_f26), .ZN(n15228) );
  OAI211_X1 U16742 ( .C1(n15228), .C2(n15227), .A(SI_6_), .B(keyinput_g26), 
        .ZN(n15229) );
  NAND2_X1 U16743 ( .A1(n15230), .A2(n15229), .ZN(n15231) );
  OAI21_X1 U16744 ( .B1(n15233), .B2(n15232), .A(n15231), .ZN(n15241) );
  NAND2_X1 U16745 ( .A1(n15235), .A2(n15234), .ZN(n15236) );
  OAI21_X1 U16746 ( .B1(n12259), .B2(P1_ADDR_REG_18__SCAN_IN), .A(n15236), 
        .ZN(n15239) );
  XNOR2_X1 U16747 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n15237) );
  XNOR2_X1 U16748 ( .A(n15237), .B(P3_ADDR_REG_19__SCAN_IN), .ZN(n15238) );
  XNOR2_X1 U16749 ( .A(n15239), .B(n15238), .ZN(n15240) );
  XNOR2_X1 U16750 ( .A(n15241), .B(n15240), .ZN(n15242) );
  XNOR2_X1 U16751 ( .A(n15243), .B(n15242), .ZN(SUB_1596_U4) );
  XOR2_X1 U16752 ( .A(n15245), .B(n15244), .Z(SUB_1596_U59) );
  XNOR2_X1 U16753 ( .A(n15246), .B(P2_ADDR_REG_5__SCAN_IN), .ZN(SUB_1596_U58)
         );
  AOI21_X1 U16754 ( .B1(n15248), .B2(n15247), .A(n15253), .ZN(SUB_1596_U53) );
  XNOR2_X1 U16755 ( .A(n15250), .B(n15249), .ZN(SUB_1596_U56) );
  XOR2_X1 U16756 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(n15251), .Z(SUB_1596_U60) );
  XOR2_X1 U16757 ( .A(n15253), .B(n15252), .Z(SUB_1596_U5) );
  AOI211_X1 U7276 ( .C1(n14037), .C2(n14523), .A(n13832), .B(n13831), .ZN(
        n14041) );
  CLKBUF_X2 U7218 ( .A(n9336), .Z(n11750) );
  CLKBUF_X1 U7244 ( .A(n9097), .Z(n11862) );
  INV_X1 U7257 ( .A(n9021), .ZN(n12732) );
  NAND2_X1 U7271 ( .A1(n7435), .A2(n10700), .ZN(n10704) );
  XNOR2_X1 U7277 ( .A(n7934), .B(P3_IR_REG_21__SCAN_IN), .ZN(n10112) );
  CLKBUF_X1 U7297 ( .A(n9593), .Z(n6483) );
  CLKBUF_X2 U7502 ( .A(n11447), .Z(n6487) );
  CLKBUF_X2 U7524 ( .A(n6476), .Z(n6468) );
endmodule

