

module b17_C_AntiSAT_k_128_9 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, U355, U356, U357, U358, U359, U360, U361, 
        U362, U363, U364, U366, U367, U368, U369, U370, U371, U372, U373, U374, 
        U375, U347, U348, U349, U350, U351, U352, U353, U354, U365, U376, U247, 
        U246, U245, U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, 
        U234, U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223, 
        U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254, U255, 
        U256, U257, U258, U259, U260, U261, U262, U263, U264, U265, U266, U267, 
        U268, U269, U270, U271, U272, U273, U274, U275, U276, U277, U278, U279, 
        U280, U281, U282, U212, U215, U213, U214, P3_U3274, P3_U3275, P3_U3276, 
        P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058, P3_U3057, P3_U3056, 
        P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051, P3_U3050, P3_U3049, 
        P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044, P3_U3043, P3_U3042, 
        P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037, P3_U3036, P3_U3035, 
        P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030, P3_U3029, P3_U3280, 
        P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025, P3_U3024, P3_U3023, 
        P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018, P3_U3017, P3_U3016, 
        P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011, P3_U3010, P3_U3009, 
        P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004, P3_U3003, P3_U3002, 
        P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998, P3_U2997, P3_U2996, 
        P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991, P3_U2990, P3_U2989, 
        P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984, P3_U2983, P3_U2982, 
        P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977, P3_U2976, P3_U2975, 
        P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970, P3_U2969, P3_U2968, 
        P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963, P3_U2962, P3_U2961, 
        P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956, P3_U2955, P3_U2954, 
        P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949, P3_U2948, P3_U2947, 
        P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942, P3_U2941, P3_U2940, 
        P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935, P3_U2934, P3_U2933, 
        P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928, P3_U2927, P3_U2926, 
        P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921, P3_U2920, P3_U2919, 
        P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914, P3_U2913, P3_U2912, 
        P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907, P3_U2906, P3_U2905, 
        P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900, P3_U2899, P3_U2898, 
        P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893, P3_U2892, P3_U2891, 
        P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886, P3_U2885, P3_U2884, 
        P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879, P3_U2878, P3_U2877, 
        P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872, P3_U2871, P3_U2870, 
        P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288, P3_U3289, P3_U3290, 
        P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863, P3_U2862, P3_U2861, 
        P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856, P3_U2855, P3_U2854, 
        P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849, P3_U2848, P3_U2847, 
        P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842, P3_U2841, P3_U2840, 
        P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835, P3_U2834, P3_U2833, 
        P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828, P3_U2827, P3_U2826, 
        P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821, P3_U2820, P3_U2819, 
        P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814, P3_U2813, P3_U2812, 
        P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807, P3_U2806, P3_U2805, 
        P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800, P3_U2799, P3_U2798, 
        P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793, P3_U2792, P3_U2791, 
        P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786, P3_U2785, P3_U2784, 
        P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779, P3_U2778, P3_U2777, 
        P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772, P3_U2771, P3_U2770, 
        P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765, P3_U2764, P3_U2763, 
        P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758, P3_U2757, P3_U2756, 
        P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751, P3_U2750, P3_U2749, 
        P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744, P3_U2743, P3_U2742, 
        P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737, P3_U2736, P3_U2735, 
        P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730, P3_U2729, P3_U2728, 
        P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723, P3_U2722, P3_U2721, 
        P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716, P3_U2715, P3_U2714, 
        P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709, P3_U2708, P3_U2707, 
        P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702, P3_U2701, P3_U2700, 
        P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695, P3_U2694, P3_U2693, 
        P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688, P3_U2687, P3_U2686, 
        P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681, P3_U2680, P3_U2679, 
        P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674, P3_U2673, P3_U2672, 
        P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667, P3_U2666, P3_U2665, 
        P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660, P3_U2659, P3_U2658, 
        P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653, P3_U2652, P3_U2651, 
        P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646, P3_U2645, P3_U2644, 
        P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639, P3_U3292, P3_U2638, 
        P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636, P3_U3296, P3_U2635, 
        P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299, P2_U3585, P2_U3586, 
        P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211, P2_U3210, P2_U3209, 
        P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206, P2_U3205, P2_U3204, 
        P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199, P2_U3198, P2_U3197, 
        P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192, P2_U3191, P2_U3190, 
        P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185, P2_U3184, P2_U3183, 
        P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593, P2_U3178, P2_U3177, 
        P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172, P2_U3171, P2_U3170, 
        P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165, P2_U3164, P2_U3163, 
        P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158, P2_U3157, P2_U3156, 
        P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151, P2_U3150, P2_U3149, 
        P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144, P2_U3143, P2_U3142, 
        P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137, P2_U3136, P2_U3135, 
        P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130, P2_U3129, P2_U3128, 
        P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123, P2_U3122, P2_U3121, 
        P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116, P2_U3115, P2_U3114, 
        P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109, P2_U3108, P2_U3107, 
        P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102, P2_U3101, P2_U3100, 
        P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095, P2_U3094, P2_U3093, 
        P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088, P2_U3087, P2_U3086, 
        P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081, P2_U3080, P2_U3079, 
        P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074, P2_U3073, P2_U3072, 
        P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067, P2_U3066, P2_U3065, 
        P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060, P2_U3059, P2_U3058, 
        P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053, P2_U3052, P2_U3051, 
        P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596, P2_U3599, P2_U3600, 
        P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604, P2_U3605, P2_U3046, 
        P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041, P2_U3040, P2_U3039, 
        P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034, P2_U3033, P2_U3032, 
        P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027, P2_U3026, P2_U3025, 
        P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020, P2_U3019, P2_U3018, 
        P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013, P2_U3012, P2_U3011, 
        P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006, P2_U3005, P2_U3004, 
        P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999, P2_U2998, P2_U2997, 
        P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992, P2_U2991, P2_U2990, 
        P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985, P2_U2984, P2_U2983, 
        P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978, P2_U2977, P2_U2976, 
        P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971, P2_U2970, P2_U2969, 
        P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964, P2_U2963, P2_U2962, 
        P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957, P2_U2956, P2_U2955, 
        P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950, P2_U2949, P2_U2948, 
        P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943, P2_U2942, P2_U2941, 
        P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936, P2_U2935, P2_U2934, 
        P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929, P2_U2928, P2_U2927, 
        P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922, P2_U2921, P2_U2920, 
        P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915, P2_U2914, P2_U2913, 
        P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908, P2_U2907, P2_U2906, 
        P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901, P2_U2900, P2_U2899, 
        P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894, P2_U2893, P2_U2892, 
        P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887, P2_U2886, P2_U2885, 
        P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880, P2_U2879, P2_U2878, 
        P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873, P2_U2872, P2_U2871, 
        P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866, P2_U2865, P2_U2864, 
        P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859, P2_U2858, P2_U2857, 
        P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852, P2_U2851, P2_U2850, 
        P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845, P2_U2844, P2_U2843, 
        P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838, P2_U2837, P2_U2836, 
        P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831, P2_U2830, P2_U2829, 
        P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824, P2_U2823, P2_U2822, 
        P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609, P2_U2818, P2_U3610, 
        P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612, P2_U2814, P1_U3458, 
        P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225, P1_U3224, P1_U3223, 
        P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217, P1_U3216, 
        P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3210, P1_U3209, 
        P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204, P1_U3203, P1_U3202, 
        P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197, P1_U3196, P1_U3195, 
        P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192, P1_U3191, P1_U3190, 
        P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185, P1_U3184, P1_U3183, 
        P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178, P1_U3177, P1_U3176, 
        P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171, P1_U3170, P1_U3169, 
        P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164, P1_U3466, P1_U3163, 
        P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158, P1_U3157, P1_U3156, 
        P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151, P1_U3150, P1_U3149, 
        P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144, P1_U3143, P1_U3142, 
        P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137, P1_U3136, P1_U3135, 
        P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130, P1_U3129, P1_U3128, 
        P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123, P1_U3122, P1_U3121, 
        P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116, P1_U3115, P1_U3114, 
        P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109, P1_U3108, P1_U3107, 
        P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102, P1_U3101, P1_U3100, 
        P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095, P1_U3094, P1_U3093, 
        P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088, P1_U3087, P1_U3086, 
        P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081, P1_U3080, P1_U3079, 
        P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074, P1_U3073, P1_U3072, 
        P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067, P1_U3066, P1_U3065, 
        P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060, P1_U3059, P1_U3058, 
        P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053, P1_U3052, P1_U3051, 
        P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046, P1_U3045, P1_U3044, 
        P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039, P1_U3038, P1_U3037, 
        P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468, P1_U3469, P1_U3472, 
        P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476, P1_U3477, P1_U3478, 
        P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027, P1_U3026, P1_U3025, 
        P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020, P1_U3019, P1_U3018, 
        P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013, P1_U3012, P1_U3011, 
        P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006, P1_U3005, P1_U3004, 
        P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999, P1_U2998, P1_U2997, 
        P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992, P1_U2991, P1_U2990, 
        P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985, P1_U2984, P1_U2983, 
        P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978, P1_U2977, P1_U2976, 
        P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971, P1_U2970, P1_U2969, 
        P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964, P1_U2963, P1_U2962, 
        P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957, P1_U2956, P1_U2955, 
        P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950, P1_U2949, P1_U2948, 
        P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943, P1_U2942, P1_U2941, 
        P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936, P1_U2935, P1_U2934, 
        P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929, P1_U2928, P1_U2927, 
        P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922, P1_U2921, P1_U2920, 
        P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915, P1_U2914, P1_U2913, 
        P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908, P1_U2907, P1_U2906, 
        P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901, P1_U2900, P1_U2899, 
        P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894, P1_U2893, P1_U2892, 
        P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887, P1_U2886, P1_U2885, 
        P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880, P1_U2879, P1_U2878, 
        P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873, P1_U2872, P1_U2871, 
        P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866, P1_U2865, P1_U2864, 
        P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859, P1_U2858, P1_U2857, 
        P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852, P1_U2851, P1_U2850, 
        P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845, P1_U2844, P1_U2843, 
        P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838, P1_U2837, P1_U2836, 
        P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831, P1_U2830, P1_U2829, 
        P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824, P1_U2823, P1_U2822, 
        P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817, P1_U2816, P1_U2815, 
        P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810, P1_U2809, P1_U2808, 
        P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806, P1_U3484, P1_U2805, 
        P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802, P1_U3487, P1_U2801
 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9637,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
         n17417, n17418, n17419, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969;

  NAND2_X1 U11071 ( .A1(n10823), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15021) );
  NOR2_X1 U11072 ( .A1(n16030), .A2(n14716), .ZN(n20164) );
  NOR2_X1 U11073 ( .A1(n14981), .A2(n14970), .ZN(n14960) );
  NAND2_X1 U11074 ( .A1(n11980), .A2(n11979), .ZN(n13161) );
  INV_X1 U11075 ( .A(n13423), .ZN(n14155) );
  INV_X1 U11076 ( .A(n19906), .ZN(n19839) );
  XNOR2_X1 U11077 ( .A(n11302), .B(n11300), .ZN(n12872) );
  INV_X1 U11078 ( .A(n18834), .ZN(n18204) );
  AND2_X1 U11079 ( .A1(n10262), .A2(n12860), .ZN(n19351) );
  NAND2_X1 U11080 ( .A1(n11287), .A2(n11286), .ZN(n11302) );
  NAND2_X1 U11081 ( .A1(n10067), .A2(n10266), .ZN(n10524) );
  INV_X1 U11082 ( .A(n13985), .ZN(n18228) );
  OR2_X1 U11083 ( .A1(n11280), .A2(n16315), .ZN(n10256) );
  INV_X1 U11084 ( .A(n11137), .ZN(n10940) );
  NAND3_X1 U11085 ( .A1(n10827), .A2(n10830), .A3(n10249), .ZN(n10254) );
  AND2_X1 U11088 ( .A1(n10305), .A2(n13269), .ZN(n11473) );
  INV_X1 U11090 ( .A(n15595), .ZN(n17157) );
  OR2_X1 U11091 ( .A1(n11668), .A2(n13269), .ZN(n11470) );
  NAND2_X1 U11093 ( .A1(n11658), .A2(n13269), .ZN(n10480) );
  INV_X1 U11094 ( .A(n13266), .ZN(n11464) );
  AND2_X1 U11095 ( .A1(n13300), .A2(n11492), .ZN(n11478) );
  AND2_X1 U11096 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10306), .ZN(
        n10448) );
  AND2_X1 U11097 ( .A1(n11492), .A2(n10311), .ZN(n10351) );
  NAND2_X1 U11098 ( .A1(n10066), .A2(n13269), .ZN(n11469) );
  CLKBUF_X2 U11099 ( .A(n12169), .Z(n9646) );
  CLKBUF_X2 U11100 ( .A(n11760), .Z(n12454) );
  CLKBUF_X2 U11101 ( .A(n11825), .Z(n12251) );
  INV_X1 U11102 ( .A(n11850), .ZN(n13639) );
  NOR2_X1 U11103 ( .A1(n13352), .A2(n13360), .ZN(n13402) );
  NAND2_X1 U11104 ( .A1(n10197), .A2(n10196), .ZN(n10204) );
  CLKBUF_X1 U11105 ( .A(n12169), .Z(n9647) );
  CLKBUF_X1 U11106 ( .A(n12169), .Z(n9648) );
  CLKBUF_X2 U11107 ( .A(n11737), .Z(n9652) );
  AND2_X1 U11108 ( .A1(n11714), .A2(n9768), .ZN(n12103) );
  AND2_X1 U11109 ( .A1(n11708), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9976) );
  AND2_X1 U11110 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13179) );
  AND2_X2 U11111 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13257) );
  INV_X2 U11112 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13280) );
  NOR2_X2 U11113 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10311) );
  AND2_X1 U11114 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13181) );
  BUF_X1 U11115 ( .A(n12419), .Z(n9629) );
  CLKBUF_X2 U11116 ( .A(n11772), .Z(n12504) );
  AND2_X1 U11117 ( .A1(n10297), .A2(n11492), .ZN(n10350) );
  AND2_X1 U11118 ( .A1(n10767), .A2(n10180), .ZN(n11180) );
  AND2_X1 U11119 ( .A1(n9976), .A2(n13201), .ZN(n11825) );
  AND2_X1 U11120 ( .A1(n11802), .A2(n11801), .ZN(n11852) );
  XNOR2_X1 U11121 ( .A(n9979), .B(n11939), .ZN(n11920) );
  AND3_X1 U11122 ( .A1(n13759), .A2(n11848), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n12580) );
  AND2_X1 U11123 ( .A1(n11492), .A2(n10307), .ZN(n10380) );
  INV_X1 U11124 ( .A(n11250), .ZN(n10909) );
  OAI22_X1 U11125 ( .A1(n10244), .A2(n13269), .B1(n13251), .B2(n19856), .ZN(
        n10833) );
  AND2_X1 U11126 ( .A1(n10811), .A2(n9854), .ZN(n9851) );
  AND2_X1 U11127 ( .A1(n9976), .A2(n13179), .ZN(n12169) );
  CLKBUF_X2 U11128 ( .A(n10214), .Z(n10863) );
  OAI22_X1 U11129 ( .A1(n13543), .A2(n13542), .B1(n13539), .B2(n19087), .ZN(
        n13711) );
  NAND2_X1 U11130 ( .A1(n10267), .A2(n9674), .ZN(n10421) );
  AND2_X1 U11131 ( .A1(n10305), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11368) );
  NAND2_X1 U11132 ( .A1(n9898), .A2(n17587), .ZN(n17744) );
  CLKBUF_X2 U11133 ( .A(n14068), .Z(n17174) );
  AND3_X1 U11134 ( .A1(n14524), .A2(n9716), .A3(n9997), .ZN(n14487) );
  INV_X1 U11135 ( .A(n15955), .ZN(n9985) );
  AND2_X1 U11136 ( .A1(n14535), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14544) );
  INV_X2 U11137 ( .A(n15808), .ZN(n15955) );
  NOR2_X2 U11138 ( .A1(n14913), .A2(n14901), .ZN(n14903) );
  AND2_X1 U11139 ( .A1(n14951), .A2(n14942), .ZN(n14933) );
  OR2_X1 U11140 ( .A1(n14923), .A2(n14911), .ZN(n14913) );
  NAND2_X1 U11141 ( .A1(n10930), .A2(n19897), .ZN(n19884) );
  OR2_X1 U11143 ( .A1(n13881), .A2(n18656), .ZN(n9675) );
  NAND2_X1 U11144 ( .A1(n18806), .A2(n18813), .ZN(n16907) );
  AND2_X1 U11145 ( .A1(n13648), .A2(n13647), .ZN(n20026) );
  NAND2_X1 U11146 ( .A1(n12689), .A2(n14577), .ZN(n14571) );
  NAND2_X1 U11147 ( .A1(n15435), .A2(n9739), .ZN(n15404) );
  AND2_X1 U11148 ( .A1(n15333), .A2(n15329), .ZN(n16319) );
  AOI211_X1 U11149 ( .C1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(n17516), .A(
        n17515), .B(n17514), .ZN(n17517) );
  INV_X1 U11150 ( .A(n14027), .ZN(n9633) );
  NAND2_X2 U11151 ( .A1(n13326), .A2(n10735), .ZN(n10207) );
  INV_X2 U11152 ( .A(n10764), .ZN(n13326) );
  NAND2_X2 U11153 ( .A1(n20112), .A2(n12630), .ZN(n20106) );
  NAND2_X2 U11154 ( .A1(n20114), .A2(n20113), .ZN(n20112) );
  CLKBUF_X1 U11155 ( .A(n12419), .Z(n9627) );
  BUF_X4 U11156 ( .A(n12419), .Z(n9628) );
  NAND2_X1 U11157 ( .A1(n11488), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10473) );
  BUF_X1 U11158 ( .A(n13888), .Z(n9630) );
  CLKBUF_X1 U11159 ( .A(n12169), .Z(n9631) );
  NAND2_X2 U11160 ( .A1(n13109), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13110) );
  AND2_X4 U11161 ( .A1(n13257), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9632) );
  INV_X2 U11162 ( .A(n9633), .ZN(n9634) );
  INV_X2 U11163 ( .A(n9633), .ZN(n9635) );
  NOR2_X1 U11164 ( .A1(n13875), .A2(n13880), .ZN(n14027) );
  NOR2_X2 U11165 ( .A1(n17836), .A2(n15629), .ZN(n15632) );
  AOI21_X2 U11166 ( .B1(n15164), .B2(n15163), .A(n15082), .ZN(n15153) );
  NOR2_X4 U11167 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13201) );
  NOR2_X4 U11168 ( .A1(n13902), .A2(n13901), .ZN(n18834) );
  XNOR2_X2 U11169 ( .A(n12629), .B(n20150), .ZN(n20114) );
  NAND2_X2 U11170 ( .A1(n20121), .A2(n12622), .ZN(n12629) );
  NOR2_X2 U11171 ( .A1(n13875), .A2(n18656), .ZN(n14026) );
  NAND2_X1 U11172 ( .A1(n18799), .A2(n18789), .ZN(n13875) );
  AND2_X1 U11173 ( .A1(n11713), .A2(n13181), .ZN(n11760) );
  NAND2_X1 U11174 ( .A1(n9817), .A2(n9823), .ZN(n9822) );
  AND2_X1 U11175 ( .A1(n9848), .A2(n9847), .ZN(n9846) );
  AND2_X1 U11176 ( .A1(n13795), .A2(n9733), .ZN(n13836) );
  OR2_X1 U11177 ( .A1(n13661), .A2(n12152), .ZN(n12153) );
  AND2_X1 U11178 ( .A1(n10812), .A2(n10559), .ZN(n10809) );
  NAND2_X1 U11179 ( .A1(n9676), .A2(n10685), .ZN(n10689) );
  AND2_X1 U11180 ( .A1(n14963), .A2(n14950), .ZN(n14951) );
  NAND2_X1 U11181 ( .A1(n20123), .A2(n20122), .ZN(n20121) );
  INV_X1 U11182 ( .A(n17851), .ZN(n17842) );
  NOR2_X1 U11183 ( .A1(n17744), .A2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17723) );
  NAND2_X1 U11184 ( .A1(n9899), .A2(n18092), .ZN(n15715) );
  OR2_X1 U11185 ( .A1(n12000), .A2(n13239), .ZN(n12039) );
  NAND2_X1 U11186 ( .A1(n12000), .A2(n11971), .ZN(n13235) );
  NAND2_X2 U11187 ( .A1(n10067), .A2(n9674), .ZN(n10422) );
  NAND2_X1 U11188 ( .A1(n9763), .A2(n11945), .ZN(n12926) );
  OAI211_X1 U11189 ( .C1(n13474), .C2(n12597), .A(n11944), .B(n11943), .ZN(
        n11945) );
  INV_X2 U11190 ( .A(n18176), .ZN(n18655) );
  NOR2_X1 U11191 ( .A1(n14001), .A2(n15652), .ZN(n15651) );
  NOR2_X1 U11192 ( .A1(n18834), .A2(n17485), .ZN(n17486) );
  NOR2_X1 U11193 ( .A1(n17424), .A2(n14015), .ZN(n16515) );
  NAND2_X1 U11194 ( .A1(n18228), .A2(n18223), .ZN(n13990) );
  NAND2_X1 U11195 ( .A1(n18223), .A2(n13985), .ZN(n18634) );
  AND2_X1 U11196 ( .A1(n11841), .A2(n11840), .ZN(n14185) );
  NAND2_X1 U11197 ( .A1(n11845), .A2(n11844), .ZN(n13760) );
  INV_X1 U11198 ( .A(n15791), .ZN(n20762) );
  NAND2_X2 U11199 ( .A1(n13639), .A2(n11848), .ZN(n15791) );
  NAND2_X1 U11200 ( .A1(n13638), .A2(n13734), .ZN(n13637) );
  INV_X1 U11201 ( .A(n10180), .ZN(n11189) );
  INV_X4 U11202 ( .A(n10930), .ZN(n11518) );
  BUF_X2 U11203 ( .A(n11850), .Z(n13734) );
  NOR2_X2 U11204 ( .A1(n11850), .A2(n11848), .ZN(n13740) );
  AND4_X1 U11205 ( .A1(n11781), .A2(n11780), .A3(n11779), .A4(n11778), .ZN(
        n11787) );
  CLKBUF_X2 U11206 ( .A(n13903), .Z(n17173) );
  CLKBUF_X2 U11207 ( .A(n11777), .Z(n12513) );
  CLKBUF_X2 U11208 ( .A(n11887), .Z(n12503) );
  CLKBUF_X2 U11209 ( .A(n11754), .Z(n12306) );
  BUF_X1 U11210 ( .A(n14068), .Z(n9645) );
  CLKBUF_X2 U11211 ( .A(n11869), .Z(n12506) );
  BUF_X4 U11212 ( .A(n13932), .Z(n9637) );
  INV_X4 U11213 ( .A(n9675), .ZN(n17181) );
  OR2_X1 U11214 ( .A1(n13881), .A2(n13880), .ZN(n17058) );
  NAND2_X4 U11215 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18656) );
  XNOR2_X1 U11216 ( .A(n9772), .B(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14111) );
  NAND2_X1 U11217 ( .A1(n12695), .A2(n12696), .ZN(n9772) );
  AOI21_X1 U11218 ( .B1(n10046), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n10045), .ZN(n15342) );
  AOI21_X1 U11219 ( .B1(n14232), .B2(n14230), .A(n14231), .ZN(n14493) );
  AND2_X1 U11220 ( .A1(n10049), .A2(n10048), .ZN(n15353) );
  OR2_X1 U11221 ( .A1(n15341), .A2(n15340), .ZN(n10045) );
  OAI21_X1 U11222 ( .B1(n10028), .B2(n10031), .A(n10065), .ZN(n11681) );
  OR2_X1 U11223 ( .A1(n10050), .A2(n15332), .ZN(n10049) );
  NOR2_X1 U11224 ( .A1(n15150), .A2(n15352), .ZN(n15332) );
  NAND2_X1 U11225 ( .A1(n10026), .A2(n10025), .ZN(n10031) );
  NOR2_X1 U11226 ( .A1(n15404), .A2(n15335), .ZN(n15336) );
  NAND2_X1 U11227 ( .A1(n15075), .A2(n9688), .ZN(n9787) );
  AND2_X1 U11228 ( .A1(n9956), .A2(n9953), .ZN(n15075) );
  NAND2_X1 U11229 ( .A1(n9849), .A2(n9846), .ZN(n10818) );
  INV_X1 U11230 ( .A(n14777), .ZN(n16157) );
  INV_X1 U11231 ( .A(n16170), .ZN(n15210) );
  AND2_X1 U11232 ( .A1(n9684), .A2(n14785), .ZN(n16170) );
  OR3_X1 U11233 ( .A1(n16133), .A2(n10693), .A3(n11257), .ZN(n11238) );
  NOR2_X1 U11234 ( .A1(n9852), .A2(n16275), .ZN(n9847) );
  NOR2_X1 U11235 ( .A1(n10699), .A2(n15233), .ZN(n15052) );
  NOR2_X1 U11236 ( .A1(n11170), .A2(n11171), .ZN(n11255) );
  OR2_X1 U11237 ( .A1(n16167), .A2(n10693), .ZN(n15016) );
  AND2_X1 U11238 ( .A1(n11243), .A2(n10687), .ZN(n16177) );
  NOR2_X1 U11239 ( .A1(n10704), .A2(n10703), .ZN(n10707) );
  NAND2_X1 U11240 ( .A1(n9770), .A2(n9989), .ZN(n15973) );
  XNOR2_X1 U11241 ( .A(n10564), .B(n13717), .ZN(n13710) );
  NAND2_X1 U11242 ( .A1(n9905), .A2(n9902), .ZN(n17539) );
  NOR2_X1 U11243 ( .A1(n9992), .A2(n9740), .ZN(n9991) );
  NAND2_X1 U11244 ( .A1(n10557), .A2(n10556), .ZN(n10812) );
  OR2_X1 U11245 ( .A1(n10800), .A2(n13717), .ZN(n10807) );
  NAND2_X1 U11246 ( .A1(n10689), .A2(n10690), .ZN(n10704) );
  OAI21_X1 U11247 ( .B1(n10800), .B2(n10506), .A(n19067), .ZN(n10564) );
  NOR2_X1 U11248 ( .A1(n9968), .A2(n15067), .ZN(n9967) );
  NOR2_X1 U11249 ( .A1(n10662), .A2(n10661), .ZN(n10663) );
  NOR2_X1 U11250 ( .A1(n9996), .A2(n9995), .ZN(n9994) );
  NOR2_X1 U11251 ( .A1(n9985), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15929) );
  NAND2_X1 U11252 ( .A1(n14933), .A2(n11154), .ZN(n14923) );
  OAI21_X1 U11253 ( .B1(n10043), .B2(n10042), .A(n10794), .ZN(n10784) );
  AOI21_X1 U11254 ( .B1(n15977), .B2(n9990), .A(n9693), .ZN(n9989) );
  OR2_X1 U11255 ( .A1(n15808), .A2(n12674), .ZN(n13725) );
  XNOR2_X1 U11256 ( .A(n9769), .B(n16105), .ZN(n15977) );
  OR2_X1 U11257 ( .A1(n14845), .A2(n14846), .ZN(n14848) );
  AND2_X2 U11258 ( .A1(n12647), .A2(n12670), .ZN(n15808) );
  NAND2_X1 U11259 ( .A1(n12646), .A2(n12645), .ZN(n9769) );
  AND2_X1 U11260 ( .A1(n14960), .A2(n14961), .ZN(n14963) );
  XNOR2_X1 U11261 ( .A(n12647), .B(n12082), .ZN(n12658) );
  AND2_X1 U11262 ( .A1(n10461), .A2(n10460), .ZN(n10464) );
  NAND2_X1 U11263 ( .A1(n10555), .A2(n10554), .ZN(n10802) );
  OR2_X1 U11264 ( .A1(n12079), .A2(n12078), .ZN(n12649) );
  NAND2_X1 U11265 ( .A1(n12079), .A2(n12078), .ZN(n12647) );
  OR3_X1 U11266 ( .A1(n10537), .A2(n10536), .A3(n10535), .ZN(n10555) );
  NOR2_X1 U11267 ( .A1(n13143), .A2(n9880), .ZN(n13518) );
  NAND2_X1 U11268 ( .A1(n11317), .A2(n11316), .ZN(n12953) );
  NOR2_X1 U11269 ( .A1(n12058), .A2(n12057), .ZN(n12079) );
  NAND2_X1 U11270 ( .A1(n9935), .A2(n9934), .ZN(n14981) );
  AND4_X1 U11271 ( .A1(n10336), .A2(n10335), .A3(n10334), .A4(n10333), .ZN(
        n10339) );
  NAND2_X1 U11272 ( .A1(n12002), .A2(n12039), .ZN(n20171) );
  NOR2_X1 U11273 ( .A1(n13063), .A2(n13064), .ZN(n13049) );
  NAND2_X1 U11274 ( .A1(n17349), .A2(n17852), .ZN(n17773) );
  INV_X1 U11275 ( .A(n10439), .ZN(n10332) );
  INV_X1 U11276 ( .A(n17848), .ZN(n17863) );
  NAND2_X2 U11277 ( .A1(n14179), .A2(n13122), .ZN(n14476) );
  CLKBUF_X1 U11278 ( .A(n13210), .Z(n9655) );
  NOR2_X2 U11280 ( .A1(n10282), .A2(n10277), .ZN(n19381) );
  AND2_X1 U11281 ( .A1(n12958), .A2(n9699), .ZN(n13073) );
  AND2_X1 U11282 ( .A1(n9767), .A2(n11999), .ZN(n13239) );
  OR2_X1 U11283 ( .A1(n10285), .A2(n10275), .ZN(n10283) );
  AND2_X1 U11284 ( .A1(n11924), .A2(n11923), .ZN(n12602) );
  AND2_X1 U11285 ( .A1(n9973), .A2(n9720), .ZN(n10626) );
  NAND2_X1 U11286 ( .A1(n9939), .A2(n9690), .ZN(n13047) );
  AND2_X1 U11287 ( .A1(n11298), .A2(n11294), .ZN(n12856) );
  OR2_X1 U11288 ( .A1(n10607), .A2(n10605), .ZN(n9973) );
  INV_X1 U11289 ( .A(n18054), .ZN(n18630) );
  NOR2_X2 U11290 ( .A1(n19227), .A2(n19614), .ZN(n19228) );
  NOR2_X2 U11291 ( .A1(n19223), .A2(n19614), .ZN(n19224) );
  NOR2_X2 U11292 ( .A1(n19170), .A2(n19614), .ZN(n15506) );
  INV_X1 U11293 ( .A(n11297), .ZN(n12860) );
  NAND2_X1 U11294 ( .A1(n10001), .A2(n11895), .ZN(n11931) );
  NAND2_X1 U11295 ( .A1(n9978), .A2(n9980), .ZN(n20340) );
  NAND2_X1 U11296 ( .A1(n10000), .A2(n9999), .ZN(n11966) );
  CLKBUF_X2 U11297 ( .A(n16911), .Z(n9653) );
  INV_X1 U11298 ( .A(n10569), .ZN(n9975) );
  NAND2_X1 U11299 ( .A1(n10234), .A2(n10233), .ZN(n10825) );
  AND2_X1 U11300 ( .A1(n10258), .A2(n10273), .ZN(n16315) );
  INV_X2 U11301 ( .A(n18636), .ZN(n18635) );
  XNOR2_X1 U11302 ( .A(n10832), .B(n10833), .ZN(n10252) );
  OR2_X1 U11303 ( .A1(n10240), .A2(n10239), .ZN(n10273) );
  NOR2_X1 U11304 ( .A1(n18174), .A2(n18175), .ZN(n18168) );
  OAI22_X1 U11305 ( .A1(n17825), .A2(n9912), .B1(n9913), .B2(n15636), .ZN(
        n15639) );
  OR2_X1 U11306 ( .A1(n11939), .A2(n11938), .ZN(n11947) );
  NAND2_X1 U11307 ( .A1(n9757), .A2(n11915), .ZN(n9979) );
  NAND3_X1 U11308 ( .A1(n10243), .A2(n10242), .A3(n10054), .ZN(n10832) );
  NOR2_X1 U11309 ( .A1(n10957), .A2(n10956), .ZN(n10964) );
  OR2_X1 U11310 ( .A1(n10836), .A2(n12918), .ZN(n10054) );
  NAND2_X2 U11311 ( .A1(n17423), .A2(n18676), .ZN(n17488) );
  AND4_X1 U11312 ( .A1(n11864), .A2(n11855), .A3(n9749), .A4(n11863), .ZN(
        n12946) );
  NOR2_X1 U11313 ( .A1(n9964), .A2(n9965), .ZN(n9963) );
  INV_X1 U11314 ( .A(n9783), .ZN(n9782) );
  AND2_X1 U11315 ( .A1(n12988), .A2(n12987), .ZN(n12990) );
  NOR2_X1 U11316 ( .A1(n15626), .A2(n17849), .ZN(n17838) );
  NOR2_X1 U11317 ( .A1(n17364), .A2(n15630), .ZN(n15634) );
  AND3_X1 U11318 ( .A1(n11178), .A2(n10174), .A3(n10173), .ZN(n10925) );
  NAND2_X1 U11319 ( .A1(n14185), .A2(n14192), .ZN(n12751) );
  AND2_X1 U11320 ( .A1(n10492), .A2(n10491), .ZN(n10514) );
  AND2_X1 U11321 ( .A1(n10931), .A2(n10951), .ZN(n10947) );
  NOR2_X1 U11322 ( .A1(n10926), .A2(n19884), .ZN(n10222) );
  CLKBUF_X1 U11323 ( .A(n11178), .Z(n19899) );
  AND4_X1 U11324 ( .A1(n15580), .A2(n15579), .A3(n15578), .A4(n15577), .ZN(
        n15581) );
  OR2_X1 U11325 ( .A1(n11846), .A2(n9643), .ZN(n13748) );
  INV_X1 U11326 ( .A(n12937), .ZN(n12648) );
  INV_X1 U11327 ( .A(n11180), .ZN(n10926) );
  NAND3_X1 U11328 ( .A1(n13958), .A2(n13957), .A3(n13956), .ZN(n18223) );
  AND2_X1 U11329 ( .A1(n11180), .A2(n10178), .ZN(n11683) );
  INV_X1 U11330 ( .A(n10178), .ZN(n12802) );
  AOI211_X1 U11331 ( .C1(n17174), .C2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A(
        n13955), .B(n13954), .ZN(n13956) );
  NAND2_X1 U11332 ( .A1(n13340), .A2(n11842), .ZN(n11843) );
  INV_X1 U11333 ( .A(n13402), .ZN(n13191) );
  CLKBUF_X1 U11334 ( .A(n11836), .Z(n11932) );
  INV_X1 U11335 ( .A(n13352), .ZN(n13747) );
  AND2_X2 U11336 ( .A1(n11848), .A2(n11850), .ZN(n14162) );
  CLKBUF_X1 U11337 ( .A(n11842), .Z(n14192) );
  NAND2_X2 U11338 ( .A1(n13360), .A2(n11850), .ZN(n13423) );
  CLKBUF_X1 U11339 ( .A(n11881), .Z(n13759) );
  NAND4_X2 U11340 ( .A1(n11789), .A2(n11788), .A3(n11787), .A4(n11786), .ZN(
        n11881) );
  AND4_X1 U11341 ( .A1(n15574), .A2(n15573), .A3(n15572), .A4(n15571), .ZN(
        n15582) );
  NAND2_X1 U11342 ( .A1(n10081), .A2(n10080), .ZN(n10177) );
  NAND2_X2 U11343 ( .A1(n9777), .A2(n9776), .ZN(n10930) );
  OR2_X2 U11344 ( .A1(n11721), .A2(n11720), .ZN(n13344) );
  AND4_X1 U11345 ( .A1(n11814), .A2(n11813), .A3(n11812), .A4(n11811), .ZN(
        n11820) );
  AND4_X1 U11346 ( .A1(n11770), .A2(n11769), .A3(n11768), .A4(n11767), .ZN(
        n11789) );
  AND4_X1 U11347 ( .A1(n11776), .A2(n11775), .A3(n11774), .A4(n11773), .ZN(
        n11788) );
  AND4_X1 U11348 ( .A1(n11806), .A2(n11805), .A3(n11804), .A4(n11803), .ZN(
        n11822) );
  AND4_X1 U11349 ( .A1(n11810), .A2(n11809), .A3(n11808), .A4(n11807), .ZN(
        n11821) );
  AND4_X1 U11350 ( .A1(n11818), .A2(n11817), .A3(n11816), .A4(n11815), .ZN(
        n11819) );
  AND4_X1 U11351 ( .A1(n11741), .A2(n11740), .A3(n11739), .A4(n11738), .ZN(
        n11752) );
  AND4_X1 U11352 ( .A1(n11745), .A2(n11744), .A3(n11743), .A4(n11742), .ZN(
        n11751) );
  AND4_X1 U11353 ( .A1(n11785), .A2(n11784), .A3(n11783), .A4(n11782), .ZN(
        n11786) );
  NAND2_X2 U11354 ( .A1(n19839), .A2(n19776), .ZN(n19835) );
  INV_X4 U11355 ( .A(n16931), .ZN(n17002) );
  AND4_X1 U11356 ( .A1(n11736), .A2(n11735), .A3(n11734), .A4(n11733), .ZN(
        n11753) );
  INV_X1 U11357 ( .A(n17056), .ZN(n17016) );
  BUF_X1 U11358 ( .A(n10407), .Z(n11399) );
  AND4_X1 U11359 ( .A1(n10159), .A2(n10158), .A3(n13269), .A4(n10157), .ZN(
        n10160) );
  INV_X2 U11360 ( .A(n16503), .ZN(U215) );
  NAND2_X2 U11361 ( .A1(n18712), .A2(n20776), .ZN(n18765) );
  BUF_X4 U11362 ( .A(n11882), .Z(n12479) );
  NAND2_X2 U11363 ( .A1(n20776), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18769) );
  NAND2_X1 U11364 ( .A1(n9933), .A2(n9810), .ZN(n16931) );
  CLKBUF_X2 U11365 ( .A(n11755), .Z(n12512) );
  BUF_X2 U11366 ( .A(n13903), .Z(n17144) );
  BUF_X2 U11367 ( .A(n14026), .Z(n17158) );
  NAND2_X1 U11368 ( .A1(n9933), .A2(n9932), .ZN(n17056) );
  OR2_X1 U11369 ( .A1(n18656), .A2(n13877), .ZN(n15595) );
  NOR2_X1 U11370 ( .A1(n13879), .A2(n13880), .ZN(n16929) );
  CLKBUF_X3 U11371 ( .A(n11737), .Z(n9651) );
  BUF_X4 U11372 ( .A(n15559), .Z(n9639) );
  INV_X2 U11373 ( .A(n16506), .ZN(n16508) );
  CLKBUF_X2 U11374 ( .A(n11874), .Z(n12514) );
  BUF_X4 U11375 ( .A(n13970), .Z(n9640) );
  CLKBUF_X1 U11376 ( .A(n10316), .Z(n11645) );
  BUF_X4 U11377 ( .A(n13971), .Z(n9641) );
  INV_X2 U11378 ( .A(n16412), .ZN(n9642) );
  AND2_X2 U11379 ( .A1(n11714), .A2(n11713), .ZN(n11882) );
  AND2_X2 U11380 ( .A1(n10307), .A2(n13280), .ZN(n11488) );
  NOR2_X1 U11381 ( .A1(n19083), .A2(n9839), .ZN(n9838) );
  NOR3_X1 U11382 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18789), .A3(
        n18659), .ZN(n13892) );
  NAND2_X1 U11383 ( .A1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n13395), .ZN(
        n13544) );
  NAND2_X1 U11384 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18799), .ZN(
        n13877) );
  NAND2_X1 U11385 ( .A1(n18806), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13880) );
  AND2_X1 U11386 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n13395) );
  NOR2_X1 U11387 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13634) );
  NOR2_X2 U11388 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13255) );
  INV_X1 U11389 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10147) );
  AND2_X1 U11390 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10307) );
  CLKBUF_X1 U11391 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15761) );
  INV_X2 U11392 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18799) );
  AOI21_X1 U11393 ( .B1(n14495), .B2(n14653), .A(n14497), .ZN(n14514) );
  NOR2_X1 U11394 ( .A1(n11732), .A2(n13352), .ZN(n12604) );
  OR2_X2 U11395 ( .A1(n10286), .A2(n9657), .ZN(n10425) );
  NAND2_X2 U11396 ( .A1(n13627), .A2(n14858), .ZN(n14851) );
  NAND2_X1 U11397 ( .A1(n9756), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11981) );
  AND2_X1 U11398 ( .A1(n11713), .A2(n9976), .ZN(n11887) );
  OR2_X1 U11399 ( .A1(n11981), .A2(n20903), .ZN(n11944) );
  NOR2_X2 U11400 ( .A1(n13569), .A2(n13614), .ZN(n13613) );
  INV_X2 U11401 ( .A(n17859), .ZN(n17817) );
  AND2_X1 U11402 ( .A1(n11714), .A2(n13179), .ZN(n11755) );
  AND4_X2 U11403 ( .A1(n11752), .A2(n11751), .A3(n11753), .A4(n11750), .ZN(
        n11836) );
  XNOR2_X2 U11404 ( .A(n11562), .B(n11563), .ZN(n14798) );
  NOR2_X2 U11405 ( .A1(n17826), .A2(n17827), .ZN(n17825) );
  NAND2_X1 U11406 ( .A1(n13360), .A2(n11850), .ZN(n9643) );
  NAND2_X1 U11407 ( .A1(n13360), .A2(n11850), .ZN(n9644) );
  AND2_X1 U11408 ( .A1(n11715), .A2(n13179), .ZN(n11772) );
  OAI211_X2 U11409 ( .C1(n14819), .C2(n10020), .A(n10019), .B(n10022), .ZN(
        n11562) );
  AOI21_X2 U11410 ( .B1(n15153), .B2(n15151), .A(n15083), .ZN(n15141) );
  NAND2_X2 U11411 ( .A1(n12928), .A2(n11838), .ZN(n13745) );
  NAND2_X2 U11412 ( .A1(n12743), .A2(n13639), .ZN(n12928) );
  XNOR2_X2 U11413 ( .A(n12621), .B(n20152), .ZN(n20123) );
  NOR2_X1 U11414 ( .A1(n16907), .A2(n13877), .ZN(n14068) );
  NAND2_X2 U11415 ( .A1(n13462), .A2(n12615), .ZN(n12621) );
  XNOR2_X2 U11416 ( .A(n11519), .B(n9731), .ZN(n14819) );
  AND2_X2 U11417 ( .A1(n14824), .A2(n11463), .ZN(n11519) );
  OAI21_X2 U11418 ( .B1(n12612), .B2(n12937), .A(n12611), .ZN(n13109) );
  AOI21_X2 U11419 ( .B1(n12689), .B2(n9982), .A(n9696), .ZN(n9981) );
  NOR2_X2 U11420 ( .A1(n14495), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14536) );
  NAND2_X2 U11421 ( .A1(n14561), .A2(n9981), .ZN(n14495) );
  AND2_X4 U11422 ( .A1(n13300), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9649) );
  BUF_X4 U11423 ( .A(n11737), .Z(n9650) );
  AND2_X1 U11424 ( .A1(n13181), .A2(n13179), .ZN(n11869) );
  XOR2_X1 U11425 ( .A(n16345), .B(n16341), .Z(n16911) );
  AND2_X1 U11426 ( .A1(n13201), .A2(n13181), .ZN(n11874) );
  INV_X2 U11428 ( .A(n13666), .ZN(n19080) );
  NOR2_X4 U11429 ( .A1(n15262), .A2(n15249), .ZN(n15065) );
  NAND2_X2 U11430 ( .A1(n15435), .A2(n9734), .ZN(n15262) );
  OR2_X2 U11431 ( .A1(n11835), .A2(n11834), .ZN(n11850) );
  BUF_X2 U11432 ( .A(n11280), .Z(n9656) );
  BUF_X2 U11433 ( .A(n11280), .Z(n9657) );
  OAI21_X1 U11434 ( .B1(n11172), .B2(n15507), .A(n11184), .ZN(n9783) );
  NAND2_X1 U11435 ( .A1(n9787), .A2(n9687), .ZN(n15013) );
  AND3_X1 U11436 ( .A1(n10483), .A2(n10482), .A3(n10481), .ZN(n10484) );
  NOR2_X1 U11437 ( .A1(n18208), .A2(n15653), .ZN(n13998) );
  OAI21_X1 U11438 ( .B1(n13996), .B2(n13995), .A(n14016), .ZN(n15652) );
  NAND2_X1 U11439 ( .A1(n18233), .A2(n16534), .ZN(n14004) );
  NAND2_X1 U11440 ( .A1(n9753), .A2(n9752), .ZN(n12058) );
  NOR2_X1 U11441 ( .A1(n13239), .A2(n10011), .ZN(n9753) );
  INV_X1 U11442 ( .A(n12000), .ZN(n9752) );
  INV_X1 U11443 ( .A(n10057), .ZN(n10011) );
  NAND2_X1 U11444 ( .A1(n11917), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11939) );
  OR2_X1 U11445 ( .A1(n11848), .A2(n9755), .ZN(n11987) );
  OAI21_X1 U11446 ( .B1(n12677), .B2(n9993), .A(n9991), .ZN(n9751) );
  NOR2_X1 U11447 ( .A1(n9994), .A2(n9993), .ZN(n9992) );
  NOR2_X1 U11448 ( .A1(n14400), .A2(n9874), .ZN(n9873) );
  INV_X1 U11449 ( .A(n13810), .ZN(n9874) );
  AND2_X1 U11450 ( .A1(n13191), .A2(n13637), .ZN(n9749) );
  NAND2_X1 U11451 ( .A1(n14162), .A2(n13423), .ZN(n14158) );
  NAND2_X1 U11452 ( .A1(n9747), .A2(n11920), .ZN(n11949) );
  INV_X1 U11453 ( .A(n9980), .ZN(n9747) );
  NOR2_X1 U11454 ( .A1(n10190), .A2(n11518), .ZN(n10191) );
  NAND2_X1 U11455 ( .A1(n10667), .A2(n10685), .ZN(n10665) );
  NAND2_X1 U11456 ( .A1(n10561), .A2(n10560), .ZN(n10572) );
  OR2_X2 U11457 ( .A1(n10217), .A2(n18853), .ZN(n10836) );
  AND2_X1 U11458 ( .A1(n10843), .A2(n12957), .ZN(n9887) );
  INV_X1 U11459 ( .A(n13029), .ZN(n10843) );
  INV_X1 U11460 ( .A(n15050), .ZN(n9786) );
  NAND2_X1 U11461 ( .A1(n10644), .A2(n10059), .ZN(n10645) );
  AND2_X1 U11462 ( .A1(n9715), .A2(n15086), .ZN(n9819) );
  INV_X1 U11463 ( .A(n13706), .ZN(n9844) );
  NOR2_X1 U11464 ( .A1(n19897), .A2(n10930), .ZN(n10178) );
  AND2_X1 U11465 ( .A1(n15641), .A2(n15672), .ZN(n15615) );
  AOI21_X1 U11466 ( .B1(n13926), .B2(n13925), .A(n13924), .ZN(n15659) );
  NOR2_X1 U11467 ( .A1(n13968), .A2(n13967), .ZN(n14002) );
  NAND2_X1 U11468 ( .A1(n14515), .A2(n9748), .ZN(n14479) );
  AND2_X1 U11469 ( .A1(n12694), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9748) );
  NAND2_X1 U11470 ( .A1(n14524), .A2(n9997), .ZN(n14515) );
  NAND2_X1 U11472 ( .A1(n14790), .A2(n9892), .ZN(n11248) );
  NOR2_X1 U11473 ( .A1(n9894), .A2(n9893), .ZN(n9892) );
  INV_X1 U11474 ( .A(n14791), .ZN(n9893) );
  NAND2_X1 U11475 ( .A1(n9896), .A2(n9895), .ZN(n9894) );
  INV_X1 U11476 ( .A(n10677), .ZN(n9791) );
  AOI21_X1 U11477 ( .B1(n9794), .B2(n9796), .A(n15392), .ZN(n9792) );
  INV_X1 U11478 ( .A(n9794), .ZN(n9793) );
  INV_X1 U11479 ( .A(n9797), .ZN(n9796) );
  AND2_X1 U11480 ( .A1(n9819), .A2(n10660), .ZN(n9818) );
  AND2_X1 U11481 ( .A1(n10782), .A2(n12858), .ZN(n11194) );
  NOR2_X1 U11482 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n16397), .ZN(
        n17511) );
  NAND2_X1 U11483 ( .A1(n16400), .A2(n15615), .ZN(n17587) );
  OAI21_X1 U11484 ( .B1(n14004), .B2(n14003), .A(n18624), .ZN(n15655) );
  NOR2_X1 U11485 ( .A1(n18233), .A2(n9802), .ZN(n9801) );
  INV_X1 U11486 ( .A(n9803), .ZN(n9802) );
  OAI22_X1 U11487 ( .A1(n10426), .A2(n10367), .B1(n11352), .B2(n19689), .ZN(
        n10330) );
  NOR2_X1 U11488 ( .A1(n13164), .A2(n11849), .ZN(n11863) );
  NAND2_X1 U11489 ( .A1(n12538), .A2(n13743), .ZN(n12939) );
  NAND2_X1 U11490 ( .A1(n11842), .A2(n11881), .ZN(n11790) );
  NAND2_X1 U11491 ( .A1(n11836), .A2(n13344), .ZN(n11857) );
  NAND2_X1 U11492 ( .A1(n11919), .A2(n11918), .ZN(n9980) );
  NAND2_X1 U11493 ( .A1(n13743), .A2(n13344), .ZN(n11846) );
  INV_X1 U11494 ( .A(n10629), .ZN(n9972) );
  NOR2_X1 U11495 ( .A1(n10061), .A2(n10387), .ZN(n10396) );
  AND2_X1 U11496 ( .A1(n10041), .A2(n10971), .ZN(n9813) );
  NAND2_X1 U11497 ( .A1(n9781), .A2(n10205), .ZN(n9780) );
  NAND2_X1 U11498 ( .A1(n10285), .A2(n10276), .ZN(n10278) );
  INV_X1 U11499 ( .A(n10196), .ZN(n10198) );
  INV_X1 U11500 ( .A(n17800), .ZN(n9924) );
  NOR2_X1 U11501 ( .A1(n17356), .A2(n15637), .ZN(n15641) );
  NOR2_X1 U11502 ( .A1(n17360), .A2(n15690), .ZN(n15675) );
  INV_X1 U11503 ( .A(n11848), .ZN(n13638) );
  INV_X1 U11504 ( .A(n12497), .ZN(n12524) );
  INV_X1 U11505 ( .A(n14280), .ZN(n10012) );
  AND2_X1 U11506 ( .A1(n14299), .A2(n10014), .ZN(n10013) );
  NAND2_X1 U11507 ( .A1(n10010), .A2(n12269), .ZN(n10009) );
  INV_X1 U11508 ( .A(n14374), .ZN(n10010) );
  INV_X1 U11509 ( .A(n13835), .ZN(n10004) );
  INV_X1 U11510 ( .A(n12086), .ZN(n12527) );
  INV_X1 U11511 ( .A(n12533), .ZN(n12086) );
  INV_X1 U11512 ( .A(n13634), .ZN(n12500) );
  INV_X1 U11513 ( .A(n12500), .ZN(n12528) );
  OR2_X1 U11514 ( .A1(n13340), .A2(n20760), .ZN(n12215) );
  NOR2_X1 U11515 ( .A1(n9877), .A2(n14265), .ZN(n9876) );
  INV_X1 U11516 ( .A(n9878), .ZN(n9877) );
  INV_X1 U11517 ( .A(n9987), .ZN(n9986) );
  INV_X1 U11518 ( .A(n14577), .ZN(n9983) );
  AOI21_X1 U11519 ( .B1(n15955), .B2(n12688), .A(n9988), .ZN(n9987) );
  INV_X1 U11520 ( .A(n13817), .ZN(n9872) );
  INV_X1 U11521 ( .A(n13567), .ZN(n9865) );
  NOR2_X1 U11522 ( .A1(n13435), .A2(n13535), .ZN(n9866) );
  INV_X1 U11523 ( .A(n13579), .ZN(n13432) );
  NAND2_X1 U11524 ( .A1(n11848), .A2(n9713), .ZN(n9863) );
  AOI21_X1 U11525 ( .B1(n10002), .B2(n11894), .A(n11899), .ZN(n9999) );
  AND2_X1 U11526 ( .A1(n10003), .A2(n11930), .ZN(n10002) );
  AND3_X1 U11527 ( .A1(n11913), .A2(n11912), .A3(n11911), .ZN(n11964) );
  XNOR2_X1 U11528 ( .A(n11966), .B(n11964), .ZN(n11968) );
  NOR2_X1 U11529 ( .A1(n9710), .A2(n11914), .ZN(n11915) );
  NAND2_X1 U11530 ( .A1(n9756), .A2(n9754), .ZN(n9757) );
  NAND2_X1 U11531 ( .A1(n11988), .A2(n11987), .ZN(n12556) );
  NOR2_X1 U11532 ( .A1(n14197), .A2(n15826), .ZN(n15789) );
  NOR2_X1 U11533 ( .A1(n10728), .A2(n10727), .ZN(n10746) );
  OAI21_X1 U11534 ( .B1(n10171), .B2(n10934), .A(n10170), .ZN(n10172) );
  NAND3_X1 U11535 ( .A1(n10490), .A2(n10489), .A3(n9961), .ZN(n9965) );
  INV_X1 U11536 ( .A(n10514), .ZN(n9961) );
  INV_X1 U11537 ( .A(n13282), .ZN(n12736) );
  NAND2_X1 U11538 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19880), .ZN(
        n10716) );
  NAND2_X1 U11539 ( .A1(n10034), .A2(n14830), .ZN(n10033) );
  NOR2_X1 U11540 ( .A1(n10036), .A2(n10035), .ZN(n10034) );
  INV_X1 U11541 ( .A(n14837), .ZN(n10035) );
  AND2_X1 U11542 ( .A1(n11288), .A2(n10107), .ZN(n12954) );
  INV_X1 U11543 ( .A(n10187), .ZN(n11701) );
  INV_X1 U11544 ( .A(n13142), .ZN(n9885) );
  NAND2_X1 U11545 ( .A1(n10241), .A2(n10828), .ZN(n10248) );
  NAND2_X1 U11546 ( .A1(n10223), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10244) );
  AND2_X1 U11547 ( .A1(n16187), .A2(n10506), .ZN(n10698) );
  AND2_X1 U11548 ( .A1(n10632), .A2(n15140), .ZN(n9960) );
  AND2_X1 U11549 ( .A1(n9890), .A2(n9889), .ZN(n9888) );
  INV_X1 U11550 ( .A(n14861), .ZN(n9889) );
  AND2_X1 U11551 ( .A1(n9706), .A2(n9883), .ZN(n9882) );
  INV_X1 U11552 ( .A(n13225), .ZN(n9883) );
  NAND2_X1 U11553 ( .A1(n10930), .A2(n19697), .ZN(n11035) );
  INV_X1 U11554 ( .A(n10947), .ZN(n10980) );
  AOI21_X1 U11555 ( .B1(n9658), .B2(n12924), .A(n9941), .ZN(n9940) );
  INV_X1 U11556 ( .A(n12920), .ZN(n9941) );
  INV_X1 U11557 ( .A(n13553), .ZN(n9937) );
  NAND2_X1 U11558 ( .A1(n10837), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10243) );
  AND2_X1 U11559 ( .A1(n10176), .A2(n19697), .ZN(n10951) );
  AND2_X1 U11560 ( .A1(n10934), .A2(n19697), .ZN(n10935) );
  NAND2_X1 U11561 ( .A1(n10285), .A2(n11305), .ZN(n11311) );
  NOR2_X1 U11562 ( .A1(n10256), .A2(n10285), .ZN(n10260) );
  AND3_X1 U11563 ( .A1(n9657), .A2(n9695), .A3(n10255), .ZN(n10262) );
  OR2_X2 U11564 ( .A1(n10285), .A2(n10271), .ZN(n10282) );
  NAND2_X1 U11565 ( .A1(n10262), .A2(n11297), .ZN(n10439) );
  INV_X1 U11566 ( .A(n10256), .ZN(n10266) );
  AND2_X1 U11567 ( .A1(n10285), .A2(n11297), .ZN(n10267) );
  NAND2_X1 U11568 ( .A1(n9656), .A2(n9814), .ZN(n19689) );
  INV_X1 U11569 ( .A(n10278), .ZN(n9814) );
  NAND2_X1 U11570 ( .A1(n15645), .A2(n10052), .ZN(n15711) );
  INV_X1 U11571 ( .A(n10051), .ZN(n9900) );
  OR2_X1 U11572 ( .A1(n9677), .A2(n9903), .ZN(n9902) );
  NAND2_X1 U11573 ( .A1(n9904), .A2(n9906), .ZN(n9903) );
  INV_X1 U11574 ( .A(n17586), .ZN(n9904) );
  OR2_X1 U11575 ( .A1(n17604), .A2(n9907), .ZN(n9905) );
  NOR2_X1 U11576 ( .A1(n17993), .A2(n17690), .ZN(n15720) );
  OR2_X1 U11577 ( .A1(n15633), .A2(n15636), .ZN(n9912) );
  AND2_X1 U11578 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n15635), .ZN(
        n15636) );
  NOR2_X1 U11579 ( .A1(n13948), .A2(n13947), .ZN(n13987) );
  NOR2_X1 U11580 ( .A1(n13938), .A2(n13937), .ZN(n13985) );
  AND2_X1 U11581 ( .A1(n15649), .A2(n18631), .ZN(n14020) );
  OAI21_X1 U11582 ( .B1(n15660), .B2(n13927), .A(n15659), .ZN(n16331) );
  NAND2_X1 U11583 ( .A1(n20029), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13656) );
  NOR2_X1 U11584 ( .A1(n14382), .A2(n9867), .ZN(n14319) );
  OR3_X1 U11585 ( .A1(n9869), .A2(n14139), .A3(n14145), .ZN(n9867) );
  OR2_X1 U11586 ( .A1(n13868), .A2(n13869), .ZN(n14382) );
  AND2_X1 U11587 ( .A1(n13777), .A2(n13776), .ZN(n13778) );
  AND2_X1 U11588 ( .A1(n13779), .A2(n13778), .ZN(n13811) );
  NOR2_X1 U11589 ( .A1(n13701), .A2(n13700), .ZN(n13779) );
  NAND2_X1 U11590 ( .A1(n13613), .A2(n13662), .ZN(n13661) );
  NOR2_X1 U11591 ( .A1(n14232), .A2(n10016), .ZN(n10015) );
  INV_X1 U11592 ( .A(n14243), .ZN(n10016) );
  NAND2_X1 U11593 ( .A1(n12434), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12473) );
  NOR2_X1 U11594 ( .A1(n12321), .A2(n15845), .ZN(n12322) );
  NAND2_X1 U11595 ( .A1(n12322), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12368) );
  INV_X1 U11596 ( .A(n14380), .ZN(n12269) );
  INV_X1 U11597 ( .A(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19976) );
  NAND2_X1 U11598 ( .A1(n13427), .A2(n13423), .ZN(n14163) );
  NAND2_X1 U11599 ( .A1(n14256), .A2(n14244), .ZN(n14246) );
  NAND2_X1 U11600 ( .A1(n12692), .A2(n15808), .ZN(n14524) );
  INV_X1 U11601 ( .A(n14583), .ZN(n9765) );
  NAND2_X1 U11602 ( .A1(n14391), .A2(n13845), .ZN(n13868) );
  NAND2_X1 U11603 ( .A1(n13811), .A2(n9873), .ZN(n14398) );
  OR2_X1 U11604 ( .A1(n13621), .A2(n13622), .ZN(n13701) );
  NAND2_X1 U11605 ( .A1(n20106), .A2(n20105), .ZN(n20104) );
  INV_X1 U11606 ( .A(n20154), .ZN(n14685) );
  NOR2_X1 U11607 ( .A1(n13420), .A2(n9861), .ZN(n13577) );
  OR2_X1 U11608 ( .A1(n13529), .A2(n13421), .ZN(n9861) );
  INV_X1 U11609 ( .A(n13165), .ZN(n11845) );
  NAND2_X1 U11610 ( .A1(n13738), .A2(n13737), .ZN(n13739) );
  AND2_X1 U11611 ( .A1(n13736), .A2(n13735), .ZN(n13737) );
  XNOR2_X1 U11612 ( .A(n9746), .B(n11963), .ZN(n11970) );
  NAND2_X1 U11613 ( .A1(n9745), .A2(n9744), .ZN(n9746) );
  NAND2_X1 U11614 ( .A1(n11961), .A2(n11922), .ZN(n9744) );
  OR2_X1 U11615 ( .A1(n13235), .A2(n12001), .ZN(n20311) );
  INV_X1 U11616 ( .A(n13239), .ZN(n12001) );
  AND2_X1 U11617 ( .A1(n20587), .A2(n20178), .ZN(n20433) );
  OR2_X1 U11618 ( .A1(n9655), .A2(n12612), .ZN(n20552) );
  OR2_X1 U11619 ( .A1(n13235), .A2(n13239), .ZN(n20559) );
  INV_X1 U11620 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20501) );
  NAND2_X1 U11621 ( .A1(n10730), .A2(n10729), .ZN(n10751) );
  MUX2_X1 U11622 ( .A(n10960), .B(n10747), .S(n19884), .Z(n10741) );
  NAND2_X1 U11623 ( .A1(n15076), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15068) );
  OR2_X1 U11624 ( .A1(n10665), .A2(n10614), .ZN(n18881) );
  NOR2_X1 U11625 ( .A1(n10633), .A2(n9726), .ZN(n10614) );
  NAND2_X1 U11626 ( .A1(n9975), .A2(n9974), .ZN(n10597) );
  INV_X1 U11627 ( .A(n10572), .ZN(n10566) );
  NAND2_X1 U11628 ( .A1(n11687), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10489) );
  NAND2_X1 U11629 ( .A1(n10741), .A2(n10671), .ZN(n10490) );
  AOI21_X1 U11630 ( .B1(n11614), .B2(n14781), .A(n9735), .ZN(n10025) );
  INV_X1 U11631 ( .A(n14773), .ZN(n10024) );
  NAND2_X1 U11632 ( .A1(n11613), .A2(n11614), .ZN(n10030) );
  OR2_X1 U11633 ( .A1(n14819), .A2(n14820), .ZN(n10023) );
  NAND2_X1 U11634 ( .A1(n14989), .A2(n14988), .ZN(n14990) );
  INV_X1 U11635 ( .A(n13050), .ZN(n10855) );
  NOR2_X1 U11636 ( .A1(n10812), .A2(n10693), .ZN(n10815) );
  NAND2_X1 U11637 ( .A1(n10811), .A2(n9853), .ZN(n9848) );
  NOR2_X1 U11638 ( .A1(n15174), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9853) );
  INV_X1 U11639 ( .A(n15462), .ZN(n9850) );
  INV_X1 U11640 ( .A(n15174), .ZN(n9854) );
  INV_X1 U11641 ( .A(n13021), .ZN(n9886) );
  NAND2_X1 U11642 ( .A1(n12958), .A2(n9887), .ZN(n13032) );
  AND2_X1 U11643 ( .A1(n18853), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n11305) );
  AND2_X1 U11644 ( .A1(n15065), .A2(n9738), .ZN(n15057) );
  NAND2_X1 U11645 ( .A1(n9968), .A2(n15067), .ZN(n9966) );
  OR2_X1 U11646 ( .A1(n9967), .A2(n9790), .ZN(n9789) );
  NAND2_X1 U11647 ( .A1(n15074), .A2(n10677), .ZN(n9790) );
  NOR2_X1 U11648 ( .A1(n10698), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15050) );
  INV_X1 U11649 ( .A(n9954), .ZN(n9953) );
  OAI21_X1 U11650 ( .B1(n10663), .B2(n9955), .A(n9707), .ZN(n9954) );
  NOR2_X2 U11651 ( .A1(n14839), .A2(n14832), .ZN(n14833) );
  NAND2_X1 U11652 ( .A1(n10615), .A2(n15260), .ZN(n15088) );
  OR2_X1 U11653 ( .A1(n18881), .A2(n10693), .ZN(n10615) );
  AOI21_X1 U11654 ( .B1(n9818), .B2(n15128), .A(n9714), .ZN(n9815) );
  AND2_X1 U11655 ( .A1(n10644), .A2(n10059), .ZN(n9820) );
  AND2_X1 U11656 ( .A1(n10596), .A2(n9697), .ZN(n9797) );
  NOR2_X1 U11657 ( .A1(n9727), .A2(n10595), .ZN(n10596) );
  NAND2_X1 U11658 ( .A1(n9800), .A2(n9799), .ZN(n9798) );
  INV_X1 U11659 ( .A(n15420), .ZN(n9800) );
  NAND2_X1 U11660 ( .A1(n9939), .A2(n9940), .ZN(n16290) );
  INV_X1 U11661 ( .A(n10257), .ZN(n10270) );
  NAND2_X1 U11662 ( .A1(n10240), .A2(n10239), .ZN(n10258) );
  NAND2_X1 U11663 ( .A1(n10127), .A2(n13269), .ZN(n10134) );
  AND2_X1 U11664 ( .A1(n19484), .A2(n19210), .ZN(n19347) );
  INV_X1 U11665 ( .A(n10421), .ZN(n19654) );
  INV_X1 U11666 ( .A(n19645), .ZN(n19701) );
  OR2_X1 U11667 ( .A1(n15501), .A2(n15500), .ZN(n19695) );
  NOR2_X1 U11668 ( .A1(n16326), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15501) );
  INV_X1 U11669 ( .A(n19695), .ZN(n19614) );
  INV_X1 U11670 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19697) );
  INV_X1 U11671 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19691) );
  AND2_X1 U11672 ( .A1(n17511), .A2(n9916), .ZN(n16332) );
  NAND2_X1 U11673 ( .A1(n17604), .A2(n17586), .ZN(n17588) );
  NOR2_X1 U11674 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n15717), .ZN(
        n17589) );
  NAND2_X1 U11675 ( .A1(n9928), .A2(n9925), .ZN(n17632) );
  NAND2_X1 U11676 ( .A1(n17587), .A2(n9930), .ZN(n9927) );
  AND2_X1 U11677 ( .A1(n17723), .A2(n15713), .ZN(n17707) );
  NOR2_X1 U11678 ( .A1(n17801), .A2(n17802), .ZN(n15640) );
  NOR2_X1 U11679 ( .A1(n15639), .A2(n15638), .ZN(n17800) );
  AND2_X1 U11680 ( .A1(n15639), .A2(n15638), .ZN(n17801) );
  XNOR2_X1 U11681 ( .A(n15632), .B(n15631), .ZN(n17826) );
  NOR2_X1 U11682 ( .A1(n14018), .A2(n14017), .ZN(n15671) );
  INV_X1 U11683 ( .A(n16331), .ZN(n18631) );
  CLKBUF_X1 U11684 ( .A(n13209), .Z(n20372) );
  NOR2_X1 U11685 ( .A1(n13292), .A2(n18857), .ZN(n19892) );
  NAND2_X1 U11686 ( .A1(n11268), .A2(n11267), .ZN(n18859) );
  AND2_X1 U11687 ( .A1(n19152), .A2(n11688), .ZN(n15000) );
  NAND2_X1 U11688 ( .A1(n11686), .A2(n12858), .ZN(n19162) );
  INV_X1 U11689 ( .A(n16284), .ZN(n16260) );
  AND2_X1 U11690 ( .A1(n16288), .A2(n19864), .ZN(n16281) );
  NAND2_X1 U11691 ( .A1(n9859), .A2(n9858), .ZN(n9857) );
  AND2_X1 U11692 ( .A1(n11248), .A2(n11227), .ZN(n16145) );
  OR2_X1 U11693 ( .A1(n16319), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10047) );
  INV_X1 U11694 ( .A(n16306), .ZN(n15476) );
  NAND2_X1 U11695 ( .A1(n11194), .A2(n10783), .ZN(n16310) );
  INV_X1 U11696 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19856) );
  AND2_X1 U11697 ( .A1(n19425), .A2(n19617), .ZN(n19414) );
  NOR2_X1 U11698 ( .A1(n14024), .A2(n16999), .ZN(n16978) );
  NAND2_X1 U11699 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n17012), .ZN(n16999) );
  NOR2_X1 U11700 ( .A1(n17069), .A2(n17070), .ZN(n17054) );
  NOR2_X1 U11701 ( .A1(n17124), .A2(n16763), .ZN(n17111) );
  AOI211_X1 U11702 ( .C1(n17002), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n13887), .B(n13886), .ZN(n13888) );
  OR2_X1 U11703 ( .A1(n15833), .A2(n9805), .ZN(n17225) );
  NAND2_X1 U11704 ( .A1(n18196), .A2(n18204), .ZN(n9805) );
  INV_X1 U11705 ( .A(n16413), .ZN(n16414) );
  OR2_X1 U11706 ( .A1(n15721), .A2(n9724), .ZN(n15722) );
  INV_X1 U11707 ( .A(n18175), .ZN(n18166) );
  AOI21_X1 U11708 ( .B1(n11839), .B2(n13340), .A(n9773), .ZN(n11858) );
  INV_X1 U11709 ( .A(n19351), .ZN(n10440) );
  NAND2_X1 U11710 ( .A1(n9785), .A2(n9784), .ZN(n10327) );
  NAND2_X1 U11711 ( .A1(n10260), .A2(n9689), .ZN(n9785) );
  NAND2_X1 U11712 ( .A1(n19351), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n9784) );
  AND2_X1 U11713 ( .A1(n10399), .A2(n10322), .ZN(n10041) );
  NOR2_X1 U11714 ( .A1(n10206), .A2(n18853), .ZN(n9812) );
  AND2_X1 U11715 ( .A1(n11518), .A2(n10204), .ZN(n11177) );
  NOR2_X1 U11716 ( .A1(n18813), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n13914) );
  INV_X1 U11717 ( .A(n12678), .ZN(n9993) );
  OR2_X1 U11718 ( .A1(n12022), .A2(n12021), .ZN(n12639) );
  OR2_X1 U11719 ( .A1(n11910), .A2(n11909), .ZN(n12603) );
  NOR2_X1 U11720 ( .A1(n14741), .A2(n9755), .ZN(n9754) );
  AND2_X2 U11721 ( .A1(n11705), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11714) );
  INV_X1 U11722 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11705) );
  AND2_X2 U11723 ( .A1(n11706), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11713) );
  NOR2_X1 U11724 ( .A1(n11837), .A2(n13171), .ZN(n11841) );
  INV_X1 U11725 ( .A(n10301), .ZN(n11668) );
  INV_X1 U11726 ( .A(n11658), .ZN(n11664) );
  INV_X1 U11727 ( .A(n10463), .ZN(n10465) );
  AND2_X1 U11728 ( .A1(n10766), .A2(n10176), .ZN(n10201) );
  AOI22_X1 U11729 ( .A1(n10301), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9632), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10143) );
  NOR2_X1 U11730 ( .A1(n13877), .A2(n13878), .ZN(n15561) );
  NAND2_X1 U11731 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18813), .ZN(
        n13878) );
  OAI21_X1 U11732 ( .B1(n13987), .B2(n15834), .A(n13998), .ZN(n14012) );
  INV_X1 U11733 ( .A(n13344), .ZN(n11839) );
  NOR2_X1 U11734 ( .A1(n14308), .A2(n14325), .ZN(n10014) );
  NAND2_X1 U11735 ( .A1(n10007), .A2(n12304), .ZN(n10006) );
  INV_X1 U11736 ( .A(n10009), .ZN(n10007) );
  AND2_X1 U11737 ( .A1(n10058), .A2(n13794), .ZN(n10005) );
  NOR2_X1 U11738 ( .A1(n12164), .A2(n13783), .ZN(n12168) );
  NOR2_X1 U11739 ( .A1(n14283), .A2(n9879), .ZN(n9878) );
  INV_X1 U11740 ( .A(n14295), .ZN(n9879) );
  NAND2_X1 U11741 ( .A1(n14512), .A2(n15955), .ZN(n14535) );
  NAND2_X1 U11742 ( .A1(n9870), .A2(n14365), .ZN(n9869) );
  INV_X1 U11743 ( .A(n14340), .ZN(n9870) );
  NOR2_X1 U11744 ( .A1(n12683), .A2(n14595), .ZN(n14583) );
  OR2_X1 U11745 ( .A1(n15808), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12678) );
  INV_X1 U11746 ( .A(n12676), .ZN(n9995) );
  NOR2_X1 U11747 ( .A1(n15955), .A2(n16075), .ZN(n9996) );
  OR2_X1 U11748 ( .A1(n11880), .A2(n11879), .ZN(n12672) );
  INV_X1 U11749 ( .A(n12637), .ZN(n9990) );
  NAND2_X1 U11750 ( .A1(n13734), .A2(n13344), .ZN(n12937) );
  OAI211_X1 U11751 ( .C1(n11867), .C2(n11866), .A(n11865), .B(n11864), .ZN(
        n11918) );
  OR2_X1 U11752 ( .A1(n11998), .A2(n11997), .ZN(n12640) );
  INV_X1 U11753 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n20903) );
  NAND2_X1 U11754 ( .A1(n11986), .A2(n11985), .ZN(n13328) );
  OR2_X1 U11755 ( .A1(n11981), .A2(n13198), .ZN(n11986) );
  OAI21_X1 U11756 ( .B1(n15800), .B2(n14733), .A(n20744), .ZN(n13333) );
  NOR2_X1 U11757 ( .A1(n16166), .A2(n9842), .ZN(n9841) );
  INV_X1 U11758 ( .A(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n9842) );
  NAND2_X1 U11759 ( .A1(n10665), .A2(n10664), .ZN(n10673) );
  NOR2_X1 U11760 ( .A1(n10612), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n9969) );
  NAND2_X1 U11761 ( .A1(n10622), .A2(n10621), .ZN(n10620) );
  INV_X1 U11762 ( .A(n9723), .ZN(n9971) );
  NAND2_X1 U11763 ( .A1(n9970), .A2(n10606), .ZN(n10630) );
  NAND2_X1 U11764 ( .A1(n9975), .A2(n9711), .ZN(n10599) );
  NOR2_X1 U11765 ( .A1(n10568), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n9974) );
  NOR2_X1 U11766 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11492) );
  INV_X1 U11767 ( .A(n11470), .ZN(n11129) );
  CLKBUF_X1 U11768 ( .A(n11489), .Z(n11672) );
  CLKBUF_X1 U11769 ( .A(n11488), .Z(n11671) );
  NAND2_X1 U11770 ( .A1(n9731), .A2(n9670), .ZN(n10022) );
  OR2_X1 U11771 ( .A1(n14804), .A2(n14820), .ZN(n10020) );
  NAND2_X1 U11772 ( .A1(n14853), .A2(n11404), .ZN(n10036) );
  INV_X1 U11773 ( .A(n15366), .ZN(n9943) );
  NOR2_X1 U11774 ( .A1(n18904), .A2(n9830), .ZN(n9829) );
  INV_X1 U11775 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n9830) );
  NOR2_X1 U11776 ( .A1(n16251), .A2(n9834), .ZN(n9833) );
  INV_X1 U11777 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n9834) );
  INV_X1 U11778 ( .A(n13143), .ZN(n9884) );
  INV_X1 U11779 ( .A(n13544), .ZN(n9837) );
  INV_X1 U11780 ( .A(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n19102) );
  AND4_X1 U11781 ( .A1(n10398), .A2(n10397), .A3(n10396), .A4(n10395), .ZN(
        n10960) );
  NAND2_X1 U11782 ( .A1(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n9860) );
  NOR2_X1 U11783 ( .A1(n9897), .A2(n14784), .ZN(n9895) );
  INV_X1 U11784 ( .A(n11226), .ZN(n9897) );
  INV_X1 U11785 ( .A(n14776), .ZN(n9896) );
  INV_X1 U11786 ( .A(n15062), .ZN(n9968) );
  INV_X1 U11787 ( .A(n15264), .ZN(n9955) );
  NOR2_X1 U11788 ( .A1(n10645), .A2(n9950), .ZN(n9949) );
  AND2_X1 U11789 ( .A1(n9795), .A2(n9824), .ZN(n9794) );
  NOR2_X1 U11790 ( .A1(n9826), .A2(n9825), .ZN(n9824) );
  NAND2_X1 U11791 ( .A1(n9797), .A2(n15421), .ZN(n9795) );
  INV_X1 U11792 ( .A(n10604), .ZN(n9825) );
  AND2_X1 U11793 ( .A1(n10822), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9855) );
  NOR2_X1 U11794 ( .A1(n13630), .A2(n9891), .ZN(n9890) );
  INV_X1 U11795 ( .A(n13678), .ZN(n9891) );
  NOR2_X1 U11796 ( .A1(n9946), .A2(n13217), .ZN(n9945) );
  INV_X1 U11797 ( .A(n13247), .ZN(n9946) );
  INV_X1 U11798 ( .A(n13216), .ZN(n9944) );
  NOR2_X1 U11799 ( .A1(n15419), .A2(n15442), .ZN(n10044) );
  AND3_X1 U11800 ( .A1(n10859), .A2(n10858), .A3(n10857), .ZN(n13142) );
  INV_X1 U11801 ( .A(n16291), .ZN(n9938) );
  NAND2_X1 U11802 ( .A1(n10564), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15177) );
  OAI22_X1 U11803 ( .A1(n10225), .A2(n10224), .B1(n10223), .B2(n10222), .ZN(
        n10230) );
  NAND2_X1 U11804 ( .A1(n19846), .A2(n19695), .ZN(n15509) );
  AND4_X1 U11805 ( .A1(n10774), .A2(n10773), .A3(n10772), .A4(n11183), .ZN(
        n12796) );
  AND3_X1 U11806 ( .A1(n10176), .A2(n10198), .A3(n10197), .ZN(n10168) );
  NAND2_X1 U11807 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18789), .ZN(
        n13879) );
  NOR2_X1 U11808 ( .A1(n16907), .A2(n13879), .ZN(n13970) );
  INV_X1 U11809 ( .A(n13875), .ZN(n9932) );
  NOR2_X1 U11810 ( .A1(n13879), .A2(n13878), .ZN(n15559) );
  NOR2_X1 U11811 ( .A1(n13875), .A2(n13878), .ZN(n13932) );
  INV_X1 U11812 ( .A(n13881), .ZN(n9810) );
  NAND2_X1 U11813 ( .A1(n15714), .A2(n9931), .ZN(n9930) );
  OAI21_X1 U11814 ( .B1(n15640), .B2(n9923), .A(n9922), .ZN(n15644) );
  NAND2_X1 U11815 ( .A1(n17787), .A2(n9678), .ZN(n9922) );
  NAND2_X1 U11816 ( .A1(n9924), .A2(n9678), .ZN(n9923) );
  OAI21_X1 U11817 ( .B1(n15615), .B2(n16400), .A(n17587), .ZN(n15643) );
  NOR2_X1 U11818 ( .A1(n15692), .A2(n17797), .ZN(n15694) );
  XNOR2_X1 U11819 ( .A(n15680), .B(n17375), .ZN(n15628) );
  NOR2_X1 U11820 ( .A1(n13986), .A2(n18646), .ZN(n13997) );
  AOI21_X1 U11821 ( .B1(n13996), .B2(n14004), .A(n13994), .ZN(n14016) );
  NOR2_X1 U11822 ( .A1(n18647), .A2(n14012), .ZN(n15649) );
  NOR2_X1 U11823 ( .A1(n18807), .A2(n18693), .ZN(n18195) );
  INV_X1 U11824 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n19953) );
  AND2_X1 U11825 ( .A1(n13699), .A2(n13698), .ZN(n13700) );
  AND2_X1 U11826 ( .A1(n14547), .A2(n13634), .ZN(n12391) );
  NAND2_X1 U11827 ( .A1(n12933), .A2(n12932), .ZN(n13118) );
  INV_X1 U11828 ( .A(n13862), .ZN(n13858) );
  AND2_X1 U11829 ( .A1(n12964), .A2(n12963), .ZN(n20043) );
  INV_X1 U11830 ( .A(n14410), .ZN(n13861) );
  NOR2_X1 U11831 ( .A1(n14192), .A2(n20760), .ZN(n12533) );
  AND2_X1 U11832 ( .A1(n20760), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12532) );
  AND2_X1 U11833 ( .A1(n12433), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12434) );
  OAI21_X1 U11834 ( .B1(n12500), .B2(n14520), .A(n12453), .ZN(n14255) );
  NAND2_X1 U11835 ( .A1(n12396), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12432) );
  INV_X1 U11836 ( .A(n12368), .ZN(n12369) );
  NAND2_X1 U11837 ( .A1(n12370), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12395) );
  AND2_X1 U11838 ( .A1(n12324), .A2(n12323), .ZN(n14339) );
  CLKBUF_X1 U11839 ( .A(n14322), .Z(n14323) );
  CLKBUF_X1 U11840 ( .A(n14337), .Z(n14338) );
  NOR2_X1 U11841 ( .A1(n12284), .A2(n14579), .ZN(n12285) );
  NAND2_X1 U11842 ( .A1(n12285), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12321) );
  AND2_X1 U11843 ( .A1(n12237), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12250) );
  CLKBUF_X1 U11844 ( .A(n13836), .Z(n13837) );
  NOR2_X1 U11845 ( .A1(n12185), .A2(n12199), .ZN(n12219) );
  NAND2_X1 U11846 ( .A1(n12201), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12185) );
  INV_X1 U11847 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n12199) );
  NAND2_X1 U11848 ( .A1(n12136), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12164) );
  NOR2_X1 U11849 ( .A1(n12121), .A2(n19940), .ZN(n12136) );
  OR2_X1 U11850 ( .A1(n12114), .A2(n19953), .ZN(n12121) );
  AND2_X1 U11851 ( .A1(n12120), .A2(n12119), .ZN(n13614) );
  NOR2_X1 U11852 ( .A1(n12071), .A2(n19976), .ZN(n12083) );
  NAND2_X1 U11853 ( .A1(n12077), .A2(n12076), .ZN(n13375) );
  NAND2_X1 U11854 ( .A1(n12649), .A2(n12194), .ZN(n12077) );
  CLKBUF_X1 U11855 ( .A(n13373), .Z(n13374) );
  NAND2_X1 U11856 ( .A1(n12053), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n12071) );
  AOI21_X1 U11857 ( .B1(n12631), .B2(n12194), .A(n12037), .ZN(n13232) );
  NAND2_X1 U11858 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12005) );
  INV_X1 U11859 ( .A(n14162), .ZN(n14198) );
  OR2_X1 U11860 ( .A1(n14246), .A2(n14227), .ZN(n14229) );
  NOR2_X1 U11861 ( .A1(n15808), .A2(n14636), .ZN(n12694) );
  AND2_X1 U11862 ( .A1(n14312), .A2(n9725), .ZN(n14256) );
  INV_X1 U11863 ( .A(n14257), .ZN(n9875) );
  NAND2_X1 U11864 ( .A1(n9984), .A2(n9987), .ZN(n14512) );
  NAND2_X1 U11865 ( .A1(n14571), .A2(n15955), .ZN(n9984) );
  NAND2_X1 U11866 ( .A1(n14312), .A2(n9876), .ZN(n14267) );
  AND2_X1 U11867 ( .A1(n13762), .A2(n13752), .ZN(n14716) );
  NAND2_X1 U11868 ( .A1(n14312), .A2(n9878), .ZN(n14281) );
  AND2_X1 U11869 ( .A1(n14319), .A2(n14310), .ZN(n14312) );
  NAND2_X1 U11870 ( .A1(n14312), .A2(n14295), .ZN(n14297) );
  NOR2_X1 U11871 ( .A1(n9986), .A2(n9983), .ZN(n9982) );
  NOR2_X1 U11872 ( .A1(n14382), .A2(n14139), .ZN(n14372) );
  INV_X1 U11873 ( .A(n14365), .ZN(n9868) );
  AND2_X1 U11874 ( .A1(n13811), .A2(n9712), .ZN(n14391) );
  INV_X1 U11875 ( .A(n14392), .ZN(n9871) );
  NAND2_X1 U11876 ( .A1(n13811), .A2(n9702), .ZN(n14393) );
  NOR2_X1 U11877 ( .A1(n15943), .A2(n9758), .ZN(n14597) );
  NAND2_X1 U11878 ( .A1(n9760), .A2(n9759), .ZN(n9758) );
  INV_X1 U11879 ( .A(n15939), .ZN(n9760) );
  NAND2_X1 U11880 ( .A1(n15808), .A2(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n14598) );
  NAND2_X1 U11881 ( .A1(n14598), .A2(n9761), .ZN(n15943) );
  NAND2_X1 U11882 ( .A1(n15955), .A2(n9762), .ZN(n9761) );
  INV_X1 U11883 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n9762) );
  AND2_X1 U11884 ( .A1(n9705), .A2(n13588), .ZN(n9864) );
  NAND2_X1 U11885 ( .A1(n13432), .A2(n9866), .ZN(n13566) );
  NAND2_X1 U11886 ( .A1(n13432), .A2(n13431), .ZN(n13533) );
  NAND2_X1 U11887 ( .A1(n13577), .A2(n13576), .ZN(n13579) );
  NAND2_X1 U11888 ( .A1(n13418), .A2(n13417), .ZN(n13420) );
  OR2_X1 U11889 ( .A1(n13420), .A2(n13421), .ZN(n13530) );
  INV_X2 U11890 ( .A(n11881), .ZN(n13743) );
  NAND2_X1 U11891 ( .A1(n12929), .A2(n14162), .ZN(n11838) );
  AOI21_X1 U11892 ( .B1(n12602), .B2(n11968), .A(n11967), .ZN(n11969) );
  CLKBUF_X1 U11893 ( .A(n12743), .Z(n12744) );
  INV_X1 U11894 ( .A(n19911), .ZN(n14201) );
  CLKBUF_X1 U11895 ( .A(n13179), .Z(n14745) );
  CLKBUF_X1 U11896 ( .A(n13201), .Z(n13202) );
  INV_X1 U11897 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n14741) );
  NAND2_X1 U11898 ( .A1(n11949), .A2(n11947), .ZN(n9763) );
  INV_X1 U11899 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20553) );
  AND3_X1 U11900 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n9755), .A3(n13333), 
        .ZN(n13361) );
  AOI21_X1 U11901 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20553), .A(n13359), 
        .ZN(n20561) );
  AND2_X1 U11902 ( .A1(n12589), .A2(n12588), .ZN(n14197) );
  NAND2_X1 U11903 ( .A1(n9778), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n9777) );
  NAND2_X1 U11904 ( .A1(n9779), .A2(n13269), .ZN(n9776) );
  OR2_X1 U11905 ( .A1(n10751), .A2(n10750), .ZN(n13282) );
  AND2_X1 U11906 ( .A1(n15042), .A2(n9840), .ZN(n15004) );
  AND2_X1 U11907 ( .A1(n9668), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n9840) );
  AND2_X1 U11908 ( .A1(n9669), .A2(n9736), .ZN(n9947) );
  NAND2_X1 U11909 ( .A1(n15042), .A2(n9841), .ZN(n15031) );
  NAND2_X1 U11910 ( .A1(n15042), .A2(n9668), .ZN(n15025) );
  INV_X1 U11911 ( .A(n10605), .ZN(n10685) );
  NOR2_X2 U11912 ( .A1(n9673), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10684) );
  AND2_X1 U11913 ( .A1(n15167), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15155) );
  INV_X1 U11914 ( .A(n10522), .ZN(n9964) );
  INV_X1 U11915 ( .A(n19884), .ZN(n10731) );
  NAND2_X1 U11916 ( .A1(n10038), .A2(n13224), .ZN(n10037) );
  INV_X1 U11917 ( .A(n10040), .ZN(n10038) );
  NAND2_X1 U11918 ( .A1(n13147), .A2(n13153), .ZN(n10040) );
  INV_X1 U11919 ( .A(n10177), .ZN(n10197) );
  NAND2_X1 U11920 ( .A1(n10030), .A2(n10029), .ZN(n10028) );
  AND2_X1 U11921 ( .A1(n14890), .A2(n14883), .ZN(n9948) );
  AND2_X1 U11922 ( .A1(n14934), .A2(n14919), .ZN(n11154) );
  INV_X1 U11923 ( .A(n14933), .ZN(n14943) );
  INV_X1 U11924 ( .A(n14979), .ZN(n9934) );
  INV_X1 U11925 ( .A(n14990), .ZN(n9935) );
  NOR2_X1 U11926 ( .A1(n13216), .A2(n9942), .ZN(n14989) );
  NAND2_X1 U11927 ( .A1(n9703), .A2(n13583), .ZN(n9942) );
  NOR2_X1 U11928 ( .A1(n13047), .A2(n13046), .ZN(n13158) );
  AOI21_X1 U11929 ( .B1(n11312), .B2(n11315), .A(n11314), .ZN(n11316) );
  NAND2_X1 U11930 ( .A1(n10941), .A2(n10940), .ZN(n10942) );
  OAI21_X1 U11931 ( .B1(n11697), .B2(n11696), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n12902) );
  NAND2_X1 U11932 ( .A1(n19897), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12837) );
  AND2_X1 U11933 ( .A1(n13595), .A2(n12753), .ZN(n19204) );
  INV_X1 U11934 ( .A(n12902), .ZN(n15510) );
  XNOR2_X1 U11935 ( .A(n13591), .B(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14171) );
  NAND2_X1 U11936 ( .A1(n15004), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n13591) );
  NAND2_X1 U11937 ( .A1(n15042), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15044) );
  AND2_X1 U11938 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n11273), .ZN(
        n15076) );
  NAND2_X1 U11939 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n15735), .ZN(
        n15734) );
  AND2_X1 U11940 ( .A1(n15131), .A2(n9828), .ZN(n15735) );
  AND2_X1 U11941 ( .A1(n9667), .A2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9828) );
  NAND2_X1 U11942 ( .A1(n15131), .A2(n9667), .ZN(n15100) );
  AND3_X1 U11943 ( .A1(n15155), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n15131) );
  NAND2_X1 U11944 ( .A1(n15131), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15123) );
  AND3_X1 U11945 ( .A1(n10882), .A2(n10881), .A3(n10880), .ZN(n14861) );
  AND2_X1 U11946 ( .A1(n15750), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15167) );
  AND2_X1 U11947 ( .A1(n15744), .A2(n9832), .ZN(n15750) );
  AND2_X1 U11948 ( .A1(n9666), .A2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n9832) );
  NAND2_X1 U11949 ( .A1(n15744), .A2(n9666), .ZN(n15749) );
  AND3_X1 U11950 ( .A1(n10866), .A2(n10865), .A3(n10864), .ZN(n13225) );
  NAND2_X1 U11951 ( .A1(n9884), .A2(n9706), .ZN(n13226) );
  NAND2_X1 U11952 ( .A1(n15744), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15748) );
  NOR2_X1 U11953 ( .A1(n16265), .A2(n15745), .ZN(n15744) );
  AND3_X1 U11954 ( .A1(n10854), .A2(n10853), .A3(n10852), .ZN(n13050) );
  NOR2_X1 U11955 ( .A1(n13544), .A2(n9836), .ZN(n9835) );
  NOR2_X1 U11956 ( .A1(n15739), .A2(n16278), .ZN(n15738) );
  AND2_X1 U11957 ( .A1(n9837), .A2(n9661), .ZN(n15740) );
  NAND2_X1 U11958 ( .A1(n9837), .A2(n9838), .ZN(n15741) );
  NOR2_X1 U11959 ( .A1(n13544), .A2(n19083), .ZN(n15187) );
  AND3_X1 U11960 ( .A1(n10842), .A2(n10841), .A3(n10840), .ZN(n13029) );
  INV_X1 U11961 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n19083) );
  AND2_X1 U11962 ( .A1(n10248), .A2(n10252), .ZN(n10245) );
  NOR2_X1 U11963 ( .A1(n9860), .A2(n11257), .ZN(n9859) );
  INV_X1 U11964 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n9858) );
  OR2_X1 U11965 ( .A1(n15230), .A2(n11213), .ZN(n15195) );
  NOR2_X2 U11966 ( .A1(n16153), .A2(n10693), .ZN(n15018) );
  XNOR2_X1 U11967 ( .A(n15015), .B(n15014), .ZN(n15030) );
  OR2_X1 U11969 ( .A1(n14814), .A2(n14815), .ZN(n14817) );
  NOR2_X2 U11970 ( .A1(n14817), .A2(n14809), .ZN(n14810) );
  AND3_X1 U11971 ( .A1(n10894), .A2(n10893), .A3(n10892), .ZN(n14832) );
  AND3_X1 U11972 ( .A1(n10891), .A2(n10890), .A3(n10889), .ZN(n14838) );
  AND3_X1 U11973 ( .A1(n10888), .A2(n10887), .A3(n10886), .ZN(n14846) );
  AND2_X1 U11974 ( .A1(n13679), .A2(n9888), .ZN(n14859) );
  AND2_X1 U11975 ( .A1(n15333), .A2(n16312), .ZN(n10050) );
  NAND2_X1 U11976 ( .A1(n13679), .A2(n9890), .ZN(n14860) );
  NAND2_X1 U11977 ( .A1(n13679), .A2(n13678), .ZN(n13677) );
  NAND2_X1 U11978 ( .A1(n9882), .A2(n9881), .ZN(n9880) );
  INV_X1 U11979 ( .A(n13466), .ZN(n9881) );
  NAND2_X1 U11980 ( .A1(n9944), .A2(n9945), .ZN(n15365) );
  NOR2_X1 U11981 ( .A1(n18998), .A2(n10602), .ZN(n15406) );
  AND2_X1 U11982 ( .A1(n15435), .A2(n10044), .ZN(n15418) );
  NAND2_X1 U11983 ( .A1(n15435), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n15434) );
  NAND2_X1 U11984 ( .A1(n10806), .A2(n10801), .ZN(n10804) );
  NAND2_X1 U11985 ( .A1(n15462), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15461) );
  AND2_X1 U11986 ( .A1(n9683), .A2(n13714), .ZN(n9936) );
  AND3_X1 U11987 ( .A1(n10974), .A2(n10973), .A3(n10972), .ZN(n13553) );
  AND2_X1 U11988 ( .A1(n13385), .A2(n9683), .ZN(n13715) );
  AND2_X1 U11989 ( .A1(n10835), .A2(n10834), .ZN(n12958) );
  NAND2_X1 U11990 ( .A1(n12958), .A2(n12957), .ZN(n13030) );
  AND2_X1 U11991 ( .A1(n11200), .A2(n11207), .ZN(n15465) );
  AOI21_X1 U11992 ( .B1(n11297), .B2(n11305), .A(n11296), .ZN(n12855) );
  AND2_X1 U11993 ( .A1(n11291), .A2(n11290), .ZN(n12878) );
  CLKBUF_X1 U11994 ( .A(n10296), .Z(n10297) );
  INV_X1 U11995 ( .A(n18857), .ZN(n12858) );
  AND2_X1 U11996 ( .A1(n19859), .A2(n19209), .ZN(n19263) );
  AND2_X1 U11997 ( .A1(n19484), .A2(n19877), .ZN(n19425) );
  INV_X1 U11998 ( .A(n19263), .ZN(n19485) );
  OR2_X1 U11999 ( .A1(n19859), .A2(n19870), .ZN(n19608) );
  OR2_X1 U12000 ( .A1(n19484), .A2(n19210), .ZN(n19609) );
  INV_X1 U12001 ( .A(n19249), .ZN(n19242) );
  INV_X1 U12002 ( .A(n19250), .ZN(n19244) );
  OR2_X1 U12003 ( .A1(n19484), .A2(n19877), .ZN(n19646) );
  OR2_X1 U12004 ( .A1(n19859), .A2(n19209), .ZN(n19645) );
  NOR2_X2 U12005 ( .A1(n15508), .A2(n15509), .ZN(n19250) );
  OR2_X1 U12006 ( .A1(n19609), .A2(n19645), .ZN(n19211) );
  INV_X1 U12007 ( .A(n10176), .ZN(n19252) );
  NAND2_X1 U12008 ( .A1(n10737), .A2(n10736), .ZN(n15479) );
  NAND2_X1 U12009 ( .A1(n10735), .A2(n10751), .ZN(n10736) );
  NAND2_X1 U12010 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13881) );
  NOR2_X1 U12011 ( .A1(n17030), .A2(n9804), .ZN(n9803) );
  INV_X1 U12012 ( .A(P3_EBX_REG_18__SCAN_IN), .ZN(n9804) );
  NOR2_X1 U12013 ( .A1(n16734), .A2(n17110), .ZN(n17073) );
  NOR2_X1 U12014 ( .A1(n17126), .A2(n9808), .ZN(n9807) );
  INV_X1 U12015 ( .A(P3_EBX_REG_10__SCAN_IN), .ZN(n9808) );
  BUF_X1 U12016 ( .A(n13892), .Z(n17159) );
  NAND2_X1 U12017 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n15577) );
  NAND2_X1 U12018 ( .A1(n9806), .A2(n18827), .ZN(n15833) );
  OR2_X1 U12019 ( .A1(n14020), .A2(n13981), .ZN(n9806) );
  AND3_X1 U12020 ( .A1(n13987), .A2(n17074), .A3(n13997), .ZN(n13981) );
  INV_X1 U12021 ( .A(n13998), .ZN(n14000) );
  NOR2_X1 U12022 ( .A1(n18675), .A2(n18626), .ZN(n17423) );
  AND2_X1 U12023 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n16370), .ZN(
        n16343) );
  INV_X1 U12024 ( .A(n16368), .ZN(n16354) );
  NOR2_X1 U12025 ( .A1(n17492), .A2(n17491), .ZN(n16370) );
  NOR2_X1 U12026 ( .A1(n17615), .A2(n17616), .ZN(n17599) );
  NAND2_X1 U12027 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n17672), .ZN(
        n17647) );
  INV_X1 U12028 ( .A(n18051), .ZN(n17679) );
  NOR2_X1 U12029 ( .A1(n17716), .A2(n17789), .ZN(n17757) );
  INV_X1 U12030 ( .A(n16387), .ZN(n9919) );
  INV_X1 U12031 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n9918) );
  NAND2_X1 U12032 ( .A1(n17510), .A2(n17769), .ZN(n16401) );
  NAND2_X1 U12033 ( .A1(n9910), .A2(n9909), .ZN(n17520) );
  NAND2_X1 U12034 ( .A1(n9901), .A2(n9730), .ZN(n9909) );
  NOR2_X1 U12035 ( .A1(n15704), .A2(n17765), .ZN(n18053) );
  NAND2_X1 U12036 ( .A1(n17767), .A2(n15715), .ZN(n17690) );
  NOR2_X1 U12037 ( .A1(n17766), .A2(n18092), .ZN(n17765) );
  NAND2_X1 U12038 ( .A1(n17768), .A2(n17769), .ZN(n17767) );
  XNOR2_X1 U12039 ( .A(n15644), .B(n15643), .ZN(n17782) );
  NOR2_X1 U12040 ( .A1(n17793), .A2(n18113), .ZN(n17792) );
  NOR2_X1 U12041 ( .A1(n17799), .A2(n17798), .ZN(n17797) );
  INV_X1 U12042 ( .A(n18661), .ZN(n18153) );
  XNOR2_X1 U12043 ( .A(n15628), .B(n15627), .ZN(n17837) );
  NAND2_X1 U12044 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18659) );
  NAND2_X1 U12045 ( .A1(n18845), .A2(n15649), .ZN(n18661) );
  NOR2_X1 U12046 ( .A1(n14005), .A2(n15655), .ZN(n16533) );
  NOR2_X1 U12047 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18195), .ZN(n18495) );
  INV_X1 U12048 ( .A(n14002), .ZN(n18208) );
  INV_X1 U12049 ( .A(n18495), .ZN(n18399) );
  OAI22_X1 U12050 ( .A1(n18628), .A2(n16398), .B1(n16331), .B2(n18630), .ZN(
        n18632) );
  CLKBUF_X1 U12051 ( .A(n12902), .Z(n15508) );
  NAND2_X1 U12052 ( .A1(n12791), .A2(n12981), .ZN(n20765) );
  INV_X1 U12053 ( .A(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n13783) );
  OR2_X1 U12054 ( .A1(n20017), .A2(n13784), .ZN(n19941) );
  INV_X1 U12055 ( .A(n19942), .ZN(n19978) );
  AND2_X1 U12056 ( .A1(n20029), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20013) );
  AND2_X1 U12057 ( .A1(n13648), .A2(n13643), .ZN(n20034) );
  INV_X1 U12058 ( .A(n20026), .ZN(n19991) );
  NAND2_X1 U12059 ( .A1(n13811), .A2(n13810), .ZN(n14401) );
  INV_X1 U12060 ( .A(n14405), .ZN(n13820) );
  INV_X1 U12061 ( .A(n14384), .ZN(n14402) );
  CLKBUF_X1 U12062 ( .A(n14384), .Z(n14377) );
  NAND2_X1 U12063 ( .A1(n14377), .A2(n9773), .ZN(n14379) );
  INV_X1 U12064 ( .A(n13820), .ZN(n14387) );
  OR2_X1 U12065 ( .A1(n13858), .A2(n13861), .ZN(n14466) );
  INV_X1 U12066 ( .A(n14466), .ZN(n14458) );
  AND2_X1 U12067 ( .A1(n13862), .A2(n13861), .ZN(n14468) );
  AND2_X1 U12068 ( .A1(n13858), .A2(n14461), .ZN(n14475) );
  CLKBUF_X1 U12069 ( .A(n20065), .Z(n20768) );
  OR2_X1 U12070 ( .A1(n12594), .A2(n14483), .ZN(n12596) );
  XNOR2_X1 U12071 ( .A(n10017), .B(n14215), .ZN(n14485) );
  NAND2_X1 U12072 ( .A1(n10008), .A2(n12269), .ZN(n14375) );
  INV_X1 U12073 ( .A(n13865), .ZN(n10008) );
  INV_X1 U12074 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n19940) );
  INV_X1 U12075 ( .A(n20130), .ZN(n15961) );
  OAI21_X1 U12076 ( .B1(n14571), .B2(n12688), .A(n15955), .ZN(n14562) );
  NAND2_X1 U12077 ( .A1(n13762), .A2(n13753), .ZN(n20154) );
  NAND2_X1 U12078 ( .A1(n12677), .A2(n12676), .ZN(n13802) );
  NAND2_X1 U12079 ( .A1(n16051), .A2(n20146), .ZN(n16099) );
  NAND2_X1 U12080 ( .A1(n15978), .A2(n15977), .ZN(n15976) );
  NAND2_X1 U12081 ( .A1(n20104), .A2(n12637), .ZN(n15978) );
  OR2_X1 U12082 ( .A1(n12597), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20135) );
  CLKBUF_X1 U12083 ( .A(n13462), .Z(n14712) );
  AND2_X1 U12084 ( .A1(n13762), .A2(n13761), .ZN(n20157) );
  CLKBUF_X1 U12085 ( .A(n11933), .Z(n11934) );
  CLKBUF_X1 U12086 ( .A(n13163), .Z(n20371) );
  NOR2_X1 U12087 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19909) );
  OR2_X1 U12088 ( .A1(n20275), .A2(n20552), .ZN(n20267) );
  OR2_X1 U12089 ( .A1(n20275), .A2(n20466), .ZN(n20315) );
  INV_X1 U12090 ( .A(n20315), .ZN(n20336) );
  OR2_X1 U12091 ( .A1(n20311), .A2(n20429), .ZN(n13511) );
  OAI211_X1 U12092 ( .C1(n13480), .C2(n20379), .A(n20598), .B(n13478), .ZN(
        n13509) );
  OAI211_X1 U12093 ( .C1(n20394), .C2(n20379), .A(n20378), .B(n20433), .ZN(
        n20397) );
  OR2_X1 U12094 ( .A1(n20467), .A2(n20552), .ZN(n20460) );
  OR2_X1 U12095 ( .A1(n20559), .A2(n20500), .ZN(n20564) );
  INV_X1 U12096 ( .A(n20564), .ZN(n20581) );
  INV_X1 U12097 ( .A(n20516), .ZN(n20605) );
  INV_X1 U12098 ( .A(n20534), .ZN(n20625) );
  INV_X1 U12099 ( .A(n20539), .ZN(n20631) );
  OAI211_X1 U12100 ( .C1(n20637), .C2(n20599), .A(n20598), .B(n20597), .ZN(
        n20641) );
  INV_X1 U12101 ( .A(n20530), .ZN(n20652) );
  INV_X1 U12102 ( .A(n20545), .ZN(n20658) );
  NOR2_X1 U12103 ( .A1(n20379), .A2(n14197), .ZN(n15801) );
  AND2_X1 U12104 ( .A1(n20669), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15798) );
  INV_X2 U12105 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20760) );
  INV_X1 U12106 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20379) );
  NOR2_X1 U12107 ( .A1(n12738), .A2(n12737), .ZN(n13595) );
  AND2_X1 U12108 ( .A1(n10193), .A2(n10187), .ZN(n10188) );
  NAND2_X1 U12109 ( .A1(n19080), .A2(n10064), .ZN(n18890) );
  NAND2_X1 U12110 ( .A1(n18890), .A2(n18886), .ZN(n18885) );
  AND2_X1 U12111 ( .A1(n19892), .A2(n13604), .ZN(n19099) );
  OR2_X1 U12112 ( .A1(n19892), .A2(n13603), .ZN(n19110) );
  NAND2_X1 U12113 ( .A1(n16122), .A2(n13600), .ZN(n19064) );
  INV_X1 U12114 ( .A(n19099), .ZN(n19085) );
  NAND2_X1 U12115 ( .A1(n10490), .A2(n10489), .ZN(n10515) );
  NOR2_X1 U12116 ( .A1(n11248), .A2(n11247), .ZN(n11253) );
  AND2_X1 U12117 ( .A1(n10023), .A2(n10018), .ZN(n14807) );
  INV_X1 U12118 ( .A(n11520), .ZN(n10018) );
  CLKBUF_X1 U12119 ( .A(n13625), .Z(n13626) );
  CLKBUF_X1 U12120 ( .A(n13221), .Z(n13222) );
  CLKBUF_X1 U12121 ( .A(n13054), .Z(n13055) );
  CLKBUF_X1 U12122 ( .A(n13052), .Z(n13053) );
  INV_X1 U12123 ( .A(n16315), .ZN(n14760) );
  OR2_X1 U12124 ( .A1(n14856), .A2(n19252), .ZN(n14865) );
  XNOR2_X1 U12125 ( .A(n14767), .B(n14768), .ZN(n14872) );
  NOR2_X1 U12126 ( .A1(n14782), .A2(n14781), .ZN(n14780) );
  OR2_X1 U12128 ( .A1(n12923), .A2(n15000), .ZN(n19134) );
  INV_X1 U12129 ( .A(n19134), .ZN(n19169) );
  NAND2_X1 U12130 ( .A1(n19201), .A2(n12838), .ZN(n19176) );
  INV_X2 U12131 ( .A(n19176), .ZN(n19199) );
  INV_X1 U12132 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n16265) );
  INV_X1 U12133 ( .A(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n16278) );
  NAND2_X1 U12134 ( .A1(n9849), .A2(n9845), .ZN(n16274) );
  AND2_X1 U12135 ( .A1(n9848), .A2(n15173), .ZN(n9845) );
  XNOR2_X1 U12136 ( .A(n10825), .B(n10828), .ZN(n10238) );
  INV_X1 U12137 ( .A(n16281), .ZN(n15182) );
  INV_X1 U12138 ( .A(n16279), .ZN(n16257) );
  INV_X1 U12139 ( .A(n16259), .ZN(n16282) );
  INV_X1 U12140 ( .A(n16288), .ZN(n16252) );
  XNOR2_X1 U12141 ( .A(n11248), .B(n11247), .ZN(n16142) );
  INV_X1 U12142 ( .A(n15035), .ZN(n10823) );
  NAND2_X1 U12143 ( .A1(n9787), .A2(n9679), .ZN(n15049) );
  OR3_X1 U12144 ( .A1(n15283), .A2(n11205), .A3(n15067), .ZN(n15241) );
  NAND2_X1 U12145 ( .A1(n9788), .A2(n10677), .ZN(n15064) );
  OR2_X1 U12146 ( .A1(n15075), .A2(n15074), .ZN(n9788) );
  NAND2_X1 U12147 ( .A1(n9952), .A2(n10663), .ZN(n15263) );
  OAI21_X1 U12148 ( .B1(n9817), .B2(n9816), .A(n9815), .ZN(n15090) );
  INV_X1 U12149 ( .A(n9818), .ZN(n9816) );
  NAND2_X1 U12150 ( .A1(n9821), .A2(n10059), .ZN(n15096) );
  INV_X1 U12151 ( .A(n16312), .ZN(n16294) );
  AND2_X1 U12152 ( .A1(n9827), .A2(n10604), .ZN(n15394) );
  NAND2_X1 U12153 ( .A1(n9798), .A2(n9797), .ZN(n9827) );
  NOR2_X1 U12154 ( .A1(n15471), .A2(n15452), .ZN(n16299) );
  OAI21_X1 U12155 ( .B1(n12925), .B2(n12924), .A(n9658), .ZN(n12921) );
  NAND2_X1 U12156 ( .A1(n13538), .A2(n10799), .ZN(n13709) );
  INV_X1 U12157 ( .A(n15445), .ZN(n16316) );
  INV_X1 U12158 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19880) );
  INV_X1 U12159 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19873) );
  XNOR2_X1 U12160 ( .A(n12856), .B(n12855), .ZN(n19870) );
  INV_X1 U12161 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n19863) );
  INV_X1 U12162 ( .A(n12878), .ZN(n15483) );
  INV_X1 U12163 ( .A(n19870), .ZN(n19209) );
  XNOR2_X1 U12164 ( .A(n12873), .B(n12872), .ZN(n19859) );
  XNOR2_X1 U12165 ( .A(n12915), .B(n12917), .ZN(n19484) );
  CLKBUF_X1 U12166 ( .A(n12916), .Z(n12917) );
  AND2_X1 U12167 ( .A1(n10196), .A2(n10190), .ZN(n10181) );
  INV_X1 U12168 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n20796) );
  AND2_X1 U12169 ( .A1(n19425), .A2(n19548), .ZN(n19372) );
  OR3_X1 U12170 ( .A1(n15504), .A2(n19614), .A3(n15503), .ZN(n19421) );
  INV_X1 U12171 ( .A(n19483), .ZN(n19455) );
  INV_X1 U12172 ( .A(n19541), .ZN(n19518) );
  NOR2_X2 U12173 ( .A1(n19646), .A2(n19847), .ZN(n19569) );
  OR2_X1 U12174 ( .A1(n19578), .A2(n19577), .ZN(n19604) );
  INV_X1 U12175 ( .A(n19711), .ZN(n19661) );
  INV_X1 U12176 ( .A(n19734), .ZN(n19671) );
  INV_X1 U12177 ( .A(n19686), .ZN(n19675) );
  INV_X1 U12178 ( .A(n19750), .ZN(n19681) );
  OAI21_X1 U12179 ( .B1(n19657), .B2(n19656), .A(n19655), .ZN(n19682) );
  OR2_X1 U12180 ( .A1(n19609), .A2(n19608), .ZN(n19686) );
  OAI22_X1 U12181 ( .A1(n14993), .A2(n19244), .B1(n14995), .B2(n19242), .ZN(
        n19703) );
  OAI22_X1 U12182 ( .A1(n19222), .A2(n19244), .B1(n19221), .B2(n19242), .ZN(
        n19708) );
  INV_X1 U12183 ( .A(n19634), .ZN(n19725) );
  OAI22_X1 U12184 ( .A1(n19245), .A2(n19244), .B1(n19243), .B2(n19242), .ZN(
        n19737) );
  INV_X1 U12185 ( .A(n19211), .ZN(n19746) );
  INV_X1 U12186 ( .A(n19607), .ZN(n19745) );
  INV_X1 U12187 ( .A(n17423), .ZN(n17385) );
  AOI21_X1 U12188 ( .B1(n18624), .B2(n18623), .A(n17385), .ZN(n18831) );
  INV_X1 U12189 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17207) );
  INV_X1 U12190 ( .A(n16915), .ZN(n16899) );
  INV_X1 U12191 ( .A(n16909), .ZN(n16925) );
  INV_X1 U12192 ( .A(n16884), .ZN(n16921) );
  INV_X1 U12193 ( .A(n16888), .ZN(n16922) );
  NAND2_X1 U12194 ( .A1(n16977), .A2(P3_EBX_REG_26__SCAN_IN), .ZN(n16969) );
  AND2_X1 U12195 ( .A1(n16983), .A2(P3_EBX_REG_25__SCAN_IN), .ZN(n16977) );
  AND2_X1 U12196 ( .A1(n16978), .A2(n9809), .ZN(n16983) );
  NOR2_X1 U12197 ( .A1(n16640), .A2(n16628), .ZN(n9809) );
  AND2_X1 U12198 ( .A1(n17054), .A2(n9672), .ZN(n17012) );
  NAND2_X1 U12199 ( .A1(n17054), .A2(P3_EBX_REG_18__SCAN_IN), .ZN(n17053) );
  NAND2_X1 U12200 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17111), .ZN(n17110) );
  NAND2_X1 U12201 ( .A1(n17172), .A2(n9671), .ZN(n17124) );
  NAND2_X1 U12202 ( .A1(n17172), .A2(P3_EBX_REG_10__SCAN_IN), .ZN(n17152) );
  NAND2_X1 U12203 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17190), .ZN(n17154) );
  NOR2_X1 U12204 ( .A1(n17155), .A2(n17154), .ZN(n17172) );
  AND4_X1 U12205 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(P3_EBX_REG_6__SCAN_IN), 
        .A3(P3_EBX_REG_5__SCAN_IN), .A4(n17203), .ZN(n17190) );
  INV_X1 U12206 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17197) );
  NOR2_X1 U12207 ( .A1(n17225), .A2(n17192), .ZN(n17203) );
  INV_X1 U12208 ( .A(n17225), .ZN(n17222) );
  INV_X1 U12209 ( .A(n17242), .ZN(n17237) );
  NOR2_X1 U12210 ( .A1(n17450), .A2(n17251), .ZN(n17246) );
  NAND2_X1 U12211 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17254), .ZN(n17251) );
  INV_X1 U12212 ( .A(n17264), .ZN(n17260) );
  NOR2_X1 U12213 ( .A1(n18233), .A2(n17269), .ZN(n17265) );
  NOR3_X1 U12214 ( .A1(n17306), .A2(n17274), .A3(n17233), .ZN(n17270) );
  NOR2_X1 U12215 ( .A1(n17489), .A2(n17313), .ZN(n17307) );
  INV_X1 U12216 ( .A(n17303), .ZN(n17304) );
  AND2_X1 U12217 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17351), .ZN(n17340) );
  NOR2_X1 U12218 ( .A1(n15548), .A2(n15547), .ZN(n17356) );
  INV_X1 U12219 ( .A(n17374), .ZN(n17377) );
  INV_X1 U12220 ( .A(n17371), .ZN(n17376) );
  CLKBUF_X1 U12221 ( .A(n17412), .Z(n17419) );
  CLKBUF_X1 U12222 ( .A(n17486), .Z(n17482) );
  BUF_X1 U12223 ( .A(n17477), .Z(n17485) );
  OR2_X1 U12224 ( .A1(n17510), .A2(n17587), .ZN(n16399) );
  NOR2_X1 U12225 ( .A1(n17572), .A2(n17573), .ZN(n17559) );
  INV_X1 U12226 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n17789) );
  NOR2_X1 U12227 ( .A1(n17818), .A2(n17820), .ZN(n17806) );
  INV_X2 U12228 ( .A(n18571), .ZN(n18397) );
  NOR2_X1 U12229 ( .A1(n17817), .A2(n17819), .ZN(n17856) );
  INV_X1 U12230 ( .A(n17852), .ZN(n17862) );
  XNOR2_X1 U12231 ( .A(n15818), .B(n15821), .ZN(n16362) );
  NAND2_X1 U12232 ( .A1(n9921), .A2(n9920), .ZN(n15818) );
  NAND2_X1 U12233 ( .A1(n17511), .A2(n9915), .ZN(n9920) );
  NOR2_X1 U12234 ( .A1(n17769), .A2(n9917), .ZN(n9915) );
  NAND2_X1 U12235 ( .A1(n9911), .A2(n17587), .ZN(n17538) );
  NAND2_X1 U12236 ( .A1(n17604), .A2(n15719), .ZN(n17545) );
  INV_X1 U12237 ( .A(n9911), .ZN(n17544) );
  NAND2_X1 U12238 ( .A1(n17588), .A2(n16411), .ZN(n17554) );
  AND3_X1 U12239 ( .A1(n9929), .A2(n9928), .A3(n15716), .ZN(n17633) );
  INV_X1 U12240 ( .A(n9929), .ZN(n17643) );
  NOR2_X1 U12241 ( .A1(n17664), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17680) );
  NOR2_X1 U12242 ( .A1(n15640), .A2(n17800), .ZN(n17788) );
  OR2_X1 U12243 ( .A1(n17825), .A2(n15633), .ZN(n9914) );
  AOI21_X2 U12244 ( .B1(n15671), .B2(n15670), .A(n18675), .ZN(n18175) );
  INV_X1 U12245 ( .A(n18141), .ZN(n18179) );
  INV_X1 U12246 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n18639) );
  INV_X1 U12247 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18193) );
  INV_X1 U12248 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18192) );
  INV_X2 U12249 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18806) );
  INV_X2 U12250 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n18789) );
  NOR2_X1 U12251 ( .A1(n14022), .A2(n14021), .ZN(n18814) );
  AND2_X1 U12252 ( .A1(n12710), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14410)
         );
  AND2_X1 U12254 ( .A1(n11703), .A2(n11702), .ZN(n11704) );
  AOI21_X1 U12255 ( .B1(n16145), .B2(n16281), .A(n11277), .ZN(n11278) );
  NAND2_X1 U12256 ( .A1(n15353), .A2(n10047), .ZN(n10046) );
  INV_X1 U12257 ( .A(n16978), .ZN(n16987) );
  NAND2_X1 U12258 ( .A1(n17054), .A2(n9801), .ZN(n17027) );
  AOI21_X1 U12259 ( .B1(n16416), .B2(n16415), .A(n16414), .ZN(n16419) );
  INV_X1 U12260 ( .A(n17058), .ZN(n17075) );
  INV_X1 U12261 ( .A(n15561), .ZN(n15538) );
  NOR2_X2 U12262 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n10754), .ZN(
        n10408) );
  CLKBUF_X1 U12263 ( .A(n11754), .Z(n12486) );
  INV_X1 U12264 ( .A(n9657), .ZN(n10277) );
  AND2_X2 U12265 ( .A1(n10485), .A2(n10484), .ZN(n10693) );
  OAI21_X1 U12266 ( .B1(n17664), .B2(n9930), .A(n17587), .ZN(n9929) );
  OR2_X1 U12267 ( .A1(n10693), .A2(n11137), .ZN(n9658) );
  AND2_X1 U12268 ( .A1(n9787), .A2(n9680), .ZN(n15039) );
  AND2_X1 U12269 ( .A1(n12344), .A2(n10014), .ZN(n14298) );
  AND2_X1 U12270 ( .A1(n9944), .A2(n9703), .ZN(n9659) );
  AND2_X1 U12271 ( .A1(n9970), .A2(n9704), .ZN(n9660) );
  NAND2_X1 U12272 ( .A1(n15435), .A2(n9855), .ZN(n15091) );
  AND2_X1 U12273 ( .A1(n9838), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9661) );
  INV_X1 U12274 ( .A(n16907), .ZN(n9933) );
  AND2_X1 U12275 ( .A1(n9940), .A2(n9938), .ZN(n9662) );
  NAND2_X1 U12276 ( .A1(n10566), .A2(n10565), .ZN(n10569) );
  AND2_X1 U12277 ( .A1(n9902), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n9663) );
  NAND2_X1 U12278 ( .A1(n10032), .A2(n10034), .ZN(n14829) );
  OR2_X1 U12279 ( .A1(n14851), .A2(n11383), .ZN(n9664) );
  NOR3_X1 U12280 ( .A1(n14382), .A2(n9869), .A3(n14139), .ZN(n9665) );
  AND2_X1 U12281 ( .A1(n9833), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9666) );
  AND2_X1 U12282 ( .A1(n9829), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n9667) );
  INV_X1 U12283 ( .A(n15128), .ZN(n9823) );
  NAND2_X1 U12284 ( .A1(n10039), .A2(n13147), .ZN(n13146) );
  AND2_X1 U12285 ( .A1(n9841), .A2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n9668) );
  AND2_X1 U12286 ( .A1(n9948), .A2(n14874), .ZN(n9669) );
  AND2_X1 U12287 ( .A1(n11540), .A2(n11539), .ZN(n9670) );
  AND2_X1 U12288 ( .A1(n9807), .A2(P3_EBX_REG_12__SCAN_IN), .ZN(n9671) );
  AND2_X1 U12289 ( .A1(n9801), .A2(P3_EBX_REG_20__SCAN_IN), .ZN(n9672) );
  OR2_X1 U12290 ( .A1(n10673), .A2(n10672), .ZN(n9673) );
  AND2_X1 U12291 ( .A1(n9657), .A2(n14760), .ZN(n9674) );
  NAND2_X1 U12292 ( .A1(n13795), .A2(n13794), .ZN(n13793) );
  AND2_X1 U12293 ( .A1(n11489), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10407) );
  OR2_X1 U12294 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n10686), .ZN(n9676) );
  NAND2_X1 U12295 ( .A1(n12344), .A2(n10013), .ZN(n14279) );
  AND2_X1 U12296 ( .A1(n15719), .A2(n9908), .ZN(n9677) );
  NAND2_X1 U12297 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15642), .ZN(
        n9678) );
  AND2_X1 U12298 ( .A1(n9789), .A2(n9966), .ZN(n9679) );
  NAND2_X1 U12299 ( .A1(n9798), .A2(n10596), .ZN(n15405) );
  AND2_X1 U12300 ( .A1(n9679), .A2(n9786), .ZN(n9680) );
  OR2_X1 U12301 ( .A1(n10620), .A2(n10612), .ZN(n9681) );
  XNOR2_X1 U12302 ( .A(n11312), .B(n11313), .ZN(n12915) );
  NAND2_X1 U12303 ( .A1(n10287), .A2(n9656), .ZN(n10426) );
  AND2_X1 U12304 ( .A1(n20105), .A2(n15977), .ZN(n9682) );
  NOR2_X1 U12305 ( .A1(n10282), .A2(n9656), .ZN(n10430) );
  AND2_X1 U12306 ( .A1(n9937), .A2(n13384), .ZN(n9683) );
  OR2_X1 U12307 ( .A1(n14793), .A2(n14784), .ZN(n9684) );
  NAND2_X1 U12308 ( .A1(n11970), .A2(n11969), .ZN(n12000) );
  OR2_X1 U12309 ( .A1(n11269), .A2(n16260), .ZN(n9685) );
  OR2_X1 U12310 ( .A1(n13865), .A2(n10009), .ZN(n9686) );
  INV_X1 U12311 ( .A(n10247), .ZN(n10828) );
  AND2_X1 U12312 ( .A1(n9680), .A2(n15040), .ZN(n9687) );
  NOR2_X1 U12313 ( .A1(n9967), .A2(n9791), .ZN(n9688) );
  NAND2_X1 U12314 ( .A1(n11853), .A2(n13740), .ZN(n11864) );
  INV_X2 U12315 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13269) );
  AND2_X1 U12316 ( .A1(n12860), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n9689) );
  AND2_X1 U12317 ( .A1(n9662), .A2(n13045), .ZN(n9690) );
  NAND2_X1 U12318 ( .A1(n9821), .A2(n9820), .ZN(n9691) );
  OR2_X1 U12319 ( .A1(n10836), .A2(n10235), .ZN(n9692) );
  NAND2_X1 U12320 ( .A1(n13795), .A2(n10005), .ZN(n13834) );
  AND2_X1 U12321 ( .A1(n9769), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n9693) );
  NAND2_X1 U12322 ( .A1(n12344), .A2(n12343), .ZN(n14307) );
  AND2_X1 U12323 ( .A1(n15435), .A2(n10822), .ZN(n9694) );
  BUF_X1 U12324 ( .A(n10196), .Z(n10193) );
  BUF_X1 U12325 ( .A(n10196), .Z(n10934) );
  AND2_X1 U12327 ( .A1(n15065), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15056) );
  AND3_X1 U12328 ( .A1(n10254), .A2(n10253), .A3(n14760), .ZN(n9695) );
  NAND2_X1 U12329 ( .A1(n11311), .A2(n11310), .ZN(n11312) );
  AND2_X1 U12330 ( .A1(n9987), .A2(n9985), .ZN(n9696) );
  INV_X2 U12331 ( .A(n19897), .ZN(n15507) );
  AND2_X2 U12332 ( .A1(n10167), .A2(n10166), .ZN(n19897) );
  NAND2_X1 U12333 ( .A1(n15406), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9697) );
  AND2_X1 U12334 ( .A1(n9677), .A2(n10051), .ZN(n9698) );
  AND2_X1 U12335 ( .A1(n9886), .A2(n9887), .ZN(n9699) );
  NAND2_X1 U12336 ( .A1(n10935), .A2(n11518), .ZN(n11137) );
  NAND2_X1 U12337 ( .A1(n12926), .A2(n11950), .ZN(n13187) );
  BUF_X1 U12338 ( .A(n10837), .Z(n10856) );
  BUF_X1 U12339 ( .A(n10856), .Z(n10916) );
  INV_X1 U12340 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10206) );
  INV_X1 U12341 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10069) );
  AND2_X1 U12342 ( .A1(n13762), .A2(n13746), .ZN(n20160) );
  NOR2_X1 U12343 ( .A1(n14851), .A2(n10036), .ZN(n14836) );
  NOR2_X1 U12344 ( .A1(n13216), .A2(n13217), .ZN(n13215) );
  AND2_X1 U12345 ( .A1(n17054), .A2(n9803), .ZN(n9700) );
  AND2_X1 U12346 ( .A1(n15744), .A2(n9833), .ZN(n9701) );
  AND2_X1 U12347 ( .A1(n9873), .A2(n9872), .ZN(n9702) );
  AND2_X1 U12348 ( .A1(n9945), .A2(n9943), .ZN(n9703) );
  AND2_X1 U12349 ( .A1(n10606), .A2(n9972), .ZN(n9704) );
  INV_X1 U12350 ( .A(n15097), .ZN(n10644) );
  AND2_X1 U12351 ( .A1(n14810), .A2(n14799), .ZN(n14790) );
  INV_X1 U12352 ( .A(n15942), .ZN(n9759) );
  INV_X1 U12353 ( .A(n15391), .ZN(n9826) );
  AND2_X1 U12355 ( .A1(n9866), .A2(n9865), .ZN(n9705) );
  AND2_X1 U12356 ( .A1(n9885), .A2(n13150), .ZN(n9706) );
  NAND2_X1 U12357 ( .A1(n15461), .A2(n10811), .ZN(n15172) );
  NOR2_X1 U12358 ( .A1(n13143), .A2(n13142), .ZN(n13144) );
  NAND2_X1 U12359 ( .A1(n10122), .A2(n19252), .ZN(n11176) );
  OR2_X1 U12360 ( .A1(n10669), .A2(n15270), .ZN(n9707) );
  NAND2_X1 U12361 ( .A1(n10563), .A2(n19053), .ZN(n15178) );
  NAND2_X1 U12362 ( .A1(n9884), .A2(n9882), .ZN(n9708) );
  XNOR2_X1 U12363 ( .A(n13661), .B(n12151), .ZN(n13773) );
  OR3_X1 U12364 ( .A1(n14382), .A2(n14139), .A3(n9868), .ZN(n9709) );
  NOR2_X1 U12365 ( .A1(n12597), .A2(n20435), .ZN(n9710) );
  AND2_X1 U12366 ( .A1(n9974), .A2(n10598), .ZN(n9711) );
  AND2_X1 U12367 ( .A1(n9702), .A2(n9871), .ZN(n9712) );
  INV_X1 U12368 ( .A(n14851), .ZN(n10032) );
  AND2_X1 U12369 ( .A1(n11850), .A2(n13411), .ZN(n9713) );
  NAND2_X1 U12370 ( .A1(n10189), .A2(n10168), .ZN(n10764) );
  INV_X1 U12371 ( .A(n15421), .ZN(n9799) );
  INV_X1 U12372 ( .A(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n19052) );
  BUF_X1 U12373 ( .A(n10177), .Z(n11281) );
  AND2_X1 U12374 ( .A1(n10656), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15099) );
  INV_X2 U12375 ( .A(n18196), .ZN(n16534) );
  NOR2_X1 U12376 ( .A1(n9820), .A2(n15099), .ZN(n9714) );
  INV_X1 U12377 ( .A(n11961), .ZN(n12623) );
  AND2_X1 U12378 ( .A1(n15120), .A2(n15107), .ZN(n9715) );
  NOR2_X1 U12379 ( .A1(n15955), .A2(n14635), .ZN(n9716) );
  AND2_X1 U12380 ( .A1(n10621), .A2(n9969), .ZN(n9717) );
  AND2_X1 U12381 ( .A1(n9888), .A2(n14854), .ZN(n9718) );
  INV_X1 U12382 ( .A(n15173), .ZN(n9852) );
  AND2_X1 U12383 ( .A1(n10013), .A2(n10012), .ZN(n9719) );
  AND2_X1 U12384 ( .A1(n9704), .A2(n9971), .ZN(n9720) );
  INV_X1 U12385 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12808) );
  INV_X1 U12386 ( .A(n11842), .ZN(n9773) );
  NAND2_X1 U12387 ( .A1(n12925), .A2(n9658), .ZN(n9939) );
  NAND2_X1 U12388 ( .A1(n13385), .A2(n13384), .ZN(n13386) );
  NOR2_X1 U12389 ( .A1(n13054), .A2(n10040), .ZN(n13152) );
  AND2_X1 U12390 ( .A1(n9939), .A2(n9662), .ZN(n13044) );
  AND2_X1 U12391 ( .A1(n15131), .A2(n9829), .ZN(n9721) );
  AND2_X1 U12392 ( .A1(n17172), .A2(n9807), .ZN(n9722) );
  INV_X1 U12393 ( .A(n17587), .ZN(n17769) );
  AND2_X1 U12394 ( .A1(n11687), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n9723) );
  INV_X1 U12395 ( .A(n18233), .ZN(n17074) );
  AND2_X1 U12396 ( .A1(n17769), .A2(n17875), .ZN(n9724) );
  AND2_X1 U12397 ( .A1(n9876), .A2(n9875), .ZN(n9725) );
  NAND2_X1 U12398 ( .A1(n11687), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n9726) );
  NOR3_X1 U12399 ( .A1(n19009), .A2(n10693), .A3(n15419), .ZN(n9727) );
  AND2_X1 U12400 ( .A1(n13432), .A2(n9705), .ZN(n9728) );
  NOR2_X1 U12401 ( .A1(n15068), .A2(n15055), .ZN(n15042) );
  NOR2_X1 U12402 ( .A1(n17788), .A2(n17787), .ZN(n9729) );
  INV_X1 U12403 ( .A(n13054), .ZN(n10039) );
  OR2_X1 U12404 ( .A1(n17587), .A2(n9900), .ZN(n9730) );
  AND2_X1 U12405 ( .A1(n11516), .A2(n11515), .ZN(n9731) );
  AND2_X1 U12406 ( .A1(n17769), .A2(n9919), .ZN(n9732) );
  INV_X1 U12407 ( .A(n10436), .ZN(n19213) );
  AND2_X1 U12408 ( .A1(n10005), .A2(n10004), .ZN(n9733) );
  INV_X1 U12409 ( .A(n14804), .ZN(n10021) );
  INV_X1 U12410 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n9755) );
  AND2_X1 U12411 ( .A1(n9855), .A2(n10063), .ZN(n9734) );
  NAND2_X1 U12412 ( .A1(n11633), .A2(n11632), .ZN(n9735) );
  NAND2_X1 U12413 ( .A1(n11169), .A2(n11168), .ZN(n9736) );
  AND2_X1 U12414 ( .A1(n9914), .A2(n9913), .ZN(n9737) );
  INV_X1 U12415 ( .A(n9907), .ZN(n9906) );
  NAND2_X1 U12416 ( .A1(n16411), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9907) );
  AND2_X1 U12417 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n9738) );
  AND2_X1 U12418 ( .A1(n10044), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n9739) );
  NAND2_X1 U12419 ( .A1(n12601), .A2(n12600), .ZN(n9740) );
  INV_X1 U12420 ( .A(n9917), .ZN(n9916) );
  NAND2_X1 U12421 ( .A1(n16408), .A2(n9918), .ZN(n9917) );
  AND2_X1 U12422 ( .A1(n9738), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n9741) );
  INV_X1 U12423 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n9931) );
  INV_X1 U12424 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n9988) );
  INV_X1 U12425 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n9831) );
  INV_X1 U12426 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n9908) );
  INV_X1 U12427 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n9836) );
  INV_X1 U12428 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n9839) );
  OR2_X1 U12429 ( .A1(n9859), .A2(n9858), .ZN(n9742) );
  CLKBUF_X1 U12430 ( .A(n18095), .Z(n9743) );
  NOR3_X1 U12431 ( .A1(n16398), .A2(n18166), .A3(n17349), .ZN(n18095) );
  AOI22_X2 U12432 ( .A1(DATAI_23_), .A2(n13365), .B1(BUF1_REG_23__SCAN_IN), 
        .B2(n13364), .ZN(n20644) );
  AOI22_X2 U12433 ( .A1(DATAI_20_), .A2(n13365), .B1(BUF1_REG_20__SCAN_IN), 
        .B2(n13364), .ZN(n20624) );
  AOI22_X2 U12434 ( .A1(DATAI_17_), .A2(n13365), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n13364), .ZN(n20610) );
  AOI22_X2 U12435 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n13364), .B1(DATAI_22_), 
        .B2(n13365), .ZN(n20636) );
  AOI22_X2 U12436 ( .A1(DATAI_21_), .A2(n13365), .B1(BUF1_REG_21__SCAN_IN), 
        .B2(n13364), .ZN(n20630) );
  AOI22_X2 U12437 ( .A1(DATAI_19_), .A2(n13365), .B1(BUF1_REG_19__SCAN_IN), 
        .B2(n13364), .ZN(n20620) );
  AOI22_X2 U12438 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n19250), .B1(
        BUF2_REG_31__SCAN_IN), .B2(n19249), .ZN(n19751) );
  NOR2_X2 U12439 ( .A1(n15510), .A2(n15509), .ZN(n19249) );
  NOR3_X2 U12440 ( .A1(n18518), .A2(n18493), .A3(n18469), .ZN(n18463) );
  AOI22_X2 U12441 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n13364), .B1(DATAI_16_), 
        .B2(n13365), .ZN(n20604) );
  NAND3_X1 U12442 ( .A1(n12926), .A2(n11950), .A3(n9755), .ZN(n9745) );
  INV_X4 U12443 ( .A(n11836), .ZN(n13340) );
  NAND2_X1 U12444 ( .A1(n9775), .A2(n11836), .ZN(n9774) );
  AND2_X1 U12445 ( .A1(n14515), .A2(n12694), .ZN(n14488) );
  NAND2_X1 U12446 ( .A1(n14535), .A2(n14514), .ZN(n9997) );
  NAND2_X2 U12447 ( .A1(n11916), .A2(n12946), .ZN(n9756) );
  NOR2_X2 U12448 ( .A1(n13745), .A2(n9750), .ZN(n11916) );
  OAI21_X2 U12449 ( .B1(n12751), .B2(n12934), .A(n13760), .ZN(n9750) );
  AOI21_X1 U12450 ( .B1(n9751), .B2(n15808), .A(n9765), .ZN(n9764) );
  NAND2_X1 U12451 ( .A1(n14479), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12695) );
  XNOR2_X1 U12452 ( .A(n12926), .B(n13328), .ZN(n13163) );
  NAND2_X2 U12453 ( .A1(n9766), .A2(n9764), .ZN(n12689) );
  NAND3_X1 U12454 ( .A1(n12687), .A2(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n12686), .ZN(n9766) );
  NAND2_X1 U12455 ( .A1(n13163), .A2(n9755), .ZN(n9767) );
  AND2_X2 U12456 ( .A1(n9768), .A2(n13181), .ZN(n12419) );
  AND2_X2 U12457 ( .A1(n9768), .A2(n11715), .ZN(n11771) );
  AND2_X2 U12458 ( .A1(n9768), .A2(n9976), .ZN(n11754) );
  AND2_X2 U12459 ( .A1(n11707), .A2(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n9768) );
  NAND2_X1 U12460 ( .A1(n15973), .A2(n12655), .ZN(n12657) );
  NAND2_X1 U12461 ( .A1(n9682), .A2(n20106), .ZN(n9770) );
  NAND2_X2 U12462 ( .A1(n15957), .A2(n12678), .ZN(n15956) );
  NAND2_X2 U12463 ( .A1(n12677), .A2(n9994), .ZN(n15957) );
  NAND2_X2 U12464 ( .A1(n13727), .A2(n12675), .ZN(n12677) );
  NAND2_X2 U12465 ( .A1(n12668), .A2(n15965), .ZN(n13727) );
  NAND2_X1 U12466 ( .A1(n9771), .A2(n12698), .ZN(P1_U2968) );
  NAND2_X1 U12467 ( .A1(n14111), .A2(n12697), .ZN(n9771) );
  INV_X1 U12468 ( .A(n11846), .ZN(n9775) );
  AND2_X2 U12469 ( .A1(n9774), .A2(n11858), .ZN(n12538) );
  XNOR2_X2 U12470 ( .A(n10827), .B(n10238), .ZN(n11280) );
  NAND2_X2 U12471 ( .A1(n10272), .A2(n10231), .ZN(n10827) );
  NAND4_X1 U12472 ( .A1(n10155), .A2(n10154), .A3(n10153), .A4(n10152), .ZN(
        n9778) );
  NAND4_X1 U12473 ( .A1(n10151), .A2(n10149), .A3(n10148), .A4(n10150), .ZN(
        n9779) );
  NAND2_X2 U12474 ( .A1(n9782), .A2(n9780), .ZN(n10223) );
  NAND3_X1 U12475 ( .A1(n10203), .A2(n10202), .A3(n19897), .ZN(n9781) );
  NAND2_X1 U12476 ( .A1(n10260), .A2(n12860), .ZN(n10436) );
  OAI21_X2 U12477 ( .B1(n15420), .B2(n9793), .A(n9792), .ZN(n9957) );
  INV_X1 U12478 ( .A(n9957), .ZN(n15381) );
  INV_X2 U12479 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18813) );
  NAND2_X1 U12480 ( .A1(n10466), .A2(n10558), .ZN(n10800) );
  NAND2_X1 U12481 ( .A1(n10223), .A2(n9812), .ZN(n9811) );
  NAND2_X1 U12482 ( .A1(n10210), .A2(n9811), .ZN(n9843) );
  NAND4_X1 U12483 ( .A1(n10340), .A2(n10341), .A3(n10339), .A4(n10338), .ZN(
        n10400) );
  NAND3_X1 U12484 ( .A1(n10293), .A2(n10294), .A3(n10295), .ZN(n10323) );
  NAND3_X1 U12485 ( .A1(n10400), .A2(n9813), .A3(n10323), .ZN(n10463) );
  NAND3_X1 U12486 ( .A1(n10400), .A2(n10323), .A3(n10041), .ZN(n10794) );
  NAND2_X1 U12487 ( .A1(n9822), .A2(n9819), .ZN(n9821) );
  INV_X2 U12488 ( .A(n15129), .ZN(n9817) );
  NAND2_X1 U12489 ( .A1(n9822), .A2(n15086), .ZN(n15122) );
  NAND2_X1 U12490 ( .A1(n9661), .A2(n9835), .ZN(n15739) );
  OR2_X2 U12491 ( .A1(n10211), .A2(n9843), .ZN(n10231) );
  NAND2_X1 U12492 ( .A1(n10211), .A2(n9843), .ZN(n10212) );
  NAND3_X4 U12493 ( .A1(n10255), .A2(n10254), .A3(n10253), .ZN(n10285) );
  AND3_X2 U12494 ( .A1(n13538), .A2(n10799), .A3(n9844), .ZN(n10806) );
  NAND2_X2 U12495 ( .A1(n13540), .A2(n13539), .ZN(n13538) );
  NAND2_X2 U12496 ( .A1(n9851), .A2(n9850), .ZN(n9849) );
  NAND2_X1 U12497 ( .A1(n15065), .A2(n9741), .ZN(n15035) );
  NAND2_X1 U12498 ( .A1(n15021), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n9856) );
  OAI211_X1 U12499 ( .C1(n15021), .C2(n9857), .A(n9856), .B(n9742), .ZN(n14176) );
  NOR2_X1 U12500 ( .A1(n15021), .A2(n9860), .ZN(n11264) );
  NOR2_X1 U12501 ( .A1(n15021), .A2(n15200), .ZN(n15022) );
  NAND2_X1 U12502 ( .A1(n9862), .A2(n13412), .ZN(n13416) );
  NAND3_X1 U12503 ( .A1(n13410), .A2(n9863), .A3(n13423), .ZN(n9862) );
  NAND2_X1 U12504 ( .A1(n13432), .A2(n9864), .ZN(n13621) );
  NAND2_X1 U12505 ( .A1(n13679), .A2(n9718), .ZN(n14845) );
  NAND2_X1 U12506 ( .A1(n14790), .A2(n14791), .ZN(n14793) );
  NOR3_X1 U12507 ( .A1(n14793), .A2(n14784), .A3(n14776), .ZN(n14775) );
  NAND2_X2 U12508 ( .A1(n10257), .A2(n10258), .ZN(n10272) );
  AND2_X2 U12509 ( .A1(n10231), .A2(n10212), .ZN(n10257) );
  INV_X1 U12510 ( .A(n15715), .ZN(n9898) );
  INV_X1 U12511 ( .A(n15711), .ZN(n9899) );
  NAND2_X1 U12512 ( .A1(n9905), .A2(n9663), .ZN(n9910) );
  NAND2_X1 U12513 ( .A1(n17604), .A2(n9698), .ZN(n9901) );
  NAND2_X1 U12514 ( .A1(n17604), .A2(n9677), .ZN(n9911) );
  INV_X1 U12515 ( .A(n17815), .ZN(n9913) );
  INV_X1 U12516 ( .A(n9914), .ZN(n17816) );
  NAND2_X1 U12517 ( .A1(n17510), .A2(n9732), .ZN(n9921) );
  NAND2_X1 U12518 ( .A1(n17511), .A2(n16408), .ZN(n15817) );
  INV_X1 U12519 ( .A(n9921), .ZN(n16335) );
  NAND2_X1 U12520 ( .A1(n17644), .A2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n9928) );
  AOI21_X1 U12521 ( .B1(n17664), .B2(n17587), .A(n9926), .ZN(n9925) );
  NAND3_X1 U12522 ( .A1(n9927), .A2(n17983), .A3(n15716), .ZN(n9926) );
  NAND2_X1 U12523 ( .A1(n13385), .A2(n9936), .ZN(n13713) );
  INV_X1 U12524 ( .A(n13713), .ZN(n10978) );
  INV_X2 U12525 ( .A(n11035), .ZN(n11167) );
  NAND2_X1 U12526 ( .A1(n14903), .A2(n9669), .ZN(n14873) );
  NAND2_X1 U12527 ( .A1(n14903), .A2(n9947), .ZN(n11170) );
  AND2_X1 U12528 ( .A1(n14903), .A2(n14890), .ZN(n14891) );
  AND2_X1 U12529 ( .A1(n14903), .A2(n9948), .ZN(n14875) );
  NOR2_X1 U12530 ( .A1(n10645), .A2(n9959), .ZN(n9958) );
  NAND2_X1 U12531 ( .A1(n9957), .A2(n9949), .ZN(n9956) );
  NAND2_X1 U12532 ( .A1(n9951), .A2(n15264), .ZN(n9950) );
  INV_X1 U12533 ( .A(n9959), .ZN(n9951) );
  NAND2_X1 U12534 ( .A1(n15088), .A2(n9960), .ZN(n9959) );
  NAND2_X1 U12535 ( .A1(n9957), .A2(n9958), .ZN(n9952) );
  NOR2_X1 U12536 ( .A1(n9962), .A2(n9965), .ZN(n10523) );
  INV_X1 U12537 ( .A(n10508), .ZN(n9962) );
  NAND2_X1 U12538 ( .A1(n9963), .A2(n10508), .ZN(n10504) );
  INV_X1 U12539 ( .A(n9965), .ZN(n10513) );
  AND2_X2 U12540 ( .A1(n10622), .A2(n9717), .ZN(n10633) );
  CLKBUF_X1 U12541 ( .A(n9973), .Z(n9970) );
  NOR2_X1 U12542 ( .A1(n10569), .A2(n10568), .ZN(n10591) );
  AND2_X4 U12543 ( .A1(n10311), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11658) );
  NAND3_X1 U12544 ( .A1(n9977), .A2(n14169), .A3(n14168), .ZN(P1_U3000) );
  NAND2_X1 U12545 ( .A1(n14111), .A2(n20160), .ZN(n9977) );
  NAND2_X1 U12546 ( .A1(n20340), .A2(n11949), .ZN(n13209) );
  INV_X1 U12547 ( .A(n11920), .ZN(n9978) );
  NAND2_X1 U12548 ( .A1(n14487), .A2(n14630), .ZN(n14478) );
  OR2_X1 U12549 ( .A1(n13375), .A2(n9998), .ZN(n13376) );
  NAND2_X1 U12550 ( .A1(n9998), .A2(n13375), .ZN(n13373) );
  NOR2_X2 U12551 ( .A1(n13231), .A2(n13371), .ZN(n9998) );
  NOR2_X4 U12552 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11715) );
  AND2_X2 U12553 ( .A1(n13201), .A2(n11715), .ZN(n11737) );
  NAND2_X1 U12554 ( .A1(n11933), .A2(n10002), .ZN(n10000) );
  NAND2_X1 U12555 ( .A1(n11933), .A2(n9755), .ZN(n10001) );
  NAND2_X1 U12556 ( .A1(n11895), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n10003) );
  NOR2_X2 U12557 ( .A1(n13865), .A2(n10006), .ZN(n14337) );
  AND2_X2 U12558 ( .A1(n12344), .A2(n9719), .ZN(n14268) );
  NAND2_X1 U12559 ( .A1(n14241), .A2(n10015), .ZN(n10017) );
  NAND2_X1 U12560 ( .A1(n14241), .A2(n14243), .ZN(n14230) );
  INV_X1 U12561 ( .A(n10017), .ZN(n14231) );
  NAND2_X1 U12562 ( .A1(n11520), .A2(n10021), .ZN(n10019) );
  INV_X1 U12563 ( .A(n10023), .ZN(n14818) );
  NOR2_X1 U12564 ( .A1(n11613), .A2(n11614), .ZN(n14773) );
  NAND2_X1 U12565 ( .A1(n11613), .A2(n14781), .ZN(n10026) );
  NAND2_X1 U12566 ( .A1(n10024), .A2(n10030), .ZN(n14782) );
  NAND2_X1 U12567 ( .A1(n10027), .A2(n10030), .ZN(n14767) );
  INV_X1 U12568 ( .A(n10031), .ZN(n10027) );
  INV_X1 U12569 ( .A(n14768), .ZN(n10029) );
  NOR2_X2 U12570 ( .A1(n14851), .A2(n10033), .ZN(n14824) );
  NOR2_X2 U12571 ( .A1(n13054), .A2(n10037), .ZN(n13221) );
  AND2_X1 U12572 ( .A1(n10323), .A2(n10322), .ZN(n10042) );
  AND2_X1 U12573 ( .A1(n10400), .A2(n10399), .ZN(n10043) );
  NAND2_X4 U12574 ( .A1(n10818), .A2(n10817), .ZN(n15435) );
  AOI21_X1 U12575 ( .B1(n15357), .B2(n15334), .A(n15354), .ZN(n10048) );
  XOR2_X1 U12576 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B(n11264), .Z(
        n15009) );
  INV_X1 U12577 ( .A(n13052), .ZN(n11320) );
  XNOR2_X1 U12578 ( .A(n11919), .B(n11868), .ZN(n11933) );
  OAI21_X2 U12579 ( .B1(n11981), .B2(n14107), .A(n11856), .ZN(n11919) );
  NAND2_X1 U12580 ( .A1(n14176), .A2(n16294), .ZN(n11265) );
  AOI22_X1 U12581 ( .A1(n12604), .A2(n13340), .B1(n11843), .B2(n11790), .ZN(
        n11802) );
  BUF_X4 U12582 ( .A(n11824), .Z(n12459) );
  AOI21_X1 U12583 ( .B1(n12658), .B2(n12194), .A(n12087), .ZN(n13561) );
  NAND2_X1 U12584 ( .A1(n14202), .A2(n10053), .ZN(n14181) );
  NAND2_X2 U12585 ( .A1(n14796), .A2(n11565), .ZN(n11587) );
  AOI21_X1 U12586 ( .B1(n14176), .B2(n16284), .A(n14175), .ZN(n14177) );
  XNOR2_X1 U12587 ( .A(n11968), .B(n12602), .ZN(n13210) );
  INV_X2 U12588 ( .A(n10190), .ZN(n10767) );
  OR2_X1 U12589 ( .A1(n17587), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10051) );
  OR2_X1 U12590 ( .A1(n15644), .A2(n15643), .ZN(n10052) );
  NAND2_X1 U12591 ( .A1(n18233), .A2(n9654), .ZN(n17363) );
  AND2_X1 U12592 ( .A1(n14179), .A2(n9773), .ZN(n10053) );
  INV_X1 U12593 ( .A(n14179), .ZN(n14462) );
  INV_X1 U12594 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15765) );
  INV_X1 U12595 ( .A(n19833), .ZN(n19906) );
  AND2_X1 U12596 ( .A1(n10162), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10055) );
  INV_X1 U12597 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n10598) );
  INV_X1 U12598 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13198) );
  OR3_X1 U12599 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17568), .ZN(n10056) );
  INV_X1 U12600 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n15627) );
  NAND2_X1 U12601 ( .A1(n12024), .A2(n12023), .ZN(n10057) );
  NOR2_X1 U12602 ( .A1(n14390), .A2(n13807), .ZN(n10058) );
  INV_X2 U12603 ( .A(n17226), .ZN(n17220) );
  AND2_X1 U12604 ( .A1(n15119), .A2(n15108), .ZN(n10059) );
  INV_X1 U12605 ( .A(n13359), .ZN(n20178) );
  NAND2_X1 U12606 ( .A1(n9755), .A2(n13333), .ZN(n13359) );
  NOR2_X1 U12607 ( .A1(n11214), .A2(n15006), .ZN(n10060) );
  AND2_X1 U12608 ( .A1(n11368), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(
        n10061) );
  INV_X1 U12609 ( .A(n12215), .ZN(n12194) );
  INV_X1 U12610 ( .A(n13152), .ZN(n13220) );
  INV_X1 U12611 ( .A(n10571), .ZN(n10565) );
  INV_X1 U12612 ( .A(n10448), .ZN(n10377) );
  INV_X1 U12613 ( .A(n12999), .ZN(n20075) );
  OR2_X1 U12614 ( .A1(n10278), .A2(n9657), .ZN(n10062) );
  AND2_X1 U12615 ( .A1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n10063) );
  OR2_X1 U12616 ( .A1(n18891), .A2(n18892), .ZN(n10064) );
  INV_X1 U12617 ( .A(n10929), .ZN(n11093) );
  INV_X1 U12618 ( .A(n11093), .ZN(n11157) );
  AND2_X1 U12619 ( .A1(n20029), .A2(n13649), .ZN(n20014) );
  AND2_X2 U12620 ( .A1(n19918), .A2(n12591), .ZN(n20120) );
  OR2_X1 U12621 ( .A1(n11654), .A2(n11653), .ZN(n10065) );
  AND2_X4 U12622 ( .A1(n13257), .A2(n10147), .ZN(n10066) );
  INV_X1 U12623 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n15828) );
  AND2_X1 U12624 ( .A1(n10285), .A2(n12860), .ZN(n10067) );
  AND4_X1 U12625 ( .A1(n10434), .A2(n10433), .A3(n10432), .A4(n10431), .ZN(
        n10068) );
  INV_X1 U12626 ( .A(n13344), .ZN(n11732) );
  INV_X1 U12627 ( .A(n16267), .ZN(n10573) );
  INV_X1 U12628 ( .A(n12556), .ZN(n12571) );
  NOR2_X1 U12629 ( .A1(n10574), .A2(n10573), .ZN(n10575) );
  INV_X1 U12630 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n11706) );
  OR3_X1 U12631 ( .A1(n12571), .A2(n12570), .A3(n12746), .ZN(n12572) );
  INV_X1 U12632 ( .A(n11937), .ZN(n11914) );
  OAI21_X1 U12633 ( .B1(n15177), .B2(n10576), .A(n10575), .ZN(n10577) );
  AOI21_X1 U12634 ( .B1(n19490), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A(
        n11518), .ZN(n10335) );
  INV_X1 U12635 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11707) );
  OR2_X1 U12636 ( .A1(n12049), .A2(n12048), .ZN(n12650) );
  AOI21_X1 U12637 ( .B1(n12556), .B2(n13734), .A(n12551), .ZN(n12563) );
  OR2_X1 U12638 ( .A1(n11960), .A2(n11959), .ZN(n11961) );
  NAND2_X1 U12639 ( .A1(n10193), .A2(n10180), .ZN(n10170) );
  AOI22_X1 U12640 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n11615), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10129) );
  AOI22_X1 U12641 ( .A1(n10301), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10156), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10085) );
  INV_X1 U12642 ( .A(n12554), .ZN(n12549) );
  AND2_X1 U12643 ( .A1(n12051), .A2(n12050), .ZN(n12057) );
  OR2_X1 U12644 ( .A1(n12068), .A2(n12067), .ZN(n12660) );
  NAND2_X1 U12645 ( .A1(n12543), .A2(n12542), .ZN(n12548) );
  OR2_X1 U12646 ( .A1(n11893), .A2(n11892), .ZN(n12609) );
  OR2_X1 U12647 ( .A1(n13759), .A2(n9755), .ZN(n11988) );
  AND2_X1 U12648 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n11180), .ZN(n10175) );
  AND2_X1 U12649 ( .A1(n12578), .A2(n12577), .ZN(n12748) );
  AOI21_X1 U12650 ( .B1(n12548), .B2(n12547), .A(n12544), .ZN(n12578) );
  AND4_X1 U12651 ( .A1(n11749), .A2(n11748), .A3(n11747), .A4(n11746), .ZN(
        n11750) );
  INV_X1 U12652 ( .A(n12580), .ZN(n12574) );
  INV_X1 U12653 ( .A(n15437), .ZN(n10595) );
  INV_X1 U12654 ( .A(n10802), .ZN(n10556) );
  NAND2_X1 U12655 ( .A1(n11518), .A2(n10321), .ZN(n10322) );
  NAND2_X1 U12656 ( .A1(n10500), .A2(n10499), .ZN(n10728) );
  OAI21_X1 U12657 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18806), .A(
        n13915), .ZN(n13919) );
  INV_X1 U12658 ( .A(n12553), .ZN(n11840) );
  INV_X1 U12659 ( .A(n14325), .ZN(n12343) );
  NOR2_X1 U12660 ( .A1(n13561), .A2(n13570), .ZN(n12101) );
  AND2_X1 U12661 ( .A1(n12474), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12475) );
  NOR2_X1 U12662 ( .A1(n12395), .A2(n12394), .ZN(n12396) );
  INV_X1 U12663 ( .A(n12532), .ZN(n12213) );
  INV_X1 U12664 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12693) );
  OR2_X1 U12665 ( .A1(n13725), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12675) );
  INV_X1 U12666 ( .A(n13535), .ZN(n13431) );
  INV_X1 U12667 ( .A(n11843), .ZN(n11844) );
  AND2_X1 U12668 ( .A1(n12648), .A2(n12580), .ZN(n12576) );
  NOR2_X1 U12669 ( .A1(n10569), .A2(n11687), .ZN(n10605) );
  AND2_X1 U12670 ( .A1(n11587), .A2(n11586), .ZN(n11588) );
  AND2_X1 U12671 ( .A1(n14806), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11288) );
  INV_X1 U12672 ( .A(n14843), .ZN(n11404) );
  INV_X1 U12673 ( .A(n11176), .ZN(n11684) );
  AND2_X1 U12674 ( .A1(n15016), .A2(n15194), .ZN(n10694) );
  AND3_X1 U12675 ( .A1(n10903), .A2(n10902), .A3(n10901), .ZN(n14809) );
  INV_X1 U12676 ( .A(n13224), .ZN(n11322) );
  OAI21_X1 U12677 ( .B1(n10784), .B2(n10506), .A(n13609), .ZN(n10520) );
  NAND2_X1 U12678 ( .A1(n17769), .A2(n18001), .ZN(n15716) );
  INV_X1 U12679 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15712) );
  AND2_X1 U12680 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n15676), .ZN(
        n15692) );
  INV_X1 U12681 ( .A(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n20908) );
  INV_X1 U12682 ( .A(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n20948) );
  NAND2_X1 U12683 ( .A1(n14739), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12497) );
  NAND2_X1 U12684 ( .A1(n12475), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12594) );
  AND2_X1 U12685 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n12369), .ZN(
        n12370) );
  OR2_X1 U12686 ( .A1(n13809), .A2(n14397), .ZN(n13807) );
  AND3_X1 U12687 ( .A1(n12100), .A2(n12099), .A3(n12098), .ZN(n13570) );
  AND2_X1 U12688 ( .A1(n13816), .A2(n13815), .ZN(n13817) );
  AND2_X1 U12689 ( .A1(n13434), .A2(n13433), .ZN(n13435) );
  INV_X1 U12690 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20502) );
  NOR2_X1 U12691 ( .A1(n10504), .A2(n10503), .ZN(n10561) );
  AND3_X1 U12692 ( .A1(n10900), .A2(n10899), .A3(n10898), .ZN(n14815) );
  AND3_X1 U12693 ( .A1(n10870), .A2(n10869), .A3(n10868), .ZN(n13466) );
  AND3_X1 U12694 ( .A1(n10846), .A2(n10845), .A3(n10844), .ZN(n13021) );
  NAND2_X1 U12695 ( .A1(n11304), .A2(n11303), .ZN(n12916) );
  OR2_X1 U12696 ( .A1(n11564), .A2(n11563), .ZN(n11565) );
  INV_X1 U12697 ( .A(n15734), .ZN(n11273) );
  NAND2_X1 U12698 ( .A1(n11215), .A2(n10060), .ZN(n11216) );
  OR3_X1 U12699 ( .A1(n10594), .A2(n10693), .A3(n15442), .ZN(n15437) );
  AND2_X1 U12700 ( .A1(n11191), .A2(n11190), .ZN(n13252) );
  AND3_X1 U12701 ( .A1(n19687), .A2(n19844), .A3(n11308), .ZN(n19579) );
  NOR2_X1 U12702 ( .A1(n16534), .A2(n18846), .ZN(n16538) );
  NOR2_X1 U12703 ( .A1(n17533), .A2(n17534), .ZN(n17521) );
  NOR2_X1 U12704 ( .A1(n17695), .A2(n17697), .ZN(n17672) );
  AND2_X1 U12706 ( .A1(n12219), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12237) );
  INV_X1 U12707 ( .A(n19937), .ZN(n15899) );
  NAND2_X1 U12708 ( .A1(n13648), .A2(n13646), .ZN(n20017) );
  OR2_X2 U12709 ( .A1(n11766), .A2(n11765), .ZN(n11842) );
  AND2_X1 U12710 ( .A1(n14179), .A2(n11844), .ZN(n13862) );
  OAI21_X1 U12711 ( .B1(n12500), .B2(n14540), .A(n12414), .ZN(n14280) );
  NAND2_X1 U12712 ( .A1(n12250), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n12284) );
  AND2_X1 U12713 ( .A1(n12168), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n12201) );
  AND2_X1 U12714 ( .A1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n12004), .ZN(
        n12030) );
  AND2_X1 U12715 ( .A1(n20278), .A2(n20304), .ZN(n20282) );
  OR2_X1 U12716 ( .A1(n20311), .A2(n20552), .ZN(n13479) );
  OR2_X1 U12717 ( .A1(n9655), .A2(n20172), .ZN(n20500) );
  INV_X1 U12718 ( .A(n12612), .ZN(n20172) );
  AND2_X1 U12719 ( .A1(n20436), .A2(n20178), .ZN(n20598) );
  OR2_X1 U12720 ( .A1(n20559), .A2(n20466), .ZN(n20204) );
  NAND2_X1 U12721 ( .A1(n10182), .A2(n15507), .ZN(n10765) );
  OR2_X1 U12722 ( .A1(n19883), .A2(n19888), .ZN(n10758) );
  AND3_X1 U12723 ( .A1(n10879), .A2(n10878), .A3(n10877), .ZN(n13630) );
  AND3_X1 U12724 ( .A1(n10851), .A2(n10850), .A3(n10849), .ZN(n13064) );
  NAND2_X1 U12725 ( .A1(n19110), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19101) );
  INV_X1 U12726 ( .A(n19107), .ZN(n19086) );
  NAND2_X1 U12727 ( .A1(n16315), .A2(n11305), .ZN(n11291) );
  OR2_X1 U12728 ( .A1(n19162), .A2(n11701), .ZN(n12922) );
  INV_X1 U12729 ( .A(n15738), .ZN(n15745) );
  AOI211_X1 U12730 ( .C1(n19122), .C2(n16306), .A(n14170), .B(n11258), .ZN(
        n11262) );
  INV_X1 U12731 ( .A(n15016), .ZN(n15014) );
  OR2_X1 U12732 ( .A1(n16212), .A2(n10676), .ZN(n10677) );
  NAND2_X1 U12733 ( .A1(n10603), .A2(n15409), .ZN(n10604) );
  AND2_X1 U12734 ( .A1(n10813), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15174) );
  INV_X1 U12735 ( .A(n10807), .ZN(n13707) );
  INV_X1 U12736 ( .A(n19847), .ZN(n19548) );
  NAND2_X1 U12737 ( .A1(n19691), .A2(n19697), .ZN(n19650) );
  NAND2_X1 U12738 ( .A1(n19859), .A2(n19870), .ZN(n19847) );
  INV_X1 U12739 ( .A(n19608), .ZN(n19617) );
  NAND2_X1 U12740 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19695), .ZN(n19251) );
  NAND2_X1 U12741 ( .A1(n18204), .A2(n16534), .ZN(n15648) );
  NAND2_X1 U12742 ( .A1(n18677), .A2(n16538), .ZN(n16915) );
  NAND2_X1 U12743 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n17073), .ZN(n17070) );
  NOR2_X1 U12744 ( .A1(n15659), .A2(n15661), .ZN(n18626) );
  NAND2_X1 U12745 ( .A1(n17559), .A2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n17533) );
  NAND2_X1 U12746 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n17639), .ZN(
        n17615) );
  INV_X1 U12747 ( .A(n18004), .ZN(n17924) );
  INV_X1 U12748 ( .A(n17490), .ZN(n17696) );
  NAND2_X1 U12749 ( .A1(n17685), .A2(n17859), .ZN(n17598) );
  AOI21_X1 U12750 ( .B1(n17913), .B2(n17501), .A(n17500), .ZN(n16413) );
  NAND2_X1 U12751 ( .A1(n15718), .A2(n10056), .ZN(n15719) );
  NOR2_X1 U12752 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17769), .ZN(
        n17627) );
  INV_X1 U12753 ( .A(n18052), .ZN(n18031) );
  NOR2_X1 U12754 ( .A1(n17838), .A2(n17837), .ZN(n17836) );
  INV_X1 U12755 ( .A(n14197), .ZN(n13730) );
  INV_X1 U12756 ( .A(n19941), .ZN(n15895) );
  OR2_X1 U12757 ( .A1(n20765), .A2(n13636), .ZN(n20029) );
  INV_X1 U12758 ( .A(n19974), .ZN(n20001) );
  OR2_X1 U12759 ( .A1(n14191), .A2(n13730), .ZN(n13405) );
  INV_X1 U12760 ( .A(n14379), .ZN(n14403) );
  NAND2_X1 U12761 ( .A1(n13118), .A2(n14201), .ZN(n13120) );
  NAND2_X1 U12762 ( .A1(n14179), .A2(n13123), .ZN(n14461) );
  INV_X1 U12763 ( .A(n13077), .ZN(n20101) );
  NAND2_X1 U12764 ( .A1(n12083), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12114) );
  AND2_X1 U12765 ( .A1(n12030), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12053) );
  AND2_X1 U12766 ( .A1(n13762), .A2(n15762), .ZN(n16030) );
  NOR2_X1 U12767 ( .A1(n14127), .A2(n16099), .ZN(n15984) );
  NAND2_X1 U12768 ( .A1(n16055), .A2(n13763), .ZN(n20146) );
  AND2_X1 U12769 ( .A1(n20164), .A2(n20154), .ZN(n16010) );
  INV_X1 U12770 ( .A(n15801), .ZN(n20744) );
  INV_X1 U12771 ( .A(n20267), .ZN(n20237) );
  NAND2_X1 U12772 ( .A1(n20171), .A2(n13235), .ZN(n20275) );
  OAI221_X1 U12773 ( .B1(n20334), .B2(n20379), .C1(n20334), .C2(n20319), .A(
        n20598), .ZN(n20337) );
  INV_X1 U12774 ( .A(n13479), .ZN(n20365) );
  INV_X1 U12775 ( .A(n13511), .ZN(n13366) );
  INV_X1 U12776 ( .A(n20460), .ZN(n20424) );
  INV_X1 U12777 ( .A(n20500), .ZN(n20370) );
  INV_X1 U12778 ( .A(n20485), .ZN(n20496) );
  OAI22_X1 U12779 ( .A1(n20512), .A2(n20511), .B1(n20587), .B2(n20510), .ZN(
        n20547) );
  OR2_X1 U12780 ( .A1(n20171), .A2(n13240), .ZN(n20467) );
  INV_X1 U12781 ( .A(n20503), .ZN(n20591) );
  INV_X1 U12782 ( .A(n20525), .ZN(n20615) );
  INV_X1 U12783 ( .A(n20600), .ZN(n20640) );
  INV_X1 U12784 ( .A(n20521), .ZN(n20646) );
  INV_X1 U12785 ( .A(n20204), .ZN(n20663) );
  INV_X1 U12786 ( .A(P1_STATE_REG_1__SCAN_IN), .ZN(n20674) );
  INV_X1 U12787 ( .A(n20734), .ZN(n20727) );
  INV_X1 U12788 ( .A(n20729), .ZN(n20731) );
  INV_X1 U12789 ( .A(n19650), .ZN(n19844) );
  INV_X1 U12790 ( .A(n19101), .ZN(n19065) );
  INV_X1 U12791 ( .A(n19110), .ZN(n19070) );
  AND2_X1 U12792 ( .A1(n13599), .A2(n13596), .ZN(n19107) );
  INV_X1 U12793 ( .A(n14865), .ZN(n14844) );
  INV_X1 U12794 ( .A(n15002), .ZN(n19164) );
  INV_X1 U12795 ( .A(n13598), .ZN(n19206) );
  INV_X1 U12796 ( .A(n15372), .ZN(n18971) );
  AND2_X1 U12797 ( .A1(n16288), .A2(n12818), .ZN(n16279) );
  INV_X1 U12798 ( .A(n11217), .ZN(n11218) );
  INV_X1 U12799 ( .A(n16310), .ZN(n16296) );
  AND2_X1 U12800 ( .A1(n11194), .A2(n11174), .ZN(n16306) );
  INV_X1 U12801 ( .A(n19210), .ZN(n19877) );
  INV_X1 U12802 ( .A(n19267), .ZN(n19284) );
  AND2_X1 U12803 ( .A1(n19347), .A2(n19548), .ZN(n19337) );
  INV_X1 U12804 ( .A(n19355), .ZN(n19373) );
  AND2_X1 U12805 ( .A1(n19347), .A2(n19617), .ZN(n19389) );
  INV_X1 U12806 ( .A(n19453), .ZN(n19446) );
  OR3_X1 U12807 ( .A1(n19458), .A2(n19614), .A3(n19457), .ZN(n19480) );
  INV_X1 U12808 ( .A(n19513), .ZN(n19506) );
  OAI21_X1 U12809 ( .B1(n19521), .B2(n19536), .A(n19695), .ZN(n19538) );
  NOR2_X1 U12810 ( .A1(n19609), .A2(n19847), .ZN(n19603) );
  INV_X1 U12811 ( .A(n19716), .ZN(n19623) );
  NOR2_X1 U12812 ( .A1(n19646), .A2(n19608), .ZN(n19635) );
  NAND2_X1 U12813 ( .A1(n15479), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16326) );
  INV_X1 U12814 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n19759) );
  INV_X1 U12815 ( .A(n18831), .ZN(n18846) );
  AND2_X1 U12816 ( .A1(n16625), .A2(n16554), .ZN(n16597) );
  NOR2_X1 U12817 ( .A1(n16738), .A2(n16535), .ZN(n16699) );
  NOR2_X1 U12818 ( .A1(n16915), .A2(n16550), .ZN(n16744) );
  INV_X1 U12819 ( .A(n9653), .ZN(n16843) );
  INV_X1 U12820 ( .A(n16912), .ZN(n16889) );
  NAND2_X1 U12821 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17260), .ZN(n17259) );
  NOR2_X1 U12822 ( .A1(n17434), .A2(n17289), .ZN(n17283) );
  NAND2_X1 U12823 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17307), .ZN(n17306) );
  NOR2_X1 U12824 ( .A1(n17474), .A2(n17339), .ZN(n17335) );
  NAND3_X1 U12825 ( .A1(n15614), .A2(n15613), .A3(n15612), .ZN(n16400) );
  NOR2_X1 U12826 ( .A1(n17385), .A2(n17384), .ZN(n17402) );
  NAND2_X1 U12827 ( .A1(n16399), .A2(n16417), .ZN(n17505) );
  NOR2_X1 U12828 ( .A1(n17647), .A2(n17648), .ZN(n17639) );
  NOR2_X1 U12829 ( .A1(n17993), .A2(n17756), .ZN(n17636) );
  INV_X1 U12830 ( .A(n17715), .ZN(n17688) );
  INV_X1 U12831 ( .A(n17773), .ZN(n17725) );
  NOR2_X2 U12832 ( .A1(n17862), .A2(n17349), .ZN(n17770) );
  NOR2_X2 U12833 ( .A1(n18399), .A2(n18446), .ZN(n18571) );
  NOR2_X2 U12834 ( .A1(n18834), .A2(n16516), .ZN(n17852) );
  NAND2_X1 U12835 ( .A1(n18061), .A2(n18635), .ZN(n17996) );
  NOR2_X1 U12836 ( .A1(n18041), .A2(n18166), .ZN(n18081) );
  NOR2_X1 U12837 ( .A1(n18204), .A2(n17996), .ZN(n18054) );
  INV_X1 U12838 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18638) );
  NOR2_X1 U12839 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18782), .ZN(
        n18807) );
  INV_X1 U12840 ( .A(n18675), .ZN(n18827) );
  INV_X1 U12841 ( .A(U212), .ZN(n16466) );
  NAND3_X1 U12842 ( .A1(n14194), .A2(n13730), .A3(n14201), .ZN(n12981) );
  INV_X1 U12843 ( .A(n20034), .ZN(n20008) );
  NAND2_X1 U12844 ( .A1(n20029), .A2(n13655), .ZN(n19942) );
  INV_X1 U12845 ( .A(n20013), .ZN(n20031) );
  INV_X1 U12846 ( .A(n20014), .ZN(n20042) );
  OAI21_X1 U12847 ( .B1(n13405), .B2(n19911), .A(n13404), .ZN(n14384) );
  NAND2_X1 U12848 ( .A1(n14377), .A2(n14192), .ZN(n14405) );
  NAND2_X1 U12849 ( .A1(n13120), .A2(n13119), .ZN(n14179) );
  INV_X1 U12850 ( .A(n14462), .ZN(n14473) );
  INV_X1 U12851 ( .A(n20043), .ZN(n20067) );
  NOR2_X1 U12852 ( .A1(n12981), .A2(n12980), .ZN(n12999) );
  OR2_X1 U12853 ( .A1(n15778), .A2(n19911), .ZN(n19918) );
  OR2_X1 U12854 ( .A1(n20120), .A2(n13115), .ZN(n20130) );
  INV_X1 U12855 ( .A(n20157), .ZN(n20137) );
  INV_X1 U12856 ( .A(n20160), .ZN(n16082) );
  INV_X1 U12857 ( .A(n15761), .ZN(n14107) );
  NAND2_X1 U12858 ( .A1(n20173), .A2(n20370), .ZN(n20235) );
  OR2_X1 U12859 ( .A1(n20275), .A2(n20429), .ZN(n20305) );
  NAND2_X1 U12860 ( .A1(n20312), .A2(n20370), .ZN(n20369) );
  INV_X1 U12861 ( .A(n13331), .ZN(n13370) );
  NAND2_X1 U12862 ( .A1(n20474), .A2(n20370), .ZN(n20428) );
  OR2_X1 U12863 ( .A1(n20467), .A2(n20429), .ZN(n20485) );
  OR2_X1 U12864 ( .A1(n20467), .A2(n20466), .ZN(n20551) );
  OR2_X1 U12865 ( .A1(n20559), .A2(n20552), .ZN(n20600) );
  OR2_X1 U12866 ( .A1(n20559), .A2(n20429), .ZN(n20667) );
  INV_X1 U12867 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n20669) );
  INV_X1 U12868 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n18853) );
  INV_X1 U12869 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19896) );
  INV_X1 U12870 ( .A(n19112), .ZN(n19091) );
  INV_X1 U12871 ( .A(n16215), .ZN(n15253) );
  NAND2_X2 U12872 ( .A1(n12859), .A2(n12858), .ZN(n14856) );
  NAND2_X1 U12873 ( .A1(n12878), .A2(n12877), .ZN(n19210) );
  OR2_X1 U12874 ( .A1(n19162), .A2(n10204), .ZN(n15002) );
  INV_X1 U12875 ( .A(n19162), .ZN(n19152) );
  OR2_X1 U12876 ( .A1(n19162), .A2(n10176), .ZN(n19153) );
  OR2_X1 U12877 ( .A1(n19201), .A2(n12837), .ZN(n19172) );
  NAND2_X1 U12878 ( .A1(n12836), .A2(n19763), .ZN(n19201) );
  NAND2_X1 U12879 ( .A1(n13595), .A2(n11518), .ZN(n13598) );
  OR2_X1 U12880 ( .A1(n18859), .A2(n11518), .ZN(n16259) );
  INV_X1 U12881 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16251) );
  NAND2_X1 U12882 ( .A1(n18859), .A2(n11270), .ZN(n16288) );
  INV_X1 U12883 ( .A(n11235), .ZN(n11236) );
  NAND2_X1 U12884 ( .A1(n11194), .A2(n10824), .ZN(n16312) );
  NAND2_X1 U12885 ( .A1(n19263), .A2(n19347), .ZN(n19267) );
  NAND2_X1 U12886 ( .A1(n19263), .A2(n19425), .ZN(n19316) );
  INV_X1 U12887 ( .A(n19389), .ZN(n19405) );
  INV_X1 U12888 ( .A(n19414), .ZN(n19424) );
  NAND2_X1 U12889 ( .A1(n19347), .A2(n19701), .ZN(n19453) );
  NAND2_X1 U12890 ( .A1(n19701), .A2(n19425), .ZN(n19483) );
  OR2_X1 U12891 ( .A1(n19646), .A2(n19485), .ZN(n19513) );
  OR2_X1 U12892 ( .A1(n19609), .A2(n19485), .ZN(n19541) );
  INV_X1 U12893 ( .A(n19603), .ZN(n19573) );
  INV_X1 U12894 ( .A(n19635), .ZN(n19644) );
  INV_X1 U12895 ( .A(n19731), .ZN(n19674) );
  OR2_X1 U12896 ( .A1(n19646), .A2(n19645), .ZN(n19750) );
  INV_X1 U12897 ( .A(n19843), .ZN(n19758) );
  NAND2_X1 U12898 ( .A1(n18827), .A2(n18632), .ZN(n16516) );
  OR2_X1 U12899 ( .A1(n18699), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18842) );
  NAND2_X1 U12900 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(n16744), .ZN(n16738) );
  INV_X1 U12901 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17720) );
  NAND2_X1 U12902 ( .A1(n16925), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n16912) );
  NOR2_X2 U12903 ( .A1(n17225), .A2(n17074), .ZN(n17226) );
  INV_X1 U12904 ( .A(n17363), .ZN(n17368) );
  INV_X1 U12905 ( .A(n16400), .ZN(n17349) );
  NOR2_X1 U12906 ( .A1(n15558), .A2(n15557), .ZN(n17364) );
  NOR2_X1 U12907 ( .A1(n18679), .A2(n17402), .ZN(n17412) );
  INV_X1 U12908 ( .A(n17402), .ZN(n17422) );
  INV_X1 U12909 ( .A(n17770), .ZN(n17727) );
  INV_X1 U12910 ( .A(n17636), .ZN(n17655) );
  NAND2_X1 U12911 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17856), .ZN(n17715) );
  INV_X1 U12912 ( .A(n17732), .ZN(n17756) );
  OAI21_X1 U12913 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18826), .A(n16516), 
        .ZN(n17859) );
  OR3_X1 U12914 ( .A1(n16417), .A2(n18065), .A3(n17504), .ZN(n16418) );
  NOR2_X1 U12915 ( .A1(n18053), .A2(n17993), .ZN(n18015) );
  INV_X1 U12916 ( .A(n9743), .ZN(n18065) );
  INV_X1 U12917 ( .A(n17768), .ZN(n18100) );
  INV_X1 U12918 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18779) );
  INV_X1 U12919 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18782) );
  INV_X1 U12920 ( .A(n16470), .ZN(n16469) );
  OAI211_X1 U12921 ( .C1(n11279), .C2(n16259), .A(n9685), .B(n11278), .ZN(
        P2_U2985) );
  OAI211_X1 U12922 ( .C1(n15011), .C2(n16310), .A(n11221), .B(n11220), .ZN(
        P2_U3016) );
  AND2_X2 U12923 ( .A1(n10206), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n13300) );
  AND2_X4 U12924 ( .A1(n13300), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10305) );
  NOR2_X2 U12925 ( .A1(n10069), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10296) );
  AND2_X4 U12926 ( .A1(n10296), .A2(n13280), .ZN(n11489) );
  AOI22_X1 U12927 ( .A1(n9649), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11489), .B2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n10073) );
  AOI22_X1 U12928 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11488), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10072) );
  AND2_X4 U12929 ( .A1(n13255), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10301) );
  AND2_X4 U12930 ( .A1(n13257), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10156) );
  AOI22_X1 U12931 ( .A1(n10301), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10156), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n10071) );
  AND2_X4 U12932 ( .A1(n13255), .A2(n10147), .ZN(n10316) );
  AND2_X4 U12933 ( .A1(n13257), .A2(n10147), .ZN(n11615) );
  AOI22_X1 U12934 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11615), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10070) );
  NAND4_X1 U12935 ( .A1(n10073), .A2(n10072), .A3(n10071), .A4(n10070), .ZN(
        n10074) );
  NAND2_X1 U12936 ( .A1(n10074), .A2(n13269), .ZN(n10081) );
  AOI22_X1 U12937 ( .A1(n10305), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_10__6__SCAN_IN), .B2(n11489), .ZN(n10078) );
  AOI22_X1 U12938 ( .A1(n10301), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9632), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10077) );
  AOI22_X1 U12939 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11615), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10076) );
  AOI22_X1 U12940 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11488), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10075) );
  NAND4_X1 U12941 ( .A1(n10078), .A2(n10077), .A3(n10076), .A4(n10075), .ZN(
        n10079) );
  NAND2_X1 U12942 ( .A1(n10079), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10080) );
  INV_X1 U12943 ( .A(n10177), .ZN(n10107) );
  AOI22_X1 U12944 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11488), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10084) );
  AOI22_X1 U12945 ( .A1(n10305), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_10__4__SCAN_IN), .B2(n11489), .ZN(n10083) );
  AOI22_X1 U12946 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n11615), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10082) );
  NAND4_X1 U12947 ( .A1(n10085), .A2(n10084), .A3(n10083), .A4(n10082), .ZN(
        n10086) );
  NAND2_X1 U12948 ( .A1(n10086), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10093) );
  AOI22_X1 U12949 ( .A1(n10301), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n10156), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n10090) );
  AOI22_X1 U12950 ( .A1(n10305), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n11489), .ZN(n10089) );
  AOI22_X1 U12951 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11615), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10088) );
  AOI22_X1 U12952 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n11488), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10087) );
  NAND4_X1 U12953 ( .A1(n10090), .A2(n10089), .A3(n10088), .A4(n10087), .ZN(
        n10091) );
  NAND2_X1 U12954 ( .A1(n10091), .A2(n13269), .ZN(n10092) );
  NAND2_X2 U12955 ( .A1(n10093), .A2(n10092), .ZN(n10759) );
  AOI22_X1 U12956 ( .A1(n10301), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10156), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n10097) );
  AOI22_X1 U12957 ( .A1(n9649), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11489), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n10096) );
  AOI22_X1 U12958 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11488), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10095) );
  AOI22_X1 U12959 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11615), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10094) );
  NAND4_X1 U12960 ( .A1(n10097), .A2(n10096), .A3(n10095), .A4(n10094), .ZN(
        n10098) );
  NAND2_X1 U12961 ( .A1(n10098), .A2(n13269), .ZN(n10105) );
  AOI22_X1 U12962 ( .A1(n10301), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10156), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n10102) );
  AOI22_X1 U12963 ( .A1(n10305), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_10__7__SCAN_IN), .B2(n11489), .ZN(n10101) );
  AOI22_X1 U12964 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n11615), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10100) );
  AOI22_X1 U12965 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11488), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10099) );
  NAND4_X1 U12966 ( .A1(n10102), .A2(n10101), .A3(n10100), .A4(n10099), .ZN(
        n10103) );
  NAND2_X1 U12967 ( .A1(n10103), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10104) );
  NAND2_X2 U12968 ( .A1(n10105), .A2(n10104), .ZN(n10176) );
  NAND2_X1 U12969 ( .A1(n10759), .A2(n10176), .ZN(n10106) );
  OAI21_X1 U12970 ( .B1(n10107), .B2(n10759), .A(n10106), .ZN(n10121) );
  AOI22_X1 U12971 ( .A1(n9649), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11489), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n10111) );
  AOI22_X1 U12972 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11488), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10110) );
  AOI22_X1 U12973 ( .A1(n10301), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9632), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10109) );
  AOI22_X1 U12974 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11615), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10108) );
  NAND4_X1 U12975 ( .A1(n10111), .A2(n10110), .A3(n10109), .A4(n10108), .ZN(
        n10112) );
  NAND2_X1 U12976 ( .A1(n10112), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10119) );
  AOI22_X1 U12977 ( .A1(n10301), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9632), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10116) );
  AOI22_X1 U12978 ( .A1(n10305), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__5__SCAN_IN), .B2(n11489), .ZN(n10115) );
  AOI22_X1 U12979 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11615), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10114) );
  AOI22_X1 U12980 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11488), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10113) );
  NAND4_X1 U12981 ( .A1(n10116), .A2(n10115), .A3(n10114), .A4(n10113), .ZN(
        n10117) );
  NAND2_X1 U12982 ( .A1(n10117), .A2(n13269), .ZN(n10118) );
  NAND2_X2 U12983 ( .A1(n10119), .A2(n10118), .ZN(n10196) );
  NAND2_X1 U12984 ( .A1(n11281), .A2(n10196), .ZN(n10120) );
  NAND2_X1 U12985 ( .A1(n10121), .A2(n10120), .ZN(n10195) );
  INV_X1 U12986 ( .A(n10195), .ZN(n10122) );
  AOI22_X1 U12987 ( .A1(n10301), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9632), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n10126) );
  AOI22_X1 U12988 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11488), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10125) );
  AOI22_X1 U12989 ( .A1(n9649), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11489), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n10124) );
  AOI22_X1 U12990 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11615), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10123) );
  NAND4_X1 U12991 ( .A1(n10126), .A2(n10125), .A3(n10124), .A4(n10123), .ZN(
        n10127) );
  AOI22_X1 U12992 ( .A1(n10301), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9632), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10131) );
  AOI22_X1 U12993 ( .A1(n9649), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11489), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10130) );
  AOI22_X1 U12994 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11488), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10128) );
  NAND4_X1 U12995 ( .A1(n10131), .A2(n10130), .A3(n10129), .A4(n10128), .ZN(
        n10132) );
  NAND2_X1 U12996 ( .A1(n10132), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10133) );
  NAND2_X2 U12997 ( .A1(n10134), .A2(n10133), .ZN(n10190) );
  AOI22_X1 U12998 ( .A1(n10301), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10156), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10138) );
  AOI22_X1 U12999 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11488), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10137) );
  AOI22_X1 U13000 ( .A1(n9649), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11489), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10136) );
  AOI22_X1 U13001 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11615), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10135) );
  NAND4_X1 U13002 ( .A1(n10138), .A2(n10137), .A3(n10136), .A4(n10135), .ZN(
        n10139) );
  NAND2_X1 U13003 ( .A1(n10139), .A2(n13269), .ZN(n10146) );
  AOI22_X1 U13004 ( .A1(n10305), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_10__3__SCAN_IN), .B2(n11489), .ZN(n10142) );
  AOI22_X1 U13005 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11615), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10141) );
  AOI22_X1 U13006 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11488), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10140) );
  NAND4_X1 U13007 ( .A1(n10143), .A2(n10142), .A3(n10141), .A4(n10140), .ZN(
        n10144) );
  NAND2_X1 U13008 ( .A1(n10144), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10145) );
  AND2_X2 U13009 ( .A1(n10146), .A2(n10145), .ZN(n10180) );
  AOI22_X1 U13010 ( .A1(n10301), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10156), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n10151) );
  AOI22_X1 U13011 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11488), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10150) );
  AOI22_X1 U13012 ( .A1(n9649), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11489), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n10149) );
  AOI22_X1 U13013 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n10066), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10148) );
  AOI22_X1 U13014 ( .A1(n10301), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9632), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n10155) );
  AOI22_X1 U13015 ( .A1(n10305), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n11489), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10154) );
  AOI22_X1 U13016 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10066), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10153) );
  AOI22_X1 U13017 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11488), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10152) );
  AOI22_X1 U13018 ( .A1(n10301), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10156), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10161) );
  AOI22_X1 U13019 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n10066), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10159) );
  AOI22_X1 U13020 ( .A1(n10305), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11489), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n10158) );
  AOI22_X1 U13021 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n11488), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10157) );
  NAND2_X1 U13022 ( .A1(n10161), .A2(n10160), .ZN(n10167) );
  AOI22_X1 U13023 ( .A1(n11658), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11488), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10162) );
  AOI22_X1 U13024 ( .A1(n9649), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n11489), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10165) );
  AOI22_X1 U13025 ( .A1(n10316), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10066), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10164) );
  AOI22_X1 U13026 ( .A1(n10301), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10156), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10163) );
  NAND4_X1 U13027 ( .A1(n10055), .A2(n10165), .A3(n10164), .A4(n10163), .ZN(
        n10166) );
  NAND2_X1 U13028 ( .A1(n11684), .A2(n10222), .ZN(n10217) );
  INV_X2 U13029 ( .A(n10759), .ZN(n10200) );
  AND3_X2 U13030 ( .A1(n11189), .A2(n10200), .A3(n10767), .ZN(n10189) );
  NOR2_X2 U13031 ( .A1(n10207), .A2(n11518), .ZN(n10214) );
  AOI22_X1 U13032 ( .A1(n10214), .A2(P2_REIP_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10186) );
  INV_X1 U13033 ( .A(n10207), .ZN(n10169) );
  NAND2_X1 U13034 ( .A1(n10169), .A2(n11518), .ZN(n10184) );
  NAND2_X1 U13035 ( .A1(n12802), .A2(n19884), .ZN(n11178) );
  NOR2_X1 U13036 ( .A1(n10930), .A2(n11189), .ZN(n10171) );
  INV_X1 U13037 ( .A(n10172), .ZN(n10174) );
  AND3_X1 U13038 ( .A1(n10197), .A2(n10176), .A3(n10759), .ZN(n10173) );
  NAND2_X1 U13039 ( .A1(n10925), .A2(n10175), .ZN(n10228) );
  AND2_X2 U13040 ( .A1(n10177), .A2(n10176), .ZN(n10187) );
  NOR2_X1 U13041 ( .A1(n11701), .A2(n10934), .ZN(n10179) );
  NAND2_X1 U13042 ( .A1(n10179), .A2(n11683), .ZN(n10183) );
  NAND4_X2 U13043 ( .A1(n10200), .A2(n10187), .A3(n10180), .A4(n10181), .ZN(
        n12801) );
  INV_X1 U13044 ( .A(n12801), .ZN(n10182) );
  NAND2_X1 U13045 ( .A1(n10183), .A2(n10765), .ZN(n10923) );
  NAND2_X1 U13046 ( .A1(n10923), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10208) );
  NAND3_X1 U13047 ( .A1(n10184), .A2(n10228), .A3(n10208), .ZN(n10213) );
  NAND2_X1 U13048 ( .A1(n10213), .A2(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10185) );
  OAI211_X1 U13049 ( .C1(n10836), .C2(n19103), .A(n10186), .B(n10185), .ZN(
        n10211) );
  NAND2_X1 U13050 ( .A1(n10189), .A2(n10188), .ZN(n10745) );
  NAND2_X1 U13051 ( .A1(n10745), .A2(n10191), .ZN(n10192) );
  NAND2_X1 U13052 ( .A1(n10192), .A2(n10764), .ZN(n11172) );
  OAI21_X1 U13053 ( .B1(n10180), .B2(n10193), .A(n10767), .ZN(n10194) );
  OAI211_X1 U13054 ( .C1(n10195), .C2(n10194), .A(n15507), .B(n12801), .ZN(
        n11184) );
  NAND2_X1 U13055 ( .A1(n10204), .A2(n10759), .ZN(n10766) );
  NAND2_X1 U13056 ( .A1(n10198), .A2(n11281), .ZN(n10199) );
  NAND2_X1 U13057 ( .A1(n10204), .A2(n10199), .ZN(n10769) );
  NAND2_X1 U13058 ( .A1(n10769), .A2(n10200), .ZN(n10761) );
  NAND2_X1 U13059 ( .A1(n10201), .A2(n10761), .ZN(n11182) );
  NAND2_X1 U13060 ( .A1(n11182), .A2(n11189), .ZN(n10203) );
  NAND2_X1 U13061 ( .A1(n11176), .A2(n10180), .ZN(n10202) );
  NAND2_X1 U13062 ( .A1(n11177), .A2(n11176), .ZN(n10205) );
  NAND2_X1 U13063 ( .A1(n18853), .A2(n15828), .ZN(n13251) );
  OAI211_X1 U13064 ( .C1(n13251), .C2(n19873), .A(n10208), .B(n10207), .ZN(
        n10209) );
  INV_X1 U13065 ( .A(n10209), .ZN(n10210) );
  BUF_X2 U13066 ( .A(n10213), .Z(n10837) );
  INV_X1 U13067 ( .A(n10214), .ZN(n10867) );
  INV_X1 U13068 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n14759) );
  NAND2_X1 U13069 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10215) );
  OAI211_X1 U13070 ( .C1(n10867), .C2(n14759), .A(n13251), .B(n10215), .ZN(
        n10216) );
  AOI21_X1 U13071 ( .B1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n10837), .A(
        n10216), .ZN(n10221) );
  INV_X1 U13073 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n10218) );
  NOR2_X1 U13074 ( .A1(n11192), .A2(n10218), .ZN(n10219) );
  OAI21_X1 U13075 ( .B1(n10223), .B2(n10219), .A(P2_STATE2_REG_0__SCAN_IN), 
        .ZN(n10220) );
  NAND2_X1 U13076 ( .A1(n10221), .A2(n10220), .ZN(n10239) );
  INV_X1 U13077 ( .A(n10836), .ZN(n10225) );
  AND2_X1 U13078 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n10224) );
  INV_X1 U13079 ( .A(n13251), .ZN(n10226) );
  NAND2_X1 U13080 ( .A1(n10226), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n10227) );
  AND2_X1 U13081 ( .A1(n10228), .A2(n10227), .ZN(n10229) );
  NAND2_X1 U13082 ( .A1(n10230), .A2(n10229), .ZN(n10240) );
  INV_X1 U13083 ( .A(n10244), .ZN(n10232) );
  NAND2_X1 U13084 ( .A1(n10232), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10234) );
  AOI21_X1 U13085 ( .B1(n18853), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10233) );
  AOI22_X1 U13086 ( .A1(n10214), .A2(P2_REIP_REG_2__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10237) );
  NAND2_X1 U13087 ( .A1(n10837), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10236) );
  INV_X1 U13088 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n10235) );
  NAND3_X1 U13089 ( .A1(n10237), .A2(n10236), .A3(n9692), .ZN(n10247) );
  INV_X1 U13090 ( .A(n10827), .ZN(n10246) );
  INV_X1 U13091 ( .A(n10825), .ZN(n10241) );
  AOI22_X1 U13092 ( .A1(n10214), .A2(P2_REIP_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10242) );
  INV_X1 U13093 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n12918) );
  NAND2_X2 U13094 ( .A1(n10246), .A2(n10245), .ZN(n10255) );
  INV_X1 U13095 ( .A(n10252), .ZN(n10830) );
  NAND2_X1 U13096 ( .A1(n10825), .A2(n10247), .ZN(n10249) );
  INV_X1 U13097 ( .A(n10248), .ZN(n10251) );
  NAND2_X1 U13098 ( .A1(n10252), .A2(n10249), .ZN(n10250) );
  OAI21_X2 U13099 ( .B1(n10252), .B2(n10251), .A(n10250), .ZN(n10253) );
  INV_X1 U13100 ( .A(n10258), .ZN(n10259) );
  XNOR2_X2 U13101 ( .A(n10270), .B(n10259), .ZN(n11297) );
  NAND2_X1 U13102 ( .A1(n10260), .A2(n11297), .ZN(n10435) );
  INV_X1 U13103 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n10261) );
  INV_X1 U13104 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11567) );
  OAI22_X1 U13105 ( .A1(n10435), .A2(n10261), .B1(n10436), .B2(n11567), .ZN(
        n10265) );
  INV_X1 U13106 ( .A(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11040) );
  INV_X1 U13107 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10263) );
  OAI22_X1 U13108 ( .A1(n11040), .A2(n10439), .B1(n10440), .B2(n10263), .ZN(
        n10264) );
  NOR2_X1 U13109 ( .A1(n10265), .A2(n10264), .ZN(n10295) );
  INV_X1 U13110 ( .A(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11574) );
  NAND2_X1 U13111 ( .A1(n10266), .A2(n10267), .ZN(n10420) );
  INV_X1 U13112 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10302) );
  OAI22_X1 U13113 ( .A1(n11574), .A2(n10524), .B1(n10420), .B2(n10302), .ZN(
        n10269) );
  INV_X1 U13114 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11396) );
  INV_X1 U13115 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11388) );
  OAI22_X1 U13116 ( .A1(n11396), .A2(n10421), .B1(n10422), .B2(n11388), .ZN(
        n10268) );
  NOR2_X1 U13117 ( .A1(n10269), .A2(n10268), .ZN(n10294) );
  AND2_X1 U13118 ( .A1(n10270), .A2(n16315), .ZN(n10284) );
  INV_X1 U13119 ( .A(n10284), .ZN(n10271) );
  INV_X1 U13120 ( .A(n10273), .ZN(n10274) );
  NOR2_X1 U13121 ( .A1(n10272), .A2(n10274), .ZN(n10276) );
  INV_X1 U13122 ( .A(n10276), .ZN(n10275) );
  NOR2_X2 U13123 ( .A1(n10283), .A2(n9657), .ZN(n10529) );
  AOI22_X1 U13124 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19381), .B1(
        n10529), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10281) );
  INV_X1 U13125 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11393) );
  INV_X1 U13126 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11041) );
  OAI22_X1 U13127 ( .A1(n11393), .A2(n19689), .B1(n10062), .B2(n11041), .ZN(
        n10279) );
  INV_X1 U13128 ( .A(n10279), .ZN(n10280) );
  NAND3_X1 U13129 ( .A1(n10281), .A2(n10280), .A3(n14806), .ZN(n10292) );
  NOR2_X2 U13130 ( .A1(n10283), .A2(n10277), .ZN(n10429) );
  AOI22_X1 U13131 ( .A1(n10430), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n10429), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10290) );
  INV_X1 U13132 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11387) );
  NAND2_X1 U13133 ( .A1(n10285), .A2(n10284), .ZN(n10286) );
  INV_X1 U13134 ( .A(n10286), .ZN(n10287) );
  INV_X1 U13135 ( .A(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10310) );
  OAI22_X1 U13136 ( .A1(n11387), .A2(n10425), .B1(n10426), .B2(n10310), .ZN(
        n10288) );
  INV_X1 U13137 ( .A(n10288), .ZN(n10289) );
  NAND2_X1 U13138 ( .A1(n10290), .A2(n10289), .ZN(n10291) );
  NOR2_X1 U13139 ( .A1(n10292), .A2(n10291), .ZN(n10293) );
  INV_X1 U13140 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10300) );
  NAND2_X1 U13141 ( .A1(n10156), .A2(n13269), .ZN(n13266) );
  NAND2_X1 U13142 ( .A1(n11464), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10299) );
  NAND2_X1 U13143 ( .A1(n10350), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n10298) );
  OAI211_X1 U13144 ( .C1(n10480), .C2(n10300), .A(n10299), .B(n10298), .ZN(
        n10304) );
  INV_X1 U13145 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11386) );
  OAI22_X1 U13146 ( .A1(n10302), .A2(n11470), .B1(n11469), .B2(n11386), .ZN(
        n10303) );
  NOR2_X1 U13147 ( .A1(n10304), .A2(n10303), .ZN(n10320) );
  AOI22_X1 U13148 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n11473), .B1(
        n11368), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10319) );
  OR2_X2 U13149 ( .A1(n11664), .A2(n13269), .ZN(n11477) );
  NAND3_X1 U13150 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10754) );
  INV_X1 U13151 ( .A(n10754), .ZN(n10306) );
  INV_X1 U13152 ( .A(n10408), .ZN(n10364) );
  AOI22_X1 U13153 ( .A1(n10448), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__3__SCAN_IN), .B2(n10408), .ZN(n10309) );
  NAND2_X1 U13154 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n10308) );
  OAI211_X1 U13155 ( .C1(n11477), .C2(n10310), .A(n10309), .B(n10308), .ZN(
        n10315) );
  NAND2_X1 U13156 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(
        n10313) );
  NAND2_X1 U13157 ( .A1(n11478), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n10312) );
  OAI211_X1 U13158 ( .C1(n10473), .C2(n11388), .A(n10313), .B(n10312), .ZN(
        n10314) );
  NOR2_X1 U13159 ( .A1(n10315), .A2(n10314), .ZN(n10318) );
  AND2_X2 U13160 ( .A1(n11645), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10403) );
  AOI22_X1 U13161 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n11399), .B1(
        n10403), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10317) );
  NAND4_X1 U13162 ( .A1(n10320), .A2(n10319), .A3(n10318), .A4(n10317), .ZN(
        n10966) );
  INV_X1 U13163 ( .A(n10966), .ZN(n10321) );
  NAND2_X1 U13164 ( .A1(n19654), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n10326) );
  NAND2_X1 U13165 ( .A1(n10430), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10325) );
  INV_X1 U13166 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n20805) );
  NAND2_X1 U13167 ( .A1(n19381), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n10324) );
  NAND3_X1 U13168 ( .A1(n10326), .A2(n10325), .A3(n10324), .ZN(n10328) );
  NOR2_X1 U13169 ( .A1(n10328), .A2(n10327), .ZN(n10341) );
  INV_X1 U13170 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11003) );
  INV_X1 U13171 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11345) );
  NAND2_X1 U13172 ( .A1(n10429), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n10329) );
  OAI21_X1 U13173 ( .B1(n10062), .B2(n11003), .A(n10329), .ZN(n10331) );
  INV_X1 U13174 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11352) );
  INV_X1 U13175 ( .A(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10367) );
  NOR2_X1 U13176 ( .A1(n10331), .A2(n10330), .ZN(n10340) );
  NAND2_X1 U13177 ( .A1(n10529), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10336) );
  INV_X1 U13178 ( .A(n10425), .ZN(n19490) );
  NAND2_X1 U13179 ( .A1(n10332), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n10334) );
  INV_X1 U13180 ( .A(n10524), .ZN(n19459) );
  NAND2_X1 U13181 ( .A1(n19459), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10333) );
  INV_X1 U13182 ( .A(n10435), .ZN(n19288) );
  INV_X1 U13183 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n10361) );
  INV_X1 U13184 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11347) );
  OAI22_X1 U13185 ( .A1(n10420), .A2(n10361), .B1(n10422), .B2(n11347), .ZN(
        n10337) );
  AOI21_X1 U13186 ( .B1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n19288), .A(
        n10337), .ZN(n10338) );
  INV_X1 U13187 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10342) );
  INV_X1 U13188 ( .A(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11327) );
  OAI22_X1 U13189 ( .A1(n10480), .A2(n10342), .B1(n11469), .B2(n11327), .ZN(
        n10343) );
  INV_X1 U13190 ( .A(n10343), .ZN(n10349) );
  INV_X1 U13191 ( .A(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10344) );
  INV_X1 U13192 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11491) );
  OAI22_X1 U13193 ( .A1(n11470), .A2(n10344), .B1(n10377), .B2(n11491), .ZN(
        n10345) );
  INV_X1 U13194 ( .A(n10345), .ZN(n10348) );
  AOI22_X1 U13195 ( .A1(n11473), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10408), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10347) );
  AOI22_X1 U13196 ( .A1(n11399), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11464), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n10346) );
  NAND4_X1 U13197 ( .A1(n10349), .A2(n10348), .A3(n10347), .A4(n10346), .ZN(
        n10358) );
  AOI22_X1 U13198 ( .A1(n10350), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10351), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n10356) );
  AOI22_X1 U13199 ( .A1(n11478), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10380), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10355) );
  AOI22_X1 U13200 ( .A1(n11368), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n10403), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n10354) );
  INV_X1 U13201 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10990) );
  INV_X1 U13202 ( .A(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11504) );
  OAI22_X1 U13203 ( .A1(n11477), .A2(n10990), .B1(n10473), .B2(n11504), .ZN(
        n10352) );
  INV_X1 U13204 ( .A(n10352), .ZN(n10353) );
  NAND4_X1 U13205 ( .A1(n10356), .A2(n10355), .A3(n10354), .A4(n10353), .ZN(
        n10357) );
  NOR2_X1 U13206 ( .A1(n10358), .A2(n10357), .ZN(n10939) );
  OR2_X1 U13207 ( .A1(n10939), .A2(n14806), .ZN(n12817) );
  INV_X1 U13208 ( .A(n12817), .ZN(n10376) );
  NAND2_X1 U13209 ( .A1(n11464), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n10360) );
  NAND2_X1 U13210 ( .A1(n10350), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n10359) );
  OAI211_X1 U13211 ( .C1(n10480), .C2(n20805), .A(n10360), .B(n10359), .ZN(
        n10363) );
  OAI22_X1 U13212 ( .A1(n10361), .A2(n11470), .B1(n11469), .B2(n11345), .ZN(
        n10362) );
  NOR2_X1 U13213 ( .A1(n10363), .A2(n10362), .ZN(n10375) );
  AOI22_X1 U13214 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n11473), .B1(
        n11368), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10374) );
  AOI22_X1 U13215 ( .A1(n10448), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n10408), .ZN(n10366) );
  NAND2_X1 U13216 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n10365) );
  OAI211_X1 U13217 ( .C1(n11477), .C2(n10367), .A(n10366), .B(n10365), .ZN(
        n10371) );
  NAND2_X1 U13218 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n10369) );
  NAND2_X1 U13219 ( .A1(n11478), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n10368) );
  OAI211_X1 U13220 ( .C1(n10473), .C2(n11347), .A(n10369), .B(n10368), .ZN(
        n10370) );
  NOR2_X1 U13221 ( .A1(n10371), .A2(n10370), .ZN(n10373) );
  AOI22_X1 U13222 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n11399), .B1(
        n10403), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10372) );
  NAND4_X1 U13223 ( .A1(n10375), .A2(n10374), .A3(n10373), .A4(n10372), .ZN(
        n10950) );
  NAND2_X1 U13224 ( .A1(n10376), .A2(n10950), .ZN(n10788) );
  NAND2_X1 U13225 ( .A1(n11473), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n10398) );
  INV_X1 U13226 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11028) );
  AOI22_X1 U13227 ( .A1(n10448), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__2__SCAN_IN), .B2(n10408), .ZN(n10379) );
  NAND2_X1 U13228 ( .A1(n11478), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n10378) );
  OAI211_X1 U13229 ( .C1(n11477), .C2(n11028), .A(n10379), .B(n10378), .ZN(
        n10384) );
  INV_X1 U13230 ( .A(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11551) );
  NAND2_X1 U13231 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n10382) );
  NAND2_X1 U13232 ( .A1(n10350), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n10381) );
  OAI211_X1 U13233 ( .C1(n10473), .C2(n11551), .A(n10382), .B(n10381), .ZN(
        n10383) );
  NOR2_X1 U13234 ( .A1(n10384), .A2(n10383), .ZN(n10397) );
  INV_X1 U13235 ( .A(n11469), .ZN(n11127) );
  NAND2_X1 U13236 ( .A1(n11127), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(
        n10386) );
  NAND2_X1 U13237 ( .A1(n11399), .A2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n10385) );
  NAND2_X1 U13238 ( .A1(n10386), .A2(n10385), .ZN(n10387) );
  INV_X1 U13239 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n10389) );
  NAND2_X1 U13240 ( .A1(n10403), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n10388) );
  OAI21_X1 U13241 ( .B1(n11470), .B2(n10389), .A(n10388), .ZN(n10394) );
  INV_X1 U13242 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10392) );
  NAND2_X1 U13243 ( .A1(n11464), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(
        n10391) );
  NAND2_X1 U13244 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(
        n10390) );
  OAI211_X1 U13245 ( .C1(n10480), .C2(n10392), .A(n10391), .B(n10390), .ZN(
        n10393) );
  NOR2_X1 U13246 ( .A1(n10394), .A2(n10393), .ZN(n10395) );
  NAND2_X1 U13247 ( .A1(n10788), .A2(n10960), .ZN(n10399) );
  INV_X1 U13248 ( .A(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11068) );
  NAND2_X1 U13249 ( .A1(n11464), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10402) );
  NAND2_X1 U13250 ( .A1(n10350), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10401) );
  OAI211_X1 U13251 ( .C1(n11477), .C2(n11068), .A(n10402), .B(n10401), .ZN(
        n10406) );
  INV_X1 U13252 ( .A(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11408) );
  INV_X1 U13253 ( .A(n10403), .ZN(n10404) );
  INV_X1 U13254 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11407) );
  OAI22_X1 U13255 ( .A1(n11408), .A2(n10404), .B1(n11469), .B2(n11407), .ZN(
        n10405) );
  NOR2_X1 U13256 ( .A1(n10406), .A2(n10405), .ZN(n10419) );
  AOI22_X1 U13257 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n11399), .B1(
        n11368), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10418) );
  INV_X1 U13258 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10411) );
  AOI22_X1 U13259 ( .A1(n10448), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_15__4__SCAN_IN), .B2(n10408), .ZN(n10410) );
  NAND2_X1 U13260 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10409) );
  OAI211_X1 U13261 ( .C1(n10480), .C2(n10411), .A(n10410), .B(n10409), .ZN(
        n10415) );
  INV_X1 U13262 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11599) );
  NAND2_X1 U13263 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n10413) );
  NAND2_X1 U13264 ( .A1(n11478), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10412) );
  OAI211_X1 U13265 ( .C1(n10473), .C2(n11599), .A(n10413), .B(n10412), .ZN(
        n10414) );
  NOR2_X1 U13266 ( .A1(n10415), .A2(n10414), .ZN(n10417) );
  AOI22_X1 U13267 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n11473), .B1(
        n11129), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n10416) );
  NAND4_X1 U13268 ( .A1(n10419), .A2(n10418), .A3(n10417), .A4(n10416), .ZN(
        n10971) );
  INV_X1 U13269 ( .A(n10971), .ZN(n10795) );
  INV_X1 U13270 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11625) );
  INV_X1 U13271 ( .A(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11624) );
  OAI22_X1 U13272 ( .A1(n11625), .A2(n10420), .B1(n10524), .B2(n11624), .ZN(
        n10424) );
  INV_X1 U13273 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11434) );
  INV_X1 U13274 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11427) );
  OAI22_X1 U13275 ( .A1(n11434), .A2(n10421), .B1(n10422), .B2(n11427), .ZN(
        n10423) );
  NOR2_X1 U13276 ( .A1(n10424), .A2(n10423), .ZN(n10434) );
  INV_X1 U13277 ( .A(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11426) );
  INV_X1 U13278 ( .A(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11086) );
  OAI22_X1 U13279 ( .A1(n11426), .A2(n10425), .B1(n10426), .B2(n11086), .ZN(
        n10428) );
  INV_X1 U13280 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11626) );
  OAI22_X1 U13281 ( .A1(n20909), .A2(n19689), .B1(n10062), .B2(n11626), .ZN(
        n10427) );
  NOR2_X1 U13282 ( .A1(n10428), .A2(n10427), .ZN(n10433) );
  AOI22_X1 U13283 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n10529), .B1(
        n19381), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10432) );
  AOI22_X1 U13284 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n10429), .B1(
        n10430), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n10431) );
  INV_X1 U13285 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n10437) );
  INV_X1 U13286 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13020) );
  OAI22_X1 U13287 ( .A1(n10437), .A2(n10435), .B1(n10436), .B2(n13020), .ZN(
        n10438) );
  INV_X1 U13288 ( .A(n10438), .ZN(n10443) );
  INV_X1 U13289 ( .A(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n11079) );
  INV_X1 U13290 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11616) );
  OAI22_X1 U13291 ( .A1(n11079), .A2(n10439), .B1(n10440), .B2(n11616), .ZN(
        n10441) );
  INV_X1 U13292 ( .A(n10441), .ZN(n10442) );
  NAND3_X1 U13293 ( .A1(n10068), .A2(n10443), .A3(n10442), .ZN(n10461) );
  INV_X1 U13294 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11617) );
  NAND2_X1 U13295 ( .A1(n11464), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n10445) );
  NAND2_X1 U13296 ( .A1(n10350), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n10444) );
  OAI211_X1 U13297 ( .C1(n11617), .C2(n10480), .A(n10445), .B(n10444), .ZN(
        n10447) );
  INV_X1 U13298 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11425) );
  OAI22_X1 U13299 ( .A1(n11470), .A2(n11625), .B1(n11469), .B2(n11425), .ZN(
        n10446) );
  NOR2_X1 U13300 ( .A1(n10447), .A2(n10446), .ZN(n10459) );
  AOI22_X1 U13301 ( .A1(n11368), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11473), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10458) );
  INV_X1 U13302 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n20909) );
  NOR2_X1 U13303 ( .A1(n10364), .A2(n20909), .ZN(n10449) );
  AOI21_X1 U13304 ( .B1(n10448), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A(
        n10449), .ZN(n10451) );
  NAND2_X1 U13305 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n10450) );
  OAI211_X1 U13306 ( .C1(n11477), .C2(n11086), .A(n10451), .B(n10450), .ZN(
        n10455) );
  NAND2_X1 U13307 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n10453) );
  NAND2_X1 U13308 ( .A1(n11478), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n10452) );
  OAI211_X1 U13309 ( .C1(n10473), .C2(n11427), .A(n10453), .B(n10452), .ZN(
        n10454) );
  NOR2_X1 U13310 ( .A1(n10455), .A2(n10454), .ZN(n10457) );
  AOI22_X1 U13311 ( .A1(n10407), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10403), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10456) );
  NAND4_X1 U13312 ( .A1(n10459), .A2(n10458), .A3(n10457), .A4(n10456), .ZN(
        n10975) );
  INV_X1 U13313 ( .A(n10975), .ZN(n10502) );
  NAND2_X1 U13314 ( .A1(n11518), .A2(n10502), .ZN(n10460) );
  INV_X1 U13315 ( .A(n10464), .ZN(n10462) );
  NAND2_X1 U13316 ( .A1(n10463), .A2(n10462), .ZN(n10466) );
  NAND2_X1 U13317 ( .A1(n10465), .A2(n10464), .ZN(n10558) );
  NAND2_X1 U13318 ( .A1(n11473), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10470) );
  NAND2_X1 U13319 ( .A1(n11368), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10469) );
  NAND2_X1 U13320 ( .A1(n11399), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10468) );
  NAND2_X1 U13321 ( .A1(n11127), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10467) );
  NAND4_X1 U13322 ( .A1(n10470), .A2(n10469), .A3(n10468), .A4(n10467), .ZN(
        n10479) );
  AOI22_X1 U13323 ( .A1(n10350), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10380), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10477) );
  INV_X1 U13324 ( .A(n11477), .ZN(n11044) );
  NAND2_X1 U13325 ( .A1(n11044), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10476) );
  INV_X1 U13326 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11476) );
  NAND2_X1 U13327 ( .A1(n10448), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10471) );
  OAI21_X1 U13328 ( .B1(n10364), .B2(n11476), .A(n10471), .ZN(n10472) );
  AOI21_X1 U13329 ( .B1(n11478), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n10472), .ZN(n10475) );
  INV_X1 U13330 ( .A(n10473), .ZN(n11047) );
  NAND2_X1 U13331 ( .A1(n11047), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10474) );
  NAND4_X1 U13332 ( .A1(n10477), .A2(n10476), .A3(n10475), .A4(n10474), .ZN(
        n10478) );
  NOR2_X1 U13333 ( .A1(n10479), .A2(n10478), .ZN(n10485) );
  AOI22_X1 U13334 ( .A1(n10403), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11464), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n10483) );
  INV_X1 U13335 ( .A(n10480), .ZN(n11128) );
  AOI22_X1 U13336 ( .A1(n11128), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n10351), .ZN(n10482) );
  NAND2_X1 U13337 ( .A1(n11129), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10481) );
  MUX2_X1 U13338 ( .A(n19873), .B(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n10739) );
  INV_X1 U13339 ( .A(n10716), .ZN(n10486) );
  NAND2_X1 U13340 ( .A1(n10739), .A2(n10486), .ZN(n10488) );
  NAND2_X1 U13341 ( .A1(n19873), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10487) );
  NAND2_X1 U13342 ( .A1(n10488), .A2(n10487), .ZN(n10494) );
  XNOR2_X1 U13343 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n10493) );
  XNOR2_X1 U13344 ( .A(n10494), .B(n10493), .ZN(n10747) );
  NOR2_X1 U13345 ( .A1(n10671), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n10509) );
  INV_X1 U13346 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n19103) );
  NAND2_X1 U13347 ( .A1(n10509), .A2(n19103), .ZN(n10492) );
  NAND2_X1 U13348 ( .A1(n10950), .A2(n10671), .ZN(n10491) );
  NAND2_X1 U13349 ( .A1(n10494), .A2(n10493), .ZN(n10496) );
  NAND2_X1 U13350 ( .A1(n19863), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10495) );
  NAND2_X1 U13351 ( .A1(n10496), .A2(n10495), .ZN(n10498) );
  XNOR2_X1 U13352 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10497) );
  XNOR2_X1 U13353 ( .A(n10498), .B(n10497), .ZN(n10748) );
  INV_X1 U13354 ( .A(n10748), .ZN(n10723) );
  MUX2_X1 U13355 ( .A(n10966), .B(n10723), .S(n19884), .Z(n10714) );
  MUX2_X1 U13356 ( .A(n10714), .B(n12918), .S(n11687), .Z(n10508) );
  NAND2_X1 U13357 ( .A1(n10498), .A2(n10497), .ZN(n10500) );
  NAND2_X1 U13358 ( .A1(n19856), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10499) );
  NAND2_X1 U13359 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n20796), .ZN(
        n10727) );
  INV_X1 U13360 ( .A(n10746), .ZN(n10501) );
  MUX2_X1 U13361 ( .A(n10971), .B(n10501), .S(n19884), .Z(n10713) );
  INV_X1 U13362 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n19084) );
  MUX2_X1 U13363 ( .A(n10713), .B(n19084), .S(n11687), .Z(n10522) );
  MUX2_X1 U13364 ( .A(P2_EBX_REG_5__SCAN_IN), .B(n10502), .S(n10671), .Z(
        n10503) );
  AND2_X1 U13365 ( .A1(n10504), .A2(n10503), .ZN(n10505) );
  OR2_X1 U13366 ( .A1(n10505), .A2(n10561), .ZN(n19067) );
  INV_X1 U13367 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13717) );
  INV_X1 U13368 ( .A(n10693), .ZN(n10506) );
  INV_X1 U13369 ( .A(n10523), .ZN(n10507) );
  OAI21_X1 U13370 ( .B1(n10513), .B2(n10508), .A(n10507), .ZN(n13609) );
  NAND2_X1 U13371 ( .A1(n10520), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13380) );
  OAI21_X1 U13372 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19880), .A(
        n10716), .ZN(n10718) );
  MUX2_X1 U13373 ( .A(n10718), .B(n10939), .S(n10731), .Z(n10510) );
  AOI21_X1 U13374 ( .B1(n10510), .B2(n10671), .A(n10509), .ZN(n14763) );
  NAND2_X1 U13375 ( .A1(n14763), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12825) );
  NAND3_X1 U13376 ( .A1(n11687), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n10511) );
  NAND2_X1 U13377 ( .A1(n10514), .A2(n10511), .ZN(n19100) );
  NOR2_X1 U13378 ( .A1(n12825), .A2(n19100), .ZN(n10512) );
  NAND2_X1 U13379 ( .A1(n12825), .A2(n19100), .ZN(n12824) );
  OAI21_X1 U13380 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10512), .A(
        n12824), .ZN(n12724) );
  NAND2_X1 U13381 ( .A1(n10515), .A2(n10514), .ZN(n10516) );
  NAND2_X1 U13382 ( .A1(n9965), .A2(n10516), .ZN(n13673) );
  INV_X1 U13383 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n12721) );
  XNOR2_X1 U13384 ( .A(n13673), .B(n12721), .ZN(n12723) );
  OR2_X1 U13385 ( .A1(n12724), .A2(n12723), .ZN(n12807) );
  INV_X1 U13386 ( .A(n13673), .ZN(n10517) );
  NAND2_X1 U13387 ( .A1(n10517), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10518) );
  NAND2_X1 U13388 ( .A1(n12807), .A2(n10518), .ZN(n13382) );
  INV_X1 U13389 ( .A(n13382), .ZN(n10519) );
  NAND2_X1 U13390 ( .A1(n13380), .A2(n10519), .ZN(n10521) );
  OR2_X1 U13391 ( .A1(n10520), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13381) );
  NAND2_X1 U13392 ( .A1(n10521), .A2(n13381), .ZN(n13543) );
  XNOR2_X1 U13393 ( .A(n10523), .B(n10522), .ZN(n19087) );
  INV_X1 U13394 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13539) );
  XNOR2_X1 U13395 ( .A(n19087), .B(n13539), .ZN(n13542) );
  NAND2_X1 U13396 ( .A1(n13710), .A2(n13711), .ZN(n15176) );
  INV_X1 U13397 ( .A(n10558), .ZN(n10557) );
  INV_X1 U13398 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n10540) );
  INV_X1 U13399 ( .A(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11447) );
  OAI22_X1 U13400 ( .A1(n10540), .A2(n10420), .B1(n10524), .B2(n11447), .ZN(
        n10526) );
  INV_X1 U13401 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11456) );
  INV_X1 U13402 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11638) );
  OAI22_X1 U13403 ( .A1(n11456), .A2(n10421), .B1(n10422), .B2(n11638), .ZN(
        n10525) );
  NOR2_X1 U13404 ( .A1(n10526), .A2(n10525), .ZN(n10533) );
  INV_X1 U13405 ( .A(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11444) );
  INV_X1 U13406 ( .A(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11107) );
  OAI22_X1 U13407 ( .A1(n11444), .A2(n10425), .B1(n10426), .B2(n11107), .ZN(
        n10528) );
  INV_X1 U13408 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11453) );
  INV_X1 U13409 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11100) );
  OAI22_X1 U13410 ( .A1(n11453), .A2(n19689), .B1(n10062), .B2(n11100), .ZN(
        n10527) );
  NOR2_X1 U13411 ( .A1(n10528), .A2(n10527), .ZN(n10532) );
  AOI22_X1 U13412 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10429), .B1(
        n10430), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n10531) );
  AOI22_X1 U13413 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10529), .B1(
        n19381), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10530) );
  NAND4_X1 U13414 ( .A1(n10533), .A2(n10532), .A3(n10531), .A4(n10530), .ZN(
        n10537) );
  INV_X1 U13415 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11640) );
  INV_X1 U13416 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11639) );
  OAI22_X1 U13417 ( .A1(n11640), .A2(n10435), .B1(n10436), .B2(n11639), .ZN(
        n10536) );
  INV_X1 U13418 ( .A(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n11099) );
  INV_X1 U13419 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10534) );
  OAI22_X1 U13420 ( .A1(n11099), .A2(n10439), .B1(n10440), .B2(n10534), .ZN(
        n10535) );
  INV_X1 U13421 ( .A(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n11642) );
  NAND2_X1 U13422 ( .A1(n11464), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n10539) );
  NAND2_X1 U13423 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n10538) );
  OAI211_X1 U13424 ( .C1(n11642), .C2(n10480), .A(n10539), .B(n10538), .ZN(
        n10542) );
  INV_X1 U13425 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11443) );
  OAI22_X1 U13426 ( .A1(n11470), .A2(n10540), .B1(n11469), .B2(n11443), .ZN(
        n10541) );
  NOR2_X1 U13427 ( .A1(n10542), .A2(n10541), .ZN(n10552) );
  AOI22_X1 U13428 ( .A1(n11368), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11473), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10551) );
  AOI22_X1 U13429 ( .A1(n10448), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n10408), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n10544) );
  NAND2_X1 U13430 ( .A1(n11478), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n10543) );
  OAI211_X1 U13431 ( .C1(n11477), .C2(n11107), .A(n10544), .B(n10543), .ZN(
        n10548) );
  NAND2_X1 U13432 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n10546) );
  NAND2_X1 U13433 ( .A1(n10350), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n10545) );
  OAI211_X1 U13434 ( .C1(n10473), .C2(n11638), .A(n10546), .B(n10545), .ZN(
        n10547) );
  NOR2_X1 U13435 ( .A1(n10548), .A2(n10547), .ZN(n10550) );
  AOI22_X1 U13436 ( .A1(n10407), .A2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n10403), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10549) );
  NAND4_X1 U13437 ( .A1(n10552), .A2(n10551), .A3(n10550), .A4(n10549), .ZN(
        n10979) );
  INV_X1 U13438 ( .A(n10979), .ZN(n10553) );
  NAND2_X1 U13439 ( .A1(n11518), .A2(n10553), .ZN(n10554) );
  NAND2_X1 U13440 ( .A1(n10558), .A2(n10802), .ZN(n10559) );
  NAND2_X1 U13441 ( .A1(n10809), .A2(n10693), .ZN(n10563) );
  MUX2_X1 U13442 ( .A(n13023), .B(n10979), .S(n10934), .Z(n10560) );
  OR2_X1 U13443 ( .A1(n10561), .A2(n10560), .ZN(n10562) );
  NAND2_X1 U13444 ( .A1(n10572), .A2(n10562), .ZN(n19053) );
  NOR2_X1 U13445 ( .A1(n15178), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10581) );
  INV_X1 U13446 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n10576) );
  MUX2_X1 U13447 ( .A(P2_EBX_REG_7__SCAN_IN), .B(n10693), .S(n10671), .Z(
        n10571) );
  INV_X1 U13448 ( .A(P2_EBX_REG_8__SCAN_IN), .ZN(n10567) );
  NOR2_X1 U13449 ( .A1(n10671), .A2(n10567), .ZN(n10568) );
  AND2_X1 U13450 ( .A1(n10569), .A2(n10568), .ZN(n10570) );
  OR2_X1 U13451 ( .A1(n10570), .A2(n10591), .ZN(n19032) );
  NOR2_X1 U13452 ( .A1(n19032), .A2(n10693), .ZN(n10582) );
  NAND2_X1 U13453 ( .A1(n10582), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16271) );
  INV_X1 U13454 ( .A(n16271), .ZN(n10574) );
  XNOR2_X1 U13455 ( .A(n10572), .B(n10565), .ZN(n19041) );
  NAND2_X1 U13456 ( .A1(n19041), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16267) );
  INV_X1 U13457 ( .A(n10577), .ZN(n10580) );
  NAND2_X1 U13458 ( .A1(n15177), .A2(n10576), .ZN(n10578) );
  NAND2_X1 U13459 ( .A1(n10578), .A2(n15178), .ZN(n10579) );
  OAI211_X1 U13460 ( .C1(n15176), .C2(n10581), .A(n10580), .B(n10579), .ZN(
        n10587) );
  INV_X1 U13461 ( .A(n10582), .ZN(n10584) );
  INV_X1 U13462 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10583) );
  NAND2_X1 U13463 ( .A1(n10584), .A2(n10583), .ZN(n16270) );
  INV_X1 U13464 ( .A(n19041), .ZN(n10585) );
  INV_X1 U13465 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15454) );
  NAND2_X1 U13466 ( .A1(n10585), .A2(n15454), .ZN(n16266) );
  AND2_X1 U13467 ( .A1(n16270), .A2(n16266), .ZN(n10586) );
  NAND2_X1 U13468 ( .A1(n10587), .A2(n10586), .ZN(n15436) );
  INV_X1 U13469 ( .A(n15436), .ZN(n10590) );
  INV_X1 U13470 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n13060) );
  NOR2_X1 U13471 ( .A1(n10671), .A2(n13060), .ZN(n10588) );
  XNOR2_X1 U13472 ( .A(n10591), .B(n10588), .ZN(n19020) );
  AOI21_X1 U13473 ( .B1(n19020), .B2(n10506), .A(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15438) );
  INV_X1 U13474 ( .A(n15438), .ZN(n10589) );
  NAND2_X1 U13475 ( .A1(n10590), .A2(n10589), .ZN(n15420) );
  NAND3_X1 U13476 ( .A1(n10597), .A2(P2_EBX_REG_10__SCAN_IN), .A3(n11687), 
        .ZN(n10592) );
  OAI211_X1 U13477 ( .C1(n10597), .C2(P2_EBX_REG_10__SCAN_IN), .A(n10592), .B(
        n10685), .ZN(n19009) );
  OR2_X1 U13478 ( .A1(n19009), .A2(n10693), .ZN(n10593) );
  INV_X1 U13479 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15419) );
  AND2_X1 U13480 ( .A1(n10593), .A2(n15419), .ZN(n15421) );
  INV_X1 U13481 ( .A(n19020), .ZN(n10594) );
  INV_X1 U13482 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15442) );
  NOR2_X2 U13483 ( .A1(n10599), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10607) );
  NAND2_X1 U13484 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n10599), .ZN(n10600) );
  NOR2_X1 U13485 ( .A1(n10934), .A2(n10600), .ZN(n10601) );
  OR2_X1 U13486 ( .A1(n10607), .A2(n10601), .ZN(n18998) );
  OR2_X1 U13487 ( .A1(n10605), .A2(n10693), .ZN(n10602) );
  INV_X1 U13488 ( .A(n15406), .ZN(n10603) );
  INV_X1 U13489 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15409) );
  NAND2_X1 U13490 ( .A1(n11687), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10606) );
  OR2_X1 U13491 ( .A1(n10607), .A2(n10606), .ZN(n10608) );
  NAND2_X1 U13492 ( .A1(n10630), .A2(n10608), .ZN(n18990) );
  INV_X1 U13493 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n20933) );
  OAI21_X1 U13494 ( .B1(n18990), .B2(n10693), .A(n20933), .ZN(n15391) );
  NOR3_X1 U13495 ( .A1(n18990), .A2(n10693), .A3(n20933), .ZN(n15392) );
  INV_X1 U13496 ( .A(P2_EBX_REG_13__SCAN_IN), .ZN(n10609) );
  NOR2_X1 U13497 ( .A1(n10671), .A2(n10609), .ZN(n10629) );
  NAND2_X1 U13498 ( .A1(n11687), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10624) );
  AND2_X2 U13499 ( .A1(n10626), .A2(n10624), .ZN(n10618) );
  INV_X1 U13500 ( .A(P2_EBX_REG_16__SCAN_IN), .ZN(n10610) );
  NAND2_X1 U13501 ( .A1(n10618), .A2(n10610), .ZN(n10616) );
  NAND2_X2 U13502 ( .A1(n10616), .A2(n10685), .ZN(n10622) );
  NAND2_X1 U13503 ( .A1(n11687), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10621) );
  NOR2_X1 U13504 ( .A1(P2_EBX_REG_19__SCAN_IN), .A2(P2_EBX_REG_18__SCAN_IN), 
        .ZN(n10611) );
  NOR2_X1 U13505 ( .A1(n10671), .A2(n10611), .ZN(n10612) );
  INV_X1 U13506 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n10613) );
  NAND2_X1 U13507 ( .A1(n10633), .A2(n10613), .ZN(n10667) );
  INV_X1 U13508 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15260) );
  NAND2_X1 U13509 ( .A1(n11687), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10617) );
  OAI211_X1 U13510 ( .C1(n10618), .C2(n10617), .A(n10685), .B(n10616), .ZN(
        n18942) );
  OR2_X1 U13511 ( .A1(n18942), .A2(n10693), .ZN(n10619) );
  XNOR2_X1 U13512 ( .A(n10619), .B(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15140) );
  OR2_X1 U13513 ( .A1(n10622), .A2(n10621), .ZN(n10623) );
  AND2_X1 U13514 ( .A1(n10620), .A2(n10623), .ZN(n18927) );
  NAND2_X1 U13515 ( .A1(n18927), .A2(n10506), .ZN(n10653) );
  INV_X1 U13516 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n10819) );
  NAND2_X1 U13517 ( .A1(n10653), .A2(n10819), .ZN(n15085) );
  INV_X1 U13518 ( .A(n10624), .ZN(n10625) );
  XNOR2_X1 U13519 ( .A(n10626), .B(n10625), .ZN(n18954) );
  NAND2_X1 U13520 ( .A1(n18954), .A2(n10506), .ZN(n10627) );
  INV_X1 U13521 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15357) );
  NAND2_X1 U13522 ( .A1(n10627), .A2(n15357), .ZN(n15152) );
  XNOR2_X1 U13523 ( .A(n9660), .B(n9723), .ZN(n18968) );
  NAND2_X1 U13524 ( .A1(n18968), .A2(n10506), .ZN(n10628) );
  INV_X1 U13525 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n15367) );
  NAND2_X1 U13526 ( .A1(n10628), .A2(n15367), .ZN(n15163) );
  AND2_X1 U13527 ( .A1(n10630), .A2(n10629), .ZN(n10631) );
  OR2_X1 U13528 ( .A1(n10631), .A2(n9660), .ZN(n18976) );
  INV_X1 U13529 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n10650) );
  OAI21_X1 U13530 ( .B1(n18976), .B2(n10693), .A(n10650), .ZN(n15380) );
  AND4_X1 U13531 ( .A1(n15085), .A2(n15152), .A3(n15163), .A4(n15380), .ZN(
        n10632) );
  INV_X1 U13532 ( .A(n10633), .ZN(n10636) );
  NAND2_X1 U13533 ( .A1(n9681), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10634) );
  MUX2_X1 U13534 ( .A(n10634), .B(n9681), .S(n10671), .Z(n10635) );
  NAND2_X1 U13535 ( .A1(n10636), .A2(n10635), .ZN(n18898) );
  NOR2_X1 U13536 ( .A1(n18898), .A2(n10693), .ZN(n10656) );
  NOR2_X1 U13537 ( .A1(n10656), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15097) );
  NAND2_X1 U13538 ( .A1(n10620), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10637) );
  MUX2_X1 U13539 ( .A(n10620), .B(n10637), .S(n11687), .Z(n10638) );
  OR2_X1 U13540 ( .A1(n10620), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10641) );
  AND2_X1 U13541 ( .A1(n10638), .A2(n10641), .ZN(n18918) );
  NAND2_X1 U13542 ( .A1(n18918), .A2(n10506), .ZN(n10657) );
  INV_X1 U13543 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15317) );
  NAND2_X1 U13544 ( .A1(n10657), .A2(n15317), .ZN(n15119) );
  INV_X1 U13545 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n10639) );
  NOR2_X1 U13546 ( .A1(n10934), .A2(n10639), .ZN(n10640) );
  NAND2_X1 U13547 ( .A1(n10641), .A2(n10640), .ZN(n10642) );
  NAND2_X1 U13548 ( .A1(n10642), .A2(n9681), .ZN(n18905) );
  OR2_X1 U13549 ( .A1(n18905), .A2(n10693), .ZN(n10643) );
  INV_X1 U13550 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15293) );
  NAND2_X1 U13551 ( .A1(n10643), .A2(n15293), .ZN(n15108) );
  OR2_X1 U13552 ( .A1(n10693), .A2(n15260), .ZN(n10646) );
  OR2_X1 U13553 ( .A1(n18881), .A2(n10646), .ZN(n15087) );
  INV_X1 U13554 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15352) );
  OR2_X1 U13555 ( .A1(n10693), .A2(n15352), .ZN(n10647) );
  OR2_X1 U13556 ( .A1(n18942), .A2(n10647), .ZN(n15084) );
  NOR2_X1 U13557 ( .A1(n10693), .A2(n15357), .ZN(n10648) );
  NAND2_X1 U13558 ( .A1(n18954), .A2(n10648), .ZN(n15151) );
  NOR2_X1 U13559 ( .A1(n10693), .A2(n15367), .ZN(n10649) );
  NAND2_X1 U13560 ( .A1(n18968), .A2(n10649), .ZN(n15162) );
  INV_X1 U13561 ( .A(n18976), .ZN(n10652) );
  NOR2_X1 U13562 ( .A1(n10693), .A2(n10650), .ZN(n10651) );
  NAND2_X1 U13563 ( .A1(n10652), .A2(n10651), .ZN(n15379) );
  AND4_X1 U13564 ( .A1(n15084), .A2(n15151), .A3(n15162), .A4(n15379), .ZN(
        n10655) );
  INV_X1 U13565 ( .A(n10653), .ZN(n10654) );
  NAND2_X1 U13566 ( .A1(n10654), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15086) );
  NAND3_X1 U13567 ( .A1(n15087), .A2(n10655), .A3(n15086), .ZN(n10662) );
  INV_X1 U13568 ( .A(n15099), .ZN(n10660) );
  INV_X1 U13569 ( .A(n10657), .ZN(n10658) );
  NAND2_X1 U13570 ( .A1(n10658), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15120) );
  OR2_X1 U13571 ( .A1(n10693), .A2(n15293), .ZN(n10659) );
  OR2_X1 U13572 ( .A1(n18905), .A2(n10659), .ZN(n15107) );
  NAND2_X1 U13573 ( .A1(n10660), .A2(n9715), .ZN(n10661) );
  NAND2_X1 U13574 ( .A1(n11687), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10664) );
  INV_X1 U13575 ( .A(n10664), .ZN(n10668) );
  INV_X1 U13576 ( .A(n10673), .ZN(n10666) );
  AOI21_X1 U13577 ( .B1(n10668), .B2(n10667), .A(n10666), .ZN(n15728) );
  NAND2_X1 U13578 ( .A1(n15728), .A2(n10506), .ZN(n10669) );
  INV_X1 U13579 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15270) );
  NAND2_X1 U13580 ( .A1(n10669), .A2(n15270), .ZN(n15264) );
  INV_X1 U13581 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n10670) );
  NOR2_X1 U13582 ( .A1(n10671), .A2(n10670), .ZN(n10672) );
  NAND2_X1 U13583 ( .A1(n10673), .A2(n10672), .ZN(n10674) );
  NAND2_X1 U13584 ( .A1(n9673), .A2(n10674), .ZN(n16212) );
  OR2_X1 U13585 ( .A1(n16212), .A2(n10693), .ZN(n10675) );
  INV_X1 U13586 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15249) );
  XNOR2_X1 U13587 ( .A(n10675), .B(n15249), .ZN(n15074) );
  NAND2_X1 U13588 ( .A1(n10506), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10676) );
  NAND2_X1 U13589 ( .A1(n11687), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10678) );
  MUX2_X1 U13590 ( .A(P2_EBX_REG_24__SCAN_IN), .B(n10678), .S(n9673), .Z(
        n10679) );
  NAND2_X1 U13591 ( .A1(n10679), .A2(n10685), .ZN(n16198) );
  NOR2_X1 U13592 ( .A1(n16198), .A2(n10693), .ZN(n15062) );
  INV_X1 U13593 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n10683) );
  NOR2_X1 U13594 ( .A1(n10684), .A2(n10683), .ZN(n10680) );
  NAND2_X1 U13595 ( .A1(n11687), .A2(n10680), .ZN(n10681) );
  NAND2_X1 U13596 ( .A1(n10685), .A2(n10681), .ZN(n10682) );
  AOI21_X1 U13597 ( .B1(n10684), .B2(n10683), .A(n10682), .ZN(n16187) );
  NAND2_X1 U13598 ( .A1(n10684), .A2(n10683), .ZN(n10686) );
  INV_X1 U13599 ( .A(n10689), .ZN(n11243) );
  NAND3_X1 U13600 ( .A1(n11687), .A2(P2_EBX_REG_26__SCAN_IN), .A3(n10686), 
        .ZN(n10687) );
  AND3_X2 U13601 ( .A1(n16177), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n10506), .ZN(n10700) );
  AOI21_X1 U13602 ( .B1(n16177), .B2(n10506), .A(
        P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10688) );
  NOR2_X1 U13603 ( .A1(n10700), .A2(n10688), .ZN(n15040) );
  NAND2_X1 U13604 ( .A1(n11687), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10690) );
  INV_X1 U13605 ( .A(n10690), .ZN(n10691) );
  NAND2_X1 U13606 ( .A1(n10691), .A2(n9676), .ZN(n10692) );
  NAND2_X1 U13607 ( .A1(n10704), .A2(n10692), .ZN(n16167) );
  INV_X1 U13608 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n15194) );
  NOR2_X1 U13609 ( .A1(n15013), .A2(n10694), .ZN(n10697) );
  INV_X1 U13610 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15200) );
  NAND2_X1 U13611 ( .A1(n11687), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n10702) );
  XOR2_X1 U13612 ( .A(n10702), .B(n10704), .Z(n16153) );
  INV_X1 U13613 ( .A(n15018), .ZN(n10695) );
  AOI21_X1 U13614 ( .B1(n15200), .B2(n15194), .A(n10695), .ZN(n10696) );
  OAI22_X1 U13615 ( .A1(n10697), .A2(n10696), .B1(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n15018), .ZN(n10701) );
  INV_X1 U13616 ( .A(n10698), .ZN(n10699) );
  INV_X1 U13617 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15233) );
  NOR2_X1 U13618 ( .A1(n15052), .A2(n10700), .ZN(n15012) );
  NAND2_X1 U13619 ( .A1(n10701), .A2(n15012), .ZN(n11223) );
  INV_X1 U13620 ( .A(n10702), .ZN(n10703) );
  NAND2_X1 U13621 ( .A1(n11687), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n10706) );
  XNOR2_X1 U13622 ( .A(n10707), .B(n10706), .ZN(n10705) );
  INV_X1 U13623 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11232) );
  OAI21_X1 U13624 ( .B1(n10705), .B2(n10693), .A(n11232), .ZN(n11222) );
  NAND2_X1 U13625 ( .A1(n11223), .A2(n11222), .ZN(n11240) );
  INV_X1 U13626 ( .A(n10705), .ZN(n16143) );
  NAND3_X1 U13627 ( .A1(n16143), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n10506), .ZN(n11237) );
  NAND2_X1 U13628 ( .A1(n11240), .A2(n11237), .ZN(n10712) );
  NAND2_X1 U13629 ( .A1(n10707), .A2(n10706), .ZN(n11241) );
  NAND2_X1 U13630 ( .A1(n11687), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n10708) );
  XNOR2_X1 U13631 ( .A(n11241), .B(n10708), .ZN(n10709) );
  AOI21_X1 U13632 ( .B1(n10709), .B2(n10506), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11239) );
  INV_X1 U13633 ( .A(n10709), .ZN(n16133) );
  INV_X1 U13634 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n11257) );
  INV_X1 U13635 ( .A(n11238), .ZN(n10710) );
  NOR2_X1 U13636 ( .A1(n11239), .A2(n10710), .ZN(n10711) );
  XNOR2_X1 U13637 ( .A(n10712), .B(n10711), .ZN(n15011) );
  NAND2_X1 U13638 ( .A1(n10714), .A2(n10713), .ZN(n10744) );
  NAND2_X1 U13639 ( .A1(n10744), .A2(n19884), .ZN(n10726) );
  NAND2_X1 U13640 ( .A1(n12837), .A2(n14806), .ZN(n10715) );
  MUX2_X1 U13641 ( .A(n19884), .B(n10715), .S(n10747), .Z(n10722) );
  INV_X1 U13642 ( .A(n10718), .ZN(n10753) );
  XNOR2_X1 U13643 ( .A(n10739), .B(n10716), .ZN(n10749) );
  OAI211_X1 U13644 ( .C1(n14806), .C2(n10753), .A(n15507), .B(n10749), .ZN(
        n10720) );
  INV_X1 U13645 ( .A(n10739), .ZN(n10717) );
  OAI21_X1 U13646 ( .B1(n10718), .B2(n10717), .A(n10731), .ZN(n10719) );
  OAI211_X1 U13647 ( .C1(n12802), .C2(n10747), .A(n10720), .B(n10719), .ZN(
        n10721) );
  NAND2_X1 U13648 ( .A1(n10722), .A2(n10721), .ZN(n10724) );
  NAND2_X1 U13649 ( .A1(n10724), .A2(n10723), .ZN(n10725) );
  NAND2_X1 U13650 ( .A1(n10726), .A2(n10725), .ZN(n10733) );
  NAND2_X1 U13651 ( .A1(n10728), .A2(n10727), .ZN(n10730) );
  INV_X1 U13652 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n15830) );
  NAND2_X1 U13653 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n15830), .ZN(
        n10729) );
  AOI21_X1 U13654 ( .B1(n10731), .B2(n10746), .A(n10751), .ZN(n10732) );
  NAND2_X1 U13655 ( .A1(n10733), .A2(n10732), .ZN(n10734) );
  MUX2_X1 U13656 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n10734), .S(
        P2_STATE2_REG_0__SCAN_IN), .Z(n10737) );
  INV_X1 U13657 ( .A(n12837), .ZN(n10735) );
  NAND2_X1 U13658 ( .A1(n15479), .A2(n14806), .ZN(n12795) );
  INV_X1 U13659 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n19764) );
  NOR2_X2 U13660 ( .A1(n19759), .A2(P2_STATE_REG_0__SCAN_IN), .ZN(n19833) );
  NAND2_X2 U13661 ( .A1(n19839), .A2(P2_STATE_REG_2__SCAN_IN), .ZN(n19831) );
  INV_X1 U13662 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19776) );
  NAND2_X1 U13663 ( .A1(n19759), .A2(n19776), .ZN(n19770) );
  NAND3_X1 U13664 ( .A1(n19764), .A2(n19831), .A3(n19770), .ZN(n19895) );
  NAND2_X1 U13665 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19898) );
  INV_X1 U13666 ( .A(n19898), .ZN(n16324) );
  NOR2_X1 U13667 ( .A1(n19895), .A2(n16324), .ZN(n13288) );
  NAND2_X1 U13668 ( .A1(n10190), .A2(n13288), .ZN(n10780) );
  AOI21_X1 U13669 ( .B1(n10737), .B2(n15507), .A(n10200), .ZN(n10738) );
  NAND2_X1 U13670 ( .A1(n12795), .A2(n10738), .ZN(n10779) );
  NAND2_X1 U13671 ( .A1(n10753), .A2(n10739), .ZN(n10740) );
  AND2_X1 U13672 ( .A1(n10741), .A2(n10740), .ZN(n10743) );
  INV_X1 U13673 ( .A(n10751), .ZN(n10742) );
  OAI21_X1 U13674 ( .B1(n10744), .B2(n10743), .A(n10742), .ZN(n19883) );
  NAND2_X1 U13675 ( .A1(n19897), .A2(n11518), .ZN(n13250) );
  OR2_X1 U13676 ( .A1(n10745), .A2(n13250), .ZN(n19888) );
  NOR3_X1 U13677 ( .A1(n10748), .A2(n10747), .A3(n10746), .ZN(n10752) );
  AND2_X1 U13678 ( .A1(n10749), .A2(n10752), .ZN(n10750) );
  AOI21_X1 U13679 ( .B1(n10753), .B2(n10752), .A(n13282), .ZN(n10755) );
  NAND2_X1 U13680 ( .A1(n20796), .A2(n10754), .ZN(n12803) );
  INV_X1 U13681 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n18860) );
  OAI21_X1 U13682 ( .B1(n11368), .B2(n12803), .A(n18860), .ZN(n16321) );
  MUX2_X1 U13683 ( .A(n10755), .B(n16321), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n19885) );
  NAND2_X1 U13684 ( .A1(n19885), .A2(n14806), .ZN(n10756) );
  OR2_X1 U13685 ( .A1(n10745), .A2(n10756), .ZN(n10757) );
  NAND2_X1 U13686 ( .A1(n10758), .A2(n10757), .ZN(n11268) );
  NAND2_X1 U13687 ( .A1(n11518), .A2(n10759), .ZN(n10760) );
  AOI21_X1 U13688 ( .B1(n10760), .B2(n15507), .A(n19252), .ZN(n10762) );
  OAI211_X1 U13689 ( .C1(n10762), .C2(n10190), .A(n10761), .B(n10926), .ZN(
        n10763) );
  INV_X1 U13690 ( .A(n10763), .ZN(n10774) );
  NAND3_X1 U13691 ( .A1(n13326), .A2(n12736), .A3(n13288), .ZN(n10773) );
  NAND2_X1 U13692 ( .A1(n10766), .A2(n10767), .ZN(n10768) );
  NAND2_X1 U13693 ( .A1(n10765), .A2(n10768), .ZN(n10772) );
  OR2_X1 U13694 ( .A1(n10769), .A2(n19252), .ZN(n10771) );
  INV_X1 U13695 ( .A(n13250), .ZN(n10770) );
  NAND2_X1 U13696 ( .A1(n10771), .A2(n10770), .ZN(n11183) );
  MUX2_X1 U13697 ( .A(n13326), .B(n10190), .S(n11518), .Z(n10775) );
  NAND3_X1 U13698 ( .A1(n10775), .A2(n12736), .A3(n19898), .ZN(n10776) );
  NAND2_X1 U13699 ( .A1(n12796), .A2(n10776), .ZN(n10777) );
  NOR2_X1 U13700 ( .A1(n11268), .A2(n10777), .ZN(n10778) );
  OAI211_X1 U13701 ( .C1(n12795), .C2(n10780), .A(n10779), .B(n10778), .ZN(
        n10782) );
  NAND2_X1 U13702 ( .A1(n15828), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n19754) );
  INV_X1 U13703 ( .A(n19754), .ZN(n10781) );
  NAND2_X1 U13704 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10781), .ZN(n18857) );
  NOR2_X1 U13705 ( .A1(n10745), .A2(n19884), .ZN(n10783) );
  INV_X1 U13706 ( .A(n10784), .ZN(n13379) );
  NAND2_X1 U13707 ( .A1(n12817), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12816) );
  INV_X1 U13708 ( .A(n12816), .ZN(n10785) );
  XNOR2_X1 U13709 ( .A(n10939), .B(n10950), .ZN(n10786) );
  NAND2_X1 U13710 ( .A1(n10785), .A2(n10786), .ZN(n10787) );
  XOR2_X1 U13711 ( .A(n10786), .B(n10785), .Z(n12828) );
  NAND2_X1 U13712 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n12828), .ZN(
        n12827) );
  NAND2_X1 U13713 ( .A1(n10787), .A2(n12827), .ZN(n10789) );
  XNOR2_X1 U13714 ( .A(n12721), .B(n10789), .ZN(n12728) );
  XNOR2_X1 U13715 ( .A(n10960), .B(n10788), .ZN(n12727) );
  NAND2_X1 U13716 ( .A1(n12728), .A2(n12727), .ZN(n12726) );
  NAND2_X1 U13717 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10789), .ZN(
        n10790) );
  NAND2_X1 U13718 ( .A1(n12726), .A2(n10790), .ZN(n10791) );
  INV_X1 U13719 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13550) );
  XNOR2_X1 U13720 ( .A(n10791), .B(n13550), .ZN(n13378) );
  NAND2_X1 U13721 ( .A1(n13379), .A2(n13378), .ZN(n10793) );
  NAND2_X1 U13722 ( .A1(n10791), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10792) );
  NAND2_X1 U13723 ( .A1(n10793), .A2(n10792), .ZN(n10796) );
  XNOR2_X1 U13724 ( .A(n10794), .B(n10795), .ZN(n10797) );
  XNOR2_X1 U13725 ( .A(n10796), .B(n10797), .ZN(n13540) );
  INV_X1 U13726 ( .A(n10796), .ZN(n10798) );
  NAND2_X1 U13727 ( .A1(n10798), .A2(n10797), .ZN(n10799) );
  AND2_X1 U13728 ( .A1(n10800), .A2(n13717), .ZN(n13706) );
  NAND2_X1 U13729 ( .A1(n10809), .A2(n10807), .ZN(n10805) );
  INV_X1 U13730 ( .A(n10809), .ZN(n10801) );
  NAND2_X1 U13731 ( .A1(n13707), .A2(n10802), .ZN(n10803) );
  OAI211_X2 U13732 ( .C1(n10806), .C2(n10805), .A(n10804), .B(n10803), .ZN(
        n15462) );
  INV_X1 U13733 ( .A(n10806), .ZN(n10808) );
  NAND2_X1 U13734 ( .A1(n10808), .A2(n10807), .ZN(n10810) );
  NAND2_X1 U13735 ( .A1(n10810), .A2(n10809), .ZN(n10811) );
  XNOR2_X1 U13736 ( .A(n10812), .B(n10506), .ZN(n10813) );
  INV_X1 U13737 ( .A(n10813), .ZN(n10814) );
  NAND2_X1 U13738 ( .A1(n10814), .A2(n15454), .ZN(n15173) );
  XNOR2_X1 U13739 ( .A(n10815), .B(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n16275) );
  INV_X1 U13740 ( .A(n10812), .ZN(n10816) );
  NAND3_X1 U13741 ( .A1(n10816), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A3(
        n10506), .ZN(n10817) );
  AND2_X1 U13742 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15384) );
  AND2_X1 U13743 ( .A1(n15384), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15331) );
  NAND2_X1 U13744 ( .A1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15337) );
  NOR2_X1 U13745 ( .A1(n15337), .A2(n10819), .ZN(n10820) );
  AND2_X1 U13746 ( .A1(n15331), .A2(n10820), .ZN(n15318) );
  NAND3_X1 U13747 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15330) );
  NOR2_X1 U13748 ( .A1(n15330), .A2(n15317), .ZN(n10821) );
  NAND2_X1 U13749 ( .A1(n15318), .A2(n10821), .ZN(n11201) );
  NOR2_X1 U13750 ( .A1(n11201), .A2(n15293), .ZN(n10822) );
  INV_X1 U13751 ( .A(n19888), .ZN(n10824) );
  NAND2_X1 U13752 ( .A1(n15009), .A2(n16294), .ZN(n11221) );
  NAND2_X1 U13753 ( .A1(n10827), .A2(n10828), .ZN(n10826) );
  NAND2_X1 U13754 ( .A1(n10826), .A2(n10825), .ZN(n10831) );
  NAND2_X1 U13755 ( .A1(n10246), .A2(n10247), .ZN(n10829) );
  NAND3_X1 U13756 ( .A1(n10831), .A2(n10830), .A3(n10829), .ZN(n10835) );
  OR2_X1 U13757 ( .A1(n10833), .A2(n10832), .ZN(n10834) );
  NAND2_X1 U13758 ( .A1(n10856), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10839) );
  AOI22_X1 U13759 ( .A1(n10863), .A2(P2_REIP_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10838) );
  OAI211_X1 U13760 ( .C1(n11250), .C2(n19084), .A(n10839), .B(n10838), .ZN(
        n12957) );
  NAND2_X1 U13761 ( .A1(n10856), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10842) );
  NAND2_X1 U13762 ( .A1(n10909), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n10841) );
  AOI22_X1 U13763 ( .A1(n10863), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10840) );
  NAND2_X1 U13764 ( .A1(n10916), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10846) );
  NAND2_X1 U13765 ( .A1(n10909), .A2(P2_EBX_REG_6__SCAN_IN), .ZN(n10845) );
  AOI22_X1 U13766 ( .A1(n10863), .A2(P2_REIP_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10844) );
  INV_X1 U13767 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n13076) );
  NAND2_X1 U13768 ( .A1(n10916), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10848) );
  AOI22_X1 U13769 ( .A1(n10863), .A2(P2_REIP_REG_7__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10847) );
  OAI211_X1 U13770 ( .C1(n11250), .C2(n13076), .A(n10848), .B(n10847), .ZN(
        n13072) );
  NAND2_X1 U13771 ( .A1(n13073), .A2(n13072), .ZN(n13063) );
  NAND2_X1 U13772 ( .A1(n10916), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10851) );
  NAND2_X1 U13773 ( .A1(n10909), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10850) );
  AOI22_X1 U13774 ( .A1(n10863), .A2(P2_REIP_REG_8__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10849) );
  NAND2_X1 U13775 ( .A1(n10916), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10854) );
  NAND2_X1 U13776 ( .A1(n10909), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10853) );
  AOI22_X1 U13777 ( .A1(n10863), .A2(P2_REIP_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10852) );
  NAND2_X1 U13778 ( .A1(n13049), .A2(n10855), .ZN(n13143) );
  NAND2_X1 U13779 ( .A1(n10916), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10859) );
  NAND2_X1 U13780 ( .A1(n10909), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n10858) );
  AOI22_X1 U13781 ( .A1(n10863), .A2(P2_REIP_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n10857) );
  INV_X1 U13782 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n10862) );
  NAND2_X1 U13783 ( .A1(n10856), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n10861) );
  AOI22_X1 U13784 ( .A1(n10863), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_11__SCAN_IN), 
        .ZN(n10860) );
  OAI211_X1 U13785 ( .C1(n11250), .C2(n10862), .A(n10861), .B(n10860), .ZN(
        n13150) );
  NAND2_X1 U13786 ( .A1(n10856), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10866) );
  NAND2_X1 U13787 ( .A1(n10909), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10865) );
  AOI22_X1 U13788 ( .A1(n10863), .A2(P2_REIP_REG_12__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), 
        .ZN(n10864) );
  NAND2_X1 U13789 ( .A1(n10856), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10870) );
  NAND2_X1 U13790 ( .A1(n10909), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10869) );
  AOI22_X1 U13791 ( .A1(n10863), .A2(P2_REIP_REG_13__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n10868) );
  INV_X1 U13792 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n10873) );
  NAND2_X1 U13793 ( .A1(n10856), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10872) );
  AOI22_X1 U13794 ( .A1(n10863), .A2(P2_REIP_REG_14__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n10871) );
  OAI211_X1 U13795 ( .C1(n11250), .C2(n10873), .A(n10872), .B(n10871), .ZN(
        n13517) );
  AND2_X2 U13796 ( .A1(n13518), .A2(n13517), .ZN(n13679) );
  INV_X1 U13797 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n10876) );
  NAND2_X1 U13798 ( .A1(n10856), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10875) );
  AOI22_X1 U13799 ( .A1(n10863), .A2(P2_REIP_REG_15__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), 
        .ZN(n10874) );
  OAI211_X1 U13800 ( .C1(n11250), .C2(n10876), .A(n10875), .B(n10874), .ZN(
        n13678) );
  NAND2_X1 U13801 ( .A1(n10856), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10879) );
  NAND2_X1 U13802 ( .A1(n10909), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10878) );
  AOI22_X1 U13803 ( .A1(n10863), .A2(P2_REIP_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n10877) );
  NAND2_X1 U13804 ( .A1(n10856), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n10882) );
  NAND2_X1 U13805 ( .A1(n10909), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10881) );
  AOI22_X1 U13806 ( .A1(n10863), .A2(P2_REIP_REG_17__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), 
        .ZN(n10880) );
  INV_X1 U13807 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n10885) );
  NAND2_X1 U13808 ( .A1(n10856), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n10884) );
  AOI22_X1 U13809 ( .A1(n10863), .A2(P2_REIP_REG_18__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), 
        .ZN(n10883) );
  OAI211_X1 U13810 ( .C1(n11250), .C2(n10885), .A(n10884), .B(n10883), .ZN(
        n14854) );
  NAND2_X1 U13811 ( .A1(n10856), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10888) );
  NAND2_X1 U13812 ( .A1(n10909), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n10887) );
  AOI22_X1 U13813 ( .A1(n10863), .A2(P2_REIP_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n10886) );
  NAND2_X1 U13814 ( .A1(n10916), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10891) );
  NAND2_X1 U13815 ( .A1(n10909), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10890) );
  AOI22_X1 U13816 ( .A1(n10863), .A2(P2_REIP_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n10889) );
  OR2_X2 U13817 ( .A1(n14848), .A2(n14838), .ZN(n14839) );
  NAND2_X1 U13818 ( .A1(n10916), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n10894) );
  NAND2_X1 U13819 ( .A1(n10909), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10893) );
  AOI22_X1 U13820 ( .A1(n10863), .A2(P2_REIP_REG_21__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_21__SCAN_IN), 
        .ZN(n10892) );
  INV_X1 U13821 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n10897) );
  NAND2_X1 U13822 ( .A1(n10916), .A2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n10896) );
  AOI22_X1 U13823 ( .A1(n10863), .A2(P2_REIP_REG_22__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), 
        .ZN(n10895) );
  OAI211_X1 U13824 ( .C1(n11250), .C2(n10897), .A(n10896), .B(n10895), .ZN(
        n14823) );
  NAND2_X1 U13825 ( .A1(n14833), .A2(n14823), .ZN(n14814) );
  NAND2_X1 U13826 ( .A1(n10916), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10900) );
  NAND2_X1 U13827 ( .A1(n10909), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10899) );
  AOI22_X1 U13828 ( .A1(n10863), .A2(P2_REIP_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n10898) );
  NAND2_X1 U13829 ( .A1(n10916), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n10903) );
  NAND2_X1 U13830 ( .A1(n10909), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10902) );
  AOI22_X1 U13831 ( .A1(n10863), .A2(P2_REIP_REG_24__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), 
        .ZN(n10901) );
  NAND2_X1 U13832 ( .A1(n10916), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n10905) );
  AOI22_X1 U13833 ( .A1(n10863), .A2(P2_REIP_REG_25__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_25__SCAN_IN), 
        .ZN(n10904) );
  OAI211_X1 U13834 ( .C1(n11250), .C2(n10683), .A(n10905), .B(n10904), .ZN(
        n14799) );
  INV_X1 U13835 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n10908) );
  NAND2_X1 U13836 ( .A1(n10916), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n10907) );
  AOI22_X1 U13837 ( .A1(n10863), .A2(P2_REIP_REG_26__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n10906) );
  OAI211_X1 U13838 ( .C1(n11250), .C2(n10908), .A(n10907), .B(n10906), .ZN(
        n14791) );
  NAND2_X1 U13839 ( .A1(n10916), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10912) );
  NAND2_X1 U13840 ( .A1(n10909), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10911) );
  AOI22_X1 U13841 ( .A1(n10863), .A2(P2_REIP_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n10910) );
  AND3_X1 U13842 ( .A1(n10912), .A2(n10911), .A3(n10910), .ZN(n14784) );
  NAND2_X1 U13843 ( .A1(n10856), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10915) );
  NAND2_X1 U13844 ( .A1(n10909), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n10914) );
  AOI22_X1 U13845 ( .A1(n10863), .A2(P2_REIP_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n10913) );
  AND3_X1 U13846 ( .A1(n10915), .A2(n10914), .A3(n10913), .ZN(n14776) );
  INV_X1 U13847 ( .A(P2_EBX_REG_29__SCAN_IN), .ZN(n10919) );
  NAND2_X1 U13848 ( .A1(n10916), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10918) );
  AOI22_X1 U13849 ( .A1(n10863), .A2(P2_REIP_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n10917) );
  OAI211_X1 U13850 ( .C1(n11250), .C2(n10919), .A(n10918), .B(n10917), .ZN(
        n11226) );
  INV_X1 U13851 ( .A(P2_EBX_REG_30__SCAN_IN), .ZN(n10921) );
  AOI22_X1 U13852 ( .A1(n10863), .A2(P2_REIP_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n10920) );
  OAI21_X1 U13853 ( .B1(n11250), .B2(n10921), .A(n10920), .ZN(n10922) );
  AOI21_X1 U13854 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n10856), .A(
        n10922), .ZN(n11247) );
  INV_X1 U13855 ( .A(n10923), .ZN(n10924) );
  OR2_X1 U13856 ( .A1(n10764), .A2(n15507), .ZN(n12738) );
  NAND2_X1 U13857 ( .A1(n10924), .A2(n12738), .ZN(n13304) );
  NAND2_X1 U13858 ( .A1(n13304), .A2(n11518), .ZN(n10927) );
  INV_X1 U13859 ( .A(n10925), .ZN(n13299) );
  OR2_X1 U13860 ( .A1(n13299), .A2(n10926), .ZN(n13259) );
  NAND2_X1 U13861 ( .A1(n10927), .A2(n13259), .ZN(n10928) );
  NAND2_X1 U13862 ( .A1(n11194), .A2(n10928), .ZN(n15445) );
  NOR2_X1 U13863 ( .A1(n16142), .A2(n15445), .ZN(n11219) );
  NOR2_X1 U13864 ( .A1(n10176), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n10929) );
  AOI22_X1 U13865 ( .A1(n11157), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n11167), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10933) );
  NOR2_X1 U13866 ( .A1(n10930), .A2(n10671), .ZN(n10931) );
  NAND2_X1 U13867 ( .A1(n11158), .A2(P2_REIP_REG_30__SCAN_IN), .ZN(n10932) );
  AND2_X1 U13868 ( .A1(n10933), .A2(n10932), .ZN(n11171) );
  INV_X1 U13869 ( .A(n10204), .ZN(n10936) );
  NAND2_X1 U13870 ( .A1(n10936), .A2(n11167), .ZN(n10959) );
  INV_X1 U13871 ( .A(n10951), .ZN(n10944) );
  NOR2_X1 U13872 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19697), .ZN(
        n19874) );
  INV_X1 U13873 ( .A(n19874), .ZN(n10937) );
  NAND2_X1 U13874 ( .A1(n10944), .A2(n10937), .ZN(n10938) );
  AND2_X1 U13875 ( .A1(n10959), .A2(n10938), .ZN(n10943) );
  INV_X1 U13876 ( .A(n10939), .ZN(n10941) );
  NAND2_X1 U13877 ( .A1(n10943), .A2(n10942), .ZN(n12988) );
  INV_X1 U13878 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n16304) );
  NAND2_X1 U13879 ( .A1(n10947), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10946) );
  OAI21_X1 U13880 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(P2_EAX_REG_0__SCAN_IN), 
        .A(n10944), .ZN(n10945) );
  OAI211_X1 U13881 ( .C1(n11518), .C2(n16304), .A(n10946), .B(n10945), .ZN(
        n12987) );
  AOI22_X1 U13882 ( .A1(n10929), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n11167), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n10949) );
  NAND2_X1 U13883 ( .A1(n10947), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10948) );
  NAND2_X1 U13884 ( .A1(n10949), .A2(n10948), .ZN(n10955) );
  XNOR2_X1 U13885 ( .A(n12990), .B(n10955), .ZN(n12863) );
  INV_X1 U13886 ( .A(n10950), .ZN(n10954) );
  NAND2_X1 U13887 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10953) );
  NAND2_X1 U13888 ( .A1(n10204), .A2(n10951), .ZN(n10952) );
  OAI211_X1 U13889 ( .C1(n11137), .C2(n10954), .A(n10953), .B(n10952), .ZN(
        n12862) );
  NOR2_X1 U13890 ( .A1(n12863), .A2(n12862), .ZN(n10957) );
  NOR2_X1 U13891 ( .A1(n12990), .A2(n10955), .ZN(n10956) );
  NAND2_X1 U13892 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n10958) );
  OAI211_X1 U13893 ( .C1(n10960), .C2(n11137), .A(n10959), .B(n10958), .ZN(
        n10963) );
  XNOR2_X1 U13894 ( .A(n10964), .B(n10963), .ZN(n12715) );
  AOI22_X1 U13895 ( .A1(n11157), .A2(P2_EAX_REG_2__SCAN_IN), .B1(n11167), .B2(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n10962) );
  INV_X2 U13896 ( .A(n10980), .ZN(n11158) );
  NAND2_X1 U13897 ( .A1(n11158), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n10961) );
  NAND2_X1 U13898 ( .A1(n10962), .A2(n10961), .ZN(n12714) );
  NOR2_X1 U13899 ( .A1(n12715), .A2(n12714), .ZN(n12716) );
  NOR2_X1 U13900 ( .A1(n10964), .A2(n10963), .ZN(n10965) );
  NOR2_X2 U13901 ( .A1(n12716), .A2(n10965), .ZN(n13385) );
  NAND2_X1 U13902 ( .A1(n11158), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n10970) );
  NAND2_X1 U13903 ( .A1(n10940), .A2(n10966), .ZN(n10969) );
  AOI22_X1 U13904 ( .A1(n11167), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n10968) );
  NAND2_X1 U13905 ( .A1(n11157), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n10967) );
  NAND4_X1 U13906 ( .A1(n10970), .A2(n10969), .A3(n10968), .A4(n10967), .ZN(
        n13384) );
  AOI22_X1 U13907 ( .A1(n11157), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n11167), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n10974) );
  NAND2_X1 U13908 ( .A1(n11158), .A2(P2_REIP_REG_4__SCAN_IN), .ZN(n10973) );
  NAND2_X1 U13909 ( .A1(n10940), .A2(n10971), .ZN(n10972) );
  AOI22_X1 U13910 ( .A1(n11158), .A2(P2_REIP_REG_5__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n11167), .ZN(n10977) );
  AOI22_X1 U13911 ( .A1(n10940), .A2(n10975), .B1(n11157), .B2(
        P2_EAX_REG_5__SCAN_IN), .ZN(n10976) );
  NAND2_X1 U13912 ( .A1(n10977), .A2(n10976), .ZN(n13714) );
  AOI21_X1 U13913 ( .B1(n10940), .B2(n10979), .A(n10978), .ZN(n12925) );
  AOI222_X1 U13914 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n11158), .B1(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n11167), .C1(
        P2_EAX_REG_6__SCAN_IN), .C2(n11157), .ZN(n12924) );
  INV_X1 U13915 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19189) );
  INV_X1 U13916 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n19787) );
  OAI222_X1 U13917 ( .A1(n11035), .A2(n15454), .B1(n11093), .B2(n19189), .C1(
        n10980), .C2(n19787), .ZN(n12920) );
  INV_X1 U13918 ( .A(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15516) );
  NAND2_X1 U13919 ( .A1(n11464), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n10982) );
  NAND2_X1 U13920 ( .A1(n10350), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n10981) );
  OAI211_X1 U13921 ( .C1(n15516), .C2(n10480), .A(n10982), .B(n10981), .ZN(
        n10985) );
  INV_X1 U13922 ( .A(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10983) );
  INV_X1 U13923 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11502) );
  OAI22_X1 U13924 ( .A1(n11470), .A2(n10983), .B1(n11469), .B2(n11502), .ZN(
        n10984) );
  NOR2_X1 U13925 ( .A1(n10985), .A2(n10984), .ZN(n10996) );
  AOI22_X1 U13926 ( .A1(n11368), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11473), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10995) );
  INV_X1 U13927 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11336) );
  AOI22_X1 U13928 ( .A1(n10448), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10408), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10987) );
  NAND2_X1 U13929 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n10986) );
  OAI211_X1 U13930 ( .C1(n11477), .C2(n11336), .A(n10987), .B(n10986), .ZN(
        n10992) );
  NAND2_X1 U13931 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n10989) );
  NAND2_X1 U13932 ( .A1(n11478), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n10988) );
  OAI211_X1 U13933 ( .C1(n10473), .C2(n10990), .A(n10989), .B(n10988), .ZN(
        n10991) );
  NOR2_X1 U13934 ( .A1(n10992), .A2(n10991), .ZN(n10994) );
  AOI22_X1 U13935 ( .A1(n10407), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n10403), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10993) );
  NAND4_X1 U13936 ( .A1(n10996), .A2(n10995), .A3(n10994), .A4(n10993), .ZN(
        n13062) );
  INV_X1 U13937 ( .A(n13062), .ZN(n10998) );
  AOI22_X1 U13938 ( .A1(n11157), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n11167), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n10997) );
  OAI21_X1 U13939 ( .B1(n10998), .B2(n11137), .A(n10997), .ZN(n10999) );
  AOI21_X1 U13940 ( .B1(P2_REIP_REG_8__SCAN_IN), .B2(n11158), .A(n10999), .ZN(
        n16291) );
  AOI22_X1 U13941 ( .A1(n11158), .A2(P2_REIP_REG_9__SCAN_IN), .B1(n10929), 
        .B2(P2_EAX_REG_9__SCAN_IN), .ZN(n11017) );
  INV_X1 U13942 ( .A(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11002) );
  NAND2_X1 U13943 ( .A1(n11464), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11001) );
  NAND2_X1 U13944 ( .A1(n10350), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11000) );
  OAI211_X1 U13945 ( .C1(n10480), .C2(n11002), .A(n11001), .B(n11000), .ZN(
        n11005) );
  INV_X1 U13946 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11529) );
  OAI22_X1 U13947 ( .A1(n11003), .A2(n11470), .B1(n11469), .B2(n11529), .ZN(
        n11004) );
  NOR2_X1 U13948 ( .A1(n11005), .A2(n11004), .ZN(n11015) );
  AOI22_X1 U13949 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n11473), .B1(
        n11368), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11014) );
  AOI22_X1 U13950 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n11478), .B1(
        n10351), .B2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11011) );
  NAND2_X1 U13951 ( .A1(n11044), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11010) );
  INV_X1 U13952 ( .A(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11006) );
  INV_X1 U13953 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11522) );
  OAI22_X1 U13954 ( .A1(n11006), .A2(n10377), .B1(n11522), .B2(n10364), .ZN(
        n11007) );
  AOI21_X1 U13955 ( .B1(n10380), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A(
        n11007), .ZN(n11009) );
  NAND2_X1 U13956 ( .A1(n11047), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11008) );
  AND4_X1 U13957 ( .A1(n11011), .A2(n11010), .A3(n11009), .A4(n11008), .ZN(
        n11013) );
  AOI22_X1 U13958 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n11399), .B1(
        n10403), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11012) );
  NAND4_X1 U13959 ( .A1(n11015), .A2(n11014), .A3(n11013), .A4(n11012), .ZN(
        n13056) );
  AOI22_X1 U13960 ( .A1(n10940), .A2(n13056), .B1(n11167), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n11016) );
  NAND2_X1 U13961 ( .A1(n11017), .A2(n11016), .ZN(n13045) );
  INV_X1 U13962 ( .A(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11020) );
  NAND2_X1 U13963 ( .A1(n11464), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(
        n11019) );
  NAND2_X1 U13964 ( .A1(n10350), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11018) );
  OAI211_X1 U13965 ( .C1(n10480), .C2(n11020), .A(n11019), .B(n11018), .ZN(
        n11023) );
  INV_X1 U13966 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11021) );
  INV_X1 U13967 ( .A(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11549) );
  OAI22_X1 U13968 ( .A1(n11021), .A2(n11470), .B1(n11469), .B2(n11549), .ZN(
        n11022) );
  NOR2_X1 U13969 ( .A1(n11023), .A2(n11022), .ZN(n11034) );
  AOI22_X1 U13970 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n11473), .B1(
        n11368), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11033) );
  INV_X1 U13971 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11376) );
  AOI22_X1 U13972 ( .A1(n10448), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n10408), .ZN(n11025) );
  NAND2_X1 U13973 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n11024) );
  OAI211_X1 U13974 ( .C1(n11477), .C2(n11376), .A(n11025), .B(n11024), .ZN(
        n11030) );
  NAND2_X1 U13975 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(
        n11027) );
  NAND2_X1 U13976 ( .A1(n11478), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11026) );
  OAI211_X1 U13977 ( .C1(n10473), .C2(n11028), .A(n11027), .B(n11026), .ZN(
        n11029) );
  NOR2_X1 U13978 ( .A1(n11030), .A2(n11029), .ZN(n11032) );
  AOI22_X1 U13979 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n10407), .B1(
        n10403), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11031) );
  NAND4_X1 U13980 ( .A1(n11034), .A2(n11033), .A3(n11032), .A4(n11031), .ZN(
        n13147) );
  INV_X1 U13981 ( .A(n13147), .ZN(n11321) );
  AOI22_X1 U13982 ( .A1(n10929), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n11167), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11036) );
  OAI21_X1 U13983 ( .B1(n11321), .B2(n11137), .A(n11036), .ZN(n11037) );
  AOI21_X1 U13984 ( .B1(P2_REIP_REG_10__SCAN_IN), .B2(n11158), .A(n11037), 
        .ZN(n13046) );
  NAND2_X1 U13985 ( .A1(n11464), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(
        n11039) );
  NAND2_X1 U13986 ( .A1(n10350), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n11038) );
  OAI211_X1 U13987 ( .C1(n10480), .C2(n11040), .A(n11039), .B(n11038), .ZN(
        n11043) );
  OAI22_X1 U13988 ( .A1(n11041), .A2(n11470), .B1(n11469), .B2(n11574), .ZN(
        n11042) );
  NOR2_X1 U13989 ( .A1(n11043), .A2(n11042), .ZN(n11055) );
  AOI22_X1 U13990 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n11473), .B1(
        n11368), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11054) );
  AOI22_X1 U13991 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n11478), .B1(
        n10351), .B2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11051) );
  NAND2_X1 U13992 ( .A1(n11044), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(
        n11050) );
  INV_X1 U13993 ( .A(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11045) );
  OAI22_X1 U13994 ( .A1(n11045), .A2(n10377), .B1(n11567), .B2(n10364), .ZN(
        n11046) );
  AOI21_X1 U13995 ( .B1(n10380), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n11046), .ZN(n11049) );
  NAND2_X1 U13996 ( .A1(n11047), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n11048) );
  AND4_X1 U13997 ( .A1(n11051), .A2(n11050), .A3(n11049), .A4(n11048), .ZN(
        n11053) );
  AOI22_X1 U13998 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n10407), .B1(
        n10403), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11052) );
  NAND4_X1 U13999 ( .A1(n11055), .A2(n11054), .A3(n11053), .A4(n11052), .ZN(
        n13153) );
  AOI22_X1 U14000 ( .A1(n11158), .A2(P2_REIP_REG_11__SCAN_IN), .B1(n10940), 
        .B2(n13153), .ZN(n11057) );
  AOI22_X1 U14001 ( .A1(n10929), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n11167), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n11056) );
  NAND2_X1 U14002 ( .A1(n11057), .A2(n11056), .ZN(n13157) );
  NAND2_X1 U14003 ( .A1(n13158), .A2(n13157), .ZN(n13216) );
  INV_X1 U14004 ( .A(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n11060) );
  NAND2_X1 U14005 ( .A1(n11464), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11059) );
  NAND2_X1 U14006 ( .A1(n10350), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11058) );
  OAI211_X1 U14007 ( .C1(n10480), .C2(n11060), .A(n11059), .B(n11058), .ZN(
        n11063) );
  INV_X1 U14008 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11061) );
  INV_X1 U14009 ( .A(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n11597) );
  OAI22_X1 U14010 ( .A1(n11061), .A2(n11470), .B1(n11469), .B2(n11597), .ZN(
        n11062) );
  NOR2_X1 U14011 ( .A1(n11063), .A2(n11062), .ZN(n11074) );
  AOI22_X1 U14012 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n11473), .B1(
        n11368), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11073) );
  INV_X1 U14013 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11416) );
  AOI22_X1 U14014 ( .A1(n10448), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n10408), .ZN(n11065) );
  NAND2_X1 U14015 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11064) );
  OAI211_X1 U14016 ( .C1(n11477), .C2(n11416), .A(n11065), .B(n11064), .ZN(
        n11070) );
  NAND2_X1 U14017 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11067) );
  NAND2_X1 U14018 ( .A1(n11478), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11066) );
  OAI211_X1 U14019 ( .C1(n10473), .C2(n11068), .A(n11067), .B(n11066), .ZN(
        n11069) );
  NOR2_X1 U14020 ( .A1(n11070), .A2(n11069), .ZN(n11072) );
  AOI22_X1 U14021 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n11399), .B1(
        n10403), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11071) );
  NAND4_X1 U14022 ( .A1(n11074), .A2(n11073), .A3(n11072), .A4(n11071), .ZN(
        n13224) );
  AOI22_X1 U14023 ( .A1(n10929), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n11167), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11075) );
  OAI21_X1 U14024 ( .B1(n11322), .B2(n11137), .A(n11075), .ZN(n11076) );
  AOI21_X1 U14025 ( .B1(P2_REIP_REG_12__SCAN_IN), .B2(n11158), .A(n11076), 
        .ZN(n13217) );
  NAND2_X1 U14026 ( .A1(n11464), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11078) );
  NAND2_X1 U14027 ( .A1(n10350), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11077) );
  OAI211_X1 U14028 ( .C1(n11079), .C2(n10480), .A(n11078), .B(n11077), .ZN(
        n11081) );
  OAI22_X1 U14029 ( .A1(n11470), .A2(n11626), .B1(n11469), .B2(n11624), .ZN(
        n11080) );
  NOR2_X1 U14030 ( .A1(n11081), .A2(n11080), .ZN(n11092) );
  AOI22_X1 U14031 ( .A1(n11368), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11473), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11091) );
  AOI22_X1 U14032 ( .A1(n10448), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10408), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11083) );
  NAND2_X1 U14033 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11082) );
  OAI211_X1 U14034 ( .C1(n11477), .C2(n11434), .A(n11083), .B(n11082), .ZN(
        n11088) );
  NAND2_X1 U14035 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11085) );
  NAND2_X1 U14036 ( .A1(n11478), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11084) );
  OAI211_X1 U14037 ( .C1(n10473), .C2(n11086), .A(n11085), .B(n11084), .ZN(
        n11087) );
  NOR2_X1 U14038 ( .A1(n11088), .A2(n11087), .ZN(n11090) );
  AOI22_X1 U14039 ( .A1(n10407), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10403), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11089) );
  NAND4_X1 U14040 ( .A1(n11092), .A2(n11091), .A3(n11090), .A4(n11089), .ZN(
        n13465) );
  INV_X1 U14041 ( .A(n13465), .ZN(n11096) );
  AOI22_X1 U14042 ( .A1(n11157), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n11167), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n11095) );
  NAND2_X1 U14043 ( .A1(n11158), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n11094) );
  OAI211_X1 U14044 ( .C1(n11096), .C2(n11137), .A(n11095), .B(n11094), .ZN(
        n13247) );
  NAND2_X1 U14045 ( .A1(n11464), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11098) );
  NAND2_X1 U14046 ( .A1(n10350), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11097) );
  OAI211_X1 U14047 ( .C1(n11099), .C2(n10480), .A(n11098), .B(n11097), .ZN(
        n11102) );
  OAI22_X1 U14048 ( .A1(n11470), .A2(n11100), .B1(n11469), .B2(n11447), .ZN(
        n11101) );
  NOR2_X1 U14049 ( .A1(n11102), .A2(n11101), .ZN(n11113) );
  AOI22_X1 U14050 ( .A1(n11368), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n11473), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11112) );
  AOI22_X1 U14051 ( .A1(n10448), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10408), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11104) );
  NAND2_X1 U14052 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11103) );
  OAI211_X1 U14053 ( .C1(n11477), .C2(n11456), .A(n11104), .B(n11103), .ZN(
        n11109) );
  NAND2_X1 U14054 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11106) );
  NAND2_X1 U14055 ( .A1(n11478), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11105) );
  OAI211_X1 U14056 ( .C1(n10473), .C2(n11107), .A(n11106), .B(n11105), .ZN(
        n11108) );
  NOR2_X1 U14057 ( .A1(n11109), .A2(n11108), .ZN(n11111) );
  AOI22_X1 U14058 ( .A1(n10407), .A2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n10403), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11110) );
  NAND4_X1 U14059 ( .A1(n11113), .A2(n11112), .A3(n11111), .A4(n11110), .ZN(
        n13524) );
  INV_X1 U14060 ( .A(n13524), .ZN(n11323) );
  AOI22_X1 U14061 ( .A1(n11157), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n11167), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11114) );
  OAI21_X1 U14062 ( .B1(n11323), .B2(n11137), .A(n11114), .ZN(n11115) );
  AOI21_X1 U14063 ( .B1(P2_REIP_REG_14__SCAN_IN), .B2(n11158), .A(n11115), 
        .ZN(n15366) );
  INV_X1 U14064 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11481) );
  AOI22_X1 U14065 ( .A1(n10448), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n10408), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11117) );
  NAND2_X1 U14066 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11116) );
  OAI211_X1 U14067 ( .C1(n11477), .C2(n11481), .A(n11117), .B(n11116), .ZN(
        n11122) );
  INV_X1 U14068 ( .A(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11120) );
  NAND2_X1 U14069 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n11119) );
  NAND2_X1 U14070 ( .A1(n11478), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11118) );
  OAI211_X1 U14071 ( .C1(n10473), .C2(n11120), .A(n11119), .B(n11118), .ZN(
        n11121) );
  NOR2_X1 U14072 ( .A1(n11122), .A2(n11121), .ZN(n11126) );
  AOI22_X1 U14073 ( .A1(n11473), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11464), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11125) );
  NAND2_X1 U14074 ( .A1(n10407), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n11124) );
  NAND2_X1 U14075 ( .A1(n11368), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n11123) );
  NAND4_X1 U14076 ( .A1(n11126), .A2(n11125), .A3(n11124), .A4(n11123), .ZN(
        n11134) );
  AOI22_X1 U14077 ( .A1(n10403), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11127), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11132) );
  AOI22_X1 U14078 ( .A1(n11128), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10350), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11131) );
  NAND2_X1 U14079 ( .A1(n11129), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n11130) );
  NAND3_X1 U14080 ( .A1(n11132), .A2(n11131), .A3(n11130), .ZN(n11133) );
  NOR2_X1 U14081 ( .A1(n11134), .A2(n11133), .ZN(n13680) );
  AOI22_X1 U14082 ( .A1(n11157), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n11167), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11136) );
  NAND2_X1 U14083 ( .A1(n11158), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n11135) );
  OAI211_X1 U14084 ( .C1(n13680), .C2(n11137), .A(n11136), .B(n11135), .ZN(
        n13583) );
  AOI22_X1 U14085 ( .A1(n11157), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n11167), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n11139) );
  NAND2_X1 U14086 ( .A1(n11158), .A2(P2_REIP_REG_16__SCAN_IN), .ZN(n11138) );
  NAND2_X1 U14087 ( .A1(n11139), .A2(n11138), .ZN(n14988) );
  AOI22_X1 U14088 ( .A1(n11157), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n11167), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11141) );
  NAND2_X1 U14089 ( .A1(n11158), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n11140) );
  AND2_X1 U14090 ( .A1(n11141), .A2(n11140), .ZN(n14979) );
  AOI22_X1 U14091 ( .A1(n11157), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n11167), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11143) );
  NAND2_X1 U14092 ( .A1(n11158), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n11142) );
  AND2_X1 U14093 ( .A1(n11143), .A2(n11142), .ZN(n14970) );
  AOI22_X1 U14094 ( .A1(n11157), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n11167), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n11145) );
  NAND2_X1 U14095 ( .A1(n11158), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n11144) );
  NAND2_X1 U14096 ( .A1(n11145), .A2(n11144), .ZN(n14961) );
  AOI22_X1 U14097 ( .A1(n11157), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n11167), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11147) );
  NAND2_X1 U14098 ( .A1(n11158), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n11146) );
  NAND2_X1 U14099 ( .A1(n11147), .A2(n11146), .ZN(n14950) );
  AOI22_X1 U14100 ( .A1(n11157), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n11167), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11149) );
  NAND2_X1 U14101 ( .A1(n11158), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n11148) );
  NAND2_X1 U14102 ( .A1(n11149), .A2(n11148), .ZN(n14942) );
  AOI22_X1 U14103 ( .A1(n11157), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n11167), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11151) );
  NAND2_X1 U14104 ( .A1(n11158), .A2(P2_REIP_REG_22__SCAN_IN), .ZN(n11150) );
  NAND2_X1 U14105 ( .A1(n11151), .A2(n11150), .ZN(n14934) );
  AOI22_X1 U14106 ( .A1(n11157), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n11167), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n11153) );
  NAND2_X1 U14107 ( .A1(n11158), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n11152) );
  NAND2_X1 U14108 ( .A1(n11153), .A2(n11152), .ZN(n14919) );
  AOI22_X1 U14109 ( .A1(n11157), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n11167), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n11156) );
  NAND2_X1 U14110 ( .A1(n11158), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n11155) );
  AND2_X1 U14111 ( .A1(n11156), .A2(n11155), .ZN(n14911) );
  AOI22_X1 U14112 ( .A1(n11157), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n11167), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11160) );
  NAND2_X1 U14113 ( .A1(n11158), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n11159) );
  AND2_X1 U14114 ( .A1(n11160), .A2(n11159), .ZN(n14901) );
  AOI22_X1 U14115 ( .A1(n11157), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n11167), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11162) );
  NAND2_X1 U14116 ( .A1(n11158), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n11161) );
  NAND2_X1 U14117 ( .A1(n11162), .A2(n11161), .ZN(n14890) );
  AOI22_X1 U14118 ( .A1(n11157), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n11167), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11164) );
  NAND2_X1 U14119 ( .A1(n11158), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n11163) );
  NAND2_X1 U14120 ( .A1(n11164), .A2(n11163), .ZN(n14883) );
  AOI22_X1 U14121 ( .A1(n11157), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n11167), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11166) );
  NAND2_X1 U14122 ( .A1(n11158), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n11165) );
  NAND2_X1 U14123 ( .A1(n11166), .A2(n11165), .ZN(n14874) );
  AOI22_X1 U14124 ( .A1(n11157), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n11167), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n11169) );
  NAND2_X1 U14125 ( .A1(n11158), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11168) );
  AOI21_X1 U14126 ( .B1(n11171), .B2(n11170), .A(n11255), .ZN(n16136) );
  AND2_X1 U14127 ( .A1(n11172), .A2(n10925), .ZN(n13283) );
  INV_X1 U14128 ( .A(n13283), .ZN(n13254) );
  NAND2_X1 U14129 ( .A1(n12738), .A2(n10765), .ZN(n13281) );
  NAND2_X1 U14130 ( .A1(n13281), .A2(n14806), .ZN(n11173) );
  NAND2_X1 U14131 ( .A1(n13254), .A2(n11173), .ZN(n11174) );
  AND3_X1 U14132 ( .A1(n10671), .A2(n10767), .A3(n11518), .ZN(n11175) );
  AND2_X1 U14133 ( .A1(n10925), .A2(n11175), .ZN(n13284) );
  NAND2_X1 U14134 ( .A1(n11194), .A2(n13284), .ZN(n15333) );
  MUX2_X1 U14135 ( .A(n12802), .B(n11177), .S(n11176), .Z(n11179) );
  NAND2_X1 U14136 ( .A1(n11179), .A2(n19899), .ZN(n11181) );
  NAND2_X1 U14137 ( .A1(n11181), .A2(n11180), .ZN(n11191) );
  NAND2_X1 U14138 ( .A1(n11182), .A2(n14806), .ZN(n13298) );
  NAND2_X1 U14139 ( .A1(n13298), .A2(n11183), .ZN(n11188) );
  OAI22_X1 U14140 ( .A1(n19899), .A2(n10200), .B1(n15507), .B2(n10767), .ZN(
        n11185) );
  INV_X1 U14141 ( .A(n11185), .ZN(n11186) );
  NAND2_X1 U14142 ( .A1(n11184), .A2(n11186), .ZN(n11187) );
  AOI21_X1 U14143 ( .B1(n11189), .B2(n11188), .A(n11187), .ZN(n11190) );
  NAND2_X1 U14144 ( .A1(n13252), .A2(n11192), .ZN(n11193) );
  NAND2_X1 U14145 ( .A1(n11194), .A2(n11193), .ZN(n15329) );
  INV_X1 U14146 ( .A(n11194), .ZN(n11196) );
  NAND2_X1 U14147 ( .A1(n15828), .A2(n19697), .ZN(n19848) );
  NAND2_X1 U14148 ( .A1(n18853), .A2(n19691), .ZN(n11195) );
  OR2_X2 U14149 ( .A1(n19848), .A2(n11195), .ZN(n19089) );
  NAND2_X1 U14150 ( .A1(n11196), .A2(n19089), .ZN(n16305) );
  NAND2_X1 U14151 ( .A1(n16319), .A2(n16305), .ZN(n11207) );
  NAND3_X1 U14152 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n11256) );
  NAND2_X1 U14153 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16298) );
  NOR3_X1 U14154 ( .A1(n13550), .A2(n13717), .A3(n13539), .ZN(n15469) );
  NAND2_X1 U14155 ( .A1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n15469), .ZN(
        n15452) );
  NAND2_X1 U14156 ( .A1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n11198) );
  INV_X1 U14157 ( .A(n11198), .ZN(n12864) );
  OR2_X1 U14158 ( .A1(n15329), .A2(n12864), .ZN(n11197) );
  AND2_X1 U14159 ( .A1(n11197), .A2(n16305), .ZN(n12722) );
  NAND2_X1 U14160 ( .A1(n12721), .A2(n11198), .ZN(n12729) );
  INV_X1 U14161 ( .A(n12729), .ZN(n11209) );
  NOR2_X1 U14162 ( .A1(n15329), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12719) );
  NOR2_X1 U14163 ( .A1(n11209), .A2(n12719), .ZN(n11199) );
  NAND2_X1 U14164 ( .A1(n12722), .A2(n11199), .ZN(n11200) );
  AOI221_X1 U14165 ( .B1(n16298), .B2(n11207), .C1(n15452), .C2(n11207), .A(
        n15465), .ZN(n15408) );
  INV_X1 U14166 ( .A(n11201), .ZN(n15296) );
  NAND2_X1 U14167 ( .A1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15277) );
  NOR2_X1 U14168 ( .A1(n15277), .A2(n15260), .ZN(n11202) );
  NAND2_X1 U14169 ( .A1(n15296), .A2(n11202), .ZN(n11210) );
  INV_X1 U14170 ( .A(n11210), .ZN(n11203) );
  OR2_X1 U14171 ( .A1(n16319), .A2(n11203), .ZN(n11204) );
  NAND2_X1 U14172 ( .A1(n15408), .A2(n11204), .ZN(n15283) );
  AND2_X1 U14173 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11208) );
  NOR2_X1 U14174 ( .A1(n16319), .A2(n11208), .ZN(n11205) );
  INV_X1 U14175 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15067) );
  NAND2_X1 U14176 ( .A1(n15241), .A2(n11207), .ZN(n15234) );
  NAND2_X1 U14177 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n11213) );
  NAND2_X1 U14178 ( .A1(n11207), .A2(n11213), .ZN(n11206) );
  NAND2_X1 U14179 ( .A1(n15234), .A2(n11206), .ZN(n15213) );
  AOI21_X1 U14180 ( .B1(n11207), .B2(n11256), .A(n15213), .ZN(n11259) );
  OR2_X1 U14181 ( .A1(n11259), .A2(n11257), .ZN(n11215) );
  INV_X1 U14182 ( .A(n11208), .ZN(n11212) );
  NAND2_X1 U14183 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n12864), .ZN(
        n12730) );
  AOI211_X1 U14184 ( .C1(n12730), .C2(n15333), .A(n11209), .B(n16319), .ZN(
        n13389) );
  INV_X1 U14185 ( .A(n13389), .ZN(n15471) );
  NAND3_X1 U14186 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A3(n16299), .ZN(n15291) );
  NOR2_X1 U14187 ( .A1(n15291), .A2(n11210), .ZN(n15267) );
  INV_X1 U14188 ( .A(n15267), .ZN(n11211) );
  NOR2_X1 U14189 ( .A1(n11212), .A2(n11211), .ZN(n15242) );
  NAND2_X1 U14190 ( .A1(n15242), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15230) );
  NOR3_X1 U14191 ( .A1(n15195), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n11256), .ZN(n11214) );
  INV_X1 U14192 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n19832) );
  NOR2_X1 U14193 ( .A1(n19089), .A2(n19832), .ZN(n15006) );
  AOI21_X1 U14194 ( .B1(n16136), .B2(n16306), .A(n11216), .ZN(n11217) );
  NOR2_X1 U14195 ( .A1(n11219), .A2(n11218), .ZN(n11220) );
  NAND2_X1 U14196 ( .A1(n11237), .A2(n11222), .ZN(n11224) );
  XOR2_X1 U14197 ( .A(n11224), .B(n11223), .Z(n11279) );
  NOR2_X1 U14198 ( .A1(n15022), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11225) );
  OR2_X2 U14199 ( .A1(n11264), .A2(n11225), .ZN(n11269) );
  OR2_X1 U14200 ( .A1(n14775), .A2(n11226), .ZN(n11227) );
  NOR2_X1 U14201 ( .A1(n15195), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15207) );
  NOR2_X1 U14202 ( .A1(n15213), .A2(n15207), .ZN(n15201) );
  XNOR2_X1 U14203 ( .A(n14873), .B(n9736), .ZN(n16144) );
  OAI21_X1 U14204 ( .B1(n15194), .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n11228) );
  OAI21_X1 U14205 ( .B1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A(n11228), .ZN(n11229) );
  INV_X2 U14206 ( .A(n19089), .ZN(n19069) );
  NAND2_X1 U14207 ( .A1(n19069), .A2(P2_REIP_REG_29__SCAN_IN), .ZN(n11274) );
  OAI21_X1 U14208 ( .B1(n15195), .B2(n11229), .A(n11274), .ZN(n11230) );
  AOI21_X1 U14209 ( .B1(n16306), .B2(n16144), .A(n11230), .ZN(n11231) );
  OAI21_X1 U14210 ( .B1(n15201), .B2(n11232), .A(n11231), .ZN(n11233) );
  AOI21_X1 U14211 ( .B1(n16145), .B2(n16316), .A(n11233), .ZN(n11234) );
  OAI21_X1 U14212 ( .B1(n11269), .B2(n16312), .A(n11234), .ZN(n11235) );
  OAI21_X1 U14213 ( .B1(n11279), .B2(n16310), .A(n11236), .ZN(P2_U3017) );
  OAI211_X2 U14214 ( .C1(n11240), .C2(n11239), .A(n11238), .B(n11237), .ZN(
        n11246) );
  NOR2_X1 U14215 ( .A1(n11241), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n11242) );
  MUX2_X1 U14216 ( .A(n11243), .B(n11242), .S(n11687), .Z(n16121) );
  NAND2_X1 U14217 ( .A1(n16121), .A2(n10506), .ZN(n11244) );
  XNOR2_X1 U14218 ( .A(n11244), .B(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11245) );
  XNOR2_X1 U14219 ( .A(n11246), .B(n11245), .ZN(n14178) );
  INV_X1 U14220 ( .A(P2_EBX_REG_31__SCAN_IN), .ZN(n16123) );
  AOI22_X1 U14221 ( .A1(n10863), .A2(P2_REIP_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n11249) );
  OAI21_X1 U14222 ( .B1(n11250), .B2(n16123), .A(n11249), .ZN(n11251) );
  AOI21_X1 U14223 ( .B1(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n10856), .A(
        n11251), .ZN(n11252) );
  XNOR2_X1 U14224 ( .A(n11253), .B(n11252), .ZN(n16127) );
  INV_X1 U14225 ( .A(n16127), .ZN(n14174) );
  AOI222_X1 U14226 ( .A1(n11158), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n10929), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n11167), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n11254) );
  XNOR2_X1 U14227 ( .A(n11255), .B(n11254), .ZN(n19122) );
  INV_X1 U14228 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n16125) );
  NOR2_X1 U14229 ( .A1(n19089), .A2(n16125), .ZN(n14170) );
  NOR4_X1 U14230 ( .A1(n15195), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n11257), .A4(n11256), .ZN(n11258) );
  OAI21_X1 U14231 ( .B1(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16319), .A(
        n11259), .ZN(n11260) );
  NAND2_X1 U14232 ( .A1(n11260), .A2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n11261) );
  OAI211_X1 U14233 ( .C1(n14174), .C2(n15445), .A(n11262), .B(n11261), .ZN(
        n11263) );
  INV_X1 U14234 ( .A(n11263), .ZN(n11266) );
  OAI211_X1 U14235 ( .C1(n14178), .C2(n16310), .A(n11266), .B(n11265), .ZN(
        P2_U3015) );
  NOR2_X1 U14236 ( .A1(n15507), .A2(n18857), .ZN(n11267) );
  NOR2_X2 U14237 ( .A1(n18859), .A2(n14806), .ZN(n16284) );
  NAND2_X1 U14238 ( .A1(n19650), .A2(n19848), .ZN(n19876) );
  NAND2_X1 U14239 ( .A1(n19876), .A2(n18853), .ZN(n11270) );
  AND2_X1 U14240 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19864) );
  INV_X1 U14241 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n11276) );
  INV_X1 U14242 ( .A(n11305), .ZN(n11272) );
  NAND2_X1 U14243 ( .A1(n19896), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n11271) );
  NAND2_X1 U14244 ( .A1(n11272), .A2(n11271), .ZN(n12818) );
  INV_X1 U14245 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16236) );
  INV_X1 U14246 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18904) );
  INV_X1 U14247 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n20917) );
  INV_X1 U14248 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15055) );
  INV_X1 U14249 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16166) );
  INV_X1 U14250 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15023) );
  AOI21_X1 U14251 ( .B1(n11276), .B2(n15025), .A(n15004), .ZN(n16120) );
  NAND2_X1 U14252 ( .A1(n16279), .A2(n16120), .ZN(n11275) );
  OAI211_X1 U14253 ( .C1(n16288), .C2(n11276), .A(n11275), .B(n11274), .ZN(
        n11277) );
  NAND2_X1 U14254 ( .A1(n9656), .A2(n11305), .ZN(n11287) );
  NAND2_X1 U14255 ( .A1(n11281), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n11282) );
  NAND2_X1 U14256 ( .A1(n11282), .A2(n19697), .ZN(n11309) );
  NAND2_X1 U14257 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19544) );
  NAND2_X1 U14258 ( .A1(n19544), .A2(n19863), .ZN(n11284) );
  NAND2_X1 U14259 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19690) );
  INV_X1 U14260 ( .A(n19690), .ZN(n11283) );
  NAND2_X1 U14261 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11283), .ZN(
        n11307) );
  NAND2_X1 U14262 ( .A1(n11284), .A2(n11307), .ZN(n19349) );
  NOR2_X1 U14263 ( .A1(n19349), .A2(n19650), .ZN(n11285) );
  AOI21_X1 U14264 ( .B1(n11309), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n11285), .ZN(n11286) );
  NAND2_X1 U14265 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(
        n11300) );
  NOR2_X1 U14266 ( .A1(n19650), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n11289) );
  AOI21_X1 U14267 ( .B1(n11309), .B2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n11289), .ZN(n11290) );
  NAND2_X1 U14268 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11292) );
  NAND2_X1 U14269 ( .A1(n12878), .A2(n11292), .ZN(n11298) );
  INV_X1 U14270 ( .A(n11292), .ZN(n11293) );
  NAND2_X1 U14271 ( .A1(n15483), .A2(n11293), .ZN(n11294) );
  NAND2_X1 U14272 ( .A1(n11309), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11295) );
  NAND2_X1 U14273 ( .A1(n19873), .A2(n19880), .ZN(n19454) );
  AND2_X1 U14274 ( .A1(n19544), .A2(n19454), .ZN(n19348) );
  NAND2_X1 U14275 ( .A1(n19348), .A2(n19844), .ZN(n19516) );
  NAND2_X1 U14276 ( .A1(n11295), .A2(n19516), .ZN(n11296) );
  INV_X1 U14277 ( .A(n11298), .ZN(n11299) );
  AOI21_X2 U14278 ( .B1(n12856), .B2(n12855), .A(n11299), .ZN(n12873) );
  NAND2_X1 U14279 ( .A1(n12872), .A2(n12873), .ZN(n11304) );
  INV_X1 U14280 ( .A(n11300), .ZN(n11301) );
  NAND2_X1 U14281 ( .A1(n11302), .A2(n11301), .ZN(n11303) );
  INV_X1 U14282 ( .A(n11307), .ZN(n11306) );
  NAND2_X1 U14283 ( .A1(n11306), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19687) );
  NAND2_X1 U14284 ( .A1(n19856), .A2(n11307), .ZN(n11308) );
  AOI21_X1 U14285 ( .B1(n11309), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19579), .ZN(n11310) );
  NAND2_X1 U14286 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n11313) );
  NAND2_X1 U14287 ( .A1(n12916), .A2(n12915), .ZN(n11317) );
  INV_X1 U14288 ( .A(n11313), .ZN(n11315) );
  AND2_X1 U14289 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n11281), .ZN(
        n11314) );
  INV_X1 U14290 ( .A(n12954), .ZN(n11607) );
  AND2_X1 U14291 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13061) );
  NAND4_X1 U14292 ( .A1(n13062), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A3(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .A4(n13061), .ZN(n11318) );
  NOR2_X1 U14293 ( .A1(n11607), .A2(n11318), .ZN(n11319) );
  NAND2_X1 U14294 ( .A1(n12953), .A2(n11319), .ZN(n13052) );
  NAND2_X1 U14295 ( .A1(n11320), .A2(n13056), .ZN(n13054) );
  NAND2_X1 U14296 ( .A1(n13221), .A2(n13465), .ZN(n13521) );
  NOR2_X2 U14297 ( .A1(n13521), .A2(n11323), .ZN(n13522) );
  INV_X1 U14298 ( .A(n13680), .ZN(n11324) );
  AND2_X2 U14299 ( .A1(n13522), .A2(n11324), .ZN(n13625) );
  NAND2_X1 U14300 ( .A1(n11464), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11326) );
  NAND2_X1 U14301 ( .A1(n10350), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11325) );
  OAI211_X1 U14302 ( .C1(n11327), .C2(n10480), .A(n11326), .B(n11325), .ZN(
        n11330) );
  INV_X1 U14303 ( .A(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11328) );
  OAI22_X1 U14304 ( .A1(n11470), .A2(n11504), .B1(n11469), .B2(n11328), .ZN(
        n11329) );
  NOR2_X1 U14305 ( .A1(n11330), .A2(n11329), .ZN(n11342) );
  AOI22_X1 U14306 ( .A1(n11368), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n11473), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11341) );
  INV_X1 U14307 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11333) );
  AOI22_X1 U14308 ( .A1(n10448), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10408), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11332) );
  NAND2_X1 U14309 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11331) );
  OAI211_X1 U14310 ( .C1(n11477), .C2(n11333), .A(n11332), .B(n11331), .ZN(
        n11338) );
  NAND2_X1 U14311 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11335) );
  NAND2_X1 U14312 ( .A1(n11478), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11334) );
  OAI211_X1 U14313 ( .C1(n10473), .C2(n11336), .A(n11335), .B(n11334), .ZN(
        n11337) );
  NOR2_X1 U14314 ( .A1(n11338), .A2(n11337), .ZN(n11340) );
  AOI22_X1 U14315 ( .A1(n10407), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10403), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11339) );
  NAND4_X1 U14316 ( .A1(n11342), .A2(n11341), .A3(n11340), .A4(n11339), .ZN(
        n13629) );
  AND2_X2 U14317 ( .A1(n13625), .A2(n13629), .ZN(n13627) );
  NAND2_X1 U14318 ( .A1(n11464), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11344) );
  NAND2_X1 U14319 ( .A1(n10350), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11343) );
  OAI211_X1 U14320 ( .C1(n10480), .C2(n11345), .A(n11344), .B(n11343), .ZN(
        n11349) );
  INV_X1 U14321 ( .A(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11346) );
  OAI22_X1 U14322 ( .A1(n11347), .A2(n11470), .B1(n11469), .B2(n11346), .ZN(
        n11348) );
  NOR2_X1 U14323 ( .A1(n11349), .A2(n11348), .ZN(n11361) );
  AOI22_X1 U14324 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11368), .B1(
        n11473), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11360) );
  AOI22_X1 U14325 ( .A1(n10448), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n10408), .ZN(n11351) );
  NAND2_X1 U14326 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11350) );
  OAI211_X1 U14327 ( .C1(n11477), .C2(n11352), .A(n11351), .B(n11350), .ZN(
        n11357) );
  INV_X1 U14328 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11355) );
  NAND2_X1 U14329 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11354) );
  NAND2_X1 U14330 ( .A1(n11478), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11353) );
  OAI211_X1 U14331 ( .C1(n10473), .C2(n11355), .A(n11354), .B(n11353), .ZN(
        n11356) );
  NOR2_X1 U14332 ( .A1(n11357), .A2(n11356), .ZN(n11359) );
  AOI22_X1 U14333 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n10407), .B1(
        n10403), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11358) );
  NAND4_X1 U14334 ( .A1(n11361), .A2(n11360), .A3(n11359), .A4(n11358), .ZN(
        n14858) );
  INV_X1 U14335 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11364) );
  NAND2_X1 U14336 ( .A1(n11464), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(
        n11363) );
  NAND2_X1 U14337 ( .A1(n10350), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(
        n11362) );
  OAI211_X1 U14338 ( .C1(n10480), .C2(n11364), .A(n11363), .B(n11362), .ZN(
        n11367) );
  INV_X1 U14339 ( .A(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11365) );
  OAI22_X1 U14340 ( .A1(n11551), .A2(n11470), .B1(n11469), .B2(n11365), .ZN(
        n11366) );
  NOR2_X1 U14341 ( .A1(n11367), .A2(n11366), .ZN(n11382) );
  INV_X1 U14342 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11369) );
  INV_X1 U14343 ( .A(n11368), .ZN(n11449) );
  INV_X1 U14344 ( .A(n11473), .ZN(n11448) );
  OAI22_X1 U14345 ( .A1(n11369), .A2(n11449), .B1(n11448), .B2(n11549), .ZN(
        n11370) );
  INV_X1 U14346 ( .A(n11370), .ZN(n11381) );
  INV_X1 U14347 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11373) );
  AOI22_X1 U14348 ( .A1(n10448), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n10408), .ZN(n11372) );
  NAND2_X1 U14349 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n11371) );
  OAI211_X1 U14350 ( .C1(n11477), .C2(n11373), .A(n11372), .B(n11371), .ZN(
        n11378) );
  NAND2_X1 U14351 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(
        n11375) );
  NAND2_X1 U14352 ( .A1(n11478), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(
        n11374) );
  OAI211_X1 U14353 ( .C1(n10473), .C2(n11376), .A(n11375), .B(n11374), .ZN(
        n11377) );
  NOR2_X1 U14354 ( .A1(n11378), .A2(n11377), .ZN(n11380) );
  AOI22_X1 U14355 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n11399), .B1(
        n10403), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11379) );
  NAND4_X1 U14356 ( .A1(n11382), .A2(n11381), .A3(n11380), .A4(n11379), .ZN(
        n14853) );
  INV_X1 U14357 ( .A(n14853), .ZN(n11383) );
  NAND2_X1 U14358 ( .A1(n11464), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11385) );
  NAND2_X1 U14359 ( .A1(n10350), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(
        n11384) );
  OAI211_X1 U14360 ( .C1(n10480), .C2(n11386), .A(n11385), .B(n11384), .ZN(
        n11390) );
  OAI22_X1 U14361 ( .A1(n11388), .A2(n11470), .B1(n11469), .B2(n11387), .ZN(
        n11389) );
  NOR2_X1 U14362 ( .A1(n11390), .A2(n11389), .ZN(n11403) );
  AOI22_X1 U14363 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11368), .B1(
        n11473), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11402) );
  AOI22_X1 U14364 ( .A1(n10448), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n10408), .ZN(n11392) );
  NAND2_X1 U14365 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n11391) );
  OAI211_X1 U14366 ( .C1(n11477), .C2(n11393), .A(n11392), .B(n11391), .ZN(
        n11398) );
  NAND2_X1 U14367 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(
        n11395) );
  NAND2_X1 U14368 ( .A1(n11478), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(
        n11394) );
  OAI211_X1 U14369 ( .C1(n10473), .C2(n11396), .A(n11395), .B(n11394), .ZN(
        n11397) );
  NOR2_X1 U14370 ( .A1(n11398), .A2(n11397), .ZN(n11401) );
  AOI22_X1 U14371 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n11399), .B1(
        n10403), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11400) );
  AND4_X1 U14372 ( .A1(n11403), .A2(n11402), .A3(n11401), .A4(n11400), .ZN(
        n14843) );
  NAND2_X1 U14373 ( .A1(n11464), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11406) );
  NAND2_X1 U14374 ( .A1(n10350), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11405) );
  OAI211_X1 U14375 ( .C1(n10480), .C2(n11407), .A(n11406), .B(n11405), .ZN(
        n11410) );
  OAI22_X1 U14376 ( .A1(n11599), .A2(n11470), .B1(n11469), .B2(n11408), .ZN(
        n11409) );
  NOR2_X1 U14377 ( .A1(n11410), .A2(n11409), .ZN(n11422) );
  AOI22_X1 U14378 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11473), .B1(
        n11368), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11421) );
  INV_X1 U14379 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11413) );
  AOI22_X1 U14380 ( .A1(n10448), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n10408), .ZN(n11412) );
  NAND2_X1 U14381 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11411) );
  OAI211_X1 U14382 ( .C1(n11477), .C2(n11413), .A(n11412), .B(n11411), .ZN(
        n11418) );
  NAND2_X1 U14383 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11415) );
  NAND2_X1 U14384 ( .A1(n11478), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11414) );
  OAI211_X1 U14385 ( .C1(n10473), .C2(n11416), .A(n11415), .B(n11414), .ZN(
        n11417) );
  NOR2_X1 U14386 ( .A1(n11418), .A2(n11417), .ZN(n11420) );
  AOI22_X1 U14387 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10407), .B1(
        n10403), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11419) );
  NAND4_X1 U14388 ( .A1(n11422), .A2(n11421), .A3(n11420), .A4(n11419), .ZN(
        n14837) );
  NAND2_X1 U14389 ( .A1(n11464), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11424) );
  NAND2_X1 U14390 ( .A1(n10350), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11423) );
  OAI211_X1 U14391 ( .C1(n11425), .C2(n10480), .A(n11424), .B(n11423), .ZN(
        n11429) );
  OAI22_X1 U14392 ( .A1(n11470), .A2(n11427), .B1(n11469), .B2(n11426), .ZN(
        n11428) );
  NOR2_X1 U14393 ( .A1(n11429), .A2(n11428), .ZN(n11440) );
  AOI22_X1 U14394 ( .A1(n11368), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11473), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11439) );
  AOI22_X1 U14395 ( .A1(n10448), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10408), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11431) );
  NAND2_X1 U14396 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11430) );
  OAI211_X1 U14397 ( .C1(n11477), .C2(n20909), .A(n11431), .B(n11430), .ZN(
        n11436) );
  NAND2_X1 U14398 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11433) );
  NAND2_X1 U14399 ( .A1(n11478), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11432) );
  OAI211_X1 U14400 ( .C1(n10473), .C2(n11434), .A(n11433), .B(n11432), .ZN(
        n11435) );
  NOR2_X1 U14401 ( .A1(n11436), .A2(n11435), .ZN(n11438) );
  AOI22_X1 U14402 ( .A1(n10407), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10403), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11437) );
  NAND4_X1 U14403 ( .A1(n11440), .A2(n11439), .A3(n11438), .A4(n11437), .ZN(
        n14830) );
  NAND2_X1 U14404 ( .A1(n11464), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11442) );
  NAND2_X1 U14405 ( .A1(n10350), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11441) );
  OAI211_X1 U14406 ( .C1(n11443), .C2(n10480), .A(n11442), .B(n11441), .ZN(
        n11446) );
  OAI22_X1 U14407 ( .A1(n11470), .A2(n11638), .B1(n11469), .B2(n11444), .ZN(
        n11445) );
  NOR2_X1 U14408 ( .A1(n11446), .A2(n11445), .ZN(n11462) );
  OAI22_X1 U14409 ( .A1(n11639), .A2(n11449), .B1(n11448), .B2(n11447), .ZN(
        n11450) );
  INV_X1 U14410 ( .A(n11450), .ZN(n11461) );
  AOI22_X1 U14411 ( .A1(n10448), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10408), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11452) );
  NAND2_X1 U14412 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11451) );
  OAI211_X1 U14413 ( .C1(n11477), .C2(n11453), .A(n11452), .B(n11451), .ZN(
        n11458) );
  NAND2_X1 U14414 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11455) );
  NAND2_X1 U14415 ( .A1(n11478), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11454) );
  OAI211_X1 U14416 ( .C1(n10473), .C2(n11456), .A(n11455), .B(n11454), .ZN(
        n11457) );
  NOR2_X1 U14417 ( .A1(n11458), .A2(n11457), .ZN(n11460) );
  AOI22_X1 U14418 ( .A1(n10407), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10403), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11459) );
  AND4_X1 U14419 ( .A1(n11462), .A2(n11461), .A3(n11460), .A4(n11459), .ZN(
        n14826) );
  INV_X1 U14420 ( .A(n14826), .ZN(n11463) );
  INV_X1 U14421 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11467) );
  NAND2_X1 U14422 ( .A1(n11464), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n11466) );
  NAND2_X1 U14423 ( .A1(n10350), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n11465) );
  OAI211_X1 U14424 ( .C1(n11467), .C2(n10480), .A(n11466), .B(n11465), .ZN(
        n11472) );
  INV_X1 U14425 ( .A(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11661) );
  INV_X1 U14426 ( .A(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11468) );
  OAI22_X1 U14427 ( .A1(n11661), .A2(n11470), .B1(n11469), .B2(n11468), .ZN(
        n11471) );
  NOR2_X1 U14428 ( .A1(n11472), .A2(n11471), .ZN(n11487) );
  AOI22_X1 U14429 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n11368), .B1(
        n11473), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11486) );
  AOI22_X1 U14430 ( .A1(n10448), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n10408), .ZN(n11475) );
  NAND2_X1 U14431 ( .A1(n10380), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n11474) );
  OAI211_X1 U14432 ( .C1(n11477), .C2(n11476), .A(n11475), .B(n11474), .ZN(
        n11483) );
  NAND2_X1 U14433 ( .A1(n10351), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n11480) );
  NAND2_X1 U14434 ( .A1(n11478), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n11479) );
  OAI211_X1 U14435 ( .C1(n10473), .C2(n11481), .A(n11480), .B(n11479), .ZN(
        n11482) );
  NOR2_X1 U14436 ( .A1(n11483), .A2(n11482), .ZN(n11485) );
  AOI22_X1 U14437 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n10407), .B1(
        n10403), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11484) );
  NAND4_X1 U14438 ( .A1(n11487), .A2(n11486), .A3(n11485), .A4(n11484), .ZN(
        n11512) );
  AOI22_X1 U14439 ( .A1(n9649), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11671), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11501) );
  INV_X1 U14440 ( .A(n10156), .ZN(n11490) );
  AOI22_X1 U14441 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n9632), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11500) );
  INV_X1 U14442 ( .A(n11645), .ZN(n11666) );
  INV_X1 U14443 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11496) );
  OR2_X1 U14444 ( .A1(n11664), .A2(n11491), .ZN(n11495) );
  INV_X1 U14445 ( .A(n11492), .ZN(n11494) );
  NAND2_X1 U14446 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11493) );
  NAND2_X1 U14447 ( .A1(n11494), .A2(n11493), .ZN(n11662) );
  OAI211_X1 U14448 ( .C1(n11666), .C2(n11496), .A(n11495), .B(n11662), .ZN(
        n11497) );
  INV_X1 U14449 ( .A(n11497), .ZN(n11499) );
  INV_X1 U14450 ( .A(n11668), .ZN(n11657) );
  AOI22_X1 U14451 ( .A1(n11657), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10066), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n11498) );
  NAND4_X1 U14452 ( .A1(n11501), .A2(n11500), .A3(n11499), .A4(n11498), .ZN(
        n11511) );
  AOI22_X1 U14453 ( .A1(n9649), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n11671), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11509) );
  AOI22_X1 U14454 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9632), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11508) );
  OR2_X1 U14455 ( .A1(n11664), .A2(n11502), .ZN(n11503) );
  INV_X1 U14456 ( .A(n11662), .ZN(n11623) );
  OAI211_X1 U14457 ( .C1(n11666), .C2(n11504), .A(n11503), .B(n11623), .ZN(
        n11505) );
  INV_X1 U14458 ( .A(n11505), .ZN(n11507) );
  AOI22_X1 U14459 ( .A1(n11657), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10066), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11506) );
  NAND4_X1 U14460 ( .A1(n11509), .A2(n11508), .A3(n11507), .A4(n11506), .ZN(
        n11510) );
  AND2_X1 U14461 ( .A1(n11511), .A2(n11510), .ZN(n11517) );
  AND2_X1 U14462 ( .A1(n11512), .A2(n11517), .ZN(n11538) );
  NAND2_X1 U14463 ( .A1(n11538), .A2(n14806), .ZN(n11516) );
  INV_X1 U14464 ( .A(n11512), .ZN(n11514) );
  NAND2_X1 U14465 ( .A1(n14806), .A2(n11517), .ZN(n11513) );
  NAND2_X1 U14466 ( .A1(n11514), .A2(n11513), .ZN(n11515) );
  NAND2_X1 U14467 ( .A1(n11518), .A2(n11517), .ZN(n14820) );
  AND2_X2 U14468 ( .A1(n11519), .A2(n9731), .ZN(n11520) );
  AOI22_X1 U14469 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11527) );
  AOI22_X1 U14470 ( .A1(n10305), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11671), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n11526) );
  AOI22_X1 U14471 ( .A1(n11657), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n9632), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11525) );
  NAND2_X1 U14472 ( .A1(n10066), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11521) );
  OAI211_X1 U14473 ( .C1(n11664), .C2(n11522), .A(n11521), .B(n11662), .ZN(
        n11523) );
  INV_X1 U14474 ( .A(n11523), .ZN(n11524) );
  NAND4_X1 U14475 ( .A1(n11527), .A2(n11526), .A3(n11525), .A4(n11524), .ZN(
        n11536) );
  AOI22_X1 U14476 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11534) );
  AOI22_X1 U14477 ( .A1(n9649), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n11671), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11533) );
  AOI22_X1 U14478 ( .A1(n11657), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9632), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11532) );
  NAND2_X1 U14479 ( .A1(n10066), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11528) );
  OAI211_X1 U14480 ( .C1(n11664), .C2(n11529), .A(n11528), .B(n11623), .ZN(
        n11530) );
  INV_X1 U14481 ( .A(n11530), .ZN(n11531) );
  NAND4_X1 U14482 ( .A1(n11534), .A2(n11533), .A3(n11532), .A4(n11531), .ZN(
        n11535) );
  NAND2_X1 U14483 ( .A1(n11536), .A2(n11535), .ZN(n14805) );
  INV_X1 U14484 ( .A(n14805), .ZN(n11539) );
  INV_X1 U14485 ( .A(n11538), .ZN(n11537) );
  OR2_X1 U14486 ( .A1(n11537), .A2(n14805), .ZN(n11541) );
  OAI211_X1 U14487 ( .C1(n11538), .C2(n11539), .A(n12954), .B(n11541), .ZN(
        n14804) );
  INV_X1 U14488 ( .A(n14820), .ZN(n11540) );
  INV_X1 U14489 ( .A(n11541), .ZN(n11559) );
  AOI22_X1 U14490 ( .A1(n10305), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11671), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11548) );
  AOI22_X1 U14491 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9632), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11547) );
  INV_X1 U14492 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11543) );
  OR2_X1 U14493 ( .A1(n11664), .A2(n11369), .ZN(n11542) );
  OAI211_X1 U14494 ( .C1(n11666), .C2(n11543), .A(n11542), .B(n11662), .ZN(
        n11544) );
  INV_X1 U14495 ( .A(n11544), .ZN(n11546) );
  AOI22_X1 U14496 ( .A1(n11657), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10066), .B2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11545) );
  NAND4_X1 U14497 ( .A1(n11548), .A2(n11547), .A3(n11546), .A4(n11545), .ZN(
        n11558) );
  AOI22_X1 U14498 ( .A1(n9649), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11671), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11556) );
  AOI22_X1 U14499 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10156), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11555) );
  OR2_X1 U14500 ( .A1(n11664), .A2(n11549), .ZN(n11550) );
  OAI211_X1 U14501 ( .C1(n11666), .C2(n11551), .A(n11550), .B(n11623), .ZN(
        n11552) );
  INV_X1 U14502 ( .A(n11552), .ZN(n11554) );
  AOI22_X1 U14503 ( .A1(n11657), .A2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n10066), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11553) );
  NAND4_X1 U14504 ( .A1(n11556), .A2(n11555), .A3(n11554), .A4(n11553), .ZN(
        n11557) );
  AND2_X1 U14505 ( .A1(n11558), .A2(n11557), .ZN(n11560) );
  NAND2_X1 U14506 ( .A1(n11559), .A2(n11560), .ZN(n11582) );
  OAI211_X1 U14507 ( .C1(n11559), .C2(n11560), .A(n12954), .B(n11582), .ZN(
        n11563) );
  INV_X1 U14508 ( .A(n11560), .ZN(n11561) );
  NOR2_X1 U14509 ( .A1(n14806), .A2(n11561), .ZN(n14797) );
  NAND2_X1 U14510 ( .A1(n14798), .A2(n14797), .ZN(n14796) );
  INV_X1 U14511 ( .A(n11562), .ZN(n11564) );
  AOI22_X1 U14512 ( .A1(n10305), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11657), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n11572) );
  AOI22_X1 U14513 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11671), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11571) );
  AOI22_X1 U14514 ( .A1(n11645), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10156), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11570) );
  NAND2_X1 U14515 ( .A1(n10066), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(
        n11566) );
  OAI211_X1 U14516 ( .C1(n11664), .C2(n11567), .A(n11566), .B(n11662), .ZN(
        n11568) );
  INV_X1 U14517 ( .A(n11568), .ZN(n11569) );
  NAND4_X1 U14518 ( .A1(n11572), .A2(n11571), .A3(n11570), .A4(n11569), .ZN(
        n11581) );
  AOI22_X1 U14519 ( .A1(n11657), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11645), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11579) );
  AOI22_X1 U14520 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11671), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11578) );
  AOI22_X1 U14521 ( .A1(n9649), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10156), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11577) );
  NAND2_X1 U14522 ( .A1(n10066), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(
        n11573) );
  OAI211_X1 U14523 ( .C1(n11664), .C2(n11574), .A(n11573), .B(n11623), .ZN(
        n11575) );
  INV_X1 U14524 ( .A(n11575), .ZN(n11576) );
  NAND4_X1 U14525 ( .A1(n11579), .A2(n11578), .A3(n11577), .A4(n11576), .ZN(
        n11580) );
  NAND2_X1 U14526 ( .A1(n11581), .A2(n11580), .ZN(n11584) );
  AOI21_X1 U14527 ( .B1(n11582), .B2(n11584), .A(n11607), .ZN(n11583) );
  OR2_X1 U14528 ( .A1(n11582), .A2(n11584), .ZN(n11608) );
  NAND2_X1 U14529 ( .A1(n11583), .A2(n11608), .ZN(n11585) );
  XNOR2_X2 U14530 ( .A(n11587), .B(n11585), .ZN(n14789) );
  NOR2_X1 U14531 ( .A1(n14806), .A2(n11584), .ZN(n14788) );
  INV_X1 U14532 ( .A(n11585), .ZN(n11586) );
  AOI21_X2 U14533 ( .B1(n14789), .B2(n14788), .A(n11588), .ZN(n11613) );
  AOI22_X1 U14534 ( .A1(n10305), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n11671), .B2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n11596) );
  AOI22_X1 U14535 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10156), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11595) );
  INV_X1 U14536 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11591) );
  INV_X1 U14537 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11589) );
  OR2_X1 U14538 ( .A1(n11664), .A2(n11589), .ZN(n11590) );
  OAI211_X1 U14539 ( .C1(n11666), .C2(n11591), .A(n11590), .B(n11662), .ZN(
        n11592) );
  INV_X1 U14540 ( .A(n11592), .ZN(n11594) );
  AOI22_X1 U14541 ( .A1(n11657), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10066), .B2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11593) );
  NAND4_X1 U14542 ( .A1(n11596), .A2(n11595), .A3(n11594), .A4(n11593), .ZN(
        n11606) );
  AOI22_X1 U14543 ( .A1(n9649), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11671), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11604) );
  AOI22_X1 U14544 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9632), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11603) );
  OR2_X1 U14545 ( .A1(n11664), .A2(n11597), .ZN(n11598) );
  OAI211_X1 U14546 ( .C1(n11666), .C2(n11599), .A(n11598), .B(n11623), .ZN(
        n11600) );
  INV_X1 U14547 ( .A(n11600), .ZN(n11602) );
  AOI22_X1 U14548 ( .A1(n11657), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10066), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n11601) );
  NAND4_X1 U14549 ( .A1(n11604), .A2(n11603), .A3(n11602), .A4(n11601), .ZN(
        n11605) );
  NAND2_X1 U14550 ( .A1(n11606), .A2(n11605), .ZN(n11609) );
  AOI21_X1 U14551 ( .B1(n11608), .B2(n11609), .A(n11607), .ZN(n11611) );
  INV_X1 U14552 ( .A(n11608), .ZN(n11610) );
  INV_X1 U14553 ( .A(n11609), .ZN(n11612) );
  NAND2_X1 U14554 ( .A1(n11610), .A2(n11612), .ZN(n14771) );
  NAND2_X1 U14555 ( .A1(n11611), .A2(n14771), .ZN(n11614) );
  NAND2_X1 U14556 ( .A1(n11518), .A2(n11612), .ZN(n14781) );
  INV_X1 U14557 ( .A(n11615), .ZN(n11641) );
  OAI21_X1 U14558 ( .B1(n11664), .B2(n13020), .A(n11662), .ZN(n11619) );
  OAI22_X1 U14559 ( .A1(n11668), .A2(n11617), .B1(n11666), .B2(n11616), .ZN(
        n11618) );
  AOI211_X1 U14560 ( .C1(n10066), .C2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A(
        n11619), .B(n11618), .ZN(n11622) );
  AOI22_X1 U14561 ( .A1(n10305), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11671), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n11621) );
  AOI22_X1 U14562 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9632), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11620) );
  NAND3_X1 U14563 ( .A1(n11622), .A2(n11621), .A3(n11620), .ZN(n11633) );
  OAI21_X1 U14564 ( .B1(n11664), .B2(n11624), .A(n11623), .ZN(n11628) );
  OAI22_X1 U14565 ( .A1(n11490), .A2(n11626), .B1(n11641), .B2(n11625), .ZN(
        n11627) );
  AOI211_X1 U14566 ( .C1(n11645), .C2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A(
        n11628), .B(n11627), .ZN(n11631) );
  AOI22_X1 U14567 ( .A1(n9649), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11671), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11630) );
  AOI22_X1 U14568 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11657), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11629) );
  NAND3_X1 U14569 ( .A1(n11631), .A2(n11630), .A3(n11629), .ZN(n11632) );
  AOI22_X1 U14570 ( .A1(n9649), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11671), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11635) );
  AOI22_X1 U14571 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10156), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11634) );
  NAND2_X1 U14572 ( .A1(n11635), .A2(n11634), .ZN(n11651) );
  AOI22_X1 U14573 ( .A1(n11657), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10066), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11637) );
  AOI21_X1 U14574 ( .B1(n11658), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n11662), .ZN(n11636) );
  OAI211_X1 U14575 ( .C1(n11666), .C2(n11638), .A(n11637), .B(n11636), .ZN(
        n11650) );
  OAI21_X1 U14576 ( .B1(n11664), .B2(n11639), .A(n11662), .ZN(n11644) );
  OAI22_X1 U14577 ( .A1(n11668), .A2(n11642), .B1(n11641), .B2(n11640), .ZN(
        n11643) );
  AOI211_X1 U14578 ( .C1(n11645), .C2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A(
        n11644), .B(n11643), .ZN(n11648) );
  AOI22_X1 U14579 ( .A1(n10305), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n11671), .B2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11647) );
  AOI22_X1 U14580 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9632), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11646) );
  NAND3_X1 U14581 ( .A1(n11648), .A2(n11647), .A3(n11646), .ZN(n11649) );
  OAI21_X1 U14582 ( .B1(n11651), .B2(n11650), .A(n11649), .ZN(n11653) );
  NOR3_X1 U14583 ( .A1(n14771), .A2(n11518), .A3(n9735), .ZN(n11652) );
  XOR2_X1 U14584 ( .A(n11653), .B(n11652), .Z(n14768) );
  INV_X1 U14585 ( .A(n11652), .ZN(n11654) );
  AOI22_X1 U14586 ( .A1(n10305), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11671), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11656) );
  AOI22_X1 U14587 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n10156), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11655) );
  NAND2_X1 U14588 ( .A1(n11656), .A2(n11655), .ZN(n11678) );
  AOI22_X1 U14589 ( .A1(n11657), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n10066), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11660) );
  AOI21_X1 U14590 ( .B1(n11658), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A(
        n11662), .ZN(n11659) );
  OAI211_X1 U14591 ( .C1(n11666), .C2(n11661), .A(n11660), .B(n11659), .ZN(
        n11677) );
  INV_X1 U14592 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11663) );
  OAI21_X1 U14593 ( .B1(n11664), .B2(n11663), .A(n11662), .ZN(n11670) );
  INV_X1 U14594 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11667) );
  INV_X1 U14595 ( .A(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11665) );
  OAI22_X1 U14596 ( .A1(n11668), .A2(n11667), .B1(n11666), .B2(n11665), .ZN(
        n11669) );
  AOI211_X1 U14597 ( .C1(n10066), .C2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A(
        n11670), .B(n11669), .ZN(n11675) );
  AOI22_X1 U14598 ( .A1(n9649), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11671), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11674) );
  AOI22_X1 U14599 ( .A1(n11672), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9632), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11673) );
  NAND3_X1 U14600 ( .A1(n11675), .A2(n11674), .A3(n11673), .ZN(n11676) );
  OAI21_X1 U14601 ( .B1(n11678), .B2(n11677), .A(n11676), .ZN(n11679) );
  INV_X1 U14602 ( .A(n11679), .ZN(n11680) );
  XNOR2_X1 U14603 ( .A(n11681), .B(n11680), .ZN(n14184) );
  NAND2_X1 U14604 ( .A1(n13281), .A2(n12736), .ZN(n13292) );
  NAND2_X1 U14605 ( .A1(n19899), .A2(n19898), .ZN(n13290) );
  NOR2_X1 U14606 ( .A1(n13292), .A2(n13290), .ZN(n11682) );
  AOI21_X1 U14607 ( .B1(n15479), .B2(n13284), .A(n11682), .ZN(n12797) );
  NAND2_X1 U14608 ( .A1(n11684), .A2(n11683), .ZN(n11685) );
  NAND2_X1 U14609 ( .A1(n12797), .A2(n11685), .ZN(n11686) );
  AND2_X1 U14610 ( .A1(n11687), .A2(n10176), .ZN(n11688) );
  NOR4_X1 U14611 ( .A1(P2_ADDRESS_REG_15__SCAN_IN), .A2(
        P2_ADDRESS_REG_14__SCAN_IN), .A3(P2_ADDRESS_REG_13__SCAN_IN), .A4(
        P2_ADDRESS_REG_12__SCAN_IN), .ZN(n11692) );
  NOR4_X1 U14612 ( .A1(P2_ADDRESS_REG_19__SCAN_IN), .A2(
        P2_ADDRESS_REG_18__SCAN_IN), .A3(P2_ADDRESS_REG_17__SCAN_IN), .A4(
        P2_ADDRESS_REG_16__SCAN_IN), .ZN(n11691) );
  NOR4_X1 U14613 ( .A1(P2_ADDRESS_REG_7__SCAN_IN), .A2(
        P2_ADDRESS_REG_6__SCAN_IN), .A3(P2_ADDRESS_REG_4__SCAN_IN), .A4(
        P2_ADDRESS_REG_3__SCAN_IN), .ZN(n11690) );
  NOR4_X1 U14614 ( .A1(P2_ADDRESS_REG_11__SCAN_IN), .A2(
        P2_ADDRESS_REG_10__SCAN_IN), .A3(P2_ADDRESS_REG_9__SCAN_IN), .A4(
        P2_ADDRESS_REG_8__SCAN_IN), .ZN(n11689) );
  NAND4_X1 U14615 ( .A1(n11692), .A2(n11691), .A3(n11690), .A4(n11689), .ZN(
        n11697) );
  NOR4_X1 U14616 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_5__SCAN_IN), .A4(
        P2_ADDRESS_REG_28__SCAN_IN), .ZN(n11695) );
  NOR4_X1 U14617 ( .A1(P2_ADDRESS_REG_23__SCAN_IN), .A2(
        P2_ADDRESS_REG_22__SCAN_IN), .A3(P2_ADDRESS_REG_21__SCAN_IN), .A4(
        P2_ADDRESS_REG_20__SCAN_IN), .ZN(n11694) );
  NOR4_X1 U14618 ( .A1(P2_ADDRESS_REG_27__SCAN_IN), .A2(
        P2_ADDRESS_REG_26__SCAN_IN), .A3(P2_ADDRESS_REG_25__SCAN_IN), .A4(
        P2_ADDRESS_REG_24__SCAN_IN), .ZN(n11693) );
  INV_X1 U14619 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19782) );
  NAND4_X1 U14620 ( .A1(n11695), .A2(n11694), .A3(n11693), .A4(n19782), .ZN(
        n11696) );
  MUX2_X1 U14621 ( .A(BUF1_REG_14__SCAN_IN), .B(BUF2_REG_14__SCAN_IN), .S(
        n15508), .Z(n19203) );
  INV_X1 U14622 ( .A(n16136), .ZN(n11699) );
  INV_X1 U14623 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n11698) );
  OAI22_X1 U14624 ( .A1(n11699), .A2(n19153), .B1(n19152), .B2(n11698), .ZN(
        n11700) );
  AOI21_X1 U14625 ( .B1(n15000), .B2(n19203), .A(n11700), .ZN(n11703) );
  NOR2_X2 U14626 ( .A1(n12922), .A2(n15510), .ZN(n19121) );
  NOR2_X2 U14627 ( .A1(n12922), .A2(n15508), .ZN(n19123) );
  AOI22_X1 U14628 ( .A1(n19121), .A2(BUF2_REG_30__SCAN_IN), .B1(n19123), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n11702) );
  OAI21_X1 U14629 ( .B1(n14184), .B2(n15002), .A(n11704), .ZN(P2_U2889) );
  AOI22_X1 U14630 ( .A1(n11755), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11712) );
  AOI22_X1 U14631 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n11771), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11711) );
  INV_X1 U14632 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11708) );
  AOI22_X1 U14633 ( .A1(n12169), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n11869), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11710) );
  AND2_X2 U14634 ( .A1(n11713), .A2(n11715), .ZN(n11777) );
  BUF_X2 U14635 ( .A(n11777), .Z(n12441) );
  AOI22_X1 U14636 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12441), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11709) );
  NAND4_X1 U14637 ( .A1(n11712), .A2(n11711), .A3(n11710), .A4(n11709), .ZN(
        n11721) );
  AOI22_X1 U14638 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11719) );
  AND2_X2 U14639 ( .A1(n11714), .A2(n13201), .ZN(n11824) );
  AOI22_X1 U14640 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n11718) );
  AOI22_X1 U14641 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9650), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11717) );
  AOI22_X1 U14642 ( .A1(n11825), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11874), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11716) );
  NAND4_X1 U14643 ( .A1(n11719), .A2(n11718), .A3(n11717), .A4(n11716), .ZN(
        n11720) );
  BUF_X2 U14644 ( .A(n11882), .Z(n12505) );
  AOI22_X1 U14645 ( .A1(n12505), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11755), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11725) );
  AOI22_X1 U14646 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11887), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n11724) );
  AOI22_X1 U14647 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11723) );
  BUF_X4 U14648 ( .A(n11771), .Z(n12485) );
  AOI22_X1 U14649 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9651), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11722) );
  NAND4_X1 U14650 ( .A1(n11725), .A2(n11724), .A3(n11723), .A4(n11722), .ZN(
        n11731) );
  AOI22_X1 U14651 ( .A1(n9628), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11729) );
  AOI22_X1 U14652 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12169), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n11728) );
  BUF_X4 U14653 ( .A(n11777), .Z(n12484) );
  AOI22_X1 U14654 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11727) );
  AOI22_X1 U14655 ( .A1(n11874), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11869), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11726) );
  NAND4_X1 U14656 ( .A1(n11729), .A2(n11728), .A3(n11727), .A4(n11726), .ZN(
        n11730) );
  OR2_X2 U14657 ( .A1(n11731), .A2(n11730), .ZN(n13352) );
  NAND2_X1 U14658 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(
        n11736) );
  NAND2_X1 U14659 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n11735) );
  NAND2_X1 U14660 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n11734) );
  NAND2_X1 U14661 ( .A1(n9627), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n11733) );
  BUF_X4 U14662 ( .A(n11824), .Z(n12325) );
  NAND2_X1 U14663 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(
        n11741) );
  NAND2_X1 U14664 ( .A1(n11825), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(
        n11740) );
  NAND2_X1 U14665 ( .A1(n11874), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(
        n11739) );
  NAND2_X1 U14666 ( .A1(n9650), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11738) );
  NAND2_X1 U14667 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(
        n11745) );
  NAND2_X1 U14668 ( .A1(n12441), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(
        n11744) );
  NAND2_X1 U14669 ( .A1(n11771), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(
        n11743) );
  NAND2_X1 U14670 ( .A1(n11772), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(
        n11742) );
  NAND2_X1 U14671 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(
        n11749) );
  NAND2_X1 U14672 ( .A1(n11755), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(
        n11748) );
  NAND2_X1 U14673 ( .A1(n12169), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(
        n11747) );
  NAND2_X1 U14674 ( .A1(n11869), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(
        n11746) );
  AOI22_X1 U14675 ( .A1(n12505), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12513), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11759) );
  AOI22_X1 U14676 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11754), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11758) );
  AOI22_X1 U14677 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11824), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11757) );
  AOI22_X1 U14678 ( .A1(n11755), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11756) );
  NAND4_X1 U14679 ( .A1(n11759), .A2(n11758), .A3(n11757), .A4(n11756), .ZN(
        n11766) );
  AOI22_X1 U14680 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n11760), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11764) );
  AOI22_X1 U14681 ( .A1(n12169), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n11869), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11763) );
  AOI22_X1 U14682 ( .A1(n9628), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11762) );
  AOI22_X1 U14683 ( .A1(n9652), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11874), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11761) );
  NAND4_X1 U14684 ( .A1(n11764), .A2(n11763), .A3(n11762), .A4(n11761), .ZN(
        n11765) );
  NAND2_X1 U14685 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11770) );
  NAND2_X1 U14686 ( .A1(n9629), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n11769) );
  NAND2_X1 U14687 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11768) );
  NAND2_X1 U14688 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n11767) );
  NAND2_X1 U14689 ( .A1(n11755), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n11776) );
  NAND2_X1 U14690 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11775) );
  BUF_X2 U14691 ( .A(n11771), .Z(n12511) );
  NAND2_X1 U14692 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11774) );
  NAND2_X1 U14693 ( .A1(n11772), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n11773) );
  NAND2_X1 U14694 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11781) );
  NAND2_X1 U14695 ( .A1(n11777), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n11780) );
  NAND2_X1 U14696 ( .A1(n12169), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n11779) );
  NAND2_X1 U14697 ( .A1(n11869), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11778) );
  NAND2_X1 U14698 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n11785) );
  NAND2_X1 U14699 ( .A1(n11825), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n11784) );
  NAND2_X1 U14700 ( .A1(n9651), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11783) );
  NAND2_X1 U14701 ( .A1(n11874), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11782) );
  OR2_X2 U14702 ( .A1(n11857), .A2(n11790), .ZN(n11854) );
  AOI22_X1 U14703 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11760), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11794) );
  AOI22_X1 U14704 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11793) );
  AOI22_X1 U14705 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11792) );
  AOI22_X1 U14706 ( .A1(n9631), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n11869), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11791) );
  NAND4_X1 U14707 ( .A1(n11794), .A2(n11793), .A3(n11792), .A4(n11791), .ZN(
        n11800) );
  AOI22_X1 U14708 ( .A1(n12505), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12513), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11798) );
  AOI22_X1 U14709 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11797) );
  AOI22_X1 U14710 ( .A1(n11755), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11796) );
  AOI22_X1 U14711 ( .A1(n9652), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n11874), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11795) );
  NAND4_X1 U14712 ( .A1(n11798), .A2(n11797), .A3(n11796), .A4(n11795), .ZN(
        n11799) );
  OR2_X2 U14713 ( .A1(n11800), .A2(n11799), .ZN(n13360) );
  NAND2_X1 U14714 ( .A1(n11854), .A2(n13360), .ZN(n11801) );
  NAND2_X1 U14715 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11806) );
  NAND2_X1 U14716 ( .A1(n9628), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11805) );
  NAND2_X1 U14717 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11804) );
  NAND2_X1 U14718 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11803) );
  NAND2_X1 U14719 ( .A1(n11755), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11810) );
  NAND2_X1 U14720 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11809) );
  NAND2_X1 U14721 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11808) );
  NAND2_X1 U14722 ( .A1(n11772), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11807) );
  NAND2_X1 U14723 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11814) );
  NAND2_X1 U14724 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11813) );
  NAND2_X1 U14725 ( .A1(n9648), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11812) );
  NAND2_X1 U14726 ( .A1(n11869), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11811) );
  NAND2_X1 U14727 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11818) );
  NAND2_X1 U14728 ( .A1(n11825), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11817) );
  NAND2_X1 U14729 ( .A1(n9651), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11816) );
  NAND2_X1 U14730 ( .A1(n11874), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11815) );
  NAND4_X4 U14731 ( .A1(n11822), .A2(n11821), .A3(n11820), .A4(n11819), .ZN(
        n11848) );
  NOR2_X1 U14732 ( .A1(n13169), .A2(n11848), .ZN(n11823) );
  AND2_X2 U14733 ( .A1(n11852), .A2(n11823), .ZN(n12743) );
  AOI22_X1 U14734 ( .A1(n11760), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U14735 ( .A1(n11887), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11828) );
  AOI22_X1 U14736 ( .A1(n11754), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n11825), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11827) );
  AOI22_X1 U14737 ( .A1(n9647), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11869), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11826) );
  NAND4_X1 U14738 ( .A1(n11829), .A2(n11828), .A3(n11827), .A4(n11826), .ZN(
        n11835) );
  AOI22_X1 U14739 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11833) );
  AOI22_X1 U14740 ( .A1(n12103), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9629), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11832) );
  AOI22_X1 U14741 ( .A1(n11755), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11772), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11831) );
  AOI22_X1 U14742 ( .A1(n9650), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11874), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11830) );
  NAND4_X1 U14743 ( .A1(n11833), .A2(n11832), .A3(n11831), .A4(n11830), .ZN(
        n11834) );
  NAND2_X1 U14744 ( .A1(n11932), .A2(n13743), .ZN(n11837) );
  NAND2_X1 U14745 ( .A1(n13747), .A2(n13360), .ZN(n13171) );
  AND2_X2 U14746 ( .A1(n12538), .A2(n11841), .ZN(n12929) );
  NAND2_X1 U14747 ( .A1(n11839), .A2(n11848), .ZN(n12553) );
  XNOR2_X1 U14748 ( .A(P1_STATE_REG_1__SCAN_IN), .B(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n12934) );
  NAND3_X1 U14749 ( .A1(n13740), .A2(n13402), .A3(n11839), .ZN(n13165) );
  NAND2_X1 U14750 ( .A1(n13352), .A2(n11848), .ZN(n11847) );
  NAND2_X1 U14751 ( .A1(n13748), .A2(n11847), .ZN(n13164) );
  NOR2_X1 U14752 ( .A1(n15791), .A2(n13743), .ZN(n11849) );
  NAND2_X1 U14753 ( .A1(n13169), .A2(n13352), .ZN(n11851) );
  NAND2_X1 U14754 ( .A1(n11852), .A2(n11851), .ZN(n11853) );
  NAND2_X1 U14755 ( .A1(n12939), .A2(n11854), .ZN(n11855) );
  NAND2_X1 U14756 ( .A1(n19909), .A2(n9755), .ZN(n12597) );
  MUX2_X1 U14757 ( .A(n12597), .B(n15798), .S(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .Z(n11856) );
  INV_X1 U14758 ( .A(n12939), .ZN(n11867) );
  NAND2_X1 U14759 ( .A1(n11854), .A2(n13734), .ZN(n11866) );
  NAND2_X1 U14760 ( .A1(n13402), .A2(n11932), .ZN(n13750) );
  AND4_X1 U14761 ( .A1(n13750), .A2(P1_STATE2_REG_0__SCAN_IN), .A3(n19909), 
        .A4(n13637), .ZN(n11862) );
  INV_X1 U14762 ( .A(n13740), .ZN(n14199) );
  AND2_X1 U14763 ( .A1(n14199), .A2(n9644), .ZN(n12794) );
  NAND2_X1 U14764 ( .A1(n11857), .A2(n13360), .ZN(n11860) );
  INV_X1 U14765 ( .A(n11858), .ZN(n11859) );
  AOI22_X1 U14766 ( .A1(n12794), .A2(n11860), .B1(n11859), .B2(n20762), .ZN(
        n11861) );
  AND3_X1 U14767 ( .A1(n11863), .A2(n11862), .A3(n11861), .ZN(n11865) );
  INV_X1 U14768 ( .A(n11918), .ZN(n11868) );
  AOI22_X1 U14769 ( .A1(n12505), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11873) );
  AOI22_X1 U14770 ( .A1(n12454), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12513), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11872) );
  AOI22_X1 U14771 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11871) );
  AOI22_X1 U14772 ( .A1(n9646), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11870) );
  NAND4_X1 U14773 ( .A1(n11873), .A2(n11872), .A3(n11871), .A4(n11870), .ZN(
        n11880) );
  AOI22_X1 U14774 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9629), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11878) );
  AOI22_X1 U14775 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11877) );
  AOI22_X1 U14776 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11876) );
  AOI22_X1 U14777 ( .A1(n12251), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11875) );
  NAND4_X1 U14778 ( .A1(n11878), .A2(n11877), .A3(n11876), .A4(n11875), .ZN(
        n11879) );
  NAND2_X1 U14779 ( .A1(n13743), .A2(n12672), .ZN(n11896) );
  NOR2_X1 U14780 ( .A1(n11896), .A2(n9755), .ZN(n11899) );
  NOR2_X1 U14781 ( .A1(n11988), .A2(n12672), .ZN(n11900) );
  AOI22_X1 U14782 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12512), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11886) );
  AOI22_X1 U14783 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12441), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n11885) );
  AOI22_X1 U14784 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11884) );
  AOI22_X1 U14785 ( .A1(n12251), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11883) );
  NAND4_X1 U14786 ( .A1(n11886), .A2(n11885), .A3(n11884), .A4(n11883), .ZN(
        n11893) );
  AOI22_X1 U14787 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12503), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n11891) );
  AOI22_X1 U14788 ( .A1(n12454), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9646), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11890) );
  AOI22_X1 U14789 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11889) );
  AOI22_X1 U14790 ( .A1(n9650), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11888) );
  NAND4_X1 U14791 ( .A1(n11891), .A2(n11890), .A3(n11889), .A4(n11888), .ZN(
        n11892) );
  MUX2_X1 U14792 ( .A(n11899), .B(n11900), .S(n12609), .Z(n11894) );
  INV_X1 U14793 ( .A(n11894), .ZN(n11895) );
  INV_X1 U14794 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11898) );
  AOI21_X1 U14795 ( .B1(n13638), .B2(n12609), .A(n9755), .ZN(n11897) );
  OAI211_X1 U14796 ( .C1(n12574), .C2(n11898), .A(n11897), .B(n11896), .ZN(
        n11930) );
  INV_X1 U14797 ( .A(n11899), .ZN(n12669) );
  INV_X1 U14798 ( .A(n11900), .ZN(n11913) );
  NAND2_X1 U14799 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11912) );
  INV_X1 U14800 ( .A(n11987), .ZN(n11962) );
  AOI22_X1 U14801 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11904) );
  AOI22_X1 U14802 ( .A1(n12454), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12441), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11903) );
  AOI22_X1 U14803 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11902) );
  AOI22_X1 U14804 ( .A1(n9646), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11901) );
  NAND4_X1 U14805 ( .A1(n11904), .A2(n11903), .A3(n11902), .A4(n11901), .ZN(
        n11910) );
  AOI22_X1 U14806 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12515), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11908) );
  AOI22_X1 U14807 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n11907) );
  AOI22_X1 U14808 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n9651), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11906) );
  AOI22_X1 U14809 ( .A1(n12251), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11905) );
  NAND4_X1 U14810 ( .A1(n11908), .A2(n11907), .A3(n11906), .A4(n11905), .ZN(
        n11909) );
  NAND2_X1 U14811 ( .A1(n11962), .A2(n12603), .ZN(n11911) );
  NAND2_X1 U14812 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n11940) );
  OAI21_X1 U14813 ( .B1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(n11940), .ZN(n20435) );
  INV_X1 U14814 ( .A(n15798), .ZN(n11942) );
  NAND2_X1 U14815 ( .A1(n11942), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11937) );
  INV_X1 U14816 ( .A(n11916), .ZN(n11917) );
  INV_X1 U14817 ( .A(n13209), .ZN(n11921) );
  NAND2_X1 U14818 ( .A1(n11921), .A2(n9755), .ZN(n11924) );
  INV_X1 U14819 ( .A(n11988), .ZN(n11922) );
  NAND2_X1 U14820 ( .A1(n11922), .A2(n12603), .ZN(n11923) );
  NAND2_X1 U14821 ( .A1(n13210), .A2(n12194), .ZN(n11929) );
  OR2_X1 U14822 ( .A1(n11843), .A2(n20760), .ZN(n12028) );
  NAND2_X1 U14823 ( .A1(n12533), .A2(P1_EAX_REG_1__SCAN_IN), .ZN(n11926) );
  NAND2_X1 U14824 ( .A1(n20760), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11925) );
  OAI211_X1 U14825 ( .C1(n12028), .C2(n14741), .A(n11926), .B(n11925), .ZN(
        n11927) );
  INV_X1 U14826 ( .A(n11927), .ZN(n11928) );
  NAND2_X1 U14827 ( .A1(n11929), .A2(n11928), .ZN(n13127) );
  XNOR2_X2 U14828 ( .A(n11931), .B(n11930), .ZN(n12612) );
  AOI21_X1 U14829 ( .B1(n12612), .B2(n11932), .A(n20760), .ZN(n13108) );
  NAND2_X1 U14830 ( .A1(n11934), .A2(n12194), .ZN(n11936) );
  AOI22_X1 U14831 ( .A1(n12533), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n20760), .ZN(n11935) );
  OAI211_X1 U14832 ( .C1(n12028), .C2(n14107), .A(n11936), .B(n11935), .ZN(
        n13107) );
  MUX2_X1 U14833 ( .A(n13634), .B(n13108), .S(n13107), .Z(n13126) );
  NAND2_X1 U14834 ( .A1(n13127), .A2(n13126), .ZN(n13124) );
  INV_X1 U14835 ( .A(n13124), .ZN(n11978) );
  AND2_X1 U14836 ( .A1(n11937), .A2(n14741), .ZN(n11938) );
  INV_X1 U14837 ( .A(n11940), .ZN(n15768) );
  NAND2_X1 U14838 ( .A1(n15768), .A2(n20502), .ZN(n20468) );
  NAND2_X1 U14839 ( .A1(n11940), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11941) );
  AND2_X1 U14840 ( .A1(n20468), .A2(n11941), .ZN(n13474) );
  NAND2_X1 U14841 ( .A1(n11942), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11943) );
  INV_X1 U14842 ( .A(n11945), .ZN(n11946) );
  AND2_X1 U14843 ( .A1(n11947), .A2(n11946), .ZN(n11948) );
  NAND2_X1 U14844 ( .A1(n11949), .A2(n11948), .ZN(n11950) );
  AOI22_X1 U14845 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12485), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11954) );
  AOI22_X1 U14846 ( .A1(n12454), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n12441), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11953) );
  INV_X1 U14847 ( .A(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n20930) );
  AOI22_X1 U14848 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11952) );
  AOI22_X1 U14849 ( .A1(n9646), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11951) );
  NAND4_X1 U14850 ( .A1(n11954), .A2(n11953), .A3(n11952), .A4(n11951), .ZN(
        n11960) );
  AOI22_X1 U14851 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12515), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11958) );
  AOI22_X1 U14852 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11957) );
  AOI22_X1 U14853 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11956) );
  AOI22_X1 U14854 ( .A1(n12251), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11955) );
  NAND4_X1 U14855 ( .A1(n11958), .A2(n11957), .A3(n11956), .A4(n11955), .ZN(
        n11959) );
  AOI22_X1 U14856 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n11962), .B2(n11961), .ZN(n11963) );
  INV_X1 U14857 ( .A(n11964), .ZN(n11965) );
  NOR2_X1 U14858 ( .A1(n11966), .A2(n11965), .ZN(n11967) );
  OR2_X1 U14859 ( .A1(n11970), .A2(n11969), .ZN(n11971) );
  NAND2_X1 U14860 ( .A1(n12533), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11973) );
  OAI21_X1 U14861 ( .B1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n12005), .ZN(n20129) );
  OAI21_X1 U14862 ( .B1(n20129), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20760), 
        .ZN(n11972) );
  OAI211_X1 U14863 ( .C1(n12028), .C2(n20903), .A(n11973), .B(n11972), .ZN(
        n11974) );
  INV_X1 U14864 ( .A(n11974), .ZN(n11975) );
  OAI21_X1 U14865 ( .B1(n13235), .B2(n12215), .A(n11975), .ZN(n11976) );
  NAND2_X1 U14866 ( .A1(n12532), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11979) );
  NAND2_X1 U14867 ( .A1(n11976), .A2(n11979), .ZN(n13125) );
  INV_X1 U14868 ( .A(n13125), .ZN(n11977) );
  NAND2_X1 U14869 ( .A1(n11978), .A2(n11977), .ZN(n11980) );
  NAND3_X1 U14870 ( .A1(n20501), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n13473) );
  INV_X1 U14871 ( .A(n13473), .ZN(n11982) );
  NAND2_X1 U14872 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n11982), .ZN(
        n13329) );
  NAND2_X1 U14873 ( .A1(n20501), .A2(n13329), .ZN(n11983) );
  NOR3_X1 U14874 ( .A1(n20501), .A2(n20502), .A3(n15765), .ZN(n20589) );
  NAND2_X1 U14875 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20589), .ZN(
        n13456) );
  NAND2_X1 U14876 ( .A1(n11983), .A2(n13456), .ZN(n20373) );
  OAI22_X1 U14877 ( .A1(n12597), .A2(n20373), .B1(n15798), .B2(n20501), .ZN(
        n11984) );
  INV_X1 U14878 ( .A(n11984), .ZN(n11985) );
  AOI22_X1 U14879 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11992) );
  AOI22_X1 U14880 ( .A1(n12454), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12513), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11991) );
  AOI22_X1 U14881 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11990) );
  AOI22_X1 U14882 ( .A1(n9646), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11989) );
  NAND4_X1 U14883 ( .A1(n11992), .A2(n11991), .A3(n11990), .A4(n11989), .ZN(
        n11998) );
  AOI22_X1 U14884 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9629), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11996) );
  AOI22_X1 U14885 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11995) );
  AOI22_X1 U14886 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9650), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11994) );
  AOI22_X1 U14887 ( .A1(n12251), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11993) );
  NAND4_X1 U14888 ( .A1(n11996), .A2(n11995), .A3(n11994), .A4(n11993), .ZN(
        n11997) );
  AOI22_X1 U14889 ( .A1(n12556), .A2(n12640), .B1(n12580), .B2(
        P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11999) );
  NAND2_X1 U14890 ( .A1(n12000), .A2(n13239), .ZN(n12002) );
  INV_X1 U14891 ( .A(n20171), .ZN(n12003) );
  NAND2_X1 U14892 ( .A1(n12003), .A2(n12194), .ZN(n12012) );
  NAND2_X1 U14893 ( .A1(n12533), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n12009) );
  INV_X1 U14894 ( .A(n12005), .ZN(n12004) );
  INV_X1 U14895 ( .A(n12030), .ZN(n12032) );
  INV_X1 U14896 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12006) );
  NAND2_X1 U14897 ( .A1(n12006), .A2(n12005), .ZN(n12007) );
  NAND2_X1 U14898 ( .A1(n12032), .A2(n12007), .ZN(n20119) );
  AOI22_X1 U14899 ( .A1(n20119), .A2(n12528), .B1(n12532), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12008) );
  OAI211_X1 U14900 ( .C1(n12028), .C2(n13198), .A(n12009), .B(n12008), .ZN(
        n12010) );
  INV_X1 U14901 ( .A(n12010), .ZN(n12011) );
  NAND2_X1 U14902 ( .A1(n12012), .A2(n12011), .ZN(n13160) );
  AOI22_X1 U14903 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12515), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12016) );
  AOI22_X1 U14904 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n12325), .B1(
        n12503), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12015) );
  AOI22_X1 U14905 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9651), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12014) );
  AOI22_X1 U14906 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12251), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12013) );
  NAND4_X1 U14907 ( .A1(n12016), .A2(n12015), .A3(n12014), .A4(n12013), .ZN(
        n12022) );
  AOI22_X1 U14908 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n12479), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12020) );
  AOI22_X1 U14909 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12484), .B1(
        n12454), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12019) );
  AOI22_X1 U14910 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12512), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12018) );
  AOI22_X1 U14911 ( .A1(n9646), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12017) );
  NAND4_X1 U14912 ( .A1(n12020), .A2(n12019), .A3(n12018), .A4(n12017), .ZN(
        n12021) );
  NAND2_X1 U14913 ( .A1(n12556), .A2(n12639), .ZN(n12024) );
  NAND2_X1 U14914 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12023) );
  INV_X1 U14916 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n12027) );
  NAND2_X1 U14917 ( .A1(n12533), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12026) );
  NAND2_X1 U14918 ( .A1(n20760), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12025) );
  OAI211_X1 U14919 ( .C1(n12028), .C2(n12027), .A(n12026), .B(n12025), .ZN(
        n12029) );
  NAND2_X1 U14920 ( .A1(n12029), .A2(n12500), .ZN(n12036) );
  INV_X1 U14921 ( .A(n12053), .ZN(n12034) );
  INV_X1 U14922 ( .A(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n12031) );
  NAND2_X1 U14923 ( .A1(n12032), .A2(n12031), .ZN(n12033) );
  NAND2_X1 U14924 ( .A1(n12034), .A2(n12033), .ZN(n20111) );
  NAND2_X1 U14925 ( .A1(n20111), .A2(n12528), .ZN(n12035) );
  NAND2_X1 U14926 ( .A1(n12036), .A2(n12035), .ZN(n12037) );
  INV_X1 U14927 ( .A(n13232), .ZN(n12038) );
  NAND3_X1 U14928 ( .A1(n13161), .A2(n13160), .A3(n12038), .ZN(n13231) );
  AOI22_X1 U14929 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12513), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12043) );
  AOI22_X1 U14930 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12042) );
  AOI22_X1 U14931 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12041) );
  AOI22_X1 U14932 ( .A1(n12251), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12040) );
  NAND4_X1 U14933 ( .A1(n12043), .A2(n12042), .A3(n12041), .A4(n12040), .ZN(
        n12049) );
  AOI22_X1 U14934 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12454), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12047) );
  AOI22_X1 U14935 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12046) );
  AOI22_X1 U14936 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12045) );
  AOI22_X1 U14937 ( .A1(n9646), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12044) );
  NAND4_X1 U14938 ( .A1(n12047), .A2(n12046), .A3(n12045), .A4(n12044), .ZN(
        n12048) );
  NAND2_X1 U14939 ( .A1(n12556), .A2(n12650), .ZN(n12051) );
  NAND2_X1 U14940 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n12050) );
  INV_X1 U14941 ( .A(n12057), .ZN(n12052) );
  XNOR2_X1 U14942 ( .A(n12058), .B(n12052), .ZN(n12638) );
  INV_X1 U14943 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n12055) );
  OAI21_X1 U14944 ( .B1(n12053), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n12071), .ZN(n19986) );
  AOI22_X1 U14945 ( .A1(n19986), .A2(n12528), .B1(n12532), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12054) );
  OAI21_X1 U14946 ( .B1(n12086), .B2(n12055), .A(n12054), .ZN(n12056) );
  AOI21_X1 U14947 ( .B1(n12638), .B2(n12194), .A(n12056), .ZN(n13371) );
  AOI22_X1 U14948 ( .A1(n12505), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12062) );
  AOI22_X1 U14949 ( .A1(n12454), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12513), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12061) );
  AOI22_X1 U14950 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12060) );
  AOI22_X1 U14951 ( .A1(n9646), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12059) );
  NAND4_X1 U14952 ( .A1(n12062), .A2(n12061), .A3(n12060), .A4(n12059), .ZN(
        n12068) );
  AOI22_X1 U14953 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12515), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12066) );
  AOI22_X1 U14954 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12065) );
  AOI22_X1 U14955 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n9650), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12064) );
  AOI22_X1 U14956 ( .A1(n12251), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12063) );
  NAND4_X1 U14957 ( .A1(n12066), .A2(n12065), .A3(n12064), .A4(n12063), .ZN(
        n12067) );
  NAND2_X1 U14958 ( .A1(n12556), .A2(n12660), .ZN(n12070) );
  NAND2_X1 U14959 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n12069) );
  NAND2_X1 U14960 ( .A1(n12070), .A2(n12069), .ZN(n12078) );
  NAND2_X1 U14961 ( .A1(n12071), .A2(n19976), .ZN(n12073) );
  INV_X1 U14962 ( .A(n12083), .ZN(n12072) );
  NAND2_X1 U14963 ( .A1(n12073), .A2(n12072), .ZN(n19971) );
  NAND2_X1 U14964 ( .A1(n19971), .A2(n12528), .ZN(n12074) );
  OAI21_X1 U14965 ( .B1(n19976), .B2(n12213), .A(n12074), .ZN(n12075) );
  AOI21_X1 U14966 ( .B1(n12527), .B2(P1_EAX_REG_6__SCAN_IN), .A(n12075), .ZN(
        n12076) );
  INV_X1 U14967 ( .A(n13373), .ZN(n12102) );
  NAND2_X1 U14968 ( .A1(n12556), .A2(n12672), .ZN(n12081) );
  NAND2_X1 U14969 ( .A1(n12580), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n12080) );
  NAND2_X1 U14970 ( .A1(n12081), .A2(n12080), .ZN(n12082) );
  INV_X1 U14971 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n12085) );
  OAI21_X1 U14972 ( .B1(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n12083), .A(
        n12114), .ZN(n19962) );
  AOI22_X1 U14973 ( .A1(n12528), .A2(n19962), .B1(n12532), .B2(
        P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12084) );
  OAI21_X1 U14974 ( .B1(n12086), .B2(n12085), .A(n12084), .ZN(n12087) );
  NAND2_X1 U14975 ( .A1(n12527), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12100) );
  AOI22_X1 U14976 ( .A1(n12505), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12306), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12091) );
  AOI22_X1 U14977 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12503), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12090) );
  AOI22_X1 U14978 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12251), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12089) );
  AOI22_X1 U14979 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12088) );
  NAND4_X1 U14980 ( .A1(n12091), .A2(n12090), .A3(n12089), .A4(n12088), .ZN(
        n12097) );
  AOI22_X1 U14981 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12513), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12095) );
  AOI22_X1 U14982 ( .A1(n12454), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9646), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12094) );
  AOI22_X1 U14983 ( .A1(n9652), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12093) );
  AOI22_X1 U14984 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12092) );
  NAND4_X1 U14985 ( .A1(n12095), .A2(n12094), .A3(n12093), .A4(n12092), .ZN(
        n12096) );
  OAI21_X1 U14986 ( .B1(n12097), .B2(n12096), .A(n12194), .ZN(n12099) );
  XOR2_X1 U14987 ( .A(n19953), .B(n12114), .Z(n19951) );
  INV_X1 U14988 ( .A(n19951), .ZN(n13769) );
  AOI22_X1 U14989 ( .A1(n12532), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n13634), .B2(n13769), .ZN(n12098) );
  NAND2_X1 U14990 ( .A1(n12102), .A2(n12101), .ZN(n13569) );
  BUF_X2 U14991 ( .A(n12103), .Z(n12305) );
  AOI22_X1 U14992 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12107) );
  AOI22_X1 U14993 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12106) );
  AOI22_X1 U14994 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12105) );
  AOI22_X1 U14995 ( .A1(n12251), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12104) );
  NAND4_X1 U14996 ( .A1(n12107), .A2(n12106), .A3(n12105), .A4(n12104), .ZN(
        n12113) );
  AOI22_X1 U14997 ( .A1(n12505), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12485), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12111) );
  AOI22_X1 U14998 ( .A1(n12454), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12110) );
  AOI22_X1 U14999 ( .A1(n9646), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12109) );
  AOI22_X1 U15000 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9650), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12108) );
  NAND4_X1 U15001 ( .A1(n12111), .A2(n12110), .A3(n12109), .A4(n12108), .ZN(
        n12112) );
  NOR2_X1 U15002 ( .A1(n12113), .A2(n12112), .ZN(n12117) );
  XNOR2_X1 U15003 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .B(n12121), .ZN(
        n19946) );
  OAI22_X1 U15004 ( .A1(n19946), .A2(n12500), .B1(n12213), .B2(n19940), .ZN(
        n12115) );
  INV_X1 U15005 ( .A(n12115), .ZN(n12116) );
  OAI21_X1 U15006 ( .B1(n12215), .B2(n12117), .A(n12116), .ZN(n12118) );
  INV_X1 U15007 ( .A(n12118), .ZN(n12120) );
  NAND2_X1 U15008 ( .A1(n12527), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12119) );
  XOR2_X1 U15009 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B(n12136), .Z(
        n15960) );
  AOI22_X1 U15010 ( .A1(n12505), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12513), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12125) );
  AOI22_X1 U15011 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12124) );
  AOI22_X1 U15012 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12251), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12123) );
  AOI22_X1 U15013 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12122) );
  NAND4_X1 U15014 ( .A1(n12125), .A2(n12124), .A3(n12123), .A4(n12122), .ZN(
        n12131) );
  AOI22_X1 U15015 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n12454), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12129) );
  AOI22_X1 U15016 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9629), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12128) );
  AOI22_X1 U15017 ( .A1(n9646), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12127) );
  AOI22_X1 U15018 ( .A1(n9651), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12126) );
  NAND4_X1 U15019 ( .A1(n12129), .A2(n12128), .A3(n12127), .A4(n12126), .ZN(
        n12130) );
  NOR2_X1 U15020 ( .A1(n12131), .A2(n12130), .ZN(n12133) );
  INV_X1 U15021 ( .A(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12132) );
  OAI22_X1 U15022 ( .A1(n12215), .A2(n12133), .B1(n12213), .B2(n12132), .ZN(
        n12134) );
  AOI21_X1 U15023 ( .B1(n12527), .B2(P1_EAX_REG_10__SCAN_IN), .A(n12134), .ZN(
        n12135) );
  OAI21_X1 U15024 ( .B1(n15960), .B2(n12500), .A(n12135), .ZN(n13662) );
  XNOR2_X1 U15025 ( .A(n12164), .B(n13783), .ZN(n14611) );
  NAND2_X1 U15026 ( .A1(n14611), .A2(n12528), .ZN(n12139) );
  NOR2_X1 U15027 ( .A1(n12213), .A2(n13783), .ZN(n12137) );
  AOI21_X1 U15028 ( .B1(n12527), .B2(P1_EAX_REG_11__SCAN_IN), .A(n12137), .ZN(
        n12138) );
  NAND2_X1 U15029 ( .A1(n12139), .A2(n12138), .ZN(n12151) );
  AOI22_X1 U15030 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12143) );
  AOI22_X1 U15031 ( .A1(n12505), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12142) );
  AOI22_X1 U15032 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9646), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12141) );
  AOI22_X1 U15033 ( .A1(n12454), .A2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12140) );
  NAND4_X1 U15034 ( .A1(n12143), .A2(n12142), .A3(n12141), .A4(n12140), .ZN(
        n12149) );
  AOI22_X1 U15035 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12512), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12147) );
  AOI22_X1 U15036 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12146) );
  AOI22_X1 U15037 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9650), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12145) );
  AOI22_X1 U15038 ( .A1(n12251), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12144) );
  NAND4_X1 U15039 ( .A1(n12147), .A2(n12146), .A3(n12145), .A4(n12144), .ZN(
        n12148) );
  NOR2_X1 U15040 ( .A1(n12149), .A2(n12148), .ZN(n12150) );
  NOR2_X1 U15041 ( .A1(n12215), .A2(n12150), .ZN(n13775) );
  NAND2_X1 U15042 ( .A1(n13773), .A2(n13775), .ZN(n13774) );
  INV_X1 U15043 ( .A(n12151), .ZN(n12152) );
  NAND2_X2 U15044 ( .A1(n13774), .A2(n12153), .ZN(n13795) );
  AOI22_X1 U15045 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12484), .B1(
        n12512), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12157) );
  AOI22_X1 U15046 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n12454), .B1(
        n9646), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12156) );
  AOI22_X1 U15047 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12251), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12155) );
  AOI22_X1 U15048 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12154) );
  NAND4_X1 U15049 ( .A1(n12157), .A2(n12156), .A3(n12155), .A4(n12154), .ZN(
        n12163) );
  AOI22_X1 U15050 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12161) );
  AOI22_X1 U15051 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12160) );
  AOI22_X1 U15052 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n12485), .B1(
        n9650), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12159) );
  AOI22_X1 U15053 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12158) );
  NAND4_X1 U15054 ( .A1(n12161), .A2(n12160), .A3(n12159), .A4(n12158), .ZN(
        n12162) );
  NOR2_X1 U15055 ( .A1(n12163), .A2(n12162), .ZN(n12167) );
  NAND2_X1 U15056 ( .A1(n12527), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n12166) );
  XNOR2_X1 U15057 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12168), .ZN(
        n15884) );
  AOI22_X1 U15058 ( .A1(n13634), .A2(n15884), .B1(n12532), .B2(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12165) );
  OAI211_X1 U15059 ( .C1(n12167), .C2(n12215), .A(n12166), .B(n12165), .ZN(
        n13794) );
  XOR2_X1 U15060 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B(n12219), .Z(
        n15934) );
  AOI22_X1 U15061 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12485), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12173) );
  AOI22_X1 U15062 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n12515), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12172) );
  AOI22_X1 U15063 ( .A1(n12454), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9646), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12171) );
  AOI22_X1 U15064 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12170) );
  NAND4_X1 U15065 ( .A1(n12173), .A2(n12172), .A3(n12171), .A4(n12170), .ZN(
        n12179) );
  AOI22_X1 U15066 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12177) );
  AOI22_X1 U15067 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12176) );
  AOI22_X1 U15068 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12175) );
  AOI22_X1 U15069 ( .A1(n12251), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12174) );
  NAND4_X1 U15070 ( .A1(n12177), .A2(n12176), .A3(n12175), .A4(n12174), .ZN(
        n12178) );
  NOR2_X1 U15071 ( .A1(n12179), .A2(n12178), .ZN(n12181) );
  INV_X1 U15072 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12180) );
  OAI22_X1 U15073 ( .A1(n12215), .A2(n12181), .B1(n12213), .B2(n12180), .ZN(
        n12182) );
  AOI21_X1 U15074 ( .B1(n12527), .B2(P1_EAX_REG_15__SCAN_IN), .A(n12182), .ZN(
        n12183) );
  OAI21_X1 U15075 ( .B1(n15934), .B2(n12500), .A(n12183), .ZN(n12184) );
  INV_X1 U15076 ( .A(n12184), .ZN(n14390) );
  XNOR2_X1 U15077 ( .A(n12185), .B(n12199), .ZN(n14603) );
  AOI22_X1 U15078 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12512), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12189) );
  AOI22_X1 U15079 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9629), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12188) );
  AOI22_X1 U15080 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12251), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12187) );
  AOI22_X1 U15081 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9650), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12186) );
  NAND4_X1 U15082 ( .A1(n12189), .A2(n12188), .A3(n12187), .A4(n12186), .ZN(
        n12196) );
  AOI22_X1 U15083 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12193) );
  AOI22_X1 U15084 ( .A1(n12454), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9646), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12192) );
  AOI22_X1 U15085 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12191) );
  AOI22_X1 U15086 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12190) );
  NAND4_X1 U15087 ( .A1(n12193), .A2(n12192), .A3(n12191), .A4(n12190), .ZN(
        n12195) );
  OAI21_X1 U15088 ( .B1(n12196), .B2(n12195), .A(n12194), .ZN(n12198) );
  NAND2_X1 U15089 ( .A1(n12527), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12197) );
  OAI211_X1 U15090 ( .C1(n12213), .C2(n12199), .A(n12198), .B(n12197), .ZN(
        n12200) );
  AOI21_X1 U15091 ( .B1(n14603), .B2(n12528), .A(n12200), .ZN(n13809) );
  XOR2_X1 U15092 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n12201), .Z(
        n15945) );
  AOI22_X1 U15093 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12205) );
  AOI22_X1 U15094 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12503), .B2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12204) );
  AOI22_X1 U15095 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12251), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12203) );
  AOI22_X1 U15096 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12202) );
  NAND4_X1 U15097 ( .A1(n12205), .A2(n12204), .A3(n12203), .A4(n12202), .ZN(
        n12211) );
  AOI22_X1 U15098 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12454), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12209) );
  AOI22_X1 U15099 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12208) );
  AOI22_X1 U15100 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9651), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12207) );
  AOI22_X1 U15101 ( .A1(n9646), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12206) );
  NAND4_X1 U15102 ( .A1(n12209), .A2(n12208), .A3(n12207), .A4(n12206), .ZN(
        n12210) );
  NOR2_X1 U15103 ( .A1(n12211), .A2(n12210), .ZN(n12214) );
  INV_X1 U15104 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12212) );
  OAI22_X1 U15105 ( .A1(n12215), .A2(n12214), .B1(n12213), .B2(n12212), .ZN(
        n12216) );
  AOI21_X1 U15106 ( .B1(n12527), .B2(P1_EAX_REG_13__SCAN_IN), .A(n12216), .ZN(
        n12217) );
  OAI21_X1 U15107 ( .B1(n15945), .B2(n12500), .A(n12217), .ZN(n12218) );
  INV_X1 U15108 ( .A(n12218), .ZN(n14397) );
  INV_X1 U15109 ( .A(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n12220) );
  XNOR2_X1 U15110 ( .A(n12237), .B(n12220), .ZN(n14589) );
  NAND2_X1 U15111 ( .A1(n14589), .A2(n12528), .ZN(n12236) );
  AOI22_X1 U15112 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12224) );
  AOI22_X1 U15113 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12251), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12223) );
  AOI22_X1 U15114 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12222) );
  AOI22_X1 U15115 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12221) );
  NAND4_X1 U15116 ( .A1(n12224), .A2(n12223), .A3(n12222), .A4(n12221), .ZN(
        n12232) );
  NAND2_X1 U15117 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12226) );
  NAND2_X1 U15118 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12225) );
  AND3_X1 U15119 ( .A1(n12226), .A2(n12225), .A3(n12500), .ZN(n12230) );
  AOI22_X1 U15120 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9646), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12229) );
  AOI22_X1 U15121 ( .A1(n12454), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U15122 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12227) );
  NAND4_X1 U15123 ( .A1(n12230), .A2(n12229), .A3(n12228), .A4(n12227), .ZN(
        n12231) );
  INV_X1 U15124 ( .A(n11854), .ZN(n14739) );
  NAND2_X1 U15125 ( .A1(n12497), .A2(n12500), .ZN(n12336) );
  OAI21_X1 U15126 ( .B1(n12232), .B2(n12231), .A(n12336), .ZN(n12234) );
  AOI22_X1 U15127 ( .A1(n12527), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n20760), .ZN(n12233) );
  NAND2_X1 U15128 ( .A1(n12234), .A2(n12233), .ZN(n12235) );
  NAND2_X1 U15129 ( .A1(n12236), .A2(n12235), .ZN(n13835) );
  XOR2_X1 U15130 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12250), .Z(
        n15925) );
  AOI22_X1 U15131 ( .A1(n12527), .A2(P1_EAX_REG_17__SCAN_IN), .B1(n12532), 
        .B2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n12249) );
  AOI22_X1 U15132 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12241) );
  AOI22_X1 U15133 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12240) );
  AOI22_X1 U15134 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12239) );
  AOI22_X1 U15135 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12238) );
  NAND4_X1 U15136 ( .A1(n12241), .A2(n12240), .A3(n12239), .A4(n12238), .ZN(
        n12247) );
  AOI22_X1 U15137 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12485), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12245) );
  AOI22_X1 U15138 ( .A1(n12454), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9646), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12244) );
  AOI22_X1 U15139 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n12251), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12243) );
  AOI22_X1 U15140 ( .A1(n9652), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12242) );
  NAND4_X1 U15141 ( .A1(n12245), .A2(n12244), .A3(n12243), .A4(n12242), .ZN(
        n12246) );
  OAI21_X1 U15142 ( .B1(n12247), .B2(n12246), .A(n12524), .ZN(n12248) );
  OAI211_X1 U15143 ( .C1(n15925), .C2(n12500), .A(n12249), .B(n12248), .ZN(
        n13866) );
  NAND2_X1 U15144 ( .A1(n13836), .A2(n13866), .ZN(n13865) );
  XNOR2_X1 U15145 ( .A(n12284), .B(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15855) );
  NAND2_X1 U15146 ( .A1(n15855), .A2(n12528), .ZN(n12268) );
  AOI22_X1 U15147 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12512), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12255) );
  AOI22_X1 U15148 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12254) );
  AOI22_X1 U15149 ( .A1(n12511), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n12251), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12253) );
  AOI22_X1 U15150 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12252) );
  NAND4_X1 U15151 ( .A1(n12255), .A2(n12254), .A3(n12253), .A4(n12252), .ZN(
        n12263) );
  NAND2_X1 U15152 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(
        n12257) );
  NAND2_X1 U15153 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(
        n12256) );
  AND3_X1 U15154 ( .A1(n12257), .A2(n12256), .A3(n12500), .ZN(n12261) );
  AOI22_X1 U15155 ( .A1(n9646), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12260) );
  AOI22_X1 U15156 ( .A1(n12454), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12259) );
  AOI22_X1 U15157 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12258) );
  NAND4_X1 U15158 ( .A1(n12261), .A2(n12260), .A3(n12259), .A4(n12258), .ZN(
        n12262) );
  OAI21_X1 U15159 ( .B1(n12263), .B2(n12262), .A(n12336), .ZN(n12266) );
  INV_X1 U15160 ( .A(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n14579) );
  NOR2_X1 U15161 ( .A1(n14579), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12264) );
  AOI21_X1 U15162 ( .B1(n12527), .B2(P1_EAX_REG_18__SCAN_IN), .A(n12264), .ZN(
        n12265) );
  NAND2_X1 U15163 ( .A1(n12266), .A2(n12265), .ZN(n12267) );
  NAND2_X1 U15164 ( .A1(n12268), .A2(n12267), .ZN(n14380) );
  AOI22_X1 U15165 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12273) );
  AOI22_X1 U15166 ( .A1(n12454), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9646), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12272) );
  AOI22_X1 U15167 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12251), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12271) );
  AOI22_X1 U15168 ( .A1(n12514), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12270) );
  NAND4_X1 U15169 ( .A1(n12273), .A2(n12272), .A3(n12271), .A4(n12270), .ZN(
        n12279) );
  AOI22_X1 U15170 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9629), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12277) );
  AOI22_X1 U15171 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12503), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12276) );
  AOI22_X1 U15172 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12275) );
  AOI22_X1 U15173 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9650), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12274) );
  NAND4_X1 U15174 ( .A1(n12277), .A2(n12276), .A3(n12275), .A4(n12274), .ZN(
        n12278) );
  NOR2_X1 U15175 ( .A1(n12279), .A2(n12278), .ZN(n12283) );
  NAND2_X1 U15176 ( .A1(n20760), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n12280) );
  NAND2_X1 U15177 ( .A1(n12500), .A2(n12280), .ZN(n12281) );
  AOI21_X1 U15178 ( .B1(n12527), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12281), .ZN(
        n12282) );
  OAI21_X1 U15179 ( .B1(n12497), .B2(n12283), .A(n12282), .ZN(n12287) );
  OAI21_X1 U15180 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n12285), .A(
        n12321), .ZN(n15918) );
  OR2_X1 U15181 ( .A1(n12500), .A2(n15918), .ZN(n12286) );
  NAND2_X1 U15182 ( .A1(n12287), .A2(n12286), .ZN(n14374) );
  AOI22_X1 U15183 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12484), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12291) );
  AOI22_X1 U15184 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n12479), .B1(
        n12251), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12290) );
  AOI22_X1 U15185 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12289) );
  AOI22_X1 U15186 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12288) );
  NAND4_X1 U15187 ( .A1(n12291), .A2(n12290), .A3(n12289), .A4(n12288), .ZN(
        n12299) );
  NAND2_X1 U15188 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n12293) );
  NAND2_X1 U15189 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n12292) );
  AND3_X1 U15190 ( .A1(n12293), .A2(n12292), .A3(n12500), .ZN(n12297) );
  AOI22_X1 U15191 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12511), .B1(
        n9646), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12296) );
  AOI22_X1 U15192 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n12454), .B1(
        n9650), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12295) );
  AOI22_X1 U15193 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12294) );
  NAND4_X1 U15194 ( .A1(n12297), .A2(n12296), .A3(n12295), .A4(n12294), .ZN(
        n12298) );
  OAI21_X1 U15195 ( .B1(n12299), .B2(n12298), .A(n12336), .ZN(n12301) );
  AOI22_X1 U15196 ( .A1(n12527), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20760), .ZN(n12300) );
  NAND2_X1 U15197 ( .A1(n12301), .A2(n12300), .ZN(n12303) );
  XNOR2_X1 U15198 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B(n12321), .ZN(
        n15836) );
  NAND2_X1 U15199 ( .A1(n13634), .A2(n15836), .ZN(n12302) );
  NAND2_X1 U15200 ( .A1(n12303), .A2(n12302), .ZN(n14367) );
  INV_X1 U15201 ( .A(n14367), .ZN(n12304) );
  AOI22_X1 U15202 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12310) );
  AOI22_X1 U15203 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12325), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12309) );
  AOI22_X1 U15204 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9651), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12308) );
  AOI22_X1 U15205 ( .A1(n12251), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12307) );
  NAND4_X1 U15206 ( .A1(n12310), .A2(n12309), .A3(n12308), .A4(n12307), .ZN(
        n12316) );
  AOI22_X1 U15207 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12454), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12314) );
  AOI22_X1 U15208 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12503), .B2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12313) );
  AOI22_X1 U15209 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12312) );
  AOI22_X1 U15210 ( .A1(n9646), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12311) );
  NAND4_X1 U15211 ( .A1(n12314), .A2(n12313), .A3(n12312), .A4(n12311), .ZN(
        n12315) );
  NOR2_X1 U15212 ( .A1(n12316), .A2(n12315), .ZN(n12320) );
  NAND2_X1 U15213 ( .A1(n20760), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12317) );
  NAND2_X1 U15214 ( .A1(n12500), .A2(n12317), .ZN(n12318) );
  AOI21_X1 U15215 ( .B1(n12527), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12318), .ZN(
        n12319) );
  OAI21_X1 U15216 ( .B1(n12497), .B2(n12320), .A(n12319), .ZN(n12324) );
  INV_X1 U15217 ( .A(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n15845) );
  OAI21_X1 U15218 ( .B1(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n12322), .A(
        n12368), .ZN(n15910) );
  OR2_X1 U15219 ( .A1(n12500), .A2(n15910), .ZN(n12323) );
  NAND2_X1 U15220 ( .A1(n14337), .A2(n14339), .ZN(n14322) );
  INV_X2 U15221 ( .A(n14322), .ZN(n12344) );
  AOI22_X1 U15222 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12513), .B2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n12329) );
  AOI22_X1 U15223 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n12454), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12328) );
  AOI22_X1 U15224 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12251), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12327) );
  AOI22_X1 U15225 ( .A1(n12325), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12326) );
  NAND4_X1 U15226 ( .A1(n12329), .A2(n12328), .A3(n12327), .A4(n12326), .ZN(
        n12338) );
  NAND2_X1 U15227 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(
        n12331) );
  NAND2_X1 U15228 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(
        n12330) );
  AND3_X1 U15229 ( .A1(n12331), .A2(n12330), .A3(n12500), .ZN(n12335) );
  AOI22_X1 U15230 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n9646), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12334) );
  AOI22_X1 U15231 ( .A1(n12504), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12333) );
  AOI22_X1 U15232 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9651), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12332) );
  NAND4_X1 U15233 ( .A1(n12335), .A2(n12334), .A3(n12333), .A4(n12332), .ZN(
        n12337) );
  OAI21_X1 U15234 ( .B1(n12338), .B2(n12337), .A(n12336), .ZN(n12340) );
  AOI22_X1 U15235 ( .A1(n12527), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n20760), .ZN(n12339) );
  NAND2_X1 U15236 ( .A1(n12340), .A2(n12339), .ZN(n12342) );
  XNOR2_X1 U15237 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B(n12368), .ZN(
        n14564) );
  NAND2_X1 U15238 ( .A1(n13634), .A2(n14564), .ZN(n12341) );
  NAND2_X1 U15239 ( .A1(n12342), .A2(n12341), .ZN(n14325) );
  AOI22_X1 U15240 ( .A1(n12454), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12441), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12348) );
  AOI22_X1 U15241 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12347) );
  AOI22_X1 U15242 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9652), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12346) );
  AOI22_X1 U15243 ( .A1(n9646), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12345) );
  NAND4_X1 U15244 ( .A1(n12348), .A2(n12347), .A3(n12346), .A4(n12345), .ZN(
        n12354) );
  AOI22_X1 U15245 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12485), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12352) );
  AOI22_X1 U15246 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12351) );
  AOI22_X1 U15247 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12251), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12350) );
  AOI22_X1 U15248 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12349) );
  NAND4_X1 U15249 ( .A1(n12352), .A2(n12351), .A3(n12350), .A4(n12349), .ZN(
        n12353) );
  NOR2_X1 U15250 ( .A1(n12354), .A2(n12353), .ZN(n12377) );
  AOI22_X1 U15251 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12454), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12358) );
  AOI22_X1 U15252 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12357) );
  AOI22_X1 U15253 ( .A1(n9646), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12356) );
  AOI22_X1 U15254 ( .A1(n9651), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12355) );
  NAND4_X1 U15255 ( .A1(n12358), .A2(n12357), .A3(n12356), .A4(n12355), .ZN(
        n12364) );
  AOI22_X1 U15256 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12441), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12362) );
  AOI22_X1 U15257 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12503), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12361) );
  AOI22_X1 U15258 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12251), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12360) );
  AOI22_X1 U15259 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12359) );
  NAND4_X1 U15260 ( .A1(n12362), .A2(n12361), .A3(n12360), .A4(n12359), .ZN(
        n12363) );
  NOR2_X1 U15261 ( .A1(n12364), .A2(n12363), .ZN(n12376) );
  XNOR2_X1 U15262 ( .A(n12377), .B(n12376), .ZN(n12367) );
  INV_X1 U15263 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n12371) );
  AOI21_X1 U15264 ( .B1(n12371), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12365) );
  AOI21_X1 U15265 ( .B1(n12527), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12365), .ZN(
        n12366) );
  OAI21_X1 U15266 ( .B1(n12497), .B2(n12367), .A(n12366), .ZN(n12375) );
  INV_X1 U15267 ( .A(n12370), .ZN(n12372) );
  NAND2_X1 U15268 ( .A1(n12372), .A2(n12371), .ZN(n12373) );
  AND2_X1 U15269 ( .A1(n12395), .A2(n12373), .ZN(n14559) );
  NAND2_X1 U15270 ( .A1(n14559), .A2(n12528), .ZN(n12374) );
  NAND2_X1 U15271 ( .A1(n12375), .A2(n12374), .ZN(n14308) );
  NOR2_X1 U15272 ( .A1(n12377), .A2(n12376), .ZN(n12410) );
  AOI22_X1 U15273 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n12485), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12381) );
  AOI22_X1 U15274 ( .A1(n12454), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12380) );
  AOI22_X1 U15275 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12379) );
  AOI22_X1 U15276 ( .A1(n9646), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12378) );
  NAND4_X1 U15277 ( .A1(n12381), .A2(n12380), .A3(n12379), .A4(n12378), .ZN(
        n12387) );
  AOI22_X1 U15278 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12385) );
  AOI22_X1 U15279 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12384) );
  AOI22_X1 U15280 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9651), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12383) );
  AOI22_X1 U15281 ( .A1(n12251), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12382) );
  NAND4_X1 U15282 ( .A1(n12385), .A2(n12384), .A3(n12383), .A4(n12382), .ZN(
        n12386) );
  OR2_X1 U15283 ( .A1(n12387), .A2(n12386), .ZN(n12409) );
  INV_X1 U15284 ( .A(n12409), .ZN(n12388) );
  XNOR2_X1 U15285 ( .A(n12410), .B(n12388), .ZN(n12389) );
  NAND2_X1 U15286 ( .A1(n12389), .A2(n12524), .ZN(n12393) );
  INV_X1 U15287 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12394) );
  AOI21_X1 U15288 ( .B1(n12394), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12390) );
  AOI21_X1 U15289 ( .B1(n12527), .B2(P1_EAX_REG_24__SCAN_IN), .A(n12390), .ZN(
        n12392) );
  XNOR2_X1 U15290 ( .A(n12395), .B(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14547) );
  AOI21_X1 U15291 ( .B1(n12393), .B2(n12392), .A(n12391), .ZN(n14299) );
  INV_X1 U15292 ( .A(n12396), .ZN(n12397) );
  INV_X1 U15293 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n14285) );
  NAND2_X1 U15294 ( .A1(n12397), .A2(n14285), .ZN(n12398) );
  NAND2_X1 U15295 ( .A1(n12432), .A2(n12398), .ZN(n14540) );
  AOI22_X1 U15296 ( .A1(n11882), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12512), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12402) );
  AOI22_X1 U15297 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12454), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12401) );
  AOI22_X1 U15298 ( .A1(n9646), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12400) );
  AOI22_X1 U15299 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n9651), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12399) );
  NAND4_X1 U15300 ( .A1(n12402), .A2(n12401), .A3(n12400), .A4(n12399), .ZN(
        n12408) );
  AOI22_X1 U15301 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n12406) );
  AOI22_X1 U15302 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n12251), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12405) );
  AOI22_X1 U15303 ( .A1(n12484), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12404) );
  AOI22_X1 U15304 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12403) );
  NAND4_X1 U15305 ( .A1(n12406), .A2(n12405), .A3(n12404), .A4(n12403), .ZN(
        n12407) );
  NOR2_X1 U15306 ( .A1(n12408), .A2(n12407), .ZN(n12427) );
  NAND2_X1 U15307 ( .A1(n12410), .A2(n12409), .ZN(n12426) );
  XNOR2_X1 U15308 ( .A(n12427), .B(n12426), .ZN(n12413) );
  AOI21_X1 U15309 ( .B1(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n20760), .A(
        n12528), .ZN(n12412) );
  NAND2_X1 U15310 ( .A1(n12527), .A2(P1_EAX_REG_25__SCAN_IN), .ZN(n12411) );
  OAI211_X1 U15311 ( .C1(n12413), .C2(n12497), .A(n12412), .B(n12411), .ZN(
        n12414) );
  AOI22_X1 U15312 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12485), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12418) );
  AOI22_X1 U15313 ( .A1(n12454), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12417) );
  AOI22_X1 U15314 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12416) );
  AOI22_X1 U15315 ( .A1(n9646), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12415) );
  NAND4_X1 U15316 ( .A1(n12418), .A2(n12417), .A3(n12416), .A4(n12415), .ZN(
        n12425) );
  AOI22_X1 U15317 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9628), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12423) );
  AOI22_X1 U15318 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12422) );
  AOI22_X1 U15319 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9651), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12421) );
  AOI22_X1 U15320 ( .A1(n12251), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12420) );
  NAND4_X1 U15321 ( .A1(n12423), .A2(n12422), .A3(n12421), .A4(n12420), .ZN(
        n12424) );
  OR2_X1 U15322 ( .A1(n12425), .A2(n12424), .ZN(n12448) );
  NOR2_X1 U15323 ( .A1(n12427), .A2(n12426), .ZN(n12449) );
  XOR2_X1 U15324 ( .A(n12448), .B(n12449), .Z(n12428) );
  NAND2_X1 U15325 ( .A1(n12428), .A2(n12524), .ZN(n12431) );
  INV_X1 U15326 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n14271) );
  NOR2_X1 U15327 ( .A1(n14271), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12429) );
  AOI211_X1 U15328 ( .C1(n12527), .C2(P1_EAX_REG_26__SCAN_IN), .A(n12528), .B(
        n12429), .ZN(n12430) );
  XNOR2_X1 U15329 ( .A(n12432), .B(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14270) );
  AOI22_X1 U15330 ( .A1(n12431), .A2(n12430), .B1(n13634), .B2(n14270), .ZN(
        n14269) );
  NAND2_X1 U15331 ( .A1(n14268), .A2(n14269), .ZN(n14254) );
  INV_X1 U15332 ( .A(n12432), .ZN(n12433) );
  INV_X1 U15333 ( .A(n12434), .ZN(n12435) );
  INV_X1 U15334 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n14258) );
  NAND2_X1 U15335 ( .A1(n12435), .A2(n14258), .ZN(n12436) );
  NAND2_X1 U15336 ( .A1(n12473), .A2(n12436), .ZN(n14520) );
  AOI22_X1 U15337 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12440) );
  AOI22_X1 U15338 ( .A1(n12454), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n9646), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12439) );
  AOI22_X1 U15339 ( .A1(n9652), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12438) );
  AOI22_X1 U15340 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12437) );
  NAND4_X1 U15341 ( .A1(n12440), .A2(n12439), .A3(n12438), .A4(n12437), .ZN(
        n12447) );
  AOI22_X1 U15342 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n12485), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12445) );
  AOI22_X1 U15343 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12441), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12444) );
  AOI22_X1 U15344 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12251), .B2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12443) );
  AOI22_X1 U15345 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12442) );
  NAND4_X1 U15346 ( .A1(n12445), .A2(n12444), .A3(n12443), .A4(n12442), .ZN(
        n12446) );
  NOR2_X1 U15347 ( .A1(n12447), .A2(n12446), .ZN(n12467) );
  NAND2_X1 U15348 ( .A1(n12449), .A2(n12448), .ZN(n12466) );
  XNOR2_X1 U15349 ( .A(n12467), .B(n12466), .ZN(n12452) );
  AOI21_X1 U15350 ( .B1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(n20760), .A(
        n13634), .ZN(n12451) );
  NAND2_X1 U15351 ( .A1(n12527), .A2(P1_EAX_REG_27__SCAN_IN), .ZN(n12450) );
  OAI211_X1 U15352 ( .C1(n12452), .C2(n12497), .A(n12451), .B(n12450), .ZN(
        n12453) );
  NOR2_X2 U15353 ( .A1(n14254), .A2(n14255), .ZN(n14241) );
  AOI22_X1 U15354 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12458) );
  AOI22_X1 U15355 ( .A1(n12454), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12457) );
  AOI22_X1 U15356 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12456) );
  AOI22_X1 U15357 ( .A1(n9646), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12455) );
  NAND4_X1 U15358 ( .A1(n12458), .A2(n12457), .A3(n12456), .A4(n12455), .ZN(
        n12465) );
  AOI22_X1 U15359 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12515), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12463) );
  AOI22_X1 U15360 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12462) );
  AOI22_X1 U15361 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9650), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12461) );
  AOI22_X1 U15362 ( .A1(n12251), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12460) );
  NAND4_X1 U15363 ( .A1(n12463), .A2(n12462), .A3(n12461), .A4(n12460), .ZN(
        n12464) );
  OR2_X1 U15364 ( .A1(n12465), .A2(n12464), .ZN(n12493) );
  NOR2_X1 U15365 ( .A1(n12467), .A2(n12466), .ZN(n12494) );
  XOR2_X1 U15366 ( .A(n12493), .B(n12494), .Z(n12468) );
  NAND2_X1 U15367 ( .A1(n12468), .A2(n12524), .ZN(n12472) );
  INV_X1 U15368 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n12469) );
  NOR2_X1 U15369 ( .A1(n12469), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12470) );
  AOI211_X1 U15370 ( .C1(n12527), .C2(P1_EAX_REG_28__SCAN_IN), .A(n12528), .B(
        n12470), .ZN(n12471) );
  XNOR2_X1 U15371 ( .A(n12473), .B(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14505) );
  AOI22_X1 U15372 ( .A1(n12472), .A2(n12471), .B1(n13634), .B2(n14505), .ZN(
        n14243) );
  INV_X1 U15373 ( .A(n12473), .ZN(n12474) );
  INV_X1 U15374 ( .A(n12475), .ZN(n12477) );
  INV_X1 U15375 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n12476) );
  NAND2_X1 U15376 ( .A1(n12477), .A2(n12476), .ZN(n12478) );
  NAND2_X1 U15377 ( .A1(n12594), .A2(n12478), .ZN(n14491) );
  AOI22_X1 U15378 ( .A1(n12479), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12454), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12483) );
  AOI22_X1 U15379 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12482) );
  AOI22_X1 U15380 ( .A1(n9646), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12481) );
  AOI22_X1 U15381 ( .A1(n9652), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12480) );
  NAND4_X1 U15382 ( .A1(n12483), .A2(n12482), .A3(n12481), .A4(n12480), .ZN(
        n12492) );
  AOI22_X1 U15383 ( .A1(n12485), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12484), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12490) );
  AOI22_X1 U15384 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12503), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12489) );
  AOI22_X1 U15385 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12251), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12488) );
  AOI22_X1 U15386 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12487) );
  NAND4_X1 U15387 ( .A1(n12490), .A2(n12489), .A3(n12488), .A4(n12487), .ZN(
        n12491) );
  NOR2_X1 U15388 ( .A1(n12492), .A2(n12491), .ZN(n12502) );
  NAND2_X1 U15389 ( .A1(n12494), .A2(n12493), .ZN(n12501) );
  XNOR2_X1 U15390 ( .A(n12502), .B(n12501), .ZN(n12498) );
  AOI21_X1 U15391 ( .B1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n20760), .A(
        n13634), .ZN(n12496) );
  NAND2_X1 U15392 ( .A1(n12527), .A2(P1_EAX_REG_29__SCAN_IN), .ZN(n12495) );
  OAI211_X1 U15393 ( .C1(n12498), .C2(n12497), .A(n12496), .B(n12495), .ZN(
        n12499) );
  OAI21_X1 U15394 ( .B1(n12500), .B2(n14491), .A(n12499), .ZN(n14232) );
  NOR2_X1 U15395 ( .A1(n12502), .A2(n12501), .ZN(n12523) );
  AOI22_X1 U15396 ( .A1(n12454), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9646), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12510) );
  AOI22_X1 U15397 ( .A1(n12503), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12251), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12509) );
  AOI22_X1 U15398 ( .A1(n12505), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12504), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12508) );
  AOI22_X1 U15399 ( .A1(n9650), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12506), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12507) );
  NAND4_X1 U15400 ( .A1(n12510), .A2(n12509), .A3(n12508), .A4(n12507), .ZN(
        n12521) );
  AOI22_X1 U15401 ( .A1(n12512), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n12511), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12519) );
  AOI22_X1 U15402 ( .A1(n12486), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12513), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12518) );
  AOI22_X1 U15403 ( .A1(n12305), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n12517) );
  AOI22_X1 U15404 ( .A1(n12515), .A2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n12514), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12516) );
  NAND4_X1 U15405 ( .A1(n12519), .A2(n12518), .A3(n12517), .A4(n12516), .ZN(
        n12520) );
  NOR2_X1 U15406 ( .A1(n12521), .A2(n12520), .ZN(n12522) );
  XNOR2_X1 U15407 ( .A(n12523), .B(n12522), .ZN(n12525) );
  NAND2_X1 U15408 ( .A1(n12525), .A2(n12524), .ZN(n12531) );
  INV_X1 U15409 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14483) );
  AOI21_X1 U15410 ( .B1(n14483), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12526) );
  AOI21_X1 U15411 ( .B1(n12527), .B2(P1_EAX_REG_30__SCAN_IN), .A(n12526), .ZN(
        n12530) );
  XNOR2_X1 U15412 ( .A(n12594), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14481) );
  AND2_X1 U15413 ( .A1(n14481), .A2(n12528), .ZN(n12529) );
  AOI21_X1 U15414 ( .B1(n12531), .B2(n12530), .A(n12529), .ZN(n14215) );
  NAND2_X1 U15415 ( .A1(n14231), .A2(n14215), .ZN(n12536) );
  AOI22_X1 U15416 ( .A1(n12533), .A2(P1_EAX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n12532), .ZN(n12534) );
  INV_X1 U15417 ( .A(n12534), .ZN(n12535) );
  XNOR2_X2 U15418 ( .A(n12536), .B(n12535), .ZN(n14202) );
  NAND3_X1 U15419 ( .A1(n9755), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16108) );
  INV_X1 U15420 ( .A(n16108), .ZN(n12537) );
  NOR2_X2 U15421 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20585) );
  NAND2_X1 U15422 ( .A1(n12537), .A2(n20585), .ZN(n14616) );
  INV_X2 U15423 ( .A(n14616), .ZN(n20125) );
  AOI21_X1 U15424 ( .B1(n11854), .B2(n13638), .A(n13171), .ZN(n12539) );
  NAND2_X1 U15425 ( .A1(n12539), .A2(n12538), .ZN(n12930) );
  NOR2_X1 U15426 ( .A1(n12930), .A2(n13169), .ZN(n12590) );
  MUX2_X1 U15427 ( .A(n15765), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n12550) );
  NAND2_X1 U15428 ( .A1(n20553), .A2(n15761), .ZN(n12554) );
  NAND2_X1 U15429 ( .A1(n12550), .A2(n12549), .ZN(n12541) );
  NAND2_X1 U15430 ( .A1(n15765), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12540) );
  NAND2_X1 U15431 ( .A1(n12541), .A2(n12540), .ZN(n12565) );
  MUX2_X1 U15432 ( .A(n20502), .B(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n12564) );
  NAND2_X1 U15433 ( .A1(n12565), .A2(n12564), .ZN(n12543) );
  NAND2_X1 U15434 ( .A1(n20502), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n12542) );
  XNOR2_X1 U15435 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n12547) );
  NOR2_X1 U15436 ( .A1(n13198), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12544) );
  INV_X1 U15437 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n12545) );
  NAND2_X1 U15438 ( .A1(n12545), .A2(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n12546) );
  NOR2_X1 U15439 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n12545), .ZN(
        n12577) );
  AOI21_X1 U15440 ( .B1(n12578), .B2(n12546), .A(n12577), .ZN(n12750) );
  NAND2_X1 U15441 ( .A1(n12576), .A2(n12750), .ZN(n12589) );
  NAND2_X1 U15442 ( .A1(n12750), .A2(n12556), .ZN(n12587) );
  XNOR2_X1 U15443 ( .A(n12548), .B(n12547), .ZN(n12747) );
  XNOR2_X1 U15444 ( .A(n12550), .B(n12549), .ZN(n12745) );
  NOR2_X1 U15445 ( .A1(n13344), .A2(n9755), .ZN(n12551) );
  INV_X1 U15446 ( .A(n12563), .ZN(n12552) );
  NOR2_X1 U15447 ( .A1(n12745), .A2(n12552), .ZN(n12561) );
  NAND2_X1 U15448 ( .A1(n12553), .A2(n13639), .ZN(n12570) );
  OAI21_X1 U15449 ( .B1(n15761), .B2(n20553), .A(n12554), .ZN(n12558) );
  INV_X1 U15450 ( .A(n12558), .ZN(n12555) );
  OAI211_X1 U15451 ( .C1(n13638), .C2(n13169), .A(n12570), .B(n12555), .ZN(
        n12560) );
  INV_X1 U15452 ( .A(n12576), .ZN(n12557) );
  OAI21_X1 U15453 ( .B1(n12571), .B2(n12558), .A(n12557), .ZN(n12559) );
  NAND2_X1 U15454 ( .A1(n12560), .A2(n12559), .ZN(n12562) );
  NAND2_X1 U15455 ( .A1(n12561), .A2(n12562), .ZN(n12569) );
  NAND2_X1 U15456 ( .A1(n12563), .A2(n13734), .ZN(n12582) );
  OAI211_X1 U15457 ( .C1(n12563), .C2(n12562), .A(n12745), .B(n12582), .ZN(
        n12568) );
  XNOR2_X1 U15458 ( .A(n12565), .B(n12564), .ZN(n12746) );
  NAND2_X1 U15459 ( .A1(n12580), .A2(n12746), .ZN(n12566) );
  OAI211_X1 U15460 ( .C1(n12571), .C2(n12746), .A(n12566), .B(n12570), .ZN(
        n12567) );
  NAND3_X1 U15461 ( .A1(n12569), .A2(n12568), .A3(n12567), .ZN(n12573) );
  AOI22_X1 U15462 ( .A1(n12574), .A2(n12747), .B1(n12573), .B2(n12572), .ZN(
        n12575) );
  AOI21_X1 U15463 ( .B1(n12576), .B2(n12747), .A(n12575), .ZN(n12584) );
  INV_X1 U15464 ( .A(n12748), .ZN(n12579) );
  NOR2_X1 U15465 ( .A1(n12580), .A2(n12579), .ZN(n12583) );
  NAND2_X1 U15466 ( .A1(n12580), .A2(n12748), .ZN(n12581) );
  OAI22_X1 U15467 ( .A1(n12584), .A2(n12583), .B1(n12582), .B2(n12581), .ZN(
        n12585) );
  AOI21_X1 U15468 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n9755), .A(
        n12585), .ZN(n12586) );
  NAND2_X1 U15469 ( .A1(n12587), .A2(n12586), .ZN(n12588) );
  NAND2_X1 U15470 ( .A1(n12590), .A2(n13730), .ZN(n15778) );
  NAND2_X1 U15471 ( .A1(n15798), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n19911) );
  INV_X1 U15472 ( .A(n20585), .ZN(n20556) );
  NAND2_X1 U15473 ( .A1(n20556), .A2(n12597), .ZN(n20766) );
  NAND2_X1 U15474 ( .A1(n20766), .A2(n9755), .ZN(n12591) );
  NAND2_X1 U15475 ( .A1(n9755), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12593) );
  INV_X1 U15476 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20761) );
  NAND2_X1 U15477 ( .A1(n20761), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n12592) );
  AND2_X1 U15478 ( .A1(n12593), .A2(n12592), .ZN(n13115) );
  INV_X1 U15479 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12595) );
  XNOR2_X1 U15480 ( .A(n12596), .B(n12595), .ZN(n13654) );
  INV_X1 U15481 ( .A(P1_REIP_REG_31__SCAN_IN), .ZN(n20735) );
  NOR2_X1 U15482 ( .A1(n20135), .A2(n20735), .ZN(n14129) );
  AOI21_X1 U15483 ( .B1(n20120), .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14129), .ZN(n12598) );
  OAI21_X1 U15484 ( .B1(n20130), .B2(n13654), .A(n12598), .ZN(n12599) );
  AOI21_X1 U15485 ( .B1(n14202), .B2(n20125), .A(n12599), .ZN(n12698) );
  NOR2_X1 U15486 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12601) );
  INV_X1 U15487 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12600) );
  NAND2_X1 U15488 ( .A1(n12602), .A2(n13734), .ZN(n12608) );
  NAND2_X1 U15489 ( .A1(n12609), .A2(n12603), .ZN(n12624) );
  OAI21_X1 U15490 ( .B1(n12603), .B2(n12609), .A(n12624), .ZN(n12605) );
  OAI21_X1 U15491 ( .B1(n12605), .B2(n15791), .A(n12604), .ZN(n12606) );
  INV_X1 U15492 ( .A(n12606), .ZN(n12607) );
  NAND2_X1 U15493 ( .A1(n12608), .A2(n12607), .ZN(n12613) );
  NAND2_X1 U15494 ( .A1(n13638), .A2(n13360), .ZN(n12616) );
  OAI21_X1 U15495 ( .B1(n15791), .B2(n12609), .A(n12616), .ZN(n12610) );
  INV_X1 U15496 ( .A(n12610), .ZN(n12611) );
  XNOR2_X1 U15497 ( .A(n12613), .B(n13110), .ZN(n13461) );
  NAND2_X1 U15498 ( .A1(n13461), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13462) );
  INV_X1 U15499 ( .A(n12613), .ZN(n12614) );
  OR2_X1 U15500 ( .A1(n13110), .A2(n12614), .ZN(n12615) );
  INV_X1 U15501 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20152) );
  OR2_X1 U15502 ( .A1(n13235), .A2(n12937), .ZN(n12620) );
  XNOR2_X1 U15503 ( .A(n12624), .B(n12623), .ZN(n12618) );
  INV_X1 U15504 ( .A(n12616), .ZN(n12617) );
  AOI21_X1 U15505 ( .B1(n12618), .B2(n20762), .A(n12617), .ZN(n12619) );
  NAND2_X1 U15506 ( .A1(n12620), .A2(n12619), .ZN(n20122) );
  NAND2_X1 U15507 ( .A1(n12621), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12622) );
  INV_X1 U15508 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20150) );
  OR2_X1 U15509 ( .A1(n20171), .A2(n12937), .ZN(n12628) );
  NAND2_X1 U15510 ( .A1(n12624), .A2(n12623), .ZN(n12642) );
  INV_X1 U15511 ( .A(n12640), .ZN(n12625) );
  XNOR2_X1 U15512 ( .A(n12642), .B(n12625), .ZN(n12626) );
  NAND2_X1 U15513 ( .A1(n12626), .A2(n20762), .ZN(n12627) );
  NAND2_X1 U15514 ( .A1(n12628), .A2(n12627), .ZN(n20113) );
  NAND2_X1 U15515 ( .A1(n12629), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n12630) );
  NAND2_X1 U15516 ( .A1(n12631), .A2(n12648), .ZN(n12635) );
  NAND2_X1 U15517 ( .A1(n12642), .A2(n12640), .ZN(n12632) );
  XNOR2_X1 U15518 ( .A(n12632), .B(n12639), .ZN(n12633) );
  NAND2_X1 U15519 ( .A1(n12633), .A2(n20762), .ZN(n12634) );
  NAND2_X1 U15520 ( .A1(n12635), .A2(n12634), .ZN(n12636) );
  INV_X1 U15521 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n20144) );
  XNOR2_X1 U15522 ( .A(n12636), .B(n20144), .ZN(n20105) );
  NAND2_X1 U15523 ( .A1(n12636), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12637) );
  NAND2_X1 U15524 ( .A1(n12638), .A2(n12648), .ZN(n12646) );
  AND2_X1 U15525 ( .A1(n12640), .A2(n12639), .ZN(n12641) );
  AND2_X1 U15526 ( .A1(n12642), .A2(n12641), .ZN(n12651) );
  INV_X1 U15527 ( .A(n12650), .ZN(n12643) );
  XNOR2_X1 U15528 ( .A(n12651), .B(n12643), .ZN(n12644) );
  NAND2_X1 U15529 ( .A1(n12644), .A2(n20762), .ZN(n12645) );
  INV_X1 U15530 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n16105) );
  NAND3_X1 U15531 ( .A1(n12647), .A2(n12649), .A3(n12648), .ZN(n12654) );
  NAND2_X1 U15532 ( .A1(n12651), .A2(n12650), .ZN(n12661) );
  XNOR2_X1 U15533 ( .A(n12660), .B(n12661), .ZN(n12652) );
  NAND2_X1 U15534 ( .A1(n20762), .A2(n12652), .ZN(n12653) );
  NAND2_X1 U15535 ( .A1(n12654), .A2(n12653), .ZN(n15971) );
  OR2_X1 U15536 ( .A1(n15971), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12655) );
  NAND2_X1 U15537 ( .A1(n15971), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12656) );
  NAND2_X1 U15538 ( .A1(n12657), .A2(n12656), .ZN(n15968) );
  INV_X1 U15539 ( .A(n12658), .ZN(n12659) );
  OR2_X1 U15540 ( .A1(n12659), .A2(n12937), .ZN(n12666) );
  INV_X1 U15541 ( .A(n12660), .ZN(n12662) );
  NOR2_X1 U15542 ( .A1(n12662), .A2(n12661), .ZN(n12671) );
  INV_X1 U15543 ( .A(n12671), .ZN(n12663) );
  XNOR2_X1 U15544 ( .A(n12672), .B(n12663), .ZN(n12664) );
  NAND2_X1 U15545 ( .A1(n20762), .A2(n12664), .ZN(n12665) );
  NAND2_X1 U15546 ( .A1(n12666), .A2(n12665), .ZN(n12667) );
  OR2_X1 U15547 ( .A1(n12667), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15966) );
  NAND2_X1 U15548 ( .A1(n15968), .A2(n15966), .ZN(n12668) );
  NAND2_X1 U15549 ( .A1(n12667), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15965) );
  NOR2_X1 U15550 ( .A1(n12669), .A2(n12937), .ZN(n12670) );
  NAND2_X1 U15551 ( .A1(n12672), .A2(n12671), .ZN(n12673) );
  NOR2_X1 U15552 ( .A1(n15791), .A2(n12673), .ZN(n12674) );
  NAND2_X1 U15553 ( .A1(n13725), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12676) );
  NAND2_X1 U15554 ( .A1(n15808), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12679) );
  NAND2_X1 U15555 ( .A1(n14598), .A2(n12679), .ZN(n12683) );
  NOR2_X1 U15556 ( .A1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15938) );
  INV_X1 U15557 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12680) );
  NAND2_X1 U15558 ( .A1(n15938), .A2(n12680), .ZN(n12681) );
  AND2_X1 U15559 ( .A1(n15808), .A2(n12681), .ZN(n14595) );
  INV_X1 U15560 ( .A(n15956), .ZN(n12687) );
  NOR2_X1 U15561 ( .A1(n15808), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15942) );
  AOI21_X1 U15562 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A(n15808), .ZN(n15939) );
  OR2_X1 U15563 ( .A1(n15808), .A2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12682) );
  NAND2_X1 U15564 ( .A1(n14597), .A2(n12682), .ZN(n14584) );
  AND2_X1 U15565 ( .A1(n15808), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14585) );
  NOR2_X1 U15566 ( .A1(n12683), .A2(n14585), .ZN(n15920) );
  NAND2_X1 U15567 ( .A1(n14584), .A2(n15920), .ZN(n12685) );
  XNOR2_X1 U15568 ( .A(n15808), .B(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n14587) );
  NOR2_X1 U15569 ( .A1(n14587), .A2(n15929), .ZN(n12684) );
  NAND2_X1 U15570 ( .A1(n12685), .A2(n12684), .ZN(n15919) );
  INV_X1 U15571 ( .A(n15919), .ZN(n12686) );
  INV_X1 U15572 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n14134) );
  XNOR2_X1 U15573 ( .A(n15808), .B(n14134), .ZN(n14577) );
  AND2_X1 U15574 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14693) );
  NAND2_X1 U15575 ( .A1(n14693), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n12688) );
  INV_X1 U15576 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12690) );
  INV_X1 U15577 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15810) );
  INV_X1 U15578 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15912) );
  NAND4_X1 U15579 ( .A1(n12690), .A2(n14134), .A3(n15810), .A4(n15912), .ZN(
        n12691) );
  OAI21_X2 U15580 ( .B1(n12689), .B2(n12691), .A(n15808), .ZN(n14561) );
  NOR2_X1 U15581 ( .A1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14496) );
  NAND2_X1 U15582 ( .A1(n14536), .A2(n14496), .ZN(n12692) );
  AND2_X1 U15583 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14119) );
  NAND2_X1 U15584 ( .A1(n14119), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14653) );
  INV_X1 U15585 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14497) );
  INV_X1 U15586 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14517) );
  INV_X1 U15587 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14502) );
  NAND2_X1 U15588 ( .A1(n14517), .A2(n14502), .ZN(n14635) );
  INV_X1 U15589 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14630) );
  NAND2_X1 U15590 ( .A1(n14478), .A2(n12693), .ZN(n12696) );
  NAND2_X1 U15591 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14636) );
  INV_X1 U15592 ( .A(n19918), .ZN(n12697) );
  NOR2_X1 U15593 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_0__SCAN_IN), 
        .ZN(n12700) );
  NOR4_X1 U15594 ( .A1(P2_BE_N_REG_1__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n12699) );
  NAND4_X1 U15595 ( .A1(n12700), .A2(P2_M_IO_N_REG_SCAN_IN), .A3(
        P2_W_R_N_REG_SCAN_IN), .A4(n12699), .ZN(n12713) );
  NOR2_X1 U15596 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n12713), .ZN(n16497)
         );
  NOR4_X1 U15597 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(
        P1_ADDRESS_REG_14__SCAN_IN), .A3(P1_ADDRESS_REG_13__SCAN_IN), .A4(
        P1_ADDRESS_REG_12__SCAN_IN), .ZN(n12704) );
  NOR4_X1 U15598 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_17__SCAN_IN), .A4(
        P1_ADDRESS_REG_16__SCAN_IN), .ZN(n12703) );
  NOR4_X1 U15599 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n12702) );
  NOR4_X1 U15600 ( .A1(P1_ADDRESS_REG_11__SCAN_IN), .A2(
        P1_ADDRESS_REG_10__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n12701) );
  AND4_X1 U15601 ( .A1(n12704), .A2(n12703), .A3(n12702), .A4(n12701), .ZN(
        n12709) );
  NOR4_X1 U15602 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_9__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n12707) );
  NOR4_X1 U15603 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n12706) );
  NOR4_X1 U15604 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n12705) );
  INV_X1 U15605 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20692) );
  AND4_X1 U15606 ( .A1(n12707), .A2(n12706), .A3(n12705), .A4(n20692), .ZN(
        n12708) );
  NAND2_X1 U15607 ( .A1(n12709), .A2(n12708), .ZN(n12710) );
  INV_X1 U15608 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20758) );
  NOR3_X1 U15609 ( .A1(P1_BE_N_REG_0__SCAN_IN), .A2(P1_BE_N_REG_1__SCAN_IN), 
        .A3(n20758), .ZN(n12712) );
  NOR4_X1 U15610 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n12711) );
  NAND4_X1 U15611 ( .A1(n14410), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n12712), .A4(
        n12711), .ZN(U214) );
  NOR2_X1 U15612 ( .A1(n15508), .A2(n12713), .ZN(n16423) );
  NAND2_X1 U15613 ( .A1(n16423), .A2(U214), .ZN(U212) );
  NAND2_X1 U15614 ( .A1(n12715), .A2(n12714), .ZN(n12718) );
  INV_X1 U15615 ( .A(n12716), .ZN(n12717) );
  NAND2_X1 U15616 ( .A1(n12718), .A2(n12717), .ZN(n19861) );
  AOI22_X1 U15617 ( .A1(n19861), .A2(n16306), .B1(n12719), .B2(n12864), .ZN(
        n12720) );
  OAI21_X1 U15618 ( .B1(n10277), .B2(n15445), .A(n12720), .ZN(n12735) );
  NOR2_X1 U15619 ( .A1(n12722), .A2(n12721), .ZN(n12734) );
  NAND2_X1 U15620 ( .A1(n12724), .A2(n12723), .ZN(n12806) );
  NAND3_X1 U15621 ( .A1(n12807), .A2(n16296), .A3(n12806), .ZN(n12725) );
  NAND2_X1 U15622 ( .A1(n19069), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n12809) );
  NAND2_X1 U15623 ( .A1(n12725), .A2(n12809), .ZN(n12733) );
  OAI21_X1 U15624 ( .B1(n12728), .B2(n12727), .A(n12726), .ZN(n12813) );
  AND2_X1 U15625 ( .A1(n12730), .A2(n12729), .ZN(n12731) );
  OAI22_X1 U15626 ( .A1(n12813), .A2(n16312), .B1(n12731), .B2(n15333), .ZN(
        n12732) );
  OR4_X1 U15627 ( .A1(n12735), .A2(n12734), .A3(n12733), .A4(n12732), .ZN(
        P2_U3044) );
  NAND2_X1 U15628 ( .A1(n12736), .A2(n12858), .ZN(n12737) );
  NOR2_X1 U15629 ( .A1(n10765), .A2(n12737), .ZN(n19113) );
  INV_X1 U15630 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n12740) );
  INV_X1 U15631 ( .A(n13595), .ZN(n12739) );
  NAND2_X1 U15632 ( .A1(n19844), .A2(n15828), .ZN(n18852) );
  OAI211_X1 U15633 ( .C1(n19113), .C2(n12740), .A(n12739), .B(n18852), .ZN(
        P2_U2814) );
  NOR2_X1 U15634 ( .A1(n19892), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n12742)
         );
  INV_X1 U15635 ( .A(n19899), .ZN(n12741) );
  AOI22_X1 U15636 ( .A1(n12742), .A2(n18852), .B1(n12741), .B2(n19892), .ZN(
        P2_U3612) );
  NOR4_X1 U15637 ( .A1(n12748), .A2(n12747), .A3(n12746), .A4(n12745), .ZN(
        n12749) );
  OR2_X1 U15638 ( .A1(n12750), .A2(n12749), .ZN(n14188) );
  INV_X1 U15639 ( .A(n14188), .ZN(n14195) );
  NAND3_X1 U15640 ( .A1(n12744), .A2(n14201), .A3(n14195), .ZN(n12791) );
  AND2_X1 U15641 ( .A1(n20585), .A2(n20669), .ZN(n13781) );
  AOI21_X1 U15642 ( .B1(n12791), .B2(P1_MEMORYFETCH_REG_SCAN_IN), .A(n13781), 
        .ZN(n12752) );
  INV_X1 U15643 ( .A(n12751), .ZN(n14194) );
  NAND2_X1 U15644 ( .A1(n12752), .A2(n12981), .ZN(P1_U2801) );
  INV_X1 U15645 ( .A(P2_EAX_REG_10__SCAN_IN), .ZN(n12755) );
  AND2_X1 U15646 ( .A1(n14806), .A2(n19898), .ZN(n12753) );
  NOR2_X2 U15647 ( .A1(n19206), .A2(n19204), .ZN(n19202) );
  NAND2_X1 U15648 ( .A1(n19202), .A2(P2_LWORD_REG_10__SCAN_IN), .ZN(n12754) );
  AOI22_X1 U15649 ( .A1(n15510), .A2(BUF1_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n12902), .ZN(n13048) );
  INV_X1 U15650 ( .A(n13048), .ZN(n14897) );
  NAND2_X1 U15651 ( .A1(n19204), .A2(n14897), .ZN(n12882) );
  OAI211_X1 U15652 ( .C1(n13598), .C2(n12755), .A(n12754), .B(n12882), .ZN(
        P2_U2977) );
  INV_X1 U15653 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n12757) );
  NAND2_X1 U15654 ( .A1(n19202), .A2(P2_UWORD_REG_0__SCAN_IN), .ZN(n12756) );
  AOI22_X1 U15655 ( .A1(n15510), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n12902), .ZN(n19170) );
  INV_X1 U15656 ( .A(n19170), .ZN(n14999) );
  NAND2_X1 U15657 ( .A1(n19204), .A2(n14999), .ZN(n12890) );
  OAI211_X1 U15658 ( .C1(n13598), .C2(n12757), .A(n12756), .B(n12890), .ZN(
        P2_U2952) );
  INV_X1 U15659 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n12759) );
  NAND2_X1 U15660 ( .A1(n19202), .A2(P2_LWORD_REG_11__SCAN_IN), .ZN(n12758) );
  AOI22_X1 U15661 ( .A1(n15510), .A2(BUF1_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n15508), .ZN(n13159) );
  INV_X1 U15662 ( .A(n13159), .ZN(n14886) );
  NAND2_X1 U15663 ( .A1(n19204), .A2(n14886), .ZN(n12886) );
  OAI211_X1 U15664 ( .C1(n13598), .C2(n12759), .A(n12758), .B(n12886), .ZN(
        P2_U2978) );
  INV_X1 U15665 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n12761) );
  NAND2_X1 U15666 ( .A1(n19202), .A2(P2_LWORD_REG_1__SCAN_IN), .ZN(n12760) );
  AOI22_X1 U15667 ( .A1(n15510), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n12902), .ZN(n19223) );
  INV_X1 U15668 ( .A(n19223), .ZN(n14984) );
  NAND2_X1 U15669 ( .A1(n19204), .A2(n14984), .ZN(n12884) );
  OAI211_X1 U15670 ( .C1(n13598), .C2(n12761), .A(n12760), .B(n12884), .ZN(
        P2_U2968) );
  INV_X1 U15671 ( .A(n19202), .ZN(n12790) );
  INV_X1 U15672 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n12763) );
  INV_X1 U15673 ( .A(n19204), .ZN(n12788) );
  AOI22_X1 U15674 ( .A1(n15510), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n12902), .ZN(n19239) );
  NOR2_X1 U15675 ( .A1(n12788), .A2(n19239), .ZN(n12778) );
  AOI21_X1 U15676 ( .B1(n19206), .B2(P2_EAX_REG_21__SCAN_IN), .A(n12778), .ZN(
        n12762) );
  OAI21_X1 U15677 ( .B1(n12790), .B2(n12763), .A(n12762), .ZN(P2_U2957) );
  INV_X1 U15678 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n12765) );
  AOI22_X1 U15679 ( .A1(n15510), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n12902), .ZN(n19254) );
  NOR2_X1 U15680 ( .A1(n12788), .A2(n19254), .ZN(n12768) );
  AOI21_X1 U15681 ( .B1(n19206), .B2(P2_EAX_REG_23__SCAN_IN), .A(n12768), .ZN(
        n12764) );
  OAI21_X1 U15682 ( .B1(n12790), .B2(n12765), .A(n12764), .ZN(P2_U2959) );
  INV_X1 U15683 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n12767) );
  AOI22_X1 U15684 ( .A1(n15510), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n15508), .ZN(n19246) );
  NOR2_X1 U15685 ( .A1(n12788), .A2(n19246), .ZN(n12771) );
  AOI21_X1 U15686 ( .B1(n19206), .B2(P2_EAX_REG_22__SCAN_IN), .A(n12771), .ZN(
        n12766) );
  OAI21_X1 U15687 ( .B1(n12790), .B2(n12767), .A(n12766), .ZN(P2_U2958) );
  INV_X1 U15688 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n12770) );
  AOI21_X1 U15689 ( .B1(n19206), .B2(P2_EAX_REG_7__SCAN_IN), .A(n12768), .ZN(
        n12769) );
  OAI21_X1 U15690 ( .B1(n12790), .B2(n12770), .A(n12769), .ZN(P2_U2974) );
  INV_X1 U15691 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n12773) );
  AOI21_X1 U15692 ( .B1(n19206), .B2(P2_EAX_REG_6__SCAN_IN), .A(n12771), .ZN(
        n12772) );
  OAI21_X1 U15693 ( .B1(n12790), .B2(n12773), .A(n12772), .ZN(P2_U2973) );
  INV_X1 U15694 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n12775) );
  AOI22_X1 U15695 ( .A1(n15510), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n12902), .ZN(n19234) );
  NOR2_X1 U15696 ( .A1(n12788), .A2(n19234), .ZN(n12781) );
  AOI21_X1 U15697 ( .B1(n19206), .B2(P2_EAX_REG_20__SCAN_IN), .A(n12781), .ZN(
        n12774) );
  OAI21_X1 U15698 ( .B1(n12790), .B2(n12775), .A(n12774), .ZN(P2_U2956) );
  INV_X1 U15699 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n12777) );
  AOI22_X1 U15700 ( .A1(n15510), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n15508), .ZN(n19231) );
  NOR2_X1 U15701 ( .A1(n12788), .A2(n19231), .ZN(n12784) );
  AOI21_X1 U15702 ( .B1(n19206), .B2(P2_EAX_REG_19__SCAN_IN), .A(n12784), .ZN(
        n12776) );
  OAI21_X1 U15703 ( .B1(n12790), .B2(n12777), .A(n12776), .ZN(P2_U2955) );
  INV_X1 U15704 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n12780) );
  AOI21_X1 U15705 ( .B1(P2_EAX_REG_5__SCAN_IN), .B2(n19206), .A(n12778), .ZN(
        n12779) );
  OAI21_X1 U15706 ( .B1(n12790), .B2(n12780), .A(n12779), .ZN(P2_U2972) );
  INV_X1 U15707 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n12783) );
  AOI21_X1 U15708 ( .B1(n19206), .B2(P2_EAX_REG_4__SCAN_IN), .A(n12781), .ZN(
        n12782) );
  OAI21_X1 U15709 ( .B1(n12790), .B2(n12783), .A(n12782), .ZN(P2_U2971) );
  INV_X1 U15710 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n12786) );
  AOI21_X1 U15711 ( .B1(n19206), .B2(P2_EAX_REG_3__SCAN_IN), .A(n12784), .ZN(
        n12785) );
  OAI21_X1 U15712 ( .B1(n12790), .B2(n12786), .A(n12785), .ZN(P2_U2970) );
  INV_X1 U15713 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n12789) );
  AOI22_X1 U15714 ( .A1(n15510), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n15508), .ZN(n13584) );
  INV_X1 U15715 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n12787) );
  OAI222_X1 U15716 ( .A1(n12790), .A2(n12789), .B1(n12788), .B2(n13584), .C1(
        n12787), .C2(n13598), .ZN(P2_U2982) );
  INV_X1 U15717 ( .A(n20765), .ZN(n12793) );
  OAI21_X1 U15718 ( .B1(n13781), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n12793), 
        .ZN(n12792) );
  OAI21_X1 U15719 ( .B1(n12794), .B2(n12793), .A(n12792), .ZN(P1_U3487) );
  NOR2_X1 U15720 ( .A1(n12795), .A2(n10765), .ZN(n12834) );
  NAND2_X1 U15721 ( .A1(n12834), .A2(n13288), .ZN(n12799) );
  INV_X1 U15722 ( .A(n15479), .ZN(n13285) );
  NAND2_X1 U15723 ( .A1(n13285), .A2(n13283), .ZN(n12857) );
  AND3_X1 U15724 ( .A1(n12797), .A2(n12857), .A3(n12796), .ZN(n12798) );
  NAND2_X1 U15725 ( .A1(n12799), .A2(n12798), .ZN(n13308) );
  NOR2_X1 U15726 ( .A1(n15828), .A2(n19691), .ZN(n16320) );
  NAND2_X1 U15727 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16320), .ZN(n15829) );
  OAI22_X1 U15728 ( .A1(n19697), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n18860), 
        .B2(n15829), .ZN(n12800) );
  AOI21_X1 U15729 ( .B1(n13308), .B2(n12858), .A(n12800), .ZN(n15498) );
  INV_X1 U15730 ( .A(n15498), .ZN(n12805) );
  NAND2_X1 U15731 ( .A1(n10178), .A2(n12803), .ZN(n13294) );
  OR4_X1 U15732 ( .A1(n15498), .A2(n19848), .A3(n12801), .A4(n13294), .ZN(
        n12804) );
  OAI21_X1 U15733 ( .B1(n12805), .B2(n20796), .A(n12804), .ZN(P2_U3595) );
  NAND3_X1 U15734 ( .A1(n12807), .A2(n16282), .A3(n12806), .ZN(n12812) );
  AOI21_X1 U15735 ( .B1(n19102), .B2(n12808), .A(n13395), .ZN(n13668) );
  OAI21_X1 U15736 ( .B1(n16288), .B2(n12808), .A(n12809), .ZN(n12810) );
  AOI21_X1 U15737 ( .B1(n16279), .B2(n13668), .A(n12810), .ZN(n12811) );
  OAI211_X1 U15738 ( .C1(n12813), .C2(n16260), .A(n12812), .B(n12811), .ZN(
        n12814) );
  AOI21_X1 U15739 ( .B1(n9656), .B2(n16281), .A(n12814), .ZN(n12815) );
  INV_X1 U15740 ( .A(n12815), .ZN(P2_U3012) );
  OAI21_X1 U15741 ( .B1(n12817), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12816), .ZN(n16311) );
  OAI21_X1 U15742 ( .B1(n16252), .B2(n12818), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n12821) );
  OAI21_X1 U15743 ( .B1(n14763), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n12825), .ZN(n16309) );
  INV_X1 U15744 ( .A(n16309), .ZN(n12819) );
  NOR2_X1 U15745 ( .A1(n19089), .A2(n14759), .ZN(n16314) );
  AOI21_X1 U15746 ( .B1(n16282), .B2(n12819), .A(n16314), .ZN(n12820) );
  OAI211_X1 U15747 ( .C1(n16260), .C2(n16311), .A(n12821), .B(n12820), .ZN(
        n12822) );
  AOI21_X1 U15748 ( .B1(n16315), .B2(n16281), .A(n12822), .ZN(n12823) );
  INV_X1 U15749 ( .A(n12823), .ZN(P2_U3014) );
  OAI21_X1 U15750 ( .B1(n12825), .B2(n19100), .A(n12824), .ZN(n12826) );
  XOR2_X1 U15751 ( .A(n12826), .B(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n12871) );
  INV_X1 U15752 ( .A(n12871), .ZN(n12832) );
  AND2_X1 U15753 ( .A1(n19069), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n12868) );
  OAI21_X1 U15754 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n12828), .A(
        n12827), .ZN(n12865) );
  NOR2_X1 U15755 ( .A1(n16260), .A2(n12865), .ZN(n12829) );
  AOI211_X1 U15756 ( .C1(n16252), .C2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n12868), .B(n12829), .ZN(n12830) );
  OAI21_X1 U15757 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n16257), .A(
        n12830), .ZN(n12831) );
  AOI21_X1 U15758 ( .B1(n16282), .B2(n12832), .A(n12831), .ZN(n12833) );
  OAI21_X1 U15759 ( .B1(n12860), .B2(n15182), .A(n12833), .ZN(P2_U3013) );
  INV_X1 U15760 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n12840) );
  NAND2_X1 U15761 ( .A1(n12834), .A2(n12858), .ZN(n12835) );
  NAND2_X1 U15762 ( .A1(n12835), .A2(n13598), .ZN(n12836) );
  INV_X1 U15763 ( .A(n19895), .ZN(n19763) );
  NAND2_X1 U15764 ( .A1(n16320), .A2(n18853), .ZN(n12838) );
  INV_X2 U15765 ( .A(n12838), .ZN(n19181) );
  AOI22_X1 U15766 ( .A1(n19181), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n12839) );
  OAI21_X1 U15767 ( .B1(n12840), .B2(n19172), .A(n12839), .ZN(P2_U2932) );
  INV_X1 U15768 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n14945) );
  AOI22_X1 U15769 ( .A1(n19181), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n12841) );
  OAI21_X1 U15770 ( .B1(n14945), .B2(n19172), .A(n12841), .ZN(P2_U2930) );
  INV_X1 U15771 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n14972) );
  AOI22_X1 U15772 ( .A1(n19181), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n12842) );
  OAI21_X1 U15773 ( .B1(n14972), .B2(n19172), .A(n12842), .ZN(P2_U2933) );
  INV_X1 U15774 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n20911) );
  AOI22_X1 U15775 ( .A1(n19181), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n12843) );
  OAI21_X1 U15776 ( .B1(n20911), .B2(n19172), .A(n12843), .ZN(P2_U2931) );
  INV_X1 U15777 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n12845) );
  AOI22_X1 U15778 ( .A1(n19181), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n12844) );
  OAI21_X1 U15779 ( .B1(n12845), .B2(n19172), .A(n12844), .ZN(P2_U2928) );
  INV_X1 U15780 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n12911) );
  AOI22_X1 U15781 ( .A1(n19181), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n12846) );
  OAI21_X1 U15782 ( .B1(n12911), .B2(n19172), .A(n12846), .ZN(P2_U2927) );
  INV_X1 U15783 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n14935) );
  AOI22_X1 U15784 ( .A1(n19181), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n12847) );
  OAI21_X1 U15785 ( .B1(n14935), .B2(n19172), .A(n12847), .ZN(P2_U2929) );
  INV_X1 U15786 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n14894) );
  AOI22_X1 U15787 ( .A1(n19181), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n12848) );
  OAI21_X1 U15788 ( .B1(n14894), .B2(n19172), .A(n12848), .ZN(P2_U2925) );
  INV_X1 U15789 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n14884) );
  AOI22_X1 U15790 ( .A1(n19181), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n12849) );
  OAI21_X1 U15791 ( .B1(n14884), .B2(n19172), .A(n12849), .ZN(P2_U2924) );
  INV_X1 U15792 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n12905) );
  AOI22_X1 U15793 ( .A1(n19181), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n12850) );
  OAI21_X1 U15794 ( .B1(n12905), .B2(n19172), .A(n12850), .ZN(P2_U2926) );
  INV_X1 U15795 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n14866) );
  AOI22_X1 U15796 ( .A1(n19181), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n12851) );
  OAI21_X1 U15797 ( .B1(n14866), .B2(n19172), .A(n12851), .ZN(P2_U2922) );
  AOI22_X1 U15798 ( .A1(n19181), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n12852) );
  OAI21_X1 U15799 ( .B1(n12757), .B2(n19172), .A(n12852), .ZN(P2_U2935) );
  INV_X1 U15800 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n14982) );
  AOI22_X1 U15801 ( .A1(n19181), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n12853) );
  OAI21_X1 U15802 ( .B1(n14982), .B2(n19172), .A(n12853), .ZN(P2_U2934) );
  INV_X1 U15803 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n14877) );
  AOI22_X1 U15804 ( .A1(n19181), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n12854) );
  OAI21_X1 U15805 ( .B1(n14877), .B2(n19172), .A(n12854), .ZN(P2_U2923) );
  NAND2_X1 U15806 ( .A1(n12857), .A2(n11192), .ZN(n12859) );
  MUX2_X1 U15807 ( .A(n19103), .B(n12860), .S(n13520), .Z(n12861) );
  OAI21_X1 U15808 ( .B1(n19209), .B2(n14865), .A(n12861), .ZN(P2_U2886) );
  XNOR2_X1 U15809 ( .A(n12863), .B(n12862), .ZN(n19866) );
  AOI22_X1 U15810 ( .A1(n11297), .A2(n16316), .B1(n16306), .B2(n19866), .ZN(
        n12870) );
  INV_X1 U15811 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15489) );
  AOI211_X1 U15812 ( .C1(n16304), .C2(n15489), .A(n12864), .B(n16319), .ZN(
        n12867) );
  OAI22_X1 U15813 ( .A1(n15489), .A2(n16305), .B1(n16312), .B2(n12865), .ZN(
        n12866) );
  NOR3_X1 U15814 ( .A1(n12868), .A2(n12867), .A3(n12866), .ZN(n12869) );
  OAI211_X1 U15815 ( .C1(n12871), .C2(n16310), .A(n12870), .B(n12869), .ZN(
        P2_U3045) );
  MUX2_X1 U15816 ( .A(n9656), .B(P2_EBX_REG_2__SCAN_IN), .S(n14856), .Z(n12874) );
  INV_X1 U15817 ( .A(n12874), .ZN(n12875) );
  OAI21_X1 U15818 ( .B1(n19859), .B2(n14865), .A(n12875), .ZN(P2_U2885) );
  NAND2_X1 U15819 ( .A1(n14806), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n12876) );
  NAND4_X1 U15820 ( .A1(n10197), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n12876), 
        .A4(n19697), .ZN(n12877) );
  NOR2_X1 U15821 ( .A1(n14760), .A2(n14856), .ZN(n12879) );
  AOI21_X1 U15822 ( .B1(P2_EBX_REG_0__SCAN_IN), .B2(n14856), .A(n12879), .ZN(
        n12880) );
  OAI21_X1 U15823 ( .B1(n14865), .B2(n19210), .A(n12880), .ZN(P2_U2887) );
  NAND2_X1 U15824 ( .A1(n19202), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n12881) );
  AOI22_X1 U15825 ( .A1(n15510), .A2(BUF1_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n12902), .ZN(n13248) );
  INV_X1 U15826 ( .A(n13248), .ZN(n14869) );
  NAND2_X1 U15827 ( .A1(n19204), .A2(n14869), .ZN(n12906) );
  OAI211_X1 U15828 ( .C1(n13598), .C2(n14866), .A(n12881), .B(n12906), .ZN(
        P2_U2965) );
  NAND2_X1 U15829 ( .A1(n19202), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n12883) );
  OAI211_X1 U15830 ( .C1(n13598), .C2(n14894), .A(n12883), .B(n12882), .ZN(
        P2_U2962) );
  NAND2_X1 U15831 ( .A1(n19202), .A2(P2_UWORD_REG_1__SCAN_IN), .ZN(n12885) );
  OAI211_X1 U15832 ( .C1(n13598), .C2(n14982), .A(n12885), .B(n12884), .ZN(
        P2_U2953) );
  NAND2_X1 U15833 ( .A1(n19202), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n12887) );
  OAI211_X1 U15834 ( .C1(n13598), .C2(n14884), .A(n12887), .B(n12886), .ZN(
        P2_U2963) );
  INV_X1 U15835 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n12889) );
  NAND2_X1 U15836 ( .A1(n19202), .A2(P2_LWORD_REG_2__SCAN_IN), .ZN(n12888) );
  AOI22_X1 U15837 ( .A1(n15510), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n12902), .ZN(n19227) );
  INV_X1 U15838 ( .A(n19227), .ZN(n14976) );
  NAND2_X1 U15839 ( .A1(n19204), .A2(n14976), .ZN(n12896) );
  OAI211_X1 U15840 ( .C1(n13598), .C2(n12889), .A(n12888), .B(n12896), .ZN(
        P2_U2969) );
  INV_X1 U15841 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n12892) );
  NAND2_X1 U15842 ( .A1(n19202), .A2(P2_LWORD_REG_0__SCAN_IN), .ZN(n12891) );
  OAI211_X1 U15843 ( .C1(n12892), .C2(n13598), .A(n12891), .B(n12890), .ZN(
        P2_U2967) );
  INV_X1 U15844 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19187) );
  NAND2_X1 U15845 ( .A1(n19202), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n12895) );
  INV_X1 U15846 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16459) );
  OR2_X1 U15847 ( .A1(n15508), .A2(n16459), .ZN(n12894) );
  NAND2_X1 U15848 ( .A1(n15508), .A2(BUF2_REG_8__SCAN_IN), .ZN(n12893) );
  NAND2_X1 U15849 ( .A1(n12894), .A2(n12893), .ZN(n19130) );
  NAND2_X1 U15850 ( .A1(n19204), .A2(n19130), .ZN(n12909) );
  OAI211_X1 U15851 ( .C1(n19187), .C2(n13598), .A(n12895), .B(n12909), .ZN(
        P2_U2975) );
  NAND2_X1 U15852 ( .A1(n19202), .A2(P2_UWORD_REG_2__SCAN_IN), .ZN(n12897) );
  OAI211_X1 U15853 ( .C1(n13598), .C2(n14972), .A(n12897), .B(n12896), .ZN(
        P2_U2954) );
  NAND2_X1 U15854 ( .A1(n19202), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n12898) );
  MUX2_X1 U15855 ( .A(BUF1_REG_12__SCAN_IN), .B(BUF2_REG_12__SCAN_IN), .S(
        n15508), .Z(n14879) );
  NAND2_X1 U15856 ( .A1(n19204), .A2(n14879), .ZN(n12899) );
  OAI211_X1 U15857 ( .C1(n13598), .C2(n14877), .A(n12898), .B(n12899), .ZN(
        P2_U2964) );
  INV_X1 U15858 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n12901) );
  NAND2_X1 U15859 ( .A1(n19202), .A2(P2_LWORD_REG_12__SCAN_IN), .ZN(n12900) );
  OAI211_X1 U15860 ( .C1(n13598), .C2(n12901), .A(n12900), .B(n12899), .ZN(
        P2_U2979) );
  NAND2_X1 U15861 ( .A1(n19202), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n12904) );
  AOI22_X1 U15862 ( .A1(n15510), .A2(BUF1_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n12902), .ZN(n14906) );
  INV_X1 U15863 ( .A(n14906), .ZN(n12903) );
  NAND2_X1 U15864 ( .A1(n19204), .A2(n12903), .ZN(n12912) );
  OAI211_X1 U15865 ( .C1(n13598), .C2(n12905), .A(n12904), .B(n12912), .ZN(
        P2_U2961) );
  INV_X1 U15866 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n12908) );
  NAND2_X1 U15867 ( .A1(n19202), .A2(P2_LWORD_REG_13__SCAN_IN), .ZN(n12907) );
  OAI211_X1 U15868 ( .C1(n13598), .C2(n12908), .A(n12907), .B(n12906), .ZN(
        P2_U2980) );
  NAND2_X1 U15869 ( .A1(n19202), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n12910) );
  OAI211_X1 U15870 ( .C1(n12911), .C2(n13598), .A(n12910), .B(n12909), .ZN(
        P2_U2960) );
  INV_X1 U15871 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n12914) );
  NAND2_X1 U15872 ( .A1(n19202), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n12913) );
  OAI211_X1 U15873 ( .C1(n13598), .C2(n12914), .A(n12913), .B(n12912), .ZN(
        P2_U2976) );
  INV_X1 U15874 ( .A(n10285), .ZN(n13388) );
  MUX2_X1 U15875 ( .A(n13388), .B(n12918), .S(n14856), .Z(n12919) );
  OAI21_X1 U15876 ( .B1(n19484), .B2(n14865), .A(n12919), .ZN(P2_U2884) );
  OAI21_X1 U15877 ( .B1(n12921), .B2(n12920), .A(n16290), .ZN(n19051) );
  AND2_X1 U15878 ( .A1(n15002), .A2(n19153), .ZN(n19143) );
  INV_X1 U15879 ( .A(n12922), .ZN(n12923) );
  OAI222_X1 U15880 ( .A1(n19051), .A2(n19143), .B1(n19152), .B2(n19189), .C1(
        n19169), .C2(n19254), .ZN(P2_U2912) );
  XNOR2_X1 U15881 ( .A(n12925), .B(n12924), .ZN(n19063) );
  INV_X1 U15882 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19191) );
  OAI222_X1 U15883 ( .A1(n19063), .A2(n19143), .B1(n19152), .B2(n19191), .C1(
        n19169), .C2(n19246), .ZN(P2_U2913) );
  INV_X1 U15884 ( .A(n13328), .ZN(n13440) );
  NOR2_X1 U15885 ( .A1(n12926), .A2(n13440), .ZN(n12927) );
  XNOR2_X1 U15886 ( .A(n12927), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n19998) );
  NAND2_X1 U15887 ( .A1(READY11_REG_SCAN_IN), .A2(READY1), .ZN(n20767) );
  INV_X1 U15888 ( .A(n20767), .ZN(n12979) );
  NOR2_X1 U15889 ( .A1(n12979), .A2(n14188), .ZN(n13729) );
  INV_X1 U15890 ( .A(n12928), .ZN(n12951) );
  NAND2_X1 U15891 ( .A1(n13729), .A2(n12951), .ZN(n12933) );
  NAND2_X1 U15892 ( .A1(n12929), .A2(n20767), .ZN(n15788) );
  INV_X1 U15893 ( .A(n12930), .ZN(n13742) );
  NAND2_X1 U15894 ( .A1(n13742), .A2(n13740), .ZN(n13178) );
  OAI21_X1 U15895 ( .B1(n15788), .B2(n14198), .A(n13178), .ZN(n12931) );
  NAND2_X1 U15896 ( .A1(n12931), .A2(n13730), .ZN(n12932) );
  INV_X1 U15897 ( .A(n13118), .ZN(n12948) );
  AND2_X1 U15898 ( .A1(n12744), .A2(n13734), .ZN(n15762) );
  INV_X1 U15899 ( .A(n12934), .ZN(n12936) );
  INV_X1 U15900 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n12935) );
  NAND2_X1 U15901 ( .A1(n12936), .A2(n12935), .ZN(n15826) );
  OAI211_X1 U15902 ( .C1(n15762), .C2(n12929), .A(n20767), .B(n15789), .ZN(
        n12944) );
  INV_X1 U15903 ( .A(n12744), .ZN(n12941) );
  NOR2_X1 U15904 ( .A1(n12937), .A2(n13340), .ZN(n12945) );
  NOR2_X1 U15905 ( .A1(n12945), .A2(n13638), .ZN(n12938) );
  NAND2_X1 U15906 ( .A1(n12939), .A2(n12938), .ZN(n13175) );
  NAND2_X1 U15907 ( .A1(n13742), .A2(n13175), .ZN(n12940) );
  NAND2_X1 U15908 ( .A1(n12941), .A2(n12940), .ZN(n13736) );
  OR2_X1 U15909 ( .A1(n13637), .A2(n13352), .ZN(n12942) );
  AND2_X1 U15910 ( .A1(n13736), .A2(n12942), .ZN(n12943) );
  AND2_X1 U15911 ( .A1(n12944), .A2(n12943), .ZN(n12947) );
  NAND2_X1 U15912 ( .A1(n12946), .A2(n12945), .ZN(n14191) );
  NAND3_X1 U15913 ( .A1(n12948), .A2(n12947), .A3(n13405), .ZN(n15759) );
  INV_X1 U15914 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19919) );
  NAND2_X1 U15915 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n16110) );
  INV_X1 U15916 ( .A(n16110), .ZN(n14733) );
  NAND2_X1 U15917 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n14733), .ZN(n16114) );
  NOR2_X1 U15918 ( .A1(n19919), .A2(n16114), .ZN(n12950) );
  NOR2_X1 U15919 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20379), .ZN(n12949) );
  AOI211_X1 U15920 ( .C1(n15759), .C2(n14201), .A(n12950), .B(n12949), .ZN(
        n14109) );
  INV_X1 U15921 ( .A(n14109), .ZN(n20748) );
  NAND3_X1 U15922 ( .A1(n20748), .A2(n19909), .A3(n12951), .ZN(n12952) );
  OAI22_X1 U15923 ( .A1(n19998), .A2(n12952), .B1(n12027), .B2(n20748), .ZN(
        P1_U3468) );
  AND2_X1 U15924 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n12955) );
  NAND2_X1 U15925 ( .A1(n12953), .A2(n12955), .ZN(n13026) );
  OR2_X1 U15926 ( .A1(n12953), .A2(n12955), .ZN(n12956) );
  NAND2_X1 U15927 ( .A1(n13026), .A2(n12956), .ZN(n19146) );
  OR2_X1 U15928 ( .A1(n12958), .A2(n12957), .ZN(n12959) );
  NAND2_X1 U15929 ( .A1(n13030), .A2(n12959), .ZN(n19092) );
  MUX2_X1 U15930 ( .A(n19092), .B(n19084), .S(n14856), .Z(n12960) );
  OAI21_X1 U15931 ( .B1(n19146), .B2(n14865), .A(n12960), .ZN(P2_U2883) );
  INV_X1 U15932 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n12966) );
  INV_X1 U15933 ( .A(n15762), .ZN(n12961) );
  NAND2_X1 U15934 ( .A1(n12929), .A2(n20762), .ZN(n13758) );
  NAND2_X1 U15935 ( .A1(n12961), .A2(n13758), .ZN(n12964) );
  INV_X1 U15936 ( .A(n15789), .ZN(n12962) );
  NOR2_X1 U15937 ( .A1(n19911), .A2(n12962), .ZN(n12963) );
  NAND2_X1 U15938 ( .A1(n20043), .A2(n11848), .ZN(n13141) );
  NOR2_X1 U15939 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16110), .ZN(n20065) );
  NOR2_X4 U15940 ( .A1(n20043), .A2(n20768), .ZN(n20064) );
  AOI22_X1 U15941 ( .A1(P1_UWORD_REG_8__SCAN_IN), .A2(n20768), .B1(n20064), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n12965) );
  OAI21_X1 U15942 ( .B1(n12966), .B2(n13141), .A(n12965), .ZN(P1_U2912) );
  INV_X1 U15943 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n12968) );
  AOI22_X1 U15944 ( .A1(P1_UWORD_REG_14__SCAN_IN), .A2(n20768), .B1(n20064), 
        .B2(P1_DATAO_REG_30__SCAN_IN), .ZN(n12967) );
  OAI21_X1 U15945 ( .B1(n12968), .B2(n13141), .A(n12967), .ZN(P1_U2906) );
  INV_X1 U15946 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n12970) );
  AOI22_X1 U15947 ( .A1(P1_UWORD_REG_10__SCAN_IN), .A2(n20768), .B1(n20064), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n12969) );
  OAI21_X1 U15948 ( .B1(n12970), .B2(n13141), .A(n12969), .ZN(P1_U2910) );
  INV_X1 U15949 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n12972) );
  AOI22_X1 U15950 ( .A1(P1_UWORD_REG_9__SCAN_IN), .A2(n20768), .B1(n20064), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n12971) );
  OAI21_X1 U15951 ( .B1(n12972), .B2(n13141), .A(n12971), .ZN(P1_U2911) );
  INV_X1 U15952 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n12974) );
  AOI22_X1 U15953 ( .A1(P1_UWORD_REG_13__SCAN_IN), .A2(n20768), .B1(n20064), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n12973) );
  OAI21_X1 U15954 ( .B1(n12974), .B2(n13141), .A(n12973), .ZN(P1_U2907) );
  INV_X1 U15955 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n12976) );
  AOI22_X1 U15956 ( .A1(P1_UWORD_REG_11__SCAN_IN), .A2(n20768), .B1(n20064), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n12975) );
  OAI21_X1 U15957 ( .B1(n12976), .B2(n13141), .A(n12975), .ZN(P1_U2909) );
  INV_X1 U15958 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n12978) );
  AOI22_X1 U15959 ( .A1(P1_UWORD_REG_12__SCAN_IN), .A2(n20768), .B1(n20064), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n12977) );
  OAI21_X1 U15960 ( .B1(n12978), .B2(n13141), .A(n12977), .ZN(P1_U2908) );
  AND2_X1 U15961 ( .A1(n15791), .A2(n12979), .ZN(n12980) );
  OR2_X1 U15962 ( .A1(n20075), .A2(n13734), .ZN(n13077) );
  INV_X1 U15963 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n12986) );
  NOR2_X2 U15964 ( .A1(n20075), .A2(n13639), .ZN(n20088) );
  INV_X1 U15965 ( .A(n20088), .ZN(n12985) );
  INV_X1 U15966 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n12982) );
  NOR2_X1 U15967 ( .A1(n13861), .A2(n12982), .ZN(n12983) );
  AOI21_X1 U15968 ( .B1(DATAI_15_), .B2(n13861), .A(n12983), .ZN(n14471) );
  INV_X1 U15969 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n12984) );
  OAI222_X1 U15970 ( .A1(n13077), .A2(n12986), .B1(n12985), .B2(n14471), .C1(
        n12984), .C2(n12999), .ZN(P1_U2967) );
  XNOR2_X1 U15971 ( .A(n19209), .B(n19866), .ZN(n12991) );
  NOR2_X1 U15972 ( .A1(n12988), .A2(n12987), .ZN(n12989) );
  NOR2_X1 U15973 ( .A1(n12990), .A2(n12989), .ZN(n19166) );
  NAND2_X1 U15974 ( .A1(n19877), .A2(n19166), .ZN(n19165) );
  NAND2_X1 U15975 ( .A1(n12991), .A2(n19165), .ZN(n13037) );
  OAI21_X1 U15976 ( .B1(n12991), .B2(n19165), .A(n13037), .ZN(n12992) );
  NAND2_X1 U15977 ( .A1(n12992), .A2(n19164), .ZN(n12994) );
  INV_X1 U15978 ( .A(n19153), .ZN(n19163) );
  AOI22_X1 U15979 ( .A1(n19163), .A2(n19866), .B1(n19162), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n12993) );
  OAI211_X1 U15980 ( .C1(n19223), .C2(n19169), .A(n12994), .B(n12993), .ZN(
        P2_U2918) );
  INV_X1 U15981 ( .A(n13077), .ZN(n20076) );
  AOI22_X1 U15982 ( .A1(n20076), .A2(P1_EAX_REG_11__SCAN_IN), .B1(
        P1_LWORD_REG_11__SCAN_IN), .B2(n20100), .ZN(n12998) );
  INV_X1 U15983 ( .A(DATAI_11_), .ZN(n12996) );
  INV_X1 U15984 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n12995) );
  MUX2_X1 U15985 ( .A(n12996), .B(n12995), .S(n14410), .Z(n14420) );
  INV_X1 U15986 ( .A(n14420), .ZN(n12997) );
  NAND2_X1 U15987 ( .A1(n20088), .A2(n12997), .ZN(n13086) );
  NAND2_X1 U15988 ( .A1(n12998), .A2(n13086), .ZN(P1_U2963) );
  INV_X1 U15989 ( .A(n12999), .ZN(n20100) );
  AOI22_X1 U15990 ( .A1(n20076), .A2(P1_EAX_REG_5__SCAN_IN), .B1(
        P1_LWORD_REG_5__SCAN_IN), .B2(n20100), .ZN(n13003) );
  NAND2_X1 U15991 ( .A1(n13861), .A2(DATAI_5_), .ZN(n13001) );
  NAND2_X1 U15992 ( .A1(n14410), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13000) );
  AND2_X1 U15993 ( .A1(n13001), .A2(n13000), .ZN(n14447) );
  INV_X1 U15994 ( .A(n14447), .ZN(n13002) );
  NAND2_X1 U15995 ( .A1(n20088), .A2(n13002), .ZN(n13078) );
  NAND2_X1 U15996 ( .A1(n13003), .A2(n13078), .ZN(P1_U2957) );
  AOI22_X1 U15997 ( .A1(n20076), .A2(P1_EAX_REG_7__SCAN_IN), .B1(
        P1_LWORD_REG_7__SCAN_IN), .B2(n20100), .ZN(n13007) );
  NAND2_X1 U15998 ( .A1(n13861), .A2(DATAI_7_), .ZN(n13005) );
  NAND2_X1 U15999 ( .A1(n14410), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13004) );
  AND2_X1 U16000 ( .A1(n13005), .A2(n13004), .ZN(n14438) );
  INV_X1 U16001 ( .A(n14438), .ZN(n13006) );
  NAND2_X1 U16002 ( .A1(n20088), .A2(n13006), .ZN(n13080) );
  NAND2_X1 U16003 ( .A1(n13007), .A2(n13080), .ZN(P1_U2959) );
  AOI22_X1 U16004 ( .A1(n20076), .A2(P1_EAX_REG_6__SCAN_IN), .B1(
        P1_LWORD_REG_6__SCAN_IN), .B2(n20100), .ZN(n13011) );
  NAND2_X1 U16005 ( .A1(n13861), .A2(DATAI_6_), .ZN(n13009) );
  NAND2_X1 U16006 ( .A1(n14410), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13008) );
  AND2_X1 U16007 ( .A1(n13009), .A2(n13008), .ZN(n14442) );
  INV_X1 U16008 ( .A(n14442), .ZN(n13010) );
  NAND2_X1 U16009 ( .A1(n20088), .A2(n13010), .ZN(n13084) );
  NAND2_X1 U16010 ( .A1(n13011), .A2(n13084), .ZN(P1_U2958) );
  AOI22_X1 U16011 ( .A1(n20076), .A2(P1_EAX_REG_3__SCAN_IN), .B1(
        P1_LWORD_REG_3__SCAN_IN), .B2(n20100), .ZN(n13015) );
  NAND2_X1 U16012 ( .A1(n13861), .A2(DATAI_3_), .ZN(n13013) );
  NAND2_X1 U16013 ( .A1(n14410), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13012) );
  AND2_X1 U16014 ( .A1(n13013), .A2(n13012), .ZN(n14456) );
  INV_X1 U16015 ( .A(n14456), .ZN(n13014) );
  NAND2_X1 U16016 ( .A1(n20088), .A2(n13014), .ZN(n13082) );
  NAND2_X1 U16017 ( .A1(n13015), .A2(n13082), .ZN(P1_U2955) );
  AOI22_X1 U16018 ( .A1(n20076), .A2(P1_EAX_REG_4__SCAN_IN), .B1(
        P1_LWORD_REG_4__SCAN_IN), .B2(n20100), .ZN(n13019) );
  NAND2_X1 U16019 ( .A1(n13861), .A2(DATAI_4_), .ZN(n13017) );
  NAND2_X1 U16020 ( .A1(n14410), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13016) );
  AND2_X1 U16021 ( .A1(n13017), .A2(n13016), .ZN(n14451) );
  INV_X1 U16022 ( .A(n14451), .ZN(n13018) );
  NAND2_X1 U16023 ( .A1(n20088), .A2(n13018), .ZN(n13088) );
  NAND2_X1 U16024 ( .A1(n13019), .A2(n13088), .ZN(P1_U2956) );
  NOR2_X1 U16025 ( .A1(n13026), .A2(n13020), .ZN(n13069) );
  XNOR2_X1 U16026 ( .A(n13069), .B(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13025) );
  AND2_X1 U16027 ( .A1(n13032), .A2(n13021), .ZN(n13022) );
  OR2_X1 U16028 ( .A1(n13022), .A2(n13073), .ZN(n15468) );
  INV_X1 U16029 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13023) );
  MUX2_X1 U16030 ( .A(n15468), .B(n13023), .S(n14856), .Z(n13024) );
  OAI21_X1 U16031 ( .B1(n13025), .B2(n14865), .A(n13024), .ZN(P2_U2881) );
  INV_X1 U16032 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n13035) );
  INV_X1 U16033 ( .A(n13026), .ZN(n13028) );
  INV_X1 U16034 ( .A(n13069), .ZN(n13027) );
  OAI211_X1 U16035 ( .C1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .C2(n13028), .A(
        n13027), .B(n14844), .ZN(n13034) );
  NAND2_X1 U16036 ( .A1(n13030), .A2(n13029), .ZN(n13031) );
  AND2_X1 U16037 ( .A1(n13032), .A2(n13031), .ZN(n19074) );
  NAND2_X1 U16038 ( .A1(n19074), .A2(n13520), .ZN(n13033) );
  OAI211_X1 U16039 ( .C1(n13520), .C2(n13035), .A(n13034), .B(n13033), .ZN(
        P2_U2882) );
  INV_X1 U16040 ( .A(n19861), .ZN(n19135) );
  XNOR2_X1 U16041 ( .A(n19859), .B(n19861), .ZN(n13040) );
  INV_X1 U16042 ( .A(n19866), .ZN(n13036) );
  NAND2_X1 U16043 ( .A1(n19209), .A2(n13036), .ZN(n13038) );
  NAND2_X1 U16044 ( .A1(n13038), .A2(n13037), .ZN(n13039) );
  NAND2_X1 U16045 ( .A1(n13040), .A2(n13039), .ZN(n19136) );
  OAI21_X1 U16046 ( .B1(n13040), .B2(n13039), .A(n19136), .ZN(n13041) );
  NAND2_X1 U16047 ( .A1(n13041), .A2(n19164), .ZN(n13043) );
  AOI22_X1 U16048 ( .A1(n19134), .A2(n14976), .B1(n19162), .B2(
        P2_EAX_REG_2__SCAN_IN), .ZN(n13042) );
  OAI211_X1 U16049 ( .C1(n19135), .C2(n19153), .A(n13043), .B(n13042), .ZN(
        P2_U2917) );
  OAI21_X1 U16050 ( .B1(n13044), .B2(n13045), .A(n13047), .ZN(n19030) );
  OAI222_X1 U16051 ( .A1(n19152), .A2(n12914), .B1(n14906), .B2(n19169), .C1(
        n19030), .C2(n19143), .ZN(P2_U2910) );
  XNOR2_X1 U16052 ( .A(n13047), .B(n13046), .ZN(n19019) );
  OAI222_X1 U16053 ( .A1(n19019), .A2(n19143), .B1(n13048), .B2(n19169), .C1(
        n12755), .C2(n19152), .ZN(P2_U2909) );
  INV_X1 U16054 ( .A(n13049), .ZN(n13066) );
  NAND2_X1 U16055 ( .A1(n13066), .A2(n13050), .ZN(n13051) );
  AND2_X1 U16056 ( .A1(n13143), .A2(n13051), .ZN(n19027) );
  NAND2_X1 U16057 ( .A1(n19027), .A2(n13520), .ZN(n13059) );
  INV_X1 U16058 ( .A(n13053), .ZN(n13057) );
  OAI211_X1 U16059 ( .C1(n13057), .C2(n13056), .A(n14844), .B(n13055), .ZN(
        n13058) );
  OAI211_X1 U16060 ( .C1(n13520), .C2(n13060), .A(n13059), .B(n13058), .ZN(
        P2_U2878) );
  AND2_X1 U16061 ( .A1(n13069), .A2(n13061), .ZN(n13070) );
  OAI211_X1 U16062 ( .C1(n13070), .C2(n13062), .A(n14844), .B(n13053), .ZN(
        n13068) );
  NAND2_X1 U16063 ( .A1(n13063), .A2(n13064), .ZN(n13065) );
  NAND2_X1 U16064 ( .A1(n13066), .A2(n13065), .ZN(n19040) );
  INV_X1 U16065 ( .A(n19040), .ZN(n16295) );
  NAND2_X1 U16066 ( .A1(n16295), .A2(n13520), .ZN(n13067) );
  OAI211_X1 U16067 ( .C1(n13520), .C2(n10567), .A(n13068), .B(n13067), .ZN(
        P2_U2879) );
  AOI21_X1 U16068 ( .B1(n13069), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13071) );
  OR3_X1 U16069 ( .A1(n13071), .A2(n13070), .A3(n14865), .ZN(n13075) );
  OAI21_X1 U16070 ( .B1(n13073), .B2(n13072), .A(n13063), .ZN(n15183) );
  INV_X1 U16071 ( .A(n15183), .ZN(n19047) );
  NAND2_X1 U16072 ( .A1(n19047), .A2(n13520), .ZN(n13074) );
  OAI211_X1 U16073 ( .C1(n13520), .C2(n13076), .A(n13075), .B(n13074), .ZN(
        P2_U2880) );
  AOI22_X1 U16074 ( .A1(n20101), .A2(P1_EAX_REG_21__SCAN_IN), .B1(
        P1_UWORD_REG_5__SCAN_IN), .B2(n20100), .ZN(n13079) );
  NAND2_X1 U16075 ( .A1(n13079), .A2(n13078), .ZN(P1_U2942) );
  AOI22_X1 U16076 ( .A1(n20101), .A2(P1_EAX_REG_23__SCAN_IN), .B1(
        P1_UWORD_REG_7__SCAN_IN), .B2(n20100), .ZN(n13081) );
  NAND2_X1 U16077 ( .A1(n13081), .A2(n13080), .ZN(P1_U2944) );
  AOI22_X1 U16078 ( .A1(n20101), .A2(P1_EAX_REG_19__SCAN_IN), .B1(
        P1_UWORD_REG_3__SCAN_IN), .B2(n20100), .ZN(n13083) );
  NAND2_X1 U16079 ( .A1(n13083), .A2(n13082), .ZN(P1_U2940) );
  AOI22_X1 U16080 ( .A1(n20101), .A2(P1_EAX_REG_22__SCAN_IN), .B1(
        P1_UWORD_REG_6__SCAN_IN), .B2(n20100), .ZN(n13085) );
  NAND2_X1 U16081 ( .A1(n13085), .A2(n13084), .ZN(P1_U2943) );
  AOI22_X1 U16082 ( .A1(n20101), .A2(P1_EAX_REG_27__SCAN_IN), .B1(
        P1_UWORD_REG_11__SCAN_IN), .B2(n20100), .ZN(n13087) );
  NAND2_X1 U16083 ( .A1(n13087), .A2(n13086), .ZN(P1_U2948) );
  AOI22_X1 U16084 ( .A1(n20101), .A2(P1_EAX_REG_20__SCAN_IN), .B1(
        P1_UWORD_REG_4__SCAN_IN), .B2(n20100), .ZN(n13089) );
  NAND2_X1 U16085 ( .A1(n13089), .A2(n13088), .ZN(P1_U2941) );
  AOI22_X1 U16086 ( .A1(n20101), .A2(P1_EAX_REG_16__SCAN_IN), .B1(
        P1_UWORD_REG_0__SCAN_IN), .B2(n20100), .ZN(n13093) );
  NAND2_X1 U16087 ( .A1(n13861), .A2(DATAI_0_), .ZN(n13091) );
  NAND2_X1 U16088 ( .A1(n14410), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13090) );
  AND2_X1 U16089 ( .A1(n13091), .A2(n13090), .ZN(n13859) );
  INV_X1 U16090 ( .A(n13859), .ZN(n13092) );
  NAND2_X1 U16091 ( .A1(n20088), .A2(n13092), .ZN(n13097) );
  NAND2_X1 U16092 ( .A1(n13093), .A2(n13097), .ZN(P1_U2937) );
  AOI22_X1 U16093 ( .A1(n20101), .A2(P1_EAX_REG_18__SCAN_IN), .B1(
        P1_UWORD_REG_2__SCAN_IN), .B2(n20100), .ZN(n13096) );
  NAND2_X1 U16094 ( .A1(n13861), .A2(DATAI_2_), .ZN(n13095) );
  NAND2_X1 U16095 ( .A1(n14410), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13094) );
  AND2_X1 U16096 ( .A1(n13095), .A2(n13094), .ZN(n13351) );
  INV_X1 U16097 ( .A(n13351), .ZN(n14463) );
  NAND2_X1 U16098 ( .A1(n20088), .A2(n14463), .ZN(n13103) );
  NAND2_X1 U16099 ( .A1(n13096), .A2(n13103), .ZN(P1_U2939) );
  AOI22_X1 U16100 ( .A1(n20101), .A2(P1_EAX_REG_0__SCAN_IN), .B1(
        P1_LWORD_REG_0__SCAN_IN), .B2(n20100), .ZN(n13098) );
  NAND2_X1 U16101 ( .A1(n13098), .A2(n13097), .ZN(P1_U2952) );
  AOI22_X1 U16102 ( .A1(n20101), .A2(P1_EAX_REG_17__SCAN_IN), .B1(
        P1_UWORD_REG_1__SCAN_IN), .B2(n20100), .ZN(n13102) );
  NAND2_X1 U16103 ( .A1(n13861), .A2(DATAI_1_), .ZN(n13100) );
  NAND2_X1 U16104 ( .A1(n14410), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13099) );
  AND2_X1 U16105 ( .A1(n13100), .A2(n13099), .ZN(n13871) );
  INV_X1 U16106 ( .A(n13871), .ZN(n13101) );
  NAND2_X1 U16107 ( .A1(n20088), .A2(n13101), .ZN(n13105) );
  NAND2_X1 U16108 ( .A1(n13102), .A2(n13105), .ZN(P1_U2938) );
  AOI22_X1 U16109 ( .A1(n20101), .A2(P1_EAX_REG_2__SCAN_IN), .B1(
        P1_LWORD_REG_2__SCAN_IN), .B2(n20100), .ZN(n13104) );
  NAND2_X1 U16110 ( .A1(n13104), .A2(n13103), .ZN(P1_U2954) );
  AOI22_X1 U16111 ( .A1(n20101), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_LWORD_REG_1__SCAN_IN), .B2(n20100), .ZN(n13106) );
  NAND2_X1 U16112 ( .A1(n13106), .A2(n13105), .ZN(P1_U2953) );
  XNOR2_X1 U16113 ( .A(n13108), .B(n13107), .ZN(n13657) );
  INV_X1 U16114 ( .A(n13109), .ZN(n13112) );
  INV_X1 U16115 ( .A(n13110), .ZN(n13111) );
  AOI21_X1 U16116 ( .B1(n13112), .B2(n20153), .A(n13111), .ZN(n14723) );
  INV_X1 U16117 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n13113) );
  NOR2_X1 U16118 ( .A1(n20135), .A2(n13113), .ZN(n14724) );
  INV_X1 U16119 ( .A(n20120), .ZN(n14580) );
  INV_X1 U16120 ( .A(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13114) );
  AOI21_X1 U16121 ( .B1(n14580), .B2(n13115), .A(n13114), .ZN(n13116) );
  AOI211_X1 U16122 ( .C1(n14723), .C2(n12697), .A(n14724), .B(n13116), .ZN(
        n13117) );
  OAI21_X1 U16123 ( .B1(n13657), .B2(n14616), .A(n13117), .ZN(P1_U2999) );
  NAND4_X1 U16124 ( .A1(n9773), .A2(n13743), .A3(n14201), .A4(n13340), .ZN(
        n13401) );
  OR2_X1 U16125 ( .A1(n13165), .A2(n13401), .ZN(n13119) );
  AND2_X1 U16126 ( .A1(n11839), .A2(n14192), .ZN(n13123) );
  INV_X1 U16127 ( .A(n13123), .ZN(n13121) );
  AND2_X1 U16128 ( .A1(n13121), .A2(n11843), .ZN(n13122) );
  INV_X1 U16129 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n20068) );
  OAI222_X1 U16130 ( .A1(n14476), .A2(n13657), .B1(n14179), .B2(n20068), .C1(
        n14475), .C2(n13859), .ZN(P1_U2904) );
  XOR2_X1 U16131 ( .A(n13124), .B(n13125), .Z(n20126) );
  INV_X1 U16132 ( .A(n20126), .ZN(n13694) );
  INV_X1 U16133 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n20061) );
  OAI222_X1 U16134 ( .A1(n13694), .A2(n14476), .B1(n13351), .B2(n14475), .C1(
        n14473), .C2(n20061), .ZN(P1_U2902) );
  OAI21_X1 U16135 ( .B1(n13127), .B2(n13126), .A(n13124), .ZN(n20027) );
  INV_X1 U16136 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n20063) );
  OAI222_X1 U16137 ( .A1(n20027), .A2(n14476), .B1(n13871), .B2(n14475), .C1(
        n14473), .C2(n20063), .ZN(P1_U2903) );
  INV_X1 U16138 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13129) );
  AOI22_X1 U16139 ( .A1(P1_UWORD_REG_5__SCAN_IN), .A2(n20768), .B1(n20064), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13128) );
  OAI21_X1 U16140 ( .B1(n13129), .B2(n13141), .A(n13128), .ZN(P1_U2915) );
  INV_X1 U16141 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n14437) );
  AOI22_X1 U16142 ( .A1(P1_UWORD_REG_7__SCAN_IN), .A2(n20768), .B1(n20064), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13130) );
  OAI21_X1 U16143 ( .B1(n14437), .B2(n13141), .A(n13130), .ZN(P1_U2913) );
  INV_X1 U16144 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13132) );
  AOI22_X1 U16145 ( .A1(P1_UWORD_REG_6__SCAN_IN), .A2(n20768), .B1(n20064), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13131) );
  OAI21_X1 U16146 ( .B1(n13132), .B2(n13141), .A(n13131), .ZN(P1_U2914) );
  AOI22_X1 U16147 ( .A1(P1_UWORD_REG_3__SCAN_IN), .A2(n20768), .B1(n20064), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13133) );
  OAI21_X1 U16148 ( .B1(n14455), .B2(n13141), .A(n13133), .ZN(P1_U2917) );
  INV_X1 U16149 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n13135) );
  AOI22_X1 U16150 ( .A1(P1_UWORD_REG_0__SCAN_IN), .A2(n20065), .B1(n20064), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13134) );
  OAI21_X1 U16151 ( .B1(n13135), .B2(n13141), .A(n13134), .ZN(P1_U2920) );
  INV_X1 U16152 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13137) );
  AOI22_X1 U16153 ( .A1(P1_UWORD_REG_4__SCAN_IN), .A2(n20768), .B1(n20064), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13136) );
  OAI21_X1 U16154 ( .B1(n13137), .B2(n13141), .A(n13136), .ZN(P1_U2916) );
  INV_X1 U16155 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13139) );
  AOI22_X1 U16156 ( .A1(P1_UWORD_REG_2__SCAN_IN), .A2(n20065), .B1(n20064), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13138) );
  OAI21_X1 U16157 ( .B1(n13139), .B2(n13141), .A(n13138), .ZN(P1_U2918) );
  INV_X1 U16158 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n20901) );
  AOI22_X1 U16159 ( .A1(P1_UWORD_REG_1__SCAN_IN), .A2(n20065), .B1(n20064), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13140) );
  OAI21_X1 U16160 ( .B1(n20901), .B2(n13141), .A(n13140), .ZN(P1_U2919) );
  AND2_X1 U16161 ( .A1(n13143), .A2(n13142), .ZN(n13145) );
  OR2_X1 U16162 ( .A1(n13145), .A2(n13144), .ZN(n15424) );
  INV_X1 U16163 ( .A(n15424), .ZN(n19016) );
  NAND2_X1 U16164 ( .A1(n19016), .A2(n13520), .ZN(n13149) );
  OAI211_X1 U16165 ( .C1(n10039), .C2(n13147), .A(n14844), .B(n13146), .ZN(
        n13148) );
  OAI211_X1 U16166 ( .C1(n13520), .C2(n10598), .A(n13149), .B(n13148), .ZN(
        P2_U2877) );
  OR2_X1 U16167 ( .A1(n13144), .A2(n13150), .ZN(n13151) );
  AND2_X1 U16168 ( .A1(n13151), .A2(n13226), .ZN(n19002) );
  INV_X1 U16169 ( .A(n19002), .ZN(n15412) );
  INV_X1 U16170 ( .A(n13146), .ZN(n13154) );
  OAI211_X1 U16171 ( .C1(n13154), .C2(n13153), .A(n14844), .B(n13220), .ZN(
        n13156) );
  NAND2_X1 U16172 ( .A1(n14856), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n13155) );
  OAI211_X1 U16173 ( .C1(n15412), .C2(n14856), .A(n13156), .B(n13155), .ZN(
        P2_U2876) );
  OAI21_X1 U16174 ( .B1(n13158), .B2(n13157), .A(n13216), .ZN(n18999) );
  OAI222_X1 U16175 ( .A1(n19152), .A2(n12759), .B1(n13159), .B2(n19169), .C1(
        n18999), .C2(n19143), .ZN(P2_U2908) );
  NAND2_X1 U16176 ( .A1(n13161), .A2(n13160), .ZN(n13233) );
  OR2_X1 U16177 ( .A1(n13161), .A2(n13160), .ZN(n13162) );
  AND2_X1 U16178 ( .A1(n13233), .A2(n13162), .ZN(n20116) );
  INV_X1 U16179 ( .A(n20116), .ZN(n13532) );
  INV_X1 U16180 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n20059) );
  OAI222_X1 U16181 ( .A1(n13532), .A2(n14476), .B1(n14456), .B2(n14475), .C1(
        n14473), .C2(n20059), .ZN(P1_U2901) );
  INV_X1 U16182 ( .A(n13164), .ZN(n13166) );
  NAND2_X1 U16183 ( .A1(n13166), .A2(n13165), .ZN(n13167) );
  NOR2_X1 U16184 ( .A1(n12929), .A2(n13167), .ZN(n13168) );
  AND2_X1 U16185 ( .A1(n12928), .A2(n13168), .ZN(n13177) );
  NAND2_X1 U16186 ( .A1(n12538), .A2(n13191), .ZN(n13174) );
  INV_X1 U16187 ( .A(n13360), .ZN(n13170) );
  NAND2_X1 U16188 ( .A1(n13170), .A2(n11848), .ZN(n13427) );
  NAND2_X1 U16189 ( .A1(n14163), .A2(n13171), .ZN(n13172) );
  OAI21_X1 U16190 ( .B1(n9775), .B2(n13637), .A(n13172), .ZN(n13173) );
  AOI21_X1 U16191 ( .B1(n13174), .B2(n13734), .A(n13173), .ZN(n13176) );
  AND3_X1 U16192 ( .A1(n11864), .A2(n13176), .A3(n13175), .ZN(n13751) );
  NAND2_X1 U16193 ( .A1(n13177), .A2(n13751), .ZN(n14102) );
  AND2_X1 U16194 ( .A1(n14191), .A2(n13178), .ZN(n13194) );
  NOR2_X1 U16195 ( .A1(n14745), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13188) );
  XNOR2_X1 U16196 ( .A(n13188), .B(n13198), .ZN(n13185) );
  NAND2_X1 U16197 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13180) );
  AOI22_X1 U16198 ( .A1(n13181), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B1(
        n13198), .B2(n13180), .ZN(n13183) );
  NAND2_X1 U16199 ( .A1(n14745), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13189) );
  AOI21_X1 U16200 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13189), .A(
        n9646), .ZN(n20745) );
  NOR3_X1 U16201 ( .A1(n14102), .A2(n20745), .A3(n13191), .ZN(n13182) );
  AOI21_X1 U16202 ( .B1(n15762), .B2(n13183), .A(n13182), .ZN(n13184) );
  OAI21_X1 U16203 ( .B1(n13194), .B2(n13185), .A(n13184), .ZN(n13186) );
  AOI21_X1 U16204 ( .B1(n20371), .B2(n14102), .A(n13186), .ZN(n20747) );
  MUX2_X1 U16205 ( .A(n13198), .B(n20747), .S(n15759), .Z(n15775) );
  INV_X1 U16206 ( .A(n15775), .ZN(n15777) );
  INV_X1 U16207 ( .A(n14102), .ZN(n14738) );
  XNOR2_X1 U16208 ( .A(n20903), .B(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n13193) );
  INV_X1 U16209 ( .A(n13188), .ZN(n13190) );
  NAND2_X1 U16210 ( .A1(n13190), .A2(n13189), .ZN(n14755) );
  NOR3_X1 U16211 ( .A1(n14102), .A2(n13191), .A3(n14755), .ZN(n13192) );
  AOI21_X1 U16212 ( .B1(n15762), .B2(n13193), .A(n13192), .ZN(n13197) );
  INV_X1 U16213 ( .A(n13194), .ZN(n13195) );
  NAND2_X1 U16214 ( .A1(n13195), .A2(n14755), .ZN(n13196) );
  OAI211_X1 U16215 ( .C1(n13187), .C2(n14738), .A(n13197), .B(n13196), .ZN(
        n14751) );
  MUX2_X1 U16216 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14751), .S(
        n15759), .Z(n15771) );
  NAND2_X1 U16217 ( .A1(n15771), .A2(n20669), .ZN(n13200) );
  NOR2_X1 U16218 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n20669), .ZN(n13205) );
  NAND3_X1 U16219 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13205), .A3(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13199) );
  OAI21_X1 U16220 ( .B1(n15775), .B2(n13200), .A(n13199), .ZN(n15784) );
  INV_X1 U16221 ( .A(n13202), .ZN(n13203) );
  NAND2_X1 U16222 ( .A1(n15784), .A2(n13203), .ZN(n14734) );
  OAI21_X1 U16223 ( .B1(n19998), .B2(n12928), .A(n15759), .ZN(n13207) );
  INV_X1 U16224 ( .A(n15759), .ZN(n13204) );
  AOI21_X1 U16225 ( .B1(n13204), .B2(n12027), .A(P1_STATE2_REG_1__SCAN_IN), 
        .ZN(n13206) );
  AOI22_X1 U16226 ( .A1(n13207), .A2(n13206), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n13205), .ZN(n15786) );
  AND3_X1 U16227 ( .A1(n14734), .A2(n19919), .A3(n15786), .ZN(n13208) );
  NOR2_X1 U16228 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n15800) );
  OAI21_X1 U16229 ( .B1(n13208), .B2(n16114), .A(n13359), .ZN(n20170) );
  NAND2_X1 U16230 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20379), .ZN(n14735) );
  INV_X1 U16231 ( .A(n14735), .ZN(n13212) );
  AND2_X1 U16232 ( .A1(n9655), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n13439) );
  NOR2_X1 U16233 ( .A1(n13439), .A2(n20556), .ZN(n20558) );
  OAI21_X1 U16234 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n9655), .A(n20558), 
        .ZN(n13211) );
  OAI21_X1 U16235 ( .B1(n13212), .B2(n20372), .A(n13211), .ZN(n13213) );
  NAND2_X1 U16236 ( .A1(n20170), .A2(n13213), .ZN(n13214) );
  OAI21_X1 U16237 ( .B1(n20170), .B2(n15765), .A(n13214), .ZN(P1_U3477) );
  AOI21_X1 U16238 ( .B1(n13217), .B2(n13216), .A(n13215), .ZN(n18992) );
  INV_X1 U16239 ( .A(n18992), .ZN(n13219) );
  INV_X1 U16240 ( .A(n14879), .ZN(n13218) );
  OAI222_X1 U16241 ( .A1(n13219), .A2(n19143), .B1(n13218), .B2(n19169), .C1(
        n12901), .C2(n19152), .ZN(P2_U2907) );
  INV_X1 U16242 ( .A(P2_EBX_REG_12__SCAN_IN), .ZN(n13230) );
  INV_X1 U16243 ( .A(n13222), .ZN(n13223) );
  OAI211_X1 U16244 ( .C1(n13152), .C2(n13224), .A(n13223), .B(n14844), .ZN(
        n13229) );
  NAND2_X1 U16245 ( .A1(n13226), .A2(n13225), .ZN(n13227) );
  AND2_X1 U16246 ( .A1(n9708), .A2(n13227), .ZN(n18993) );
  INV_X1 U16247 ( .A(n14856), .ZN(n13520) );
  NAND2_X1 U16248 ( .A1(n18993), .A2(n13520), .ZN(n13228) );
  OAI211_X1 U16249 ( .C1(n13520), .C2(n13230), .A(n13229), .B(n13228), .ZN(
        P2_U2875) );
  NAND2_X1 U16250 ( .A1(n13233), .A2(n13232), .ZN(n13234) );
  AND2_X1 U16251 ( .A1(n13231), .A2(n13234), .ZN(n20108) );
  INV_X1 U16252 ( .A(n20108), .ZN(n13580) );
  INV_X1 U16253 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n20057) );
  OAI222_X1 U16254 ( .A1(n13580), .A2(n14476), .B1(n14451), .B2(n14475), .C1(
        n14473), .C2(n20057), .ZN(P1_U2900) );
  INV_X1 U16255 ( .A(n20170), .ZN(n13246) );
  INV_X1 U16256 ( .A(n13187), .ZN(n20177) );
  AND2_X1 U16257 ( .A1(n13439), .A2(n20585), .ZN(n20473) );
  MUX2_X1 U16258 ( .A(n20558), .B(n20473), .S(n13235), .Z(n13236) );
  AOI21_X1 U16259 ( .B1(n14735), .B2(n20177), .A(n13236), .ZN(n13238) );
  NAND2_X1 U16260 ( .A1(n13246), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n13237) );
  OAI21_X1 U16261 ( .B1(n13246), .B2(n13238), .A(n13237), .ZN(P1_U3476) );
  MUX2_X1 U16262 ( .A(n20559), .B(n20311), .S(n9655), .Z(n13241) );
  INV_X1 U16263 ( .A(n13235), .ZN(n13240) );
  NAND3_X1 U16264 ( .A1(n13241), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(n20467), 
        .ZN(n13242) );
  NAND2_X1 U16265 ( .A1(n13242), .A2(n20585), .ZN(n20343) );
  AOI21_X1 U16266 ( .B1(n20171), .B2(n20761), .A(n20343), .ZN(n13243) );
  AOI21_X1 U16267 ( .B1(n14735), .B2(n20371), .A(n13243), .ZN(n13245) );
  NAND2_X1 U16268 ( .A1(n13246), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13244) );
  OAI21_X1 U16269 ( .B1(n13246), .B2(n13245), .A(n13244), .ZN(P1_U3475) );
  OAI21_X1 U16270 ( .B1(n13215), .B2(n13247), .A(n15365), .ZN(n18986) );
  OAI222_X1 U16271 ( .A1(n18986), .A2(n19143), .B1(n13248), .B2(n19169), .C1(
        n12908), .C2(n19152), .ZN(P2_U2906) );
  AND2_X1 U16272 ( .A1(n13288), .A2(n19896), .ZN(n13597) );
  INV_X1 U16273 ( .A(n13597), .ZN(n13249) );
  NOR2_X1 U16274 ( .A1(n13250), .A2(n13249), .ZN(n13604) );
  AND2_X1 U16275 ( .A1(n13251), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19894) );
  INV_X1 U16276 ( .A(n19894), .ZN(n13325) );
  INV_X1 U16277 ( .A(n13252), .ZN(n13307) );
  INV_X1 U16278 ( .A(n13284), .ZN(n13253) );
  NAND2_X1 U16279 ( .A1(n13254), .A2(n13253), .ZN(n13271) );
  NOR2_X1 U16280 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13256) );
  OR2_X1 U16281 ( .A1(n13255), .A2(n13256), .ZN(n13258) );
  INV_X1 U16282 ( .A(n13258), .ZN(n13270) );
  AOI22_X1 U16283 ( .A1(n13271), .A2(n13270), .B1(n13257), .B2(n13304), .ZN(
        n13265) );
  INV_X1 U16284 ( .A(n13304), .ZN(n13262) );
  NAND2_X1 U16285 ( .A1(n13271), .A2(n13258), .ZN(n13261) );
  NAND2_X1 U16286 ( .A1(n13259), .A2(n11192), .ZN(n13274) );
  NAND2_X1 U16287 ( .A1(n13274), .A2(n11490), .ZN(n13260) );
  OAI211_X1 U16288 ( .C1(n13257), .C2(n13262), .A(n13261), .B(n13260), .ZN(
        n13263) );
  INV_X1 U16289 ( .A(n13263), .ZN(n13264) );
  MUX2_X1 U16290 ( .A(n13265), .B(n13264), .S(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13267) );
  NAND2_X1 U16291 ( .A1(n13267), .A2(n13266), .ZN(n13268) );
  AOI21_X1 U16292 ( .B1(n10285), .B2(n13307), .A(n13268), .ZN(n15497) );
  MUX2_X1 U16293 ( .A(n13269), .B(n15497), .S(n13308), .Z(n13314) );
  INV_X1 U16294 ( .A(n13314), .ZN(n13323) );
  NAND2_X1 U16295 ( .A1(n13270), .A2(n11490), .ZN(n13272) );
  NAND2_X1 U16296 ( .A1(n13271), .A2(n13272), .ZN(n13278) );
  INV_X1 U16297 ( .A(n13272), .ZN(n13273) );
  NAND2_X1 U16298 ( .A1(n13274), .A2(n13273), .ZN(n13277) );
  NOR2_X1 U16299 ( .A1(n13255), .A2(n13257), .ZN(n13275) );
  NAND2_X1 U16300 ( .A1(n13304), .A2(n13275), .ZN(n13276) );
  NAND3_X1 U16301 ( .A1(n13278), .A2(n13277), .A3(n13276), .ZN(n13279) );
  AOI21_X1 U16302 ( .B1(n9657), .B2(n13307), .A(n13279), .ZN(n15493) );
  MUX2_X1 U16303 ( .A(n13280), .B(n15493), .S(n13308), .Z(n13316) );
  INV_X1 U16304 ( .A(n13316), .ZN(n13322) );
  AOI22_X1 U16305 ( .A1(n15479), .A2(n13283), .B1(n13282), .B2(n13281), .ZN(
        n13287) );
  NAND2_X1 U16306 ( .A1(n13285), .A2(n13284), .ZN(n13286) );
  AND2_X1 U16307 ( .A1(n13287), .A2(n13286), .ZN(n19887) );
  INV_X1 U16308 ( .A(n13288), .ZN(n13289) );
  NAND2_X1 U16309 ( .A1(n13290), .A2(n13289), .ZN(n13291) );
  NOR2_X1 U16310 ( .A1(n13292), .A2(n13291), .ZN(n18858) );
  INV_X1 U16311 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n13293) );
  NAND2_X1 U16312 ( .A1(n18860), .A2(n13293), .ZN(n13296) );
  OAI22_X1 U16313 ( .A1(n15507), .A2(n10745), .B1(n13294), .B2(n12801), .ZN(
        n13295) );
  AOI21_X1 U16314 ( .B1(n18858), .B2(n13296), .A(n13295), .ZN(n13297) );
  OAI211_X1 U16315 ( .C1(n13308), .C2(n20796), .A(n19887), .B(n13297), .ZN(
        n13321) );
  NAND2_X1 U16316 ( .A1(n15497), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n13313) );
  NAND2_X1 U16317 ( .A1(n13304), .A2(n10069), .ZN(n13302) );
  NAND2_X1 U16318 ( .A1(n13299), .A2(n13298), .ZN(n13305) );
  OAI21_X1 U16319 ( .B1(n13300), .B2(n10297), .A(n13305), .ZN(n13301) );
  NAND2_X1 U16320 ( .A1(n13302), .A2(n13301), .ZN(n13303) );
  AOI21_X1 U16321 ( .B1(n11297), .B2(n13307), .A(n13303), .ZN(n15490) );
  MUX2_X1 U16322 ( .A(n13305), .B(n13304), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n13306) );
  AOI21_X1 U16323 ( .B1(n16315), .B2(n13307), .A(n13306), .ZN(n15482) );
  OAI211_X1 U16324 ( .C1(n15490), .C2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n15482), .ZN(n13311) );
  INV_X1 U16325 ( .A(n13308), .ZN(n13309) );
  AOI21_X1 U16326 ( .B1(n15490), .B2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A(
        n13309), .ZN(n13310) );
  AND2_X1 U16327 ( .A1(n13311), .A2(n13310), .ZN(n13312) );
  AND2_X1 U16328 ( .A1(n13313), .A2(n13312), .ZN(n13318) );
  INV_X1 U16329 ( .A(n13318), .ZN(n13315) );
  OAI221_X1 U16330 ( .B1(n13316), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), 
        .C1(n13316), .C2(n13315), .A(n13314), .ZN(n13317) );
  AOI22_X1 U16331 ( .A1(n13318), .A2(n19863), .B1(n19856), .B2(n13317), .ZN(
        n13319) );
  NOR2_X1 U16332 ( .A1(n13319), .A2(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(
        n13320) );
  AOI211_X1 U16333 ( .C1(n13323), .C2(n13322), .A(n13321), .B(n13320), .ZN(
        n16330) );
  AOI21_X1 U16334 ( .B1(n16330), .B2(n15828), .A(n18853), .ZN(n13324) );
  AOI211_X1 U16335 ( .C1(n13326), .C2(n13604), .A(n13325), .B(n13324), .ZN(
        n16325) );
  OAI21_X1 U16336 ( .B1(n16325), .B2(n18853), .A(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n13327) );
  NAND2_X1 U16337 ( .A1(n13327), .A2(n15829), .ZN(P2_U3593) );
  AND2_X1 U16338 ( .A1(n20311), .A2(n20585), .ZN(n20345) );
  OR2_X1 U16339 ( .A1(n13187), .A2(n13328), .ZN(n20318) );
  INV_X1 U16340 ( .A(n20318), .ZN(n20341) );
  AND2_X1 U16341 ( .A1(n11920), .A2(n11934), .ZN(n20469) );
  INV_X1 U16342 ( .A(n13329), .ZN(n13362) );
  AOI21_X1 U16343 ( .B1(n20341), .B2(n20469), .A(n13362), .ZN(n13332) );
  OAI21_X1 U16344 ( .B1(n20345), .B2(n20558), .A(n13332), .ZN(n13330) );
  OAI211_X1 U16345 ( .C1(n20585), .C2(n11982), .A(n20561), .B(n13330), .ZN(
        n13331) );
  INV_X1 U16346 ( .A(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13336) );
  NOR2_X2 U16347 ( .A1(n13871), .A2(n13359), .ZN(n20606) );
  OAI22_X1 U16348 ( .A1(n13332), .A2(n20556), .B1(n13473), .B2(n20760), .ZN(
        n13363) );
  NAND2_X1 U16349 ( .A1(n13361), .A2(n13734), .ZN(n20516) );
  AOI22_X1 U16350 ( .A1(n20606), .A2(n13363), .B1(n13362), .B2(n20605), .ZN(
        n13335) );
  NAND2_X1 U16351 ( .A1(n9655), .A2(n12612), .ZN(n20429) );
  NOR2_X2 U16352 ( .A1(n14616), .A2(n13861), .ZN(n13364) );
  NOR2_X2 U16353 ( .A1(n14410), .A2(n14616), .ZN(n13365) );
  AOI22_X1 U16354 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n13364), .B1(DATAI_25_), 
        .B2(n13365), .ZN(n20520) );
  INV_X1 U16355 ( .A(n20520), .ZN(n20607) );
  NAND2_X1 U16356 ( .A1(n9655), .A2(n20172), .ZN(n20466) );
  NOR2_X2 U16357 ( .A1(n20311), .A2(n20466), .ZN(n20396) );
  INV_X1 U16358 ( .A(n20610), .ZN(n20479) );
  AOI22_X1 U16359 ( .A1(n13366), .A2(n20607), .B1(n20396), .B2(n20479), .ZN(
        n13334) );
  OAI211_X1 U16360 ( .C1(n13370), .C2(n13336), .A(n13335), .B(n13334), .ZN(
        P1_U3090) );
  INV_X1 U16361 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13339) );
  NOR2_X2 U16362 ( .A1(n13859), .A2(n13359), .ZN(n20592) );
  NAND2_X1 U16363 ( .A1(n13361), .A2(n11848), .ZN(n20503) );
  AOI22_X1 U16364 ( .A1(n20592), .A2(n13363), .B1(n13362), .B2(n20591), .ZN(
        n13338) );
  AOI22_X1 U16365 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n13364), .B1(DATAI_24_), 
        .B2(n13365), .ZN(n20515) );
  INV_X1 U16366 ( .A(n20515), .ZN(n20601) );
  INV_X1 U16367 ( .A(n20604), .ZN(n20404) );
  AOI22_X1 U16368 ( .A1(n13366), .A2(n20601), .B1(n20396), .B2(n20404), .ZN(
        n13337) );
  OAI211_X1 U16369 ( .C1(n13370), .C2(n13339), .A(n13338), .B(n13337), .ZN(
        P1_U3089) );
  INV_X1 U16370 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13343) );
  NOR2_X2 U16371 ( .A1(n14442), .A2(n13359), .ZN(n20632) );
  NAND2_X1 U16372 ( .A1(n13361), .A2(n13340), .ZN(n20539) );
  AOI22_X1 U16373 ( .A1(n20632), .A2(n13363), .B1(n13362), .B2(n20631), .ZN(
        n13342) );
  AOI22_X1 U16374 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n13364), .B1(DATAI_30_), 
        .B2(n13365), .ZN(n20543) );
  INV_X1 U16375 ( .A(n20543), .ZN(n20633) );
  INV_X1 U16376 ( .A(n20636), .ZN(n20419) );
  AOI22_X1 U16377 ( .A1(n13366), .A2(n20633), .B1(n20396), .B2(n20419), .ZN(
        n13341) );
  OAI211_X1 U16378 ( .C1(n13370), .C2(n13343), .A(n13342), .B(n13341), .ZN(
        P1_U3095) );
  INV_X1 U16379 ( .A(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13347) );
  NOR2_X2 U16380 ( .A1(n14447), .A2(n13359), .ZN(n20626) );
  NAND2_X1 U16381 ( .A1(n13361), .A2(n13344), .ZN(n20534) );
  AOI22_X1 U16382 ( .A1(n20626), .A2(n13363), .B1(n13362), .B2(n20625), .ZN(
        n13346) );
  AOI22_X1 U16383 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n13364), .B1(DATAI_29_), 
        .B2(n13365), .ZN(n20538) );
  INV_X1 U16384 ( .A(n20538), .ZN(n20627) );
  INV_X1 U16385 ( .A(n20630), .ZN(n20416) );
  AOI22_X1 U16386 ( .A1(n13366), .A2(n20627), .B1(n20396), .B2(n20416), .ZN(
        n13345) );
  OAI211_X1 U16387 ( .C1(n13370), .C2(n13347), .A(n13346), .B(n13345), .ZN(
        P1_U3094) );
  INV_X1 U16388 ( .A(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13350) );
  NOR2_X2 U16389 ( .A1(n14438), .A2(n13359), .ZN(n20661) );
  NAND2_X1 U16390 ( .A1(n13361), .A2(n14192), .ZN(n20545) );
  AOI22_X1 U16391 ( .A1(n20661), .A2(n13363), .B1(n13362), .B2(n20658), .ZN(
        n13349) );
  AOI22_X1 U16392 ( .A1(BUF1_REG_31__SCAN_IN), .A2(n13364), .B1(DATAI_31_), 
        .B2(n13365), .ZN(n20668) );
  INV_X1 U16393 ( .A(n20668), .ZN(n20639) );
  INV_X1 U16394 ( .A(n20644), .ZN(n20662) );
  AOI22_X1 U16395 ( .A1(n13366), .A2(n20639), .B1(n20396), .B2(n20662), .ZN(
        n13348) );
  OAI211_X1 U16396 ( .C1(n13370), .C2(n13350), .A(n13349), .B(n13348), .ZN(
        P1_U3096) );
  INV_X1 U16397 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13355) );
  NOR2_X2 U16398 ( .A1(n13351), .A2(n13359), .ZN(n20647) );
  NAND2_X1 U16399 ( .A1(n13361), .A2(n13352), .ZN(n20521) );
  AOI22_X1 U16400 ( .A1(n20647), .A2(n13363), .B1(n13362), .B2(n20646), .ZN(
        n13354) );
  AOI22_X1 U16401 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n13364), .B1(DATAI_26_), 
        .B2(n13365), .ZN(n20651) );
  INV_X1 U16402 ( .A(n20651), .ZN(n20611) );
  AOI22_X1 U16403 ( .A1(DATAI_18_), .A2(n13365), .B1(BUF1_REG_18__SCAN_IN), 
        .B2(n13364), .ZN(n20614) );
  INV_X1 U16404 ( .A(n20614), .ZN(n20648) );
  AOI22_X1 U16405 ( .A1(n13366), .A2(n20611), .B1(n20396), .B2(n20648), .ZN(
        n13353) );
  OAI211_X1 U16406 ( .C1(n13370), .C2(n13355), .A(n13354), .B(n13353), .ZN(
        P1_U3091) );
  INV_X1 U16407 ( .A(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13358) );
  NOR2_X2 U16408 ( .A1(n14451), .A2(n13359), .ZN(n20653) );
  NAND2_X1 U16409 ( .A1(n13361), .A2(n13759), .ZN(n20530) );
  AOI22_X1 U16410 ( .A1(n20653), .A2(n13363), .B1(n13362), .B2(n20652), .ZN(
        n13357) );
  AOI22_X1 U16411 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n13364), .B1(DATAI_28_), 
        .B2(n13365), .ZN(n20657) );
  INV_X1 U16412 ( .A(n20657), .ZN(n20621) );
  INV_X1 U16413 ( .A(n20624), .ZN(n20654) );
  AOI22_X1 U16414 ( .A1(n13366), .A2(n20621), .B1(n20396), .B2(n20654), .ZN(
        n13356) );
  OAI211_X1 U16415 ( .C1(n13370), .C2(n13358), .A(n13357), .B(n13356), .ZN(
        P1_U3093) );
  INV_X1 U16416 ( .A(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13369) );
  NOR2_X2 U16417 ( .A1(n14456), .A2(n13359), .ZN(n20616) );
  NAND2_X1 U16418 ( .A1(n13361), .A2(n13360), .ZN(n20525) );
  AOI22_X1 U16419 ( .A1(n20616), .A2(n13363), .B1(n13362), .B2(n20615), .ZN(
        n13368) );
  AOI22_X1 U16420 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n13364), .B1(DATAI_27_), 
        .B2(n13365), .ZN(n20529) );
  INV_X1 U16421 ( .A(n20529), .ZN(n20617) );
  INV_X1 U16422 ( .A(n20620), .ZN(n20411) );
  AOI22_X1 U16423 ( .A1(n13366), .A2(n20617), .B1(n20396), .B2(n20411), .ZN(
        n13367) );
  OAI211_X1 U16424 ( .C1(n13370), .C2(n13369), .A(n13368), .B(n13367), .ZN(
        P1_U3092) );
  INV_X1 U16425 ( .A(n13371), .ZN(n13372) );
  XNOR2_X1 U16426 ( .A(n13231), .B(n13372), .ZN(n19993) );
  INV_X1 U16427 ( .A(n19993), .ZN(n13537) );
  OAI222_X1 U16428 ( .A1(n14476), .A2(n13537), .B1(n14179), .B2(n12055), .C1(
        n14475), .C2(n14447), .ZN(P1_U2899) );
  AND2_X1 U16429 ( .A1(n13374), .A2(n13376), .ZN(n19979) );
  INV_X1 U16430 ( .A(n19979), .ZN(n13438) );
  INV_X1 U16431 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n13377) );
  OAI222_X1 U16432 ( .A1(n13438), .A2(n14476), .B1(n14442), .B2(n14475), .C1(
        n13377), .C2(n14179), .ZN(P1_U2898) );
  XNOR2_X1 U16433 ( .A(n13379), .B(n13378), .ZN(n13400) );
  NAND2_X1 U16434 ( .A1(n13381), .A2(n13380), .ZN(n13383) );
  XNOR2_X1 U16435 ( .A(n13383), .B(n13382), .ZN(n13394) );
  NAND2_X1 U16436 ( .A1(n13394), .A2(n16296), .ZN(n13393) );
  OR2_X1 U16437 ( .A1(n13385), .A2(n13384), .ZN(n13387) );
  NAND2_X1 U16438 ( .A1(n13387), .A2(n13386), .ZN(n19154) );
  INV_X1 U16439 ( .A(n19154), .ZN(n19850) );
  INV_X1 U16440 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n19781) );
  OAI22_X1 U16441 ( .A1(n13388), .A2(n15445), .B1(n19781), .B2(n19089), .ZN(
        n13391) );
  MUX2_X1 U16442 ( .A(n15465), .B(n13389), .S(n13550), .Z(n13390) );
  AOI211_X1 U16443 ( .C1(n19850), .C2(n16306), .A(n13391), .B(n13390), .ZN(
        n13392) );
  OAI211_X1 U16444 ( .C1(n13400), .C2(n16312), .A(n13393), .B(n13392), .ZN(
        P2_U3043) );
  NAND2_X1 U16445 ( .A1(n13394), .A2(n16282), .ZN(n13399) );
  OAI21_X1 U16446 ( .B1(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n13395), .A(
        n13544), .ZN(n15742) );
  NOR2_X1 U16447 ( .A1(n16257), .A2(n15742), .ZN(n13397) );
  INV_X1 U16448 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n13605) );
  OAI22_X1 U16449 ( .A1(n16288), .A2(n13605), .B1(n19781), .B2(n19089), .ZN(
        n13396) );
  AOI211_X1 U16450 ( .C1(n10285), .C2(n16281), .A(n13397), .B(n13396), .ZN(
        n13398) );
  OAI211_X1 U16451 ( .C1(n13400), .C2(n16260), .A(n13399), .B(n13398), .ZN(
        P2_U3011) );
  INV_X1 U16452 ( .A(n13401), .ZN(n13403) );
  NAND4_X1 U16453 ( .A1(n13403), .A2(n11732), .A3(n13402), .A4(n14162), .ZN(
        n13404) );
  NAND2_X1 U16454 ( .A1(n13427), .A2(n20152), .ZN(n13407) );
  INV_X1 U16455 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13689) );
  NAND2_X1 U16456 ( .A1(n14162), .A2(n13689), .ZN(n13406) );
  NAND3_X1 U16457 ( .A1(n13407), .A2(n13423), .A3(n13406), .ZN(n13409) );
  NAND2_X1 U16458 ( .A1(n14155), .A2(n13689), .ZN(n13408) );
  AND2_X1 U16459 ( .A1(n13409), .A2(n13408), .ZN(n13421) );
  INV_X1 U16460 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20165) );
  NAND2_X1 U16461 ( .A1(n13427), .A2(n20165), .ZN(n13410) );
  INV_X1 U16462 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n13411) );
  NAND2_X1 U16463 ( .A1(n14155), .A2(n13411), .ZN(n13412) );
  NAND2_X1 U16464 ( .A1(n13427), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13414) );
  INV_X1 U16465 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n13575) );
  NAND2_X1 U16466 ( .A1(n13423), .A2(n13575), .ZN(n13413) );
  NAND2_X1 U16467 ( .A1(n13414), .A2(n13413), .ZN(n13573) );
  XNOR2_X1 U16468 ( .A(n13416), .B(n13573), .ZN(n20033) );
  NAND2_X1 U16469 ( .A1(n20033), .A2(n14162), .ZN(n13418) );
  INV_X1 U16470 ( .A(n13573), .ZN(n13415) );
  OR2_X1 U16471 ( .A1(n13416), .A2(n13415), .ZN(n13417) );
  INV_X1 U16472 ( .A(n13530), .ZN(n13419) );
  AOI21_X1 U16473 ( .B1(n13421), .B2(n13420), .A(n13419), .ZN(n20158) );
  AOI22_X1 U16474 ( .A1(n14403), .A2(n20158), .B1(n14402), .B2(
        P1_EBX_REG_2__SCAN_IN), .ZN(n13422) );
  OAI21_X1 U16475 ( .B1(n13694), .B2(n14405), .A(n13422), .ZN(P1_U2870) );
  MUX2_X1 U16476 ( .A(n14158), .B(n13423), .S(P1_EBX_REG_3__SCAN_IN), .Z(
        n13424) );
  OAI21_X1 U16477 ( .B1(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .B2(n14163), .A(
        n13424), .ZN(n13529) );
  MUX2_X1 U16478 ( .A(n13423), .B(n13427), .S(P1_EBX_REG_4__SCAN_IN), .Z(
        n13426) );
  NAND2_X1 U16479 ( .A1(n14198), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13425) );
  NAND2_X1 U16480 ( .A1(n13426), .A2(n13425), .ZN(n13576) );
  INV_X1 U16481 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n19990) );
  NAND2_X1 U16482 ( .A1(n14162), .A2(n19990), .ZN(n13429) );
  NAND2_X1 U16483 ( .A1(n13423), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13428) );
  NAND3_X1 U16484 ( .A1(n13429), .A2(n13427), .A3(n13428), .ZN(n13430) );
  OAI21_X1 U16485 ( .B1(n14158), .B2(P1_EBX_REG_5__SCAN_IN), .A(n13430), .ZN(
        n13535) );
  MUX2_X1 U16486 ( .A(n13423), .B(n13427), .S(P1_EBX_REG_6__SCAN_IN), .Z(
        n13434) );
  NAND2_X1 U16487 ( .A1(n14198), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13433) );
  NAND2_X1 U16488 ( .A1(n13533), .A2(n13435), .ZN(n13436) );
  AND2_X1 U16489 ( .A1(n13566), .A2(n13436), .ZN(n19973) );
  AOI22_X1 U16490 ( .A1(n19973), .A2(n14403), .B1(n14402), .B2(
        P1_EBX_REG_6__SCAN_IN), .ZN(n13437) );
  OAI21_X1 U16491 ( .B1(n13438), .B2(n14405), .A(n13437), .ZN(P1_U2866) );
  INV_X1 U16492 ( .A(n13439), .ZN(n20274) );
  OR2_X1 U16493 ( .A1(n13187), .A2(n13440), .ZN(n20506) );
  INV_X1 U16494 ( .A(n20506), .ZN(n20595) );
  INV_X1 U16495 ( .A(n13456), .ZN(n20659) );
  AOI21_X1 U16496 ( .B1(n20595), .B2(n20469), .A(n20659), .ZN(n13442) );
  OAI211_X1 U16497 ( .C1(n20559), .C2(n20274), .A(n20585), .B(n13442), .ZN(
        n13441) );
  OAI211_X1 U16498 ( .C1(n20589), .C2(n20585), .A(n20561), .B(n13441), .ZN(
        n20664) );
  OAI22_X1 U16499 ( .A1(n20529), .A2(n20667), .B1(n20204), .B2(n20620), .ZN(
        n13445) );
  INV_X1 U16500 ( .A(n20616), .ZN(n13515) );
  INV_X1 U16501 ( .A(n13442), .ZN(n13443) );
  AOI22_X1 U16502 ( .A1(n13443), .A2(n20585), .B1(n20589), .B2(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20645) );
  OAI22_X1 U16503 ( .A1(n13515), .A2(n20645), .B1(n13456), .B2(n20525), .ZN(
        n13444) );
  AOI211_X1 U16504 ( .C1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .C2(n20664), .A(
        n13445), .B(n13444), .ZN(n13446) );
  INV_X1 U16505 ( .A(n13446), .ZN(P1_U3156) );
  OAI22_X1 U16506 ( .A1(n20543), .A2(n20667), .B1(n20204), .B2(n20636), .ZN(
        n13448) );
  INV_X1 U16507 ( .A(n20632), .ZN(n13496) );
  OAI22_X1 U16508 ( .A1(n13496), .A2(n20645), .B1(n13456), .B2(n20539), .ZN(
        n13447) );
  AOI211_X1 U16509 ( .C1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .C2(n20664), .A(
        n13448), .B(n13447), .ZN(n13449) );
  INV_X1 U16510 ( .A(n13449), .ZN(P1_U3159) );
  OAI22_X1 U16511 ( .A1(n20520), .A2(n20667), .B1(n20204), .B2(n20610), .ZN(
        n13451) );
  INV_X1 U16512 ( .A(n20606), .ZN(n13488) );
  OAI22_X1 U16513 ( .A1(n13488), .A2(n20645), .B1(n13456), .B2(n20516), .ZN(
        n13450) );
  AOI211_X1 U16514 ( .C1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .C2(n20664), .A(
        n13451), .B(n13450), .ZN(n13452) );
  INV_X1 U16515 ( .A(n13452), .ZN(P1_U3154) );
  OAI22_X1 U16516 ( .A1(n20538), .A2(n20667), .B1(n20204), .B2(n20630), .ZN(
        n13454) );
  INV_X1 U16517 ( .A(n20626), .ZN(n13508) );
  OAI22_X1 U16518 ( .A1(n13508), .A2(n20645), .B1(n13456), .B2(n20534), .ZN(
        n13453) );
  AOI211_X1 U16519 ( .C1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .C2(n20664), .A(
        n13454), .B(n13453), .ZN(n13455) );
  INV_X1 U16520 ( .A(n13455), .ZN(P1_U3158) );
  OAI22_X1 U16521 ( .A1(n20515), .A2(n20667), .B1(n20204), .B2(n20604), .ZN(
        n13458) );
  INV_X1 U16522 ( .A(n20592), .ZN(n13504) );
  OAI22_X1 U16523 ( .A1(n13504), .A2(n20645), .B1(n13456), .B2(n20503), .ZN(
        n13457) );
  AOI211_X1 U16524 ( .C1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .C2(n20664), .A(
        n13458), .B(n13457), .ZN(n13459) );
  INV_X1 U16525 ( .A(n13459), .ZN(P1_U3153) );
  INV_X1 U16526 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n20030) );
  NOR2_X1 U16527 ( .A1(n20135), .A2(n20750), .ZN(n14714) );
  AND2_X1 U16528 ( .A1(n20120), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13460) );
  AOI211_X1 U16529 ( .C1(n20030), .C2(n15961), .A(n14714), .B(n13460), .ZN(
        n13464) );
  OR2_X1 U16530 ( .A1(n13461), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n14713) );
  NAND3_X1 U16531 ( .A1(n14713), .A2(n14712), .A3(n12697), .ZN(n13463) );
  OAI211_X1 U16532 ( .C1(n20027), .C2(n14616), .A(n13464), .B(n13463), .ZN(
        P1_U2998) );
  XNOR2_X1 U16533 ( .A(n13222), .B(n13465), .ZN(n13469) );
  AND2_X1 U16534 ( .A1(n9708), .A2(n13466), .ZN(n13467) );
  OR2_X1 U16535 ( .A1(n13467), .A2(n13518), .ZN(n16230) );
  MUX2_X1 U16536 ( .A(n16230), .B(n10609), .S(n14856), .Z(n13468) );
  OAI21_X1 U16537 ( .B1(n13469), .B2(n14865), .A(n13468), .ZN(P2_U2874) );
  AOI21_X1 U16538 ( .B1(n13479), .B2(n13511), .A(n20761), .ZN(n13470) );
  NOR2_X1 U16539 ( .A1(n13470), .A2(n20556), .ZN(n13477) );
  NOR2_X1 U16540 ( .A1(n20318), .A2(n20372), .ZN(n13475) );
  OR2_X1 U16541 ( .A1(n20435), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20243) );
  INV_X1 U16542 ( .A(n20243), .ZN(n13472) );
  OR2_X1 U16543 ( .A1(n13474), .A2(n20760), .ZN(n20587) );
  INV_X1 U16544 ( .A(n20587), .ZN(n13471) );
  AOI22_X1 U16545 ( .A1(n13477), .A2(n13475), .B1(n13472), .B2(n13471), .ZN(
        n13516) );
  INV_X1 U16546 ( .A(n20653), .ZN(n13484) );
  NOR2_X1 U16547 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n13473), .ZN(
        n13480) );
  NAND2_X1 U16548 ( .A1(n13474), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20436) );
  INV_X1 U16549 ( .A(n13475), .ZN(n13476) );
  AND2_X1 U16550 ( .A1(n20243), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20240) );
  AOI21_X1 U16551 ( .B1(n13477), .B2(n13476), .A(n20240), .ZN(n13478) );
  NAND2_X1 U16552 ( .A1(n13509), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n13483) );
  INV_X1 U16553 ( .A(n13480), .ZN(n13510) );
  OAI22_X1 U16554 ( .A1(n13511), .A2(n20624), .B1(n13510), .B2(n20530), .ZN(
        n13481) );
  AOI21_X1 U16555 ( .B1(n20365), .B2(n20621), .A(n13481), .ZN(n13482) );
  OAI211_X1 U16556 ( .C1(n13516), .C2(n13484), .A(n13483), .B(n13482), .ZN(
        P1_U3085) );
  NAND2_X1 U16557 ( .A1(n13509), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n13487) );
  OAI22_X1 U16558 ( .A1(n13511), .A2(n20610), .B1(n13510), .B2(n20516), .ZN(
        n13485) );
  AOI21_X1 U16559 ( .B1(n20365), .B2(n20607), .A(n13485), .ZN(n13486) );
  OAI211_X1 U16560 ( .C1(n13516), .C2(n13488), .A(n13487), .B(n13486), .ZN(
        P1_U3082) );
  INV_X1 U16561 ( .A(n20647), .ZN(n13492) );
  NAND2_X1 U16562 ( .A1(n13509), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(
        n13491) );
  OAI22_X1 U16563 ( .A1(n13511), .A2(n20614), .B1(n13510), .B2(n20521), .ZN(
        n13489) );
  AOI21_X1 U16564 ( .B1(n20365), .B2(n20611), .A(n13489), .ZN(n13490) );
  OAI211_X1 U16565 ( .C1(n13516), .C2(n13492), .A(n13491), .B(n13490), .ZN(
        P1_U3083) );
  NAND2_X1 U16566 ( .A1(n13509), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(
        n13495) );
  OAI22_X1 U16567 ( .A1(n13511), .A2(n20636), .B1(n13510), .B2(n20539), .ZN(
        n13493) );
  AOI21_X1 U16568 ( .B1(n20365), .B2(n20633), .A(n13493), .ZN(n13494) );
  OAI211_X1 U16569 ( .C1(n13516), .C2(n13496), .A(n13495), .B(n13494), .ZN(
        P1_U3087) );
  INV_X1 U16570 ( .A(n20661), .ZN(n13500) );
  NAND2_X1 U16571 ( .A1(n13509), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n13499) );
  OAI22_X1 U16572 ( .A1(n13511), .A2(n20644), .B1(n13510), .B2(n20545), .ZN(
        n13497) );
  AOI21_X1 U16573 ( .B1(n20365), .B2(n20639), .A(n13497), .ZN(n13498) );
  OAI211_X1 U16574 ( .C1(n13516), .C2(n13500), .A(n13499), .B(n13498), .ZN(
        P1_U3088) );
  NAND2_X1 U16575 ( .A1(n13509), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n13503) );
  OAI22_X1 U16576 ( .A1(n13511), .A2(n20604), .B1(n13510), .B2(n20503), .ZN(
        n13501) );
  AOI21_X1 U16577 ( .B1(n20365), .B2(n20601), .A(n13501), .ZN(n13502) );
  OAI211_X1 U16578 ( .C1(n13516), .C2(n13504), .A(n13503), .B(n13502), .ZN(
        P1_U3081) );
  NAND2_X1 U16579 ( .A1(n13509), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n13507) );
  OAI22_X1 U16580 ( .A1(n13511), .A2(n20630), .B1(n13510), .B2(n20534), .ZN(
        n13505) );
  AOI21_X1 U16581 ( .B1(n20365), .B2(n20627), .A(n13505), .ZN(n13506) );
  OAI211_X1 U16582 ( .C1(n13516), .C2(n13508), .A(n13507), .B(n13506), .ZN(
        P1_U3086) );
  NAND2_X1 U16583 ( .A1(n13509), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(
        n13514) );
  OAI22_X1 U16584 ( .A1(n13511), .A2(n20620), .B1(n13510), .B2(n20525), .ZN(
        n13512) );
  AOI21_X1 U16585 ( .B1(n20365), .B2(n20617), .A(n13512), .ZN(n13513) );
  OAI211_X1 U16586 ( .C1(n13516), .C2(n13515), .A(n13514), .B(n13513), .ZN(
        P1_U3084) );
  NOR2_X1 U16587 ( .A1(n13518), .A2(n13517), .ZN(n13519) );
  OR2_X1 U16588 ( .A1(n13679), .A2(n13519), .ZN(n15372) );
  NAND2_X1 U16589 ( .A1(n18971), .A2(n13520), .ZN(n13527) );
  INV_X1 U16590 ( .A(n13521), .ZN(n13525) );
  INV_X1 U16591 ( .A(n13522), .ZN(n13523) );
  OAI211_X1 U16592 ( .C1(n13525), .C2(n13524), .A(n14844), .B(n13523), .ZN(
        n13526) );
  OAI211_X1 U16593 ( .C1(n13520), .C2(n10873), .A(n13527), .B(n13526), .ZN(
        P2_U2873) );
  XNOR2_X1 U16594 ( .A(n20033), .B(n14162), .ZN(n14715) );
  AOI22_X1 U16595 ( .A1(n14403), .A2(n14715), .B1(n14402), .B2(
        P1_EBX_REG_1__SCAN_IN), .ZN(n13528) );
  OAI21_X1 U16596 ( .B1(n20027), .B2(n14387), .A(n13528), .ZN(P1_U2871) );
  AOI21_X1 U16597 ( .B1(n13530), .B2(n13529), .A(n13577), .ZN(n20145) );
  AOI22_X1 U16598 ( .A1(n14403), .A2(n20145), .B1(n14402), .B2(
        P1_EBX_REG_3__SCAN_IN), .ZN(n13531) );
  OAI21_X1 U16599 ( .B1(n13532), .B2(n14387), .A(n13531), .ZN(P1_U2869) );
  INV_X1 U16600 ( .A(n13533), .ZN(n13534) );
  AOI21_X1 U16601 ( .B1(n13535), .B2(n13579), .A(n13534), .ZN(n19988) );
  AOI22_X1 U16602 ( .A1(n19988), .A2(n14403), .B1(n14402), .B2(
        P1_EBX_REG_5__SCAN_IN), .ZN(n13536) );
  OAI21_X1 U16603 ( .B1(n13537), .B2(n14387), .A(n13536), .ZN(P1_U2867) );
  OAI21_X1 U16604 ( .B1(n13540), .B2(n13539), .A(n13538), .ZN(n13541) );
  INV_X1 U16605 ( .A(n13541), .ZN(n13560) );
  XOR2_X1 U16606 ( .A(n13543), .B(n13542), .Z(n13558) );
  INV_X1 U16607 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n19783) );
  OAI22_X1 U16608 ( .A1(n16288), .A2(n19083), .B1(n19783), .B2(n19089), .ZN(
        n13546) );
  AOI21_X1 U16609 ( .B1(n19083), .B2(n13544), .A(n15187), .ZN(n19081) );
  AND2_X1 U16610 ( .A1(n16279), .A2(n19081), .ZN(n13545) );
  NOR2_X1 U16611 ( .A1(n13546), .A2(n13545), .ZN(n13547) );
  OAI21_X1 U16612 ( .B1(n19092), .B2(n15182), .A(n13547), .ZN(n13548) );
  AOI21_X1 U16613 ( .B1(n13558), .B2(n16282), .A(n13548), .ZN(n13549) );
  OAI21_X1 U16614 ( .B1(n13560), .B2(n16260), .A(n13549), .ZN(P2_U3010) );
  OR2_X1 U16615 ( .A1(n13550), .A2(n15471), .ZN(n13712) );
  NOR2_X1 U16616 ( .A1(n16319), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13551) );
  NOR2_X1 U16617 ( .A1(n15465), .A2(n13551), .ZN(n13718) );
  NAND2_X1 U16618 ( .A1(P2_REIP_REG_4__SCAN_IN), .A2(n19069), .ZN(n13552) );
  OAI221_X1 U16619 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n13712), .C1(
        n13539), .C2(n13718), .A(n13552), .ZN(n13557) );
  NAND2_X1 U16620 ( .A1(n13553), .A2(n13386), .ZN(n13555) );
  INV_X1 U16621 ( .A(n13715), .ZN(n13554) );
  NAND2_X1 U16622 ( .A1(n13555), .A2(n13554), .ZN(n19144) );
  OAI22_X1 U16623 ( .A1(n19092), .A2(n15445), .B1(n15476), .B2(n19144), .ZN(
        n13556) );
  AOI211_X1 U16624 ( .C1(n13558), .C2(n16296), .A(n13557), .B(n13556), .ZN(
        n13559) );
  OAI21_X1 U16625 ( .B1(n13560), .B2(n16312), .A(n13559), .ZN(P2_U3042) );
  XOR2_X1 U16626 ( .A(n13561), .B(n13374), .Z(n19967) );
  INV_X1 U16627 ( .A(n19967), .ZN(n13585) );
  INV_X1 U16628 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n13562) );
  NAND2_X1 U16629 ( .A1(n14162), .A2(n13562), .ZN(n13564) );
  NAND2_X1 U16630 ( .A1(n13423), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n13563) );
  NAND3_X1 U16631 ( .A1(n13564), .A2(n13427), .A3(n13563), .ZN(n13565) );
  OAI21_X1 U16632 ( .B1(n14158), .B2(P1_EBX_REG_7__SCAN_IN), .A(n13565), .ZN(
        n13567) );
  AOI21_X1 U16633 ( .B1(n13567), .B2(n13566), .A(n9728), .ZN(n19961) );
  AOI22_X1 U16634 ( .A1(n19961), .A2(n14403), .B1(n14402), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n13568) );
  OAI21_X1 U16635 ( .B1(n13585), .B2(n14405), .A(n13568), .ZN(P1_U2865) );
  OAI21_X1 U16636 ( .B1(n13374), .B2(n13561), .A(n13570), .ZN(n13571) );
  AND2_X1 U16637 ( .A1(n13569), .A2(n13571), .ZN(n19956) );
  INV_X1 U16638 ( .A(n19956), .ZN(n13589) );
  INV_X1 U16639 ( .A(DATAI_8_), .ZN(n13572) );
  MUX2_X1 U16640 ( .A(n13572), .B(n16459), .S(n14410), .Z(n20069) );
  INV_X1 U16641 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n20802) );
  OAI222_X1 U16642 ( .A1(n13589), .A2(n14476), .B1(n20069), .B2(n14475), .C1(
        n14179), .C2(n20802), .ZN(P1_U2896) );
  OR2_X1 U16643 ( .A1(n14163), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13574) );
  NAND2_X1 U16644 ( .A1(n13574), .A2(n13573), .ZN(n13644) );
  OAI222_X1 U16645 ( .A1(n13644), .A2(n14379), .B1(n14377), .B2(n13575), .C1(
        n14387), .C2(n13657), .ZN(P1_U2872) );
  OR2_X1 U16646 ( .A1(n13577), .A2(n13576), .ZN(n13578) );
  NAND2_X1 U16647 ( .A1(n13579), .A2(n13578), .ZN(n20136) );
  INV_X1 U16648 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n13581) );
  OAI222_X1 U16649 ( .A1(n20136), .A2(n14379), .B1(n14377), .B2(n13581), .C1(
        n14387), .C2(n13580), .ZN(P1_U2868) );
  INV_X1 U16650 ( .A(n14989), .ZN(n13582) );
  OAI21_X1 U16651 ( .B1(n9659), .B2(n13583), .A(n13582), .ZN(n18965) );
  OAI222_X1 U16652 ( .A1(n18965), .A2(n19143), .B1(n19152), .B2(n12787), .C1(
        n13584), .C2(n19169), .ZN(P2_U2904) );
  OAI222_X1 U16653 ( .A1(n14476), .A2(n13585), .B1(n14179), .B2(n12085), .C1(
        n14475), .C2(n14438), .ZN(P1_U2897) );
  MUX2_X1 U16654 ( .A(n13423), .B(n13427), .S(P1_EBX_REG_8__SCAN_IN), .Z(
        n13587) );
  NAND2_X1 U16655 ( .A1(n14198), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13586) );
  NAND2_X1 U16656 ( .A1(n13587), .A2(n13586), .ZN(n13588) );
  OAI21_X1 U16657 ( .B1(n9728), .B2(n13588), .A(n13621), .ZN(n19952) );
  INV_X1 U16658 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n13590) );
  OAI222_X1 U16659 ( .A1(n19952), .A2(n14379), .B1(n13590), .B2(n14377), .C1(
        n13589), .C2(n14387), .ZN(P1_U2864) );
  INV_X1 U16660 ( .A(n19113), .ZN(n19093) );
  OAI22_X2 U16661 ( .A1(n14171), .A2(P2_STATE2_REG_0__SCAN_IN), .B1(n18853), 
        .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n13666) );
  AOI22_X1 U16662 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n18853), .ZN(n15488) );
  AOI22_X1 U16663 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(n19102), .B2(n18853), .ZN(
        n15487) );
  NAND2_X1 U16664 ( .A1(n15488), .A2(n15487), .ZN(n15486) );
  NOR2_X1 U16665 ( .A1(n13668), .A2(n15486), .ZN(n15743) );
  NOR2_X1 U16666 ( .A1(n13666), .A2(n15743), .ZN(n13592) );
  XNOR2_X1 U16667 ( .A(n13592), .B(n15742), .ZN(n13593) );
  NAND4_X1 U16668 ( .A1(n18853), .A2(n19691), .A3(n19896), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19116) );
  INV_X1 U16669 ( .A(n19116), .ZN(n19076) );
  NAND2_X1 U16670 ( .A1(n13593), .A2(n19076), .ZN(n13612) );
  AND2_X2 U16671 ( .A1(n19204), .A2(n19896), .ZN(n19112) );
  NAND2_X1 U16672 ( .A1(n19898), .A2(n19896), .ZN(n13594) );
  AND2_X1 U16673 ( .A1(n13595), .A2(n13594), .ZN(n13599) );
  AND2_X1 U16674 ( .A1(n14806), .A2(P2_EBX_REG_31__SCAN_IN), .ZN(n13596) );
  OR2_X1 U16675 ( .A1(n13598), .A2(n13597), .ZN(n16122) );
  NAND2_X1 U16676 ( .A1(n13599), .A2(n16123), .ZN(n13600) );
  NOR2_X1 U16677 ( .A1(n19697), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19752) );
  INV_X1 U16678 ( .A(n19752), .ZN(n13601) );
  NOR2_X1 U16679 ( .A1(n19754), .A2(n13601), .ZN(n16323) );
  NAND2_X1 U16680 ( .A1(n19089), .A2(n19116), .ZN(n13602) );
  OR2_X1 U16681 ( .A1(n16323), .A2(n13602), .ZN(n13603) );
  OAI22_X1 U16682 ( .A1(n13605), .A2(n19101), .B1(n19085), .B2(n19154), .ZN(
        n13607) );
  NOR2_X1 U16683 ( .A1(n19110), .A2(n19781), .ZN(n13606) );
  AOI211_X1 U16684 ( .C1(P2_EBX_REG_3__SCAN_IN), .C2(n19064), .A(n13607), .B(
        n13606), .ZN(n13608) );
  OAI21_X1 U16685 ( .B1(n13609), .B2(n19086), .A(n13608), .ZN(n13610) );
  AOI21_X1 U16686 ( .B1(n10285), .B2(n19112), .A(n13610), .ZN(n13611) );
  OAI211_X1 U16687 ( .C1(n19484), .C2(n19093), .A(n13612), .B(n13611), .ZN(
        P2_U2852) );
  AND2_X1 U16688 ( .A1(n13569), .A2(n13614), .ZN(n13615) );
  OR2_X1 U16689 ( .A1(n13613), .A2(n13615), .ZN(n19943) );
  INV_X1 U16690 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n13616) );
  NAND2_X1 U16691 ( .A1(n14162), .A2(n13616), .ZN(n13618) );
  NAND2_X1 U16692 ( .A1(n13423), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n13617) );
  NAND3_X1 U16693 ( .A1(n13618), .A2(n13427), .A3(n13617), .ZN(n13619) );
  OAI21_X1 U16694 ( .B1(n14158), .B2(P1_EBX_REG_9__SCAN_IN), .A(n13619), .ZN(
        n13622) );
  INV_X1 U16695 ( .A(n13701), .ZN(n13620) );
  AOI21_X1 U16696 ( .B1(n13622), .B2(n13621), .A(n13620), .ZN(n19938) );
  AOI22_X1 U16697 ( .A1(n19938), .A2(n14403), .B1(n14402), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n13623) );
  OAI21_X1 U16698 ( .B1(n19943), .B2(n14405), .A(n13623), .ZN(P1_U2863) );
  INV_X1 U16699 ( .A(DATAI_9_), .ZN(n20900) );
  INV_X1 U16700 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16457) );
  MUX2_X1 U16701 ( .A(n20900), .B(n16457), .S(n14410), .Z(n20072) );
  INV_X1 U16702 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n13624) );
  OAI222_X1 U16703 ( .A1(n19943), .A2(n14476), .B1(n20072), .B2(n14475), .C1(
        n13624), .C2(n14473), .ZN(P1_U2895) );
  INV_X1 U16704 ( .A(n13627), .ZN(n13628) );
  OAI21_X1 U16705 ( .B1(n13626), .B2(n13629), .A(n13628), .ZN(n15003) );
  NAND2_X1 U16706 ( .A1(n13677), .A2(n13630), .ZN(n13631) );
  NAND2_X1 U16707 ( .A1(n14860), .A2(n13631), .ZN(n18953) );
  MUX2_X1 U16708 ( .A(n18953), .B(n10610), .S(n14856), .Z(n13632) );
  OAI21_X1 U16709 ( .B1(n15003), .B2(n14865), .A(n13632), .ZN(P2_U2871) );
  AND2_X1 U16710 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n9755), .ZN(n13633) );
  INV_X1 U16711 ( .A(n15800), .ZN(n20763) );
  NOR2_X1 U16712 ( .A1(n20379), .A2(n20763), .ZN(n16111) );
  AOI22_X1 U16713 ( .A1(n13634), .A2(n13633), .B1(P1_STATE2_REG_0__SCAN_IN), 
        .B2(n16111), .ZN(n13635) );
  NAND2_X1 U16714 ( .A1(n20135), .A2(n13635), .ZN(n13636) );
  NOR2_X1 U16715 ( .A1(n13656), .A2(n13637), .ZN(n20028) );
  NOR2_X1 U16716 ( .A1(n13656), .A2(n13638), .ZN(n13648) );
  NAND2_X1 U16717 ( .A1(n20767), .A2(n20761), .ZN(n13640) );
  AOI21_X1 U16718 ( .B1(n13639), .B2(n15826), .A(n13640), .ZN(n13646) );
  NAND2_X1 U16719 ( .A1(n20017), .A2(n20029), .ZN(n19937) );
  NAND2_X1 U16720 ( .A1(n19937), .A2(P1_REIP_REG_0__SCAN_IN), .ZN(n13653) );
  AND2_X1 U16721 ( .A1(n13734), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n13645) );
  INV_X1 U16722 ( .A(n13645), .ZN(n13642) );
  INV_X1 U16723 ( .A(n13640), .ZN(n13641) );
  NOR2_X1 U16724 ( .A1(n13642), .A2(n13641), .ZN(n13643) );
  INV_X1 U16725 ( .A(n13644), .ZN(n14725) );
  NAND2_X1 U16726 ( .A1(n20034), .A2(n14725), .ZN(n13652) );
  NOR2_X1 U16727 ( .A1(n13646), .A2(n13645), .ZN(n13647) );
  NAND2_X1 U16728 ( .A1(n20026), .A2(P1_EBX_REG_0__SCAN_IN), .ZN(n13651) );
  AND2_X1 U16729 ( .A1(n13654), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13649) );
  OAI21_X1 U16730 ( .B1(n20013), .B2(n20014), .A(
        P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13650) );
  NAND4_X1 U16731 ( .A1(n13653), .A2(n13652), .A3(n13651), .A4(n13650), .ZN(
        n13659) );
  NOR2_X1 U16732 ( .A1(n13654), .A2(n20669), .ZN(n13655) );
  OAI21_X1 U16733 ( .B1(n13656), .B2(n14199), .A(n19942), .ZN(n20038) );
  INV_X1 U16734 ( .A(n20038), .ZN(n13693) );
  NOR2_X1 U16735 ( .A1(n13657), .A2(n13693), .ZN(n13658) );
  AOI211_X1 U16736 ( .C1(n20028), .C2(n11934), .A(n13659), .B(n13658), .ZN(
        n13660) );
  INV_X1 U16737 ( .A(n13660), .ZN(P1_U2840) );
  OAI21_X1 U16738 ( .B1(n13613), .B2(n13662), .A(n13661), .ZN(n13695) );
  INV_X1 U16739 ( .A(DATAI_10_), .ZN(n13664) );
  INV_X1 U16740 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n13663) );
  MUX2_X1 U16741 ( .A(n13664), .B(n13663), .S(n14410), .Z(n20077) );
  INV_X1 U16742 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n13665) );
  OAI222_X1 U16743 ( .A1(n13695), .A2(n14476), .B1(n20077), .B2(n14475), .C1(
        n13665), .C2(n14473), .ZN(P1_U2894) );
  NAND2_X1 U16744 ( .A1(n19080), .A2(n15486), .ZN(n13667) );
  XNOR2_X1 U16745 ( .A(n13668), .B(n13667), .ZN(n13669) );
  NAND2_X1 U16746 ( .A1(n13669), .A2(n19076), .ZN(n13676) );
  NAND2_X1 U16747 ( .A1(n19861), .A2(n19099), .ZN(n13672) );
  INV_X1 U16748 ( .A(n19064), .ZN(n19104) );
  OAI22_X1 U16749 ( .A1(n19104), .A2(n10235), .B1(n12808), .B2(n19101), .ZN(
        n13670) );
  AOI21_X1 U16750 ( .B1(n19070), .B2(P2_REIP_REG_2__SCAN_IN), .A(n13670), .ZN(
        n13671) );
  OAI211_X1 U16751 ( .C1(n19086), .C2(n13673), .A(n13672), .B(n13671), .ZN(
        n13674) );
  AOI21_X1 U16752 ( .B1(n9657), .B2(n19112), .A(n13674), .ZN(n13675) );
  OAI211_X1 U16753 ( .C1(n19859), .C2(n19093), .A(n13676), .B(n13675), .ZN(
        P2_U2853) );
  OAI21_X1 U16754 ( .B1(n13679), .B2(n13678), .A(n13677), .ZN(n18957) );
  NOR2_X1 U16755 ( .A1(n18957), .A2(n14856), .ZN(n13682) );
  AOI211_X1 U16756 ( .C1(n13680), .C2(n13523), .A(n14865), .B(n13626), .ZN(
        n13681) );
  AOI211_X1 U16757 ( .C1(P2_EBX_REG_15__SCAN_IN), .C2(n14856), .A(n13682), .B(
        n13681), .ZN(n13683) );
  INV_X1 U16758 ( .A(n13683), .ZN(P2_U2872) );
  INV_X1 U16759 ( .A(n20017), .ZN(n20019) );
  INV_X1 U16760 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20750) );
  NAND2_X1 U16761 ( .A1(n20019), .A2(n20750), .ZN(n20024) );
  INV_X1 U16762 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n13684) );
  AOI21_X1 U16763 ( .B1(n20024), .B2(n20029), .A(n13684), .ZN(n13691) );
  NOR3_X1 U16764 ( .A1(n20017), .A2(n20750), .A3(P1_REIP_REG_2__SCAN_IN), .ZN(
        n13685) );
  AOI21_X1 U16765 ( .B1(n20158), .B2(n20034), .A(n13685), .ZN(n13688) );
  INV_X1 U16766 ( .A(n20129), .ZN(n13686) );
  AOI22_X1 U16767 ( .A1(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n20013), .B1(
        n20014), .B2(n13686), .ZN(n13687) );
  OAI211_X1 U16768 ( .C1(n13689), .C2(n19991), .A(n13688), .B(n13687), .ZN(
        n13690) );
  AOI211_X1 U16769 ( .C1(n20028), .C2(n20177), .A(n13691), .B(n13690), .ZN(
        n13692) );
  OAI21_X1 U16770 ( .B1(n13694), .B2(n13693), .A(n13692), .ZN(P1_U2838) );
  INV_X1 U16771 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n13705) );
  INV_X1 U16772 ( .A(n13695), .ZN(n15962) );
  NAND2_X1 U16773 ( .A1(n15962), .A2(n13820), .ZN(n13704) );
  INV_X1 U16774 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15958) );
  NAND2_X1 U16775 ( .A1(n13427), .A2(n15958), .ZN(n13697) );
  NAND2_X1 U16776 ( .A1(n14162), .A2(n13705), .ZN(n13696) );
  NAND3_X1 U16777 ( .A1(n13697), .A2(n13423), .A3(n13696), .ZN(n13699) );
  NAND2_X1 U16778 ( .A1(n14155), .A2(n13705), .ZN(n13698) );
  AND2_X1 U16779 ( .A1(n13701), .A2(n13700), .ZN(n13702) );
  NOR2_X1 U16780 ( .A1(n13779), .A2(n13702), .ZN(n15896) );
  NAND2_X1 U16781 ( .A1(n15896), .A2(n14403), .ZN(n13703) );
  OAI211_X1 U16782 ( .C1(n13705), .C2(n14377), .A(n13704), .B(n13703), .ZN(
        P1_U2862) );
  NOR2_X1 U16783 ( .A1(n13707), .A2(n13706), .ZN(n13708) );
  XOR2_X1 U16784 ( .A(n13709), .B(n13708), .Z(n15193) );
  XNOR2_X1 U16785 ( .A(n13710), .B(n13711), .ZN(n15186) );
  INV_X1 U16786 ( .A(n15186), .ZN(n13723) );
  AOI221_X1 U16787 ( .B1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C1(n13717), .C2(n13539), .A(
        n13712), .ZN(n13722) );
  OAI21_X1 U16788 ( .B1(n13715), .B2(n13714), .A(n13713), .ZN(n19142) );
  INV_X1 U16789 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n13716) );
  NOR2_X1 U16790 ( .A1(n19089), .A2(n13716), .ZN(n15189) );
  AOI21_X1 U16791 ( .B1(n19074), .B2(n16316), .A(n15189), .ZN(n13720) );
  OR2_X1 U16792 ( .A1(n13718), .A2(n13717), .ZN(n13719) );
  OAI211_X1 U16793 ( .C1(n19142), .C2(n15476), .A(n13720), .B(n13719), .ZN(
        n13721) );
  AOI211_X1 U16794 ( .C1(n13723), .C2(n16296), .A(n13722), .B(n13721), .ZN(
        n13724) );
  OAI21_X1 U16795 ( .B1(n16312), .B2(n15193), .A(n13724), .ZN(P2_U3041) );
  XOR2_X1 U16796 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B(n13725), .Z(
        n13726) );
  XNOR2_X1 U16797 ( .A(n13727), .B(n13726), .ZN(n13772) );
  NAND2_X1 U16798 ( .A1(n13734), .A2(n15826), .ZN(n13728) );
  NAND2_X1 U16799 ( .A1(n13729), .A2(n13728), .ZN(n13733) );
  AOI22_X1 U16800 ( .A1(n15788), .A2(n11848), .B1(n20762), .B2(n15826), .ZN(
        n13731) );
  OAI21_X1 U16801 ( .B1(n13731), .B2(n11844), .A(n13730), .ZN(n13732) );
  MUX2_X1 U16802 ( .A(n13733), .B(n13732), .S(n13747), .Z(n13738) );
  NAND3_X1 U16803 ( .A1(n14197), .A2(n14739), .A3(n13734), .ZN(n13735) );
  OR2_X1 U16804 ( .A1(n9775), .A2(n13740), .ZN(n13741) );
  NAND2_X1 U16805 ( .A1(n13742), .A2(n13741), .ZN(n14187) );
  OAI21_X1 U16806 ( .B1(n13743), .B2(n13760), .A(n14187), .ZN(n13744) );
  OR2_X1 U16807 ( .A1(n13745), .A2(n13744), .ZN(n13746) );
  MUX2_X1 U16808 ( .A(n13748), .B(n13747), .S(n11848), .Z(n13749) );
  NAND3_X1 U16809 ( .A1(n13751), .A2(n13750), .A3(n13749), .ZN(n13752) );
  INV_X1 U16810 ( .A(n14191), .ZN(n13753) );
  NOR2_X1 U16811 ( .A1(n20152), .A2(n20165), .ZN(n14112) );
  NOR2_X1 U16812 ( .A1(n16030), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n20163) );
  NOR2_X1 U16813 ( .A1(n20164), .A2(n20163), .ZN(n14670) );
  NAND2_X1 U16814 ( .A1(n14112), .A2(n14670), .ZN(n16055) );
  INV_X1 U16815 ( .A(n16055), .ZN(n13757) );
  NOR2_X1 U16816 ( .A1(n20144), .A2(n20150), .ZN(n20138) );
  INV_X1 U16817 ( .A(n20138), .ZN(n13754) );
  NOR2_X1 U16818 ( .A1(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n13754), .ZN(
        n16101) );
  NOR2_X1 U16819 ( .A1(n16105), .A2(n13754), .ZN(n16051) );
  INV_X1 U16820 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20153) );
  OAI21_X1 U16821 ( .B1(n20153), .B2(n20165), .A(n20152), .ZN(n20131) );
  NAND2_X1 U16822 ( .A1(n16051), .A2(n20131), .ZN(n14113) );
  NAND2_X1 U16823 ( .A1(n14716), .A2(n20153), .ZN(n13756) );
  INV_X1 U16824 ( .A(n13762), .ZN(n13755) );
  NAND2_X1 U16825 ( .A1(n13755), .A2(n20135), .ZN(n16040) );
  NAND2_X1 U16826 ( .A1(n13756), .A2(n16040), .ZN(n20132) );
  AOI21_X1 U16827 ( .B1(n14685), .B2(n14113), .A(n20132), .ZN(n16072) );
  OAI221_X1 U16828 ( .B1(n20164), .B2(n14112), .C1(n20164), .C2(n20138), .A(
        n16072), .ZN(n16100) );
  AOI21_X1 U16829 ( .B1(n13757), .B2(n16101), .A(n16100), .ZN(n16097) );
  OAI21_X1 U16830 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16010), .A(
        n16097), .ZN(n16090) );
  OAI21_X1 U16831 ( .B1(n13760), .B2(n13759), .A(n13758), .ZN(n13761) );
  INV_X1 U16832 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20699) );
  OAI22_X1 U16833 ( .A1(n19952), .A2(n20137), .B1(n20699), .B2(n20135), .ZN(
        n13766) );
  INV_X1 U16834 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n16098) );
  NAND2_X1 U16835 ( .A1(n14685), .A2(n20131), .ZN(n13763) );
  NOR2_X1 U16836 ( .A1(n16098), .A2(n16099), .ZN(n16073) );
  NAND2_X1 U16837 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16074) );
  OAI211_X1 U16838 ( .C1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16073), .B(n16074), .ZN(n13764) );
  INV_X1 U16839 ( .A(n13764), .ZN(n13765) );
  AOI211_X1 U16840 ( .C1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(n16090), .A(
        n13766), .B(n13765), .ZN(n13767) );
  OAI21_X1 U16841 ( .B1(n13772), .B2(n16082), .A(n13767), .ZN(P1_U3023) );
  INV_X2 U16842 ( .A(n20135), .ZN(n20162) );
  AOI22_X1 U16843 ( .A1(n20120), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        n20162), .B2(P1_REIP_REG_8__SCAN_IN), .ZN(n13768) );
  OAI21_X1 U16844 ( .B1(n20130), .B2(n13769), .A(n13768), .ZN(n13770) );
  AOI21_X1 U16845 ( .B1(n19956), .B2(n20125), .A(n13770), .ZN(n13771) );
  OAI21_X1 U16846 ( .B1(n13772), .B2(n19918), .A(n13771), .ZN(P1_U2991) );
  OAI21_X1 U16847 ( .B1(n13773), .B2(n13775), .A(n13774), .ZN(n14615) );
  INV_X1 U16848 ( .A(n14611), .ZN(n13789) );
  MUX2_X1 U16849 ( .A(n14158), .B(n13423), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n13777) );
  OR2_X1 U16850 ( .A1(n14163), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n13776) );
  NOR2_X1 U16851 ( .A1(n13779), .A2(n13778), .ZN(n13780) );
  OR2_X1 U16852 ( .A1(n13811), .A2(n13780), .ZN(n13792) );
  INV_X1 U16853 ( .A(n13792), .ZN(n16063) );
  AOI22_X1 U16854 ( .A1(n20034), .A2(n16063), .B1(n20026), .B2(
        P1_EBX_REG_11__SCAN_IN), .ZN(n13782) );
  NAND2_X1 U16855 ( .A1(n20029), .A2(n13781), .ZN(n19974) );
  OAI211_X1 U16856 ( .C1(n20031), .C2(n13783), .A(n13782), .B(n19974), .ZN(
        n13788) );
  INV_X1 U16857 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n20697) );
  INV_X1 U16858 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n19980) );
  NAND4_X1 U16859 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_1__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n20004)
         );
  NOR3_X1 U16860 ( .A1(n20697), .A2(n19980), .A3(n20004), .ZN(n19966) );
  NAND2_X1 U16861 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n19966), .ZN(n19949) );
  NOR2_X1 U16862 ( .A1(n20699), .A2(n19949), .ZN(n14341) );
  INV_X1 U16863 ( .A(n14341), .ZN(n13784) );
  NAND3_X1 U16864 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .A3(n15895), .ZN(n15888) );
  INV_X1 U16865 ( .A(n15888), .ZN(n13786) );
  INV_X1 U16866 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n16076) );
  INV_X1 U16867 ( .A(P1_REIP_REG_9__SCAN_IN), .ZN(n19948) );
  AND2_X1 U16868 ( .A1(n20029), .A2(n14341), .ZN(n15848) );
  INV_X1 U16869 ( .A(n15848), .ZN(n19936) );
  NOR3_X1 U16870 ( .A1(n16076), .A2(n19948), .A3(n19936), .ZN(n15900) );
  NOR2_X1 U16871 ( .A1(n15899), .A2(n15900), .ZN(n13785) );
  MUX2_X1 U16872 ( .A(n13786), .B(n13785), .S(P1_REIP_REG_11__SCAN_IN), .Z(
        n13787) );
  AOI211_X1 U16873 ( .C1(n20014), .C2(n13789), .A(n13788), .B(n13787), .ZN(
        n13790) );
  OAI21_X1 U16874 ( .B1(n14615), .B2(n19942), .A(n13790), .ZN(P1_U2829) );
  INV_X1 U16875 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n20049) );
  OAI222_X1 U16876 ( .A1(n14615), .A2(n14476), .B1(n14420), .B2(n14475), .C1(
        n20049), .C2(n14473), .ZN(P1_U2893) );
  INV_X1 U16877 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n13791) );
  OAI222_X1 U16878 ( .A1(n13792), .A2(n14379), .B1(n13791), .B2(n14384), .C1(
        n14387), .C2(n14615), .ZN(P1_U2861) );
  OAI21_X1 U16879 ( .B1(n13795), .B2(n13794), .A(n13793), .ZN(n15886) );
  MUX2_X1 U16880 ( .A(n13423), .B(n13427), .S(P1_EBX_REG_12__SCAN_IN), .Z(
        n13797) );
  NAND2_X1 U16881 ( .A1(n14198), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n13796) );
  NAND2_X1 U16882 ( .A1(n13797), .A2(n13796), .ZN(n13810) );
  XNOR2_X1 U16883 ( .A(n13811), .B(n13810), .ZN(n15885) );
  INV_X1 U16884 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n13798) );
  OAI222_X1 U16885 ( .A1(n15886), .A2(n14405), .B1(n14379), .B2(n15885), .C1(
        n14377), .C2(n13798), .ZN(P1_U2860) );
  INV_X1 U16886 ( .A(DATAI_12_), .ZN(n13800) );
  INV_X1 U16887 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n13799) );
  MUX2_X1 U16888 ( .A(n13800), .B(n13799), .S(n14410), .Z(n20080) );
  INV_X1 U16889 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n13801) );
  OAI222_X1 U16890 ( .A1(n15886), .A2(n14476), .B1(n20080), .B2(n14475), .C1(
        n13801), .C2(n14179), .ZN(P1_U2892) );
  INV_X1 U16891 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n16075) );
  MUX2_X1 U16892 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B(n16075), .S(n9985), .Z(n13803) );
  XOR2_X1 U16893 ( .A(n13803), .B(n13802), .Z(n16086) );
  NAND2_X1 U16894 ( .A1(n16086), .A2(n12697), .ZN(n13806) );
  NAND2_X1 U16895 ( .A1(n20162), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n16083) );
  OAI21_X1 U16896 ( .B1(n14580), .B2(n19940), .A(n16083), .ZN(n13804) );
  AOI21_X1 U16897 ( .B1(n15961), .B2(n19946), .A(n13804), .ZN(n13805) );
  OAI211_X1 U16898 ( .C1(n14616), .C2(n19943), .A(n13806), .B(n13805), .ZN(
        P1_U2990) );
  OR2_X1 U16899 ( .A1(n13793), .A2(n14397), .ZN(n14395) );
  OR2_X1 U16900 ( .A1(n13793), .A2(n13807), .ZN(n14389) );
  INV_X1 U16901 ( .A(n14389), .ZN(n13808) );
  AOI21_X1 U16902 ( .B1(n13809), .B2(n14395), .A(n13808), .ZN(n14605) );
  MUX2_X1 U16903 ( .A(n14158), .B(n13423), .S(P1_EBX_REG_13__SCAN_IN), .Z(
        n13812) );
  OAI21_X1 U16904 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n14163), .A(
        n13812), .ZN(n14400) );
  INV_X1 U16905 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16027) );
  NAND2_X1 U16906 ( .A1(n13427), .A2(n16027), .ZN(n13814) );
  INV_X1 U16907 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n13823) );
  NAND2_X1 U16908 ( .A1(n14162), .A2(n13823), .ZN(n13813) );
  NAND3_X1 U16909 ( .A1(n13814), .A2(n13423), .A3(n13813), .ZN(n13816) );
  NAND2_X1 U16910 ( .A1(n14155), .A2(n13823), .ZN(n13815) );
  NAND2_X1 U16911 ( .A1(n14398), .A2(n13817), .ZN(n13818) );
  NAND2_X1 U16912 ( .A1(n14393), .A2(n13818), .ZN(n16022) );
  OAI22_X1 U16913 ( .A1(n16022), .A2(n14379), .B1(n13823), .B2(n14377), .ZN(
        n13819) );
  AOI21_X1 U16914 ( .B1(n14605), .B2(n13820), .A(n13819), .ZN(n13821) );
  INV_X1 U16915 ( .A(n13821), .ZN(P1_U2858) );
  INV_X1 U16916 ( .A(n14605), .ZN(n13833) );
  INV_X1 U16917 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n16021) );
  INV_X1 U16918 ( .A(P1_REIP_REG_12__SCAN_IN), .ZN(n15887) );
  INV_X1 U16919 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n15889) );
  NOR2_X1 U16920 ( .A1(n15887), .A2(n15889), .ZN(n15880) );
  NAND4_X1 U16921 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .A3(P1_REIP_REG_9__SCAN_IN), .A4(n15880), .ZN(n13822) );
  NOR2_X1 U16922 ( .A1(n16021), .A2(n13822), .ZN(n14203) );
  AOI21_X1 U16923 ( .B1(n14203), .B2(n15848), .A(n15899), .ZN(n15871) );
  OAI21_X1 U16924 ( .B1(n13822), .B2(n19941), .A(n16021), .ZN(n13828) );
  NOR2_X1 U16925 ( .A1(n16022), .A2(n20008), .ZN(n13827) );
  NOR2_X1 U16926 ( .A1(n19991), .A2(n13823), .ZN(n13824) );
  AOI211_X1 U16927 ( .C1(n20013), .C2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n20001), .B(n13824), .ZN(n13825) );
  OAI21_X1 U16928 ( .B1(n14603), .B2(n20042), .A(n13825), .ZN(n13826) );
  AOI211_X1 U16929 ( .C1(n15871), .C2(n13828), .A(n13827), .B(n13826), .ZN(
        n13829) );
  OAI21_X1 U16930 ( .B1(n13833), .B2(n19942), .A(n13829), .ZN(P1_U2826) );
  INV_X1 U16931 ( .A(DATAI_14_), .ZN(n13831) );
  INV_X1 U16932 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n13830) );
  MUX2_X1 U16933 ( .A(n13831), .B(n13830), .S(n14410), .Z(n20086) );
  INV_X1 U16934 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n13832) );
  OAI222_X1 U16935 ( .A1(n13833), .A2(n14476), .B1(n20086), .B2(n14475), .C1(
        n13832), .C2(n14473), .ZN(P1_U2890) );
  AND2_X1 U16936 ( .A1(n13834), .A2(n13835), .ZN(n13838) );
  OR2_X1 U16937 ( .A1(n13838), .A2(n13837), .ZN(n14592) );
  MUX2_X1 U16938 ( .A(n14158), .B(n13423), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n13839) );
  OAI21_X1 U16939 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n14163), .A(
        n13839), .ZN(n14392) );
  INV_X1 U16940 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n13840) );
  NAND2_X1 U16941 ( .A1(n13427), .A2(n13840), .ZN(n13842) );
  INV_X1 U16942 ( .A(P1_EBX_REG_16__SCAN_IN), .ZN(n13852) );
  NAND2_X1 U16943 ( .A1(n14162), .A2(n13852), .ZN(n13841) );
  NAND3_X1 U16944 ( .A1(n13842), .A2(n13423), .A3(n13841), .ZN(n13844) );
  NAND2_X1 U16945 ( .A1(n14155), .A2(n13852), .ZN(n13843) );
  NAND2_X1 U16946 ( .A1(n13844), .A2(n13843), .ZN(n13845) );
  OAI21_X1 U16947 ( .B1(n14391), .B2(n13845), .A(n13868), .ZN(n13853) );
  INV_X1 U16948 ( .A(n13853), .ZN(n16009) );
  AOI22_X1 U16949 ( .A1(n16009), .A2(n14403), .B1(n14402), .B2(
        P1_EBX_REG_16__SCAN_IN), .ZN(n13846) );
  OAI21_X1 U16950 ( .B1(n14592), .B2(n14387), .A(n13846), .ZN(P1_U2856) );
  INV_X1 U16951 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n13847) );
  NAND2_X1 U16952 ( .A1(n14203), .A2(n15895), .ZN(n13848) );
  NOR2_X1 U16953 ( .A1(n13847), .A2(n13848), .ZN(n15866) );
  INV_X1 U16954 ( .A(n15866), .ZN(n13850) );
  NOR2_X1 U16955 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n13848), .ZN(n15872) );
  NOR2_X1 U16956 ( .A1(n15871), .A2(n15872), .ZN(n13849) );
  MUX2_X1 U16957 ( .A(n13850), .B(n13849), .S(P1_REIP_REG_16__SCAN_IN), .Z(
        n13857) );
  AOI21_X1 U16958 ( .B1(n20013), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n20001), .ZN(n13851) );
  OAI21_X1 U16959 ( .B1(n19991), .B2(n13852), .A(n13851), .ZN(n13855) );
  NOR2_X1 U16960 ( .A1(n13853), .A2(n20008), .ZN(n13854) );
  AOI211_X1 U16961 ( .C1(n20014), .C2(n14589), .A(n13855), .B(n13854), .ZN(
        n13856) );
  OAI211_X1 U16962 ( .C1(n14592), .C2(n19942), .A(n13857), .B(n13856), .ZN(
        P1_U2824) );
  OAI22_X1 U16963 ( .A1(n14461), .A2(n13859), .B1(n13135), .B2(n14179), .ZN(
        n13860) );
  AOI21_X1 U16964 ( .B1(n14458), .B2(BUF1_REG_16__SCAN_IN), .A(n13860), .ZN(
        n13864) );
  NAND2_X1 U16965 ( .A1(n14468), .A2(DATAI_16_), .ZN(n13863) );
  OAI211_X1 U16966 ( .C1(n14592), .C2(n14476), .A(n13864), .B(n13863), .ZN(
        P1_U2888) );
  OAI21_X1 U16967 ( .B1(n13837), .B2(n13866), .A(n13865), .ZN(n15864) );
  MUX2_X1 U16968 ( .A(n14158), .B(n13423), .S(P1_EBX_REG_17__SCAN_IN), .Z(
        n13867) );
  OAI21_X1 U16969 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n14163), .A(
        n13867), .ZN(n13869) );
  INV_X1 U16970 ( .A(n14382), .ZN(n14371) );
  AOI21_X1 U16971 ( .B1(n13869), .B2(n13868), .A(n14371), .ZN(n16002) );
  AOI22_X1 U16972 ( .A1(n16002), .A2(n14403), .B1(n14402), .B2(
        P1_EBX_REG_17__SCAN_IN), .ZN(n13870) );
  OAI21_X1 U16973 ( .B1(n15864), .B2(n14387), .A(n13870), .ZN(P1_U2855) );
  OAI22_X1 U16974 ( .A1(n14461), .A2(n13871), .B1(n20901), .B2(n14179), .ZN(
        n13872) );
  AOI21_X1 U16975 ( .B1(n14458), .B2(BUF1_REG_17__SCAN_IN), .A(n13872), .ZN(
        n13874) );
  NAND2_X1 U16976 ( .A1(n14468), .A2(DATAI_17_), .ZN(n13873) );
  OAI211_X1 U16977 ( .C1(n15864), .C2(n14476), .A(n13874), .B(n13873), .ZN(
        P1_U2887) );
  AOI22_X1 U16978 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9634), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13890) );
  INV_X2 U16979 ( .A(n15538), .ZN(n17164) );
  AOI22_X1 U16980 ( .A1(n9645), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13889) );
  AOI22_X1 U16981 ( .A1(n9637), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n13876) );
  OAI21_X1 U16982 ( .B1(n17056), .B2(n17197), .A(n13876), .ZN(n13887) );
  INV_X2 U16983 ( .A(n15595), .ZN(n17128) );
  NOR2_X2 U16984 ( .A1(n13880), .A2(n13877), .ZN(n13971) );
  AOI22_X1 U16985 ( .A1(n17128), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13885) );
  NOR2_X2 U16986 ( .A1(n18656), .A2(n13879), .ZN(n13903) );
  AOI22_X1 U16987 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n13884) );
  AOI22_X1 U16988 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(n9639), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n13883) );
  INV_X2 U16989 ( .A(n17058), .ZN(n15584) );
  AOI22_X1 U16990 ( .A1(n15584), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n13882) );
  NAND4_X1 U16991 ( .A1(n13885), .A2(n13884), .A3(n13883), .A4(n13882), .ZN(
        n13886) );
  NAND3_X2 U16992 ( .A1(n13890), .A2(n13889), .A3(n9630), .ZN(n18233) );
  INV_X1 U16993 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16955) );
  AND2_X1 U16994 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(P3_EBX_REG_27__SCAN_IN), 
        .ZN(n14025) );
  INV_X1 U16995 ( .A(P3_EBX_REG_26__SCAN_IN), .ZN(n16606) );
  INV_X1 U16996 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16623) );
  INV_X1 U16997 ( .A(P3_EBX_REG_22__SCAN_IN), .ZN(n14024) );
  INV_X1 U16998 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n17014) );
  NOR4_X1 U16999 ( .A1(n16606), .A2(n16623), .A3(n14024), .A4(n17014), .ZN(
        n13891) );
  NAND4_X1 U17000 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(n14025), .A4(n13891), .ZN(n16963) );
  INV_X1 U17001 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n17030) );
  INV_X1 U17002 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n17069) );
  INV_X1 U17003 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16734) );
  INV_X1 U17004 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16763) );
  INV_X1 U17005 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n17126) );
  INV_X1 U17006 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n17155) );
  AOI22_X1 U17007 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13896) );
  BUF_X4 U17008 ( .A(n16929), .Z(n17180) );
  AOI22_X1 U17009 ( .A1(n9637), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n13895) );
  AOI22_X1 U17010 ( .A1(n17164), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n13894) );
  AOI22_X1 U17011 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(n9639), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n13893) );
  NAND4_X1 U17012 ( .A1(n13896), .A2(n13895), .A3(n13894), .A4(n13893), .ZN(
        n13902) );
  AOI22_X1 U17013 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13900) );
  AOI22_X1 U17014 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n17016), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13899) );
  AOI22_X1 U17015 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13898) );
  AOI22_X1 U17016 ( .A1(n15584), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13897) );
  NAND4_X1 U17017 ( .A1(n13900), .A2(n13899), .A3(n13898), .A4(n13897), .ZN(
        n13901) );
  AOI22_X1 U17018 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n13913) );
  AOI22_X1 U17019 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n13912) );
  AOI22_X1 U17020 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(n9639), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n13904) );
  OAI21_X1 U17021 ( .B1(n15595), .B2(n20908), .A(n13904), .ZN(n13910) );
  INV_X2 U17022 ( .A(n15538), .ZN(n15519) );
  AOI22_X1 U17023 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n15519), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n13908) );
  AOI22_X1 U17024 ( .A1(n9645), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n14027), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n13907) );
  AOI22_X1 U17025 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n13906) );
  AOI22_X1 U17026 ( .A1(n9637), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n13905) );
  NAND4_X1 U17027 ( .A1(n13908), .A2(n13907), .A3(n13906), .A4(n13905), .ZN(
        n13909) );
  AOI211_X2 U17028 ( .C1(n17180), .C2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A(
        n13910), .B(n13909), .ZN(n13911) );
  NAND3_X2 U17029 ( .A1(n13913), .A2(n13912), .A3(n13911), .ZN(n18196) );
  INV_X1 U17030 ( .A(n13914), .ZN(n14008) );
  OAI21_X1 U17031 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18638), .A(
        n14008), .ZN(n15660) );
  AOI22_X1 U17032 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18639), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18806), .ZN(n14009) );
  AOI22_X1 U17033 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18193), .B1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18799), .ZN(n13920) );
  NAND2_X1 U17034 ( .A1(n14009), .A2(n13914), .ZN(n13915) );
  NAND2_X1 U17035 ( .A1(n13920), .A2(n13919), .ZN(n13916) );
  OAI21_X1 U17036 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18799), .A(
        n13916), .ZN(n13917) );
  OAI22_X1 U17037 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18192), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n13917), .ZN(n13921) );
  NOR2_X1 U17038 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18192), .ZN(
        n13918) );
  NAND2_X1 U17039 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n13917), .ZN(
        n13922) );
  AOI22_X1 U17040 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n13921), .B1(
        n13918), .B2(n13922), .ZN(n13925) );
  NAND2_X1 U17041 ( .A1(n14009), .A2(n13925), .ZN(n13927) );
  XOR2_X1 U17042 ( .A(n13920), .B(n13919), .Z(n13926) );
  AOI21_X1 U17043 ( .B1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n13922), .A(
        n13921), .ZN(n13923) );
  AOI21_X1 U17044 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18192), .A(
        n13923), .ZN(n14006) );
  INV_X1 U17045 ( .A(n14006), .ZN(n13924) );
  AOI22_X1 U17046 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n13931) );
  AOI22_X1 U17047 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13930) );
  AOI22_X1 U17048 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9639), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n13929) );
  AOI22_X1 U17049 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n13928) );
  NAND4_X1 U17050 ( .A1(n13931), .A2(n13930), .A3(n13929), .A4(n13928), .ZN(
        n13938) );
  AOI22_X1 U17051 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n15519), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13936) );
  AOI22_X1 U17052 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13935) );
  AOI22_X1 U17053 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n9637), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13934) );
  AOI22_X1 U17054 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17128), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13933) );
  NAND4_X1 U17055 ( .A1(n13936), .A2(n13935), .A3(n13934), .A4(n13933), .ZN(
        n13937) );
  AOI22_X1 U17056 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n15519), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13942) );
  AOI22_X1 U17057 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n13971), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13941) );
  AOI22_X1 U17058 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13940) );
  AOI22_X1 U17059 ( .A1(n9637), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n13939) );
  NAND4_X1 U17060 ( .A1(n13942), .A2(n13941), .A3(n13940), .A4(n13939), .ZN(
        n13948) );
  AOI22_X1 U17061 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n13946) );
  AOI22_X1 U17062 ( .A1(n9645), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(n9639), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n13945) );
  AOI22_X1 U17063 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13944) );
  AOI22_X1 U17064 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13943) );
  NAND4_X1 U17065 ( .A1(n13946), .A2(n13945), .A3(n13944), .A4(n13943), .ZN(
        n13947) );
  INV_X1 U17066 ( .A(n13987), .ZN(n18218) );
  NAND2_X1 U17067 ( .A1(n13985), .A2(n18218), .ZN(n18647) );
  AOI22_X1 U17068 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(n9639), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n13958) );
  AOI22_X1 U17069 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13957) );
  INV_X1 U17070 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n17204) );
  AOI22_X1 U17071 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n15519), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13949) );
  OAI21_X1 U17072 ( .B1(n17056), .B2(n17204), .A(n13949), .ZN(n13955) );
  AOI22_X1 U17073 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13953) );
  AOI22_X1 U17074 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n13952) );
  AOI22_X1 U17075 ( .A1(n9637), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(n9641), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13951) );
  AOI22_X1 U17076 ( .A1(n17180), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n13950) );
  NAND4_X1 U17077 ( .A1(n13953), .A2(n13952), .A3(n13951), .A4(n13950), .ZN(
        n13954) );
  INV_X1 U17078 ( .A(n18634), .ZN(n15834) );
  AOI22_X1 U17079 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17016), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13962) );
  AOI22_X1 U17080 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13961) );
  AOI22_X1 U17081 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17128), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13960) );
  AOI22_X1 U17082 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n13959) );
  NAND4_X1 U17083 ( .A1(n13962), .A2(n13961), .A3(n13960), .A4(n13959), .ZN(
        n13968) );
  AOI22_X1 U17084 ( .A1(n9637), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(n9639), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n13966) );
  AOI22_X1 U17085 ( .A1(n17180), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13965) );
  AOI22_X1 U17086 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13964) );
  AOI22_X1 U17087 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15519), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13963) );
  NAND4_X1 U17088 ( .A1(n13966), .A2(n13965), .A3(n13964), .A4(n13963), .ZN(
        n13967) );
  AOI22_X1 U17089 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13980) );
  AOI22_X1 U17090 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9639), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n13979) );
  INV_X1 U17091 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17212) );
  AOI22_X1 U17092 ( .A1(n17180), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13969) );
  OAI21_X1 U17093 ( .B1(n17056), .B2(n17212), .A(n13969), .ZN(n13977) );
  AOI22_X1 U17094 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13975) );
  AOI22_X1 U17095 ( .A1(n9637), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n15519), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13974) );
  AOI22_X1 U17096 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n13973) );
  AOI22_X1 U17097 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13972) );
  NAND4_X1 U17098 ( .A1(n13975), .A2(n13974), .A3(n13973), .A4(n13972), .ZN(
        n13976) );
  AOI211_X1 U17099 ( .C1(n15584), .C2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A(
        n13977), .B(n13976), .ZN(n13978) );
  NAND3_X1 U17100 ( .A1(n13980), .A2(n13979), .A3(n13978), .ZN(n18213) );
  NAND2_X1 U17101 ( .A1(n18233), .A2(n18213), .ZN(n15653) );
  NOR2_X1 U17102 ( .A1(n13985), .A2(n18223), .ZN(n14013) );
  INV_X1 U17103 ( .A(n14013), .ZN(n13986) );
  INV_X1 U17104 ( .A(n18213), .ZN(n13996) );
  NAND2_X1 U17105 ( .A1(n14002), .A2(n13996), .ZN(n18646) );
  NOR2_X1 U17106 ( .A1(n18779), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n18688) );
  NAND2_X1 U17107 ( .A1(n18688), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18675) );
  INV_X1 U17108 ( .A(P3_EBX_REG_4__SCAN_IN), .ZN(n16865) );
  NAND3_X1 U17109 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n17211) );
  OR3_X1 U17110 ( .A1(n16865), .A2(n17207), .A3(n17211), .ZN(n17192) );
  NAND2_X1 U17111 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n9700), .ZN(n17000) );
  NOR3_X1 U17112 ( .A1(n16955), .A2(n16963), .A3(n17000), .ZN(n16928) );
  NAND2_X1 U17113 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16928), .ZN(n13982) );
  NOR2_X1 U17114 ( .A1(n18233), .A2(n13982), .ZN(n13984) );
  NAND2_X1 U17115 ( .A1(n17220), .A2(n13982), .ZN(n16953) );
  INV_X1 U17116 ( .A(n16953), .ZN(n13983) );
  MUX2_X1 U17117 ( .A(n13984), .B(n13983), .S(P3_EBX_REG_31__SCAN_IN), .Z(
        P3_U2672) );
  INV_X1 U17118 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18792) );
  NAND2_X1 U17119 ( .A1(n18792), .A2(n18782), .ZN(n18844) );
  OR4_X2 U17120 ( .A1(n18218), .A2(n18213), .A3(n14004), .A4(n13990), .ZN(
        n14001) );
  NAND3_X1 U17121 ( .A1(n14002), .A2(n18647), .A3(n13986), .ZN(n13993) );
  NAND2_X1 U17122 ( .A1(n14002), .A2(n18223), .ZN(n15665) );
  NAND2_X1 U17123 ( .A1(n18834), .A2(n18196), .ZN(n15647) );
  AOI21_X1 U17124 ( .B1(n18233), .B2(n18634), .A(n15647), .ZN(n14018) );
  AOI21_X1 U17125 ( .B1(n13993), .B2(n15665), .A(n14018), .ZN(n13995) );
  NAND2_X1 U17126 ( .A1(n13987), .A2(n18634), .ZN(n13999) );
  NOR2_X1 U17127 ( .A1(n13987), .A2(n17074), .ZN(n13988) );
  NAND2_X1 U17128 ( .A1(n13990), .A2(n13988), .ZN(n13991) );
  NAND2_X1 U17129 ( .A1(n14002), .A2(n15648), .ZN(n13989) );
  AOI22_X1 U17130 ( .A1(n13999), .A2(n13991), .B1(n13990), .B2(n13989), .ZN(
        n13992) );
  OAI21_X1 U17131 ( .B1(n18196), .B2(n13993), .A(n13992), .ZN(n13994) );
  INV_X1 U17132 ( .A(n15651), .ZN(n14005) );
  NAND2_X1 U17133 ( .A1(n18834), .A2(n13997), .ZN(n14003) );
  NOR4_X4 U17134 ( .A1(n16534), .A2(n18228), .A3(n14000), .A4(n13999), .ZN(
        n17424) );
  NOR2_X2 U17135 ( .A1(n14002), .A2(n14001), .ZN(n14015) );
  NOR2_X2 U17136 ( .A1(n16515), .A2(n15648), .ZN(n14010) );
  NOR2_X2 U17137 ( .A1(n17424), .A2(n14010), .ZN(n18624) );
  INV_X1 U17138 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n16864) );
  OAI21_X1 U17139 ( .B1(n18659), .B2(n18789), .A(n16864), .ZN(n15531) );
  NAND2_X1 U17140 ( .A1(n16533), .A2(n15531), .ZN(n18671) );
  NOR2_X1 U17141 ( .A1(n18844), .A2(n18671), .ZN(n14023) );
  NAND2_X1 U17142 ( .A1(n18779), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18194) );
  INV_X1 U17143 ( .A(n18194), .ZN(n14022) );
  OAI21_X1 U17144 ( .B1(n14009), .B2(n14008), .A(n14006), .ZN(n14007) );
  AOI21_X1 U17145 ( .B1(n14009), .B2(n14008), .A(n14007), .ZN(n15661) );
  NAND2_X1 U17146 ( .A1(READY22_REG_SCAN_IN), .A2(READY2), .ZN(n18835) );
  INV_X1 U17147 ( .A(n18835), .ZN(n18829) );
  OR2_X1 U17148 ( .A1(n18626), .A2(n18829), .ZN(n15832) );
  AOI21_X1 U17149 ( .B1(n17424), .B2(n18204), .A(n16533), .ZN(n15831) );
  NOR2_X1 U17150 ( .A1(n18834), .A2(n14010), .ZN(n15654) );
  INV_X1 U17151 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18710) );
  INV_X1 U17152 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n18699) );
  INV_X2 U17153 ( .A(n18842), .ZN(n20776) );
  NOR2_X1 U17154 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18697) );
  INV_X1 U17155 ( .A(n18697), .ZN(n14011) );
  NAND3_X1 U17156 ( .A1(n18710), .A2(n18769), .A3(n14011), .ZN(n18832) );
  OR3_X1 U17157 ( .A1(n18624), .A2(n15654), .A3(n18832), .ZN(n17384) );
  INV_X1 U17158 ( .A(n15648), .ZN(n14014) );
  NOR3_X1 U17159 ( .A1(n14014), .A2(n14013), .A3(n14012), .ZN(n15658) );
  AOI21_X1 U17160 ( .B1(n15658), .B2(n14016), .A(n14015), .ZN(n14017) );
  OAI221_X1 U17161 ( .B1(n15832), .B2(n15831), .C1(n15832), .C2(n17384), .A(
        n15671), .ZN(n14019) );
  NOR2_X1 U17162 ( .A1(n14020), .A2(n14019), .ZN(n18664) );
  INV_X1 U17163 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n16517) );
  NAND3_X1 U17164 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18781)
         );
  OAI22_X1 U17165 ( .A1(n18664), .A2(n18675), .B1(n16517), .B2(n18781), .ZN(
        n14021) );
  MUX2_X1 U17166 ( .A(n14023), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18814), .Z(P3_U3284) );
  NAND2_X1 U17167 ( .A1(n17074), .A2(n17222), .ZN(n17228) );
  INV_X1 U17168 ( .A(P3_EBX_REG_24__SCAN_IN), .ZN(n16628) );
  INV_X1 U17169 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16640) );
  INV_X1 U17170 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n17028) );
  NAND2_X1 U17171 ( .A1(n17220), .A2(n16969), .ZN(n16967) );
  OAI21_X1 U17172 ( .B1(n14025), .B2(n17228), .A(n16967), .ZN(n16960) );
  AOI22_X1 U17173 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(n9639), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n14031) );
  AOI22_X1 U17174 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n14030) );
  AOI22_X1 U17175 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9637), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n14029) );
  AOI22_X1 U17176 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n14028) );
  NAND4_X1 U17177 ( .A1(n14031), .A2(n14030), .A3(n14029), .A4(n14028), .ZN(
        n14037) );
  AOI22_X1 U17178 ( .A1(n15584), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n15519), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n14035) );
  AOI22_X1 U17179 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n14034) );
  AOI22_X1 U17180 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n14033) );
  AOI22_X1 U17181 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n14032) );
  NAND4_X1 U17182 ( .A1(n14035), .A2(n14034), .A3(n14033), .A4(n14032), .ZN(
        n14036) );
  NOR2_X1 U17183 ( .A1(n14037), .A2(n14036), .ZN(n16965) );
  AOI22_X1 U17184 ( .A1(n9645), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9639), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n14041) );
  AOI22_X1 U17185 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15519), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n14040) );
  AOI22_X1 U17186 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17128), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n14039) );
  AOI22_X1 U17187 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n14038) );
  NAND4_X1 U17188 ( .A1(n14041), .A2(n14040), .A3(n14039), .A4(n14038), .ZN(
        n14047) );
  AOI22_X1 U17189 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n9637), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n14045) );
  AOI22_X1 U17190 ( .A1(n14026), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n14044) );
  AOI22_X1 U17191 ( .A1(n17180), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n14043) );
  AOI22_X1 U17192 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n14042) );
  NAND4_X1 U17193 ( .A1(n14045), .A2(n14044), .A3(n14043), .A4(n14042), .ZN(
        n14046) );
  NOR2_X1 U17194 ( .A1(n14047), .A2(n14046), .ZN(n16975) );
  AOI22_X1 U17195 ( .A1(n15584), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n14051) );
  AOI22_X1 U17196 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13971), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n14050) );
  AOI22_X1 U17197 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n14049) );
  AOI22_X1 U17198 ( .A1(n9645), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n14048) );
  NAND4_X1 U17199 ( .A1(n14051), .A2(n14050), .A3(n14049), .A4(n14048), .ZN(
        n14057) );
  AOI22_X1 U17200 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15519), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n14055) );
  AOI22_X1 U17201 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n9639), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n14054) );
  AOI22_X1 U17202 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n14053) );
  AOI22_X1 U17203 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9637), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n14052) );
  NAND4_X1 U17204 ( .A1(n14055), .A2(n14054), .A3(n14053), .A4(n14052), .ZN(
        n14056) );
  NOR2_X1 U17205 ( .A1(n14057), .A2(n14056), .ZN(n16985) );
  AOI22_X1 U17206 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n17128), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n14061) );
  AOI22_X1 U17207 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(n9634), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n14060) );
  AOI22_X1 U17208 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n14059) );
  AOI22_X1 U17209 ( .A1(n9645), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n14058) );
  NAND4_X1 U17210 ( .A1(n14061), .A2(n14060), .A3(n14059), .A4(n14058), .ZN(
        n14067) );
  AOI22_X1 U17211 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n14065) );
  AOI22_X1 U17212 ( .A1(n9639), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n15519), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n14064) );
  AOI22_X1 U17213 ( .A1(n15584), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n14063) );
  AOI22_X1 U17214 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9637), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n14062) );
  NAND4_X1 U17215 ( .A1(n14065), .A2(n14064), .A3(n14063), .A4(n14062), .ZN(
        n14066) );
  NOR2_X1 U17216 ( .A1(n14067), .A2(n14066), .ZN(n16984) );
  NOR2_X1 U17217 ( .A1(n16985), .A2(n16984), .ZN(n16981) );
  AOI22_X1 U17218 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17144), .B1(
        n9639), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n14078) );
  AOI22_X1 U17219 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17174), .B1(
        n9637), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n14077) );
  INV_X1 U17220 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n17221) );
  AOI22_X1 U17221 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n17181), .B1(
        n17128), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n14069) );
  OAI21_X1 U17222 ( .B1(n16931), .B2(n17221), .A(n14069), .ZN(n14075) );
  AOI22_X1 U17223 ( .A1(n17180), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n9635), .ZN(n14073) );
  INV_X2 U17224 ( .A(n17056), .ZN(n17182) );
  AOI22_X1 U17225 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n14072) );
  AOI22_X1 U17226 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n9641), .ZN(n14071) );
  AOI22_X1 U17227 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17159), .B1(
        n15519), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n14070) );
  NAND4_X1 U17228 ( .A1(n14073), .A2(n14072), .A3(n14071), .A4(n14070), .ZN(
        n14074) );
  AOI211_X1 U17229 ( .C1(n17145), .C2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A(
        n14075), .B(n14074), .ZN(n14076) );
  NAND3_X1 U17230 ( .A1(n14078), .A2(n14077), .A3(n14076), .ZN(n16980) );
  NAND2_X1 U17231 ( .A1(n16981), .A2(n16980), .ZN(n16979) );
  NOR2_X1 U17232 ( .A1(n16975), .A2(n16979), .ZN(n16972) );
  AOI22_X1 U17233 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9639), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n14088) );
  AOI22_X1 U17234 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n15519), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n14087) );
  AOI22_X1 U17235 ( .A1(n15584), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17128), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n14079) );
  OAI21_X1 U17236 ( .B1(n16931), .B2(n17212), .A(n14079), .ZN(n14085) );
  AOI22_X1 U17237 ( .A1(n9645), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n13903), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n14083) );
  AOI22_X1 U17238 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n14082) );
  AOI22_X1 U17239 ( .A1(n9634), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n14081) );
  AOI22_X1 U17240 ( .A1(n9637), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n9641), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n14080) );
  NAND4_X1 U17241 ( .A1(n14083), .A2(n14082), .A3(n14081), .A4(n14080), .ZN(
        n14084) );
  AOI211_X1 U17242 ( .C1(n17145), .C2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A(
        n14085), .B(n14084), .ZN(n14086) );
  NAND3_X1 U17243 ( .A1(n14088), .A2(n14087), .A3(n14086), .ZN(n16971) );
  NAND2_X1 U17244 ( .A1(n16972), .A2(n16971), .ZN(n16970) );
  NOR2_X1 U17245 ( .A1(n16965), .A2(n16970), .ZN(n16964) );
  INV_X1 U17246 ( .A(n16964), .ZN(n16957) );
  AOI22_X1 U17247 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n14092) );
  AOI22_X1 U17248 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(n9639), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n14091) );
  AOI22_X1 U17249 ( .A1(n9634), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n15519), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n14090) );
  AOI22_X1 U17250 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n14089) );
  NAND4_X1 U17251 ( .A1(n14092), .A2(n14091), .A3(n14090), .A4(n14089), .ZN(
        n14098) );
  AOI22_X1 U17252 ( .A1(n15584), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17128), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n14096) );
  AOI22_X1 U17253 ( .A1(n9637), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n14095) );
  AOI22_X1 U17254 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n14094) );
  AOI22_X1 U17255 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n13903), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n14093) );
  NAND4_X1 U17256 ( .A1(n14096), .A2(n14095), .A3(n14094), .A4(n14093), .ZN(
        n14097) );
  NOR2_X1 U17257 ( .A1(n14098), .A2(n14097), .ZN(n16956) );
  XOR2_X1 U17258 ( .A(n16957), .B(n16956), .Z(n17245) );
  AOI22_X1 U17259 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16960), .B1(n17226), 
        .B2(n17245), .ZN(n14101) );
  INV_X1 U17260 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n14099) );
  INV_X1 U17261 ( .A(n16969), .ZN(n16974) );
  NAND3_X1 U17262 ( .A1(P3_EBX_REG_27__SCAN_IN), .A2(n14099), .A3(n16974), 
        .ZN(n14100) );
  NAND2_X1 U17263 ( .A1(n14101), .A2(n14100), .ZN(P3_U2675) );
  NAND2_X1 U17264 ( .A1(n11934), .A2(n14102), .ZN(n14104) );
  NAND2_X1 U17265 ( .A1(n14739), .A2(n14107), .ZN(n14103) );
  NAND2_X1 U17266 ( .A1(n14104), .A2(n14103), .ZN(n15764) );
  INV_X1 U17267 ( .A(n15764), .ZN(n14105) );
  OAI21_X1 U17268 ( .B1(n14105), .B2(P1_STATE2_REG_3__SCAN_IN), .A(n20669), 
        .ZN(n14106) );
  NOR2_X1 U17269 ( .A1(n20669), .A2(n20153), .ZN(n14747) );
  INV_X1 U17270 ( .A(n14747), .ZN(n14753) );
  AOI22_X1 U17271 ( .A1(n14106), .A2(n14753), .B1(n15801), .B2(n14107), .ZN(
        n14110) );
  AOI21_X1 U17272 ( .B1(n15762), .B2(n19909), .A(n14109), .ZN(n14108) );
  OAI22_X1 U17273 ( .A1(n14110), .A2(n14109), .B1(n14108), .B2(n14107), .ZN(
        P1_U3474) );
  INV_X1 U17274 ( .A(n20164), .ZN(n20134) );
  NAND2_X1 U17275 ( .A1(n14112), .A2(n16051), .ZN(n16069) );
  INV_X1 U17276 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n16049) );
  NOR4_X1 U17277 ( .A1(n15958), .A2(n16075), .A3(n16098), .A4(n16074), .ZN(
        n16050) );
  INV_X1 U17278 ( .A(n16050), .ZN(n16052) );
  NOR2_X1 U17279 ( .A1(n16049), .A2(n16052), .ZN(n16057) );
  NAND2_X1 U17280 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16057), .ZN(
        n14127) );
  NOR2_X1 U17281 ( .A1(n16069), .A2(n14127), .ZN(n16037) );
  INV_X1 U17282 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n16000) );
  NAND3_X1 U17283 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n16001) );
  NOR2_X1 U17284 ( .A1(n16000), .A2(n16001), .ZN(n14709) );
  NAND3_X1 U17285 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n14709), .ZN(n14686) );
  INV_X1 U17286 ( .A(n14686), .ZN(n14114) );
  NAND2_X1 U17287 ( .A1(n16037), .A2(n14114), .ZN(n14684) );
  NOR2_X1 U17288 ( .A1(n14127), .A2(n14113), .ZN(n16038) );
  AOI21_X1 U17289 ( .B1(n14114), .B2(n16038), .A(n20154), .ZN(n14115) );
  AOI211_X1 U17290 ( .C1(n20134), .C2(n14684), .A(n14115), .B(n20132), .ZN(
        n15992) );
  INV_X1 U17291 ( .A(n16010), .ZN(n14122) );
  NOR2_X1 U17292 ( .A1(n14122), .A2(n20132), .ZN(n16070) );
  AOI21_X1 U17293 ( .B1(n14693), .B2(n15992), .A(n16070), .ZN(n15806) );
  NAND2_X1 U17294 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n14688) );
  INV_X1 U17295 ( .A(n14688), .ZN(n14116) );
  NOR2_X1 U17296 ( .A1(n16010), .A2(n14116), .ZN(n14117) );
  OR2_X1 U17297 ( .A1(n15806), .A2(n14117), .ZN(n15982) );
  NOR2_X1 U17298 ( .A1(n20154), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14118) );
  NOR2_X1 U17299 ( .A1(n15982), .A2(n14118), .ZN(n14673) );
  INV_X1 U17300 ( .A(n16030), .ZN(n14727) );
  NAND2_X1 U17301 ( .A1(n14727), .A2(n20154), .ZN(n14120) );
  INV_X1 U17302 ( .A(n14119), .ZN(n14657) );
  AOI22_X1 U17303 ( .A1(n14120), .A2(n14653), .B1(n14716), .B2(n14657), .ZN(
        n14121) );
  NAND2_X1 U17304 ( .A1(n14673), .A2(n14121), .ZN(n14664) );
  NOR2_X1 U17305 ( .A1(n14664), .A2(n14122), .ZN(n14126) );
  INV_X1 U17306 ( .A(n14126), .ZN(n14125) );
  INV_X1 U17307 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14123) );
  NOR3_X1 U17308 ( .A1(n14664), .A2(n14123), .A3(n14497), .ZN(n14124) );
  NOR2_X1 U17309 ( .A1(n14124), .A2(n14126), .ZN(n14649) );
  AOI21_X1 U17310 ( .B1(n14636), .B2(n14125), .A(n14649), .ZN(n14631) );
  OAI211_X1 U17311 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16010), .A(
        n14631), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14621) );
  INV_X1 U17312 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14744) );
  NOR2_X1 U17313 ( .A1(n14126), .A2(n14744), .ZN(n14131) );
  NOR2_X1 U17314 ( .A1(n14688), .A2(n14686), .ZN(n14669) );
  NAND3_X1 U17315 ( .A1(n15984), .A2(n14693), .A3(n14669), .ZN(n14668) );
  NOR3_X1 U17316 ( .A1(n14668), .A2(n14653), .A3(n14497), .ZN(n14637) );
  INV_X1 U17317 ( .A(n14636), .ZN(n14128) );
  NAND3_X1 U17318 ( .A1(n14637), .A2(n14128), .A3(
        P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14620) );
  NOR3_X1 U17319 ( .A1(n14620), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n12693), .ZN(n14130) );
  AOI211_X1 U17320 ( .C1(n14621), .C2(n14131), .A(n14130), .B(n14129), .ZN(
        n14169) );
  AOI22_X1 U17321 ( .A1(n14163), .A2(P1_EBX_REG_31__SCAN_IN), .B1(n14198), 
        .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14167) );
  AOI22_X1 U17322 ( .A1(n14163), .A2(P1_EBX_REG_30__SCAN_IN), .B1(n14198), 
        .B2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14219) );
  MUX2_X1 U17323 ( .A(n14158), .B(n13423), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n14133) );
  OR2_X1 U17324 ( .A1(n14163), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n14132) );
  AND2_X1 U17325 ( .A1(n14133), .A2(n14132), .ZN(n14370) );
  NAND2_X1 U17326 ( .A1(n13427), .A2(n14134), .ZN(n14136) );
  INV_X1 U17327 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14383) );
  NAND2_X1 U17328 ( .A1(n14162), .A2(n14383), .ZN(n14135) );
  NAND3_X1 U17329 ( .A1(n14136), .A2(n13423), .A3(n14135), .ZN(n14138) );
  NAND2_X1 U17330 ( .A1(n14155), .A2(n14383), .ZN(n14137) );
  NAND2_X1 U17331 ( .A1(n14138), .A2(n14137), .ZN(n14381) );
  NAND2_X1 U17332 ( .A1(n14370), .A2(n14381), .ZN(n14139) );
  MUX2_X1 U17333 ( .A(n13423), .B(n13427), .S(P1_EBX_REG_20__SCAN_IN), .Z(
        n14141) );
  NAND2_X1 U17334 ( .A1(n14198), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14140) );
  NAND2_X1 U17335 ( .A1(n14141), .A2(n14140), .ZN(n14365) );
  MUX2_X1 U17336 ( .A(n14158), .B(n13423), .S(P1_EBX_REG_21__SCAN_IN), .Z(
        n14142) );
  OAI21_X1 U17337 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n14163), .A(
        n14142), .ZN(n14340) );
  MUX2_X1 U17338 ( .A(n13423), .B(n13427), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n14144) );
  NAND2_X1 U17339 ( .A1(n14198), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14143) );
  NAND2_X1 U17340 ( .A1(n14144), .A2(n14143), .ZN(n14321) );
  INV_X1 U17341 ( .A(n14321), .ZN(n14145) );
  MUX2_X1 U17342 ( .A(n14158), .B(n13423), .S(P1_EBX_REG_23__SCAN_IN), .Z(
        n14147) );
  OR2_X1 U17343 ( .A1(n14163), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14146) );
  AND2_X1 U17344 ( .A1(n14147), .A2(n14146), .ZN(n14310) );
  INV_X1 U17345 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14671) );
  NAND2_X1 U17346 ( .A1(n13427), .A2(n14671), .ZN(n14149) );
  INV_X1 U17347 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14361) );
  NAND2_X1 U17348 ( .A1(n14162), .A2(n14361), .ZN(n14148) );
  NAND3_X1 U17349 ( .A1(n14149), .A2(n13423), .A3(n14148), .ZN(n14151) );
  NAND2_X1 U17350 ( .A1(n14155), .A2(n14361), .ZN(n14150) );
  NAND2_X1 U17351 ( .A1(n14151), .A2(n14150), .ZN(n14295) );
  MUX2_X1 U17352 ( .A(n14158), .B(n13423), .S(P1_EBX_REG_25__SCAN_IN), .Z(
        n14152) );
  OAI21_X1 U17353 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n14163), .A(
        n14152), .ZN(n14283) );
  NAND2_X1 U17354 ( .A1(n13427), .A2(n14497), .ZN(n14154) );
  INV_X1 U17355 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14359) );
  NAND2_X1 U17356 ( .A1(n14162), .A2(n14359), .ZN(n14153) );
  NAND3_X1 U17357 ( .A1(n14154), .A2(n13423), .A3(n14153), .ZN(n14157) );
  NAND2_X1 U17358 ( .A1(n14155), .A2(n14359), .ZN(n14156) );
  AND2_X1 U17359 ( .A1(n14157), .A2(n14156), .ZN(n14265) );
  MUX2_X1 U17360 ( .A(n14158), .B(n13423), .S(P1_EBX_REG_27__SCAN_IN), .Z(
        n14159) );
  OAI21_X1 U17361 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14163), .A(
        n14159), .ZN(n14257) );
  MUX2_X1 U17362 ( .A(n13423), .B(n13427), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n14161) );
  NAND2_X1 U17363 ( .A1(n14198), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14160) );
  NAND2_X1 U17364 ( .A1(n14161), .A2(n14160), .ZN(n14244) );
  INV_X1 U17365 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14355) );
  NAND2_X1 U17366 ( .A1(n14162), .A2(n14355), .ZN(n14165) );
  OR2_X1 U17367 ( .A1(n14163), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14164) );
  NAND2_X1 U17368 ( .A1(n14164), .A2(n14165), .ZN(n14216) );
  MUX2_X1 U17369 ( .A(n14165), .B(n14216), .S(n13423), .Z(n14227) );
  MUX2_X1 U17370 ( .A(n14219), .B(n13423), .S(n14229), .Z(n14166) );
  XOR2_X1 U17371 ( .A(n14167), .B(n14166), .Z(n14350) );
  NAND2_X1 U17372 ( .A1(n14350), .A2(n20157), .ZN(n14168) );
  AOI21_X1 U17373 ( .B1(n16252), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A(
        n14170), .ZN(n14173) );
  NAND2_X1 U17374 ( .A1(n16279), .A2(n14171), .ZN(n14172) );
  OAI211_X1 U17375 ( .C1(n14174), .C2(n15182), .A(n14173), .B(n14172), .ZN(
        n14175) );
  OAI21_X1 U17376 ( .B1(n14178), .B2(n16259), .A(n14177), .ZN(P2_U2983) );
  INV_X1 U17377 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n16424) );
  AOI22_X1 U17378 ( .A1(n14468), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14462), .ZN(n14180) );
  OAI211_X1 U17379 ( .C1(n14466), .C2(n16424), .A(n14181), .B(n14180), .ZN(
        P1_U2873) );
  NOR2_X1 U17380 ( .A1(n16142), .A2(n14856), .ZN(n14182) );
  AOI21_X1 U17381 ( .B1(P2_EBX_REG_30__SCAN_IN), .B2(n14856), .A(n14182), .ZN(
        n14183) );
  OAI21_X1 U17382 ( .B1(n14184), .B2(n14865), .A(n14183), .ZN(P2_U2857) );
  INV_X1 U17383 ( .A(n14185), .ZN(n14186) );
  NAND2_X1 U17384 ( .A1(n14187), .A2(n14186), .ZN(n14189) );
  AOI22_X1 U17385 ( .A1(n14189), .A2(n14197), .B1(n12744), .B2(n14188), .ZN(
        n14190) );
  OAI21_X1 U17386 ( .B1(n14191), .B2(n14197), .A(n14190), .ZN(n14193) );
  AND2_X1 U17387 ( .A1(n14193), .A2(n14192), .ZN(n15782) );
  AOI21_X1 U17388 ( .B1(n12744), .B2(n14195), .A(n14194), .ZN(n14196) );
  AOI21_X1 U17389 ( .B1(n14197), .B2(n14199), .A(n14196), .ZN(n19910) );
  NAND3_X1 U17390 ( .A1(n14199), .A2(n14198), .A3(n15826), .ZN(n14200) );
  NAND2_X1 U17391 ( .A1(n14200), .A2(n20767), .ZN(n20759) );
  NAND2_X1 U17392 ( .A1(n19910), .A2(n20759), .ZN(n15779) );
  AND2_X1 U17393 ( .A1(n15779), .A2(n14201), .ZN(n19920) );
  MUX2_X1 U17394 ( .A(P1_MORE_REG_SCAN_IN), .B(n15782), .S(n19920), .Z(
        P1_U3484) );
  INV_X1 U17395 ( .A(n14202), .ZN(n14214) );
  NAND4_X1 U17396 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_16__SCAN_IN), 
        .A3(P1_REIP_REG_15__SCAN_IN), .A4(n14203), .ZN(n15837) );
  NAND2_X1 U17397 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(P1_REIP_REG_18__SCAN_IN), 
        .ZN(n15846) );
  NOR2_X1 U17398 ( .A1(n15837), .A2(n15846), .ZN(n14342) );
  AND3_X1 U17399 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(P1_REIP_REG_21__SCAN_IN), 
        .A3(n14341), .ZN(n14204) );
  NAND2_X1 U17400 ( .A1(n14342), .A2(n14204), .ZN(n14328) );
  NAND2_X1 U17401 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14205) );
  OR2_X1 U17402 ( .A1(n14328), .A2(n14205), .ZN(n14287) );
  INV_X1 U17403 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n14548) );
  NOR2_X1 U17404 ( .A1(n14287), .A2(n14548), .ZN(n14272) );
  AND2_X1 U17405 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .ZN(n14206) );
  AND2_X1 U17406 ( .A1(n14272), .A2(n14206), .ZN(n14247) );
  AND2_X1 U17407 ( .A1(P1_REIP_REG_27__SCAN_IN), .A2(P1_REIP_REG_28__SCAN_IN), 
        .ZN(n14207) );
  NAND2_X1 U17408 ( .A1(n14247), .A2(n14207), .ZN(n14234) );
  INV_X1 U17409 ( .A(n14234), .ZN(n14208) );
  AND2_X1 U17410 ( .A1(n20029), .A2(n14208), .ZN(n14233) );
  NAND3_X1 U17411 ( .A1(n14233), .A2(P1_REIP_REG_30__SCAN_IN), .A3(
        P1_REIP_REG_29__SCAN_IN), .ZN(n14209) );
  NAND2_X1 U17412 ( .A1(n19937), .A2(n14209), .ZN(n14220) );
  INV_X1 U17413 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n20730) );
  NOR3_X1 U17414 ( .A1(n20017), .A2(n20730), .A3(n14234), .ZN(n14222) );
  NAND3_X1 U17415 ( .A1(n14222), .A2(P1_REIP_REG_30__SCAN_IN), .A3(n20735), 
        .ZN(n14211) );
  AOI22_X1 U17416 ( .A1(n20026), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n20013), .ZN(n14210) );
  OAI211_X1 U17417 ( .C1(n14220), .C2(n20735), .A(n14211), .B(n14210), .ZN(
        n14212) );
  AOI21_X1 U17418 ( .B1(n14350), .B2(n20034), .A(n14212), .ZN(n14213) );
  OAI21_X1 U17419 ( .B1(n14214), .B2(n19942), .A(n14213), .ZN(P1_U2809) );
  INV_X1 U17420 ( .A(n14485), .ZN(n14409) );
  INV_X1 U17421 ( .A(n14229), .ZN(n14217) );
  OAI22_X1 U17422 ( .A1(n14217), .A2(n13423), .B1(n14216), .B2(n14246), .ZN(
        n14218) );
  XOR2_X1 U17423 ( .A(n14219), .B(n14218), .Z(n14353) );
  INV_X1 U17424 ( .A(n14353), .ZN(n14619) );
  INV_X1 U17425 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14354) );
  INV_X1 U17426 ( .A(n14220), .ZN(n14221) );
  OAI21_X1 U17427 ( .B1(n14222), .B2(P1_REIP_REG_30__SCAN_IN), .A(n14221), 
        .ZN(n14224) );
  AOI22_X1 U17428 ( .A1(n14481), .A2(n20014), .B1(n20013), .B2(
        P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14223) );
  OAI211_X1 U17429 ( .C1(n19991), .C2(n14354), .A(n14224), .B(n14223), .ZN(
        n14225) );
  AOI21_X1 U17430 ( .B1(n14619), .B2(n20034), .A(n14225), .ZN(n14226) );
  OAI21_X1 U17431 ( .B1(n14409), .B2(n19942), .A(n14226), .ZN(P1_U2810) );
  NAND2_X1 U17432 ( .A1(n14246), .A2(n14227), .ZN(n14228) );
  NAND2_X1 U17433 ( .A1(n14229), .A2(n14228), .ZN(n14626) );
  NAND2_X1 U17434 ( .A1(n14493), .A2(n19978), .ZN(n14240) );
  NOR2_X1 U17435 ( .A1(n15899), .A2(n14233), .ZN(n14248) );
  NOR3_X1 U17436 ( .A1(n20017), .A2(P1_REIP_REG_29__SCAN_IN), .A3(n14234), 
        .ZN(n14238) );
  INV_X1 U17437 ( .A(n14491), .ZN(n14235) );
  AOI22_X1 U17438 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n20013), .B1(
        n20014), .B2(n14235), .ZN(n14236) );
  OAI21_X1 U17439 ( .B1(n19991), .B2(n14355), .A(n14236), .ZN(n14237) );
  AOI211_X1 U17440 ( .C1(n14248), .C2(P1_REIP_REG_29__SCAN_IN), .A(n14238), 
        .B(n14237), .ZN(n14239) );
  OAI211_X1 U17441 ( .C1(n20008), .C2(n14626), .A(n14240), .B(n14239), .ZN(
        P1_U2811) );
  OAI21_X1 U17443 ( .B1(n14242), .B2(n14243), .A(n14230), .ZN(n14504) );
  OR2_X1 U17444 ( .A1(n14256), .A2(n14244), .ZN(n14245) );
  NAND2_X1 U17445 ( .A1(n14246), .A2(n14245), .ZN(n14356) );
  INV_X1 U17446 ( .A(n14356), .ZN(n14640) );
  INV_X1 U17447 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14357) );
  INV_X1 U17448 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n20724) );
  INV_X1 U17449 ( .A(n14247), .ZN(n14259) );
  NOR3_X1 U17450 ( .A1(n20017), .A2(n20724), .A3(n14259), .ZN(n14249) );
  OAI21_X1 U17451 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(n14249), .A(n14248), 
        .ZN(n14251) );
  AOI22_X1 U17452 ( .A1(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n20013), .B1(
        n20014), .B2(n14505), .ZN(n14250) );
  OAI211_X1 U17453 ( .C1(n14357), .C2(n19991), .A(n14251), .B(n14250), .ZN(
        n14252) );
  AOI21_X1 U17454 ( .B1(n14640), .B2(n20034), .A(n14252), .ZN(n14253) );
  OAI21_X1 U17455 ( .B1(n14504), .B2(n19942), .A(n14253), .ZN(P1_U2812) );
  AOI21_X1 U17456 ( .B1(n14255), .B2(n14254), .A(n14242), .ZN(n14522) );
  INV_X1 U17457 ( .A(n14522), .ZN(n14424) );
  AOI21_X1 U17458 ( .B1(n14257), .B2(n14267), .A(n14256), .ZN(n14645) );
  INV_X1 U17459 ( .A(n20029), .ZN(n20003) );
  OAI21_X1 U17460 ( .B1(n20003), .B2(n14259), .A(n19937), .ZN(n14273) );
  OAI22_X1 U17461 ( .A1(n14258), .A2(n20031), .B1(n20042), .B2(n14520), .ZN(
        n14261) );
  NOR3_X1 U17462 ( .A1(n20017), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n14259), 
        .ZN(n14260) );
  AOI211_X1 U17463 ( .C1(P1_EBX_REG_27__SCAN_IN), .C2(n20026), .A(n14261), .B(
        n14260), .ZN(n14262) );
  OAI21_X1 U17464 ( .B1(n20724), .B2(n14273), .A(n14262), .ZN(n14263) );
  AOI21_X1 U17465 ( .B1(n14645), .B2(n20034), .A(n14263), .ZN(n14264) );
  OAI21_X1 U17466 ( .B1(n14424), .B2(n19942), .A(n14264), .ZN(P1_U2813) );
  NAND2_X1 U17467 ( .A1(n14281), .A2(n14265), .ZN(n14266) );
  NAND2_X1 U17468 ( .A1(n14267), .A2(n14266), .ZN(n14652) );
  OAI21_X1 U17469 ( .B1(n14268), .B2(n14269), .A(n14254), .ZN(n14428) );
  INV_X1 U17470 ( .A(n14428), .ZN(n14533) );
  NAND2_X1 U17471 ( .A1(n14533), .A2(n19978), .ZN(n14278) );
  INV_X1 U17472 ( .A(n14270), .ZN(n14531) );
  OAI22_X1 U17473 ( .A1(n14271), .A2(n20031), .B1(n20042), .B2(n14531), .ZN(
        n14276) );
  AND2_X1 U17474 ( .A1(n20019), .A2(n14272), .ZN(n14284) );
  AOI21_X1 U17475 ( .B1(n14284), .B2(P1_REIP_REG_25__SCAN_IN), .A(
        P1_REIP_REG_26__SCAN_IN), .ZN(n14274) );
  NOR2_X1 U17476 ( .A1(n14274), .A2(n14273), .ZN(n14275) );
  AOI211_X1 U17477 ( .C1(P1_EBX_REG_26__SCAN_IN), .C2(n20026), .A(n14276), .B(
        n14275), .ZN(n14277) );
  OAI211_X1 U17478 ( .C1(n20008), .C2(n14652), .A(n14278), .B(n14277), .ZN(
        P1_U2814) );
  AOI21_X1 U17479 ( .B1(n14280), .B2(n14279), .A(n14268), .ZN(n14542) );
  INV_X1 U17480 ( .A(n14542), .ZN(n14432) );
  INV_X1 U17481 ( .A(n14281), .ZN(n14282) );
  AOI21_X1 U17482 ( .B1(n14283), .B2(n14297), .A(n14282), .ZN(n14663) );
  INV_X1 U17483 ( .A(n14284), .ZN(n14292) );
  OAI22_X1 U17484 ( .A1(n14285), .A2(n20031), .B1(n20042), .B2(n14540), .ZN(
        n14286) );
  AOI21_X1 U17485 ( .B1(n20026), .B2(P1_EBX_REG_25__SCAN_IN), .A(n14286), .ZN(
        n14291) );
  INV_X1 U17486 ( .A(n14287), .ZN(n14300) );
  OR2_X1 U17487 ( .A1(n20017), .A2(n14300), .ZN(n14288) );
  NAND2_X1 U17488 ( .A1(n14288), .A2(n20029), .ZN(n14313) );
  NOR2_X1 U17489 ( .A1(n20017), .A2(P1_REIP_REG_24__SCAN_IN), .ZN(n14289) );
  OAI21_X1 U17490 ( .B1(n14313), .B2(n14289), .A(P1_REIP_REG_25__SCAN_IN), 
        .ZN(n14290) );
  OAI211_X1 U17491 ( .C1(n14292), .C2(P1_REIP_REG_25__SCAN_IN), .A(n14291), 
        .B(n14290), .ZN(n14293) );
  AOI21_X1 U17492 ( .B1(n14663), .B2(n20034), .A(n14293), .ZN(n14294) );
  OAI21_X1 U17493 ( .B1(n14432), .B2(n19942), .A(n14294), .ZN(P1_U2815) );
  OR2_X1 U17494 ( .A1(n14312), .A2(n14295), .ZN(n14296) );
  NAND2_X1 U17495 ( .A1(n14297), .A2(n14296), .ZN(n14674) );
  OAI21_X1 U17496 ( .B1(n14298), .B2(n14299), .A(n14279), .ZN(n14436) );
  INV_X1 U17497 ( .A(n14436), .ZN(n14552) );
  NAND2_X1 U17498 ( .A1(n14552), .A2(n19978), .ZN(n14306) );
  NAND2_X1 U17499 ( .A1(n14300), .A2(n14548), .ZN(n14303) );
  NAND2_X1 U17500 ( .A1(n20026), .A2(P1_EBX_REG_24__SCAN_IN), .ZN(n14302) );
  AOI22_X1 U17501 ( .A1(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n20013), .B1(
        n20014), .B2(n14547), .ZN(n14301) );
  OAI211_X1 U17502 ( .C1(n14303), .C2(n20017), .A(n14302), .B(n14301), .ZN(
        n14304) );
  AOI21_X1 U17503 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n14313), .A(n14304), 
        .ZN(n14305) );
  OAI211_X1 U17504 ( .C1(n20008), .C2(n14674), .A(n14306), .B(n14305), .ZN(
        P1_U2816) );
  AOI21_X1 U17505 ( .B1(n14308), .B2(n14307), .A(n14298), .ZN(n14309) );
  INV_X1 U17506 ( .A(n14309), .ZN(n14556) );
  NOR2_X1 U17507 ( .A1(n14319), .A2(n14310), .ZN(n14311) );
  OR2_X1 U17508 ( .A1(n14312), .A2(n14311), .ZN(n14363) );
  INV_X1 U17509 ( .A(n14363), .ZN(n15986) );
  INV_X1 U17510 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14362) );
  INV_X1 U17511 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n14565) );
  NOR3_X1 U17512 ( .A1(n20017), .A2(n14328), .A3(n14565), .ZN(n14314) );
  OAI21_X1 U17513 ( .B1(n14314), .B2(P1_REIP_REG_23__SCAN_IN), .A(n14313), 
        .ZN(n14316) );
  AOI22_X1 U17514 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n20013), .B1(
        n20014), .B2(n14559), .ZN(n14315) );
  OAI211_X1 U17515 ( .C1(n14362), .C2(n19991), .A(n14316), .B(n14315), .ZN(
        n14317) );
  AOI21_X1 U17516 ( .B1(n15986), .B2(n20034), .A(n14317), .ZN(n14318) );
  OAI21_X1 U17517 ( .B1(n14556), .B2(n19942), .A(n14318), .ZN(P1_U2817) );
  INV_X1 U17518 ( .A(n14319), .ZN(n14320) );
  OAI21_X1 U17519 ( .B1(n9665), .B2(n14321), .A(n14320), .ZN(n14681) );
  INV_X1 U17520 ( .A(n14307), .ZN(n14324) );
  AOI21_X1 U17521 ( .B1(n14325), .B2(n14323), .A(n14324), .ZN(n14569) );
  NAND2_X1 U17522 ( .A1(n14569), .A2(n19978), .ZN(n14336) );
  INV_X1 U17523 ( .A(n14342), .ZN(n14326) );
  INV_X1 U17524 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n20713) );
  NOR3_X1 U17525 ( .A1(n19936), .A2(n14326), .A3(n20713), .ZN(n14327) );
  NOR2_X1 U17526 ( .A1(n15899), .A2(n14327), .ZN(n15842) );
  INV_X1 U17527 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n14333) );
  INV_X1 U17528 ( .A(n14328), .ZN(n14330) );
  NAND2_X1 U17529 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_22__SCAN_IN), 
        .ZN(n14329) );
  OAI211_X1 U17530 ( .C1(n14330), .C2(P1_REIP_REG_22__SCAN_IN), .A(n20019), 
        .B(n14329), .ZN(n14332) );
  AOI22_X1 U17531 ( .A1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n20013), .B1(
        n20014), .B2(n14564), .ZN(n14331) );
  OAI211_X1 U17532 ( .C1(n19991), .C2(n14333), .A(n14332), .B(n14331), .ZN(
        n14334) );
  AOI21_X1 U17533 ( .B1(n15842), .B2(P1_REIP_REG_22__SCAN_IN), .A(n14334), 
        .ZN(n14335) );
  OAI211_X1 U17534 ( .C1(n14681), .C2(n20008), .A(n14336), .B(n14335), .ZN(
        P1_U2818) );
  OAI21_X1 U17535 ( .B1(n14338), .B2(n14339), .A(n14323), .ZN(n15905) );
  AOI21_X1 U17536 ( .B1(n14340), .B2(n9709), .A(n9665), .ZN(n15813) );
  INV_X1 U17537 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n20716) );
  NAND4_X1 U17538 ( .A1(n14342), .A2(P1_REIP_REG_20__SCAN_IN), .A3(n14341), 
        .A4(n20716), .ZN(n14347) );
  NAND2_X1 U17539 ( .A1(n15842), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14346) );
  INV_X1 U17540 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n14343) );
  OAI22_X1 U17541 ( .A1(n14343), .A2(n20031), .B1(n20042), .B2(n15910), .ZN(
        n14344) );
  AOI21_X1 U17542 ( .B1(n20026), .B2(P1_EBX_REG_21__SCAN_IN), .A(n14344), .ZN(
        n14345) );
  OAI211_X1 U17543 ( .C1(n20017), .C2(n14347), .A(n14346), .B(n14345), .ZN(
        n14348) );
  AOI21_X1 U17544 ( .B1(n15813), .B2(n20034), .A(n14348), .ZN(n14349) );
  OAI21_X1 U17545 ( .B1(n15905), .B2(n19942), .A(n14349), .ZN(P1_U2819) );
  INV_X1 U17546 ( .A(n14350), .ZN(n14352) );
  INV_X1 U17547 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14351) );
  OAI22_X1 U17548 ( .A1(n14352), .A2(n14379), .B1(n14351), .B2(n14377), .ZN(
        P1_U2841) );
  OAI222_X1 U17549 ( .A1(n14387), .A2(n14409), .B1(n14384), .B2(n14354), .C1(
        n14353), .C2(n14379), .ZN(P1_U2842) );
  INV_X1 U17550 ( .A(n14493), .ZN(n14416) );
  OAI222_X1 U17551 ( .A1(n14355), .A2(n14384), .B1(n14379), .B2(n14626), .C1(
        n14416), .C2(n14387), .ZN(P1_U2843) );
  OAI222_X1 U17552 ( .A1(n14357), .A2(n14384), .B1(n14379), .B2(n14356), .C1(
        n14504), .C2(n14405), .ZN(P1_U2844) );
  AOI22_X1 U17553 ( .A1(n14645), .A2(n14403), .B1(n14402), .B2(
        P1_EBX_REG_27__SCAN_IN), .ZN(n14358) );
  OAI21_X1 U17554 ( .B1(n14424), .B2(n14405), .A(n14358), .ZN(P1_U2845) );
  OAI222_X1 U17555 ( .A1(n14359), .A2(n14377), .B1(n14379), .B2(n14652), .C1(
        n14428), .C2(n14387), .ZN(P1_U2846) );
  AOI22_X1 U17556 ( .A1(n14663), .A2(n14403), .B1(n14402), .B2(
        P1_EBX_REG_25__SCAN_IN), .ZN(n14360) );
  OAI21_X1 U17557 ( .B1(n14432), .B2(n14405), .A(n14360), .ZN(P1_U2847) );
  OAI222_X1 U17558 ( .A1(n14361), .A2(n14384), .B1(n14379), .B2(n14674), .C1(
        n14436), .C2(n14387), .ZN(P1_U2848) );
  OAI222_X1 U17559 ( .A1(n14363), .A2(n14379), .B1(n14362), .B2(n14377), .C1(
        n14556), .C2(n14387), .ZN(P1_U2849) );
  INV_X1 U17560 ( .A(n14569), .ZN(n14446) );
  OAI222_X1 U17561 ( .A1(n14681), .A2(n14379), .B1(n14384), .B2(n14333), .C1(
        n14387), .C2(n14446), .ZN(P1_U2850) );
  AOI22_X1 U17562 ( .A1(n15813), .A2(n14403), .B1(n14402), .B2(
        P1_EBX_REG_21__SCAN_IN), .ZN(n14364) );
  OAI21_X1 U17563 ( .B1(n15905), .B2(n14405), .A(n14364), .ZN(P1_U2851) );
  OR2_X1 U17564 ( .A1(n14372), .A2(n14365), .ZN(n14366) );
  NAND2_X1 U17565 ( .A1(n9709), .A2(n14366), .ZN(n15838) );
  INV_X1 U17566 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n14369) );
  AOI21_X1 U17567 ( .B1(n14367), .B2(n9686), .A(n14338), .ZN(n14368) );
  INV_X1 U17568 ( .A(n14368), .ZN(n15839) );
  OAI222_X1 U17569 ( .A1(n15838), .A2(n14379), .B1(n14384), .B2(n14369), .C1(
        n14387), .C2(n15839), .ZN(P1_U2852) );
  AOI21_X1 U17570 ( .B1(n14371), .B2(n14381), .A(n14370), .ZN(n14373) );
  OR2_X1 U17571 ( .A1(n14373), .A2(n14372), .ZN(n15994) );
  INV_X1 U17572 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n14378) );
  NAND2_X1 U17573 ( .A1(n14375), .A2(n14374), .ZN(n14376) );
  NAND2_X1 U17574 ( .A1(n9686), .A2(n14376), .ZN(n15914) );
  OAI222_X1 U17575 ( .A1(n15994), .A2(n14379), .B1(n14378), .B2(n14377), .C1(
        n15914), .C2(n14387), .ZN(P1_U2853) );
  XOR2_X1 U17576 ( .A(n14380), .B(n13865), .Z(n15860) );
  INV_X1 U17577 ( .A(n15860), .ZN(n14470) );
  XNOR2_X1 U17578 ( .A(n14382), .B(n14381), .ZN(n15859) );
  NOR2_X1 U17579 ( .A1(n14384), .A2(n14383), .ZN(n14385) );
  AOI21_X1 U17580 ( .B1(n15859), .B2(n14403), .A(n14385), .ZN(n14386) );
  OAI21_X1 U17581 ( .B1(n14470), .B2(n14387), .A(n14386), .ZN(P1_U2854) );
  INV_X1 U17582 ( .A(n13834), .ZN(n14388) );
  AOI21_X1 U17583 ( .B1(n14390), .B2(n14389), .A(n14388), .ZN(n15935) );
  INV_X1 U17584 ( .A(n15935), .ZN(n14472) );
  AOI21_X1 U17585 ( .B1(n14393), .B2(n14392), .A(n14391), .ZN(n16015) );
  AOI22_X1 U17586 ( .A1(n16015), .A2(n14403), .B1(n14402), .B2(
        P1_EBX_REG_15__SCAN_IN), .ZN(n14394) );
  OAI21_X1 U17587 ( .B1(n14472), .B2(n14405), .A(n14394), .ZN(P1_U2857) );
  INV_X1 U17588 ( .A(n14395), .ZN(n14396) );
  AOI21_X1 U17589 ( .B1(n14397), .B2(n13793), .A(n14396), .ZN(n15946) );
  INV_X1 U17590 ( .A(n15946), .ZN(n14477) );
  INV_X1 U17591 ( .A(n14398), .ZN(n14399) );
  AOI21_X1 U17592 ( .B1(n14401), .B2(n14400), .A(n14399), .ZN(n15877) );
  AOI22_X1 U17593 ( .A1(n15877), .A2(n14403), .B1(n14402), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14404) );
  OAI21_X1 U17594 ( .B1(n14477), .B2(n14405), .A(n14404), .ZN(P1_U2859) );
  OAI22_X1 U17595 ( .A1(n14461), .A2(n20086), .B1(n12968), .B2(n14473), .ZN(
        n14406) );
  AOI21_X1 U17596 ( .B1(BUF1_REG_30__SCAN_IN), .B2(n14458), .A(n14406), .ZN(
        n14408) );
  NAND2_X1 U17597 ( .A1(n14468), .A2(DATAI_30_), .ZN(n14407) );
  OAI211_X1 U17598 ( .C1(n14409), .C2(n14476), .A(n14408), .B(n14407), .ZN(
        P1_U2874) );
  INV_X1 U17599 ( .A(DATAI_13_), .ZN(n14412) );
  INV_X1 U17600 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n14411) );
  MUX2_X1 U17601 ( .A(n14412), .B(n14411), .S(n14410), .Z(n20083) );
  OAI22_X1 U17602 ( .A1(n14461), .A2(n20083), .B1(n12974), .B2(n14179), .ZN(
        n14413) );
  AOI21_X1 U17603 ( .B1(BUF1_REG_29__SCAN_IN), .B2(n14458), .A(n14413), .ZN(
        n14415) );
  NAND2_X1 U17604 ( .A1(n14468), .A2(DATAI_29_), .ZN(n14414) );
  OAI211_X1 U17605 ( .C1(n14416), .C2(n14476), .A(n14415), .B(n14414), .ZN(
        P1_U2875) );
  OAI22_X1 U17606 ( .A1(n14461), .A2(n20080), .B1(n12978), .B2(n14179), .ZN(
        n14417) );
  AOI21_X1 U17607 ( .B1(BUF1_REG_28__SCAN_IN), .B2(n14458), .A(n14417), .ZN(
        n14419) );
  NAND2_X1 U17608 ( .A1(n14468), .A2(DATAI_28_), .ZN(n14418) );
  OAI211_X1 U17609 ( .C1(n14504), .C2(n14476), .A(n14419), .B(n14418), .ZN(
        P1_U2876) );
  OAI22_X1 U17610 ( .A1(n14461), .A2(n14420), .B1(n12976), .B2(n14179), .ZN(
        n14421) );
  AOI21_X1 U17611 ( .B1(BUF1_REG_27__SCAN_IN), .B2(n14458), .A(n14421), .ZN(
        n14423) );
  NAND2_X1 U17612 ( .A1(n14468), .A2(DATAI_27_), .ZN(n14422) );
  OAI211_X1 U17613 ( .C1(n14424), .C2(n14476), .A(n14423), .B(n14422), .ZN(
        P1_U2877) );
  OAI22_X1 U17614 ( .A1(n14461), .A2(n20077), .B1(n12970), .B2(n14179), .ZN(
        n14425) );
  AOI21_X1 U17615 ( .B1(BUF1_REG_26__SCAN_IN), .B2(n14458), .A(n14425), .ZN(
        n14427) );
  NAND2_X1 U17616 ( .A1(n14468), .A2(DATAI_26_), .ZN(n14426) );
  OAI211_X1 U17617 ( .C1(n14428), .C2(n14476), .A(n14427), .B(n14426), .ZN(
        P1_U2878) );
  OAI22_X1 U17618 ( .A1(n14461), .A2(n20072), .B1(n12972), .B2(n14473), .ZN(
        n14429) );
  AOI21_X1 U17619 ( .B1(n14458), .B2(BUF1_REG_25__SCAN_IN), .A(n14429), .ZN(
        n14431) );
  NAND2_X1 U17620 ( .A1(n14468), .A2(DATAI_25_), .ZN(n14430) );
  OAI211_X1 U17621 ( .C1(n14432), .C2(n14476), .A(n14431), .B(n14430), .ZN(
        P1_U2879) );
  OAI22_X1 U17622 ( .A1(n14461), .A2(n20069), .B1(n12966), .B2(n14179), .ZN(
        n14433) );
  AOI21_X1 U17623 ( .B1(n14458), .B2(BUF1_REG_24__SCAN_IN), .A(n14433), .ZN(
        n14435) );
  NAND2_X1 U17624 ( .A1(n14468), .A2(DATAI_24_), .ZN(n14434) );
  OAI211_X1 U17625 ( .C1(n14436), .C2(n14476), .A(n14435), .B(n14434), .ZN(
        P1_U2880) );
  OAI22_X1 U17626 ( .A1(n14461), .A2(n14438), .B1(n14437), .B2(n14473), .ZN(
        n14439) );
  AOI21_X1 U17627 ( .B1(n14458), .B2(BUF1_REG_23__SCAN_IN), .A(n14439), .ZN(
        n14441) );
  NAND2_X1 U17628 ( .A1(n14468), .A2(DATAI_23_), .ZN(n14440) );
  OAI211_X1 U17629 ( .C1(n14556), .C2(n14476), .A(n14441), .B(n14440), .ZN(
        P1_U2881) );
  OAI22_X1 U17630 ( .A1(n14461), .A2(n14442), .B1(n13132), .B2(n14473), .ZN(
        n14443) );
  AOI21_X1 U17631 ( .B1(n14458), .B2(BUF1_REG_22__SCAN_IN), .A(n14443), .ZN(
        n14445) );
  NAND2_X1 U17632 ( .A1(n14468), .A2(DATAI_22_), .ZN(n14444) );
  OAI211_X1 U17633 ( .C1(n14446), .C2(n14476), .A(n14445), .B(n14444), .ZN(
        P1_U2882) );
  OAI22_X1 U17634 ( .A1(n14461), .A2(n14447), .B1(n13129), .B2(n14179), .ZN(
        n14448) );
  AOI21_X1 U17635 ( .B1(n14458), .B2(BUF1_REG_21__SCAN_IN), .A(n14448), .ZN(
        n14450) );
  NAND2_X1 U17636 ( .A1(n14468), .A2(DATAI_21_), .ZN(n14449) );
  OAI211_X1 U17637 ( .C1(n15905), .C2(n14476), .A(n14450), .B(n14449), .ZN(
        P1_U2883) );
  OAI22_X1 U17638 ( .A1(n14461), .A2(n14451), .B1(n13137), .B2(n14473), .ZN(
        n14452) );
  AOI21_X1 U17639 ( .B1(n14458), .B2(BUF1_REG_20__SCAN_IN), .A(n14452), .ZN(
        n14454) );
  NAND2_X1 U17640 ( .A1(n14468), .A2(DATAI_20_), .ZN(n14453) );
  OAI211_X1 U17641 ( .C1(n15839), .C2(n14476), .A(n14454), .B(n14453), .ZN(
        P1_U2884) );
  INV_X1 U17642 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n14455) );
  OAI22_X1 U17643 ( .A1(n14461), .A2(n14456), .B1(n14455), .B2(n14473), .ZN(
        n14457) );
  AOI21_X1 U17644 ( .B1(n14458), .B2(BUF1_REG_19__SCAN_IN), .A(n14457), .ZN(
        n14460) );
  NAND2_X1 U17645 ( .A1(n14468), .A2(DATAI_19_), .ZN(n14459) );
  OAI211_X1 U17646 ( .C1(n15914), .C2(n14476), .A(n14460), .B(n14459), .ZN(
        P1_U2885) );
  INV_X1 U17647 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n16446) );
  INV_X1 U17648 ( .A(n14461), .ZN(n14464) );
  AOI22_X1 U17649 ( .A1(n14464), .A2(n14463), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n14462), .ZN(n14465) );
  OAI21_X1 U17650 ( .B1(n16446), .B2(n14466), .A(n14465), .ZN(n14467) );
  AOI21_X1 U17651 ( .B1(n14468), .B2(DATAI_18_), .A(n14467), .ZN(n14469) );
  OAI21_X1 U17652 ( .B1(n14470), .B2(n14476), .A(n14469), .ZN(P1_U2886) );
  OAI222_X1 U17653 ( .A1(n14472), .A2(n14476), .B1(n14471), .B2(n14475), .C1(
        n14473), .C2(n12986), .ZN(P1_U2889) );
  INV_X1 U17654 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n14474) );
  OAI222_X1 U17655 ( .A1(n14477), .A2(n14476), .B1(n20083), .B2(n14475), .C1(
        n14474), .C2(n14473), .ZN(P1_U2891) );
  NAND2_X1 U17656 ( .A1(n14479), .A2(n14478), .ZN(n14480) );
  XNOR2_X1 U17657 ( .A(n14480), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14625) );
  NAND2_X1 U17658 ( .A1(n15961), .A2(n14481), .ZN(n14482) );
  NAND2_X1 U17659 ( .A1(n20162), .A2(P1_REIP_REG_30__SCAN_IN), .ZN(n14617) );
  OAI211_X1 U17660 ( .C1(n14483), .C2(n14580), .A(n14482), .B(n14617), .ZN(
        n14484) );
  AOI21_X1 U17661 ( .B1(n14485), .B2(n20125), .A(n14484), .ZN(n14486) );
  OAI21_X1 U17662 ( .B1(n14625), .B2(n19918), .A(n14486), .ZN(P1_U2969) );
  NOR2_X1 U17663 ( .A1(n14488), .A2(n14487), .ZN(n14489) );
  XNOR2_X1 U17664 ( .A(n14489), .B(n14630), .ZN(n14634) );
  NOR2_X1 U17665 ( .A1(n20135), .A2(n20730), .ZN(n14628) );
  AOI21_X1 U17666 ( .B1(n20120), .B2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14628), .ZN(n14490) );
  OAI21_X1 U17667 ( .B1(n20130), .B2(n14491), .A(n14490), .ZN(n14492) );
  AOI21_X1 U17668 ( .B1(n14493), .B2(n20125), .A(n14492), .ZN(n14494) );
  OAI21_X1 U17669 ( .B1(n14634), .B2(n19918), .A(n14494), .ZN(P1_U2970) );
  INV_X1 U17670 ( .A(n14653), .ZN(n14525) );
  OAI21_X1 U17671 ( .B1(n9985), .B2(n14525), .A(n14495), .ZN(n14501) );
  INV_X1 U17672 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15990) );
  NAND3_X1 U17673 ( .A1(n14496), .A2(n15990), .A3(n14497), .ZN(n14499) );
  MUX2_X1 U17674 ( .A(n14497), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .S(
        n9985), .Z(n14498) );
  AOI21_X1 U17675 ( .B1(n14501), .B2(n14499), .A(n14498), .ZN(n14500) );
  OAI21_X1 U17676 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14501), .A(
        n14500), .ZN(n14503) );
  XNOR2_X1 U17677 ( .A(n14503), .B(n14502), .ZN(n14643) );
  INV_X1 U17678 ( .A(n14504), .ZN(n14510) );
  INV_X1 U17679 ( .A(n14505), .ZN(n14508) );
  INV_X1 U17680 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14506) );
  NOR2_X1 U17681 ( .A1(n20135), .A2(n14506), .ZN(n14639) );
  AOI21_X1 U17682 ( .B1(n20120), .B2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n14639), .ZN(n14507) );
  OAI21_X1 U17683 ( .B1(n20130), .B2(n14508), .A(n14507), .ZN(n14509) );
  AOI21_X1 U17684 ( .B1(n14510), .B2(n20125), .A(n14509), .ZN(n14511) );
  OAI21_X1 U17685 ( .B1(n19918), .B2(n14643), .A(n14511), .ZN(P1_U2971) );
  INV_X1 U17686 ( .A(n14512), .ZN(n14513) );
  NAND2_X1 U17687 ( .A1(n14514), .A2(n14513), .ZN(n14516) );
  MUX2_X1 U17688 ( .A(n14516), .B(n14515), .S(n9985), .Z(n14518) );
  XNOR2_X1 U17689 ( .A(n14518), .B(n14517), .ZN(n14651) );
  NOR2_X1 U17690 ( .A1(n20135), .A2(n20724), .ZN(n14644) );
  AOI21_X1 U17691 ( .B1(n20120), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14644), .ZN(n14519) );
  OAI21_X1 U17692 ( .B1(n20130), .B2(n14520), .A(n14519), .ZN(n14521) );
  AOI21_X1 U17693 ( .B1(n14522), .B2(n20125), .A(n14521), .ZN(n14523) );
  OAI21_X1 U17694 ( .B1(n19918), .B2(n14651), .A(n14523), .ZN(P1_U2972) );
  INV_X1 U17695 ( .A(n14524), .ZN(n14527) );
  AOI21_X1 U17696 ( .B1(n14495), .B2(n14525), .A(n15808), .ZN(n14526) );
  NOR2_X1 U17697 ( .A1(n14527), .A2(n14526), .ZN(n14528) );
  XNOR2_X1 U17698 ( .A(n14528), .B(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14660) );
  INV_X1 U17699 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n14529) );
  NOR2_X1 U17700 ( .A1(n20135), .A2(n14529), .ZN(n14655) );
  AOI21_X1 U17701 ( .B1(n20120), .B2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A(
        n14655), .ZN(n14530) );
  OAI21_X1 U17702 ( .B1(n20130), .B2(n14531), .A(n14530), .ZN(n14532) );
  AOI21_X1 U17703 ( .B1(n14533), .B2(n20125), .A(n14532), .ZN(n14534) );
  OAI21_X1 U17704 ( .B1(n19918), .B2(n14660), .A(n14534), .ZN(P1_U2973) );
  MUX2_X1 U17705 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n14536), .S(
        n9985), .Z(n14537) );
  OAI21_X1 U17706 ( .B1(n14544), .B2(n14671), .A(n14537), .ZN(n14538) );
  XOR2_X1 U17707 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B(n14538), .Z(
        n14667) );
  INV_X1 U17708 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n20722) );
  NOR2_X1 U17709 ( .A1(n20135), .A2(n20722), .ZN(n14662) );
  AOI21_X1 U17710 ( .B1(n20120), .B2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .A(
        n14662), .ZN(n14539) );
  OAI21_X1 U17711 ( .B1(n20130), .B2(n14540), .A(n14539), .ZN(n14541) );
  AOI21_X1 U17712 ( .B1(n14542), .B2(n20125), .A(n14541), .ZN(n14543) );
  OAI21_X1 U17713 ( .B1(n19918), .B2(n14667), .A(n14543), .ZN(P1_U2974) );
  NOR2_X1 U17714 ( .A1(n14544), .A2(n14495), .ZN(n14545) );
  MUX2_X1 U17715 ( .A(n14545), .B(n14544), .S(n15955), .Z(n14546) );
  XNOR2_X1 U17716 ( .A(n14546), .B(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14680) );
  INV_X1 U17717 ( .A(n14547), .ZN(n14550) );
  NOR2_X1 U17718 ( .A1(n20135), .A2(n14548), .ZN(n14675) );
  AOI21_X1 U17719 ( .B1(n20120), .B2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n14675), .ZN(n14549) );
  OAI21_X1 U17720 ( .B1(n20130), .B2(n14550), .A(n14549), .ZN(n14551) );
  AOI21_X1 U17721 ( .B1(n14552), .B2(n20125), .A(n14551), .ZN(n14553) );
  OAI21_X1 U17722 ( .B1(n19918), .B2(n14680), .A(n14553), .ZN(P1_U2975) );
  XNOR2_X1 U17723 ( .A(n15808), .B(n15990), .ZN(n14554) );
  XNOR2_X1 U17724 ( .A(n14495), .B(n14554), .ZN(n15985) );
  INV_X1 U17725 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n20718) );
  NAND2_X1 U17726 ( .A1(n20120), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14555) );
  OAI21_X1 U17727 ( .B1(n20718), .B2(n20135), .A(n14555), .ZN(n14558) );
  NOR2_X1 U17728 ( .A1(n14556), .A2(n14616), .ZN(n14557) );
  AOI211_X1 U17729 ( .C1(n15961), .C2(n14559), .A(n14558), .B(n14557), .ZN(
        n14560) );
  OAI21_X1 U17730 ( .B1(n15985), .B2(n19918), .A(n14560), .ZN(P1_U2976) );
  NAND2_X1 U17731 ( .A1(n14562), .A2(n14561), .ZN(n14563) );
  XOR2_X1 U17732 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B(n14563), .Z(
        n14692) );
  INV_X1 U17733 ( .A(n14564), .ZN(n14567) );
  NOR2_X1 U17734 ( .A1(n20135), .A2(n14565), .ZN(n14683) );
  AOI21_X1 U17735 ( .B1(n20120), .B2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .A(
        n14683), .ZN(n14566) );
  OAI21_X1 U17736 ( .B1(n20130), .B2(n14567), .A(n14566), .ZN(n14568) );
  AOI21_X1 U17737 ( .B1(n14569), .B2(n20125), .A(n14568), .ZN(n14570) );
  OAI21_X1 U17738 ( .B1(n19918), .B2(n14692), .A(n14570), .ZN(P1_U2977) );
  NOR4_X1 U17739 ( .A1(n12689), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A4(n15955), .ZN(n15811) );
  NOR3_X1 U17740 ( .A1(n9985), .A2(n14571), .A3(n15912), .ZN(n14572) );
  OR2_X1 U17741 ( .A1(n15811), .A2(n14572), .ZN(n14573) );
  XOR2_X1 U17742 ( .A(n14573), .B(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .Z(
        n14700) );
  AOI22_X1 U17743 ( .A1(n12697), .A2(n14700), .B1(n20162), .B2(
        P1_REIP_REG_20__SCAN_IN), .ZN(n14574) );
  OAI21_X1 U17744 ( .B1(n14580), .B2(n15845), .A(n14574), .ZN(n14575) );
  AOI21_X1 U17745 ( .B1(n15961), .B2(n15836), .A(n14575), .ZN(n14576) );
  OAI21_X1 U17746 ( .B1(n15839), .B2(n14616), .A(n14576), .ZN(P1_U2979) );
  OAI21_X1 U17747 ( .B1(n12689), .B2(n14577), .A(n14571), .ZN(n14711) );
  NAND2_X1 U17748 ( .A1(n15855), .A2(n15961), .ZN(n14578) );
  NAND2_X1 U17749 ( .A1(n20162), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n14704) );
  OAI211_X1 U17750 ( .C1(n14580), .C2(n14579), .A(n14578), .B(n14704), .ZN(
        n14581) );
  AOI21_X1 U17751 ( .B1(n15860), .B2(n20125), .A(n14581), .ZN(n14582) );
  OAI21_X1 U17752 ( .B1(n19918), .B2(n14711), .A(n14582), .ZN(P1_U2981) );
  OAI21_X1 U17753 ( .B1(n15956), .B2(n14584), .A(n14583), .ZN(n15933) );
  NOR3_X1 U17754 ( .A1(n15933), .A2(n14585), .A3(n15929), .ZN(n15931) );
  NOR2_X1 U17755 ( .A1(n15929), .A2(n15931), .ZN(n14586) );
  XNOR2_X1 U17756 ( .A(n14587), .B(n14586), .ZN(n16011) );
  INV_X1 U17757 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n14588) );
  NOR2_X1 U17758 ( .A1(n20135), .A2(n14588), .ZN(n16008) );
  AOI21_X1 U17759 ( .B1(n20120), .B2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n16008), .ZN(n14591) );
  NAND2_X1 U17760 ( .A1(n14589), .A2(n15961), .ZN(n14590) );
  OAI211_X1 U17761 ( .C1(n14592), .C2(n14616), .A(n14591), .B(n14590), .ZN(
        n14593) );
  AOI21_X1 U17762 ( .B1(n16011), .B2(n12697), .A(n14593), .ZN(n14594) );
  INV_X1 U17763 ( .A(n14594), .ZN(P1_U2983) );
  INV_X1 U17764 ( .A(n14595), .ZN(n14596) );
  AND2_X1 U17765 ( .A1(n15956), .A2(n14596), .ZN(n15921) );
  INV_X1 U17766 ( .A(n14597), .ZN(n14599) );
  OAI21_X1 U17767 ( .B1(n15921), .B2(n14599), .A(n14598), .ZN(n14601) );
  AOI22_X1 U17768 ( .A1(n15808), .A2(n16027), .B1(
        P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n15955), .ZN(n14600) );
  XNOR2_X1 U17769 ( .A(n14601), .B(n14600), .ZN(n16024) );
  INV_X1 U17770 ( .A(n16024), .ZN(n14607) );
  AOI22_X1 U17771 ( .A1(n20120), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n20162), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n14602) );
  OAI21_X1 U17772 ( .B1(n20130), .B2(n14603), .A(n14602), .ZN(n14604) );
  AOI21_X1 U17773 ( .B1(n14605), .B2(n20125), .A(n14604), .ZN(n14606) );
  OAI21_X1 U17774 ( .B1(n14607), .B2(n19918), .A(n14606), .ZN(P1_U2985) );
  NOR2_X1 U17775 ( .A1(n15957), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14609) );
  NOR2_X1 U17776 ( .A1(n15956), .A2(n15958), .ZN(n14608) );
  MUX2_X1 U17777 ( .A(n14609), .B(n14608), .S(n15955), .Z(n14610) );
  XOR2_X1 U17778 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n14610), .Z(
        n16064) );
  NAND2_X1 U17779 ( .A1(n16064), .A2(n12697), .ZN(n14614) );
  NOR2_X1 U17780 ( .A1(n20135), .A2(n15889), .ZN(n16062) );
  NOR2_X1 U17781 ( .A1(n20130), .A2(n14611), .ZN(n14612) );
  AOI211_X1 U17782 ( .C1(n20120), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n16062), .B(n14612), .ZN(n14613) );
  OAI211_X1 U17783 ( .C1(n14616), .C2(n14615), .A(n14614), .B(n14613), .ZN(
        P1_U2988) );
  INV_X1 U17784 ( .A(n14617), .ZN(n14618) );
  AOI21_X1 U17785 ( .B1(n14619), .B2(n20157), .A(n14618), .ZN(n14624) );
  INV_X1 U17786 ( .A(n14620), .ZN(n14622) );
  OAI21_X1 U17787 ( .B1(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n14622), .A(
        n14621), .ZN(n14623) );
  OAI211_X1 U17788 ( .C1(n14625), .C2(n16082), .A(n14624), .B(n14623), .ZN(
        P1_U3001) );
  INV_X1 U17789 ( .A(n14626), .ZN(n14629) );
  INV_X1 U17790 ( .A(n14637), .ZN(n14647) );
  NOR3_X1 U17791 ( .A1(n14647), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n14636), .ZN(n14627) );
  AOI211_X1 U17792 ( .C1(n20157), .C2(n14629), .A(n14628), .B(n14627), .ZN(
        n14633) );
  OR2_X1 U17793 ( .A1(n14631), .A2(n14630), .ZN(n14632) );
  OAI211_X1 U17794 ( .C1(n14634), .C2(n16082), .A(n14633), .B(n14632), .ZN(
        P1_U3002) );
  AND3_X1 U17795 ( .A1(n14637), .A2(n14636), .A3(n14635), .ZN(n14638) );
  AOI211_X1 U17796 ( .C1(n20157), .C2(n14640), .A(n14639), .B(n14638), .ZN(
        n14642) );
  NAND2_X1 U17797 ( .A1(n14649), .A2(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14641) );
  OAI211_X1 U17798 ( .C1(n14643), .C2(n16082), .A(n14642), .B(n14641), .ZN(
        P1_U3003) );
  AOI21_X1 U17799 ( .B1(n14645), .B2(n20157), .A(n14644), .ZN(n14646) );
  OAI21_X1 U17800 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14647), .A(
        n14646), .ZN(n14648) );
  AOI21_X1 U17801 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14649), .A(
        n14648), .ZN(n14650) );
  OAI21_X1 U17802 ( .B1(n14651), .B2(n16082), .A(n14650), .ZN(P1_U3004) );
  INV_X1 U17803 ( .A(n14652), .ZN(n14656) );
  NOR3_X1 U17804 ( .A1(n14668), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A3(
        n14653), .ZN(n14654) );
  AOI211_X1 U17805 ( .C1(n20157), .C2(n14656), .A(n14655), .B(n14654), .ZN(
        n14659) );
  NOR3_X1 U17806 ( .A1(n14668), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n14657), .ZN(n14661) );
  OAI21_X1 U17807 ( .B1(n14661), .B2(n14664), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14658) );
  OAI211_X1 U17808 ( .C1(n14660), .C2(n16082), .A(n14659), .B(n14658), .ZN(
        P1_U3005) );
  AOI211_X1 U17809 ( .C1(n20157), .C2(n14663), .A(n14662), .B(n14661), .ZN(
        n14666) );
  NAND2_X1 U17810 ( .A1(n14664), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14665) );
  OAI211_X1 U17811 ( .C1(n14667), .C2(n16082), .A(n14666), .B(n14665), .ZN(
        P1_U3006) );
  NOR3_X1 U17812 ( .A1(n14668), .A2(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        n15990), .ZN(n14678) );
  AND3_X1 U17813 ( .A1(n14693), .A2(n14669), .A3(n15990), .ZN(n15983) );
  NAND2_X1 U17814 ( .A1(n14670), .A2(n15983), .ZN(n14672) );
  AOI21_X1 U17815 ( .B1(n14673), .B2(n14672), .A(n14671), .ZN(n14677) );
  NOR2_X1 U17816 ( .A1(n14674), .A2(n20137), .ZN(n14676) );
  NOR4_X1 U17817 ( .A1(n14678), .A2(n14677), .A3(n14676), .A4(n14675), .ZN(
        n14679) );
  OAI21_X1 U17818 ( .B1(n14680), .B2(n16082), .A(n14679), .ZN(P1_U3007) );
  NOR2_X1 U17819 ( .A1(n14681), .A2(n20137), .ZN(n14682) );
  AOI211_X1 U17820 ( .C1(n15806), .C2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n14683), .B(n14682), .ZN(n14691) );
  INV_X1 U17821 ( .A(n14684), .ZN(n14687) );
  AND2_X1 U17822 ( .A1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n16037), .ZN(
        n16041) );
  AOI22_X1 U17823 ( .A1(n14685), .A2(n16038), .B1(n14716), .B2(n16041), .ZN(
        n16032) );
  NOR2_X1 U17824 ( .A1(n16032), .A2(n14686), .ZN(n14694) );
  AOI21_X1 U17825 ( .B1(n14687), .B2(n16030), .A(n14694), .ZN(n15999) );
  NOR2_X1 U17826 ( .A1(n15999), .A2(n15912), .ZN(n14695) );
  NAND2_X1 U17827 ( .A1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n14695), .ZN(
        n15816) );
  AOI21_X1 U17828 ( .B1(n12690), .B2(n9988), .A(n15816), .ZN(n14689) );
  NAND2_X1 U17829 ( .A1(n14689), .A2(n14688), .ZN(n14690) );
  OAI211_X1 U17830 ( .C1(n14692), .C2(n16082), .A(n14691), .B(n14690), .ZN(
        P1_U3009) );
  INV_X1 U17831 ( .A(n14693), .ZN(n15807) );
  OAI21_X1 U17832 ( .B1(n16030), .B2(n14694), .A(n15807), .ZN(n14697) );
  INV_X1 U17833 ( .A(n14695), .ZN(n14696) );
  AOI22_X1 U17834 ( .A1(n15992), .A2(n14697), .B1(n15810), .B2(n14696), .ZN(
        n14698) );
  INV_X1 U17835 ( .A(n14698), .ZN(n14702) );
  NOR2_X1 U17836 ( .A1(n20135), .A2(n20713), .ZN(n14699) );
  AOI21_X1 U17837 ( .B1(n20160), .B2(n14700), .A(n14699), .ZN(n14701) );
  OAI211_X1 U17838 ( .C1(n15838), .C2(n20137), .A(n14702), .B(n14701), .ZN(
        P1_U3011) );
  NAND2_X1 U17839 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n15984), .ZN(
        n16028) );
  NOR2_X1 U17840 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n16028), .ZN(
        n14708) );
  INV_X1 U17841 ( .A(n15859), .ZN(n14706) );
  NAND2_X1 U17842 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n16037), .ZN(
        n16029) );
  AOI21_X1 U17843 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16038), .A(
        n20154), .ZN(n14703) );
  AOI211_X1 U17844 ( .C1(n20134), .C2(n16029), .A(n20132), .B(n14703), .ZN(
        n16026) );
  OAI21_X1 U17845 ( .B1(n16010), .B2(n14709), .A(n16026), .ZN(n16003) );
  NAND2_X1 U17846 ( .A1(n16003), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14705) );
  OAI211_X1 U17847 ( .C1(n14706), .C2(n20137), .A(n14705), .B(n14704), .ZN(
        n14707) );
  AOI21_X1 U17848 ( .B1(n14709), .B2(n14708), .A(n14707), .ZN(n14710) );
  OAI21_X1 U17849 ( .B1(n14711), .B2(n16082), .A(n14710), .ZN(P1_U3013) );
  NAND3_X1 U17850 ( .A1(n14713), .A2(n14712), .A3(n20160), .ZN(n14722) );
  AOI21_X1 U17851 ( .B1(n20157), .B2(n14715), .A(n14714), .ZN(n14721) );
  INV_X1 U17852 ( .A(n14716), .ZN(n16042) );
  NAND2_X1 U17853 ( .A1(n16042), .A2(n20154), .ZN(n14726) );
  INV_X1 U17854 ( .A(n16040), .ZN(n14717) );
  AOI21_X1 U17855 ( .B1(n14726), .B2(n20153), .A(n14717), .ZN(n14718) );
  OR2_X1 U17856 ( .A1(n14718), .A2(n20165), .ZN(n14720) );
  OR3_X1 U17857 ( .A1(n16010), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(
        n20163), .ZN(n14719) );
  NAND4_X1 U17858 ( .A1(n14722), .A2(n14721), .A3(n14720), .A4(n14719), .ZN(
        P1_U3030) );
  NAND2_X1 U17859 ( .A1(n14723), .A2(n20160), .ZN(n14732) );
  AOI21_X1 U17860 ( .B1(n20157), .B2(n14725), .A(n14724), .ZN(n14731) );
  NAND2_X1 U17861 ( .A1(n14726), .A2(n20153), .ZN(n14730) );
  NAND2_X1 U17862 ( .A1(n14727), .A2(n16040), .ZN(n14728) );
  NAND2_X1 U17863 ( .A1(n14728), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n14729) );
  NAND4_X1 U17864 ( .A1(n14732), .A2(n14731), .A3(n14730), .A4(n14729), .ZN(
        P1_U3031) );
  NAND3_X1 U17865 ( .A1(n14734), .A2(n15786), .A3(n14733), .ZN(n15804) );
  AOI22_X1 U17866 ( .A1(n20172), .A2(n20585), .B1(n11934), .B2(n14735), .ZN(
        n14736) );
  NAND2_X1 U17867 ( .A1(n15804), .A2(n14736), .ZN(n14737) );
  MUX2_X1 U17868 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B(n14737), .S(
        n20170), .Z(P1_U3478) );
  OR2_X1 U17869 ( .A1(n20372), .A2(n14738), .ZN(n14743) );
  NOR2_X1 U17870 ( .A1(n13202), .A2(n14745), .ZN(n14740) );
  AOI22_X1 U17871 ( .A1(n15762), .A2(n14741), .B1(n14740), .B2(n14739), .ZN(
        n14742) );
  NAND2_X1 U17872 ( .A1(n14743), .A2(n14742), .ZN(n15760) );
  INV_X1 U17873 ( .A(n15760), .ZN(n14749) );
  INV_X1 U17874 ( .A(n19909), .ZN(n20746) );
  AOI22_X1 U17875 ( .A1(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n20165), .B1(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n14744), .ZN(n14754) );
  NOR3_X1 U17876 ( .A1(n13202), .A2(n14745), .A3(n20744), .ZN(n14746) );
  AOI21_X1 U17877 ( .B1(n14747), .B2(n14754), .A(n14746), .ZN(n14748) );
  OAI21_X1 U17878 ( .B1(n14749), .B2(n20746), .A(n14748), .ZN(n14750) );
  MUX2_X1 U17879 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n14750), .S(
        n20748), .Z(P1_U3473) );
  INV_X1 U17880 ( .A(n14751), .ZN(n14752) );
  OAI222_X1 U17881 ( .A1(n20744), .A2(n14755), .B1(n14754), .B2(n14753), .C1(
        n20746), .C2(n14752), .ZN(n14756) );
  MUX2_X1 U17882 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(n14756), .S(
        n20748), .Z(P1_U3472) );
  NOR2_X1 U17883 ( .A1(n13666), .A2(n15488), .ZN(n15480) );
  NAND2_X1 U17884 ( .A1(n15480), .A2(n19076), .ZN(n14765) );
  AOI22_X1 U17885 ( .A1(n19099), .A2(n19166), .B1(n19064), .B2(
        P2_EBX_REG_0__SCAN_IN), .ZN(n14758) );
  NOR2_X1 U17886 ( .A1(n19080), .A2(n19116), .ZN(n18896) );
  OAI21_X1 U17887 ( .B1(n19065), .B2(n18896), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n14757) );
  OAI211_X1 U17888 ( .C1(n14759), .C2(n19110), .A(n14758), .B(n14757), .ZN(
        n14762) );
  NOR2_X1 U17889 ( .A1(n14760), .A2(n19091), .ZN(n14761) );
  AOI211_X1 U17890 ( .C1(n19107), .C2(n14763), .A(n14762), .B(n14761), .ZN(
        n14764) );
  OAI211_X1 U17891 ( .C1(n19093), .C2(n19210), .A(n14765), .B(n14764), .ZN(
        P2_U2855) );
  NAND2_X1 U17892 ( .A1(n16127), .A2(n13520), .ZN(n14766) );
  OAI21_X1 U17893 ( .B1(n13520), .B2(n16123), .A(n14766), .ZN(P2_U2856) );
  NAND2_X1 U17894 ( .A1(n14856), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14770) );
  NAND2_X1 U17895 ( .A1(n16145), .A2(n13520), .ZN(n14769) );
  OAI211_X1 U17896 ( .C1(n14872), .C2(n14865), .A(n14770), .B(n14769), .ZN(
        P2_U2858) );
  INV_X1 U17897 ( .A(n14771), .ZN(n14772) );
  NOR2_X1 U17898 ( .A1(n14773), .A2(n14772), .ZN(n14774) );
  XNOR2_X1 U17899 ( .A(n14774), .B(n9735), .ZN(n14882) );
  AOI21_X1 U17900 ( .B1(n14776), .B2(n9684), .A(n14775), .ZN(n14777) );
  NOR2_X1 U17901 ( .A1(n16157), .A2(n14856), .ZN(n14778) );
  AOI21_X1 U17902 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n14856), .A(n14778), .ZN(
        n14779) );
  OAI21_X1 U17903 ( .B1(n14882), .B2(n14865), .A(n14779), .ZN(P2_U2859) );
  AOI21_X1 U17904 ( .B1(n14782), .B2(n14781), .A(n14780), .ZN(n14783) );
  INV_X1 U17905 ( .A(n14783), .ZN(n14889) );
  NAND2_X1 U17906 ( .A1(n14793), .A2(n14784), .ZN(n14785) );
  NOR2_X1 U17907 ( .A1(n15210), .A2(n14856), .ZN(n14786) );
  AOI21_X1 U17908 ( .B1(P2_EBX_REG_27__SCAN_IN), .B2(n14856), .A(n14786), .ZN(
        n14787) );
  OAI21_X1 U17909 ( .B1(n14889), .B2(n14865), .A(n14787), .ZN(P2_U2860) );
  XNOR2_X1 U17910 ( .A(n14789), .B(n14788), .ZN(n14900) );
  OR2_X1 U17911 ( .A1(n14790), .A2(n14791), .ZN(n14792) );
  NAND2_X1 U17912 ( .A1(n14793), .A2(n14792), .ZN(n15222) );
  NOR2_X1 U17913 ( .A1(n15222), .A2(n14856), .ZN(n14794) );
  AOI21_X1 U17914 ( .B1(P2_EBX_REG_26__SCAN_IN), .B2(n14856), .A(n14794), .ZN(
        n14795) );
  OAI21_X1 U17915 ( .B1(n14900), .B2(n14865), .A(n14795), .ZN(P2_U2861) );
  OAI21_X1 U17916 ( .B1(n14798), .B2(n14797), .A(n14796), .ZN(n14909) );
  INV_X1 U17917 ( .A(n14799), .ZN(n14801) );
  INV_X1 U17918 ( .A(n14810), .ZN(n14800) );
  AOI21_X1 U17919 ( .B1(n14801), .B2(n14800), .A(n14790), .ZN(n16189) );
  NOR2_X1 U17920 ( .A1(n13520), .A2(n10683), .ZN(n14802) );
  AOI21_X1 U17921 ( .B1(n16189), .B2(n13520), .A(n14802), .ZN(n14803) );
  OAI21_X1 U17922 ( .B1(n14909), .B2(n14865), .A(n14803), .ZN(P2_U2862) );
  OAI21_X1 U17923 ( .B1(n14806), .B2(n14805), .A(n14804), .ZN(n14808) );
  XOR2_X1 U17924 ( .A(n14808), .B(n14807), .Z(n14910) );
  AND2_X1 U17925 ( .A1(n14817), .A2(n14809), .ZN(n14811) );
  OR2_X1 U17926 ( .A1(n14811), .A2(n14810), .ZN(n16200) );
  NOR2_X1 U17927 ( .A1(n16200), .A2(n14856), .ZN(n14812) );
  AOI21_X1 U17928 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n14856), .A(n14812), .ZN(
        n14813) );
  OAI21_X1 U17929 ( .B1(n14910), .B2(n14865), .A(n14813), .ZN(P2_U2863) );
  NAND2_X1 U17930 ( .A1(n14814), .A2(n14815), .ZN(n14816) );
  AND2_X1 U17931 ( .A1(n14817), .A2(n14816), .ZN(n16215) );
  AOI21_X1 U17932 ( .B1(n14820), .B2(n14819), .A(n14818), .ZN(n14918) );
  NAND2_X1 U17933 ( .A1(n14918), .A2(n14844), .ZN(n14822) );
  NAND2_X1 U17934 ( .A1(n14856), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n14821) );
  OAI211_X1 U17935 ( .C1(n15253), .C2(n14856), .A(n14822), .B(n14821), .ZN(
        P2_U2864) );
  OAI21_X1 U17936 ( .B1(n14833), .B2(n14823), .A(n14814), .ZN(n16222) );
  INV_X1 U17937 ( .A(n14824), .ZN(n14825) );
  AOI21_X1 U17938 ( .B1(n14826), .B2(n14825), .A(n11519), .ZN(n14932) );
  NAND2_X1 U17939 ( .A1(n14932), .A2(n14844), .ZN(n14828) );
  NAND2_X1 U17940 ( .A1(n14856), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n14827) );
  OAI211_X1 U17941 ( .C1(n16222), .C2(n14856), .A(n14828), .B(n14827), .ZN(
        P2_U2865) );
  INV_X1 U17942 ( .A(n14829), .ZN(n14831) );
  OAI21_X1 U17943 ( .B1(n14831), .B2(n14830), .A(n14825), .ZN(n14949) );
  AND2_X1 U17944 ( .A1(n14839), .A2(n14832), .ZN(n14834) );
  OR2_X1 U17945 ( .A1(n14834), .A2(n14833), .ZN(n18880) );
  MUX2_X1 U17946 ( .A(n18880), .B(n10613), .S(n14856), .Z(n14835) );
  OAI21_X1 U17947 ( .B1(n14865), .B2(n14949), .A(n14835), .ZN(P2_U2866) );
  OAI21_X1 U17948 ( .B1(n14836), .B2(n14837), .A(n14829), .ZN(n14959) );
  INV_X1 U17949 ( .A(n14848), .ZN(n14841) );
  INV_X1 U17950 ( .A(n14838), .ZN(n14840) );
  OAI21_X1 U17951 ( .B1(n14841), .B2(n14840), .A(n14839), .ZN(n18903) );
  INV_X1 U17952 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n18893) );
  MUX2_X1 U17953 ( .A(n18903), .B(n18893), .S(n14856), .Z(n14842) );
  OAI21_X1 U17954 ( .B1(n14865), .B2(n14959), .A(n14842), .ZN(P2_U2867) );
  AOI21_X1 U17955 ( .B1(n14843), .B2(n9664), .A(n14836), .ZN(n14968) );
  NAND2_X1 U17956 ( .A1(n14968), .A2(n14844), .ZN(n14850) );
  NAND2_X1 U17957 ( .A1(n14845), .A2(n14846), .ZN(n14847) );
  AND2_X1 U17958 ( .A1(n14848), .A2(n14847), .ZN(n18912) );
  NAND2_X1 U17959 ( .A1(n18912), .A2(n13520), .ZN(n14849) );
  OAI211_X1 U17960 ( .C1(n13520), .C2(n10639), .A(n14850), .B(n14849), .ZN(
        P2_U2868) );
  OAI21_X1 U17961 ( .B1(n10032), .B2(n14853), .A(n9664), .ZN(n14978) );
  OAI21_X1 U17962 ( .B1(n14859), .B2(n14854), .A(n14845), .ZN(n15322) );
  NOR2_X1 U17963 ( .A1(n15322), .A2(n14856), .ZN(n14855) );
  AOI21_X1 U17964 ( .B1(P2_EBX_REG_18__SCAN_IN), .B2(n14856), .A(n14855), .ZN(
        n14857) );
  OAI21_X1 U17965 ( .B1(n14865), .B2(n14978), .A(n14857), .ZN(P2_U2869) );
  OAI21_X1 U17966 ( .B1(n13627), .B2(n14858), .A(n14851), .ZN(n14987) );
  AOI21_X1 U17967 ( .B1(n14861), .B2(n14860), .A(n14859), .ZN(n18937) );
  INV_X1 U17968 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n14862) );
  NOR2_X1 U17969 ( .A1(n13520), .A2(n14862), .ZN(n14863) );
  AOI21_X1 U17970 ( .B1(n18937), .B2(n13520), .A(n14863), .ZN(n14864) );
  OAI21_X1 U17971 ( .B1(n14865), .B2(n14987), .A(n14864), .ZN(P2_U2870) );
  INV_X1 U17972 ( .A(n16144), .ZN(n14867) );
  OAI22_X1 U17973 ( .A1(n14867), .A2(n19153), .B1(n19152), .B2(n14866), .ZN(
        n14868) );
  AOI21_X1 U17974 ( .B1(n15000), .B2(n14869), .A(n14868), .ZN(n14871) );
  AOI22_X1 U17975 ( .A1(n19121), .A2(BUF2_REG_29__SCAN_IN), .B1(n19123), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n14870) );
  OAI211_X1 U17976 ( .C1(n14872), .C2(n15002), .A(n14871), .B(n14870), .ZN(
        P2_U2890) );
  OR2_X1 U17977 ( .A1(n14875), .A2(n14874), .ZN(n14876) );
  NAND2_X1 U17978 ( .A1(n14873), .A2(n14876), .ZN(n16164) );
  OAI22_X1 U17979 ( .A1(n16164), .A2(n19153), .B1(n19152), .B2(n14877), .ZN(
        n14878) );
  AOI21_X1 U17980 ( .B1(n15000), .B2(n14879), .A(n14878), .ZN(n14881) );
  AOI22_X1 U17981 ( .A1(n19121), .A2(BUF2_REG_28__SCAN_IN), .B1(n19123), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n14880) );
  OAI211_X1 U17982 ( .C1(n14882), .C2(n15002), .A(n14881), .B(n14880), .ZN(
        P2_U2891) );
  XNOR2_X1 U17983 ( .A(n14891), .B(n14883), .ZN(n16176) );
  OAI22_X1 U17984 ( .A1(n16176), .A2(n19153), .B1(n19152), .B2(n14884), .ZN(
        n14885) );
  AOI21_X1 U17985 ( .B1(n15000), .B2(n14886), .A(n14885), .ZN(n14888) );
  AOI22_X1 U17986 ( .A1(n19121), .A2(BUF2_REG_27__SCAN_IN), .B1(n19123), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n14887) );
  OAI211_X1 U17987 ( .C1(n14889), .C2(n15002), .A(n14888), .B(n14887), .ZN(
        P2_U2892) );
  INV_X1 U17988 ( .A(n14890), .ZN(n14893) );
  INV_X1 U17989 ( .A(n14903), .ZN(n14892) );
  AOI21_X1 U17990 ( .B1(n14893), .B2(n14892), .A(n14891), .ZN(n16178) );
  INV_X1 U17991 ( .A(n16178), .ZN(n14895) );
  OAI22_X1 U17992 ( .A1(n14895), .A2(n19153), .B1(n19152), .B2(n14894), .ZN(
        n14896) );
  AOI21_X1 U17993 ( .B1(n15000), .B2(n14897), .A(n14896), .ZN(n14899) );
  AOI22_X1 U17994 ( .A1(n19121), .A2(BUF2_REG_26__SCAN_IN), .B1(n19123), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n14898) );
  OAI211_X1 U17995 ( .C1(n14900), .C2(n15002), .A(n14899), .B(n14898), .ZN(
        P2_U2893) );
  INV_X1 U17996 ( .A(n15000), .ZN(n14966) );
  AOI22_X1 U17997 ( .A1(n19121), .A2(BUF2_REG_25__SCAN_IN), .B1(n19123), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n14905) );
  AND2_X1 U17998 ( .A1(n14913), .A2(n14901), .ZN(n14902) );
  NOR2_X1 U17999 ( .A1(n14903), .A2(n14902), .ZN(n16188) );
  AOI22_X1 U18000 ( .A1(n19163), .A2(n16188), .B1(P2_EAX_REG_25__SCAN_IN), 
        .B2(n19162), .ZN(n14904) );
  OAI211_X1 U18001 ( .C1(n14906), .C2(n14966), .A(n14905), .B(n14904), .ZN(
        n14907) );
  INV_X1 U18002 ( .A(n14907), .ZN(n14908) );
  OAI21_X1 U18003 ( .B1(n14909), .B2(n15002), .A(n14908), .ZN(P2_U2894) );
  OR2_X1 U18004 ( .A1(n14910), .A2(n15002), .ZN(n14917) );
  NAND2_X1 U18005 ( .A1(n14923), .A2(n14911), .ZN(n14912) );
  AND2_X1 U18006 ( .A1(n14913), .A2(n14912), .ZN(n16201) );
  AOI22_X1 U18007 ( .A1(n19163), .A2(n16201), .B1(P2_EAX_REG_24__SCAN_IN), 
        .B2(n19162), .ZN(n14916) );
  AOI22_X1 U18008 ( .A1(n19121), .A2(BUF2_REG_24__SCAN_IN), .B1(n19123), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n14915) );
  NAND2_X1 U18009 ( .A1(n15000), .A2(n19130), .ZN(n14914) );
  NAND4_X1 U18010 ( .A1(n14917), .A2(n14916), .A3(n14915), .A4(n14914), .ZN(
        P2_U2895) );
  INV_X1 U18011 ( .A(n14918), .ZN(n14931) );
  INV_X1 U18012 ( .A(n19254), .ZN(n14929) );
  INV_X1 U18013 ( .A(n14919), .ZN(n14921) );
  NAND2_X1 U18014 ( .A1(n14934), .A2(n14933), .ZN(n14920) );
  NAND2_X1 U18015 ( .A1(n14921), .A2(n14920), .ZN(n14922) );
  NAND2_X1 U18016 ( .A1(n14923), .A2(n14922), .ZN(n16221) );
  NAND2_X1 U18017 ( .A1(n19162), .A2(P2_EAX_REG_23__SCAN_IN), .ZN(n14924) );
  OAI21_X1 U18018 ( .B1(n19153), .B2(n16221), .A(n14924), .ZN(n14928) );
  INV_X1 U18019 ( .A(n19121), .ZN(n14996) );
  INV_X1 U18020 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n14926) );
  INV_X1 U18021 ( .A(n19123), .ZN(n14994) );
  INV_X1 U18022 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n14925) );
  OAI22_X1 U18023 ( .A1(n14996), .A2(n14926), .B1(n14994), .B2(n14925), .ZN(
        n14927) );
  AOI211_X1 U18024 ( .C1(n15000), .C2(n14929), .A(n14928), .B(n14927), .ZN(
        n14930) );
  OAI21_X1 U18025 ( .B1(n14931), .B2(n15002), .A(n14930), .ZN(P2_U2896) );
  INV_X1 U18026 ( .A(n14932), .ZN(n14941) );
  INV_X1 U18027 ( .A(n19246), .ZN(n14938) );
  XNOR2_X1 U18028 ( .A(n14934), .B(n14943), .ZN(n15733) );
  INV_X1 U18029 ( .A(n15733), .ZN(n14936) );
  OAI22_X1 U18030 ( .A1(n14936), .A2(n19153), .B1(n19152), .B2(n14935), .ZN(
        n14937) );
  AOI21_X1 U18031 ( .B1(n15000), .B2(n14938), .A(n14937), .ZN(n14940) );
  AOI22_X1 U18032 ( .A1(n19121), .A2(BUF2_REG_22__SCAN_IN), .B1(n19123), .B2(
        BUF1_REG_22__SCAN_IN), .ZN(n14939) );
  OAI211_X1 U18033 ( .C1(n14941), .C2(n15002), .A(n14940), .B(n14939), .ZN(
        P2_U2897) );
  INV_X1 U18034 ( .A(n19239), .ZN(n19133) );
  OR2_X1 U18035 ( .A1(n14951), .A2(n14942), .ZN(n14944) );
  NAND2_X1 U18036 ( .A1(n14944), .A2(n14943), .ZN(n18889) );
  OAI22_X1 U18037 ( .A1(n18889), .A2(n19153), .B1(n19152), .B2(n14945), .ZN(
        n14946) );
  AOI21_X1 U18038 ( .B1(n15000), .B2(n19133), .A(n14946), .ZN(n14948) );
  AOI22_X1 U18039 ( .A1(n19121), .A2(BUF2_REG_21__SCAN_IN), .B1(n19123), .B2(
        BUF1_REG_21__SCAN_IN), .ZN(n14947) );
  OAI211_X1 U18040 ( .C1(n14949), .C2(n15002), .A(n14948), .B(n14947), .ZN(
        P2_U2898) );
  INV_X1 U18041 ( .A(n19234), .ZN(n14956) );
  INV_X1 U18042 ( .A(n14950), .ZN(n14953) );
  INV_X1 U18043 ( .A(n14963), .ZN(n14952) );
  AOI21_X1 U18044 ( .B1(n14953), .B2(n14952), .A(n14951), .ZN(n18900) );
  INV_X1 U18045 ( .A(n18900), .ZN(n14954) );
  OAI22_X1 U18046 ( .A1(n14954), .A2(n19153), .B1(n19152), .B2(n20911), .ZN(
        n14955) );
  AOI21_X1 U18047 ( .B1(n15000), .B2(n14956), .A(n14955), .ZN(n14958) );
  AOI22_X1 U18048 ( .A1(n19121), .A2(BUF2_REG_20__SCAN_IN), .B1(n19123), .B2(
        BUF1_REG_20__SCAN_IN), .ZN(n14957) );
  OAI211_X1 U18049 ( .C1(n14959), .C2(n15002), .A(n14958), .B(n14957), .ZN(
        P2_U2899) );
  AOI22_X1 U18050 ( .A1(n19121), .A2(BUF2_REG_19__SCAN_IN), .B1(n19123), .B2(
        BUF1_REG_19__SCAN_IN), .ZN(n14965) );
  NOR2_X1 U18051 ( .A1(n14961), .A2(n14960), .ZN(n14962) );
  OR2_X1 U18052 ( .A1(n14963), .A2(n14962), .ZN(n18915) );
  INV_X1 U18053 ( .A(n18915), .ZN(n15305) );
  AOI22_X1 U18054 ( .A1(n19163), .A2(n15305), .B1(n19162), .B2(
        P2_EAX_REG_19__SCAN_IN), .ZN(n14964) );
  OAI211_X1 U18055 ( .C1(n19231), .C2(n14966), .A(n14965), .B(n14964), .ZN(
        n14967) );
  AOI21_X1 U18056 ( .B1(n14968), .B2(n19164), .A(n14967), .ZN(n14969) );
  INV_X1 U18057 ( .A(n14969), .ZN(P2_U2900) );
  INV_X1 U18058 ( .A(n14970), .ZN(n14971) );
  XNOR2_X1 U18059 ( .A(n14981), .B(n14971), .ZN(n18922) );
  INV_X1 U18060 ( .A(n18922), .ZN(n15321) );
  OAI22_X1 U18061 ( .A1(n15321), .A2(n19153), .B1(n19152), .B2(n14972), .ZN(
        n14975) );
  INV_X1 U18062 ( .A(BUF2_REG_18__SCAN_IN), .ZN(n14973) );
  OAI22_X1 U18063 ( .A1(n14996), .A2(n14973), .B1(n14994), .B2(n16446), .ZN(
        n14974) );
  AOI211_X1 U18064 ( .C1(n15000), .C2(n14976), .A(n14975), .B(n14974), .ZN(
        n14977) );
  OAI21_X1 U18065 ( .B1(n14978), .B2(n15002), .A(n14977), .ZN(P2_U2901) );
  NAND2_X1 U18066 ( .A1(n14990), .A2(n14979), .ZN(n14980) );
  NAND2_X1 U18067 ( .A1(n14981), .A2(n14980), .ZN(n18935) );
  OAI22_X1 U18068 ( .A1(n18935), .A2(n19153), .B1(n19152), .B2(n14982), .ZN(
        n14983) );
  AOI21_X1 U18069 ( .B1(n15000), .B2(n14984), .A(n14983), .ZN(n14986) );
  AOI22_X1 U18070 ( .A1(n19121), .A2(BUF2_REG_17__SCAN_IN), .B1(n19123), .B2(
        BUF1_REG_17__SCAN_IN), .ZN(n14985) );
  OAI211_X1 U18071 ( .C1(n14987), .C2(n15002), .A(n14986), .B(n14985), .ZN(
        P2_U2902) );
  OR2_X1 U18072 ( .A1(n14989), .A2(n14988), .ZN(n14991) );
  AND2_X1 U18073 ( .A1(n14991), .A2(n14990), .ZN(n18950) );
  INV_X1 U18074 ( .A(n18950), .ZN(n14992) );
  OAI22_X1 U18075 ( .A1(n14992), .A2(n19153), .B1(n19152), .B2(n12757), .ZN(
        n14998) );
  INV_X1 U18076 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n14995) );
  INV_X1 U18077 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n14993) );
  OAI22_X1 U18078 ( .A1(n14996), .A2(n14995), .B1(n14994), .B2(n14993), .ZN(
        n14997) );
  AOI211_X1 U18079 ( .C1(n15000), .C2(n14999), .A(n14998), .B(n14997), .ZN(
        n15001) );
  OAI21_X1 U18080 ( .B1(n15003), .B2(n15002), .A(n15001), .ZN(P2_U2903) );
  XNOR2_X1 U18081 ( .A(n15004), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16138) );
  NOR2_X1 U18082 ( .A1(n16257), .A2(n16138), .ZN(n15005) );
  AOI211_X1 U18083 ( .C1(n16252), .C2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n15006), .B(n15005), .ZN(n15007) );
  OAI21_X1 U18084 ( .B1(n16142), .B2(n15182), .A(n15007), .ZN(n15008) );
  AOI21_X1 U18085 ( .B1(n15009), .B2(n16284), .A(n15008), .ZN(n15010) );
  OAI21_X1 U18086 ( .B1(n15011), .B2(n16259), .A(n15010), .ZN(P2_U2984) );
  NAND2_X1 U18087 ( .A1(n15013), .A2(n15012), .ZN(n15015) );
  INV_X1 U18088 ( .A(n15015), .ZN(n15017) );
  OAI22_X1 U18089 ( .A1(n15030), .A2(n15194), .B1(n15017), .B2(n15016), .ZN(
        n15020) );
  XNOR2_X1 U18090 ( .A(n15018), .B(n15200), .ZN(n15019) );
  XNOR2_X1 U18091 ( .A(n15020), .B(n15019), .ZN(n15206) );
  AOI21_X1 U18092 ( .B1(n15200), .B2(n15021), .A(n15022), .ZN(n15204) );
  INV_X1 U18093 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19828) );
  NOR2_X1 U18094 ( .A1(n19089), .A2(n19828), .ZN(n15197) );
  NAND2_X1 U18095 ( .A1(n15031), .A2(n15023), .ZN(n15024) );
  NAND2_X1 U18096 ( .A1(n15025), .A2(n15024), .ZN(n16161) );
  NOR2_X1 U18097 ( .A1(n16257), .A2(n16161), .ZN(n15026) );
  AOI211_X1 U18098 ( .C1(n16252), .C2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15197), .B(n15026), .ZN(n15027) );
  OAI21_X1 U18099 ( .B1(n16157), .B2(n15182), .A(n15027), .ZN(n15028) );
  AOI21_X1 U18100 ( .B1(n15204), .B2(n16284), .A(n15028), .ZN(n15029) );
  OAI21_X1 U18101 ( .B1(n15206), .B2(n16259), .A(n15029), .ZN(P2_U2986) );
  XNOR2_X1 U18102 ( .A(n15030), .B(n15194), .ZN(n15217) );
  INV_X1 U18103 ( .A(n15031), .ZN(n15032) );
  AOI21_X1 U18104 ( .B1(n16166), .B2(n15044), .A(n15032), .ZN(n16119) );
  NAND2_X1 U18105 ( .A1(n16279), .A2(n16119), .ZN(n15033) );
  NAND2_X1 U18106 ( .A1(n19069), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15209) );
  OAI211_X1 U18107 ( .C1(n16288), .C2(n16166), .A(n15033), .B(n15209), .ZN(
        n15034) );
  AOI21_X1 U18108 ( .B1(n16170), .B2(n16281), .A(n15034), .ZN(n15037) );
  NAND2_X1 U18109 ( .A1(n15038), .A2(n15194), .ZN(n15214) );
  NAND3_X1 U18110 ( .A1(n15021), .A2(n16284), .A3(n15214), .ZN(n15036) );
  OAI211_X1 U18111 ( .C1(n15217), .C2(n16259), .A(n15037), .B(n15036), .ZN(
        P2_U2987) );
  OAI21_X1 U18112 ( .B1(n15057), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15038), .ZN(n15228) );
  NOR2_X1 U18113 ( .A1(n15039), .A2(n15052), .ZN(n15041) );
  XNOR2_X1 U18114 ( .A(n15041), .B(n15040), .ZN(n15218) );
  NAND2_X1 U18115 ( .A1(n15218), .A2(n16282), .ZN(n15048) );
  INV_X1 U18116 ( .A(n15222), .ZN(n16179) );
  OR2_X1 U18117 ( .A1(n15042), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15043) );
  NAND2_X1 U18118 ( .A1(n15044), .A2(n15043), .ZN(n16182) );
  NAND2_X1 U18119 ( .A1(n19069), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15219) );
  NAND2_X1 U18120 ( .A1(n16252), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15045) );
  OAI211_X1 U18121 ( .C1(n16257), .C2(n16182), .A(n15219), .B(n15045), .ZN(
        n15046) );
  AOI21_X1 U18122 ( .B1(n16179), .B2(n16281), .A(n15046), .ZN(n15047) );
  OAI211_X1 U18123 ( .C1(n16260), .C2(n15228), .A(n15048), .B(n15047), .ZN(
        P2_U2988) );
  INV_X1 U18124 ( .A(n15039), .ZN(n15053) );
  OAI21_X1 U18125 ( .B1(n15050), .B2(n15052), .A(n15049), .ZN(n15051) );
  OAI21_X1 U18126 ( .B1(n15053), .B2(n15052), .A(n15051), .ZN(n15239) );
  AOI21_X1 U18127 ( .B1(n15055), .B2(n15068), .A(n15042), .ZN(n16118) );
  NAND2_X1 U18128 ( .A1(n16279), .A2(n16118), .ZN(n15054) );
  NAND2_X1 U18129 ( .A1(n19069), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15229) );
  OAI211_X1 U18130 ( .C1(n16288), .C2(n15055), .A(n15054), .B(n15229), .ZN(
        n15060) );
  INV_X1 U18131 ( .A(n15057), .ZN(n15058) );
  OAI21_X1 U18132 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n15056), .A(
        n15058), .ZN(n15235) );
  NOR2_X1 U18133 ( .A1(n15235), .A2(n16260), .ZN(n15059) );
  AOI211_X1 U18134 ( .C1(n16281), .C2(n16189), .A(n15060), .B(n15059), .ZN(
        n15061) );
  OAI21_X1 U18135 ( .B1(n15239), .B2(n16259), .A(n15061), .ZN(P2_U2989) );
  XOR2_X1 U18136 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B(n15062), .Z(
        n15063) );
  XNOR2_X1 U18137 ( .A(n15064), .B(n15063), .ZN(n15248) );
  INV_X1 U18138 ( .A(n15065), .ZN(n15066) );
  AOI21_X1 U18139 ( .B1(n15067), .B2(n15066), .A(n15056), .ZN(n15246) );
  INV_X1 U18140 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n19820) );
  NOR2_X1 U18141 ( .A1(n19089), .A2(n19820), .ZN(n15240) );
  AOI21_X1 U18142 ( .B1(n16252), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15240), .ZN(n15071) );
  OAI21_X1 U18143 ( .B1(n15076), .B2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A(
        n15068), .ZN(n16205) );
  INV_X1 U18144 ( .A(n16205), .ZN(n15069) );
  NAND2_X1 U18145 ( .A1(n16279), .A2(n15069), .ZN(n15070) );
  OAI211_X1 U18146 ( .C1(n16200), .C2(n15182), .A(n15071), .B(n15070), .ZN(
        n15072) );
  AOI21_X1 U18147 ( .B1(n15246), .B2(n16284), .A(n15072), .ZN(n15073) );
  OAI21_X1 U18148 ( .B1(n15248), .B2(n16259), .A(n15073), .ZN(P2_U2990) );
  XNOR2_X1 U18149 ( .A(n15075), .B(n15074), .ZN(n15259) );
  INV_X1 U18150 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n16211) );
  AOI21_X1 U18151 ( .B1(n16211), .B2(n15734), .A(n15076), .ZN(n16117) );
  INV_X1 U18152 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n19818) );
  OAI22_X1 U18153 ( .A1(n16288), .A2(n16211), .B1(n19818), .B2(n19089), .ZN(
        n15078) );
  NOR2_X1 U18154 ( .A1(n15253), .A2(n15182), .ZN(n15077) );
  AOI211_X1 U18155 ( .C1(n16279), .C2(n16117), .A(n15078), .B(n15077), .ZN(
        n15080) );
  AOI21_X1 U18156 ( .B1(n15249), .B2(n15262), .A(n15065), .ZN(n15256) );
  NAND2_X1 U18157 ( .A1(n15256), .A2(n16284), .ZN(n15079) );
  OAI211_X1 U18158 ( .C1(n15259), .C2(n16259), .A(n15080), .B(n15079), .ZN(
        P2_U2991) );
  INV_X1 U18159 ( .A(n15380), .ZN(n15081) );
  AOI21_X2 U18160 ( .B1(n15381), .B2(n15379), .A(n15081), .ZN(n15164) );
  INV_X1 U18161 ( .A(n15162), .ZN(n15082) );
  INV_X1 U18162 ( .A(n15152), .ZN(n15083) );
  NAND2_X1 U18163 ( .A1(n15141), .A2(n15140), .ZN(n15139) );
  AND2_X2 U18164 ( .A1(n15139), .A2(n15084), .ZN(n15129) );
  NAND2_X1 U18165 ( .A1(n15086), .A2(n15085), .ZN(n15128) );
  NAND2_X1 U18166 ( .A1(n15088), .A2(n15087), .ZN(n15089) );
  XNOR2_X1 U18167 ( .A(n15090), .B(n15089), .ZN(n15288) );
  XNOR2_X1 U18168 ( .A(n15091), .B(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15286) );
  AOI21_X1 U18169 ( .B1(n20917), .B2(n15100), .A(n15735), .ZN(n15755) );
  NAND2_X1 U18170 ( .A1(n19069), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15280) );
  OAI21_X1 U18171 ( .B1(n16288), .B2(n20917), .A(n15280), .ZN(n15092) );
  AOI21_X1 U18172 ( .B1(n16279), .B2(n15755), .A(n15092), .ZN(n15093) );
  OAI21_X1 U18173 ( .B1(n18880), .B2(n15182), .A(n15093), .ZN(n15094) );
  AOI21_X1 U18174 ( .B1(n15286), .B2(n16284), .A(n15094), .ZN(n15095) );
  OAI21_X1 U18175 ( .B1(n15288), .B2(n16259), .A(n15095), .ZN(P2_U2993) );
  OAI21_X1 U18176 ( .B1(n15097), .B2(n15099), .A(n15096), .ZN(n15098) );
  OAI21_X1 U18177 ( .B1(n9691), .B2(n15099), .A(n15098), .ZN(n15304) );
  INV_X1 U18178 ( .A(n18903), .ZN(n15104) );
  OAI21_X1 U18179 ( .B1(n9721), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15100), .ZN(n18897) );
  NAND2_X1 U18180 ( .A1(n19069), .A2(P2_REIP_REG_20__SCAN_IN), .ZN(n15290) );
  NAND2_X1 U18181 ( .A1(n16252), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n15101) );
  OAI211_X1 U18182 ( .C1(n18897), .C2(n16257), .A(n15290), .B(n15101), .ZN(
        n15103) );
  OAI21_X1 U18183 ( .B1(n9694), .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n15091), .ZN(n15289) );
  NOR2_X1 U18184 ( .A1(n15289), .A2(n16260), .ZN(n15102) );
  AOI211_X1 U18185 ( .C1(n16281), .C2(n15104), .A(n15103), .B(n15102), .ZN(
        n15105) );
  OAI21_X1 U18186 ( .B1(n15304), .B2(n16259), .A(n15105), .ZN(P2_U2994) );
  INV_X1 U18187 ( .A(n15120), .ZN(n15106) );
  AOI21_X1 U18188 ( .B1(n15122), .B2(n15119), .A(n15106), .ZN(n15110) );
  NAND2_X1 U18189 ( .A1(n15108), .A2(n15107), .ZN(n15109) );
  XNOR2_X1 U18190 ( .A(n15110), .B(n15109), .ZN(n15315) );
  AOI21_X1 U18191 ( .B1(n18904), .B2(n15123), .A(n9721), .ZN(n18909) );
  NAND2_X1 U18192 ( .A1(n18909), .A2(n16279), .ZN(n15111) );
  NAND2_X1 U18193 ( .A1(n19069), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15309) );
  OAI211_X1 U18194 ( .C1(n16288), .C2(n18904), .A(n15111), .B(n15309), .ZN(
        n15115) );
  INV_X1 U18195 ( .A(n9694), .ZN(n15113) );
  NAND2_X1 U18196 ( .A1(n15435), .A2(n15296), .ZN(n15118) );
  NAND2_X1 U18197 ( .A1(n15118), .A2(n15293), .ZN(n15112) );
  NAND2_X1 U18198 ( .A1(n15113), .A2(n15112), .ZN(n15312) );
  NOR2_X1 U18199 ( .A1(n15312), .A2(n16260), .ZN(n15114) );
  AOI211_X1 U18200 ( .C1(n16281), .C2(n18912), .A(n15115), .B(n15114), .ZN(
        n15116) );
  OAI21_X1 U18201 ( .B1(n15315), .B2(n16259), .A(n15116), .ZN(P2_U2995) );
  INV_X1 U18202 ( .A(n15318), .ZN(n15117) );
  NOR2_X1 U18203 ( .A1(n15404), .A2(n15117), .ZN(n15135) );
  OAI21_X1 U18204 ( .B1(n15135), .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n15118), .ZN(n15328) );
  NAND2_X1 U18205 ( .A1(n15120), .A2(n15119), .ZN(n15121) );
  XNOR2_X1 U18206 ( .A(n15122), .B(n15121), .ZN(n15316) );
  NAND2_X1 U18207 ( .A1(n15316), .A2(n16282), .ZN(n15127) );
  INV_X1 U18208 ( .A(n15322), .ZN(n18923) );
  OAI21_X1 U18209 ( .B1(n15131), .B2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n15123), .ZN(n15736) );
  NAND2_X1 U18210 ( .A1(n19069), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n15320) );
  NAND2_X1 U18211 ( .A1(n16252), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15124) );
  OAI211_X1 U18212 ( .C1(n15736), .C2(n16257), .A(n15320), .B(n15124), .ZN(
        n15125) );
  AOI21_X1 U18213 ( .B1(n18923), .B2(n16281), .A(n15125), .ZN(n15126) );
  OAI211_X1 U18214 ( .C1(n16260), .C2(n15328), .A(n15127), .B(n15126), .ZN(
        P2_U2996) );
  XNOR2_X1 U18215 ( .A(n15129), .B(n15128), .ZN(n15343) );
  AOI21_X1 U18216 ( .B1(n15155), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15130) );
  OR2_X1 U18217 ( .A1(n15131), .A2(n15130), .ZN(n18940) );
  NOR2_X1 U18218 ( .A1(n18940), .A2(n16257), .ZN(n15134) );
  INV_X1 U18219 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15132) );
  NAND2_X1 U18220 ( .A1(n19069), .A2(P2_REIP_REG_17__SCAN_IN), .ZN(n15338) );
  OAI21_X1 U18221 ( .B1(n16288), .B2(n15132), .A(n15338), .ZN(n15133) );
  AOI211_X1 U18222 ( .C1(n18937), .C2(n16281), .A(n15134), .B(n15133), .ZN(
        n15138) );
  INV_X1 U18223 ( .A(n15331), .ZN(n15335) );
  NAND2_X1 U18224 ( .A1(n15336), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15150) );
  INV_X1 U18225 ( .A(n15135), .ZN(n15136) );
  OAI211_X1 U18226 ( .C1(n15332), .C2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n16284), .B(n15136), .ZN(n15137) );
  OAI211_X1 U18227 ( .C1(n15343), .C2(n16259), .A(n15138), .B(n15137), .ZN(
        P2_U2997) );
  OAI21_X1 U18228 ( .B1(n15141), .B2(n15140), .A(n15139), .ZN(n15344) );
  INV_X1 U18229 ( .A(n18953), .ZN(n15145) );
  INV_X1 U18230 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n18941) );
  XNOR2_X1 U18231 ( .A(n15155), .B(n18941), .ZN(n15753) );
  INV_X1 U18232 ( .A(n15753), .ZN(n18948) );
  INV_X1 U18233 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n15142) );
  NOR2_X1 U18234 ( .A1(n19089), .A2(n15142), .ZN(n15346) );
  AOI21_X1 U18235 ( .B1(n16252), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n15346), .ZN(n15143) );
  OAI21_X1 U18236 ( .B1(n18948), .B2(n16257), .A(n15143), .ZN(n15144) );
  AOI21_X1 U18237 ( .B1(n15145), .B2(n16281), .A(n15144), .ZN(n15149) );
  INV_X1 U18238 ( .A(n15150), .ZN(n15147) );
  INV_X1 U18239 ( .A(n15332), .ZN(n15146) );
  OAI211_X1 U18240 ( .C1(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .C2(n15147), .A(
        n15146), .B(n16284), .ZN(n15148) );
  OAI211_X1 U18241 ( .C1(n15344), .C2(n16259), .A(n15149), .B(n15148), .ZN(
        P2_U2998) );
  OAI21_X1 U18242 ( .B1(n15336), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n15150), .ZN(n15364) );
  NAND2_X1 U18243 ( .A1(n15152), .A2(n15151), .ZN(n15154) );
  XOR2_X1 U18244 ( .A(n15154), .B(n15153), .Z(n15362) );
  AOI22_X1 U18245 ( .A1(n16252), .A2(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        P2_REIP_REG_15__SCAN_IN), .B2(n19069), .ZN(n15159) );
  INV_X1 U18246 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15157) );
  INV_X1 U18247 ( .A(n15167), .ZN(n15156) );
  AOI21_X1 U18248 ( .B1(n15157), .B2(n15156), .A(n15155), .ZN(n18959) );
  NAND2_X1 U18249 ( .A1(n18959), .A2(n16279), .ZN(n15158) );
  OAI211_X1 U18250 ( .C1(n18957), .C2(n15182), .A(n15159), .B(n15158), .ZN(
        n15160) );
  AOI21_X1 U18251 ( .B1(n15362), .B2(n16282), .A(n15160), .ZN(n15161) );
  OAI21_X1 U18252 ( .B1(n16260), .B2(n15364), .A(n15161), .ZN(P2_U2999) );
  NAND2_X1 U18253 ( .A1(n15163), .A2(n15162), .ZN(n15165) );
  XOR2_X1 U18254 ( .A(n15165), .B(n15164), .Z(n15377) );
  NOR2_X1 U18255 ( .A1(n15750), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n15166) );
  OR2_X1 U18256 ( .A1(n15167), .A2(n15166), .ZN(n15737) );
  AOI22_X1 U18257 ( .A1(n16252), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19069), .ZN(n15168) );
  OAI21_X1 U18258 ( .B1(n16257), .B2(n15737), .A(n15168), .ZN(n15169) );
  AOI21_X1 U18259 ( .B1(n18971), .B2(n16281), .A(n15169), .ZN(n15171) );
  INV_X1 U18260 ( .A(n15404), .ZN(n15395) );
  NAND2_X1 U18261 ( .A1(n15395), .A2(n15384), .ZN(n15378) );
  AOI21_X1 U18262 ( .B1(n15367), .B2(n15378), .A(n15336), .ZN(n15374) );
  NAND2_X1 U18263 ( .A1(n15374), .A2(n16284), .ZN(n15170) );
  OAI211_X1 U18264 ( .C1(n15377), .C2(n16259), .A(n15171), .B(n15170), .ZN(
        P2_U3000) );
  NOR2_X1 U18265 ( .A1(n9852), .A2(n15174), .ZN(n15175) );
  XNOR2_X1 U18266 ( .A(n15172), .B(n15175), .ZN(n15460) );
  NAND2_X1 U18267 ( .A1(n16267), .A2(n16266), .ZN(n15179) );
  NAND2_X1 U18268 ( .A1(n15176), .A2(n15177), .ZN(n15463) );
  XNOR2_X1 U18269 ( .A(n15178), .B(n10576), .ZN(n15464) );
  AOI22_X1 U18270 ( .A1(n15463), .A2(n15464), .B1(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15178), .ZN(n16269) );
  XOR2_X1 U18271 ( .A(n15179), .B(n16269), .Z(n15458) );
  OAI21_X1 U18272 ( .B1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n15740), .A(
        n15739), .ZN(n19045) );
  OAI22_X1 U18273 ( .A1(n16288), .A2(n9836), .B1(n16257), .B2(n19045), .ZN(
        n15180) );
  AOI21_X1 U18274 ( .B1(n19069), .B2(P2_REIP_REG_7__SCAN_IN), .A(n15180), .ZN(
        n15181) );
  OAI21_X1 U18275 ( .B1(n15183), .B2(n15182), .A(n15181), .ZN(n15184) );
  AOI21_X1 U18276 ( .B1(n15458), .B2(n16282), .A(n15184), .ZN(n15185) );
  OAI21_X1 U18277 ( .B1(n15460), .B2(n16260), .A(n15185), .ZN(P2_U3007) );
  NOR2_X1 U18278 ( .A1(n15186), .A2(n16259), .ZN(n15191) );
  AND2_X1 U18279 ( .A1(n19074), .A2(n16281), .ZN(n15190) );
  OAI21_X1 U18280 ( .B1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n15187), .A(
        n15741), .ZN(n19072) );
  OAI22_X1 U18281 ( .A1(n16288), .A2(n9839), .B1(n16257), .B2(n19072), .ZN(
        n15188) );
  NOR4_X1 U18282 ( .A1(n15191), .A2(n15190), .A3(n15189), .A4(n15188), .ZN(
        n15192) );
  OAI21_X1 U18283 ( .B1(n16260), .B2(n15193), .A(n15192), .ZN(P2_U3009) );
  NOR2_X1 U18284 ( .A1(n16157), .A2(n15445), .ZN(n15203) );
  INV_X1 U18285 ( .A(n16164), .ZN(n15198) );
  NOR3_X1 U18286 ( .A1(n15195), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n15194), .ZN(n15196) );
  AOI211_X1 U18287 ( .C1(n16306), .C2(n15198), .A(n15197), .B(n15196), .ZN(
        n15199) );
  OAI21_X1 U18288 ( .B1(n15201), .B2(n15200), .A(n15199), .ZN(n15202) );
  AOI211_X1 U18289 ( .C1(n15204), .C2(n16294), .A(n15203), .B(n15202), .ZN(
        n15205) );
  OAI21_X1 U18290 ( .B1(n15206), .B2(n16310), .A(n15205), .ZN(P2_U3018) );
  INV_X1 U18291 ( .A(n15207), .ZN(n15208) );
  OAI211_X1 U18292 ( .C1(n15476), .C2(n16176), .A(n15209), .B(n15208), .ZN(
        n15212) );
  NOR2_X1 U18293 ( .A1(n15210), .A2(n15445), .ZN(n15211) );
  AOI211_X1 U18294 ( .C1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .C2(n15213), .A(
        n15212), .B(n15211), .ZN(n15216) );
  NAND3_X1 U18295 ( .A1(n15021), .A2(n16294), .A3(n15214), .ZN(n15215) );
  OAI211_X1 U18296 ( .C1(n15217), .C2(n16310), .A(n15216), .B(n15215), .ZN(
        P2_U3019) );
  NAND2_X1 U18297 ( .A1(n15218), .A2(n16296), .ZN(n15227) );
  INV_X1 U18298 ( .A(n15234), .ZN(n15225) );
  XNOR2_X1 U18299 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15221) );
  NAND2_X1 U18300 ( .A1(n16306), .A2(n16178), .ZN(n15220) );
  OAI211_X1 U18301 ( .C1(n15230), .C2(n15221), .A(n15220), .B(n15219), .ZN(
        n15224) );
  NOR2_X1 U18302 ( .A1(n15222), .A2(n15445), .ZN(n15223) );
  AOI211_X1 U18303 ( .C1(n15225), .C2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n15224), .B(n15223), .ZN(n15226) );
  OAI211_X1 U18304 ( .C1(n15228), .C2(n16312), .A(n15227), .B(n15226), .ZN(
        P2_U3020) );
  OAI21_X1 U18305 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n15230), .A(
        n15229), .ZN(n15231) );
  AOI21_X1 U18306 ( .B1(n16306), .B2(n16188), .A(n15231), .ZN(n15232) );
  OAI21_X1 U18307 ( .B1(n15234), .B2(n15233), .A(n15232), .ZN(n15237) );
  NOR2_X1 U18308 ( .A1(n15235), .A2(n16312), .ZN(n15236) );
  AOI211_X1 U18309 ( .C1(n16189), .C2(n16316), .A(n15237), .B(n15236), .ZN(
        n15238) );
  OAI21_X1 U18310 ( .B1(n15239), .B2(n16310), .A(n15238), .ZN(P2_U3021) );
  AOI21_X1 U18311 ( .B1(n16306), .B2(n16201), .A(n15240), .ZN(n15244) );
  OAI21_X1 U18312 ( .B1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n15242), .A(
        n15241), .ZN(n15243) );
  OAI211_X1 U18313 ( .C1(n16200), .C2(n15445), .A(n15244), .B(n15243), .ZN(
        n15245) );
  AOI21_X1 U18314 ( .B1(n15246), .B2(n16294), .A(n15245), .ZN(n15247) );
  OAI21_X1 U18315 ( .B1(n15248), .B2(n16310), .A(n15247), .ZN(P2_U3022) );
  NAND2_X1 U18316 ( .A1(n19069), .A2(P2_REIP_REG_23__SCAN_IN), .ZN(n15252) );
  XNOR2_X1 U18317 ( .A(n15249), .B(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15250) );
  NAND2_X1 U18318 ( .A1(n15250), .A2(n15267), .ZN(n15251) );
  OAI211_X1 U18319 ( .C1(n15476), .C2(n16221), .A(n15252), .B(n15251), .ZN(
        n15255) );
  NOR2_X1 U18320 ( .A1(n15253), .A2(n15445), .ZN(n15254) );
  AOI211_X1 U18321 ( .C1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n15283), .A(
        n15255), .B(n15254), .ZN(n15258) );
  NAND2_X1 U18322 ( .A1(n15256), .A2(n16294), .ZN(n15257) );
  OAI211_X1 U18323 ( .C1(n15259), .C2(n16310), .A(n15258), .B(n15257), .ZN(
        P2_U3023) );
  OAI21_X1 U18324 ( .B1(n15091), .B2(n15260), .A(n15270), .ZN(n15261) );
  AND2_X1 U18325 ( .A1(n15262), .A2(n15261), .ZN(n16223) );
  INV_X1 U18326 ( .A(n16223), .ZN(n15275) );
  NAND2_X1 U18327 ( .A1(n9707), .A2(n15264), .ZN(n15265) );
  XNOR2_X1 U18328 ( .A(n15263), .B(n15265), .ZN(n16225) );
  NOR2_X1 U18329 ( .A1(n16222), .A2(n15445), .ZN(n15273) );
  INV_X1 U18330 ( .A(n15283), .ZN(n15271) );
  INV_X1 U18331 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n19816) );
  NOR2_X1 U18332 ( .A1(n19816), .A2(n19089), .ZN(n15266) );
  AOI21_X1 U18333 ( .B1(n15267), .B2(n15270), .A(n15266), .ZN(n15269) );
  NAND2_X1 U18334 ( .A1(n16306), .A2(n15733), .ZN(n15268) );
  OAI211_X1 U18335 ( .C1(n15271), .C2(n15270), .A(n15269), .B(n15268), .ZN(
        n15272) );
  AOI211_X1 U18336 ( .C1(n16225), .C2(n16296), .A(n15273), .B(n15272), .ZN(
        n15274) );
  OAI21_X1 U18337 ( .B1(n16312), .B2(n15275), .A(n15274), .ZN(P2_U3024) );
  INV_X1 U18338 ( .A(n18889), .ZN(n15276) );
  NAND2_X1 U18339 ( .A1(n16306), .A2(n15276), .ZN(n15281) );
  INV_X1 U18340 ( .A(n15277), .ZN(n15278) );
  INV_X1 U18341 ( .A(n15291), .ZN(n15443) );
  NAND4_X1 U18342 ( .A1(n15296), .A2(n15260), .A3(n15278), .A4(n15443), .ZN(
        n15279) );
  NAND3_X1 U18343 ( .A1(n15281), .A2(n15280), .A3(n15279), .ZN(n15282) );
  AOI21_X1 U18344 ( .B1(n15283), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15282), .ZN(n15284) );
  OAI21_X1 U18345 ( .B1(n18880), .B2(n15445), .A(n15284), .ZN(n15285) );
  AOI21_X1 U18346 ( .B1(n15286), .B2(n16294), .A(n15285), .ZN(n15287) );
  OAI21_X1 U18347 ( .B1(n15288), .B2(n16310), .A(n15287), .ZN(P2_U3025) );
  INV_X1 U18348 ( .A(n15289), .ZN(n15302) );
  INV_X1 U18349 ( .A(n15290), .ZN(n15295) );
  NOR2_X1 U18350 ( .A1(n15330), .A2(n15291), .ZN(n15368) );
  AND2_X1 U18351 ( .A1(n15368), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15292) );
  NAND2_X1 U18352 ( .A1(n15292), .A2(n15318), .ZN(n15298) );
  NOR3_X1 U18353 ( .A1(n15298), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        n15293), .ZN(n15294) );
  AOI211_X1 U18354 ( .C1(n16306), .C2(n18900), .A(n15295), .B(n15294), .ZN(
        n15300) );
  OR2_X1 U18355 ( .A1(n16319), .A2(n15296), .ZN(n15297) );
  NAND2_X1 U18356 ( .A1(n15408), .A2(n15297), .ZN(n15325) );
  NOR2_X1 U18357 ( .A1(n15298), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15306) );
  OAI21_X1 U18358 ( .B1(n15325), .B2(n15306), .A(
        P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15299) );
  OAI211_X1 U18359 ( .C1(n18903), .C2(n15445), .A(n15300), .B(n15299), .ZN(
        n15301) );
  AOI21_X1 U18360 ( .B1(n15302), .B2(n16294), .A(n15301), .ZN(n15303) );
  OAI21_X1 U18361 ( .B1(n15304), .B2(n16310), .A(n15303), .ZN(P2_U3026) );
  NAND2_X1 U18362 ( .A1(n15325), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15310) );
  NAND2_X1 U18363 ( .A1(n16306), .A2(n15305), .ZN(n15308) );
  INV_X1 U18364 ( .A(n15306), .ZN(n15307) );
  NAND4_X1 U18365 ( .A1(n15310), .A2(n15309), .A3(n15308), .A4(n15307), .ZN(
        n15311) );
  AOI21_X1 U18366 ( .B1(n18912), .B2(n16316), .A(n15311), .ZN(n15314) );
  OR2_X1 U18367 ( .A1(n15312), .A2(n16312), .ZN(n15313) );
  OAI211_X1 U18368 ( .C1(n15315), .C2(n16310), .A(n15314), .B(n15313), .ZN(
        P2_U3027) );
  NAND2_X1 U18369 ( .A1(n15316), .A2(n16296), .ZN(n15327) );
  NAND3_X1 U18370 ( .A1(n15318), .A2(n15368), .A3(n15317), .ZN(n15319) );
  OAI211_X1 U18371 ( .C1(n15476), .C2(n15321), .A(n15320), .B(n15319), .ZN(
        n15324) );
  NOR2_X1 U18372 ( .A1(n15322), .A2(n15445), .ZN(n15323) );
  AOI211_X1 U18373 ( .C1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .C2(n15325), .A(
        n15324), .B(n15323), .ZN(n15326) );
  OAI211_X1 U18374 ( .C1(n15328), .C2(n16312), .A(n15327), .B(n15326), .ZN(
        P2_U3028) );
  INV_X1 U18375 ( .A(n15329), .ZN(n15334) );
  INV_X1 U18376 ( .A(n16319), .ZN(n15451) );
  INV_X1 U18377 ( .A(n15408), .ZN(n15441) );
  AOI21_X1 U18378 ( .B1(n15330), .B2(n15451), .A(n15441), .ZN(n15399) );
  OAI21_X1 U18379 ( .B1(n15331), .B2(n16319), .A(n15399), .ZN(n15354) );
  INV_X1 U18380 ( .A(n15368), .ZN(n15398) );
  NOR2_X1 U18381 ( .A1(n15398), .A2(n15335), .ZN(n15358) );
  AOI21_X1 U18382 ( .B1(n15336), .B2(n16294), .A(n15358), .ZN(n15345) );
  NOR3_X1 U18383 ( .A1(n15345), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15337), .ZN(n15341) );
  NAND2_X1 U18384 ( .A1(n18937), .A2(n16316), .ZN(n15339) );
  OAI211_X1 U18385 ( .C1(n15476), .C2(n18935), .A(n15339), .B(n15338), .ZN(
        n15340) );
  OAI21_X1 U18386 ( .B1(n15343), .B2(n16310), .A(n15342), .ZN(P2_U3029) );
  INV_X1 U18387 ( .A(n15344), .ZN(n15350) );
  NOR3_X1 U18388 ( .A1(n15345), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A3(
        n15357), .ZN(n15349) );
  AOI21_X1 U18389 ( .B1(n16306), .B2(n18950), .A(n15346), .ZN(n15347) );
  OAI21_X1 U18390 ( .B1(n18953), .B2(n15445), .A(n15347), .ZN(n15348) );
  AOI211_X1 U18391 ( .C1(n15350), .C2(n16296), .A(n15349), .B(n15348), .ZN(
        n15351) );
  OAI21_X1 U18392 ( .B1(n15353), .B2(n15352), .A(n15351), .ZN(P2_U3030) );
  NAND2_X1 U18393 ( .A1(n15354), .A2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15360) );
  INV_X1 U18394 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19803) );
  NOR2_X1 U18395 ( .A1(n19803), .A2(n19089), .ZN(n15356) );
  NOR2_X1 U18396 ( .A1(n15476), .A2(n18965), .ZN(n15355) );
  AOI211_X1 U18397 ( .C1(n15358), .C2(n15357), .A(n15356), .B(n15355), .ZN(
        n15359) );
  OAI211_X1 U18398 ( .C1(n18957), .C2(n15445), .A(n15360), .B(n15359), .ZN(
        n15361) );
  AOI21_X1 U18399 ( .B1(n15362), .B2(n16296), .A(n15361), .ZN(n15363) );
  OAI21_X1 U18400 ( .B1(n16312), .B2(n15364), .A(n15363), .ZN(P2_U3031) );
  OAI21_X1 U18401 ( .B1(n15384), .B2(n15398), .A(n15399), .ZN(n15383) );
  AOI21_X1 U18402 ( .B1(n15366), .B2(n15365), .A(n9659), .ZN(n19126) );
  INV_X1 U18403 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n19801) );
  NAND3_X1 U18404 ( .A1(n15368), .A2(n15384), .A3(n15367), .ZN(n15369) );
  OAI21_X1 U18405 ( .B1(n19801), .B2(n19089), .A(n15369), .ZN(n15370) );
  AOI21_X1 U18406 ( .B1(n16306), .B2(n19126), .A(n15370), .ZN(n15371) );
  OAI21_X1 U18407 ( .B1(n15372), .B2(n15445), .A(n15371), .ZN(n15373) );
  AOI21_X1 U18408 ( .B1(n15383), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n15373), .ZN(n15376) );
  NAND2_X1 U18409 ( .A1(n15374), .A2(n16294), .ZN(n15375) );
  OAI211_X1 U18410 ( .C1(n15377), .C2(n16310), .A(n15376), .B(n15375), .ZN(
        P2_U3032) );
  NOR2_X1 U18411 ( .A1(n15404), .A2(n20933), .ZN(n16238) );
  OAI21_X1 U18412 ( .B1(n16238), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15378), .ZN(n16231) );
  NAND2_X1 U18413 ( .A1(n15380), .A2(n15379), .ZN(n15382) );
  XOR2_X1 U18414 ( .A(n15382), .B(n15381), .Z(n16233) );
  NAND2_X1 U18415 ( .A1(n15383), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15388) );
  NOR3_X1 U18416 ( .A1(n15398), .A2(n15384), .A3(n20933), .ZN(n15386) );
  NOR2_X1 U18417 ( .A1(n16230), .A2(n15445), .ZN(n15385) );
  AOI211_X1 U18418 ( .C1(n19069), .C2(P2_REIP_REG_13__SCAN_IN), .A(n15386), 
        .B(n15385), .ZN(n15387) );
  OAI211_X1 U18419 ( .C1(n15476), .C2(n18986), .A(n15388), .B(n15387), .ZN(
        n15389) );
  AOI21_X1 U18420 ( .B1(n16233), .B2(n16296), .A(n15389), .ZN(n15390) );
  OAI21_X1 U18421 ( .B1(n16312), .B2(n16231), .A(n15390), .ZN(P2_U3033) );
  NOR2_X1 U18422 ( .A1(n15392), .A2(n9826), .ZN(n15393) );
  XNOR2_X1 U18423 ( .A(n15394), .B(n15393), .ZN(n16237) );
  NOR2_X1 U18424 ( .A1(n15395), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16239) );
  OR3_X1 U18425 ( .A1(n16239), .A2(n16238), .A3(n16312), .ZN(n15403) );
  NAND2_X1 U18426 ( .A1(n18993), .A2(n16316), .ZN(n15397) );
  NAND2_X1 U18427 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n19069), .ZN(n15396) );
  OAI211_X1 U18428 ( .C1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .C2(n15398), .A(
        n15397), .B(n15396), .ZN(n15401) );
  NOR2_X1 U18429 ( .A1(n15399), .A2(n20933), .ZN(n15400) );
  AOI211_X1 U18430 ( .C1(n16306), .C2(n18992), .A(n15401), .B(n15400), .ZN(
        n15402) );
  OAI211_X1 U18431 ( .C1(n16237), .C2(n16310), .A(n15403), .B(n15402), .ZN(
        P2_U3034) );
  OAI21_X1 U18432 ( .B1(n15418), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n15404), .ZN(n16247) );
  XNOR2_X1 U18433 ( .A(n15406), .B(n15409), .ZN(n15407) );
  XNOR2_X1 U18434 ( .A(n15405), .B(n15407), .ZN(n16246) );
  OAI21_X1 U18435 ( .B1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16319), .A(
        n15408), .ZN(n15427) );
  NAND2_X1 U18436 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n15443), .ZN(
        n15429) );
  AOI221_X1 U18437 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C1(n15419), .C2(n15409), .A(
        n15429), .ZN(n15411) );
  INV_X1 U18438 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n19795) );
  NOR2_X1 U18439 ( .A1(n19795), .A2(n19089), .ZN(n15410) );
  AOI211_X1 U18440 ( .C1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15427), .A(
        n15411), .B(n15410), .ZN(n15415) );
  OAI22_X1 U18441 ( .A1(n18999), .A2(n15476), .B1(n15445), .B2(n15412), .ZN(
        n15413) );
  INV_X1 U18442 ( .A(n15413), .ZN(n15414) );
  OAI211_X1 U18443 ( .C1(n16246), .C2(n16310), .A(n15415), .B(n15414), .ZN(
        n15416) );
  INV_X1 U18444 ( .A(n15416), .ZN(n15417) );
  OAI21_X1 U18445 ( .B1(n16247), .B2(n16312), .A(n15417), .ZN(P2_U3035) );
  AOI21_X1 U18446 ( .B1(n15419), .B2(n15434), .A(n15418), .ZN(n16253) );
  INV_X1 U18447 ( .A(n16253), .ZN(n15433) );
  NAND2_X1 U18448 ( .A1(n15420), .A2(n15437), .ZN(n15423) );
  OR2_X1 U18449 ( .A1(n9727), .A2(n15421), .ZN(n15422) );
  XNOR2_X1 U18450 ( .A(n15423), .B(n15422), .ZN(n16254) );
  NOR2_X1 U18451 ( .A1(n19019), .A2(n15476), .ZN(n15431) );
  INV_X1 U18452 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n19793) );
  NOR2_X1 U18453 ( .A1(n19793), .A2(n19089), .ZN(n15426) );
  NOR2_X1 U18454 ( .A1(n15424), .A2(n15445), .ZN(n15425) );
  AOI211_X1 U18455 ( .C1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n15427), .A(
        n15426), .B(n15425), .ZN(n15428) );
  OAI21_X1 U18456 ( .B1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n15429), .A(
        n15428), .ZN(n15430) );
  AOI211_X1 U18457 ( .C1(n16254), .C2(n16296), .A(n15431), .B(n15430), .ZN(
        n15432) );
  OAI21_X1 U18458 ( .B1(n15433), .B2(n16312), .A(n15432), .ZN(P2_U3036) );
  OAI21_X1 U18459 ( .B1(n15435), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n15434), .ZN(n16261) );
  OR2_X1 U18460 ( .A1(n10595), .A2(n15438), .ZN(n15439) );
  XNOR2_X1 U18461 ( .A(n15436), .B(n15439), .ZN(n16258) );
  INV_X1 U18462 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n19791) );
  NOR2_X1 U18463 ( .A1(n19791), .A2(n19089), .ZN(n15440) );
  AOI221_X1 U18464 ( .B1(n15443), .B2(n15442), .C1(n15441), .C2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(n15440), .ZN(n15448) );
  INV_X1 U18465 ( .A(n19027), .ZN(n15444) );
  OAI22_X1 U18466 ( .A1(n19030), .A2(n15476), .B1(n15445), .B2(n15444), .ZN(
        n15446) );
  INV_X1 U18467 ( .A(n15446), .ZN(n15447) );
  OAI211_X1 U18468 ( .C1(n16258), .C2(n16310), .A(n15448), .B(n15447), .ZN(
        n15449) );
  INV_X1 U18469 ( .A(n15449), .ZN(n15450) );
  OAI21_X1 U18470 ( .B1(n16261), .B2(n16312), .A(n15450), .ZN(P2_U3037) );
  AOI21_X1 U18471 ( .B1(n15452), .B2(n15451), .A(n15465), .ZN(n16289) );
  AOI22_X1 U18472 ( .A1(n19069), .A2(P2_REIP_REG_7__SCAN_IN), .B1(n16299), 
        .B2(n15454), .ZN(n15453) );
  OAI21_X1 U18473 ( .B1(n16289), .B2(n15454), .A(n15453), .ZN(n15455) );
  AOI21_X1 U18474 ( .B1(n19047), .B2(n16316), .A(n15455), .ZN(n15456) );
  OAI21_X1 U18475 ( .B1(n19051), .B2(n15476), .A(n15456), .ZN(n15457) );
  AOI21_X1 U18476 ( .B1(n15458), .B2(n16296), .A(n15457), .ZN(n15459) );
  OAI21_X1 U18477 ( .B1(n15460), .B2(n16312), .A(n15459), .ZN(P2_U3039) );
  OAI21_X1 U18478 ( .B1(n15462), .B2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A(
        n15461), .ZN(n16280) );
  XOR2_X1 U18479 ( .A(n15464), .B(n15463), .Z(n16283) );
  INV_X1 U18480 ( .A(n15465), .ZN(n15466) );
  OAI21_X1 U18481 ( .B1(n16319), .B2(n15469), .A(n15466), .ZN(n15467) );
  NAND2_X1 U18482 ( .A1(n15467), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15475) );
  INV_X1 U18483 ( .A(n15468), .ZN(n19059) );
  INV_X1 U18484 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n19786) );
  NOR2_X1 U18485 ( .A1(n19786), .A2(n19089), .ZN(n15473) );
  NAND2_X1 U18486 ( .A1(n15469), .A2(n10576), .ZN(n15470) );
  NOR2_X1 U18487 ( .A1(n15471), .A2(n15470), .ZN(n15472) );
  AOI211_X1 U18488 ( .C1(n19059), .C2(n16316), .A(n15473), .B(n15472), .ZN(
        n15474) );
  OAI211_X1 U18489 ( .C1(n15476), .C2(n19063), .A(n15475), .B(n15474), .ZN(
        n15477) );
  AOI21_X1 U18490 ( .B1(n16283), .B2(n16296), .A(n15477), .ZN(n15478) );
  OAI21_X1 U18491 ( .B1(n16280), .B2(n16312), .A(n15478), .ZN(P2_U3040) );
  AOI21_X1 U18492 ( .B1(n13666), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n15480), .ZN(n15485) );
  INV_X1 U18493 ( .A(n15485), .ZN(n15481) );
  OAI222_X1 U18494 ( .A1(n16326), .A2(n15483), .B1(n19848), .B2(n15482), .C1(
        n15828), .C2(n15481), .ZN(n15484) );
  MUX2_X1 U18495 ( .A(n15484), .B(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .S(
        n15498), .Z(P2_U3601) );
  OR2_X1 U18496 ( .A1(n15485), .A2(n15828), .ZN(n15494) );
  OAI211_X1 U18497 ( .C1(n15488), .C2(n15487), .A(n19080), .B(n15486), .ZN(
        n19117) );
  OAI21_X1 U18498 ( .B1(n19080), .B2(n15489), .A(n19117), .ZN(n15492) );
  OAI222_X1 U18499 ( .A1(n16326), .A2(n19209), .B1(n15494), .B2(n15492), .C1(
        n19848), .C2(n15490), .ZN(n15491) );
  MUX2_X1 U18500 ( .A(n15491), .B(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .S(
        n15498), .Z(P2_U3600) );
  INV_X1 U18501 ( .A(n15492), .ZN(n15495) );
  OAI222_X1 U18502 ( .A1(n15495), .A2(n15494), .B1(n19848), .B2(n15493), .C1(
        n16326), .C2(n19859), .ZN(n15496) );
  MUX2_X1 U18503 ( .A(n15496), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15498), .Z(P2_U3599) );
  OAI22_X1 U18504 ( .A1(n19484), .A2(n16326), .B1(n15497), .B2(n19848), .ZN(
        n15499) );
  MUX2_X1 U18505 ( .A(n15499), .B(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(
        n15498), .Z(P2_U3596) );
  NOR3_X2 U18506 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n19690), .ZN(n19419) );
  AOI211_X1 U18507 ( .C1(n10332), .C2(n19697), .A(n19419), .B(n19844), .ZN(
        n15504) );
  OAI21_X1 U18508 ( .B1(P2_STATE2_REG_1__SCAN_IN), .B2(
        P2_STATE2_REG_2__SCAN_IN), .A(n18853), .ZN(n19902) );
  NOR2_X1 U18509 ( .A1(n19902), .A2(n16320), .ZN(n15500) );
  NAND2_X1 U18510 ( .A1(n19856), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19426) );
  INV_X1 U18511 ( .A(n19426), .ZN(n19376) );
  AOI21_X1 U18512 ( .B1(n19424), .B2(n19453), .A(n19896), .ZN(n15502) );
  AOI21_X1 U18513 ( .B1(n19348), .B2(n19376), .A(n15502), .ZN(n15503) );
  INV_X1 U18514 ( .A(n19421), .ZN(n15517) );
  OAI21_X1 U18515 ( .B1(n10332), .B2(n19419), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n15505) );
  OAI21_X1 U18516 ( .B1(n19426), .B2(n19516), .A(n15505), .ZN(n19420) );
  NOR2_X2 U18517 ( .A1(n15507), .A2(n19251), .ZN(n19694) );
  INV_X1 U18518 ( .A(n19694), .ZN(n15513) );
  INV_X1 U18519 ( .A(n19419), .ZN(n15512) );
  NOR2_X1 U18520 ( .A1(n19650), .A2(n19896), .ZN(n19846) );
  AOI22_X1 U18521 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19250), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19249), .ZN(n19706) );
  INV_X1 U18522 ( .A(n19706), .ZN(n19647) );
  AOI22_X1 U18523 ( .A1(n19414), .A2(n19647), .B1(n19446), .B2(n19703), .ZN(
        n15511) );
  OAI21_X1 U18524 ( .B1(n15513), .B2(n15512), .A(n15511), .ZN(n15514) );
  AOI21_X1 U18525 ( .B1(n19420), .B2(n15506), .A(n15514), .ZN(n15515) );
  OAI21_X1 U18526 ( .B1(n15517), .B2(n15516), .A(n15515), .ZN(P2_U3096) );
  AOI21_X1 U18527 ( .B1(n16763), .B2(n17124), .A(n17226), .ZN(n15518) );
  INV_X1 U18528 ( .A(n15518), .ZN(n15530) );
  AOI22_X1 U18529 ( .A1(n17180), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n15519), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15523) );
  AOI22_X1 U18530 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n9637), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15522) );
  AOI22_X1 U18531 ( .A1(n9634), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n13971), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15521) );
  AOI22_X1 U18532 ( .A1(n15584), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15520) );
  NAND4_X1 U18533 ( .A1(n15523), .A2(n15522), .A3(n15521), .A4(n15520), .ZN(
        n15529) );
  AOI22_X1 U18534 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15527) );
  AOI22_X1 U18535 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15526) );
  AOI22_X1 U18536 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9639), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15525) );
  AOI22_X1 U18537 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17128), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15524) );
  NAND4_X1 U18538 ( .A1(n15527), .A2(n15526), .A3(n15525), .A4(n15524), .ZN(
        n15528) );
  NOR2_X1 U18539 ( .A1(n15529), .A2(n15528), .ZN(n17322) );
  OAI22_X1 U18540 ( .A1(n17111), .A2(n15530), .B1(n17322), .B2(n17220), .ZN(
        P3_U2690) );
  NAND2_X1 U18541 ( .A1(n18638), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18470) );
  NOR2_X1 U18542 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18837) );
  AOI21_X1 U18543 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(
        P3_STATE2_REG_1__SCAN_IN), .A(n18837), .ZN(n18693) );
  NOR2_X1 U18544 ( .A1(n17075), .A2(n15531), .ZN(n18184) );
  AOI21_X1 U18545 ( .B1(n18184), .B2(n16517), .A(n18781), .ZN(n15532) );
  NOR2_X1 U18546 ( .A1(n18495), .A2(n15532), .ZN(n18187) );
  INV_X1 U18547 ( .A(n18187), .ZN(n18191) );
  NAND2_X1 U18548 ( .A1(n18470), .A2(n18191), .ZN(n15535) );
  INV_X1 U18549 ( .A(n15535), .ZN(n15534) );
  INV_X1 U18550 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18678) );
  NAND3_X1 U18551 ( .A1(n18678), .A2(n18782), .A3(P3_STATEBS16_REG_SCAN_IN), 
        .ZN(n18446) );
  NAND2_X1 U18552 ( .A1(n18678), .A2(n18782), .ZN(n16512) );
  NAND2_X1 U18553 ( .A1(n18844), .A2(n16512), .ZN(n18185) );
  INV_X1 U18554 ( .A(n18185), .ZN(n18826) );
  INV_X1 U18555 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18833) );
  NOR2_X1 U18556 ( .A1(n18792), .A2(n18833), .ZN(n17819) );
  OAI22_X1 U18557 ( .A1(n18826), .A2(n17819), .B1(n18638), .B2(n18782), .ZN(
        n15537) );
  NAND3_X1 U18558 ( .A1(n18639), .A2(n18191), .A3(n15537), .ZN(n15533) );
  OAI221_X1 U18559 ( .B1(n18639), .B2(n15534), .C1(n18639), .C2(n18446), .A(
        n15533), .ZN(P3_U2864) );
  NAND2_X1 U18560 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18373) );
  NOR2_X1 U18561 ( .A1(n18826), .A2(n17819), .ZN(n15536) );
  AOI221_X1 U18562 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18373), .C1(n15536), 
        .C2(n18373), .A(n15535), .ZN(n18190) );
  INV_X1 U18563 ( .A(n18446), .ZN(n18544) );
  OAI221_X1 U18564 ( .B1(n18544), .B2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .C1(n18544), .C2(n15537), .A(n18191), .ZN(n18188) );
  AOI22_X1 U18565 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18190), .B1(
        n18188), .B2(n18193), .ZN(P3_U2865) );
  NAND2_X1 U18566 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16377) );
  INV_X1 U18567 ( .A(n16377), .ZN(n15709) );
  NAND2_X1 U18568 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17977) );
  INV_X1 U18569 ( .A(n17977), .ZN(n17626) );
  INV_X1 U18570 ( .A(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n17935) );
  NAND2_X1 U18571 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17591) );
  INV_X1 U18572 ( .A(n17591), .ZN(n17946) );
  NAND3_X1 U18573 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(n17946), .ZN(n17934) );
  NOR2_X1 U18574 ( .A1(n17935), .A2(n17934), .ZN(n16411) );
  NAND2_X1 U18575 ( .A1(n17626), .A2(n16411), .ZN(n16352) );
  NAND2_X1 U18576 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17869) );
  INV_X1 U18577 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17891) );
  INV_X1 U18578 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17888) );
  NOR3_X1 U18579 ( .A1(n17869), .A2(n17891), .A3(n17888), .ZN(n16353) );
  INV_X1 U18580 ( .A(n16353), .ZN(n17865) );
  NOR2_X1 U18581 ( .A1(n16352), .A2(n17865), .ZN(n15706) );
  NAND2_X1 U18582 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18058) );
  NOR2_X1 U18583 ( .A1(n18058), .A2(n15712), .ZN(n18060) );
  NAND2_X1 U18584 ( .A1(n18060), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n18038) );
  NAND2_X1 U18585 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17677) );
  NOR2_X1 U18586 ( .A1(n18038), .A2(n17677), .ZN(n18006) );
  NAND2_X1 U18587 ( .A1(n18006), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17993) );
  INV_X1 U18588 ( .A(n17993), .ZN(n17971) );
  INV_X1 U18589 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n17783) );
  AOI22_X1 U18590 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n17158), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15542) );
  AOI22_X1 U18591 ( .A1(n17180), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15541) );
  AOI22_X1 U18592 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n9637), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15540) );
  AOI22_X1 U18593 ( .A1(n9645), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n15539) );
  NAND4_X1 U18594 ( .A1(n15542), .A2(n15541), .A3(n15540), .A4(n15539), .ZN(
        n15548) );
  AOI22_X1 U18595 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n15546) );
  AOI22_X1 U18596 ( .A1(n15584), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15545) );
  AOI22_X1 U18597 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n9639), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15544) );
  AOI22_X1 U18598 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n15543) );
  NAND4_X1 U18599 ( .A1(n15546), .A2(n15545), .A3(n15544), .A4(n15543), .ZN(
        n15547) );
  AOI22_X1 U18600 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n15552) );
  AOI22_X1 U18601 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(n9635), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15551) );
  AOI22_X1 U18602 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n15550) );
  AOI22_X1 U18603 ( .A1(n9637), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n15549) );
  NAND4_X1 U18604 ( .A1(n15552), .A2(n15551), .A3(n15550), .A4(n15549), .ZN(
        n15558) );
  AOI22_X1 U18605 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n15556) );
  AOI22_X1 U18606 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15555) );
  AOI22_X1 U18607 ( .A1(n15584), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9639), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15554) );
  AOI22_X1 U18608 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15553) );
  NAND4_X1 U18609 ( .A1(n15556), .A2(n15555), .A3(n15554), .A4(n15553), .ZN(
        n15557) );
  AOI22_X1 U18610 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15570) );
  AOI22_X1 U18611 ( .A1(n9637), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(n9635), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15569) );
  INV_X1 U18612 ( .A(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n20931) );
  AOI22_X1 U18613 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n15559), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15560) );
  OAI21_X1 U18614 ( .B1(n15595), .B2(n20931), .A(n15560), .ZN(n15567) );
  AOI22_X1 U18615 ( .A1(n14026), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15565) );
  AOI22_X1 U18616 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15561), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n15564) );
  AOI22_X1 U18617 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n15563) );
  AOI22_X1 U18618 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n15562) );
  NAND4_X1 U18619 ( .A1(n15565), .A2(n15564), .A3(n15563), .A4(n15562), .ZN(
        n15566) );
  AOI211_X1 U18620 ( .C1(n9645), .C2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A(
        n15567), .B(n15566), .ZN(n15568) );
  NAND3_X1 U18621 ( .A1(n15570), .A2(n15569), .A3(n15568), .ZN(n15680) );
  AOI22_X1 U18622 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n17164), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n15574) );
  AOI22_X1 U18623 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17144), .ZN(n15573) );
  AOI22_X1 U18624 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17157), .B1(
        n17016), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n15572) );
  AOI22_X1 U18625 ( .A1(n15584), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n17159), .ZN(n15571) );
  AOI22_X1 U18626 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n9634), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n15575) );
  OAI21_X1 U18627 ( .B1(n17221), .B2(n9675), .A(n15575), .ZN(n15576) );
  INV_X1 U18628 ( .A(n15576), .ZN(n15580) );
  AOI22_X1 U18629 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_3__1__SCAN_IN), .B2(n9637), .ZN(n15579) );
  AOI22_X1 U18630 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n9639), .ZN(n15578) );
  NAND2_X2 U18631 ( .A1(n15582), .A2(n15581), .ZN(n17375) );
  NAND2_X1 U18632 ( .A1(n15680), .A2(n17375), .ZN(n15630) );
  AOI22_X1 U18633 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n15593) );
  AOI22_X1 U18634 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n15592) );
  INV_X1 U18635 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17208) );
  AOI22_X1 U18636 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n15583) );
  OAI21_X1 U18637 ( .B1(n9675), .B2(n17208), .A(n15583), .ZN(n15590) );
  AOI22_X1 U18638 ( .A1(n14026), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n15588) );
  AOI22_X1 U18639 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9639), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15587) );
  AOI22_X1 U18640 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9637), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n15586) );
  AOI22_X1 U18641 ( .A1(n15584), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9634), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15585) );
  NAND4_X1 U18642 ( .A1(n15588), .A2(n15587), .A3(n15586), .A4(n15585), .ZN(
        n15589) );
  AOI211_X1 U18643 ( .C1(n17174), .C2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A(
        n15590), .B(n15589), .ZN(n15591) );
  NAND3_X1 U18644 ( .A1(n15593), .A2(n15592), .A3(n15591), .ZN(n15673) );
  NAND2_X1 U18645 ( .A1(n15634), .A2(n15673), .ZN(n15637) );
  AOI22_X1 U18646 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n15604) );
  AOI22_X1 U18647 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n15603) );
  AOI22_X1 U18648 ( .A1(n9637), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(n9639), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n15594) );
  OAI21_X1 U18649 ( .B1(n15595), .B2(n20948), .A(n15594), .ZN(n15601) );
  AOI22_X1 U18650 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n15599) );
  AOI22_X1 U18651 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n15598) );
  AOI22_X1 U18652 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n15597) );
  AOI22_X1 U18653 ( .A1(n9634), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n15596) );
  NAND4_X1 U18654 ( .A1(n15599), .A2(n15598), .A3(n15597), .A4(n15596), .ZN(
        n15600) );
  AOI211_X1 U18655 ( .C1(n9640), .C2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A(
        n15601), .B(n15600), .ZN(n15602) );
  NAND3_X1 U18656 ( .A1(n15604), .A2(n15603), .A3(n15602), .ZN(n15672) );
  AOI22_X1 U18657 ( .A1(n15584), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15614) );
  AOI22_X1 U18658 ( .A1(n17128), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n15613) );
  AOI22_X1 U18659 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15605) );
  OAI21_X1 U18660 ( .B1(n9675), .B2(n17197), .A(n15605), .ZN(n15611) );
  AOI22_X1 U18661 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9637), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n15609) );
  AOI22_X1 U18662 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n15608) );
  AOI22_X1 U18663 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(n9639), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15607) );
  AOI22_X1 U18664 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n15606) );
  NAND4_X1 U18665 ( .A1(n15609), .A2(n15608), .A3(n15607), .A4(n15606), .ZN(
        n15610) );
  AOI211_X1 U18666 ( .C1(n17145), .C2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A(
        n15611), .B(n15610), .ZN(n15612) );
  INV_X1 U18667 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n17827) );
  INV_X1 U18668 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18793) );
  NOR2_X1 U18669 ( .A1(n17375), .A2(n18793), .ZN(n15626) );
  XOR2_X2 U18670 ( .A(n17375), .B(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .Z(
        n17850) );
  AOI22_X1 U18671 ( .A1(n9645), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17173), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n15625) );
  AOI22_X1 U18672 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9639), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15624) );
  AOI22_X1 U18673 ( .A1(n17180), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n15616) );
  OAI21_X1 U18674 ( .B1(n15538), .B2(n20908), .A(n15616), .ZN(n15622) );
  AOI22_X1 U18675 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(n9634), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15620) );
  AOI22_X1 U18676 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n15619) );
  AOI22_X1 U18677 ( .A1(n15584), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n15618) );
  AOI22_X1 U18678 ( .A1(n17016), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n17157), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n15617) );
  NAND4_X1 U18679 ( .A1(n15620), .A2(n15619), .A3(n15618), .A4(n15617), .ZN(
        n15621) );
  AOI211_X1 U18680 ( .C1(n9637), .C2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A(
        n15622), .B(n15621), .ZN(n15623) );
  NAND3_X1 U18681 ( .A1(n15625), .A2(n15624), .A3(n15623), .ZN(n17858) );
  NAND2_X1 U18682 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17858), .ZN(
        n17857) );
  NOR2_X1 U18683 ( .A1(n17850), .A2(n17857), .ZN(n17849) );
  NOR2_X1 U18684 ( .A1(n15627), .A2(n15628), .ZN(n15629) );
  XNOR2_X1 U18685 ( .A(n17364), .B(n15630), .ZN(n15631) );
  NOR2_X1 U18686 ( .A1(n15632), .A2(n15631), .ZN(n15633) );
  INV_X1 U18687 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18135) );
  XOR2_X1 U18688 ( .A(n15673), .B(n15634), .Z(n15635) );
  XOR2_X1 U18689 ( .A(n18135), .B(n15635), .Z(n17815) );
  XNOR2_X1 U18690 ( .A(n17356), .B(n15637), .ZN(n15638) );
  INV_X1 U18691 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n17802) );
  INV_X1 U18692 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18113) );
  XOR2_X1 U18693 ( .A(n15672), .B(n15641), .Z(n15642) );
  XOR2_X1 U18694 ( .A(n18113), .B(n15642), .Z(n17787) );
  NOR2_X1 U18695 ( .A1(n17783), .A2(n17782), .ZN(n17781) );
  INV_X1 U18696 ( .A(n17781), .ZN(n15645) );
  INV_X1 U18697 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n18092) );
  NAND2_X2 U18698 ( .A1(n15711), .A2(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n18051) );
  NAND2_X1 U18699 ( .A1(n17971), .A2(n17679), .ZN(n18004) );
  NAND2_X1 U18700 ( .A1(n15706), .A2(n17924), .ZN(n17870) );
  INV_X1 U18701 ( .A(n16411), .ZN(n15646) );
  NOR3_X1 U18702 ( .A1(n17802), .A2(n17827), .A3(n18135), .ZN(n17969) );
  AOI21_X1 U18703 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n18152) );
  INV_X1 U18704 ( .A(n18152), .ZN(n18132) );
  NAND2_X1 U18705 ( .A1(n17969), .A2(n18132), .ZN(n18086) );
  NAND2_X1 U18706 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18090) );
  NOR3_X1 U18707 ( .A1(n18092), .A2(n18086), .A3(n18090), .ZN(n17991) );
  NAND3_X1 U18708 ( .A1(n17971), .A2(n17626), .A3(n17991), .ZN(n17973) );
  NOR2_X1 U18709 ( .A1(n15646), .A2(n17973), .ZN(n17890) );
  INV_X1 U18710 ( .A(n17890), .ZN(n17908) );
  AND2_X1 U18711 ( .A1(n15648), .A2(n15647), .ZN(n18845) );
  NAND2_X1 U18712 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18131) );
  INV_X1 U18713 ( .A(n18131), .ZN(n15650) );
  NAND2_X1 U18714 ( .A1(n17969), .A2(n15650), .ZN(n18085) );
  NOR2_X1 U18715 ( .A1(n18090), .A2(n18085), .ZN(n17992) );
  AND2_X1 U18716 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17992), .ZN(
        n17940) );
  NAND2_X1 U18717 ( .A1(n17971), .A2(n17940), .ZN(n17972) );
  NOR2_X1 U18718 ( .A1(n17977), .A2(n17972), .ZN(n17867) );
  NAND2_X1 U18719 ( .A1(n16411), .A2(n17867), .ZN(n15657) );
  NOR2_X2 U18720 ( .A1(n15651), .A2(n15655), .ZN(n18176) );
  INV_X1 U18721 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18810) );
  NOR2_X1 U18722 ( .A1(n18810), .A2(n15657), .ZN(n17866) );
  INV_X1 U18723 ( .A(n17866), .ZN(n15656) );
  AOI21_X1 U18724 ( .B1(n15654), .B2(n15653), .A(n15652), .ZN(n18645) );
  OAI21_X2 U18725 ( .B1(n18646), .B2(n15655), .A(n18645), .ZN(n18636) );
  OAI222_X1 U18726 ( .A1(n17908), .A2(n18661), .B1(n15657), .B2(n18176), .C1(
        n15656), .C2(n18635), .ZN(n17893) );
  NAND2_X1 U18727 ( .A1(n16353), .A2(n17893), .ZN(n16385) );
  NOR2_X1 U18728 ( .A1(n18208), .A2(n18834), .ZN(n15662) );
  AND2_X1 U18729 ( .A1(n18228), .A2(n15662), .ZN(n15669) );
  NAND2_X1 U18730 ( .A1(n15669), .A2(n15658), .ZN(n16398) );
  NOR2_X1 U18731 ( .A1(n16398), .A2(n16400), .ZN(n18052) );
  AOI21_X1 U18732 ( .B1(n15661), .B2(n15660), .A(n15659), .ZN(n18628) );
  INV_X1 U18733 ( .A(n18628), .ZN(n15668) );
  AOI21_X1 U18734 ( .B1(n18208), .B2(n18834), .A(n15662), .ZN(n15663) );
  AOI21_X1 U18735 ( .B1(n18832), .B2(n15663), .A(n18829), .ZN(n16514) );
  INV_X1 U18736 ( .A(n16514), .ZN(n15664) );
  NOR2_X1 U18737 ( .A1(n18626), .A2(n15664), .ZN(n15666) );
  MUX2_X1 U18738 ( .A(n18631), .B(n15666), .S(n15665), .Z(n15667) );
  AOI21_X1 U18739 ( .B1(n15669), .B2(n15668), .A(n15667), .ZN(n15670) );
  AOI221_X1 U18740 ( .B1(n17870), .B2(n16385), .C1(n18031), .C2(n16385), .A(
        n18166), .ZN(n15705) );
  NOR2_X4 U18741 ( .A1(n18655), .A2(n18153), .ZN(n18061) );
  NAND2_X1 U18742 ( .A1(n18054), .A2(n18175), .ZN(n18141) );
  INV_X1 U18743 ( .A(n15672), .ZN(n17353) );
  INV_X1 U18744 ( .A(n15673), .ZN(n17360) );
  INV_X1 U18745 ( .A(n15680), .ZN(n17370) );
  NAND2_X1 U18746 ( .A1(n17858), .A2(n17375), .ZN(n15679) );
  NAND2_X1 U18747 ( .A1(n17370), .A2(n15679), .ZN(n15678) );
  INV_X1 U18748 ( .A(n17364), .ZN(n15677) );
  NAND2_X1 U18749 ( .A1(n15678), .A2(n15677), .ZN(n15690) );
  INV_X1 U18750 ( .A(n17356), .ZN(n15674) );
  NAND2_X1 U18751 ( .A1(n15675), .A2(n15674), .ZN(n15693) );
  NOR2_X1 U18752 ( .A1(n17353), .A2(n15693), .ZN(n15697) );
  NAND2_X1 U18753 ( .A1(n15697), .A2(n16400), .ZN(n15698) );
  XOR2_X1 U18754 ( .A(n15675), .B(n15674), .Z(n15676) );
  XOR2_X1 U18755 ( .A(n17802), .B(n15676), .Z(n17799) );
  XNOR2_X1 U18756 ( .A(n15678), .B(n15677), .ZN(n15688) );
  NOR2_X1 U18757 ( .A1(n15688), .A2(n17827), .ZN(n15689) );
  XNOR2_X1 U18758 ( .A(n15680), .B(n15679), .ZN(n15685) );
  NOR2_X1 U18759 ( .A1(n15685), .A2(n15627), .ZN(n15687) );
  INV_X1 U18760 ( .A(n17375), .ZN(n15682) );
  NOR2_X1 U18761 ( .A1(n15682), .A2(n18810), .ZN(n15684) );
  INV_X1 U18762 ( .A(n17858), .ZN(n15683) );
  NAND3_X1 U18763 ( .A1(n15683), .A2(n15682), .A3(n18810), .ZN(n15681) );
  OAI221_X1 U18764 ( .B1(n15684), .B2(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C1(
        n15683), .C2(n15682), .A(n15681), .ZN(n17840) );
  XOR2_X1 U18765 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n15685), .Z(
        n17839) );
  NOR2_X1 U18766 ( .A1(n17840), .A2(n17839), .ZN(n15686) );
  NOR2_X1 U18767 ( .A1(n15687), .A2(n15686), .ZN(n17830) );
  XOR2_X1 U18768 ( .A(n15688), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(
        n17829) );
  NOR2_X1 U18769 ( .A1(n17830), .A2(n17829), .ZN(n17828) );
  NOR2_X1 U18770 ( .A1(n15689), .A2(n17828), .ZN(n17811) );
  XNOR2_X1 U18771 ( .A(n15690), .B(n17360), .ZN(n17812) );
  NOR2_X1 U18772 ( .A1(n17811), .A2(n17812), .ZN(n15691) );
  NAND2_X1 U18773 ( .A1(n17811), .A2(n17812), .ZN(n17810) );
  OAI21_X1 U18774 ( .B1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n15691), .A(
        n17810), .ZN(n17798) );
  XNOR2_X1 U18775 ( .A(n15693), .B(n17353), .ZN(n15695) );
  NOR2_X1 U18776 ( .A1(n15694), .A2(n15695), .ZN(n15696) );
  XNOR2_X1 U18777 ( .A(n15695), .B(n15694), .ZN(n17793) );
  NOR2_X1 U18778 ( .A1(n15696), .A2(n17792), .ZN(n15699) );
  XOR2_X1 U18779 ( .A(n15697), .B(n17349), .Z(n15700) );
  NAND2_X1 U18780 ( .A1(n15699), .A2(n15700), .ZN(n17778) );
  NAND2_X1 U18781 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17778), .ZN(
        n15702) );
  NOR2_X1 U18782 ( .A1(n15698), .A2(n15702), .ZN(n15704) );
  INV_X1 U18783 ( .A(n15698), .ZN(n15703) );
  OR2_X1 U18784 ( .A1(n15700), .A2(n15699), .ZN(n17779) );
  OAI21_X1 U18785 ( .B1(n15703), .B2(n15702), .A(n17779), .ZN(n15701) );
  AOI21_X1 U18786 ( .B1(n15703), .B2(n15702), .A(n15701), .ZN(n17766) );
  NAND2_X1 U18787 ( .A1(n18015), .A2(n15706), .ZN(n17871) );
  NOR2_X1 U18788 ( .A1(n17871), .A2(n16377), .ZN(n16403) );
  AOI22_X1 U18789 ( .A1(n15709), .A2(n15705), .B1(n18179), .B2(n16403), .ZN(
        n15825) );
  NOR3_X1 U18790 ( .A1(n18844), .A2(P3_STATE2_REG_0__SCAN_IN), .A3(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n16412) );
  INV_X1 U18791 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n16408) );
  NAND3_X1 U18792 ( .A1(n16353), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        n17866), .ZN(n15708) );
  INV_X1 U18793 ( .A(n17972), .ZN(n17926) );
  AOI21_X1 U18794 ( .B1(n15706), .B2(n17926), .A(n18176), .ZN(n15707) );
  AOI21_X1 U18795 ( .B1(n16353), .B2(n17890), .A(n18661), .ZN(n17874) );
  AOI211_X1 U18796 ( .C1(n18636), .C2(n15708), .A(n15707), .B(n17874), .ZN(
        n15819) );
  OAI21_X1 U18797 ( .B1(n18061), .B2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15819), .ZN(n16405) );
  AOI211_X1 U18798 ( .C1(n17996), .C2(n16408), .A(n18166), .B(n16405), .ZN(
        n15710) );
  NAND2_X1 U18799 ( .A1(n18175), .A2(n18052), .ZN(n18099) );
  INV_X1 U18800 ( .A(n18099), .ZN(n16391) );
  NAND2_X1 U18801 ( .A1(n15709), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16387) );
  NOR2_X1 U18802 ( .A1(n16387), .A2(n17870), .ZN(n16360) );
  INV_X1 U18803 ( .A(n16360), .ZN(n16378) );
  NOR2_X1 U18804 ( .A1(n17871), .A2(n16387), .ZN(n16361) );
  INV_X1 U18805 ( .A(n16361), .ZN(n16379) );
  AOI22_X1 U18806 ( .A1(n16391), .A2(n16378), .B1(n18179), .B2(n16379), .ZN(
        n15822) );
  OAI21_X1 U18807 ( .B1(n16412), .B2(n15710), .A(n15822), .ZN(n15726) );
  INV_X1 U18808 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18072) );
  AND2_X1 U18809 ( .A1(n18072), .A2(n15712), .ZN(n15713) );
  INV_X1 U18810 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17693) );
  NAND2_X1 U18811 ( .A1(n17707), .A2(n17693), .ZN(n17664) );
  NOR2_X1 U18812 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15714) );
  AND2_X2 U18813 ( .A1(n15715), .A2(n18051), .ZN(n17768) );
  INV_X1 U18814 ( .A(n15720), .ZN(n17644) );
  INV_X1 U18815 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n18001) );
  INV_X1 U18816 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17983) );
  NAND2_X2 U18817 ( .A1(n17632), .A2(n17587), .ZN(n17604) );
  INV_X1 U18818 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17907) );
  NOR2_X1 U18819 ( .A1(n16352), .A2(n17907), .ZN(n17551) );
  NAND2_X1 U18820 ( .A1(n15720), .A2(n17551), .ZN(n15718) );
  INV_X1 U18821 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17962) );
  NAND2_X1 U18822 ( .A1(n17627), .A2(n17962), .ZN(n15717) );
  INV_X1 U18823 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17594) );
  NAND2_X1 U18824 ( .A1(n17589), .A2(n17594), .ZN(n17568) );
  NAND2_X1 U18825 ( .A1(n17626), .A2(n15720), .ZN(n17586) );
  INV_X1 U18826 ( .A(n17520), .ZN(n15723) );
  NOR2_X1 U18827 ( .A1(n17539), .A2(n17587), .ZN(n15721) );
  NAND2_X1 U18828 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17875) );
  AOI21_X2 U18829 ( .B1(n15723), .B2(n17888), .A(n15722), .ZN(n16397) );
  AND2_X2 U18830 ( .A1(n16397), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n17510) );
  NOR2_X1 U18831 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17587), .ZN(
        n15724) );
  AOI21_X1 U18832 ( .B1(n15817), .B2(n16401), .A(n15724), .ZN(n15725) );
  XOR2_X1 U18833 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B(n15725), .Z(
        n16376) );
  AOI22_X1 U18834 ( .A1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(n15726), .B1(
        n9743), .B2(n16376), .ZN(n15727) );
  INV_X2 U18835 ( .A(n9642), .ZN(n18174) );
  NAND2_X1 U18836 ( .A1(n18174), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16372) );
  OAI211_X1 U18837 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n15825), .A(
        n15727), .B(n16372), .ZN(P3_U2833) );
  OAI22_X1 U18838 ( .A1(n19104), .A2(n10897), .B1(n19816), .B2(n19110), .ZN(
        n15732) );
  INV_X1 U18839 ( .A(n15728), .ZN(n15730) );
  INV_X1 U18840 ( .A(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15729) );
  OAI22_X1 U18841 ( .A1(n15730), .A2(n19086), .B1(n19101), .B2(n15729), .ZN(
        n15731) );
  AOI211_X1 U18842 ( .C1(n15733), .C2(n19099), .A(n15732), .B(n15731), .ZN(
        n15758) );
  OAI21_X1 U18843 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n15735), .A(
        n15734), .ZN(n16228) );
  INV_X1 U18844 ( .A(n15736), .ZN(n18917) );
  INV_X1 U18845 ( .A(n15737), .ZN(n18967) );
  OAI21_X1 U18846 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n9701), .A(
        n15749), .ZN(n16244) );
  INV_X1 U18847 ( .A(n16244), .ZN(n18988) );
  OAI21_X1 U18848 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n15744), .A(
        n15748), .ZN(n19014) );
  INV_X1 U18849 ( .A(n19014), .ZN(n15747) );
  AOI21_X1 U18850 ( .B1(n16278), .B2(n15739), .A(n15738), .ZN(n19036) );
  AOI21_X1 U18851 ( .B1(n19052), .B2(n15741), .A(n15740), .ZN(n19058) );
  NAND2_X1 U18852 ( .A1(n15743), .A2(n15742), .ZN(n19079) );
  NOR2_X1 U18853 ( .A1(n19081), .A2(n19079), .ZN(n19071) );
  NAND2_X1 U18854 ( .A1(n19071), .A2(n19072), .ZN(n19056) );
  NOR2_X1 U18855 ( .A1(n19058), .A2(n19056), .ZN(n19044) );
  NAND2_X1 U18856 ( .A1(n19044), .A2(n19045), .ZN(n19034) );
  NOR2_X1 U18857 ( .A1(n19036), .A2(n19034), .ZN(n19023) );
  AOI21_X1 U18858 ( .B1(n16265), .B2(n15745), .A(n15744), .ZN(n19024) );
  INV_X1 U18859 ( .A(n19024), .ZN(n15746) );
  NAND2_X1 U18860 ( .A1(n19023), .A2(n15746), .ZN(n19012) );
  NOR2_X1 U18861 ( .A1(n15747), .A2(n19012), .ZN(n19005) );
  AOI21_X1 U18862 ( .B1(n16251), .B2(n15748), .A(n9701), .ZN(n16245) );
  INV_X1 U18863 ( .A(n16245), .ZN(n19008) );
  NAND2_X1 U18864 ( .A1(n19005), .A2(n19008), .ZN(n18987) );
  NOR2_X1 U18865 ( .A1(n18988), .A2(n18987), .ZN(n18983) );
  AND2_X1 U18866 ( .A1(n15749), .A2(n16236), .ZN(n15751) );
  OR2_X1 U18867 ( .A1(n15751), .A2(n15750), .ZN(n18982) );
  NAND2_X1 U18868 ( .A1(n18983), .A2(n18982), .ZN(n18966) );
  NOR2_X1 U18869 ( .A1(n18967), .A2(n18966), .ZN(n18958) );
  INV_X1 U18870 ( .A(n18959), .ZN(n15752) );
  NAND2_X1 U18871 ( .A1(n18958), .A2(n15752), .ZN(n18946) );
  NOR2_X1 U18872 ( .A1(n15753), .A2(n18946), .ZN(n18930) );
  NAND2_X1 U18873 ( .A1(n18930), .A2(n18940), .ZN(n18928) );
  NOR2_X1 U18874 ( .A1(n18917), .A2(n18928), .ZN(n18908) );
  INV_X1 U18875 ( .A(n18909), .ZN(n15754) );
  NAND2_X1 U18876 ( .A1(n18908), .A2(n15754), .ZN(n18891) );
  INV_X1 U18877 ( .A(n18897), .ZN(n18892) );
  INV_X1 U18878 ( .A(n15755), .ZN(n18886) );
  NAND2_X1 U18879 ( .A1(n19080), .A2(n18885), .ZN(n15756) );
  NAND2_X1 U18880 ( .A1(n16228), .A2(n15756), .ZN(n16116) );
  OAI211_X1 U18881 ( .C1(n16228), .C2(n15756), .A(n19076), .B(n16116), .ZN(
        n15757) );
  OAI211_X1 U18882 ( .C1(n19091), .C2(n16222), .A(n15758), .B(n15757), .ZN(
        P2_U2833) );
  NAND2_X1 U18883 ( .A1(n15760), .A2(n15759), .ZN(n15770) );
  AND2_X1 U18884 ( .A1(n15762), .A2(n15761), .ZN(n15763) );
  OR2_X1 U18885 ( .A1(n15764), .A2(n15763), .ZN(n15766) );
  OAI21_X1 U18886 ( .B1(n15766), .B2(n20553), .A(n15765), .ZN(n15769) );
  INV_X1 U18887 ( .A(n15766), .ZN(n15767) );
  AOI22_X1 U18888 ( .A1(n15770), .A2(n15769), .B1(n15768), .B2(n15767), .ZN(
        n15772) );
  NAND2_X1 U18889 ( .A1(n15772), .A2(n20502), .ZN(n15774) );
  OAI21_X1 U18890 ( .B1(n15772), .B2(n20502), .A(n15771), .ZN(n15773) );
  OAI211_X1 U18891 ( .C1(n15775), .C2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n15774), .B(n15773), .ZN(n15776) );
  OAI21_X1 U18892 ( .B1(n15777), .B2(n20501), .A(n15776), .ZN(n15787) );
  INV_X1 U18893 ( .A(n15778), .ZN(n15783) );
  INV_X1 U18894 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n15780) );
  AOI21_X1 U18895 ( .B1(n19919), .B2(n15780), .A(n15779), .ZN(n15781) );
  NOR4_X1 U18896 ( .A1(n15784), .A2(n15783), .A3(n15782), .A4(n15781), .ZN(
        n15785) );
  OAI211_X1 U18897 ( .C1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n15787), .A(
        n15786), .B(n15785), .ZN(n15797) );
  INV_X1 U18898 ( .A(n15788), .ZN(n15795) );
  NAND2_X1 U18899 ( .A1(n20761), .A2(n15789), .ZN(n15790) );
  NOR2_X1 U18900 ( .A1(n15791), .A2(n15790), .ZN(n15794) );
  NOR3_X1 U18901 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n20760), .A3(n20767), 
        .ZN(n15792) );
  NOR2_X1 U18902 ( .A1(n15798), .A2(n15792), .ZN(n15793) );
  AOI21_X1 U18903 ( .B1(n15795), .B2(n15794), .A(n15793), .ZN(n16109) );
  INV_X1 U18904 ( .A(n16109), .ZN(n15796) );
  AOI221_X1 U18905 ( .B1(n9755), .B2(n20669), .C1(n15797), .C2(n20669), .A(
        n15796), .ZN(n15799) );
  NOR2_X1 U18906 ( .A1(n15799), .A2(n9755), .ZN(n16115) );
  OAI21_X1 U18907 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n20767), .A(n16115), 
        .ZN(n16113) );
  AOI211_X1 U18908 ( .C1(n15798), .C2(n15797), .A(n16111), .B(n16113), .ZN(
        n15805) );
  AOI21_X1 U18909 ( .B1(n15801), .B2(n15800), .A(n15799), .ZN(n15802) );
  INV_X1 U18910 ( .A(n15802), .ZN(n15803) );
  AOI22_X1 U18911 ( .A1(n15805), .A2(n15804), .B1(n9755), .B2(n15803), .ZN(
        P1_U3161) );
  AOI22_X1 U18912 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15806), .B1(
        n20162), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15815) );
  NOR3_X1 U18913 ( .A1(n14571), .A2(n15808), .A3(n15807), .ZN(n15809) );
  AOI21_X1 U18914 ( .B1(n15811), .B2(n15810), .A(n15809), .ZN(n15812) );
  XNOR2_X1 U18915 ( .A(n15812), .B(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n15906) );
  AOI22_X1 U18916 ( .A1(n15906), .A2(n20160), .B1(n20157), .B2(n15813), .ZN(
        n15814) );
  OAI211_X1 U18917 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15816), .A(
        n15815), .B(n15814), .ZN(P1_U3010) );
  OR2_X1 U18918 ( .A1(n16387), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16366) );
  INV_X1 U18919 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n15821) );
  INV_X1 U18920 ( .A(n17996), .ZN(n18134) );
  NOR2_X1 U18921 ( .A1(n18166), .A2(n18134), .ZN(n18169) );
  INV_X1 U18922 ( .A(n18168), .ZN(n18162) );
  OAI21_X1 U18923 ( .B1(n15819), .B2(n18166), .A(n18162), .ZN(n15820) );
  AOI21_X1 U18924 ( .B1(n18169), .B2(n16387), .A(n15820), .ZN(n16383) );
  AOI21_X1 U18925 ( .B1(n16383), .B2(n15822), .A(n15821), .ZN(n15823) );
  AOI21_X1 U18926 ( .B1(n9743), .B2(n16362), .A(n15823), .ZN(n15824) );
  NAND2_X1 U18927 ( .A1(n16412), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16355) );
  OAI211_X1 U18928 ( .C1(n15825), .C2(n16366), .A(n15824), .B(n16355), .ZN(
        P3_U2832) );
  INV_X1 U18929 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n20688) );
  INV_X1 U18930 ( .A(HOLD), .ZN(n20687) );
  NOR2_X1 U18931 ( .A1(n20688), .A2(n20687), .ZN(n20676) );
  AOI22_X1 U18932 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(HOLD), .B1(
        P1_STATE_REG_0__SCAN_IN), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n15827) );
  NOR2_X1 U18933 ( .A1(n20674), .A2(n20767), .ZN(n20683) );
  INV_X1 U18934 ( .A(n20683), .ZN(n20673) );
  OAI211_X1 U18935 ( .C1(n20676), .C2(n15827), .A(n15826), .B(n20673), .ZN(
        P1_U3195) );
  AND2_X1 U18936 ( .A1(n20064), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  OAI221_X1 U18937 ( .B1(P2_STATE2_REG_0__SCAN_IN), .B2(n19896), .C1(n18853), 
        .C2(n16324), .A(n19691), .ZN(n19757) );
  NAND2_X1 U18938 ( .A1(n15828), .A2(n19691), .ZN(n16327) );
  AND3_X1 U18939 ( .A1(n19757), .A2(n16327), .A3(n15829), .ZN(P2_U3178) );
  OAI221_X1 U18940 ( .B1(n18860), .B2(n15829), .C1(n19885), .C2(n15829), .A(
        n19614), .ZN(n19878) );
  NOR2_X1 U18941 ( .A1(n15830), .A2(n19878), .ZN(P2_U3047) );
  OAI33_X1 U18942 ( .A1(n18196), .A2(n18204), .A3(n15833), .B1(n15832), .B2(
        n18675), .B3(n15831), .ZN(n17229) );
  NAND2_X1 U18943 ( .A1(n17074), .A2(n9654), .ZN(n17378) );
  INV_X1 U18944 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17455) );
  NAND2_X1 U18945 ( .A1(n18634), .A2(n17368), .ZN(n17374) );
  NAND2_X1 U18946 ( .A1(n15834), .A2(n9654), .ZN(n17371) );
  AOI22_X1 U18947 ( .A1(n17377), .A2(BUF2_REG_0__SCAN_IN), .B1(n17376), .B2(
        n17858), .ZN(n15835) );
  OAI221_X1 U18948 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17378), .C1(n17455), 
        .C2(n9654), .A(n15835), .ZN(P3_U2735) );
  AOI22_X1 U18949 ( .A1(n20026), .A2(P1_EBX_REG_20__SCAN_IN), .B1(n20014), 
        .B2(n15836), .ZN(n15844) );
  INV_X1 U18950 ( .A(n15837), .ZN(n15847) );
  NAND2_X1 U18951 ( .A1(n15847), .A2(n15895), .ZN(n15863) );
  OAI21_X1 U18952 ( .B1(n15846), .B2(n15863), .A(n20713), .ZN(n15841) );
  OAI22_X1 U18953 ( .A1(n15839), .A2(n19942), .B1(n20008), .B2(n15838), .ZN(
        n15840) );
  AOI21_X1 U18954 ( .B1(n15842), .B2(n15841), .A(n15840), .ZN(n15843) );
  OAI211_X1 U18955 ( .C1(n15845), .C2(n20031), .A(n15844), .B(n15843), .ZN(
        P1_U2820) );
  OAI21_X1 U18956 ( .B1(P1_REIP_REG_19__SCAN_IN), .B2(P1_REIP_REG_18__SCAN_IN), 
        .A(n15846), .ZN(n15854) );
  AOI21_X1 U18957 ( .B1(n15848), .B2(n15847), .A(n15899), .ZN(n15865) );
  AOI22_X1 U18958 ( .A1(n15865), .A2(P1_REIP_REG_19__SCAN_IN), .B1(n20026), 
        .B2(P1_EBX_REG_19__SCAN_IN), .ZN(n15849) );
  OAI21_X1 U18959 ( .B1(n15918), .B2(n20042), .A(n15849), .ZN(n15850) );
  AOI211_X1 U18960 ( .C1(n20013), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n20001), .B(n15850), .ZN(n15853) );
  OAI22_X1 U18961 ( .A1(n15914), .A2(n19942), .B1(n20008), .B2(n15994), .ZN(
        n15851) );
  INV_X1 U18962 ( .A(n15851), .ZN(n15852) );
  OAI211_X1 U18963 ( .C1(n15863), .C2(n15854), .A(n15853), .B(n15852), .ZN(
        P1_U2821) );
  INV_X1 U18964 ( .A(n15855), .ZN(n15857) );
  AOI22_X1 U18965 ( .A1(n15865), .A2(P1_REIP_REG_18__SCAN_IN), .B1(n20026), 
        .B2(P1_EBX_REG_18__SCAN_IN), .ZN(n15856) );
  OAI21_X1 U18966 ( .B1(n15857), .B2(n20042), .A(n15856), .ZN(n15858) );
  AOI211_X1 U18967 ( .C1(n20013), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n20001), .B(n15858), .ZN(n15862) );
  AOI22_X1 U18968 ( .A1(n15860), .A2(n19978), .B1(n20034), .B2(n15859), .ZN(
        n15861) );
  OAI211_X1 U18969 ( .C1(P1_REIP_REG_18__SCAN_IN), .C2(n15863), .A(n15862), 
        .B(n15861), .ZN(P1_U2822) );
  AOI22_X1 U18970 ( .A1(n20026), .A2(P1_EBX_REG_17__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n20013), .ZN(n15870) );
  AOI21_X1 U18971 ( .B1(n20014), .B2(n15925), .A(n20001), .ZN(n15869) );
  INV_X1 U18972 ( .A(n15864), .ZN(n15926) );
  AOI22_X1 U18973 ( .A1(n15926), .A2(n19978), .B1(n20034), .B2(n16002), .ZN(
        n15868) );
  OAI221_X1 U18974 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(P1_REIP_REG_16__SCAN_IN), .C1(P1_REIP_REG_17__SCAN_IN), .C2(n15866), .A(n15865), .ZN(n15867) );
  NAND4_X1 U18975 ( .A1(n15870), .A2(n15869), .A3(n15868), .A4(n15867), .ZN(
        P1_U2823) );
  AOI22_X1 U18976 ( .A1(n16015), .A2(n20034), .B1(n20014), .B2(n15934), .ZN(
        n15876) );
  AOI22_X1 U18977 ( .A1(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n20013), .B1(
        P1_REIP_REG_15__SCAN_IN), .B2(n15871), .ZN(n15875) );
  AOI21_X1 U18978 ( .B1(n20026), .B2(P1_EBX_REG_15__SCAN_IN), .A(n20001), .ZN(
        n15874) );
  AOI21_X1 U18979 ( .B1(n15935), .B2(n19978), .A(n15872), .ZN(n15873) );
  NAND4_X1 U18980 ( .A1(n15876), .A2(n15875), .A3(n15874), .A4(n15873), .ZN(
        P1_U2825) );
  INV_X1 U18981 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n16031) );
  NAND2_X1 U18982 ( .A1(n15880), .A2(n16031), .ZN(n15883) );
  INV_X1 U18983 ( .A(n15877), .ZN(n16033) );
  AOI22_X1 U18984 ( .A1(n20026), .A2(P1_EBX_REG_13__SCAN_IN), .B1(n20014), 
        .B2(n15945), .ZN(n15878) );
  OAI21_X1 U18985 ( .B1(n16033), .B2(n20008), .A(n15878), .ZN(n15879) );
  AOI211_X1 U18986 ( .C1(n20013), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n20001), .B(n15879), .ZN(n15882) );
  AOI21_X1 U18987 ( .B1(n15900), .B2(n15880), .A(n15899), .ZN(n15891) );
  AOI22_X1 U18988 ( .A1(n15946), .A2(n19978), .B1(n15891), .B2(
        P1_REIP_REG_13__SCAN_IN), .ZN(n15881) );
  OAI211_X1 U18989 ( .C1(n15888), .C2(n15883), .A(n15882), .B(n15881), .ZN(
        P1_U2827) );
  INV_X1 U18990 ( .A(n15884), .ZN(n15951) );
  AOI22_X1 U18991 ( .A1(n20026), .A2(P1_EBX_REG_12__SCAN_IN), .B1(n15951), 
        .B2(n20014), .ZN(n15894) );
  INV_X1 U18992 ( .A(n15885), .ZN(n16048) );
  AOI22_X1 U18993 ( .A1(n16048), .A2(n20034), .B1(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n20013), .ZN(n15893) );
  INV_X1 U18994 ( .A(n15886), .ZN(n15952) );
  OAI21_X1 U18995 ( .B1(n15889), .B2(n15888), .A(n15887), .ZN(n15890) );
  AOI22_X1 U18996 ( .A1(n15952), .A2(n19978), .B1(n15891), .B2(n15890), .ZN(
        n15892) );
  NAND4_X1 U18997 ( .A1(n15894), .A2(n15893), .A3(n15892), .A4(n19974), .ZN(
        P1_U2828) );
  NAND2_X1 U18998 ( .A1(P1_REIP_REG_9__SCAN_IN), .A2(n15895), .ZN(n15904) );
  INV_X1 U18999 ( .A(n15896), .ZN(n16077) );
  AOI22_X1 U19000 ( .A1(n20026), .A2(P1_EBX_REG_10__SCAN_IN), .B1(n20014), 
        .B2(n15960), .ZN(n15897) );
  OAI21_X1 U19001 ( .B1(n16077), .B2(n20008), .A(n15897), .ZN(n15898) );
  AOI211_X1 U19002 ( .C1(n20013), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n20001), .B(n15898), .ZN(n15903) );
  NOR3_X1 U19003 ( .A1(n15900), .A2(n15899), .A3(n16076), .ZN(n15901) );
  AOI21_X1 U19004 ( .B1(n15962), .B2(n19978), .A(n15901), .ZN(n15902) );
  OAI211_X1 U19005 ( .C1(P1_REIP_REG_10__SCAN_IN), .C2(n15904), .A(n15903), 
        .B(n15902), .ZN(P1_U2830) );
  AOI22_X1 U19006 ( .A1(n20120), .A2(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B1(
        n20162), .B2(P1_REIP_REG_21__SCAN_IN), .ZN(n15909) );
  INV_X1 U19007 ( .A(n15905), .ZN(n15907) );
  AOI22_X1 U19008 ( .A1(n15907), .A2(n20125), .B1(n15906), .B2(n12697), .ZN(
        n15908) );
  OAI211_X1 U19009 ( .C1(n20130), .C2(n15910), .A(n15909), .B(n15908), .ZN(
        P1_U2978) );
  AOI22_X1 U19010 ( .A1(n20120), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n20162), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15917) );
  NOR2_X1 U19011 ( .A1(n15955), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n15911) );
  MUX2_X1 U19012 ( .A(n15955), .B(n15911), .S(n14571), .Z(n15913) );
  XNOR2_X1 U19013 ( .A(n15913), .B(n15912), .ZN(n15996) );
  INV_X1 U19014 ( .A(n15914), .ZN(n15915) );
  AOI22_X1 U19015 ( .A1(n15996), .A2(n12697), .B1(n15915), .B2(n20125), .ZN(
        n15916) );
  OAI211_X1 U19016 ( .C1(n20130), .C2(n15918), .A(n15917), .B(n15916), .ZN(
        P1_U2980) );
  NOR2_X1 U19017 ( .A1(n15955), .A2(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15923) );
  AOI21_X1 U19018 ( .B1(n15921), .B2(n15920), .A(n15919), .ZN(n15922) );
  MUX2_X1 U19019 ( .A(n15923), .B(n15955), .S(n15922), .Z(n15924) );
  XOR2_X1 U19020 ( .A(n16000), .B(n15924), .Z(n16007) );
  AOI22_X1 U19021 ( .A1(n20120), .A2(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n20162), .B2(P1_REIP_REG_17__SCAN_IN), .ZN(n15928) );
  AOI22_X1 U19022 ( .A1(n15926), .A2(n20125), .B1(n15925), .B2(n15961), .ZN(
        n15927) );
  OAI211_X1 U19023 ( .C1(n19918), .C2(n16007), .A(n15928), .B(n15927), .ZN(
        P1_U2982) );
  INV_X1 U19024 ( .A(n15929), .ZN(n15930) );
  OAI21_X1 U19025 ( .B1(n12600), .B2(n15955), .A(n15930), .ZN(n15932) );
  AOI21_X1 U19026 ( .B1(n15933), .B2(n15932), .A(n15931), .ZN(n16020) );
  AOI22_X1 U19027 ( .A1(n20120), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n20162), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n15937) );
  AOI22_X1 U19028 ( .A1(n15935), .A2(n20125), .B1(n15961), .B2(n15934), .ZN(
        n15936) );
  OAI211_X1 U19029 ( .C1(n16020), .C2(n19918), .A(n15937), .B(n15936), .ZN(
        P1_U2984) );
  OAI22_X1 U19030 ( .A1(n15956), .A2(n15939), .B1(n15938), .B2(n15955), .ZN(
        n15949) );
  NAND2_X1 U19031 ( .A1(n9985), .A2(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n15940) );
  NAND2_X1 U19032 ( .A1(n15940), .A2(n9759), .ZN(n15950) );
  NOR2_X1 U19033 ( .A1(n15949), .A2(n15950), .ZN(n15941) );
  NOR2_X1 U19034 ( .A1(n15942), .A2(n15941), .ZN(n15944) );
  XOR2_X1 U19035 ( .A(n15944), .B(n15943), .Z(n16047) );
  AOI22_X1 U19036 ( .A1(n20120), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n20162), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n15948) );
  AOI22_X1 U19037 ( .A1(n15946), .A2(n20125), .B1(n15961), .B2(n15945), .ZN(
        n15947) );
  OAI211_X1 U19038 ( .C1(n19918), .C2(n16047), .A(n15948), .B(n15947), .ZN(
        P1_U2986) );
  XOR2_X1 U19039 ( .A(n15950), .B(n15949), .Z(n16061) );
  AOI22_X1 U19040 ( .A1(n20120), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n20162), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15954) );
  AOI22_X1 U19041 ( .A1(n15952), .A2(n20125), .B1(n15951), .B2(n15961), .ZN(
        n15953) );
  OAI211_X1 U19042 ( .C1(n16061), .C2(n19918), .A(n15954), .B(n15953), .ZN(
        P1_U2987) );
  MUX2_X1 U19043 ( .A(n15957), .B(n15956), .S(n15955), .Z(n15959) );
  XNOR2_X1 U19044 ( .A(n15959), .B(n15958), .ZN(n16081) );
  AOI22_X1 U19045 ( .A1(n20120), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        n20162), .B2(P1_REIP_REG_10__SCAN_IN), .ZN(n15964) );
  AOI22_X1 U19046 ( .A1(n15962), .A2(n20125), .B1(n15961), .B2(n15960), .ZN(
        n15963) );
  OAI211_X1 U19047 ( .C1(n19918), .C2(n16081), .A(n15964), .B(n15963), .ZN(
        P1_U2989) );
  AOI22_X1 U19048 ( .A1(n20120), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n20162), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15970) );
  NAND2_X1 U19049 ( .A1(n15966), .A2(n15965), .ZN(n15967) );
  XNOR2_X1 U19050 ( .A(n15968), .B(n15967), .ZN(n16091) );
  AOI22_X1 U19051 ( .A1(n16091), .A2(n12697), .B1(n20125), .B2(n19967), .ZN(
        n15969) );
  OAI211_X1 U19052 ( .C1(n20130), .C2(n19962), .A(n15970), .B(n15969), .ZN(
        P1_U2992) );
  AOI22_X1 U19053 ( .A1(n20120), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n20162), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15975) );
  XNOR2_X1 U19054 ( .A(n15971), .B(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15972) );
  XNOR2_X1 U19055 ( .A(n15973), .B(n15972), .ZN(n16095) );
  AOI22_X1 U19056 ( .A1(n16095), .A2(n12697), .B1(n20125), .B2(n19979), .ZN(
        n15974) );
  OAI211_X1 U19057 ( .C1(n20130), .C2(n19971), .A(n15975), .B(n15974), .ZN(
        P1_U2993) );
  AOI22_X1 U19058 ( .A1(n20120), .A2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .B1(
        n20162), .B2(P1_REIP_REG_5__SCAN_IN), .ZN(n15981) );
  OAI21_X1 U19059 ( .B1(n15978), .B2(n15977), .A(n15976), .ZN(n15979) );
  INV_X1 U19060 ( .A(n15979), .ZN(n16102) );
  AOI22_X1 U19061 ( .A1(n16102), .A2(n12697), .B1(n20125), .B2(n19993), .ZN(
        n15980) );
  OAI211_X1 U19062 ( .C1(n20130), .C2(n19986), .A(n15981), .B(n15980), .ZN(
        P1_U2994) );
  INV_X1 U19063 ( .A(n15982), .ZN(n15991) );
  AOI22_X1 U19064 ( .A1(n20162), .A2(P1_REIP_REG_23__SCAN_IN), .B1(n15984), 
        .B2(n15983), .ZN(n15989) );
  INV_X1 U19065 ( .A(n15985), .ZN(n15987) );
  AOI22_X1 U19066 ( .A1(n15987), .A2(n20160), .B1(n20157), .B2(n15986), .ZN(
        n15988) );
  OAI211_X1 U19067 ( .C1(n15991), .C2(n15990), .A(n15989), .B(n15988), .ZN(
        P1_U3008) );
  INV_X1 U19068 ( .A(n15992), .ZN(n15993) );
  AOI22_X1 U19069 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n15993), .B1(
        n20162), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n15998) );
  INV_X1 U19070 ( .A(n15994), .ZN(n15995) );
  AOI22_X1 U19071 ( .A1(n15996), .A2(n20160), .B1(n20157), .B2(n15995), .ZN(
        n15997) );
  OAI211_X1 U19072 ( .C1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n15999), .A(
        n15998), .B(n15997), .ZN(P1_U3012) );
  OAI21_X1 U19073 ( .B1(n16001), .B2(n16028), .A(n16000), .ZN(n16004) );
  AOI22_X1 U19074 ( .A1(n16004), .A2(n16003), .B1(n20157), .B2(n16002), .ZN(
        n16006) );
  NAND2_X1 U19075 ( .A1(n20162), .A2(P1_REIP_REG_17__SCAN_IN), .ZN(n16005) );
  OAI211_X1 U19076 ( .C1(n16007), .C2(n16082), .A(n16006), .B(n16005), .ZN(
        P1_U3014) );
  AOI21_X1 U19077 ( .B1(n16009), .B2(n20157), .A(n16008), .ZN(n16014) );
  OAI21_X1 U19078 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16010), .A(
        n16026), .ZN(n16017) );
  AOI22_X1 U19079 ( .A1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n16017), .B1(
        n20160), .B2(n16011), .ZN(n16013) );
  NOR2_X1 U19080 ( .A1(n16027), .A2(n16028), .ZN(n16016) );
  OAI221_X1 U19081 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(n12600), .C2(n13840), .A(
        n16016), .ZN(n16012) );
  NAND3_X1 U19082 ( .A1(n16014), .A2(n16013), .A3(n16012), .ZN(P1_U3015) );
  AOI22_X1 U19083 ( .A1(n16015), .A2(n20157), .B1(n20162), .B2(
        P1_REIP_REG_15__SCAN_IN), .ZN(n16019) );
  AOI22_X1 U19084 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n16017), .B1(
        n16016), .B2(n12600), .ZN(n16018) );
  OAI211_X1 U19085 ( .C1(n16020), .C2(n16082), .A(n16019), .B(n16018), .ZN(
        P1_U3016) );
  OAI22_X1 U19086 ( .A1(n16022), .A2(n20137), .B1(n16021), .B2(n20135), .ZN(
        n16023) );
  AOI21_X1 U19087 ( .B1(n20160), .B2(n16024), .A(n16023), .ZN(n16025) );
  OAI221_X1 U19088 ( .B1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n16028), 
        .C1(n16027), .C2(n16026), .A(n16025), .ZN(P1_U3017) );
  NAND2_X1 U19089 ( .A1(n16030), .A2(n16029), .ZN(n16039) );
  INV_X1 U19090 ( .A(n16039), .ZN(n16036) );
  NOR2_X1 U19091 ( .A1(n20135), .A2(n16031), .ZN(n16035) );
  OAI22_X1 U19092 ( .A1(n16033), .A2(n20137), .B1(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n16032), .ZN(n16034) );
  AOI211_X1 U19093 ( .C1(n16037), .C2(n16036), .A(n16035), .B(n16034), .ZN(
        n16046) );
  NOR2_X1 U19094 ( .A1(n16038), .A2(n20154), .ZN(n16044) );
  OAI211_X1 U19095 ( .C1(n16042), .C2(n16041), .A(n16040), .B(n16039), .ZN(
        n16043) );
  OAI21_X1 U19096 ( .B1(n16044), .B2(n16043), .A(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n16045) );
  OAI211_X1 U19097 ( .C1(n16047), .C2(n16082), .A(n16046), .B(n16045), .ZN(
        P1_U3018) );
  AOI22_X1 U19098 ( .A1(n16048), .A2(n20157), .B1(n20162), .B2(
        P1_REIP_REG_12__SCAN_IN), .ZN(n16060) );
  NAND3_X1 U19099 ( .A1(n16051), .A2(n16050), .A3(n16049), .ZN(n16068) );
  OAI21_X1 U19100 ( .B1(n16069), .B2(n16052), .A(n20134), .ZN(n16053) );
  OAI211_X1 U19101 ( .C1(n16057), .C2(n20154), .A(n16072), .B(n16053), .ZN(
        n16065) );
  INV_X1 U19102 ( .A(n16065), .ZN(n16054) );
  OAI21_X1 U19103 ( .B1(n16055), .B2(n16068), .A(n16054), .ZN(n16058) );
  NOR2_X1 U19104 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16099), .ZN(
        n16056) );
  AOI22_X1 U19105 ( .A1(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n16058), .B1(
        n16057), .B2(n16056), .ZN(n16059) );
  OAI211_X1 U19106 ( .C1(n16061), .C2(n16082), .A(n16060), .B(n16059), .ZN(
        P1_U3019) );
  INV_X1 U19107 ( .A(n20146), .ZN(n20139) );
  AOI21_X1 U19108 ( .B1(n16063), .B2(n20157), .A(n16062), .ZN(n16067) );
  AOI22_X1 U19109 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n16065), .B1(
        n20160), .B2(n16064), .ZN(n16066) );
  OAI211_X1 U19110 ( .C1(n20139), .C2(n16068), .A(n16067), .B(n16066), .ZN(
        P1_U3020) );
  AOI211_X1 U19111 ( .C1(n20134), .C2(n16069), .A(n16098), .B(n16074), .ZN(
        n16071) );
  AOI21_X1 U19112 ( .B1(n16072), .B2(n16071), .A(n16070), .ZN(n16085) );
  INV_X1 U19113 ( .A(n16073), .ZN(n16094) );
  OR2_X1 U19114 ( .A1(n16074), .A2(n16094), .ZN(n16089) );
  AOI221_X1 U19115 ( .B1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(n15958), .C2(n16075), .A(
        n16089), .ZN(n16079) );
  OAI22_X1 U19116 ( .A1(n16077), .A2(n20137), .B1(n16076), .B2(n20135), .ZN(
        n16078) );
  AOI211_X1 U19117 ( .C1(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .C2(n16085), .A(
        n16079), .B(n16078), .ZN(n16080) );
  OAI21_X1 U19118 ( .B1(n16082), .B2(n16081), .A(n16080), .ZN(P1_U3021) );
  INV_X1 U19119 ( .A(n16083), .ZN(n16084) );
  AOI21_X1 U19120 ( .B1(n19938), .B2(n20157), .A(n16084), .ZN(n16088) );
  AOI22_X1 U19121 ( .A1(n16086), .A2(n20160), .B1(
        P1_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n16085), .ZN(n16087) );
  OAI211_X1 U19122 ( .C1(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n16089), .A(
        n16088), .B(n16087), .ZN(P1_U3022) );
  AOI22_X1 U19123 ( .A1(n19961), .A2(n20157), .B1(n20162), .B2(
        P1_REIP_REG_7__SCAN_IN), .ZN(n16093) );
  AOI22_X1 U19124 ( .A1(n16091), .A2(n20160), .B1(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n16090), .ZN(n16092) );
  OAI211_X1 U19125 ( .C1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n16094), .A(
        n16093), .B(n16092), .ZN(P1_U3024) );
  AOI222_X1 U19126 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(n20162), .B1(n20157), 
        .B2(n19973), .C1(n20160), .C2(n16095), .ZN(n16096) );
  OAI221_X1 U19127 ( .B1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n16099), .C1(
        n16098), .C2(n16097), .A(n16096), .ZN(P1_U3025) );
  INV_X1 U19128 ( .A(n16100), .ZN(n16106) );
  AOI22_X1 U19129 ( .A1(n19988), .A2(n20157), .B1(n20162), .B2(
        P1_REIP_REG_5__SCAN_IN), .ZN(n16104) );
  AOI22_X1 U19130 ( .A1(n16102), .A2(n20160), .B1(n16101), .B2(n20146), .ZN(
        n16103) );
  OAI211_X1 U19131 ( .C1(n16106), .C2(n16105), .A(n16104), .B(n16103), .ZN(
        P1_U3026) );
  NAND4_X1 U19132 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20760), .A4(n20767), .ZN(n16107) );
  AND2_X1 U19133 ( .A1(n16108), .A2(n16107), .ZN(n20670) );
  AOI21_X1 U19134 ( .B1(n20670), .B2(n16110), .A(n16109), .ZN(n16112) );
  AOI211_X1 U19135 ( .C1(n20669), .C2(n16113), .A(n16112), .B(n16111), .ZN(
        P1_U3162) );
  OAI21_X1 U19136 ( .B1(n16115), .B2(n20379), .A(n16114), .ZN(P1_U3466) );
  NOR2_X1 U19137 ( .A1(n19116), .A2(n13666), .ZN(n18929) );
  INV_X1 U19138 ( .A(n18929), .ZN(n16130) );
  NAND2_X1 U19139 ( .A1(n19080), .A2(n16116), .ZN(n16217) );
  INV_X1 U19140 ( .A(n16117), .ZN(n16218) );
  NAND2_X1 U19141 ( .A1(n16217), .A2(n16218), .ZN(n16216) );
  NAND2_X1 U19142 ( .A1(n19080), .A2(n16216), .ZN(n16204) );
  NAND2_X1 U19143 ( .A1(n16205), .A2(n16204), .ZN(n16203) );
  NAND2_X1 U19144 ( .A1(n19080), .A2(n16203), .ZN(n16191) );
  INV_X1 U19145 ( .A(n16118), .ZN(n16192) );
  NAND2_X1 U19146 ( .A1(n16191), .A2(n16192), .ZN(n16190) );
  NAND2_X1 U19147 ( .A1(n19080), .A2(n16190), .ZN(n16181) );
  NAND2_X1 U19148 ( .A1(n16181), .A2(n16182), .ZN(n16180) );
  NAND2_X1 U19149 ( .A1(n19080), .A2(n16180), .ZN(n16172) );
  INV_X1 U19150 ( .A(n16119), .ZN(n16173) );
  NAND2_X1 U19151 ( .A1(n16172), .A2(n16173), .ZN(n16171) );
  NAND2_X1 U19152 ( .A1(n19080), .A2(n16171), .ZN(n16160) );
  NAND2_X1 U19153 ( .A1(n16160), .A2(n16161), .ZN(n16159) );
  NAND2_X1 U19154 ( .A1(n19080), .A2(n16159), .ZN(n16147) );
  INV_X1 U19155 ( .A(n16120), .ZN(n16148) );
  NAND2_X1 U19156 ( .A1(n16147), .A2(n16148), .ZN(n16146) );
  NAND2_X1 U19157 ( .A1(n19080), .A2(n16146), .ZN(n16139) );
  NAND2_X1 U19158 ( .A1(n16139), .A2(n16138), .ZN(n16137) );
  INV_X1 U19159 ( .A(n16121), .ZN(n16124) );
  OAI222_X1 U19160 ( .A1(n19110), .A2(n16125), .B1(n19086), .B2(n16124), .C1(
        n16123), .C2(n16122), .ZN(n16126) );
  AOI21_X1 U19161 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n19065), .A(
        n16126), .ZN(n16129) );
  AOI22_X1 U19162 ( .A1(n19099), .A2(n19122), .B1(n19112), .B2(n16127), .ZN(
        n16128) );
  OAI211_X1 U19163 ( .C1(n16130), .C2(n16137), .A(n16129), .B(n16128), .ZN(
        P2_U2824) );
  AOI22_X1 U19164 ( .A1(n19064), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n19070), .ZN(n16131) );
  INV_X1 U19165 ( .A(n16131), .ZN(n16135) );
  INV_X1 U19166 ( .A(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16132) );
  OAI22_X1 U19167 ( .A1(n16133), .A2(n19086), .B1(n19101), .B2(n16132), .ZN(
        n16134) );
  AOI211_X1 U19168 ( .C1(n16136), .C2(n19099), .A(n16135), .B(n16134), .ZN(
        n16141) );
  OAI211_X1 U19169 ( .C1(n16139), .C2(n16138), .A(n16137), .B(n19076), .ZN(
        n16140) );
  OAI211_X1 U19170 ( .C1(n19091), .C2(n16142), .A(n16141), .B(n16140), .ZN(
        P2_U2825) );
  AOI22_X1 U19171 ( .A1(P2_REIP_REG_29__SCAN_IN), .A2(n19070), .B1(
        P2_EBX_REG_29__SCAN_IN), .B2(n19064), .ZN(n16152) );
  AOI22_X1 U19172 ( .A1(n16143), .A2(n19107), .B1(
        P2_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n19065), .ZN(n16151) );
  AOI22_X1 U19173 ( .A1(n16145), .A2(n19112), .B1(n16144), .B2(n19099), .ZN(
        n16150) );
  OAI211_X1 U19174 ( .C1(n16148), .C2(n16147), .A(n19076), .B(n16146), .ZN(
        n16149) );
  NAND4_X1 U19175 ( .A1(n16152), .A2(n16151), .A3(n16150), .A4(n16149), .ZN(
        P2_U2826) );
  AOI22_X1 U19176 ( .A1(n19064), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n19070), .ZN(n16156) );
  INV_X1 U19177 ( .A(n16153), .ZN(n16154) );
  AOI22_X1 U19178 ( .A1(n16154), .A2(n19107), .B1(
        P2_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n19065), .ZN(n16155) );
  OAI211_X1 U19179 ( .C1(n16157), .C2(n19091), .A(n16156), .B(n16155), .ZN(
        n16158) );
  INV_X1 U19180 ( .A(n16158), .ZN(n16163) );
  OAI211_X1 U19181 ( .C1(n16161), .C2(n16160), .A(n19076), .B(n16159), .ZN(
        n16162) );
  OAI211_X1 U19182 ( .C1(n19085), .C2(n16164), .A(n16163), .B(n16162), .ZN(
        P2_U2827) );
  AOI22_X1 U19183 ( .A1(n19064), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_REIP_REG_27__SCAN_IN), .B2(n19070), .ZN(n16165) );
  INV_X1 U19184 ( .A(n16165), .ZN(n16169) );
  OAI22_X1 U19185 ( .A1(n16167), .A2(n19086), .B1(n19101), .B2(n16166), .ZN(
        n16168) );
  AOI211_X1 U19186 ( .C1(n16170), .C2(n19112), .A(n16169), .B(n16168), .ZN(
        n16175) );
  OAI211_X1 U19187 ( .C1(n16173), .C2(n16172), .A(n19076), .B(n16171), .ZN(
        n16174) );
  OAI211_X1 U19188 ( .C1(n19085), .C2(n16176), .A(n16175), .B(n16174), .ZN(
        P2_U2828) );
  AOI22_X1 U19189 ( .A1(P2_REIP_REG_26__SCAN_IN), .A2(n19070), .B1(
        P2_EBX_REG_26__SCAN_IN), .B2(n19064), .ZN(n16186) );
  AOI22_X1 U19190 ( .A1(n16177), .A2(n19107), .B1(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n19065), .ZN(n16185) );
  AOI22_X1 U19191 ( .A1(n16179), .A2(n19112), .B1(n16178), .B2(n19099), .ZN(
        n16184) );
  OAI211_X1 U19192 ( .C1(n16182), .C2(n16181), .A(n19076), .B(n16180), .ZN(
        n16183) );
  NAND4_X1 U19193 ( .A1(n16186), .A2(n16185), .A3(n16184), .A4(n16183), .ZN(
        P2_U2829) );
  AOI22_X1 U19194 ( .A1(P2_REIP_REG_25__SCAN_IN), .A2(n19070), .B1(
        P2_EBX_REG_25__SCAN_IN), .B2(n19064), .ZN(n16196) );
  AOI22_X1 U19195 ( .A1(n16187), .A2(n19107), .B1(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n19065), .ZN(n16195) );
  AOI22_X1 U19196 ( .A1(n16189), .A2(n19112), .B1(n16188), .B2(n19099), .ZN(
        n16194) );
  OAI211_X1 U19197 ( .C1(n16192), .C2(n16191), .A(n19076), .B(n16190), .ZN(
        n16193) );
  NAND4_X1 U19198 ( .A1(n16196), .A2(n16195), .A3(n16194), .A4(n16193), .ZN(
        P2_U2830) );
  AOI22_X1 U19199 ( .A1(P2_REIP_REG_24__SCAN_IN), .A2(n19070), .B1(
        P2_EBX_REG_24__SCAN_IN), .B2(n19064), .ZN(n16209) );
  INV_X1 U19200 ( .A(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n16197) );
  OAI22_X1 U19201 ( .A1(n16198), .A2(n19086), .B1(n19101), .B2(n16197), .ZN(
        n16199) );
  INV_X1 U19202 ( .A(n16199), .ZN(n16208) );
  INV_X1 U19203 ( .A(n16200), .ZN(n16202) );
  AOI22_X1 U19204 ( .A1(n16202), .A2(n19112), .B1(n16201), .B2(n19099), .ZN(
        n16207) );
  OAI211_X1 U19205 ( .C1(n16205), .C2(n16204), .A(n19076), .B(n16203), .ZN(
        n16206) );
  NAND4_X1 U19206 ( .A1(n16209), .A2(n16208), .A3(n16207), .A4(n16206), .ZN(
        P2_U2831) );
  AOI22_X1 U19207 ( .A1(n19064), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n19070), .ZN(n16210) );
  INV_X1 U19208 ( .A(n16210), .ZN(n16214) );
  OAI22_X1 U19209 ( .A1(n16212), .A2(n19086), .B1(n19101), .B2(n16211), .ZN(
        n16213) );
  AOI211_X1 U19210 ( .C1(n16215), .C2(n19112), .A(n16214), .B(n16213), .ZN(
        n16220) );
  OAI211_X1 U19211 ( .C1(n16218), .C2(n16217), .A(n19076), .B(n16216), .ZN(
        n16219) );
  OAI211_X1 U19212 ( .C1(n19085), .C2(n16221), .A(n16220), .B(n16219), .ZN(
        P2_U2832) );
  AOI22_X1 U19213 ( .A1(n16252), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19069), .ZN(n16227) );
  INV_X1 U19214 ( .A(n16222), .ZN(n16224) );
  AOI222_X1 U19215 ( .A1(n16225), .A2(n16282), .B1(n16281), .B2(n16224), .C1(
        n16284), .C2(n16223), .ZN(n16226) );
  OAI211_X1 U19216 ( .C1(n16257), .C2(n16228), .A(n16227), .B(n16226), .ZN(
        P2_U2992) );
  INV_X1 U19217 ( .A(n18982), .ZN(n16229) );
  AOI22_X1 U19218 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19069), .B1(n16279), 
        .B2(n16229), .ZN(n16235) );
  INV_X1 U19219 ( .A(n16230), .ZN(n18979) );
  INV_X1 U19220 ( .A(n16231), .ZN(n16232) );
  AOI222_X1 U19221 ( .A1(n16233), .A2(n16282), .B1(n16281), .B2(n18979), .C1(
        n16284), .C2(n16232), .ZN(n16234) );
  OAI211_X1 U19222 ( .C1(n16288), .C2(n16236), .A(n16235), .B(n16234), .ZN(
        P2_U3001) );
  AOI22_X1 U19223 ( .A1(n16252), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19069), .ZN(n16243) );
  NOR2_X1 U19224 ( .A1(n16237), .A2(n16259), .ZN(n16241) );
  NOR3_X1 U19225 ( .A1(n16239), .A2(n16238), .A3(n16260), .ZN(n16240) );
  AOI211_X1 U19226 ( .C1(n16281), .C2(n18993), .A(n16241), .B(n16240), .ZN(
        n16242) );
  OAI211_X1 U19227 ( .C1(n16257), .C2(n16244), .A(n16243), .B(n16242), .ZN(
        P2_U3002) );
  AOI22_X1 U19228 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19069), .B1(n16279), 
        .B2(n16245), .ZN(n16250) );
  OAI22_X1 U19229 ( .A1(n16247), .A2(n16260), .B1(n16246), .B2(n16259), .ZN(
        n16248) );
  AOI21_X1 U19230 ( .B1(n16281), .B2(n19002), .A(n16248), .ZN(n16249) );
  OAI211_X1 U19231 ( .C1(n16288), .C2(n16251), .A(n16250), .B(n16249), .ZN(
        P2_U3003) );
  AOI22_X1 U19232 ( .A1(n16252), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19069), .ZN(n16256) );
  AOI222_X1 U19233 ( .A1(n16254), .A2(n16282), .B1(n16281), .B2(n19016), .C1(
        n16284), .C2(n16253), .ZN(n16255) );
  OAI211_X1 U19234 ( .C1(n16257), .C2(n19014), .A(n16256), .B(n16255), .ZN(
        P2_U3004) );
  AOI22_X1 U19235 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n19069), .B1(n16279), 
        .B2(n19024), .ZN(n16264) );
  OAI22_X1 U19236 ( .A1(n16261), .A2(n16260), .B1(n16259), .B2(n16258), .ZN(
        n16262) );
  AOI21_X1 U19237 ( .B1(n16281), .B2(n19027), .A(n16262), .ZN(n16263) );
  OAI211_X1 U19238 ( .C1(n16288), .C2(n16265), .A(n16264), .B(n16263), .ZN(
        P2_U3005) );
  AOI22_X1 U19239 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19069), .B1(n16279), 
        .B2(n19036), .ZN(n16277) );
  INV_X1 U19240 ( .A(n16266), .ZN(n16268) );
  OAI21_X1 U19241 ( .B1(n16269), .B2(n16268), .A(n16267), .ZN(n16273) );
  NAND2_X1 U19242 ( .A1(n16271), .A2(n16270), .ZN(n16272) );
  XNOR2_X1 U19243 ( .A(n16273), .B(n16272), .ZN(n16297) );
  XOR2_X1 U19244 ( .A(n16275), .B(n16274), .Z(n16293) );
  AOI222_X1 U19245 ( .A1(n16297), .A2(n16282), .B1(n16281), .B2(n16295), .C1(
        n16284), .C2(n16293), .ZN(n16276) );
  OAI211_X1 U19246 ( .C1(n16288), .C2(n16278), .A(n16277), .B(n16276), .ZN(
        P2_U3006) );
  AOI22_X1 U19247 ( .A1(P2_REIP_REG_6__SCAN_IN), .A2(n19069), .B1(n16279), 
        .B2(n19058), .ZN(n16287) );
  INV_X1 U19248 ( .A(n16280), .ZN(n16285) );
  AOI222_X1 U19249 ( .A1(n16285), .A2(n16284), .B1(n16283), .B2(n16282), .C1(
        n16281), .C2(n19059), .ZN(n16286) );
  OAI211_X1 U19250 ( .C1(n16288), .C2(n19052), .A(n16287), .B(n16286), .ZN(
        P2_U3008) );
  INV_X1 U19251 ( .A(n16289), .ZN(n16292) );
  AOI21_X1 U19252 ( .B1(n16291), .B2(n16290), .A(n13044), .ZN(n19129) );
  AOI22_X1 U19253 ( .A1(n16292), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .B1(
        n16306), .B2(n19129), .ZN(n16303) );
  AOI222_X1 U19254 ( .A1(n16297), .A2(n16296), .B1(n16316), .B2(n16295), .C1(
        n16294), .C2(n16293), .ZN(n16302) );
  NAND2_X1 U19255 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19069), .ZN(n16301) );
  OAI211_X1 U19256 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16299), .B(n16298), .ZN(n16300) );
  NAND4_X1 U19257 ( .A1(n16303), .A2(n16302), .A3(n16301), .A4(n16300), .ZN(
        P2_U3038) );
  OR2_X1 U19258 ( .A1(n16305), .A2(n16304), .ZN(n16308) );
  NAND2_X1 U19259 ( .A1(n16306), .A2(n19166), .ZN(n16307) );
  AND2_X1 U19260 ( .A1(n16308), .A2(n16307), .ZN(n16318) );
  OAI22_X1 U19261 ( .A1(n16312), .A2(n16311), .B1(n16310), .B2(n16309), .ZN(
        n16313) );
  AOI211_X1 U19262 ( .C1(n16316), .C2(n16315), .A(n16314), .B(n16313), .ZN(
        n16317) );
  OAI211_X1 U19263 ( .C1(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n16319), .A(
        n16318), .B(n16317), .ZN(P2_U3046) );
  AND2_X1 U19264 ( .A1(n16321), .A2(n16320), .ZN(n19875) );
  INV_X1 U19265 ( .A(n16325), .ZN(n16322) );
  OAI21_X1 U19266 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19898), .A(n16322), 
        .ZN(n19753) );
  AOI221_X1 U19267 ( .B1(n19875), .B2(P2_STATE2_REG_0__SCAN_IN), .C1(n19753), 
        .C2(P2_STATE2_REG_0__SCAN_IN), .A(n16323), .ZN(n16329) );
  NAND2_X1 U19268 ( .A1(n16325), .A2(n16324), .ZN(n19756) );
  OAI211_X1 U19269 ( .C1(n16327), .C2(n16326), .A(n18853), .B(n19756), .ZN(
        n16328) );
  OAI211_X1 U19270 ( .C1(n16330), .C2(n18857), .A(n16329), .B(n16328), .ZN(
        P2_U3176) );
  INV_X1 U19271 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18794) );
  AOI22_X1 U19272 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n17769), .B1(
        n17587), .B2(n18794), .ZN(n16340) );
  NOR2_X1 U19273 ( .A1(n17769), .A2(n16332), .ZN(n16338) );
  AOI21_X1 U19274 ( .B1(n18794), .B2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A(
        n16335), .ZN(n16333) );
  INV_X1 U19275 ( .A(n16333), .ZN(n16334) );
  OAI22_X1 U19276 ( .A1(n16338), .A2(n16334), .B1(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n17587), .ZN(n16339) );
  OAI21_X1 U19277 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n16335), .A(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16336) );
  NAND2_X1 U19278 ( .A1(n16340), .A2(n16336), .ZN(n16337) );
  OAI22_X1 U19279 ( .A1(n16340), .A2(n16339), .B1(n16338), .B2(n16337), .ZN(
        n16396) );
  INV_X1 U19280 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16345) );
  NAND2_X1 U19281 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17818) );
  INV_X1 U19282 ( .A(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17820) );
  NAND2_X1 U19283 ( .A1(n17806), .A2(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n17716) );
  NAND2_X1 U19284 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17717) );
  INV_X1 U19285 ( .A(n17717), .ZN(n17758) );
  NAND3_X1 U19286 ( .A1(n17758), .A2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n16781) );
  NOR2_X1 U19287 ( .A1(n16781), .A2(n17720), .ZN(n16739) );
  NAND2_X1 U19288 ( .A1(n17757), .A2(n16739), .ZN(n17695) );
  NAND2_X1 U19289 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17697) );
  NAND2_X1 U19290 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n17648) );
  NAND2_X1 U19291 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17616) );
  NAND2_X1 U19292 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17599), .ZN(
        n17572) );
  NAND2_X1 U19293 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17573) );
  NAND2_X1 U19294 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17534) );
  NAND2_X1 U19295 ( .A1(n17521), .A2(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17492) );
  NAND2_X1 U19296 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17491) );
  NAND2_X1 U19297 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n16343), .ZN(
        n16368) );
  NAND2_X1 U19298 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n16354), .ZN(
        n16341) );
  INV_X1 U19299 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18766) );
  NOR2_X1 U19300 ( .A1(n18766), .A2(n9642), .ZN(n16389) );
  INV_X1 U19301 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17855) );
  NAND2_X1 U19302 ( .A1(n18779), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18696) );
  INV_X1 U19303 ( .A(n18696), .ZN(n17685) );
  OAI21_X1 U19304 ( .B1(n17855), .B2(n17598), .A(n18397), .ZN(n17490) );
  NAND2_X1 U19305 ( .A1(n16343), .A2(n17490), .ZN(n16358) );
  XNOR2_X1 U19306 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16346) );
  NOR2_X1 U19307 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17598), .ZN(
        n16367) );
  NOR2_X1 U19308 ( .A1(n17855), .A2(n17492), .ZN(n16544) );
  INV_X1 U19309 ( .A(n16544), .ZN(n16342) );
  NOR2_X1 U19310 ( .A1(n16342), .A2(n17491), .ZN(n16542) );
  NOR2_X1 U19311 ( .A1(n18397), .A2(n16343), .ZN(n16369) );
  INV_X1 U19312 ( .A(n16369), .ZN(n16344) );
  OAI211_X1 U19313 ( .C1(n16542), .C2(n18696), .A(n17859), .B(n16344), .ZN(
        n16371) );
  NOR2_X1 U19314 ( .A1(n16367), .A2(n16371), .ZN(n16356) );
  OAI22_X1 U19315 ( .A1(n16358), .A2(n16346), .B1(n16356), .B2(n16345), .ZN(
        n16347) );
  AOI211_X1 U19316 ( .C1(n17688), .C2(n9653), .A(n16389), .B(n16347), .ZN(
        n16351) );
  NOR2_X4 U19317 ( .A1(n18204), .A2(n16516), .ZN(n17848) );
  NAND2_X1 U19318 ( .A1(n16361), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16348) );
  XOR2_X1 U19319 ( .A(n18794), .B(n16348), .Z(n16393) );
  NAND2_X1 U19320 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16360), .ZN(
        n16349) );
  XOR2_X1 U19321 ( .A(n18794), .B(n16349), .Z(n16392) );
  AOI22_X1 U19322 ( .A1(n17848), .A2(n16393), .B1(n17725), .B2(n16392), .ZN(
        n16350) );
  OAI211_X1 U19323 ( .C1(n17727), .C2(n16396), .A(n16351), .B(n16350), .ZN(
        P3_U2799) );
  OAI22_X2 U19324 ( .A1(n18053), .A2(n17863), .B1(n17773), .B2(n18051), .ZN(
        n17732) );
  NOR2_X2 U19325 ( .A1(n16352), .A2(n17655), .ZN(n17565) );
  NAND2_X1 U19326 ( .A1(n16353), .A2(n17565), .ZN(n17519) );
  INV_X1 U19327 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16357) );
  XNOR2_X1 U19328 ( .A(n16357), .B(n16354), .ZN(n16565) );
  OAI221_X1 U19329 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16358), .C1(
        n16357), .C2(n16356), .A(n16355), .ZN(n16359) );
  AOI21_X1 U19330 ( .B1(n17688), .B2(n16565), .A(n16359), .ZN(n16365) );
  OAI22_X1 U19331 ( .A1(n16361), .A2(n17863), .B1(n16360), .B2(n17773), .ZN(
        n16363) );
  AOI22_X1 U19332 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16363), .B1(
        n17770), .B2(n16362), .ZN(n16364) );
  OAI211_X1 U19333 ( .C1(n16366), .C2(n17519), .A(n16365), .B(n16364), .ZN(
        P3_U2800) );
  NOR2_X1 U19334 ( .A1(n16367), .A2(n17688), .ZN(n16374) );
  OAI21_X1 U19335 ( .B1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n16542), .A(
        n16368), .ZN(n16580) );
  AOI22_X1 U19336 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n16371), .B1(
        n16370), .B2(n16369), .ZN(n16373) );
  OAI211_X1 U19337 ( .C1(n16374), .C2(n16580), .A(n16373), .B(n16372), .ZN(
        n16375) );
  AOI21_X1 U19338 ( .B1(n17770), .B2(n16376), .A(n16375), .ZN(n16382) );
  NOR2_X1 U19339 ( .A1(n16377), .A2(n17870), .ZN(n16402) );
  OAI211_X1 U19340 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16402), .A(
        n17725), .B(n16378), .ZN(n16381) );
  OAI211_X1 U19341 ( .C1(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n16403), .A(
        n17848), .B(n16379), .ZN(n16380) );
  NAND3_X1 U19342 ( .A1(n16382), .A2(n16381), .A3(n16380), .ZN(P3_U2801) );
  INV_X1 U19343 ( .A(n18169), .ZN(n16384) );
  OAI21_X1 U19344 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n16384), .A(
        n16383), .ZN(n16390) );
  NAND2_X1 U19345 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n18794), .ZN(
        n16386) );
  NOR4_X1 U19346 ( .A1(n16387), .A2(n16386), .A3(n18166), .A4(n16385), .ZN(
        n16388) );
  AOI211_X1 U19347 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16390), .A(
        n16389), .B(n16388), .ZN(n16395) );
  AOI22_X1 U19348 ( .A1(n16393), .A2(n18179), .B1(n16392), .B2(n16391), .ZN(
        n16394) );
  OAI211_X1 U19349 ( .C1(n16396), .C2(n18065), .A(n16395), .B(n16394), .ZN(
        P3_U2831) );
  NAND4_X1 U19350 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17769), .A3(
        n16397), .A4(n16408), .ZN(n16420) );
  NOR2_X1 U19351 ( .A1(n16398), .A2(n18166), .ZN(n18164) );
  INV_X1 U19352 ( .A(n18164), .ZN(n18183) );
  INV_X1 U19353 ( .A(n16398), .ZN(n18627) );
  INV_X1 U19354 ( .A(n17511), .ZN(n16417) );
  AOI22_X1 U19355 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17769), .B1(
        n17587), .B2(n16408), .ZN(n17504) );
  NAND2_X1 U19356 ( .A1(n17505), .A2(n17504), .ZN(n17503) );
  NAND4_X1 U19357 ( .A1(n18627), .A2(n16401), .A3(n16400), .A4(n17503), .ZN(
        n16407) );
  OAI22_X1 U19358 ( .A1(n16403), .A2(n18630), .B1(n16402), .B2(n18031), .ZN(
        n16404) );
  NOR3_X1 U19359 ( .A1(n18168), .A2(n16405), .A3(n16404), .ZN(n16406) );
  NAND2_X1 U19360 ( .A1(n16407), .A2(n16406), .ZN(n16416) );
  NOR2_X1 U19361 ( .A1(n18174), .A2(n16408), .ZN(n16415) );
  NOR2_X1 U19362 ( .A1(n17993), .A2(n17977), .ZN(n16409) );
  OAI22_X1 U19363 ( .A1(n18053), .A2(n18630), .B1(n18051), .B2(n18031), .ZN(
        n17970) );
  AOI21_X1 U19364 ( .B1(n18636), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n18655), .ZN(n17968) );
  INV_X1 U19365 ( .A(n17968), .ZN(n18154) );
  AOI22_X1 U19366 ( .A1(n16409), .A2(n17970), .B1(n17867), .B2(n18154), .ZN(
        n16410) );
  OAI21_X1 U19367 ( .B1(n18661), .B2(n17973), .A(n16410), .ZN(n17923) );
  NAND2_X1 U19368 ( .A1(n16411), .A2(n17923), .ZN(n17917) );
  NOR2_X1 U19369 ( .A1(n18166), .A2(n17917), .ZN(n17913) );
  INV_X1 U19370 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17518) );
  NOR3_X1 U19371 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17518), .A3(
        n17865), .ZN(n17501) );
  INV_X1 U19372 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18762) );
  NOR2_X1 U19373 ( .A1(n9642), .A2(n18762), .ZN(n17500) );
  OAI211_X1 U19374 ( .C1(n16420), .C2(n18183), .A(n16419), .B(n16418), .ZN(
        P3_U2834) );
  NOR3_X1 U19375 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16422) );
  NOR4_X1 U19376 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16421) );
  NAND4_X1 U19377 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16422), .A3(n16421), .A4(
        U215), .ZN(U213) );
  INV_X1 U19378 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19171) );
  INV_X2 U19379 ( .A(U214), .ZN(n16467) );
  NOR2_X1 U19380 ( .A1(n16467), .A2(n16423), .ZN(n16470) );
  INV_X1 U19381 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16505) );
  OAI222_X1 U19382 ( .A1(U212), .A2(n19171), .B1(n16469), .B2(n16424), .C1(
        U214), .C2(n16505), .ZN(U216) );
  AOI222_X1 U19383 ( .A1(n16466), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(n16470), 
        .B2(BUF1_REG_30__SCAN_IN), .C1(n16467), .C2(P1_DATAO_REG_30__SCAN_IN), 
        .ZN(n16425) );
  INV_X1 U19384 ( .A(n16425), .ZN(U217) );
  INV_X1 U19385 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n16427) );
  AOI22_X1 U19386 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16467), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16466), .ZN(n16426) );
  OAI21_X1 U19387 ( .B1(n16427), .B2(n16469), .A(n16426), .ZN(U218) );
  INV_X1 U19388 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16429) );
  AOI22_X1 U19389 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16467), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16466), .ZN(n16428) );
  OAI21_X1 U19390 ( .B1(n16429), .B2(n16469), .A(n16428), .ZN(U219) );
  INV_X1 U19391 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16431) );
  AOI22_X1 U19392 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16467), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16466), .ZN(n16430) );
  OAI21_X1 U19393 ( .B1(n16431), .B2(n16469), .A(n16430), .ZN(U220) );
  INV_X1 U19394 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16433) );
  AOI22_X1 U19395 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16467), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16466), .ZN(n16432) );
  OAI21_X1 U19396 ( .B1(n16433), .B2(n16469), .A(n16432), .ZN(U221) );
  INV_X1 U19397 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n16435) );
  AOI22_X1 U19398 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16467), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16466), .ZN(n16434) );
  OAI21_X1 U19399 ( .B1(n16435), .B2(n16469), .A(n16434), .ZN(U222) );
  INV_X1 U19400 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16437) );
  AOI22_X1 U19401 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16467), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16466), .ZN(n16436) );
  OAI21_X1 U19402 ( .B1(n16437), .B2(n16469), .A(n16436), .ZN(U223) );
  AOI22_X1 U19403 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16467), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16466), .ZN(n16438) );
  OAI21_X1 U19404 ( .B1(n14925), .B2(n16469), .A(n16438), .ZN(U224) );
  INV_X1 U19405 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n19245) );
  AOI22_X1 U19406 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16467), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16466), .ZN(n16439) );
  OAI21_X1 U19407 ( .B1(n19245), .B2(n16469), .A(n16439), .ZN(U225) );
  INV_X1 U19408 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n19238) );
  AOI22_X1 U19409 ( .A1(P1_DATAO_REG_21__SCAN_IN), .A2(n16467), .B1(
        P2_DATAO_REG_21__SCAN_IN), .B2(n16466), .ZN(n16440) );
  OAI21_X1 U19410 ( .B1(n19238), .B2(n16469), .A(n16440), .ZN(U226) );
  INV_X1 U19411 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16442) );
  AOI22_X1 U19412 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16467), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16466), .ZN(n16441) );
  OAI21_X1 U19413 ( .B1(n16442), .B2(n16469), .A(n16441), .ZN(U227) );
  INV_X1 U19414 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n16444) );
  AOI22_X1 U19415 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16467), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16466), .ZN(n16443) );
  OAI21_X1 U19416 ( .B1(n16444), .B2(n16469), .A(n16443), .ZN(U228) );
  AOI22_X1 U19417 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16467), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16466), .ZN(n16445) );
  OAI21_X1 U19418 ( .B1(n16446), .B2(n16469), .A(n16445), .ZN(U229) );
  INV_X1 U19419 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n19222) );
  AOI22_X1 U19420 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16467), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16466), .ZN(n16447) );
  OAI21_X1 U19421 ( .B1(n19222), .B2(n16469), .A(n16447), .ZN(U230) );
  AOI22_X1 U19422 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16467), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16466), .ZN(n16448) );
  OAI21_X1 U19423 ( .B1(n14993), .B2(n16469), .A(n16448), .ZN(U231) );
  AOI22_X1 U19424 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16467), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16466), .ZN(n16449) );
  OAI21_X1 U19425 ( .B1(n12982), .B2(n16469), .A(n16449), .ZN(U232) );
  INV_X1 U19426 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n20949) );
  AOI22_X1 U19427 ( .A1(BUF1_REG_14__SCAN_IN), .A2(n16470), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(n16467), .ZN(n16450) );
  OAI21_X1 U19428 ( .B1(n20949), .B2(U212), .A(n16450), .ZN(U233) );
  INV_X1 U19429 ( .A(P2_DATAO_REG_13__SCAN_IN), .ZN(n16486) );
  AOI22_X1 U19430 ( .A1(BUF1_REG_13__SCAN_IN), .A2(n16470), .B1(
        P1_DATAO_REG_13__SCAN_IN), .B2(n16467), .ZN(n16451) );
  OAI21_X1 U19431 ( .B1(n16486), .B2(U212), .A(n16451), .ZN(U234) );
  INV_X1 U19432 ( .A(P2_DATAO_REG_12__SCAN_IN), .ZN(n16485) );
  AOI22_X1 U19433 ( .A1(BUF1_REG_12__SCAN_IN), .A2(n16470), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n16467), .ZN(n16452) );
  OAI21_X1 U19434 ( .B1(n16485), .B2(U212), .A(n16452), .ZN(U235) );
  INV_X1 U19435 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n16484) );
  AOI22_X1 U19436 ( .A1(BUF1_REG_11__SCAN_IN), .A2(n16470), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n16467), .ZN(n16453) );
  OAI21_X1 U19437 ( .B1(n16484), .B2(U212), .A(n16453), .ZN(U236) );
  INV_X1 U19438 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n16455) );
  AOI22_X1 U19439 ( .A1(BUF1_REG_10__SCAN_IN), .A2(n16470), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n16467), .ZN(n16454) );
  OAI21_X1 U19440 ( .B1(n16455), .B2(U212), .A(n16454), .ZN(U237) );
  AOI22_X1 U19441 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16467), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16466), .ZN(n16456) );
  OAI21_X1 U19442 ( .B1(n16457), .B2(n16469), .A(n16456), .ZN(U238) );
  AOI22_X1 U19443 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16467), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16466), .ZN(n16458) );
  OAI21_X1 U19444 ( .B1(n16459), .B2(n16469), .A(n16458), .ZN(U239) );
  INV_X1 U19445 ( .A(P2_DATAO_REG_7__SCAN_IN), .ZN(n16479) );
  AOI22_X1 U19446 ( .A1(BUF1_REG_7__SCAN_IN), .A2(n16470), .B1(
        P1_DATAO_REG_7__SCAN_IN), .B2(n16467), .ZN(n16460) );
  OAI21_X1 U19447 ( .B1(n16479), .B2(U212), .A(n16460), .ZN(U240) );
  INV_X1 U19448 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n16478) );
  AOI22_X1 U19449 ( .A1(BUF1_REG_6__SCAN_IN), .A2(n16470), .B1(
        P1_DATAO_REG_6__SCAN_IN), .B2(n16467), .ZN(n16461) );
  OAI21_X1 U19450 ( .B1(n16478), .B2(U212), .A(n16461), .ZN(U241) );
  INV_X1 U19451 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n20793) );
  AOI22_X1 U19452 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16467), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16466), .ZN(n16462) );
  OAI21_X1 U19453 ( .B1(n20793), .B2(n16469), .A(n16462), .ZN(U242) );
  INV_X1 U19454 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n20955) );
  AOI22_X1 U19455 ( .A1(BUF1_REG_4__SCAN_IN), .A2(n16470), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16466), .ZN(n16463) );
  OAI21_X1 U19456 ( .B1(n20955), .B2(U214), .A(n16463), .ZN(U243) );
  INV_X1 U19457 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n16475) );
  AOI22_X1 U19458 ( .A1(BUF1_REG_3__SCAN_IN), .A2(n16470), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n16467), .ZN(n16464) );
  OAI21_X1 U19459 ( .B1(n16475), .B2(U212), .A(n16464), .ZN(U244) );
  INV_X1 U19460 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n20815) );
  AOI22_X1 U19461 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16467), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16466), .ZN(n16465) );
  OAI21_X1 U19462 ( .B1(n20815), .B2(n16469), .A(n16465), .ZN(U245) );
  INV_X1 U19463 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n20946) );
  AOI22_X1 U19464 ( .A1(P1_DATAO_REG_1__SCAN_IN), .A2(n16467), .B1(
        P2_DATAO_REG_1__SCAN_IN), .B2(n16466), .ZN(n16468) );
  OAI21_X1 U19465 ( .B1(n20946), .B2(n16469), .A(n16468), .ZN(U246) );
  INV_X1 U19466 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n16472) );
  AOI22_X1 U19467 ( .A1(BUF1_REG_0__SCAN_IN), .A2(n16470), .B1(
        P1_DATAO_REG_0__SCAN_IN), .B2(n16467), .ZN(n16471) );
  OAI21_X1 U19468 ( .B1(n16472), .B2(U212), .A(n16471), .ZN(U247) );
  INV_X1 U19469 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18198) );
  AOI22_X1 U19470 ( .A1(n16503), .A2(n16472), .B1(n18198), .B2(U215), .ZN(U251) );
  OAI22_X1 U19471 ( .A1(U215), .A2(P2_DATAO_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n16503), .ZN(n16473) );
  INV_X1 U19472 ( .A(n16473), .ZN(U252) );
  OAI22_X1 U19473 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16503), .ZN(n16474) );
  INV_X1 U19474 ( .A(n16474), .ZN(U253) );
  INV_X1 U19475 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18214) );
  AOI22_X1 U19476 ( .A1(n16503), .A2(n16475), .B1(n18214), .B2(U215), .ZN(U254) );
  OAI22_X1 U19477 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16503), .ZN(n16476) );
  INV_X1 U19478 ( .A(n16476), .ZN(U255) );
  OAI22_X1 U19479 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16503), .ZN(n16477) );
  INV_X1 U19480 ( .A(n16477), .ZN(U256) );
  INV_X1 U19481 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18230) );
  AOI22_X1 U19482 ( .A1(n16503), .A2(n16478), .B1(n18230), .B2(U215), .ZN(U257) );
  INV_X1 U19483 ( .A(BUF2_REG_7__SCAN_IN), .ZN(n18235) );
  AOI22_X1 U19484 ( .A1(n16503), .A2(n16479), .B1(n18235), .B2(U215), .ZN(U258) );
  INV_X1 U19485 ( .A(P2_DATAO_REG_8__SCAN_IN), .ZN(n16481) );
  INV_X1 U19486 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n16480) );
  AOI22_X1 U19487 ( .A1(n16503), .A2(n16481), .B1(n16480), .B2(U215), .ZN(U259) );
  OAI22_X1 U19488 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16503), .ZN(n16482) );
  INV_X1 U19489 ( .A(n16482), .ZN(U260) );
  OAI22_X1 U19490 ( .A1(U215), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(
        BUF2_REG_10__SCAN_IN), .B2(n16503), .ZN(n16483) );
  INV_X1 U19491 ( .A(n16483), .ZN(U261) );
  INV_X1 U19492 ( .A(BUF2_REG_11__SCAN_IN), .ZN(n17334) );
  AOI22_X1 U19493 ( .A1(n16497), .A2(n16484), .B1(n17334), .B2(U215), .ZN(U262) );
  INV_X1 U19494 ( .A(BUF2_REG_12__SCAN_IN), .ZN(n17330) );
  AOI22_X1 U19495 ( .A1(n16503), .A2(n16485), .B1(n17330), .B2(U215), .ZN(U263) );
  INV_X1 U19496 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n17325) );
  AOI22_X1 U19497 ( .A1(n16497), .A2(n16486), .B1(n17325), .B2(U215), .ZN(U264) );
  OAI22_X1 U19498 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16503), .ZN(n16487) );
  INV_X1 U19499 ( .A(n16487), .ZN(U265) );
  OAI22_X1 U19500 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16503), .ZN(n16488) );
  INV_X1 U19501 ( .A(n16488), .ZN(U266) );
  INV_X1 U19502 ( .A(P2_DATAO_REG_16__SCAN_IN), .ZN(n20936) );
  AOI22_X1 U19503 ( .A1(n16497), .A2(n20936), .B1(n14995), .B2(U215), .ZN(U267) );
  OAI22_X1 U19504 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16503), .ZN(n16489) );
  INV_X1 U19505 ( .A(n16489), .ZN(U268) );
  OAI22_X1 U19506 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16497), .ZN(n16490) );
  INV_X1 U19507 ( .A(n16490), .ZN(U269) );
  OAI22_X1 U19508 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16497), .ZN(n16491) );
  INV_X1 U19509 ( .A(n16491), .ZN(U270) );
  OAI22_X1 U19510 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16497), .ZN(n16492) );
  INV_X1 U19511 ( .A(n16492), .ZN(U271) );
  OAI22_X1 U19512 ( .A1(U215), .A2(P2_DATAO_REG_21__SCAN_IN), .B1(
        BUF2_REG_21__SCAN_IN), .B2(n16497), .ZN(n16493) );
  INV_X1 U19513 ( .A(n16493), .ZN(U272) );
  OAI22_X1 U19514 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16497), .ZN(n16494) );
  INV_X1 U19515 ( .A(n16494), .ZN(U273) );
  OAI22_X1 U19516 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16497), .ZN(n16495) );
  INV_X1 U19517 ( .A(n16495), .ZN(U274) );
  OAI22_X1 U19518 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16503), .ZN(n16496) );
  INV_X1 U19519 ( .A(n16496), .ZN(U275) );
  OAI22_X1 U19520 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16497), .ZN(n16498) );
  INV_X1 U19521 ( .A(n16498), .ZN(U276) );
  OAI22_X1 U19522 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16503), .ZN(n16499) );
  INV_X1 U19523 ( .A(n16499), .ZN(U277) );
  OAI22_X1 U19524 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16503), .ZN(n16500) );
  INV_X1 U19525 ( .A(n16500), .ZN(U278) );
  OAI22_X1 U19526 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16503), .ZN(n16501) );
  INV_X1 U19527 ( .A(n16501), .ZN(U279) );
  OAI22_X1 U19528 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16503), .ZN(n16502) );
  INV_X1 U19529 ( .A(n16502), .ZN(U280) );
  INV_X1 U19530 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n19175) );
  INV_X1 U19531 ( .A(BUF2_REG_30__SCAN_IN), .ZN(n18229) );
  AOI22_X1 U19532 ( .A1(n16503), .A2(n19175), .B1(n18229), .B2(U215), .ZN(U281) );
  INV_X1 U19533 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n18237) );
  AOI22_X1 U19534 ( .A1(n16503), .A2(n19171), .B1(n18237), .B2(U215), .ZN(U282) );
  INV_X1 U19535 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16504) );
  AOI222_X1 U19536 ( .A1(n16505), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n19171), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16504), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16506) );
  INV_X2 U19537 ( .A(n16508), .ZN(n16507) );
  INV_X1 U19538 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18732) );
  INV_X1 U19539 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19794) );
  AOI22_X1 U19540 ( .A1(n16507), .A2(n18732), .B1(n19794), .B2(n16508), .ZN(
        U347) );
  INV_X1 U19541 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n18730) );
  INV_X1 U19542 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19792) );
  AOI22_X1 U19543 ( .A1(n16507), .A2(n18730), .B1(n19792), .B2(n16508), .ZN(
        U348) );
  INV_X1 U19544 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18727) );
  INV_X1 U19545 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19790) );
  AOI22_X1 U19546 ( .A1(n16507), .A2(n18727), .B1(n19790), .B2(n16508), .ZN(
        U349) );
  INV_X1 U19547 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18726) );
  INV_X1 U19548 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19788) );
  AOI22_X1 U19549 ( .A1(n16507), .A2(n18726), .B1(n19788), .B2(n16508), .ZN(
        U350) );
  INV_X1 U19550 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18724) );
  INV_X1 U19551 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20951) );
  AOI22_X1 U19552 ( .A1(n16507), .A2(n18724), .B1(n20951), .B2(n16508), .ZN(
        U351) );
  INV_X1 U19553 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18721) );
  INV_X1 U19554 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19785) );
  AOI22_X1 U19555 ( .A1(n16507), .A2(n18721), .B1(n19785), .B2(n16508), .ZN(
        U352) );
  INV_X1 U19556 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18720) );
  INV_X1 U19557 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n19784) );
  AOI22_X1 U19558 ( .A1(n16507), .A2(n18720), .B1(n19784), .B2(n16508), .ZN(
        U353) );
  INV_X1 U19559 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18718) );
  AOI22_X1 U19560 ( .A1(n16507), .A2(n18718), .B1(n19782), .B2(n16508), .ZN(
        U354) );
  INV_X1 U19561 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18767) );
  INV_X1 U19562 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19834) );
  AOI22_X1 U19563 ( .A1(n16507), .A2(n18767), .B1(n19834), .B2(n16508), .ZN(
        U355) );
  INV_X1 U19564 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18764) );
  INV_X1 U19565 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19830) );
  AOI22_X1 U19566 ( .A1(n16507), .A2(n18764), .B1(n19830), .B2(n16508), .ZN(
        U356) );
  INV_X1 U19567 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18761) );
  INV_X1 U19568 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19829) );
  AOI22_X1 U19569 ( .A1(n16507), .A2(n18761), .B1(n19829), .B2(n16508), .ZN(
        U357) );
  INV_X1 U19570 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18760) );
  INV_X1 U19571 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19826) );
  AOI22_X1 U19572 ( .A1(n16507), .A2(n18760), .B1(n19826), .B2(n16508), .ZN(
        U358) );
  INV_X1 U19573 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n20795) );
  INV_X1 U19574 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19825) );
  AOI22_X1 U19575 ( .A1(n16507), .A2(n20795), .B1(n19825), .B2(n16508), .ZN(
        U359) );
  INV_X1 U19576 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18757) );
  INV_X1 U19577 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19823) );
  AOI22_X1 U19578 ( .A1(n16507), .A2(n18757), .B1(n19823), .B2(n16508), .ZN(
        U360) );
  INV_X1 U19579 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n20938) );
  INV_X1 U19580 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19821) );
  AOI22_X1 U19581 ( .A1(n16507), .A2(n20938), .B1(n19821), .B2(n16508), .ZN(
        U361) );
  INV_X1 U19582 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18753) );
  INV_X1 U19583 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19819) );
  AOI22_X1 U19584 ( .A1(n16507), .A2(n18753), .B1(n19819), .B2(n16508), .ZN(
        U362) );
  INV_X1 U19585 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18752) );
  INV_X1 U19586 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19817) );
  AOI22_X1 U19587 ( .A1(n16507), .A2(n18752), .B1(n19817), .B2(n16508), .ZN(
        U363) );
  INV_X1 U19588 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18749) );
  INV_X1 U19589 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19815) );
  AOI22_X1 U19590 ( .A1(n16507), .A2(n18749), .B1(n19815), .B2(n16508), .ZN(
        U364) );
  INV_X1 U19591 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18716) );
  INV_X1 U19592 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19780) );
  AOI22_X1 U19593 ( .A1(n16507), .A2(n18716), .B1(n19780), .B2(n16508), .ZN(
        U365) );
  INV_X1 U19594 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18748) );
  INV_X1 U19595 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19813) );
  AOI22_X1 U19596 ( .A1(n16507), .A2(n18748), .B1(n19813), .B2(n16508), .ZN(
        U366) );
  INV_X1 U19597 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18745) );
  INV_X1 U19598 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19811) );
  AOI22_X1 U19599 ( .A1(n16507), .A2(n18745), .B1(n19811), .B2(n16508), .ZN(
        U367) );
  INV_X1 U19600 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18744) );
  INV_X1 U19601 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19809) );
  AOI22_X1 U19602 ( .A1(n16507), .A2(n18744), .B1(n19809), .B2(n16508), .ZN(
        U368) );
  INV_X1 U19603 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18741) );
  INV_X1 U19604 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19807) );
  AOI22_X1 U19605 ( .A1(n16507), .A2(n18741), .B1(n19807), .B2(n16508), .ZN(
        U369) );
  INV_X1 U19606 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18740) );
  INV_X1 U19607 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19805) );
  AOI22_X1 U19608 ( .A1(n16507), .A2(n18740), .B1(n19805), .B2(n16508), .ZN(
        U370) );
  INV_X1 U19609 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18738) );
  INV_X1 U19610 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19804) );
  AOI22_X1 U19611 ( .A1(n16507), .A2(n18738), .B1(n19804), .B2(n16508), .ZN(
        U371) );
  INV_X1 U19612 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n20775) );
  INV_X1 U19613 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19802) );
  AOI22_X1 U19614 ( .A1(n16507), .A2(n20775), .B1(n19802), .B2(n16508), .ZN(
        U372) );
  INV_X1 U19615 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18737) );
  INV_X1 U19616 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19800) );
  AOI22_X1 U19617 ( .A1(n16507), .A2(n18737), .B1(n19800), .B2(n16508), .ZN(
        U373) );
  INV_X1 U19618 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18735) );
  INV_X1 U19619 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19798) );
  AOI22_X1 U19620 ( .A1(n16507), .A2(n18735), .B1(n19798), .B2(n16508), .ZN(
        U374) );
  INV_X1 U19621 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18734) );
  INV_X1 U19622 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n19796) );
  AOI22_X1 U19623 ( .A1(n16507), .A2(n18734), .B1(n19796), .B2(n16508), .ZN(
        U375) );
  INV_X1 U19624 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18713) );
  INV_X1 U19625 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19778) );
  AOI22_X1 U19626 ( .A1(n16507), .A2(n18713), .B1(n19778), .B2(n16508), .ZN(
        U376) );
  INV_X1 U19627 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18712) );
  NAND2_X1 U19628 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18712), .ZN(n16509) );
  AOI22_X1 U19629 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n16509), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18710), .ZN(n18778) );
  AOI21_X1 U19630 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18778), .ZN(n16510) );
  INV_X1 U19631 ( .A(n16510), .ZN(P3_U2633) );
  INV_X1 U19632 ( .A(n18688), .ZN(n16537) );
  OAI21_X1 U19633 ( .B1(n16515), .B2(n17385), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16511) );
  OAI21_X1 U19634 ( .B1(n16512), .B2(n16537), .A(n16511), .ZN(P3_U2634) );
  AOI21_X1 U19635 ( .B1(n18710), .B2(n18712), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16513) );
  AOI22_X1 U19636 ( .A1(n20776), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16513), 
        .B2(n18842), .ZN(P3_U2635) );
  OAI21_X1 U19637 ( .B1(n18697), .B2(BS16), .A(n18778), .ZN(n18776) );
  OAI21_X1 U19638 ( .B1(n18778), .B2(n18833), .A(n18776), .ZN(P3_U2636) );
  NOR3_X1 U19639 ( .A1(n16515), .A2(n18626), .A3(n16514), .ZN(n18633) );
  NOR2_X1 U19640 ( .A1(n18633), .A2(n18675), .ZN(n18824) );
  OAI21_X1 U19641 ( .B1(n18824), .B2(n16517), .A(n16516), .ZN(P3_U2637) );
  NOR4_X1 U19642 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_21__SCAN_IN), .A3(P3_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_23__SCAN_IN), .ZN(n16521) );
  NOR4_X1 U19643 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_17__SCAN_IN), .A3(P3_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_19__SCAN_IN), .ZN(n16520) );
  NOR4_X1 U19644 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16519) );
  NOR4_X1 U19645 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_25__SCAN_IN), .A3(P3_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16518) );
  NAND4_X1 U19646 ( .A1(n16521), .A2(n16520), .A3(n16519), .A4(n16518), .ZN(
        n16527) );
  NOR4_X1 U19647 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16525) );
  AOI211_X1 U19648 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_7__SCAN_IN), .B(
        P3_DATAWIDTH_REG_2__SCAN_IN), .ZN(n16524) );
  NOR4_X1 U19649 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_13__SCAN_IN), .A3(P3_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_15__SCAN_IN), .ZN(n16523) );
  NOR4_X1 U19650 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_9__SCAN_IN), .A3(P3_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_11__SCAN_IN), .ZN(n16522) );
  NAND4_X1 U19651 ( .A1(n16525), .A2(n16524), .A3(n16523), .A4(n16522), .ZN(
        n16526) );
  NOR2_X1 U19652 ( .A1(n16527), .A2(n16526), .ZN(n18822) );
  INV_X1 U19653 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16529) );
  NOR3_X1 U19654 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16530) );
  OAI21_X1 U19655 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16530), .A(n18822), .ZN(
        n16528) );
  OAI21_X1 U19656 ( .B1(n18822), .B2(n16529), .A(n16528), .ZN(P3_U2638) );
  INV_X1 U19657 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16532) );
  NOR2_X1 U19658 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18817) );
  OAI21_X1 U19659 ( .B1(n16530), .B2(n18817), .A(n18822), .ZN(n16531) );
  OAI21_X1 U19660 ( .B1(n18822), .B2(n16532), .A(n16531), .ZN(P3_U2639) );
  INV_X1 U19661 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18755) );
  AOI211_X1 U19662 ( .C1(n18834), .C2(n18832), .A(n18829), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n18677) );
  INV_X1 U19663 ( .A(n16533), .ZN(n18623) );
  INV_X1 U19664 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n20954) );
  INV_X1 U19665 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18722) );
  NAND4_X1 U19666 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(P3_REIP_REG_3__SCAN_IN), 
        .A3(P3_REIP_REG_1__SCAN_IN), .A4(P3_REIP_REG_2__SCAN_IN), .ZN(n16850)
         );
  NOR2_X1 U19667 ( .A1(n18722), .A2(n16850), .ZN(n16833) );
  INV_X1 U19668 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18728) );
  NAND2_X1 U19669 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .ZN(n16814) );
  NOR2_X1 U19670 ( .A1(n18728), .A2(n16814), .ZN(n16794) );
  INV_X1 U19671 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18731) );
  INV_X1 U19672 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18729) );
  NOR2_X1 U19673 ( .A1(n18731), .A2(n18729), .ZN(n16795) );
  NAND4_X1 U19674 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16833), .A3(n16794), 
        .A4(n16795), .ZN(n16773) );
  NOR2_X1 U19675 ( .A1(n20954), .A2(n16773), .ZN(n16756) );
  NAND2_X1 U19676 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16756), .ZN(n16550) );
  NAND3_X1 U19677 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .A3(P3_REIP_REG_16__SCAN_IN), .ZN(n16535) );
  NAND4_X1 U19678 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(n16699), .A3(
        P3_REIP_REG_20__SCAN_IN), .A4(P3_REIP_REG_18__SCAN_IN), .ZN(n16650) );
  INV_X1 U19679 ( .A(n16650), .ZN(n16536) );
  INV_X1 U19680 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n18754) );
  INV_X1 U19681 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18750) );
  INV_X1 U19682 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18751) );
  NOR3_X1 U19683 ( .A1(n18754), .A2(n18750), .A3(n18751), .ZN(n16552) );
  NAND2_X1 U19684 ( .A1(n16536), .A2(n16552), .ZN(n16553) );
  NOR2_X1 U19685 ( .A1(n18755), .A2(n16553), .ZN(n16625) );
  INV_X1 U19686 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18758) );
  INV_X1 U19687 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18756) );
  NOR2_X1 U19688 ( .A1(n18758), .A2(n18756), .ZN(n16554) );
  INV_X1 U19689 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18759) );
  NOR2_X1 U19690 ( .A1(n18762), .A2(n18759), .ZN(n16587) );
  NAND3_X1 U19691 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16597), .A3(n16587), 
        .ZN(n16563) );
  NAND2_X1 U19692 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n18766), .ZN(n16562) );
  NOR4_X1 U19693 ( .A1(n18792), .A2(P3_STATE2_REG_2__SCAN_IN), .A3(
        P3_STATE2_REG_0__SCAN_IN), .A4(P3_STATEBS16_REG_SCAN_IN), .ZN(n16541)
         );
  NOR2_X1 U19694 ( .A1(n18782), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n18518) );
  INV_X1 U19695 ( .A(n18518), .ZN(n18686) );
  NOR2_X1 U19696 ( .A1(n16537), .A2(n18686), .ZN(n18682) );
  NOR4_X2 U19697 ( .A1(n18174), .A2(n18831), .A3(n16541), .A4(n18682), .ZN(
        n16909) );
  INV_X1 U19698 ( .A(n16538), .ZN(n16540) );
  AOI211_X4 U19699 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n18204), .A(n18677), .B(
        n16540), .ZN(n16888) );
  AOI22_X1 U19700 ( .A1(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n16889), .B1(
        P3_EBX_REG_31__SCAN_IN), .B2(n16888), .ZN(n16561) );
  NAND2_X1 U19701 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n18204), .ZN(n16539) );
  AOI211_X4 U19702 ( .C1(n18833), .C2(n18835), .A(n16540), .B(n16539), .ZN(
        n16884) );
  NOR3_X1 U19703 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16900) );
  NAND2_X1 U19704 ( .A1(n16900), .A2(n17207), .ZN(n16883) );
  NOR2_X1 U19705 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16883), .ZN(n16863) );
  INV_X1 U19706 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n17199) );
  NAND2_X1 U19707 ( .A1(n16863), .A2(n17199), .ZN(n16854) );
  NOR2_X1 U19708 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16854), .ZN(n16842) );
  INV_X1 U19709 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17194) );
  NAND2_X1 U19710 ( .A1(n16842), .A2(n17194), .ZN(n16829) );
  NOR2_X1 U19711 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16829), .ZN(n16820) );
  NAND2_X1 U19712 ( .A1(n16820), .A2(n17155), .ZN(n16808) );
  NOR2_X1 U19713 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16808), .ZN(n16790) );
  NAND2_X1 U19714 ( .A1(n16790), .A2(n17126), .ZN(n16787) );
  NOR2_X1 U19715 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16787), .ZN(n16771) );
  NAND2_X1 U19716 ( .A1(n16771), .A2(n16763), .ZN(n16762) );
  NOR2_X1 U19717 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16762), .ZN(n16746) );
  NAND2_X1 U19718 ( .A1(n16746), .A2(n16734), .ZN(n16732) );
  NOR2_X1 U19719 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16732), .ZN(n16713) );
  NAND2_X1 U19720 ( .A1(n16713), .A2(n17069), .ZN(n16709) );
  NOR2_X1 U19721 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16709), .ZN(n16692) );
  NAND2_X1 U19722 ( .A1(n16692), .A2(n17030), .ZN(n16685) );
  NOR2_X1 U19723 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16685), .ZN(n16669) );
  NAND2_X1 U19724 ( .A1(n16669), .A2(n17014), .ZN(n16664) );
  NOR2_X1 U19725 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16664), .ZN(n16655) );
  NAND2_X1 U19726 ( .A1(n16655), .A2(n16640), .ZN(n16639) );
  NOR2_X1 U19727 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16639), .ZN(n16617) );
  NAND2_X1 U19728 ( .A1(n16617), .A2(n16623), .ZN(n16605) );
  NOR2_X1 U19729 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16605), .ZN(n16604) );
  INV_X1 U19730 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16968) );
  NAND2_X1 U19731 ( .A1(n16604), .A2(n16968), .ZN(n16598) );
  NOR2_X1 U19732 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16598), .ZN(n16584) );
  NAND2_X1 U19733 ( .A1(n16584), .A2(n16955), .ZN(n16566) );
  NOR2_X1 U19734 ( .A1(n16921), .A2(n16566), .ZN(n16569) );
  INV_X1 U19735 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16559) );
  INV_X1 U19736 ( .A(n16541), .ZN(n18692) );
  INV_X1 U19737 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16585) );
  NAND2_X1 U19738 ( .A1(n16544), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n16543) );
  AOI21_X1 U19739 ( .B1(n16585), .B2(n16543), .A(n16542), .ZN(n17496) );
  INV_X1 U19740 ( .A(n17496), .ZN(n16592) );
  OAI21_X1 U19741 ( .B1(n16544), .B2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n16543), .ZN(n17509) );
  INV_X1 U19742 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n16607) );
  NAND2_X1 U19743 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17521), .ZN(
        n17495) );
  AOI21_X1 U19744 ( .B1(n16607), .B2(n17495), .A(n16544), .ZN(n17522) );
  INV_X1 U19745 ( .A(n17522), .ZN(n16612) );
  INV_X1 U19746 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17549) );
  NOR3_X1 U19747 ( .A1(n17855), .A2(n17533), .A3(n17549), .ZN(n16545) );
  OAI21_X1 U19748 ( .B1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n16545), .A(
        n17495), .ZN(n17536) );
  NOR2_X1 U19749 ( .A1(n17855), .A2(n17533), .ZN(n16547) );
  INV_X1 U19750 ( .A(n16545), .ZN(n16546) );
  OAI21_X1 U19751 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n16547), .A(
        n16546), .ZN(n17546) );
  INV_X1 U19752 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17561) );
  NAND2_X1 U19753 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17559), .ZN(
        n17532) );
  AOI21_X1 U19754 ( .B1(n17561), .B2(n17532), .A(n16547), .ZN(n17557) );
  INV_X1 U19755 ( .A(n17557), .ZN(n16643) );
  INV_X1 U19756 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17584) );
  INV_X1 U19757 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16702) );
  NOR2_X1 U19758 ( .A1(n17855), .A2(n17647), .ZN(n17646) );
  INV_X1 U19759 ( .A(n17646), .ZN(n16740) );
  NOR2_X1 U19760 ( .A1(n17648), .A2(n16740), .ZN(n16703) );
  INV_X1 U19761 ( .A(n16703), .ZN(n16715) );
  NOR2_X1 U19762 ( .A1(n16702), .A2(n16715), .ZN(n17608) );
  NAND2_X1 U19763 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n17608), .ZN(
        n16695) );
  INV_X1 U19764 ( .A(n16695), .ZN(n16682) );
  NAND2_X1 U19765 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n16682), .ZN(
        n16680) );
  INV_X1 U19766 ( .A(n16680), .ZN(n17570) );
  NAND2_X1 U19767 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n17570), .ZN(
        n16549) );
  NOR2_X1 U19768 ( .A1(n17584), .A2(n16549), .ZN(n16548) );
  OAI21_X1 U19769 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n16548), .A(
        n17532), .ZN(n17575) );
  XNOR2_X1 U19770 ( .A(n17584), .B(n16549), .ZN(n17581) );
  OAI21_X1 U19771 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16680), .A(
        n9653), .ZN(n16675) );
  OAI21_X1 U19772 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17570), .A(
        n16549), .ZN(n17597) );
  NAND2_X1 U19773 ( .A1(n16675), .A2(n17597), .ZN(n16674) );
  NAND2_X1 U19774 ( .A1(n9653), .A2(n16674), .ZN(n16663) );
  NAND2_X1 U19775 ( .A1(n17581), .A2(n16663), .ZN(n16662) );
  NAND2_X1 U19776 ( .A1(n9653), .A2(n16662), .ZN(n16654) );
  NAND2_X1 U19777 ( .A1(n17575), .A2(n16654), .ZN(n16653) );
  NAND2_X1 U19778 ( .A1(n9653), .A2(n16653), .ZN(n16642) );
  NAND2_X1 U19779 ( .A1(n16643), .A2(n16642), .ZN(n16641) );
  NAND2_X1 U19780 ( .A1(n9653), .A2(n16641), .ZN(n16634) );
  NAND2_X1 U19781 ( .A1(n17546), .A2(n16634), .ZN(n16633) );
  NAND2_X1 U19782 ( .A1(n9653), .A2(n16633), .ZN(n16619) );
  NAND2_X1 U19783 ( .A1(n17536), .A2(n16619), .ZN(n16618) );
  NAND2_X1 U19784 ( .A1(n9653), .A2(n16618), .ZN(n16611) );
  NAND2_X1 U19785 ( .A1(n16612), .A2(n16611), .ZN(n16610) );
  NAND2_X1 U19786 ( .A1(n9653), .A2(n16610), .ZN(n16600) );
  NAND2_X1 U19787 ( .A1(n17509), .A2(n16600), .ZN(n16599) );
  NAND2_X1 U19788 ( .A1(n9653), .A2(n16599), .ZN(n16591) );
  NAND2_X1 U19789 ( .A1(n16592), .A2(n16591), .ZN(n16590) );
  NAND2_X1 U19790 ( .A1(n9653), .A2(n16590), .ZN(n16579) );
  NAND2_X1 U19791 ( .A1(n16580), .A2(n16579), .ZN(n16578) );
  NOR4_X1 U19792 ( .A1(n16565), .A2(n16843), .A3(n18692), .A4(n16578), .ZN(
        n16558) );
  NAND2_X1 U19793 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16587), .ZN(n16555) );
  NAND3_X1 U19794 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_20__SCAN_IN), 
        .A3(P3_REIP_REG_18__SCAN_IN), .ZN(n16551) );
  INV_X1 U19795 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n20774) );
  NOR3_X1 U19796 ( .A1(n16909), .A2(n20774), .A3(n16550), .ZN(n16724) );
  NAND4_X1 U19797 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(P3_REIP_REG_15__SCAN_IN), 
        .A3(P3_REIP_REG_16__SCAN_IN), .A4(n16724), .ZN(n16679) );
  NOR2_X1 U19798 ( .A1(n16551), .A2(n16679), .ZN(n16649) );
  NAND2_X1 U19799 ( .A1(n16925), .A2(n16915), .ZN(n16923) );
  INV_X1 U19800 ( .A(n16923), .ZN(n16792) );
  AOI21_X1 U19801 ( .B1(n16552), .B2(n16649), .A(n16792), .ZN(n16638) );
  NOR2_X1 U19802 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16553), .ZN(n16630) );
  NOR2_X1 U19803 ( .A1(n16638), .A2(n16630), .ZN(n16627) );
  OAI21_X1 U19804 ( .B1(n16554), .B2(n16915), .A(n16627), .ZN(n16596) );
  AOI21_X1 U19805 ( .B1(n16899), .B2(n16555), .A(n16596), .ZN(n16583) );
  NOR2_X1 U19806 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n16563), .ZN(n16568) );
  INV_X1 U19807 ( .A(n16568), .ZN(n16556) );
  AOI21_X1 U19808 ( .B1(n16583), .B2(n16556), .A(n18766), .ZN(n16557) );
  AOI211_X1 U19809 ( .C1(n16569), .C2(n16559), .A(n16558), .B(n16557), .ZN(
        n16560) );
  OAI211_X1 U19810 ( .C1(n16563), .C2(n16562), .A(n16561), .B(n16560), .ZN(
        P3_U2640) );
  NAND2_X1 U19811 ( .A1(n9653), .A2(n16578), .ZN(n16564) );
  XOR2_X1 U19812 ( .A(n16565), .B(n16564), .Z(n16572) );
  NAND2_X1 U19813 ( .A1(n16884), .A2(n16566), .ZN(n16573) );
  INV_X1 U19814 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18768) );
  OAI22_X1 U19815 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16573), .B1(n16583), 
        .B2(n18768), .ZN(n16567) );
  AOI211_X1 U19816 ( .C1(n16889), .C2(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n16568), .B(n16567), .ZN(n16571) );
  OAI21_X1 U19817 ( .B1(n16888), .B2(n16569), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16570) );
  OAI211_X1 U19818 ( .C1(n18692), .C2(n16572), .A(n16571), .B(n16570), .ZN(
        P3_U2641) );
  INV_X1 U19819 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18763) );
  INV_X1 U19820 ( .A(n16584), .ZN(n16574) );
  AOI21_X1 U19821 ( .B1(P3_EBX_REG_29__SCAN_IN), .B2(n16574), .A(n16573), .ZN(
        n16577) );
  NAND2_X1 U19822 ( .A1(n16597), .A2(n16587), .ZN(n16575) );
  OAI22_X1 U19823 ( .A1(P3_REIP_REG_29__SCAN_IN), .A2(n16575), .B1(n16955), 
        .B2(n16922), .ZN(n16576) );
  AOI211_X1 U19824 ( .C1(n16889), .C2(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n16577), .B(n16576), .ZN(n16582) );
  INV_X1 U19825 ( .A(n18692), .ZN(n16910) );
  OAI211_X1 U19826 ( .C1(n16580), .C2(n16579), .A(n16910), .B(n16578), .ZN(
        n16581) );
  OAI211_X1 U19827 ( .C1(n16583), .C2(n18763), .A(n16582), .B(n16581), .ZN(
        P3_U2642) );
  INV_X1 U19828 ( .A(n16596), .ZN(n16616) );
  AOI211_X1 U19829 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16598), .A(n16584), .B(
        n16921), .ZN(n16589) );
  OAI21_X1 U19830 ( .B1(P3_REIP_REG_28__SCAN_IN), .B2(P3_REIP_REG_27__SCAN_IN), 
        .A(n16597), .ZN(n16586) );
  OAI22_X1 U19831 ( .A1(n16587), .A2(n16586), .B1(n16585), .B2(n16912), .ZN(
        n16588) );
  AOI211_X1 U19832 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16888), .A(n16589), .B(
        n16588), .ZN(n16594) );
  OAI211_X1 U19833 ( .C1(n16592), .C2(n16591), .A(n16910), .B(n16590), .ZN(
        n16593) );
  OAI211_X1 U19834 ( .C1(n16616), .C2(n18762), .A(n16594), .B(n16593), .ZN(
        P3_U2643) );
  INV_X1 U19835 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n20912) );
  OAI22_X1 U19836 ( .A1(n20912), .A2(n16912), .B1(n16922), .B2(n16968), .ZN(
        n16595) );
  AOI221_X1 U19837 ( .B1(n16597), .B2(n18759), .C1(n16596), .C2(
        P3_REIP_REG_27__SCAN_IN), .A(n16595), .ZN(n16603) );
  OAI211_X1 U19838 ( .C1(n16604), .C2(n16968), .A(n16884), .B(n16598), .ZN(
        n16602) );
  OAI211_X1 U19839 ( .C1(n17509), .C2(n16600), .A(n16910), .B(n16599), .ZN(
        n16601) );
  NAND3_X1 U19840 ( .A1(n16603), .A2(n16602), .A3(n16601), .ZN(P3_U2644) );
  AOI21_X1 U19841 ( .B1(P3_REIP_REG_25__SCAN_IN), .B2(n16625), .A(
        P3_REIP_REG_26__SCAN_IN), .ZN(n16615) );
  AOI211_X1 U19842 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16605), .A(n16604), .B(
        n16921), .ZN(n16609) );
  OAI22_X1 U19843 ( .A1(n16607), .A2(n16912), .B1(n16922), .B2(n16606), .ZN(
        n16608) );
  NOR2_X1 U19844 ( .A1(n16609), .A2(n16608), .ZN(n16614) );
  OAI211_X1 U19845 ( .C1(n16612), .C2(n16611), .A(n16910), .B(n16610), .ZN(
        n16613) );
  OAI211_X1 U19846 ( .C1(n16616), .C2(n16615), .A(n16614), .B(n16613), .ZN(
        P3_U2645) );
  AOI21_X1 U19847 ( .B1(n16884), .B2(n16617), .A(n16888), .ZN(n16622) );
  NOR2_X1 U19848 ( .A1(n16617), .A2(n16921), .ZN(n16632) );
  AOI22_X1 U19849 ( .A1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n16889), .B1(
        n16632), .B2(n16623), .ZN(n16621) );
  OAI211_X1 U19850 ( .C1(n17536), .C2(n16619), .A(n16910), .B(n16618), .ZN(
        n16620) );
  OAI211_X1 U19851 ( .C1(n16623), .C2(n16622), .A(n16621), .B(n16620), .ZN(
        n16624) );
  AOI21_X1 U19852 ( .B1(n16625), .B2(n18756), .A(n16624), .ZN(n16626) );
  OAI21_X1 U19853 ( .B1(n16627), .B2(n18756), .A(n16626), .ZN(P3_U2646) );
  INV_X1 U19854 ( .A(n16638), .ZN(n16637) );
  NAND2_X1 U19855 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16639), .ZN(n16631) );
  OAI22_X1 U19856 ( .A1(n17549), .A2(n16912), .B1(n16922), .B2(n16628), .ZN(
        n16629) );
  AOI211_X1 U19857 ( .C1(n16632), .C2(n16631), .A(n16630), .B(n16629), .ZN(
        n16636) );
  OAI211_X1 U19858 ( .C1(n17546), .C2(n16634), .A(n16910), .B(n16633), .ZN(
        n16635) );
  OAI211_X1 U19859 ( .C1(n16637), .C2(n18755), .A(n16636), .B(n16635), .ZN(
        P3_U2647) );
  AOI22_X1 U19860 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n16889), .B1(
        n16888), .B2(P3_EBX_REG_23__SCAN_IN), .ZN(n16647) );
  NOR2_X1 U19861 ( .A1(n18750), .A2(n16650), .ZN(n16648) );
  OAI221_X1 U19862 ( .B1(P3_REIP_REG_23__SCAN_IN), .B2(P3_REIP_REG_22__SCAN_IN), .C1(P3_REIP_REG_23__SCAN_IN), .C2(n16648), .A(n16638), .ZN(n16646) );
  OAI211_X1 U19863 ( .C1(n16655), .C2(n16640), .A(n16884), .B(n16639), .ZN(
        n16645) );
  OAI211_X1 U19864 ( .C1(n16643), .C2(n16642), .A(n16910), .B(n16641), .ZN(
        n16644) );
  NAND4_X1 U19865 ( .A1(n16647), .A2(n16646), .A3(n16645), .A4(n16644), .ZN(
        P3_U2648) );
  AOI22_X1 U19866 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n16889), .B1(
        n16888), .B2(P3_EBX_REG_22__SCAN_IN), .ZN(n16660) );
  INV_X1 U19867 ( .A(n16648), .ZN(n16652) );
  NOR2_X1 U19868 ( .A1(n16792), .A2(n16649), .ZN(n16673) );
  NOR2_X1 U19869 ( .A1(P3_REIP_REG_21__SCAN_IN), .A2(n16650), .ZN(n16661) );
  NOR2_X1 U19870 ( .A1(n16673), .A2(n16661), .ZN(n16651) );
  MUX2_X1 U19871 ( .A(n16652), .B(n16651), .S(P3_REIP_REG_22__SCAN_IN), .Z(
        n16659) );
  OAI211_X1 U19872 ( .C1(n17575), .C2(n16654), .A(n16910), .B(n16653), .ZN(
        n16658) );
  AOI211_X1 U19873 ( .C1(n16664), .C2(P3_EBX_REG_22__SCAN_IN), .A(n16921), .B(
        n16655), .ZN(n16656) );
  INV_X1 U19874 ( .A(n16656), .ZN(n16657) );
  NAND4_X1 U19875 ( .A1(n16660), .A2(n16659), .A3(n16658), .A4(n16657), .ZN(
        P3_U2649) );
  AOI22_X1 U19876 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n16889), .B1(
        n16888), .B2(P3_EBX_REG_21__SCAN_IN), .ZN(n16668) );
  AOI21_X1 U19877 ( .B1(n16673), .B2(P3_REIP_REG_21__SCAN_IN), .A(n16661), 
        .ZN(n16667) );
  OAI211_X1 U19878 ( .C1(n17581), .C2(n16663), .A(n16910), .B(n16662), .ZN(
        n16666) );
  OAI211_X1 U19879 ( .C1(n16669), .C2(n17014), .A(n16884), .B(n16664), .ZN(
        n16665) );
  NAND4_X1 U19880 ( .A1(n16668), .A2(n16667), .A3(n16666), .A4(n16665), .ZN(
        P3_U2650) );
  AOI211_X1 U19881 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16685), .A(n16669), .B(
        n16921), .ZN(n16672) );
  AOI22_X1 U19882 ( .A1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n16889), .B1(
        n16888), .B2(P3_EBX_REG_20__SCAN_IN), .ZN(n16670) );
  INV_X1 U19883 ( .A(n16670), .ZN(n16671) );
  AOI211_X1 U19884 ( .C1(n16673), .C2(P3_REIP_REG_20__SCAN_IN), .A(n16672), 
        .B(n16671), .ZN(n16678) );
  OAI211_X1 U19885 ( .C1(n16675), .C2(n17597), .A(n16910), .B(n16674), .ZN(
        n16677) );
  INV_X1 U19886 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18747) );
  NAND4_X1 U19887 ( .A1(n16699), .A2(P3_REIP_REG_19__SCAN_IN), .A3(
        P3_REIP_REG_18__SCAN_IN), .A4(n18747), .ZN(n16676) );
  NAND3_X1 U19888 ( .A1(n16678), .A2(n16677), .A3(n16676), .ZN(P3_U2651) );
  INV_X1 U19889 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18746) );
  NAND2_X1 U19890 ( .A1(n16923), .A2(n16679), .ZN(n16694) );
  OAI21_X1 U19891 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16682), .A(
        n16680), .ZN(n16681) );
  INV_X1 U19892 ( .A(n16681), .ZN(n17609) );
  INV_X1 U19893 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16914) );
  INV_X1 U19894 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17659) );
  NOR2_X1 U19895 ( .A1(n17659), .A2(n16740), .ZN(n16728) );
  AOI21_X1 U19896 ( .B1(n16914), .B2(n16728), .A(n16843), .ZN(n16716) );
  INV_X1 U19897 ( .A(n16716), .ZN(n16727) );
  OAI21_X1 U19898 ( .B1(n16682), .B2(n16843), .A(n16727), .ZN(n16684) );
  OAI21_X1 U19899 ( .B1(n17609), .B2(n16684), .A(n16910), .ZN(n16683) );
  AOI21_X1 U19900 ( .B1(n17609), .B2(n16684), .A(n16683), .ZN(n16688) );
  OAI211_X1 U19901 ( .C1(n16692), .C2(n17030), .A(n16884), .B(n16685), .ZN(
        n16686) );
  OAI211_X1 U19902 ( .C1(n16922), .C2(n17030), .A(n9642), .B(n16686), .ZN(
        n16687) );
  AOI211_X1 U19903 ( .C1(n16889), .C2(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n16688), .B(n16687), .ZN(n16691) );
  NAND2_X1 U19904 ( .A1(P3_REIP_REG_19__SCAN_IN), .A2(P3_REIP_REG_18__SCAN_IN), 
        .ZN(n16689) );
  OAI211_X1 U19905 ( .C1(P3_REIP_REG_19__SCAN_IN), .C2(P3_REIP_REG_18__SCAN_IN), .A(n16699), .B(n16689), .ZN(n16690) );
  OAI211_X1 U19906 ( .C1(n18746), .C2(n16694), .A(n16691), .B(n16690), .ZN(
        P3_U2652) );
  INV_X1 U19907 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17623) );
  AOI211_X1 U19908 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16709), .A(n16692), .B(
        n16921), .ZN(n16693) );
  AOI211_X1 U19909 ( .C1(n16888), .C2(P3_EBX_REG_18__SCAN_IN), .A(n18174), .B(
        n16693), .ZN(n16701) );
  INV_X1 U19910 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18743) );
  INV_X1 U19911 ( .A(n16694), .ZN(n16708) );
  OAI21_X1 U19912 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17608), .A(
        n16695), .ZN(n17620) );
  NOR2_X1 U19913 ( .A1(n17855), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16867) );
  INV_X1 U19914 ( .A(n16867), .ZN(n16893) );
  OAI21_X1 U19915 ( .B1(n17615), .B2(n16893), .A(n9653), .ZN(n16697) );
  OAI21_X1 U19916 ( .B1(n17620), .B2(n16697), .A(n16910), .ZN(n16696) );
  AOI21_X1 U19917 ( .B1(n17620), .B2(n16697), .A(n16696), .ZN(n16698) );
  AOI221_X1 U19918 ( .B1(n16699), .B2(n18743), .C1(n16708), .C2(
        P3_REIP_REG_18__SCAN_IN), .A(n16698), .ZN(n16700) );
  OAI211_X1 U19919 ( .C1(n17623), .C2(n16912), .A(n16701), .B(n16700), .ZN(
        P3_U2653) );
  AOI22_X1 U19920 ( .A1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n16889), .B1(
        n16888), .B2(P3_EBX_REG_17__SCAN_IN), .ZN(n16712) );
  AOI21_X1 U19921 ( .B1(n16702), .B2(n16715), .A(n17608), .ZN(n17634) );
  AOI21_X1 U19922 ( .B1(n16703), .B2(n16914), .A(n16843), .ZN(n16705) );
  OAI21_X1 U19923 ( .B1(n17634), .B2(n16705), .A(n16910), .ZN(n16704) );
  AOI21_X1 U19924 ( .B1(n17634), .B2(n16705), .A(n16704), .ZN(n16707) );
  INV_X1 U19925 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n20773) );
  INV_X1 U19926 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18739) );
  NOR4_X1 U19927 ( .A1(P3_REIP_REG_17__SCAN_IN), .A2(n16738), .A3(n20773), 
        .A4(n18739), .ZN(n16706) );
  AOI211_X1 U19928 ( .C1(n16708), .C2(P3_REIP_REG_17__SCAN_IN), .A(n16707), 
        .B(n16706), .ZN(n16711) );
  OAI211_X1 U19929 ( .C1(n16713), .C2(n17069), .A(n16884), .B(n16709), .ZN(
        n16710) );
  NAND4_X1 U19930 ( .A1(n16712), .A2(n16711), .A3(n9642), .A4(n16710), .ZN(
        P3_U2654) );
  INV_X1 U19931 ( .A(P3_EBX_REG_16__SCAN_IN), .ZN(n16723) );
  AOI211_X1 U19932 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16732), .A(n16713), .B(
        n16921), .ZN(n16714) );
  AOI211_X1 U19933 ( .C1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .C2(n16889), .A(
        n18174), .B(n16714), .ZN(n16722) );
  OAI22_X1 U19934 ( .A1(P3_REIP_REG_15__SCAN_IN), .A2(n16738), .B1(n16792), 
        .B2(n16724), .ZN(n16720) );
  OAI21_X1 U19935 ( .B1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n16728), .A(
        n16715), .ZN(n17651) );
  INV_X1 U19936 ( .A(n17651), .ZN(n16717) );
  AOI221_X1 U19937 ( .B1(n16717), .B2(n16716), .C1(n17651), .C2(n16727), .A(
        n18692), .ZN(n16719) );
  NOR3_X1 U19938 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n20773), .A3(n16738), 
        .ZN(n16718) );
  AOI211_X1 U19939 ( .C1(P3_REIP_REG_16__SCAN_IN), .C2(n16720), .A(n16719), 
        .B(n16718), .ZN(n16721) );
  OAI211_X1 U19940 ( .C1(n16922), .C2(n16723), .A(n16722), .B(n16721), .ZN(
        P3_U2655) );
  INV_X1 U19941 ( .A(n16724), .ZN(n16743) );
  NAND2_X1 U19942 ( .A1(n16923), .A2(n16743), .ZN(n16752) );
  NOR2_X1 U19943 ( .A1(n16843), .A2(n16914), .ZN(n16725) );
  NOR2_X1 U19944 ( .A1(n16725), .A2(n18692), .ZN(n16918) );
  OAI21_X1 U19945 ( .B1(n17646), .B2(n16843), .A(n16918), .ZN(n16726) );
  INV_X1 U19946 ( .A(n16726), .ZN(n16731) );
  NOR2_X1 U19947 ( .A1(n16727), .A2(n18692), .ZN(n16730) );
  AOI21_X1 U19948 ( .B1(n17659), .B2(n16740), .A(n16728), .ZN(n16729) );
  INV_X1 U19949 ( .A(n16729), .ZN(n17656) );
  MUX2_X1 U19950 ( .A(n16731), .B(n16730), .S(n17656), .Z(n16736) );
  OAI211_X1 U19951 ( .C1(n16746), .C2(n16734), .A(n16884), .B(n16732), .ZN(
        n16733) );
  OAI211_X1 U19952 ( .C1(n16922), .C2(n16734), .A(n9642), .B(n16733), .ZN(
        n16735) );
  AOI211_X1 U19953 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n16889), .A(
        n16736), .B(n16735), .ZN(n16737) );
  OAI221_X1 U19954 ( .B1(P3_REIP_REG_15__SCAN_IN), .B2(n16738), .C1(n20773), 
        .C2(n16752), .A(n16737), .ZN(P3_U2656) );
  INV_X1 U19955 ( .A(n17757), .ZN(n17760) );
  NOR2_X1 U19956 ( .A1(n17855), .A2(n17760), .ZN(n16828) );
  NAND2_X1 U19957 ( .A1(n16739), .A2(n16828), .ZN(n17684) );
  NOR2_X1 U19958 ( .A1(n17697), .A2(n17684), .ZN(n16753) );
  OAI21_X1 U19959 ( .B1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n16753), .A(
        n16740), .ZN(n17673) );
  NOR2_X1 U19960 ( .A1(n18692), .A2(n17673), .ZN(n16742) );
  AOI21_X1 U19961 ( .B1(n17672), .B2(n16867), .A(n16843), .ZN(n16741) );
  INV_X1 U19962 ( .A(n16741), .ZN(n16745) );
  AOI22_X1 U19963 ( .A1(n16744), .A2(n16743), .B1(n16742), .B2(n16745), .ZN(
        n16751) );
  NOR2_X1 U19964 ( .A1(n18692), .A2(n16745), .ZN(n16755) );
  AOI211_X1 U19965 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16762), .A(n16746), .B(
        n16921), .ZN(n16749) );
  AOI22_X1 U19966 ( .A1(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n16889), .B1(
        n16888), .B2(P3_EBX_REG_14__SCAN_IN), .ZN(n16747) );
  NAND2_X1 U19967 ( .A1(n16747), .A2(n9642), .ZN(n16748) );
  AOI211_X1 U19968 ( .C1(n16755), .C2(n17673), .A(n16749), .B(n16748), .ZN(
        n16750) );
  OAI211_X1 U19969 ( .C1(n20774), .C2(n16752), .A(n16751), .B(n16750), .ZN(
        P3_U2657) );
  INV_X1 U19970 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16757) );
  INV_X1 U19971 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17704) );
  NOR2_X1 U19972 ( .A1(n17704), .A2(n17684), .ZN(n16761) );
  INV_X1 U19973 ( .A(n16761), .ZN(n16768) );
  AOI21_X1 U19974 ( .B1(n16757), .B2(n16768), .A(n16753), .ZN(n17687) );
  INV_X1 U19975 ( .A(n17687), .ZN(n16754) );
  AOI22_X1 U19976 ( .A1(n16888), .A2(P3_EBX_REG_13__SCAN_IN), .B1(n16755), 
        .B2(n16754), .ZN(n16767) );
  AOI21_X1 U19977 ( .B1(n16899), .B2(n16773), .A(n16909), .ZN(n16784) );
  OAI21_X1 U19978 ( .B1(P3_REIP_REG_12__SCAN_IN), .B2(n16915), .A(n16784), 
        .ZN(n16760) );
  NAND2_X1 U19979 ( .A1(n16899), .A2(n16756), .ZN(n16758) );
  OAI22_X1 U19980 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16758), .B1(n16757), 
        .B2(n16912), .ZN(n16759) );
  AOI211_X1 U19981 ( .C1(P3_REIP_REG_13__SCAN_IN), .C2(n16760), .A(n18174), 
        .B(n16759), .ZN(n16766) );
  OAI211_X1 U19982 ( .C1(n16761), .C2(n16843), .A(n17687), .B(n16918), .ZN(
        n16765) );
  OAI211_X1 U19983 ( .C1(n16771), .C2(n16763), .A(n16884), .B(n16762), .ZN(
        n16764) );
  NAND4_X1 U19984 ( .A1(n16767), .A2(n16766), .A3(n16765), .A4(n16764), .ZN(
        P3_U2658) );
  AOI22_X1 U19985 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n16889), .B1(
        n16888), .B2(P3_EBX_REG_12__SCAN_IN), .ZN(n16778) );
  INV_X1 U19986 ( .A(n17684), .ZN(n16769) );
  AOI21_X1 U19987 ( .B1(n16769), .B2(n16914), .A(n16843), .ZN(n16770) );
  OAI21_X1 U19988 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n16769), .A(
        n16768), .ZN(n17714) );
  XNOR2_X1 U19989 ( .A(n16770), .B(n17714), .ZN(n16776) );
  AOI211_X1 U19990 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16787), .A(n16771), .B(
        n16921), .ZN(n16775) );
  NAND2_X1 U19991 ( .A1(n16899), .A2(n20954), .ZN(n16772) );
  OAI21_X1 U19992 ( .B1(n16773), .B2(n16772), .A(n9642), .ZN(n16774) );
  AOI211_X1 U19993 ( .C1(n16776), .C2(n16910), .A(n16775), .B(n16774), .ZN(
        n16777) );
  OAI211_X1 U19994 ( .C1(n20954), .C2(n16784), .A(n16778), .B(n16777), .ZN(
        P3_U2659) );
  NAND2_X1 U19995 ( .A1(n16899), .A2(n16833), .ZN(n16834) );
  INV_X1 U19996 ( .A(n16834), .ZN(n16779) );
  NAND2_X1 U19997 ( .A1(n16794), .A2(n16779), .ZN(n16813) );
  INV_X1 U19998 ( .A(n16813), .ZN(n16780) );
  AOI21_X1 U19999 ( .B1(n16795), .B2(n16780), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16785) );
  INV_X1 U20000 ( .A(n16828), .ZN(n16838) );
  NOR2_X1 U20001 ( .A1(n16781), .A2(n16838), .ZN(n16796) );
  AOI21_X1 U20002 ( .B1(n16796), .B2(n16914), .A(n16843), .ZN(n16782) );
  OAI21_X1 U20003 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16796), .A(
        n17684), .ZN(n17731) );
  XOR2_X1 U20004 ( .A(n16782), .B(n17731), .Z(n16783) );
  OAI22_X1 U20005 ( .A1(n16785), .A2(n16784), .B1(n18692), .B2(n16783), .ZN(
        n16786) );
  AOI211_X1 U20006 ( .C1(n16888), .C2(P3_EBX_REG_11__SCAN_IN), .A(n16412), .B(
        n16786), .ZN(n16789) );
  OAI211_X1 U20007 ( .C1(n16790), .C2(n17126), .A(n16884), .B(n16787), .ZN(
        n16788) );
  OAI211_X1 U20008 ( .C1(n16912), .C2(n17720), .A(n16789), .B(n16788), .ZN(
        P3_U2660) );
  INV_X1 U20009 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17737) );
  AOI211_X1 U20010 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16808), .A(n16790), .B(
        n16921), .ZN(n16791) );
  AOI211_X1 U20011 ( .C1(n16888), .C2(P3_EBX_REG_10__SCAN_IN), .A(n18174), .B(
        n16791), .ZN(n16801) );
  AND2_X1 U20012 ( .A1(n16925), .A2(n16833), .ZN(n16793) );
  AOI21_X1 U20013 ( .B1(n16794), .B2(n16793), .A(n16792), .ZN(n16802) );
  AOI211_X1 U20014 ( .C1(n18731), .C2(n18729), .A(n16795), .B(n16813), .ZN(
        n16799) );
  NOR2_X1 U20015 ( .A1(n17717), .A2(n16838), .ZN(n16816) );
  NAND2_X1 U20016 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n16816), .ZN(
        n16803) );
  AOI21_X1 U20017 ( .B1(n17737), .B2(n16803), .A(n16796), .ZN(n17733) );
  INV_X1 U20018 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n17761) );
  NAND3_X1 U20019 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17757), .A3(
        P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n16827) );
  NOR3_X1 U20020 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n17761), .A3(
        n16827), .ZN(n16805) );
  AOI21_X1 U20021 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16805), .A(
        n16843), .ZN(n16804) );
  OAI21_X1 U20022 ( .B1(n17733), .B2(n16804), .A(n16910), .ZN(n16797) );
  AOI21_X1 U20023 ( .B1(n17733), .B2(n16804), .A(n16797), .ZN(n16798) );
  AOI211_X1 U20024 ( .C1(P3_REIP_REG_10__SCAN_IN), .C2(n16802), .A(n16799), 
        .B(n16798), .ZN(n16800) );
  OAI211_X1 U20025 ( .C1(n17737), .C2(n16912), .A(n16801), .B(n16800), .ZN(
        P3_U2661) );
  INV_X1 U20026 ( .A(n16802), .ZN(n16825) );
  OAI21_X1 U20027 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16816), .A(
        n16803), .ZN(n17749) );
  INV_X1 U20028 ( .A(n16804), .ZN(n16807) );
  NAND2_X1 U20029 ( .A1(n16910), .A2(n16843), .ZN(n16895) );
  OAI21_X1 U20030 ( .B1(n16805), .B2(n17749), .A(n16910), .ZN(n16806) );
  AOI22_X1 U20031 ( .A1(n17749), .A2(n16807), .B1(n16895), .B2(n16806), .ZN(
        n16811) );
  OAI211_X1 U20032 ( .C1(n16820), .C2(n17155), .A(n16884), .B(n16808), .ZN(
        n16809) );
  OAI211_X1 U20033 ( .C1(n16922), .C2(n17155), .A(n9642), .B(n16809), .ZN(
        n16810) );
  AOI211_X1 U20034 ( .C1(n16889), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n16811), .B(n16810), .ZN(n16812) );
  OAI221_X1 U20035 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(n16813), .C1(n18729), 
        .C2(n16825), .A(n16812), .ZN(P3_U2662) );
  NOR3_X1 U20036 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16814), .A3(n16834), .ZN(
        n16815) );
  AOI211_X1 U20037 ( .C1(n16888), .C2(P3_EBX_REG_8__SCAN_IN), .A(n18174), .B(
        n16815), .ZN(n16824) );
  AOI21_X1 U20038 ( .B1(n17761), .B2(n16827), .A(n16816), .ZN(n17764) );
  NOR2_X1 U20039 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16827), .ZN(
        n16817) );
  NOR2_X1 U20040 ( .A1(n16817), .A2(n16843), .ZN(n16819) );
  OAI21_X1 U20041 ( .B1(n17764), .B2(n16819), .A(n16910), .ZN(n16818) );
  AOI21_X1 U20042 ( .B1(n17764), .B2(n16819), .A(n16818), .ZN(n16822) );
  AOI211_X1 U20043 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16829), .A(n16820), .B(
        n16921), .ZN(n16821) );
  AOI211_X1 U20044 ( .C1(n16889), .C2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n16822), .B(n16821), .ZN(n16823) );
  OAI211_X1 U20045 ( .C1(n18728), .C2(n16825), .A(n16824), .B(n16823), .ZN(
        P3_U2663) );
  NOR2_X1 U20046 ( .A1(P3_REIP_REG_7__SCAN_IN), .A2(n16834), .ZN(n16826) );
  AOI22_X1 U20047 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n16889), .B1(
        P3_REIP_REG_6__SCAN_IN), .B2(n16826), .ZN(n16837) );
  AOI21_X1 U20048 ( .B1(n16914), .B2(n16828), .A(n16843), .ZN(n16840) );
  OAI21_X1 U20049 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n16828), .A(
        n16827), .ZN(n17786) );
  XNOR2_X1 U20050 ( .A(n16840), .B(n17786), .ZN(n16832) );
  OAI211_X1 U20051 ( .C1(n16842), .C2(n17194), .A(n16884), .B(n16829), .ZN(
        n16830) );
  OAI21_X1 U20052 ( .B1(n17194), .B2(n16922), .A(n16830), .ZN(n16831) );
  AOI21_X1 U20053 ( .B1(n16832), .B2(n16910), .A(n16831), .ZN(n16836) );
  OAI21_X1 U20054 ( .B1(n16833), .B2(n16915), .A(n16925), .ZN(n16860) );
  NOR2_X1 U20055 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16834), .ZN(n16841) );
  OAI21_X1 U20056 ( .B1(n16860), .B2(n16841), .A(P3_REIP_REG_7__SCAN_IN), .ZN(
        n16835) );
  NAND4_X1 U20057 ( .A1(n16837), .A2(n16836), .A3(n9642), .A4(n16835), .ZN(
        P3_U2664) );
  NOR2_X1 U20058 ( .A1(n17855), .A2(n17716), .ZN(n16851) );
  OAI21_X1 U20059 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16851), .A(
        n16838), .ZN(n16839) );
  INV_X1 U20060 ( .A(n16839), .ZN(n17791) );
  NAND2_X1 U20061 ( .A1(n16910), .A2(n16840), .ZN(n16849) );
  AOI211_X1 U20062 ( .C1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .C2(n16889), .A(
        n18174), .B(n16841), .ZN(n16848) );
  AOI211_X1 U20063 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16854), .A(n16842), .B(
        n16921), .ZN(n16846) );
  INV_X1 U20064 ( .A(P3_EBX_REG_6__SCAN_IN), .ZN(n17193) );
  OAI211_X1 U20065 ( .C1(n17789), .C2(n16843), .A(n17791), .B(n16918), .ZN(
        n16844) );
  OAI21_X1 U20066 ( .B1(n17193), .B2(n16922), .A(n16844), .ZN(n16845) );
  AOI211_X1 U20067 ( .C1(n16860), .C2(P3_REIP_REG_6__SCAN_IN), .A(n16846), .B(
        n16845), .ZN(n16847) );
  OAI211_X1 U20068 ( .C1(n17791), .C2(n16849), .A(n16848), .B(n16847), .ZN(
        P3_U2665) );
  OAI21_X1 U20069 ( .B1(n16915), .B2(n16850), .A(n18722), .ZN(n16859) );
  INV_X1 U20070 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16857) );
  NAND2_X1 U20071 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17806), .ZN(
        n16862) );
  AOI21_X1 U20072 ( .B1(n16857), .B2(n16862), .A(n16851), .ZN(n16853) );
  OAI21_X1 U20073 ( .B1(n16862), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n9653), .ZN(n16852) );
  INV_X1 U20074 ( .A(n16852), .ZN(n16866) );
  INV_X1 U20075 ( .A(n16853), .ZN(n17809) );
  OAI221_X1 U20076 ( .B1(n16853), .B2(n16866), .C1(n17809), .C2(n16852), .A(
        n16910), .ZN(n16856) );
  OAI211_X1 U20077 ( .C1(n16863), .C2(n17199), .A(n16884), .B(n16854), .ZN(
        n16855) );
  OAI211_X1 U20078 ( .C1(n16912), .C2(n16857), .A(n16856), .B(n16855), .ZN(
        n16858) );
  AOI21_X1 U20079 ( .B1(n16860), .B2(n16859), .A(n16858), .ZN(n16861) );
  OAI211_X1 U20080 ( .C1(n16922), .C2(n17199), .A(n16861), .B(n9642), .ZN(
        P3_U2666) );
  NOR2_X1 U20081 ( .A1(n17855), .A2(n17818), .ZN(n16876) );
  OAI21_X1 U20082 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16876), .A(
        n16862), .ZN(n17821) );
  AOI211_X1 U20083 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16883), .A(n16863), .B(
        n16921), .ZN(n16873) );
  NOR2_X1 U20084 ( .A1(n18196), .A2(n18846), .ZN(n16908) );
  INV_X1 U20085 ( .A(n16908), .ZN(n18848) );
  OAI221_X1 U20086 ( .B1(n18848), .B2(n9675), .C1(n18848), .C2(n16864), .A(
        n9642), .ZN(n16872) );
  OAI22_X1 U20087 ( .A1(n17820), .A2(n16912), .B1(n16922), .B2(n16865), .ZN(
        n16871) );
  NOR2_X1 U20088 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n17818), .ZN(
        n17814) );
  AOI22_X1 U20089 ( .A1(n16867), .A2(n17814), .B1(n16866), .B2(n17821), .ZN(
        n16869) );
  INV_X1 U20090 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18719) );
  NAND3_X1 U20091 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(P3_REIP_REG_1__SCAN_IN), 
        .A3(P3_REIP_REG_2__SCAN_IN), .ZN(n16868) );
  AOI21_X1 U20092 ( .B1(n16899), .B2(n16868), .A(n16909), .ZN(n16878) );
  OAI22_X1 U20093 ( .A1(n16869), .A2(n18692), .B1(n18719), .B2(n16878), .ZN(
        n16870) );
  NOR4_X1 U20094 ( .A1(n16873), .A2(n16872), .A3(n16871), .A4(n16870), .ZN(
        n16875) );
  NAND2_X1 U20095 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16898) );
  NOR2_X1 U20096 ( .A1(n16915), .A2(n16898), .ZN(n16877) );
  NAND3_X1 U20097 ( .A1(P3_REIP_REG_3__SCAN_IN), .A2(n16877), .A3(n18719), 
        .ZN(n16874) );
  OAI211_X1 U20098 ( .C1(n16895), .C2(n17821), .A(n16875), .B(n16874), .ZN(
        P3_U2667) );
  INV_X1 U20099 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16887) );
  NAND2_X1 U20100 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16891) );
  AOI21_X1 U20101 ( .B1(n16887), .B2(n16891), .A(n16876), .ZN(n17831) );
  OAI21_X1 U20102 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16891), .A(
        n9653), .ZN(n16892) );
  XNOR2_X1 U20103 ( .A(n17831), .B(n16892), .ZN(n16882) );
  INV_X1 U20104 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18717) );
  INV_X1 U20105 ( .A(n16877), .ZN(n16879) );
  AOI21_X1 U20106 ( .B1(n18717), .B2(n16879), .A(n16878), .ZN(n16881) );
  NOR2_X1 U20107 ( .A1(n18813), .A2(n18659), .ZN(n16890) );
  INV_X1 U20108 ( .A(n16890), .ZN(n18654) );
  AOI21_X1 U20109 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18654), .A(
        n17144), .ZN(n18784) );
  OAI22_X1 U20110 ( .A1(n18784), .A2(n18848), .B1(n16922), .B2(n17207), .ZN(
        n16880) );
  AOI211_X1 U20111 ( .C1(n16910), .C2(n16882), .A(n16881), .B(n16880), .ZN(
        n16886) );
  OAI211_X1 U20112 ( .C1(n16900), .C2(n17207), .A(n16884), .B(n16883), .ZN(
        n16885) );
  OAI211_X1 U20113 ( .C1(n16912), .C2(n16887), .A(n16886), .B(n16885), .ZN(
        P3_U2668) );
  AOI22_X1 U20114 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n16889), .B1(
        n16888), .B2(P3_EBX_REG_2__SCAN_IN), .ZN(n16906) );
  AOI21_X1 U20115 ( .B1(n18799), .B2(n18656), .A(n16890), .ZN(n18795) );
  OAI21_X1 U20116 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16891), .ZN(n17841) );
  INV_X1 U20117 ( .A(n17841), .ZN(n16894) );
  AOI211_X1 U20118 ( .C1(n16894), .C2(n16893), .A(n18692), .B(n16892), .ZN(
        n16897) );
  INV_X1 U20119 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18715) );
  OAI22_X1 U20120 ( .A1(n16925), .A2(n18715), .B1(n17841), .B2(n16895), .ZN(
        n16896) );
  AOI211_X1 U20121 ( .C1(n16908), .C2(n18795), .A(n16897), .B(n16896), .ZN(
        n16905) );
  OAI211_X1 U20122 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16899), .B(n16898), .ZN(n16904) );
  OR2_X1 U20123 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), .ZN(
        n16901) );
  AOI211_X1 U20124 ( .C1(n16901), .C2(P3_EBX_REG_2__SCAN_IN), .A(n16921), .B(
        n16900), .ZN(n16902) );
  INV_X1 U20125 ( .A(n16902), .ZN(n16903) );
  NAND4_X1 U20126 ( .A1(n16906), .A2(n16905), .A3(n16904), .A4(n16903), .ZN(
        P3_U2669) );
  NAND2_X1 U20127 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .ZN(n17215) );
  OAI21_X1 U20128 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(P3_EBX_REG_1__SCAN_IN), 
        .A(n17215), .ZN(n17224) );
  AND2_X1 U20129 ( .A1(n16907), .A2(n18656), .ZN(n18803) );
  AOI22_X1 U20130 ( .A1(n16909), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n18803), 
        .B2(n16908), .ZN(n16920) );
  NAND2_X1 U20131 ( .A1(n9653), .A2(n16910), .ZN(n16913) );
  OAI21_X1 U20132 ( .B1(n16914), .B2(n16913), .A(n16912), .ZN(n16917) );
  INV_X1 U20133 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17223) );
  OAI22_X1 U20134 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16915), .B1(n16922), 
        .B2(n17223), .ZN(n16916) );
  AOI221_X1 U20135 ( .B1(n16918), .B2(n17855), .C1(n16917), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n16916), .ZN(n16919) );
  OAI211_X1 U20136 ( .C1(n16921), .C2(n17224), .A(n16920), .B(n16919), .ZN(
        P3_U2670) );
  NAND2_X1 U20137 ( .A1(n16922), .A2(n16921), .ZN(n16924) );
  AOI22_X1 U20138 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n16924), .B1(
        P3_REIP_REG_0__SCAN_IN), .B2(n16923), .ZN(n16927) );
  NAND3_X1 U20139 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18844), .A3(
        n16925), .ZN(n16926) );
  OAI211_X1 U20140 ( .C1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n18848), .A(
        n16927), .B(n16926), .ZN(P3_U2671) );
  NOR2_X1 U20141 ( .A1(P3_EBX_REG_30__SCAN_IN), .A2(n16928), .ZN(n16954) );
  AOI22_X1 U20142 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n16940) );
  AOI22_X1 U20143 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16939) );
  AOI22_X1 U20144 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16930) );
  OAI21_X1 U20145 ( .B1(n16931), .B2(n17197), .A(n16930), .ZN(n16937) );
  AOI22_X1 U20146 ( .A1(n9634), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16935) );
  AOI22_X1 U20147 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n9639), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n16934) );
  AOI22_X1 U20148 ( .A1(n15584), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16933) );
  AOI22_X1 U20149 ( .A1(n17128), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9637), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16932) );
  NAND4_X1 U20150 ( .A1(n16935), .A2(n16934), .A3(n16933), .A4(n16932), .ZN(
        n16936) );
  AOI211_X1 U20151 ( .C1(n17174), .C2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A(
        n16937), .B(n16936), .ZN(n16938) );
  NAND3_X1 U20152 ( .A1(n16940), .A2(n16939), .A3(n16938), .ZN(n16952) );
  AOI22_X1 U20153 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(n9639), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16944) );
  AOI22_X1 U20154 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16943) );
  AOI22_X1 U20155 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17128), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16942) );
  AOI22_X1 U20156 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16941) );
  NAND4_X1 U20157 ( .A1(n16944), .A2(n16943), .A3(n16942), .A4(n16941), .ZN(
        n16950) );
  AOI22_X1 U20158 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9641), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16948) );
  AOI22_X1 U20159 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16947) );
  AOI22_X1 U20160 ( .A1(n15584), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9637), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16946) );
  AOI22_X1 U20161 ( .A1(n14026), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16945) );
  NAND4_X1 U20162 ( .A1(n16948), .A2(n16947), .A3(n16946), .A4(n16945), .ZN(
        n16949) );
  NOR2_X1 U20163 ( .A1(n16950), .A2(n16949), .ZN(n16958) );
  NOR3_X1 U20164 ( .A1(n16958), .A2(n16956), .A3(n16957), .ZN(n16951) );
  XNOR2_X1 U20165 ( .A(n16952), .B(n16951), .ZN(n17240) );
  OAI22_X1 U20166 ( .A1(n16954), .A2(n16953), .B1(n17240), .B2(n17220), .ZN(
        P3_U2673) );
  NAND2_X1 U20167 ( .A1(n17012), .A2(n16955), .ZN(n16962) );
  NOR2_X1 U20168 ( .A1(n16957), .A2(n16956), .ZN(n16959) );
  XNOR2_X1 U20169 ( .A(n16959), .B(n16958), .ZN(n17241) );
  AOI22_X1 U20170 ( .A1(P3_EBX_REG_29__SCAN_IN), .A2(n16960), .B1(n17226), 
        .B2(n17241), .ZN(n16961) );
  OAI21_X1 U20171 ( .B1(n16963), .B2(n16962), .A(n16961), .ZN(P3_U2674) );
  AOI21_X1 U20172 ( .B1(n16965), .B2(n16970), .A(n16964), .ZN(n17250) );
  NAND2_X1 U20173 ( .A1(n17226), .A2(n17250), .ZN(n16966) );
  OAI221_X1 U20174 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n16969), .C1(n16968), 
        .C2(n16967), .A(n16966), .ZN(P3_U2676) );
  AOI21_X1 U20175 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17220), .A(n16977), .ZN(
        n16973) );
  OAI21_X1 U20176 ( .B1(n16972), .B2(n16971), .A(n16970), .ZN(n17258) );
  OAI22_X1 U20177 ( .A1(n16974), .A2(n16973), .B1(n17220), .B2(n17258), .ZN(
        P3_U2677) );
  AOI21_X1 U20178 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17220), .A(n16983), .ZN(
        n16976) );
  XNOR2_X1 U20179 ( .A(n16975), .B(n16979), .ZN(n17263) );
  OAI22_X1 U20180 ( .A1(n16977), .A2(n16976), .B1(n17220), .B2(n17263), .ZN(
        P3_U2678) );
  AOI22_X1 U20181 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n17220), .B1(
        P3_EBX_REG_23__SCAN_IN), .B2(n16978), .ZN(n16982) );
  OAI21_X1 U20182 ( .B1(n16981), .B2(n16980), .A(n16979), .ZN(n17268) );
  OAI22_X1 U20183 ( .A1(n16983), .A2(n16982), .B1(n17220), .B2(n17268), .ZN(
        P3_U2679) );
  XNOR2_X1 U20184 ( .A(n16985), .B(n16984), .ZN(n17273) );
  NAND3_X1 U20185 ( .A1(n16987), .A2(P3_EBX_REG_23__SCAN_IN), .A3(n17220), 
        .ZN(n16986) );
  OAI221_X1 U20186 ( .B1(n16987), .B2(P3_EBX_REG_23__SCAN_IN), .C1(n17220), 
        .C2(n17273), .A(n16986), .ZN(P3_U2680) );
  AOI22_X1 U20187 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16991) );
  AOI22_X1 U20188 ( .A1(n17128), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16990) );
  AOI22_X1 U20189 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16989) );
  AOI22_X1 U20190 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16988) );
  NAND4_X1 U20191 ( .A1(n16991), .A2(n16990), .A3(n16989), .A4(n16988), .ZN(
        n16997) );
  AOI22_X1 U20192 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n9639), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n16995) );
  AOI22_X1 U20193 ( .A1(n9637), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16994) );
  AOI22_X1 U20194 ( .A1(n15584), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n16993) );
  AOI22_X1 U20195 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(n9641), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16992) );
  NAND4_X1 U20196 ( .A1(n16995), .A2(n16994), .A3(n16993), .A4(n16992), .ZN(
        n16996) );
  NOR2_X1 U20197 ( .A1(n16997), .A2(n16996), .ZN(n17275) );
  NAND3_X1 U20198 ( .A1(n16999), .A2(P3_EBX_REG_22__SCAN_IN), .A3(n17220), 
        .ZN(n16998) );
  OAI221_X1 U20199 ( .B1(n16999), .B2(P3_EBX_REG_22__SCAN_IN), .C1(n17220), 
        .C2(n17275), .A(n16998), .ZN(P3_U2681) );
  NAND2_X1 U20200 ( .A1(n17220), .A2(n17000), .ZN(n17029) );
  AOI22_X1 U20201 ( .A1(n17128), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n17011) );
  AOI22_X1 U20202 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n17010) );
  AOI22_X1 U20203 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n17001) );
  OAI21_X1 U20204 ( .B1(n17058), .B2(n17204), .A(n17001), .ZN(n17008) );
  AOI22_X1 U20205 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n17006) );
  AOI22_X1 U20206 ( .A1(n9637), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n9641), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n17005) );
  AOI22_X1 U20207 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n17004) );
  AOI22_X1 U20208 ( .A1(n9639), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n17003) );
  NAND4_X1 U20209 ( .A1(n17006), .A2(n17005), .A3(n17004), .A4(n17003), .ZN(
        n17007) );
  AOI211_X1 U20210 ( .C1(n17182), .C2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A(
        n17008), .B(n17007), .ZN(n17009) );
  NAND3_X1 U20211 ( .A1(n17011), .A2(n17010), .A3(n17009), .ZN(n17279) );
  AOI22_X1 U20212 ( .A1(n17226), .A2(n17279), .B1(n17012), .B2(n17014), .ZN(
        n17013) );
  OAI21_X1 U20213 ( .B1(n17014), .B2(n17029), .A(n17013), .ZN(P3_U2682) );
  AOI22_X1 U20214 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n17025) );
  AOI22_X1 U20215 ( .A1(n17128), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17024) );
  AOI22_X1 U20216 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17015) );
  OAI21_X1 U20217 ( .B1(n17058), .B2(n17208), .A(n17015), .ZN(n17022) );
  AOI22_X1 U20218 ( .A1(n9637), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n17020) );
  AOI22_X1 U20219 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17016), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17019) );
  AOI22_X1 U20220 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9639), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n17018) );
  AOI22_X1 U20221 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n17017) );
  NAND4_X1 U20222 ( .A1(n17020), .A2(n17019), .A3(n17018), .A4(n17017), .ZN(
        n17021) );
  AOI211_X1 U20223 ( .C1(n9640), .C2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n17022), .B(n17021), .ZN(n17023) );
  NAND3_X1 U20224 ( .A1(n17025), .A2(n17024), .A3(n17023), .ZN(n17286) );
  NAND2_X1 U20225 ( .A1(n17226), .A2(n17286), .ZN(n17026) );
  OAI221_X1 U20226 ( .B1(n17029), .B2(n17028), .C1(n17029), .C2(n17027), .A(
        n17026), .ZN(P3_U2683) );
  AOI21_X1 U20227 ( .B1(n17030), .B2(n17053), .A(n17226), .ZN(n17031) );
  INV_X1 U20228 ( .A(n17031), .ZN(n17042) );
  AOI22_X1 U20229 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n17035) );
  AOI22_X1 U20230 ( .A1(n9637), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17034) );
  AOI22_X1 U20231 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17033) );
  AOI22_X1 U20232 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17032) );
  NAND4_X1 U20233 ( .A1(n17035), .A2(n17034), .A3(n17033), .A4(n17032), .ZN(
        n17041) );
  AOI22_X1 U20234 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n13903), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17039) );
  AOI22_X1 U20235 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n9639), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n17038) );
  AOI22_X1 U20236 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17037) );
  AOI22_X1 U20237 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17128), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n17036) );
  NAND4_X1 U20238 ( .A1(n17039), .A2(n17038), .A3(n17037), .A4(n17036), .ZN(
        n17040) );
  NOR2_X1 U20239 ( .A1(n17041), .A2(n17040), .ZN(n17292) );
  OAI22_X1 U20240 ( .A1(n9700), .A2(n17042), .B1(n17292), .B2(n17220), .ZN(
        P3_U2684) );
  AOI22_X1 U20241 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17046) );
  AOI22_X1 U20242 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17045) );
  AOI22_X1 U20243 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(n9637), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17044) );
  AOI22_X1 U20244 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17043) );
  NAND4_X1 U20245 ( .A1(n17046), .A2(n17045), .A3(n17044), .A4(n17043), .ZN(
        n17052) );
  AOI22_X1 U20246 ( .A1(n17144), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n17050) );
  AOI22_X1 U20247 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n9634), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n17049) );
  AOI22_X1 U20248 ( .A1(n17128), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17048) );
  AOI22_X1 U20249 ( .A1(n9639), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17047) );
  NAND4_X1 U20250 ( .A1(n17050), .A2(n17049), .A3(n17048), .A4(n17047), .ZN(
        n17051) );
  NOR2_X1 U20251 ( .A1(n17052), .A2(n17051), .ZN(n17297) );
  OAI21_X1 U20252 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n17054), .A(n17053), .ZN(
        n17055) );
  AOI22_X1 U20253 ( .A1(n17226), .A2(n17297), .B1(n17055), .B2(n17220), .ZN(
        P3_U2685) );
  AOI22_X1 U20254 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_13__1__SCAN_IN), .B2(n17164), .ZN(n17067) );
  AOI22_X1 U20255 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n17180), .ZN(n17066) );
  AOI22_X1 U20256 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n17181), .ZN(n17057) );
  OAI21_X1 U20257 ( .B1(n17221), .B2(n17058), .A(n17057), .ZN(n17064) );
  AOI22_X1 U20258 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n9634), .B1(n9637), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17062) );
  AOI22_X1 U20259 ( .A1(n17157), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17061) );
  AOI22_X1 U20260 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n9641), .B1(
        P3_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n9639), .ZN(n17060) );
  AOI22_X1 U20261 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17159), .ZN(n17059) );
  NAND4_X1 U20262 ( .A1(n17062), .A2(n17061), .A3(n17060), .A4(n17059), .ZN(
        n17063) );
  AOI211_X1 U20263 ( .C1(n17182), .C2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A(
        n17064), .B(n17063), .ZN(n17065) );
  NAND3_X1 U20264 ( .A1(n17067), .A2(n17066), .A3(n17065), .ZN(n17298) );
  INV_X1 U20265 ( .A(n17070), .ZN(n17068) );
  OAI33_X1 U20266 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n18233), .A3(n17070), 
        .B1(n17069), .B2(n17226), .B3(n17068), .ZN(n17071) );
  AOI21_X1 U20267 ( .B1(n17226), .B2(n17298), .A(n17071), .ZN(n17072) );
  INV_X1 U20268 ( .A(n17072), .ZN(P3_U2686) );
  NAND2_X1 U20269 ( .A1(n17074), .A2(n17073), .ZN(n17097) );
  AOI22_X1 U20270 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9639), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n17079) );
  AOI22_X1 U20271 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n17075), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17078) );
  AOI22_X1 U20272 ( .A1(n9637), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(n9635), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n17077) );
  AOI22_X1 U20273 ( .A1(n17128), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17076) );
  NAND4_X1 U20274 ( .A1(n17079), .A2(n17078), .A3(n17077), .A4(n17076), .ZN(
        n17085) );
  AOI22_X1 U20275 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n13903), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17083) );
  AOI22_X1 U20276 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17082) );
  AOI22_X1 U20277 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17081) );
  AOI22_X1 U20278 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17080) );
  NAND4_X1 U20279 ( .A1(n17083), .A2(n17082), .A3(n17081), .A4(n17080), .ZN(
        n17084) );
  NOR2_X1 U20280 ( .A1(n17085), .A2(n17084), .ZN(n17310) );
  NAND3_X1 U20281 ( .A1(n17097), .A2(P3_EBX_REG_16__SCAN_IN), .A3(n17220), 
        .ZN(n17086) );
  OAI221_X1 U20282 ( .B1(n17097), .B2(P3_EBX_REG_16__SCAN_IN), .C1(n17220), 
        .C2(n17310), .A(n17086), .ZN(P3_U2687) );
  AOI22_X1 U20283 ( .A1(n17128), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9639), .B2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n17090) );
  AOI22_X1 U20284 ( .A1(n9637), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n17089) );
  AOI22_X1 U20285 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n17088) );
  AOI22_X1 U20286 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n9641), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n17087) );
  NAND4_X1 U20287 ( .A1(n17090), .A2(n17089), .A3(n17088), .A4(n17087), .ZN(
        n17096) );
  AOI22_X1 U20288 ( .A1(n15584), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n17094) );
  AOI22_X1 U20289 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n13903), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n17093) );
  AOI22_X1 U20290 ( .A1(n17174), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n17092) );
  AOI22_X1 U20291 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n17091) );
  NAND4_X1 U20292 ( .A1(n17094), .A2(n17093), .A3(n17092), .A4(n17091), .ZN(
        n17095) );
  NOR2_X1 U20293 ( .A1(n17096), .A2(n17095), .ZN(n17314) );
  INV_X1 U20294 ( .A(n17110), .ZN(n17098) );
  OAI211_X1 U20295 ( .C1(P3_EBX_REG_15__SCAN_IN), .C2(n17098), .A(n17097), .B(
        n17220), .ZN(n17099) );
  OAI21_X1 U20296 ( .B1(n17314), .B2(n17220), .A(n17099), .ZN(P3_U2688) );
  AOI22_X1 U20297 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n9639), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n17109) );
  AOI22_X1 U20298 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n17108) );
  AOI22_X1 U20299 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(n9641), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n17100) );
  OAI21_X1 U20300 ( .B1(n15538), .B2(n20948), .A(n17100), .ZN(n17106) );
  AOI22_X1 U20301 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9637), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n17104) );
  AOI22_X1 U20302 ( .A1(n15584), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n17103) );
  AOI22_X1 U20303 ( .A1(n17128), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n17102) );
  AOI22_X1 U20304 ( .A1(n17180), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17101) );
  NAND4_X1 U20305 ( .A1(n17104), .A2(n17103), .A3(n17102), .A4(n17101), .ZN(
        n17105) );
  AOI211_X1 U20306 ( .C1(n9640), .C2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A(
        n17106), .B(n17105), .ZN(n17107) );
  NAND3_X1 U20307 ( .A1(n17109), .A2(n17108), .A3(n17107), .ZN(n17318) );
  INV_X1 U20308 ( .A(n17318), .ZN(n17113) );
  OAI21_X1 U20309 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17111), .A(n17110), .ZN(
        n17112) );
  AOI22_X1 U20310 ( .A1(n17226), .A2(n17113), .B1(n17112), .B2(n17220), .ZN(
        P3_U2689) );
  AOI22_X1 U20311 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n15584), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17117) );
  AOI22_X1 U20312 ( .A1(n9637), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17116) );
  AOI22_X1 U20313 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(n9639), .B2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n17115) );
  AOI22_X1 U20314 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17114) );
  NAND4_X1 U20315 ( .A1(n17117), .A2(n17116), .A3(n17115), .A4(n17114), .ZN(
        n17123) );
  AOI22_X1 U20316 ( .A1(n17128), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9635), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n17121) );
  AOI22_X1 U20317 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n17120) );
  AOI22_X1 U20318 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17119) );
  AOI22_X1 U20319 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17118) );
  NAND4_X1 U20320 ( .A1(n17121), .A2(n17120), .A3(n17119), .A4(n17118), .ZN(
        n17122) );
  NOR2_X1 U20321 ( .A1(n17123), .A2(n17122), .ZN(n17327) );
  OAI21_X1 U20322 ( .B1(P3_EBX_REG_12__SCAN_IN), .B2(n9722), .A(n17124), .ZN(
        n17125) );
  AOI22_X1 U20323 ( .A1(n17226), .A2(n17327), .B1(n17125), .B2(n17220), .ZN(
        P3_U2691) );
  AOI21_X1 U20324 ( .B1(n17126), .B2(n17152), .A(n17226), .ZN(n17127) );
  INV_X1 U20325 ( .A(n17127), .ZN(n17139) );
  AOI22_X1 U20326 ( .A1(n17128), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17132) );
  AOI22_X1 U20327 ( .A1(n9637), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(n9634), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n17131) );
  AOI22_X1 U20328 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17130) );
  AOI22_X1 U20329 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17129) );
  NAND4_X1 U20330 ( .A1(n17132), .A2(n17131), .A3(n17130), .A4(n17129), .ZN(
        n17138) );
  AOI22_X1 U20331 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n17136) );
  AOI22_X1 U20332 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17135) );
  AOI22_X1 U20333 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n17134) );
  AOI22_X1 U20334 ( .A1(n15584), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9639), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n17133) );
  NAND4_X1 U20335 ( .A1(n17136), .A2(n17135), .A3(n17134), .A4(n17133), .ZN(
        n17137) );
  NOR2_X1 U20336 ( .A1(n17138), .A2(n17137), .ZN(n17331) );
  OAI22_X1 U20337 ( .A1(n9722), .A2(n17139), .B1(n17331), .B2(n17220), .ZN(
        P3_U2692) );
  AOI22_X1 U20338 ( .A1(n9641), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9639), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n17143) );
  AOI22_X1 U20339 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n17142) );
  AOI22_X1 U20340 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n17128), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n17141) );
  AOI22_X1 U20341 ( .A1(n17181), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17159), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17140) );
  NAND4_X1 U20342 ( .A1(n17143), .A2(n17142), .A3(n17141), .A4(n17140), .ZN(
        n17151) );
  AOI22_X1 U20343 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17149) );
  AOI22_X1 U20344 ( .A1(n9637), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n17148) );
  AOI22_X1 U20345 ( .A1(n17145), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n17147) );
  AOI22_X1 U20346 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n17146) );
  NAND4_X1 U20347 ( .A1(n17149), .A2(n17148), .A3(n17147), .A4(n17146), .ZN(
        n17150) );
  NOR2_X1 U20348 ( .A1(n17151), .A2(n17150), .ZN(n17338) );
  OAI21_X1 U20349 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17172), .A(n17152), .ZN(
        n17153) );
  AOI22_X1 U20350 ( .A1(n17226), .A2(n17338), .B1(n17153), .B2(n17220), .ZN(
        P3_U2693) );
  AOI21_X1 U20351 ( .B1(n17155), .B2(n17154), .A(n17226), .ZN(n17156) );
  INV_X1 U20352 ( .A(n17156), .ZN(n17171) );
  AOI22_X1 U20353 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9640), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n17163) );
  AOI22_X1 U20354 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n17157), .B1(
        P3_INSTQUEUE_REG_8__1__SCAN_IN), .B2(n9639), .ZN(n17162) );
  AOI22_X1 U20355 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n9635), .B1(
        n17144), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n17161) );
  AOI22_X1 U20356 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17159), .B1(
        n17158), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n17160) );
  NAND4_X1 U20357 ( .A1(n17163), .A2(n17162), .A3(n17161), .A4(n17160), .ZN(
        n17170) );
  AOI22_X1 U20358 ( .A1(n15584), .A2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_11__1__SCAN_IN), .B2(n9641), .ZN(n17168) );
  AOI22_X1 U20359 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17181), .ZN(n17167) );
  AOI22_X1 U20360 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n17164), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n17180), .ZN(n17166) );
  AOI22_X1 U20361 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n9637), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17165) );
  NAND4_X1 U20362 ( .A1(n17168), .A2(n17167), .A3(n17166), .A4(n17165), .ZN(
        n17169) );
  NOR2_X1 U20363 ( .A1(n17170), .A2(n17169), .ZN(n17341) );
  OAI22_X1 U20364 ( .A1(n17172), .A2(n17171), .B1(n17341), .B2(n17220), .ZN(
        P3_U2694) );
  AOI22_X1 U20365 ( .A1(n17173), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9639), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n17179) );
  AOI22_X1 U20366 ( .A1(n9637), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n17164), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17178) );
  AOI22_X1 U20367 ( .A1(n9640), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17174), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n17177) );
  AOI22_X1 U20368 ( .A1(n17158), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17175), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17176) );
  NAND4_X1 U20369 ( .A1(n17179), .A2(n17178), .A3(n17177), .A4(n17176), .ZN(
        n17188) );
  AOI22_X1 U20370 ( .A1(n17002), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9641), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n17186) );
  AOI22_X1 U20371 ( .A1(n17075), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n17180), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17185) );
  AOI22_X1 U20372 ( .A1(n9635), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17181), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17184) );
  AOI22_X1 U20373 ( .A1(n17182), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n17128), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n17183) );
  NAND4_X1 U20374 ( .A1(n17186), .A2(n17185), .A3(n17184), .A4(n17183), .ZN(
        n17187) );
  NOR2_X1 U20375 ( .A1(n17188), .A2(n17187), .ZN(n17348) );
  NOR2_X1 U20376 ( .A1(n17226), .A2(n17190), .ZN(n17195) );
  NOR2_X1 U20377 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n18233), .ZN(n17189) );
  AOI22_X1 U20378 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17195), .B1(n17190), .B2(
        n17189), .ZN(n17191) );
  OAI21_X1 U20379 ( .B1(n17348), .B2(n17220), .A(n17191), .ZN(P3_U2695) );
  NOR2_X1 U20380 ( .A1(n17192), .A2(n17228), .ZN(n17210) );
  INV_X1 U20381 ( .A(n17210), .ZN(n17198) );
  NOR3_X1 U20382 ( .A1(n17193), .A2(n17199), .A3(n17198), .ZN(n17202) );
  AOI22_X1 U20383 ( .A1(P3_EBX_REG_7__SCAN_IN), .A2(n17195), .B1(n17202), .B2(
        n17194), .ZN(n17196) );
  OAI21_X1 U20384 ( .B1(n17197), .B2(n17220), .A(n17196), .ZN(P3_U2696) );
  NOR2_X1 U20385 ( .A1(n17199), .A2(n17198), .ZN(n17206) );
  AOI21_X1 U20386 ( .B1(P3_EBX_REG_6__SCAN_IN), .B2(n17220), .A(n17206), .ZN(
        n17201) );
  INV_X1 U20387 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n17200) );
  OAI22_X1 U20388 ( .A1(n17202), .A2(n17201), .B1(n17200), .B2(n17220), .ZN(
        P3_U2697) );
  OAI21_X1 U20389 ( .B1(P3_EBX_REG_5__SCAN_IN), .B2(n17203), .A(n17220), .ZN(
        n17205) );
  OAI22_X1 U20390 ( .A1(n17206), .A2(n17205), .B1(n17204), .B2(n17220), .ZN(
        P3_U2698) );
  NOR3_X1 U20391 ( .A1(n17207), .A2(n17211), .A3(n17228), .ZN(n17214) );
  AOI21_X1 U20392 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17220), .A(n17214), .ZN(
        n17209) );
  OAI22_X1 U20393 ( .A1(n17210), .A2(n17209), .B1(n17208), .B2(n17220), .ZN(
        P3_U2699) );
  NOR2_X1 U20394 ( .A1(n17211), .A2(n17228), .ZN(n17217) );
  AOI21_X1 U20395 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17220), .A(n17217), .ZN(
        n17213) );
  OAI22_X1 U20396 ( .A1(n17214), .A2(n17213), .B1(n17212), .B2(n17220), .ZN(
        P3_U2700) );
  INV_X1 U20397 ( .A(n17215), .ZN(n17216) );
  AOI21_X1 U20398 ( .B1(n17222), .B2(n17216), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n17219) );
  INV_X1 U20399 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17218) );
  AOI221_X1 U20400 ( .B1(n17219), .B2(n17220), .C1(n17218), .C2(n17226), .A(
        n17217), .ZN(P3_U2701) );
  OAI222_X1 U20401 ( .A1(n17224), .A2(n17228), .B1(n17223), .B2(n17222), .C1(
        n17221), .C2(n17220), .ZN(P3_U2702) );
  AOI22_X1 U20402 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n17226), .B1(
        P3_EBX_REG_0__SCAN_IN), .B2(n17225), .ZN(n17227) );
  OAI21_X1 U20403 ( .B1(P3_EBX_REG_0__SCAN_IN), .B2(n17228), .A(n17227), .ZN(
        P3_U2703) );
  INV_X1 U20404 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17450) );
  INV_X1 U20405 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17446) );
  INV_X1 U20406 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17489) );
  NAND2_X1 U20407 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n9654), .ZN(n17379) );
  NAND3_X1 U20408 ( .A1(P3_EAX_REG_7__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_0__SCAN_IN), .ZN(n17231) );
  NAND4_X1 U20409 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_4__SCAN_IN), 
        .A3(P3_EAX_REG_3__SCAN_IN), .A4(P3_EAX_REG_2__SCAN_IN), .ZN(n17230) );
  NOR3_X2 U20410 ( .A1(n17379), .A2(n17231), .A3(n17230), .ZN(n17311) );
  INV_X1 U20411 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n17472) );
  INV_X1 U20412 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n20778) );
  INV_X1 U20413 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17484) );
  NAND4_X1 U20414 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(P3_EAX_REG_12__SCAN_IN), 
        .A3(P3_EAX_REG_11__SCAN_IN), .A4(P3_EAX_REG_10__SCAN_IN), .ZN(n17232)
         );
  NOR4_X1 U20415 ( .A1(n17472), .A2(n20778), .A3(n17484), .A4(n17232), .ZN(
        n17312) );
  NAND2_X1 U20416 ( .A1(n17311), .A2(n17312), .ZN(n17313) );
  NAND3_X1 U20417 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(P3_EAX_REG_18__SCAN_IN), 
        .A3(P3_EAX_REG_17__SCAN_IN), .ZN(n17274) );
  NAND3_X1 U20418 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(P3_EAX_REG_22__SCAN_IN), 
        .A3(P3_EAX_REG_21__SCAN_IN), .ZN(n17233) );
  NAND2_X1 U20419 ( .A1(P3_EAX_REG_23__SCAN_IN), .A2(n17270), .ZN(n17269) );
  NAND2_X1 U20420 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17265), .ZN(n17264) );
  NOR2_X2 U20421 ( .A1(n17446), .A2(n17259), .ZN(n17254) );
  NAND2_X1 U20422 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(n17246), .ZN(n17242) );
  NAND2_X1 U20423 ( .A1(n17237), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17236) );
  NAND2_X1 U20424 ( .A1(n18228), .A2(n17368), .ZN(n17303) );
  OAI22_X1 U20425 ( .A1(P3_EAX_REG_30__SCAN_IN), .A2(n17378), .B1(n17368), 
        .B2(n17237), .ZN(n17234) );
  AOI22_X1 U20426 ( .A1(BUF2_REG_31__SCAN_IN), .A2(n17304), .B1(
        P3_EAX_REG_31__SCAN_IN), .B2(n17234), .ZN(n17235) );
  OAI21_X1 U20427 ( .B1(P3_EAX_REG_31__SCAN_IN), .B2(n17236), .A(n17235), .ZN(
        P3_U2704) );
  NOR2_X2 U20428 ( .A1(n18223), .A2(n17363), .ZN(n17305) );
  AOI22_X1 U20429 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17305), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n17304), .ZN(n17239) );
  OAI211_X1 U20430 ( .C1(n17237), .C2(P3_EAX_REG_30__SCAN_IN), .A(n17363), .B(
        n17236), .ZN(n17238) );
  OAI211_X1 U20431 ( .C1(n17240), .C2(n17371), .A(n17239), .B(n17238), .ZN(
        P3_U2705) );
  INV_X1 U20432 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n18225) );
  AOI22_X1 U20433 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17305), .B1(n17241), .B2(
        n17376), .ZN(n17244) );
  OAI211_X1 U20434 ( .C1(n17246), .C2(P3_EAX_REG_29__SCAN_IN), .A(n17363), .B(
        n17242), .ZN(n17243) );
  OAI211_X1 U20435 ( .C1(n17303), .C2(n18225), .A(n17244), .B(n17243), .ZN(
        P3_U2706) );
  INV_X1 U20436 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n18219) );
  AOI22_X1 U20437 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17305), .B1(n17245), .B2(
        n17376), .ZN(n17249) );
  AOI211_X1 U20438 ( .C1(n17450), .C2(n17251), .A(n17246), .B(n17368), .ZN(
        n17247) );
  INV_X1 U20439 ( .A(n17247), .ZN(n17248) );
  OAI211_X1 U20440 ( .C1(n17303), .C2(n18219), .A(n17249), .B(n17248), .ZN(
        P3_U2707) );
  INV_X1 U20441 ( .A(BUF2_REG_27__SCAN_IN), .ZN(n18215) );
  AOI22_X1 U20442 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17305), .B1(n17250), .B2(
        n17376), .ZN(n17253) );
  OAI211_X1 U20443 ( .C1(n17254), .C2(P3_EAX_REG_27__SCAN_IN), .A(n17363), .B(
        n17251), .ZN(n17252) );
  OAI211_X1 U20444 ( .C1(n17303), .C2(n18215), .A(n17253), .B(n17252), .ZN(
        P3_U2708) );
  AOI22_X1 U20445 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17305), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17304), .ZN(n17257) );
  AOI211_X1 U20446 ( .C1(n17446), .C2(n17259), .A(n17254), .B(n17368), .ZN(
        n17255) );
  INV_X1 U20447 ( .A(n17255), .ZN(n17256) );
  OAI211_X1 U20448 ( .C1(n17371), .C2(n17258), .A(n17257), .B(n17256), .ZN(
        P3_U2709) );
  AOI22_X1 U20449 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17305), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n17304), .ZN(n17262) );
  OAI211_X1 U20450 ( .C1(n17260), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17363), .B(
        n17259), .ZN(n17261) );
  OAI211_X1 U20451 ( .C1(n17371), .C2(n17263), .A(n17262), .B(n17261), .ZN(
        P3_U2710) );
  AOI22_X1 U20452 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17305), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17304), .ZN(n17267) );
  OAI211_X1 U20453 ( .C1(n17265), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17363), .B(
        n17264), .ZN(n17266) );
  OAI211_X1 U20454 ( .C1(n17371), .C2(n17268), .A(n17267), .B(n17266), .ZN(
        P3_U2711) );
  AOI22_X1 U20455 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17305), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n17304), .ZN(n17272) );
  OAI211_X1 U20456 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17270), .A(n17363), .B(
        n17269), .ZN(n17271) );
  OAI211_X1 U20457 ( .C1(n17371), .C2(n17273), .A(n17272), .B(n17271), .ZN(
        P3_U2712) );
  INV_X1 U20458 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17434) );
  OR3_X1 U20459 ( .A1(n18233), .A2(n17306), .A3(n17274), .ZN(n17289) );
  NAND2_X1 U20460 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17283), .ZN(n17280) );
  NAND2_X1 U20461 ( .A1(n17280), .A2(P3_EAX_REG_22__SCAN_IN), .ZN(n17278) );
  INV_X1 U20462 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n19243) );
  OAI22_X1 U20463 ( .A1(n17275), .A2(n17371), .B1(n19243), .B2(n17303), .ZN(
        n17276) );
  AOI21_X1 U20464 ( .B1(BUF2_REG_6__SCAN_IN), .B2(n17305), .A(n17276), .ZN(
        n17277) );
  OAI221_X1 U20465 ( .B1(n17280), .B2(P3_EAX_REG_22__SCAN_IN), .C1(n17278), 
        .C2(n17368), .A(n17277), .ZN(P3_U2713) );
  INV_X1 U20466 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n19237) );
  AOI22_X1 U20467 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17305), .B1(n17376), .B2(
        n17279), .ZN(n17282) );
  OAI211_X1 U20468 ( .C1(n17283), .C2(P3_EAX_REG_21__SCAN_IN), .A(n17363), .B(
        n17280), .ZN(n17281) );
  OAI211_X1 U20469 ( .C1(n17303), .C2(n19237), .A(n17282), .B(n17281), .ZN(
        P3_U2714) );
  INV_X1 U20470 ( .A(n17283), .ZN(n17285) );
  OAI21_X1 U20471 ( .B1(n17368), .B2(n17434), .A(n17289), .ZN(n17284) );
  AOI22_X1 U20472 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n17304), .B1(n17285), .B2(
        n17284), .ZN(n17288) );
  AOI22_X1 U20473 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17305), .B1(n17376), .B2(
        n17286), .ZN(n17287) );
  NAND2_X1 U20474 ( .A1(n17288), .A2(n17287), .ZN(P3_U2715) );
  AOI22_X1 U20475 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17305), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17304), .ZN(n17291) );
  INV_X1 U20476 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17430) );
  INV_X1 U20477 ( .A(n17306), .ZN(n17300) );
  NAND2_X1 U20478 ( .A1(P3_EAX_REG_17__SCAN_IN), .A2(n17300), .ZN(n17299) );
  NOR2_X1 U20479 ( .A1(n17430), .A2(n17299), .ZN(n17293) );
  OAI211_X1 U20480 ( .C1(n17293), .C2(P3_EAX_REG_19__SCAN_IN), .A(n17363), .B(
        n17289), .ZN(n17290) );
  OAI211_X1 U20481 ( .C1(n17292), .C2(n17371), .A(n17291), .B(n17290), .ZN(
        P3_U2716) );
  AOI22_X1 U20482 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17305), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17304), .ZN(n17296) );
  AOI211_X1 U20483 ( .C1(n17430), .C2(n17299), .A(n17293), .B(n17368), .ZN(
        n17294) );
  INV_X1 U20484 ( .A(n17294), .ZN(n17295) );
  OAI211_X1 U20485 ( .C1(n17297), .C2(n17371), .A(n17296), .B(n17295), .ZN(
        P3_U2717) );
  INV_X1 U20486 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n19221) );
  AOI22_X1 U20487 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17305), .B1(n17376), .B2(
        n17298), .ZN(n17302) );
  OAI211_X1 U20488 ( .C1(n17300), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17363), .B(
        n17299), .ZN(n17301) );
  OAI211_X1 U20489 ( .C1(n17303), .C2(n19221), .A(n17302), .B(n17301), .ZN(
        P3_U2718) );
  AOI22_X1 U20490 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17305), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17304), .ZN(n17309) );
  OAI211_X1 U20491 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17307), .A(n17363), .B(
        n17306), .ZN(n17308) );
  OAI211_X1 U20492 ( .C1(n17310), .C2(n17371), .A(n17309), .B(n17308), .ZN(
        P3_U2719) );
  INV_X1 U20493 ( .A(n17311), .ZN(n17345) );
  NOR2_X1 U20494 ( .A1(n18233), .A2(n17345), .ZN(n17351) );
  NAND2_X1 U20495 ( .A1(n17312), .A2(n17351), .ZN(n17317) );
  NAND2_X1 U20496 ( .A1(n17363), .A2(n17313), .ZN(n17320) );
  INV_X1 U20497 ( .A(n17314), .ZN(n17315) );
  AOI22_X1 U20498 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17377), .B1(n17376), .B2(
        n17315), .ZN(n17316) );
  OAI221_X1 U20499 ( .B1(P3_EAX_REG_15__SCAN_IN), .B2(n17317), .C1(n17489), 
        .C2(n17320), .A(n17316), .ZN(P3_U2720) );
  INV_X1 U20500 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n17479) );
  INV_X1 U20501 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17474) );
  NAND2_X1 U20502 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17340), .ZN(n17339) );
  NAND2_X1 U20503 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(n17335), .ZN(n17326) );
  NOR2_X1 U20504 ( .A1(n17479), .A2(n17326), .ZN(n17329) );
  NAND2_X1 U20505 ( .A1(P3_EAX_REG_13__SCAN_IN), .A2(n17329), .ZN(n17321) );
  AOI22_X1 U20506 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17377), .B1(n17376), .B2(
        n17318), .ZN(n17319) );
  OAI221_X1 U20507 ( .B1(P3_EAX_REG_14__SCAN_IN), .B2(n17321), .C1(n17484), 
        .C2(n17320), .A(n17319), .ZN(P3_U2721) );
  INV_X1 U20508 ( .A(n17321), .ZN(n17324) );
  AOI21_X1 U20509 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17363), .A(n17329), .ZN(
        n17323) );
  OAI222_X1 U20510 ( .A1(n17374), .A2(n17325), .B1(n17324), .B2(n17323), .C1(
        n17371), .C2(n17322), .ZN(P3_U2722) );
  INV_X1 U20511 ( .A(n17326), .ZN(n17333) );
  AOI21_X1 U20512 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17363), .A(n17333), .ZN(
        n17328) );
  OAI222_X1 U20513 ( .A1(n17374), .A2(n17330), .B1(n17329), .B2(n17328), .C1(
        n17371), .C2(n17327), .ZN(P3_U2723) );
  AOI21_X1 U20514 ( .B1(P3_EAX_REG_11__SCAN_IN), .B2(n17363), .A(n17335), .ZN(
        n17332) );
  OAI222_X1 U20515 ( .A1(n17374), .A2(n17334), .B1(n17333), .B2(n17332), .C1(
        n17371), .C2(n17331), .ZN(P3_U2724) );
  AOI211_X1 U20516 ( .C1(n17474), .C2(n17339), .A(n17368), .B(n17335), .ZN(
        n17336) );
  AOI21_X1 U20517 ( .B1(n17377), .B2(BUF2_REG_10__SCAN_IN), .A(n17336), .ZN(
        n17337) );
  OAI21_X1 U20518 ( .B1(n17338), .B2(n17371), .A(n17337), .ZN(P3_U2725) );
  INV_X1 U20519 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17344) );
  INV_X1 U20520 ( .A(n17339), .ZN(n17343) );
  AOI21_X1 U20521 ( .B1(P3_EAX_REG_9__SCAN_IN), .B2(n17363), .A(n17340), .ZN(
        n17342) );
  OAI222_X1 U20522 ( .A1(n17374), .A2(n17344), .B1(n17343), .B2(n17342), .C1(
        n17371), .C2(n17341), .ZN(P3_U2726) );
  AOI22_X1 U20523 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17377), .B1(n17351), .B2(
        n20778), .ZN(n17347) );
  NAND3_X1 U20524 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17363), .A3(n17345), .ZN(
        n17346) );
  OAI211_X1 U20525 ( .C1(n17348), .C2(n17371), .A(n17347), .B(n17346), .ZN(
        P3_U2727) );
  INV_X1 U20526 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n17467) );
  INV_X1 U20527 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17463) );
  INV_X1 U20528 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17459) );
  NOR2_X1 U20529 ( .A1(n17455), .A2(n17378), .ZN(n17381) );
  NAND2_X1 U20530 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17381), .ZN(n17367) );
  NOR2_X1 U20531 ( .A1(n17459), .A2(n17367), .ZN(n17373) );
  NAND2_X1 U20532 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17373), .ZN(n17359) );
  NOR2_X1 U20533 ( .A1(n17463), .A2(n17359), .ZN(n17362) );
  NAND2_X1 U20534 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17362), .ZN(n17352) );
  NOR2_X1 U20535 ( .A1(n17467), .A2(n17352), .ZN(n17355) );
  AOI21_X1 U20536 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17363), .A(n17355), .ZN(
        n17350) );
  OAI222_X1 U20537 ( .A1(n17374), .A2(n18235), .B1(n17351), .B2(n17350), .C1(
        n17371), .C2(n17349), .ZN(P3_U2728) );
  INV_X1 U20538 ( .A(n17352), .ZN(n17358) );
  AOI21_X1 U20539 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17363), .A(n17358), .ZN(
        n17354) );
  OAI222_X1 U20540 ( .A1(n18230), .A2(n17374), .B1(n17355), .B2(n17354), .C1(
        n17371), .C2(n17353), .ZN(P3_U2729) );
  INV_X1 U20541 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18224) );
  AOI21_X1 U20542 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17363), .A(n17362), .ZN(
        n17357) );
  OAI222_X1 U20543 ( .A1(n18224), .A2(n17374), .B1(n17358), .B2(n17357), .C1(
        n17371), .C2(n17356), .ZN(P3_U2730) );
  INV_X1 U20544 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18220) );
  INV_X1 U20545 ( .A(n17359), .ZN(n17366) );
  AOI21_X1 U20546 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17363), .A(n17366), .ZN(
        n17361) );
  OAI222_X1 U20547 ( .A1(n18220), .A2(n17374), .B1(n17362), .B2(n17361), .C1(
        n17371), .C2(n17360), .ZN(P3_U2731) );
  AOI21_X1 U20548 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17363), .A(n17373), .ZN(
        n17365) );
  OAI222_X1 U20549 ( .A1(n18214), .A2(n17374), .B1(n17366), .B2(n17365), .C1(
        n17371), .C2(n17364), .ZN(P3_U2732) );
  INV_X1 U20550 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18209) );
  OAI21_X1 U20551 ( .B1(n17459), .B2(n17368), .A(n17367), .ZN(n17369) );
  INV_X1 U20552 ( .A(n17369), .ZN(n17372) );
  OAI222_X1 U20553 ( .A1(n18209), .A2(n17374), .B1(n17373), .B2(n17372), .C1(
        n17371), .C2(n17370), .ZN(P3_U2733) );
  AOI22_X1 U20554 ( .A1(n17377), .A2(BUF2_REG_1__SCAN_IN), .B1(n17376), .B2(
        n17375), .ZN(n17383) );
  NOR2_X1 U20555 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17378), .ZN(n17380) );
  OAI22_X1 U20556 ( .A1(P3_EAX_REG_1__SCAN_IN), .A2(n17381), .B1(n17380), .B2(
        n17379), .ZN(n17382) );
  NAND2_X1 U20557 ( .A1(n17383), .A2(n17382), .ZN(P3_U2734) );
  OR2_X1 U20558 ( .A1(n18792), .A2(n18696), .ZN(n18828) );
  AND2_X1 U20560 ( .A1(n17412), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  INV_X1 U20561 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17453) );
  NAND2_X1 U20562 ( .A1(n17402), .A2(n18196), .ZN(n17401) );
  AOI22_X1 U20563 ( .A1(n18679), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(n17419), 
        .B2(P3_DATAO_REG_30__SCAN_IN), .ZN(n17386) );
  OAI21_X1 U20564 ( .B1(n17453), .B2(n17401), .A(n17386), .ZN(P3_U2737) );
  INV_X1 U20565 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n20935) );
  AOI22_X1 U20566 ( .A1(n18679), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17419), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17387) );
  OAI21_X1 U20567 ( .B1(n20935), .B2(n17401), .A(n17387), .ZN(P3_U2738) );
  AOI22_X1 U20568 ( .A1(n18679), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17419), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17388) );
  OAI21_X1 U20569 ( .B1(n17450), .B2(n17401), .A(n17388), .ZN(P3_U2739) );
  INV_X1 U20570 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17448) );
  AOI22_X1 U20571 ( .A1(n18679), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17412), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17389) );
  OAI21_X1 U20572 ( .B1(n17448), .B2(n17401), .A(n17389), .ZN(P3_U2740) );
  AOI22_X1 U20573 ( .A1(n18679), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17412), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17390) );
  OAI21_X1 U20574 ( .B1(n17446), .B2(n17401), .A(n17390), .ZN(P3_U2741) );
  INV_X1 U20575 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17444) );
  AOI22_X1 U20576 ( .A1(n18679), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17412), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17391) );
  OAI21_X1 U20577 ( .B1(n17444), .B2(n17401), .A(n17391), .ZN(P3_U2742) );
  INV_X1 U20578 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17442) );
  AOI22_X1 U20579 ( .A1(n18679), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17412), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17392) );
  OAI21_X1 U20580 ( .B1(n17442), .B2(n17401), .A(n17392), .ZN(P3_U2743) );
  INV_X1 U20581 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17440) );
  AOI22_X1 U20583 ( .A1(n18679), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17419), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17393) );
  OAI21_X1 U20584 ( .B1(n17440), .B2(n17401), .A(n17393), .ZN(P3_U2744) );
  INV_X1 U20585 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17438) );
  AOI22_X1 U20586 ( .A1(n18679), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17419), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17394) );
  OAI21_X1 U20587 ( .B1(n17438), .B2(n17401), .A(n17394), .ZN(P3_U2745) );
  INV_X1 U20588 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17436) );
  AOI22_X1 U20589 ( .A1(n18679), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17419), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17395) );
  OAI21_X1 U20590 ( .B1(n17436), .B2(n17401), .A(n17395), .ZN(P3_U2746) );
  AOI22_X1 U20591 ( .A1(n18679), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17419), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17396) );
  OAI21_X1 U20592 ( .B1(n17434), .B2(n17401), .A(n17396), .ZN(P3_U2747) );
  INV_X1 U20593 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17432) );
  AOI22_X1 U20594 ( .A1(n18679), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17419), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17397) );
  OAI21_X1 U20595 ( .B1(n17432), .B2(n17401), .A(n17397), .ZN(P3_U2748) );
  AOI22_X1 U20596 ( .A1(n18679), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17419), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17398) );
  OAI21_X1 U20597 ( .B1(n17430), .B2(n17401), .A(n17398), .ZN(P3_U2749) );
  INV_X1 U20598 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17428) );
  AOI22_X1 U20599 ( .A1(n18679), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17419), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17399) );
  OAI21_X1 U20600 ( .B1(n17428), .B2(n17401), .A(n17399), .ZN(P3_U2750) );
  INV_X1 U20601 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17426) );
  AOI22_X1 U20602 ( .A1(n18679), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17419), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17400) );
  OAI21_X1 U20603 ( .B1(n17426), .B2(n17401), .A(n17400), .ZN(P3_U2751) );
  AOI22_X1 U20604 ( .A1(n18679), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17419), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17403) );
  OAI21_X1 U20605 ( .B1(n17489), .B2(n17422), .A(n17403), .ZN(P3_U2752) );
  AOI22_X1 U20606 ( .A1(n18679), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17419), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17404) );
  OAI21_X1 U20607 ( .B1(n17484), .B2(n17422), .A(n17404), .ZN(P3_U2753) );
  INV_X1 U20608 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17481) );
  AOI22_X1 U20609 ( .A1(n18679), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17419), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17405) );
  OAI21_X1 U20610 ( .B1(n17481), .B2(n17422), .A(n17405), .ZN(P3_U2754) );
  AOI22_X1 U20611 ( .A1(n18679), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17419), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17406) );
  OAI21_X1 U20612 ( .B1(n17479), .B2(n17422), .A(n17406), .ZN(P3_U2755) );
  INV_X1 U20613 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17476) );
  AOI22_X1 U20614 ( .A1(n18679), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17412), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17407) );
  OAI21_X1 U20615 ( .B1(n17476), .B2(n17422), .A(n17407), .ZN(P3_U2756) );
  AOI22_X1 U20616 ( .A1(n18679), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17412), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17408) );
  OAI21_X1 U20617 ( .B1(n17474), .B2(n17422), .A(n17408), .ZN(P3_U2757) );
  AOI22_X1 U20618 ( .A1(n18679), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17412), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17409) );
  OAI21_X1 U20619 ( .B1(n17472), .B2(n17422), .A(n17409), .ZN(P3_U2758) );
  AOI22_X1 U20620 ( .A1(n18679), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17412), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17410) );
  OAI21_X1 U20621 ( .B1(n20778), .B2(n17422), .A(n17410), .ZN(P3_U2759) );
  INV_X1 U20622 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17469) );
  AOI22_X1 U20623 ( .A1(n18679), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17412), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17411) );
  OAI21_X1 U20624 ( .B1(n17469), .B2(n17422), .A(n17411), .ZN(P3_U2760) );
  AOI22_X1 U20625 ( .A1(n18679), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17412), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17413) );
  OAI21_X1 U20626 ( .B1(n17467), .B2(n17422), .A(n17413), .ZN(P3_U2761) );
  INV_X1 U20627 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n17465) );
  AOI22_X1 U20628 ( .A1(n18679), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17419), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17414) );
  OAI21_X1 U20629 ( .B1(n17465), .B2(n17422), .A(n17414), .ZN(P3_U2762) );
  AOI22_X1 U20630 ( .A1(n18679), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17419), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17415) );
  OAI21_X1 U20631 ( .B1(n17463), .B2(n17422), .A(n17415), .ZN(P3_U2763) );
  INV_X1 U20632 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17461) );
  AOI22_X1 U20633 ( .A1(n18679), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17419), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17416) );
  OAI21_X1 U20634 ( .B1(n17461), .B2(n17422), .A(n17416), .ZN(P3_U2764) );
  AOI22_X1 U20635 ( .A1(n18679), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17419), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17417) );
  OAI21_X1 U20636 ( .B1(n17459), .B2(n17422), .A(n17417), .ZN(P3_U2765) );
  INV_X1 U20637 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17457) );
  AOI22_X1 U20638 ( .A1(n18679), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17419), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17418) );
  OAI21_X1 U20639 ( .B1(n17457), .B2(n17422), .A(n17418), .ZN(P3_U2766) );
  AOI22_X1 U20640 ( .A1(n18679), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17419), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17421) );
  OAI21_X1 U20641 ( .B1(n17455), .B2(n17422), .A(n17421), .ZN(P3_U2767) );
  AND2_X1 U20642 ( .A1(n18834), .A2(n17424), .ZN(n18676) );
  OAI211_X1 U20643 ( .C1(n18834), .C2(n18835), .A(n17424), .B(n17423), .ZN(
        n17477) );
  AOI22_X1 U20644 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17482), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17485), .ZN(n17425) );
  OAI21_X1 U20645 ( .B1(n17426), .B2(n17488), .A(n17425), .ZN(P3_U2768) );
  AOI22_X1 U20646 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17482), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17485), .ZN(n17427) );
  OAI21_X1 U20647 ( .B1(n17428), .B2(n17488), .A(n17427), .ZN(P3_U2769) );
  AOI22_X1 U20648 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17482), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17485), .ZN(n17429) );
  OAI21_X1 U20649 ( .B1(n17430), .B2(n17488), .A(n17429), .ZN(P3_U2770) );
  AOI22_X1 U20650 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17482), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17485), .ZN(n17431) );
  OAI21_X1 U20651 ( .B1(n17432), .B2(n17488), .A(n17431), .ZN(P3_U2771) );
  AOI22_X1 U20652 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17486), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17485), .ZN(n17433) );
  OAI21_X1 U20653 ( .B1(n17434), .B2(n17488), .A(n17433), .ZN(P3_U2772) );
  AOI22_X1 U20654 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17486), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17485), .ZN(n17435) );
  OAI21_X1 U20655 ( .B1(n17436), .B2(n17488), .A(n17435), .ZN(P3_U2773) );
  AOI22_X1 U20656 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17486), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17485), .ZN(n17437) );
  OAI21_X1 U20657 ( .B1(n17438), .B2(n17488), .A(n17437), .ZN(P3_U2774) );
  AOI22_X1 U20658 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17486), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17485), .ZN(n17439) );
  OAI21_X1 U20659 ( .B1(n17440), .B2(n17488), .A(n17439), .ZN(P3_U2775) );
  AOI22_X1 U20660 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17486), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17485), .ZN(n17441) );
  OAI21_X1 U20661 ( .B1(n17442), .B2(n17488), .A(n17441), .ZN(P3_U2776) );
  AOI22_X1 U20662 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17486), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17485), .ZN(n17443) );
  OAI21_X1 U20663 ( .B1(n17444), .B2(n17488), .A(n17443), .ZN(P3_U2777) );
  AOI22_X1 U20664 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17486), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17485), .ZN(n17445) );
  OAI21_X1 U20665 ( .B1(n17446), .B2(n17488), .A(n17445), .ZN(P3_U2778) );
  AOI22_X1 U20666 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17486), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17485), .ZN(n17447) );
  OAI21_X1 U20667 ( .B1(n17448), .B2(n17488), .A(n17447), .ZN(P3_U2779) );
  AOI22_X1 U20668 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17482), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17485), .ZN(n17449) );
  OAI21_X1 U20669 ( .B1(n17450), .B2(n17488), .A(n17449), .ZN(P3_U2780) );
  AOI22_X1 U20670 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17482), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17485), .ZN(n17451) );
  OAI21_X1 U20671 ( .B1(n20935), .B2(n17488), .A(n17451), .ZN(P3_U2781) );
  AOI22_X1 U20672 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17482), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17485), .ZN(n17452) );
  OAI21_X1 U20673 ( .B1(n17453), .B2(n17488), .A(n17452), .ZN(P3_U2782) );
  AOI22_X1 U20674 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17482), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17485), .ZN(n17454) );
  OAI21_X1 U20675 ( .B1(n17455), .B2(n17488), .A(n17454), .ZN(P3_U2783) );
  AOI22_X1 U20676 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17482), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17485), .ZN(n17456) );
  OAI21_X1 U20677 ( .B1(n17457), .B2(n17488), .A(n17456), .ZN(P3_U2784) );
  AOI22_X1 U20678 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17482), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17485), .ZN(n17458) );
  OAI21_X1 U20679 ( .B1(n17459), .B2(n17488), .A(n17458), .ZN(P3_U2785) );
  AOI22_X1 U20680 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17482), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17477), .ZN(n17460) );
  OAI21_X1 U20681 ( .B1(n17461), .B2(n17488), .A(n17460), .ZN(P3_U2786) );
  AOI22_X1 U20682 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17482), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17477), .ZN(n17462) );
  OAI21_X1 U20683 ( .B1(n17463), .B2(n17488), .A(n17462), .ZN(P3_U2787) );
  AOI22_X1 U20684 ( .A1(BUF2_REG_5__SCAN_IN), .A2(n17482), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17477), .ZN(n17464) );
  OAI21_X1 U20685 ( .B1(n17465), .B2(n17488), .A(n17464), .ZN(P3_U2788) );
  AOI22_X1 U20686 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17482), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17477), .ZN(n17466) );
  OAI21_X1 U20687 ( .B1(n17467), .B2(n17488), .A(n17466), .ZN(P3_U2789) );
  AOI22_X1 U20688 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17482), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17477), .ZN(n17468) );
  OAI21_X1 U20689 ( .B1(n17469), .B2(n17488), .A(n17468), .ZN(P3_U2790) );
  AOI22_X1 U20690 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17482), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17477), .ZN(n17470) );
  OAI21_X1 U20691 ( .B1(n20778), .B2(n17488), .A(n17470), .ZN(P3_U2791) );
  AOI22_X1 U20692 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17482), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17477), .ZN(n17471) );
  OAI21_X1 U20693 ( .B1(n17472), .B2(n17488), .A(n17471), .ZN(P3_U2792) );
  AOI22_X1 U20694 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17486), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17477), .ZN(n17473) );
  OAI21_X1 U20695 ( .B1(n17474), .B2(n17488), .A(n17473), .ZN(P3_U2793) );
  AOI22_X1 U20696 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17482), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17477), .ZN(n17475) );
  OAI21_X1 U20697 ( .B1(n17476), .B2(n17488), .A(n17475), .ZN(P3_U2794) );
  AOI22_X1 U20698 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17482), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17477), .ZN(n17478) );
  OAI21_X1 U20699 ( .B1(n17479), .B2(n17488), .A(n17478), .ZN(P3_U2795) );
  AOI22_X1 U20700 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17486), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17485), .ZN(n17480) );
  OAI21_X1 U20701 ( .B1(n17481), .B2(n17488), .A(n17480), .ZN(P3_U2796) );
  AOI22_X1 U20702 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17482), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17485), .ZN(n17483) );
  OAI21_X1 U20703 ( .B1(n17484), .B2(n17488), .A(n17483), .ZN(P3_U2797) );
  AOI22_X1 U20704 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17486), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17485), .ZN(n17487) );
  OAI21_X1 U20705 ( .B1(n17489), .B2(n17488), .A(n17487), .ZN(P3_U2798) );
  OR2_X1 U20706 ( .A1(n17492), .A2(n17696), .ZN(n17513) );
  OAI21_X1 U20707 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A(n17491), .ZN(n17498) );
  AOI21_X1 U20708 ( .B1(n17492), .B2(n17819), .A(n17817), .ZN(n17493) );
  INV_X1 U20709 ( .A(n17493), .ZN(n17494) );
  AOI21_X1 U20710 ( .B1(n17685), .B2(n17495), .A(n17494), .ZN(n17526) );
  OAI21_X1 U20711 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17598), .A(
        n17526), .ZN(n17516) );
  AOI22_X1 U20712 ( .A1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n17516), .B1(
        n17688), .B2(n17496), .ZN(n17497) );
  OAI21_X1 U20713 ( .B1(n17513), .B2(n17498), .A(n17497), .ZN(n17499) );
  AOI211_X1 U20714 ( .C1(n17501), .C2(n17565), .A(n17500), .B(n17499), .ZN(
        n17508) );
  NAND2_X1 U20715 ( .A1(n17863), .A2(n17773), .ZN(n17596) );
  AOI22_X1 U20716 ( .A1(n17848), .A2(n17871), .B1(n17725), .B2(n17870), .ZN(
        n17529) );
  NAND2_X1 U20717 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17529), .ZN(
        n17502) );
  NAND3_X1 U20718 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17596), .A3(
        n17502), .ZN(n17507) );
  OAI211_X1 U20719 ( .C1(n17505), .C2(n17504), .A(n17770), .B(n17503), .ZN(
        n17506) );
  NAND3_X1 U20720 ( .A1(n17508), .A2(n17507), .A3(n17506), .ZN(P3_U2802) );
  OAI22_X1 U20721 ( .A1(n9642), .A2(n18759), .B1(n17715), .B2(n17509), .ZN(
        n17515) );
  OR2_X2 U20722 ( .A1(n17511), .A2(n17510), .ZN(n17512) );
  XNOR2_X2 U20723 ( .A(n17512), .B(n17769), .ZN(n17881) );
  OAI22_X1 U20724 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17513), .B1(
        n17881), .B2(n17727), .ZN(n17514) );
  OAI221_X1 U20725 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17519), 
        .C1(n17518), .C2(n17529), .A(n17517), .ZN(P3_U2803) );
  INV_X1 U20726 ( .A(n17869), .ZN(n17894) );
  NAND3_X1 U20727 ( .A1(n17894), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A3(
        n17565), .ZN(n17530) );
  XOR2_X1 U20728 ( .A(n17888), .B(n17520), .Z(n17884) );
  AOI21_X1 U20729 ( .B1(n17521), .B2(n18571), .A(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17525) );
  INV_X1 U20730 ( .A(n17598), .ZN(n17523) );
  OAI21_X1 U20731 ( .B1(n17688), .B2(n17523), .A(n17522), .ZN(n17524) );
  NAND2_X1 U20732 ( .A1(n16412), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17886) );
  OAI211_X1 U20733 ( .C1(n17526), .C2(n17525), .A(n17524), .B(n17886), .ZN(
        n17527) );
  AOI21_X1 U20734 ( .B1(n17770), .B2(n17884), .A(n17527), .ZN(n17528) );
  OAI221_X1 U20735 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17530), 
        .C1(n17888), .C2(n17529), .A(n17528), .ZN(P3_U2804) );
  NAND3_X1 U20736 ( .A1(n17924), .A2(n17551), .A3(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17531) );
  XOR2_X1 U20737 ( .A(n17531), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17898) );
  AND2_X1 U20738 ( .A1(n17533), .A2(n18571), .ZN(n17558) );
  AOI211_X1 U20739 ( .C1(n17685), .C2(n17532), .A(n17817), .B(n17558), .ZN(
        n17562) );
  OAI21_X1 U20740 ( .B1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n17598), .A(
        n17562), .ZN(n17548) );
  NOR2_X1 U20741 ( .A1(n17696), .A2(n17533), .ZN(n17550) );
  OAI211_X1 U20742 ( .C1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17550), .B(n17534), .ZN(n17535) );
  NAND2_X1 U20743 ( .A1(n18174), .A2(P3_REIP_REG_25__SCAN_IN), .ZN(n17895) );
  OAI211_X1 U20744 ( .C1(n17715), .C2(n17536), .A(n17535), .B(n17895), .ZN(
        n17542) );
  NAND3_X1 U20745 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17551), .A3(
        n18015), .ZN(n17537) );
  XOR2_X1 U20746 ( .A(n17537), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17902) );
  OAI21_X1 U20747 ( .B1(n17587), .B2(n17539), .A(n17538), .ZN(n17540) );
  XOR2_X1 U20748 ( .A(n17540), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17897) );
  OAI22_X1 U20749 ( .A1(n17863), .A2(n17902), .B1(n17727), .B2(n17897), .ZN(
        n17541) );
  AOI211_X1 U20750 ( .C1(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .C2(n17548), .A(
        n17542), .B(n17541), .ZN(n17543) );
  OAI21_X1 U20751 ( .B1(n17773), .B2(n17898), .A(n17543), .ZN(P3_U2805) );
  AOI21_X1 U20752 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17545), .A(
        n17544), .ZN(n17916) );
  OAI22_X1 U20753 ( .A1(n9642), .A2(n18755), .B1(n17715), .B2(n17546), .ZN(
        n17547) );
  AOI221_X1 U20754 ( .B1(n17550), .B2(n17549), .C1(n17548), .C2(
        P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A(n17547), .ZN(n17553) );
  AND2_X1 U20755 ( .A1(n17924), .A2(n17551), .ZN(n17904) );
  AND2_X1 U20756 ( .A1(n18015), .A2(n17551), .ZN(n17903) );
  OAI22_X1 U20757 ( .A1(n17904), .A2(n17773), .B1(n17903), .B2(n17863), .ZN(
        n17564) );
  NOR2_X1 U20758 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17907), .ZN(
        n17912) );
  AOI22_X1 U20759 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17564), .B1(
        n17565), .B2(n17912), .ZN(n17552) );
  OAI211_X1 U20760 ( .C1(n17916), .C2(n17727), .A(n17553), .B(n17552), .ZN(
        P3_U2806) );
  AOI22_X1 U20761 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17587), .B1(
        n17554), .B2(n17568), .ZN(n17555) );
  NAND2_X1 U20762 ( .A1(n17604), .A2(n17555), .ZN(n17556) );
  XOR2_X1 U20763 ( .A(n17556), .B(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .Z(
        n17922) );
  NAND2_X1 U20764 ( .A1(n17715), .A2(n17598), .ZN(n17851) );
  AOI22_X1 U20765 ( .A1(n17559), .A2(n17558), .B1(n17557), .B2(n17851), .ZN(
        n17560) );
  NAND2_X1 U20766 ( .A1(n18174), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17921) );
  OAI211_X1 U20767 ( .C1(n17562), .C2(n17561), .A(n17560), .B(n17921), .ZN(
        n17563) );
  AOI221_X1 U20768 ( .B1(n17565), .B2(n17907), .C1(n17564), .C2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A(n17563), .ZN(n17566) );
  OAI21_X1 U20769 ( .B1(n17727), .B2(n17922), .A(n17566), .ZN(P3_U2807) );
  INV_X1 U20770 ( .A(n17604), .ZN(n17567) );
  AOI221_X1 U20771 ( .B1(n17934), .B2(n17568), .C1(n17586), .C2(n17568), .A(
        n17567), .ZN(n17569) );
  XOR2_X1 U20772 ( .A(n17935), .B(n17569), .Z(n17939) );
  NOR2_X1 U20773 ( .A1(n17570), .A2(n18696), .ZN(n17571) );
  AOI211_X1 U20774 ( .C1(n17819), .C2(n17572), .A(n17817), .B(n17571), .ZN(
        n17601) );
  OAI21_X1 U20775 ( .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n17598), .A(
        n17601), .ZN(n17583) );
  NAND2_X1 U20776 ( .A1(n18174), .A2(P3_REIP_REG_22__SCAN_IN), .ZN(n17937) );
  NOR2_X1 U20777 ( .A1(n17696), .A2(n17572), .ZN(n17585) );
  OAI211_X1 U20778 ( .C1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A(n17585), .B(n17573), .ZN(n17574) );
  OAI211_X1 U20779 ( .C1(n17575), .C2(n17715), .A(n17937), .B(n17574), .ZN(
        n17579) );
  NAND2_X1 U20780 ( .A1(n17626), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17941) );
  OR3_X1 U20781 ( .A1(n17594), .A2(n17591), .A3(n17941), .ZN(n17928) );
  NOR2_X1 U20782 ( .A1(n17655), .A2(n17928), .ZN(n17577) );
  OAI22_X1 U20783 ( .A1(n18015), .A2(n17863), .B1(n17924), .B2(n17773), .ZN(
        n17625) );
  AOI21_X1 U20784 ( .B1(n17596), .B2(n17928), .A(n17625), .ZN(n17595) );
  INV_X1 U20785 ( .A(n17595), .ZN(n17576) );
  MUX2_X1 U20786 ( .A(n17577), .B(n17576), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n17578) );
  AOI211_X1 U20787 ( .C1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(n17583), .A(
        n17579), .B(n17578), .ZN(n17580) );
  OAI21_X1 U20788 ( .B1(n17727), .B2(n17939), .A(n17580), .ZN(P3_U2808) );
  OAI22_X1 U20789 ( .A1(n9642), .A2(n18750), .B1(n17715), .B2(n17581), .ZN(
        n17582) );
  AOI221_X1 U20790 ( .B1(n17585), .B2(n17584), .C1(n17583), .C2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A(n17582), .ZN(n17593) );
  INV_X1 U20791 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17948) );
  NOR3_X1 U20792 ( .A1(n17948), .A2(n17587), .A3(n17586), .ZN(n17610) );
  INV_X1 U20793 ( .A(n17588), .ZN(n17628) );
  AOI22_X1 U20794 ( .A1(n17946), .A2(n17610), .B1(n17628), .B2(n17589), .ZN(
        n17590) );
  XOR2_X1 U20795 ( .A(n17594), .B(n17590), .Z(n17951) );
  NOR2_X1 U20796 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17591), .ZN(
        n17950) );
  NOR2_X1 U20797 ( .A1(n17655), .A2(n17941), .ZN(n17614) );
  AOI22_X1 U20798 ( .A1(n17770), .A2(n17951), .B1(n17950), .B2(n17614), .ZN(
        n17592) );
  OAI211_X1 U20799 ( .C1(n17595), .C2(n17594), .A(n17593), .B(n17592), .ZN(
        P3_U2809) );
  NOR2_X1 U20800 ( .A1(n17962), .A2(n17941), .ZN(n17925) );
  INV_X1 U20801 ( .A(n17925), .ZN(n17957) );
  AOI21_X1 U20802 ( .B1(n17596), .B2(n17957), .A(n17625), .ZN(n17612) );
  INV_X1 U20803 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17929) );
  INV_X1 U20804 ( .A(n17597), .ZN(n17603) );
  AOI21_X1 U20805 ( .B1(n17599), .B2(n18571), .A(
        P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n17600) );
  OAI22_X1 U20806 ( .A1(n17601), .A2(n17600), .B1(n9642), .B2(n18747), .ZN(
        n17602) );
  AOI221_X1 U20807 ( .B1(n17688), .B2(n17603), .C1(n17523), .C2(n17603), .A(
        n17602), .ZN(n17607) );
  OAI221_X1 U20808 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17627), 
        .C1(n17962), .C2(n17610), .A(n17604), .ZN(n17605) );
  XOR2_X1 U20809 ( .A(n17929), .B(n17605), .Z(n17955) );
  NOR2_X1 U20810 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17962), .ZN(
        n17954) );
  AOI22_X1 U20811 ( .A1(n17770), .A2(n17955), .B1(n17614), .B2(n17954), .ZN(
        n17606) );
  OAI211_X1 U20812 ( .C1(n17612), .C2(n17929), .A(n17607), .B(n17606), .ZN(
        P3_U2810) );
  AOI21_X1 U20813 ( .B1(n17819), .B2(n17615), .A(n17817), .ZN(n17637) );
  OAI21_X1 U20814 ( .B1(n17608), .B2(n18696), .A(n17637), .ZN(n17622) );
  AOI22_X1 U20815 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(n17622), .B1(
        n17688), .B2(n17609), .ZN(n17619) );
  AOI21_X1 U20816 ( .B1(n17628), .B2(n17627), .A(n17610), .ZN(n17611) );
  XOR2_X1 U20817 ( .A(n17611), .B(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .Z(
        n17967) );
  OAI22_X1 U20818 ( .A1(n17612), .A2(n17962), .B1(n17967), .B2(n17727), .ZN(
        n17613) );
  AOI21_X1 U20819 ( .B1(n17614), .B2(n17962), .A(n17613), .ZN(n17618) );
  NAND2_X1 U20820 ( .A1(n18174), .A2(P3_REIP_REG_19__SCAN_IN), .ZN(n17965) );
  NOR2_X1 U20821 ( .A1(n17696), .A2(n17615), .ZN(n17624) );
  OAI211_X1 U20822 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17624), .B(n17616), .ZN(n17617) );
  NAND4_X1 U20823 ( .A1(n17619), .A2(n17618), .A3(n17965), .A4(n17617), .ZN(
        P3_U2811) );
  NAND2_X1 U20824 ( .A1(n17626), .A2(n17948), .ZN(n17982) );
  OAI22_X1 U20825 ( .A1(n9642), .A2(n18743), .B1(n17715), .B2(n17620), .ZN(
        n17621) );
  AOI221_X1 U20826 ( .B1(n17624), .B2(n17623), .C1(n17622), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17621), .ZN(n17631) );
  INV_X1 U20827 ( .A(n17625), .ZN(n17654) );
  OAI21_X1 U20828 ( .B1(n17626), .B2(n17655), .A(n17654), .ZN(n17635) );
  AOI21_X1 U20829 ( .B1(n17769), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17627), .ZN(n17629) );
  XOR2_X1 U20830 ( .A(n17629), .B(n17628), .Z(n17978) );
  AOI22_X1 U20831 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17635), .B1(
        n17770), .B2(n17978), .ZN(n17630) );
  OAI211_X1 U20832 ( .C1(n17655), .C2(n17982), .A(n17631), .B(n17630), .ZN(
        P3_U2812) );
  OAI21_X1 U20833 ( .B1(n17633), .B2(n17983), .A(n17632), .ZN(n17987) );
  AOI22_X1 U20834 ( .A1(n17770), .A2(n17987), .B1(n17634), .B2(n17851), .ZN(
        n17642) );
  OAI221_X1 U20835 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .C2(n17636), .A(n17635), .ZN(
        n17641) );
  NAND2_X1 U20836 ( .A1(n18174), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n17988) );
  INV_X1 U20837 ( .A(n17637), .ZN(n17638) );
  OAI221_X1 U20838 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n17639), .C1(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .C2(n18571), .A(n17638), .ZN(
        n17640) );
  NAND4_X1 U20839 ( .A1(n17642), .A2(n17641), .A3(n17988), .A4(n17640), .ZN(
        P3_U2813) );
  AOI21_X1 U20840 ( .B1(n17769), .B2(n17644), .A(n17643), .ZN(n17645) );
  XOR2_X1 U20841 ( .A(n17645), .B(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .Z(
        n17998) );
  AOI21_X1 U20842 ( .B1(n17819), .B2(n17647), .A(n17817), .ZN(n17675) );
  OAI21_X1 U20843 ( .B1(n17646), .B2(n18696), .A(n17675), .ZN(n17658) );
  AOI22_X1 U20844 ( .A1(n18174), .A2(P3_REIP_REG_16__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n17658), .ZN(n17650) );
  NOR2_X1 U20845 ( .A1(n17696), .A2(n17647), .ZN(n17660) );
  OAI211_X1 U20846 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17660), .B(n17648), .ZN(n17649) );
  OAI211_X1 U20847 ( .C1(n17715), .C2(n17651), .A(n17650), .B(n17649), .ZN(
        n17652) );
  AOI21_X1 U20848 ( .B1(n17770), .B2(n17998), .A(n17652), .ZN(n17653) );
  OAI221_X1 U20849 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17655), 
        .C1(n18001), .C2(n17654), .A(n17653), .ZN(P3_U2814) );
  AOI21_X1 U20850 ( .B1(n18006), .B2(n17679), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n18009) );
  NAND2_X1 U20851 ( .A1(n17725), .A2(n18004), .ZN(n17670) );
  OAI22_X1 U20852 ( .A1(n9642), .A2(n20773), .B1(n17715), .B2(n17656), .ZN(
        n17657) );
  AOI221_X1 U20853 ( .B1(n17660), .B2(n17659), .C1(n17658), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17657), .ZN(n17669) );
  INV_X1 U20854 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17994) );
  INV_X1 U20855 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n18016) );
  INV_X1 U20856 ( .A(n17677), .ZN(n17662) );
  INV_X1 U20857 ( .A(n17690), .ZN(n17661) );
  NAND3_X1 U20858 ( .A1(n18060), .A2(n17662), .A3(n17661), .ZN(n17663) );
  NAND2_X1 U20859 ( .A1(n17664), .A2(n17663), .ZN(n17665) );
  OAI221_X1 U20860 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18016), 
        .C1(n9931), .C2(n17769), .A(n17665), .ZN(n17666) );
  XOR2_X1 U20861 ( .A(n17994), .B(n17666), .Z(n18010) );
  NOR2_X1 U20862 ( .A1(n18015), .A2(n17863), .ZN(n17667) );
  OR2_X1 U20863 ( .A1(n18038), .A2(n18053), .ZN(n18029) );
  OAI21_X1 U20864 ( .B1(n17677), .B2(n18029), .A(n17994), .ZN(n18003) );
  AOI22_X1 U20865 ( .A1(n17770), .A2(n18010), .B1(n17667), .B2(n18003), .ZN(
        n17668) );
  OAI211_X1 U20866 ( .C1(n18009), .C2(n17670), .A(n17669), .B(n17668), .ZN(
        P3_U2815) );
  NOR2_X1 U20867 ( .A1(n18038), .A2(n18051), .ZN(n18032) );
  NAND2_X1 U20868 ( .A1(n18006), .A2(n17679), .ZN(n17671) );
  OAI221_X1 U20869 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C1(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .C2(n18032), .A(n17671), .ZN(
        n18020) );
  AOI21_X1 U20870 ( .B1(n17672), .B2(n18571), .A(
        P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17674) );
  OAI22_X1 U20871 ( .A1(n17675), .A2(n17674), .B1(n17842), .B2(n17673), .ZN(
        n17676) );
  AOI21_X1 U20872 ( .B1(n18174), .B2(P3_REIP_REG_14__SCAN_IN), .A(n17676), 
        .ZN(n17683) );
  NOR2_X1 U20873 ( .A1(n17677), .A2(n18029), .ZN(n17678) );
  AOI221_X1 U20874 ( .B1(n17693), .B2(n18016), .C1(n18029), .C2(n18016), .A(
        n17678), .ZN(n18024) );
  NAND2_X1 U20875 ( .A1(n17769), .A2(n17679), .ZN(n17745) );
  INV_X1 U20876 ( .A(n17745), .ZN(n17706) );
  NOR2_X1 U20877 ( .A1(n18038), .A2(n17693), .ZN(n18017) );
  AOI21_X1 U20878 ( .B1(n17706), .B2(n18017), .A(n17680), .ZN(n17681) );
  XOR2_X1 U20879 ( .A(n18016), .B(n17681), .Z(n18023) );
  AOI22_X1 U20880 ( .A1(n17848), .A2(n18024), .B1(n17770), .B2(n18023), .ZN(
        n17682) );
  OAI211_X1 U20881 ( .C1(n17773), .C2(n18020), .A(n17683), .B(n17682), .ZN(
        P3_U2816) );
  AOI22_X1 U20882 ( .A1(n17685), .A2(n17684), .B1(n17819), .B2(n17695), .ZN(
        n17686) );
  NAND2_X1 U20883 ( .A1(n17686), .A2(n17859), .ZN(n17703) );
  AOI22_X1 U20884 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17703), .B1(
        n17688), .B2(n17687), .ZN(n17701) );
  NOR2_X1 U20885 ( .A1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n18038), .ZN(
        n18028) );
  INV_X1 U20886 ( .A(n18032), .ZN(n17689) );
  AOI22_X1 U20887 ( .A1(n17848), .A2(n18029), .B1(n17725), .B2(n17689), .ZN(
        n17709) );
  OAI22_X1 U20888 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17769), .B1(
        n17690), .B2(n18038), .ZN(n17691) );
  OAI21_X1 U20889 ( .B1(n17769), .B2(n17707), .A(n17691), .ZN(n17692) );
  XOR2_X1 U20890 ( .A(n17692), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n18037) );
  OAI22_X1 U20891 ( .A1(n17709), .A2(n17693), .B1(n17727), .B2(n18037), .ZN(
        n17694) );
  AOI21_X1 U20892 ( .B1(n18028), .B2(n17732), .A(n17694), .ZN(n17700) );
  NAND2_X1 U20893 ( .A1(n18174), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17699) );
  NOR2_X1 U20894 ( .A1(n17696), .A2(n17695), .ZN(n17705) );
  OAI211_X1 U20895 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17705), .B(n17697), .ZN(n17698) );
  NAND4_X1 U20896 ( .A1(n17701), .A2(n17700), .A3(n17699), .A4(n17698), .ZN(
        P3_U2817) );
  NOR2_X1 U20897 ( .A1(n9642), .A2(n20954), .ZN(n17702) );
  AOI221_X1 U20898 ( .B1(n17705), .B2(n17704), .C1(n17703), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17702), .ZN(n17713) );
  INV_X1 U20899 ( .A(n18060), .ZN(n18040) );
  NOR2_X1 U20900 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18040), .ZN(
        n17711) );
  NAND2_X1 U20901 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n17706), .ZN(
        n17734) );
  NOR2_X1 U20902 ( .A1(n18072), .A2(n17734), .ZN(n17722) );
  AOI21_X1 U20903 ( .B1(n17722), .B2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n17707), .ZN(n17708) );
  XOR2_X1 U20904 ( .A(n17708), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n18047) );
  OAI22_X1 U20905 ( .A1(n18047), .A2(n17727), .B1(n17709), .B2(n9931), .ZN(
        n17710) );
  AOI21_X1 U20906 ( .B1(n17711), .B2(n17732), .A(n17710), .ZN(n17712) );
  OAI211_X1 U20907 ( .C1(n17715), .C2(n17714), .A(n17713), .B(n17712), .ZN(
        P3_U2818) );
  NOR2_X1 U20908 ( .A1(n17716), .A2(n18397), .ZN(n17790) );
  NAND2_X1 U20909 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17790), .ZN(
        n17775) );
  NOR2_X1 U20910 ( .A1(n17717), .A2(n17775), .ZN(n17747) );
  NAND2_X1 U20911 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17747), .ZN(
        n17736) );
  INV_X1 U20912 ( .A(n17736), .ZN(n17751) );
  NAND2_X1 U20913 ( .A1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A2(n17751), .ZN(
        n17739) );
  INV_X1 U20914 ( .A(n17739), .ZN(n17721) );
  NOR2_X1 U20915 ( .A1(n17721), .A2(n17720), .ZN(n17719) );
  INV_X1 U20916 ( .A(n17856), .ZN(n17748) );
  INV_X1 U20917 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18733) );
  NOR2_X1 U20918 ( .A1(n9642), .A2(n18733), .ZN(n17718) );
  AOI221_X1 U20919 ( .B1(n17721), .B2(n17720), .C1(n17719), .C2(n17748), .A(
        n17718), .ZN(n17730) );
  NOR2_X1 U20920 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18058), .ZN(
        n18048) );
  AOI21_X1 U20921 ( .B1(n17723), .B2(n18072), .A(n17722), .ZN(n17724) );
  XOR2_X1 U20922 ( .A(n17724), .B(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .Z(
        n18066) );
  AOI22_X1 U20923 ( .A1(n18051), .A2(n17725), .B1(n17848), .B2(n18053), .ZN(
        n17755) );
  INV_X1 U20924 ( .A(n17755), .ZN(n17726) );
  AOI21_X1 U20925 ( .B1(n18058), .B2(n17732), .A(n17726), .ZN(n17743) );
  OAI22_X1 U20926 ( .A1(n18066), .A2(n17727), .B1(n17743), .B2(n15712), .ZN(
        n17728) );
  AOI21_X1 U20927 ( .B1(n18048), .B2(n17732), .A(n17728), .ZN(n17729) );
  OAI211_X1 U20928 ( .C1(n17842), .C2(n17731), .A(n17730), .B(n17729), .ZN(
        P3_U2819) );
  AOI21_X1 U20929 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17732), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17742) );
  AOI22_X1 U20930 ( .A1(n18174), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n17733), 
        .B2(n17851), .ZN(n17741) );
  OAI21_X1 U20931 ( .B1(n17744), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17734), .ZN(n17735) );
  XOR2_X1 U20932 ( .A(n17735), .B(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .Z(
        n18069) );
  OAI21_X1 U20933 ( .B1(n17856), .B2(n17737), .A(n17736), .ZN(n17738) );
  AOI22_X1 U20934 ( .A1(n17770), .A2(n18069), .B1(n17739), .B2(n17738), .ZN(
        n17740) );
  OAI211_X1 U20935 ( .C1(n17743), .C2(n17742), .A(n17741), .B(n17740), .ZN(
        P3_U2820) );
  INV_X1 U20936 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18080) );
  NAND2_X1 U20937 ( .A1(n17745), .A2(n17744), .ZN(n17746) );
  XOR2_X1 U20938 ( .A(n17746), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n18082) );
  NOR2_X1 U20939 ( .A1(n9642), .A2(n18729), .ZN(n17753) );
  AOI21_X1 U20940 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n17748), .A(
        n17747), .ZN(n17750) );
  OAI22_X1 U20941 ( .A1(n17751), .A2(n17750), .B1(n17842), .B2(n17749), .ZN(
        n17752) );
  AOI211_X1 U20942 ( .C1(n17770), .C2(n18082), .A(n17753), .B(n17752), .ZN(
        n17754) );
  OAI221_X1 U20943 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17756), .C1(
        n18080), .C2(n17755), .A(n17754), .ZN(P3_U2821) );
  NAND2_X1 U20944 ( .A1(n17757), .A2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n17759) );
  AOI211_X1 U20945 ( .C1(n17761), .C2(n17759), .A(n17758), .B(n18397), .ZN(
        n17763) );
  AOI21_X1 U20946 ( .B1(n17819), .B2(n17760), .A(n17817), .ZN(n17776) );
  OAI22_X1 U20947 ( .A1(n17776), .A2(n17761), .B1(n9642), .B2(n18728), .ZN(
        n17762) );
  AOI211_X1 U20948 ( .C1(n17764), .C2(n17851), .A(n17763), .B(n17762), .ZN(
        n17772) );
  AOI21_X1 U20949 ( .B1(n17766), .B2(n18092), .A(n17765), .ZN(n18096) );
  OAI21_X1 U20950 ( .B1(n17769), .B2(n17768), .A(n17767), .ZN(n18094) );
  AOI22_X1 U20951 ( .A1(n17848), .A2(n18096), .B1(n17770), .B2(n18094), .ZN(
        n17771) );
  OAI211_X1 U20952 ( .C1(n17773), .C2(n18100), .A(n17772), .B(n17771), .ZN(
        P3_U2822) );
  INV_X1 U20953 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17774) );
  AOI22_X1 U20954 ( .A1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A2(n17776), .B1(
        n17775), .B2(n17774), .ZN(n17777) );
  AOI21_X1 U20955 ( .B1(n18174), .B2(P3_REIP_REG_7__SCAN_IN), .A(n17777), .ZN(
        n17785) );
  NAND2_X1 U20956 ( .A1(n17779), .A2(n17778), .ZN(n17780) );
  XOR2_X1 U20957 ( .A(n17780), .B(n17783), .Z(n18107) );
  AOI21_X1 U20958 ( .B1(n17783), .B2(n17782), .A(n17781), .ZN(n18106) );
  AOI22_X1 U20959 ( .A1(n17848), .A2(n18107), .B1(n17852), .B2(n18106), .ZN(
        n17784) );
  OAI211_X1 U20960 ( .C1(n17842), .C2(n17786), .A(n17785), .B(n17784), .ZN(
        P3_U2823) );
  AOI21_X1 U20961 ( .B1(n17788), .B2(n17787), .A(n9729), .ZN(n18116) );
  AOI22_X1 U20962 ( .A1(n17852), .A2(n18116), .B1(n17790), .B2(n17789), .ZN(
        n17796) );
  NOR2_X1 U20963 ( .A1(n17856), .A2(n17790), .ZN(n17805) );
  AOI22_X1 U20964 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17805), .B1(
        n17791), .B2(n17851), .ZN(n17795) );
  AOI21_X1 U20965 ( .B1(n17793), .B2(n18113), .A(n17792), .ZN(n18110) );
  NAND2_X1 U20966 ( .A1(n17848), .A2(n18110), .ZN(n17794) );
  NAND2_X1 U20967 ( .A1(n18174), .A2(P3_REIP_REG_6__SCAN_IN), .ZN(n18112) );
  NAND4_X1 U20968 ( .A1(n17796), .A2(n17795), .A3(n17794), .A4(n18112), .ZN(
        P3_U2824) );
  AOI21_X1 U20969 ( .B1(n17799), .B2(n17798), .A(n17797), .ZN(n18125) );
  NOR2_X1 U20970 ( .A1(n17801), .A2(n17800), .ZN(n17803) );
  XOR2_X1 U20971 ( .A(n17803), .B(n17802), .Z(n18127) );
  OAI22_X1 U20972 ( .A1(n17862), .A2(n18127), .B1(n9642), .B2(n18722), .ZN(
        n17804) );
  AOI21_X1 U20973 ( .B1(n17848), .B2(n18125), .A(n17804), .ZN(n17808) );
  OAI221_X1 U20974 ( .B1(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n17806), .C1(
        P3_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n17859), .A(n17805), .ZN(n17807) );
  OAI211_X1 U20975 ( .C1(n17842), .C2(n17809), .A(n17808), .B(n17807), .ZN(
        P3_U2825) );
  OAI21_X1 U20976 ( .B1(n17812), .B2(n17811), .A(n17810), .ZN(n17813) );
  XOR2_X1 U20977 ( .A(n17813), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(
        n18140) );
  AOI22_X1 U20978 ( .A1(n18174), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18571), 
        .B2(n17814), .ZN(n17824) );
  AOI21_X1 U20979 ( .B1(n17816), .B2(n17815), .A(n9737), .ZN(n18128) );
  AOI21_X1 U20980 ( .B1(n17819), .B2(n17818), .A(n17817), .ZN(n17834) );
  OAI22_X1 U20981 ( .A1(n17842), .A2(n17821), .B1(n17820), .B2(n17834), .ZN(
        n17822) );
  AOI21_X1 U20982 ( .B1(n17852), .B2(n18128), .A(n17822), .ZN(n17823) );
  OAI211_X1 U20983 ( .C1(n17863), .C2(n18140), .A(n17824), .B(n17823), .ZN(
        P3_U2826) );
  AOI21_X1 U20984 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n17859), .A(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17835) );
  AOI21_X1 U20985 ( .B1(n17827), .B2(n17826), .A(n17825), .ZN(n18143) );
  AOI22_X1 U20986 ( .A1(n17852), .A2(n18143), .B1(n18174), .B2(
        P3_REIP_REG_3__SCAN_IN), .ZN(n17833) );
  AOI21_X1 U20987 ( .B1(n17830), .B2(n17829), .A(n17828), .ZN(n18144) );
  AOI22_X1 U20988 ( .A1(n17848), .A2(n18144), .B1(n17831), .B2(n17851), .ZN(
        n17832) );
  OAI211_X1 U20989 ( .C1(n17835), .C2(n17834), .A(n17833), .B(n17832), .ZN(
        P3_U2827) );
  INV_X1 U20990 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n17846) );
  AOI21_X1 U20991 ( .B1(n17838), .B2(n17837), .A(n17836), .ZN(n18158) );
  NAND2_X1 U20992 ( .A1(n18174), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18160) );
  INV_X1 U20993 ( .A(n18160), .ZN(n17844) );
  XNOR2_X1 U20994 ( .A(n17840), .B(n17839), .ZN(n18157) );
  OAI22_X1 U20995 ( .A1(n17842), .A2(n17841), .B1(n17863), .B2(n18157), .ZN(
        n17843) );
  AOI211_X1 U20996 ( .C1(n17852), .C2(n18158), .A(n17844), .B(n17843), .ZN(
        n17845) );
  OAI221_X1 U20997 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n18397), .C1(
        n17846), .C2(n17859), .A(n17845), .ZN(P3_U2828) );
  NOR2_X1 U20998 ( .A1(n17858), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n17847) );
  XNOR2_X1 U20999 ( .A(n17850), .B(n17847), .ZN(n18165) );
  AOI22_X1 U21000 ( .A1(n17848), .A2(n18165), .B1(n18174), .B2(
        P3_REIP_REG_1__SCAN_IN), .ZN(n17854) );
  AOI21_X1 U21001 ( .B1(n17850), .B2(n17857), .A(n17849), .ZN(n18163) );
  AOI22_X1 U21002 ( .A1(n17852), .A2(n18163), .B1(n17855), .B2(n17851), .ZN(
        n17853) );
  OAI211_X1 U21003 ( .C1(n17856), .C2(n17855), .A(n17854), .B(n17853), .ZN(
        P3_U2829) );
  OAI21_X1 U21004 ( .B1(n17858), .B2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n17857), .ZN(n18182) );
  INV_X1 U21005 ( .A(n18182), .ZN(n17864) );
  OAI21_X1 U21006 ( .B1(n18688), .B2(n18837), .A(n17859), .ZN(n17860) );
  AOI22_X1 U21007 ( .A1(n18174), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17860), .ZN(n17861) );
  OAI221_X1 U21008 ( .B1(n17864), .B2(n17863), .C1(n18182), .C2(n17862), .A(
        n17861), .ZN(P3_U2830) );
  NOR2_X1 U21009 ( .A1(n17865), .A2(n17917), .ZN(n17877) );
  NOR2_X1 U21010 ( .A1(n18655), .A2(n18636), .ZN(n18087) );
  INV_X1 U21011 ( .A(n18087), .ZN(n18130) );
  AOI21_X1 U21012 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18635), .A(
        n17866), .ZN(n17932) );
  NOR2_X1 U21013 ( .A1(n17934), .A2(n17932), .ZN(n17868) );
  AOI21_X1 U21014 ( .B1(n17868), .B2(n17867), .A(n18087), .ZN(n17906) );
  AOI21_X1 U21015 ( .B1(n17869), .B2(n18130), .A(n17906), .ZN(n17889) );
  AOI22_X1 U21016 ( .A1(n18054), .A2(n17871), .B1(n18052), .B2(n17870), .ZN(
        n17872) );
  NAND2_X1 U21017 ( .A1(n17889), .A2(n17872), .ZN(n17873) );
  AOI211_X1 U21018 ( .C1(n17875), .C2(n18130), .A(n17874), .B(n17873), .ZN(
        n17882) );
  INV_X1 U21019 ( .A(n17882), .ZN(n17876) );
  MUX2_X1 U21020 ( .A(n17877), .B(n17876), .S(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .Z(n17878) );
  AOI22_X1 U21021 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n18168), .B1(
        n18175), .B2(n17878), .ZN(n17880) );
  NAND2_X1 U21022 ( .A1(n18174), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17879) );
  OAI211_X1 U21023 ( .C1(n17881), .C2(n18065), .A(n17880), .B(n17879), .ZN(
        P3_U2835) );
  NAND2_X1 U21024 ( .A1(n17894), .A2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n17883) );
  AOI221_X1 U21025 ( .B1(n17917), .B2(n17888), .C1(n17883), .C2(n17888), .A(
        n17882), .ZN(n17885) );
  AOI22_X1 U21026 ( .A1(n18175), .A2(n17885), .B1(n9743), .B2(n17884), .ZN(
        n17887) );
  OAI211_X1 U21027 ( .C1(n18162), .C2(n17888), .A(n17887), .B(n17886), .ZN(
        P3_U2836) );
  OAI221_X1 U21028 ( .B1(n18661), .B2(n17894), .C1(n18661), .C2(n17890), .A(
        n17889), .ZN(n17892) );
  OAI222_X1 U21029 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(n17894), 
        .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17893), .C1(n17892), 
        .C2(n17891), .ZN(n17896) );
  OAI21_X1 U21030 ( .B1(n18166), .B2(n17896), .A(n17895), .ZN(n17900) );
  OAI22_X1 U21031 ( .A1(n18099), .A2(n17898), .B1(n18065), .B2(n17897), .ZN(
        n17899) );
  AOI211_X1 U21032 ( .C1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .C2(n18168), .A(
        n17900), .B(n17899), .ZN(n17901) );
  OAI21_X1 U21033 ( .B1(n18141), .B2(n17902), .A(n17901), .ZN(P3_U2837) );
  OAI22_X1 U21034 ( .A1(n17904), .A2(n18031), .B1(n17903), .B2(n18630), .ZN(
        n17905) );
  NOR3_X1 U21035 ( .A1(n18168), .A2(n17906), .A3(n17905), .ZN(n17910) );
  AOI21_X1 U21036 ( .B1(n18153), .B2(n17908), .A(n17907), .ZN(n17909) );
  AOI21_X1 U21037 ( .B1(n17910), .B2(n17909), .A(n18174), .ZN(n17918) );
  AOI21_X1 U21038 ( .B1(n18134), .B2(n17910), .A(n9908), .ZN(n17911) );
  AOI22_X1 U21039 ( .A1(n17913), .A2(n17912), .B1(n17918), .B2(n17911), .ZN(
        n17915) );
  NAND2_X1 U21040 ( .A1(n18174), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n17914) );
  OAI211_X1 U21041 ( .C1(n17916), .C2(n18065), .A(n17915), .B(n17914), .ZN(
        P3_U2838) );
  INV_X1 U21042 ( .A(n17917), .ZN(n17919) );
  OAI221_X1 U21043 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17919), 
        .C1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n18162), .A(n17918), .ZN(
        n17920) );
  OAI211_X1 U21044 ( .C1(n17922), .C2(n18065), .A(n17921), .B(n17920), .ZN(
        P3_U2839) );
  INV_X1 U21045 ( .A(n17923), .ZN(n17949) );
  NOR2_X1 U21046 ( .A1(n18061), .A2(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n17931) );
  OAI22_X1 U21047 ( .A1(n18015), .A2(n18630), .B1(n17924), .B2(n18031), .ZN(
        n17942) );
  AOI21_X1 U21048 ( .B1(n17926), .B2(n17925), .A(n18176), .ZN(n17927) );
  AOI221_X1 U21049 ( .B1(n17948), .B2(n18153), .C1(n17973), .C2(n18153), .A(
        n17927), .ZN(n17943) );
  NAND2_X1 U21050 ( .A1(n18630), .A2(n18031), .ZN(n18057) );
  AOI22_X1 U21051 ( .A1(n18655), .A2(n17929), .B1(n17928), .B2(n18057), .ZN(
        n17945) );
  OAI211_X1 U21052 ( .C1(n17946), .C2(n18661), .A(n17943), .B(n17945), .ZN(
        n17930) );
  NOR4_X1 U21053 ( .A1(n17932), .A2(n17931), .A3(n17942), .A4(n17930), .ZN(
        n17933) );
  AOI221_X1 U21054 ( .B1(n17949), .B2(n17935), .C1(n17934), .C2(n17935), .A(
        n17933), .ZN(n17936) );
  AOI22_X1 U21055 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18168), .B1(
        n18175), .B2(n17936), .ZN(n17938) );
  OAI211_X1 U21056 ( .C1(n17939), .C2(n18065), .A(n17938), .B(n17937), .ZN(
        P3_U2840) );
  NAND2_X1 U21057 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n17940), .ZN(
        n18049) );
  NOR3_X1 U21058 ( .A1(n17993), .A2(n17941), .A3(n18049), .ZN(n17944) );
  NOR2_X1 U21059 ( .A1(n18166), .A2(n17942), .ZN(n17990) );
  OAI211_X1 U21060 ( .C1(n18635), .C2(n17944), .A(n17990), .B(n17943), .ZN(
        n17956) );
  NOR2_X1 U21061 ( .A1(n18153), .A2(n18636), .ZN(n18167) );
  OAI21_X1 U21062 ( .B1(n17946), .B2(n18167), .A(n17945), .ZN(n17947) );
  OAI21_X1 U21063 ( .B1(n17956), .B2(n17947), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17953) );
  NOR3_X1 U21064 ( .A1(n17949), .A2(n18166), .A3(n17948), .ZN(n17963) );
  AOI22_X1 U21065 ( .A1(n9743), .A2(n17951), .B1(n17950), .B2(n17963), .ZN(
        n17952) );
  OAI221_X1 U21066 ( .B1(n18174), .B2(n17953), .C1(n9642), .C2(n18750), .A(
        n17952), .ZN(P3_U2841) );
  AOI22_X1 U21067 ( .A1(n9743), .A2(n17955), .B1(n17963), .B2(n17954), .ZN(
        n17961) );
  AOI21_X1 U21068 ( .B1(n18057), .B2(n17957), .A(n17956), .ZN(n17958) );
  NOR2_X1 U21069 ( .A1(n18174), .A2(n17958), .ZN(n17964) );
  NOR3_X1 U21070 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n18167), .A3(
        n18678), .ZN(n17959) );
  OAI21_X1 U21071 ( .B1(n17964), .B2(n17959), .A(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17960) );
  OAI211_X1 U21072 ( .C1(n18747), .C2(n9642), .A(n17961), .B(n17960), .ZN(
        P3_U2842) );
  AOI22_X1 U21073 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17964), .B1(
        n17963), .B2(n17962), .ZN(n17966) );
  OAI211_X1 U21074 ( .C1(n17967), .C2(n18065), .A(n17966), .B(n17965), .ZN(
        P3_U2843) );
  OAI22_X1 U21075 ( .A1(n18152), .A2(n18661), .B1(n18131), .B2(n17968), .ZN(
        n18142) );
  NAND2_X1 U21076 ( .A1(n17969), .A2(n18142), .ZN(n18101) );
  NOR3_X1 U21077 ( .A1(n18092), .A2(n18090), .A3(n18101), .ZN(n18018) );
  NOR2_X1 U21078 ( .A1(n18018), .A2(n17970), .ZN(n18041) );
  NAND2_X1 U21079 ( .A1(n17971), .A2(n18081), .ZN(n18002) );
  NOR2_X1 U21080 ( .A1(n18635), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18129) );
  NOR3_X1 U21081 ( .A1(n18129), .A2(n17972), .A3(n18001), .ZN(n17975) );
  NAND2_X1 U21082 ( .A1(n18153), .A2(n17973), .ZN(n17974) );
  OAI211_X1 U21083 ( .C1(n18087), .C2(n17975), .A(n17990), .B(n17974), .ZN(
        n17976) );
  AOI21_X1 U21084 ( .B1(n17977), .B2(n18057), .A(n17976), .ZN(n17984) );
  AOI221_X1 U21085 ( .B1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n17984), 
        .C1(n18087), .C2(n17984), .A(n18174), .ZN(n17979) );
  AOI22_X1 U21086 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17979), .B1(
        n9743), .B2(n17978), .ZN(n17981) );
  NAND2_X1 U21087 ( .A1(n18174), .A2(P3_REIP_REG_18__SCAN_IN), .ZN(n17980) );
  OAI211_X1 U21088 ( .C1(n17982), .C2(n18002), .A(n17981), .B(n17980), .ZN(
        P3_U2844) );
  NOR3_X1 U21089 ( .A1(n16412), .A2(n17984), .A3(n17983), .ZN(n17986) );
  NOR3_X1 U21090 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18001), .A3(
        n18002), .ZN(n17985) );
  AOI211_X1 U21091 ( .C1(n9743), .C2(n17987), .A(n17986), .B(n17985), .ZN(
        n17989) );
  NAND2_X1 U21092 ( .A1(n17989), .A2(n17988), .ZN(P3_U2845) );
  INV_X1 U21093 ( .A(n17990), .ZN(n17997) );
  OAI22_X1 U21094 ( .A1(n18176), .A2(n17992), .B1(n17991), .B2(n18661), .ZN(
        n18079) );
  AOI21_X1 U21095 ( .B1(n18655), .B2(n18092), .A(n18079), .ZN(n18050) );
  OAI22_X1 U21096 ( .A1(n18636), .A2(n17994), .B1(n17993), .B2(n18049), .ZN(
        n17995) );
  OAI211_X1 U21097 ( .C1(n18061), .C2(n18006), .A(n18050), .B(n17995), .ZN(
        n18005) );
  OAI221_X1 U21098 ( .B1(n17997), .B2(n17996), .C1(n17997), .C2(n18005), .A(
        n9642), .ZN(n18000) );
  AOI22_X1 U21099 ( .A1(n18174), .A2(P3_REIP_REG_16__SCAN_IN), .B1(n9743), 
        .B2(n17998), .ZN(n17999) );
  OAI221_X1 U21100 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n18002), 
        .C1(n18001), .C2(n18000), .A(n17999), .ZN(P3_U2846) );
  NAND2_X1 U21101 ( .A1(n18179), .A2(n18003), .ZN(n18014) );
  AOI22_X1 U21102 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n18168), .B1(
        n18174), .B2(P3_REIP_REG_15__SCAN_IN), .ZN(n18013) );
  NAND2_X1 U21103 ( .A1(n18052), .A2(n18004), .ZN(n18008) );
  OAI221_X1 U21104 ( .B1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18006), 
        .C1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n18018), .A(n18005), .ZN(
        n18007) );
  OAI21_X1 U21105 ( .B1(n18009), .B2(n18008), .A(n18007), .ZN(n18011) );
  AOI22_X1 U21106 ( .A1(n18175), .A2(n18011), .B1(n9743), .B2(n18010), .ZN(
        n18012) );
  OAI211_X1 U21107 ( .C1(n18015), .C2(n18014), .A(n18013), .B(n18012), .ZN(
        P3_U2847) );
  OAI21_X1 U21108 ( .B1(n18038), .B2(n18049), .A(n18636), .ZN(n18033) );
  OAI211_X1 U21109 ( .C1(n18134), .C2(n18017), .A(n18050), .B(n18033), .ZN(
        n18022) );
  NAND3_X1 U21110 ( .A1(n18018), .A2(n18017), .A3(n18016), .ZN(n18019) );
  OAI21_X1 U21111 ( .B1(n18020), .B2(n18031), .A(n18019), .ZN(n18021) );
  AOI21_X1 U21112 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n18022), .A(
        n18021), .ZN(n18027) );
  AOI22_X1 U21113 ( .A1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n18168), .B1(
        n18174), .B2(P3_REIP_REG_14__SCAN_IN), .ZN(n18026) );
  AOI22_X1 U21114 ( .A1(n18179), .A2(n18024), .B1(n9743), .B2(n18023), .ZN(
        n18025) );
  OAI211_X1 U21115 ( .C1(n18027), .C2(n18166), .A(n18026), .B(n18025), .ZN(
        P3_U2848) );
  AOI22_X1 U21116 ( .A1(n18174), .A2(P3_REIP_REG_13__SCAN_IN), .B1(n18081), 
        .B2(n18028), .ZN(n18036) );
  INV_X1 U21117 ( .A(n18061), .ZN(n18067) );
  AOI22_X1 U21118 ( .A1(n18054), .A2(n18029), .B1(n18067), .B2(n18040), .ZN(
        n18030) );
  OAI211_X1 U21119 ( .C1(n18032), .C2(n18031), .A(n18050), .B(n18030), .ZN(
        n18043) );
  OAI211_X1 U21120 ( .C1(n18061), .C2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A(
        n18175), .B(n18033), .ZN(n18034) );
  OAI211_X1 U21121 ( .C1(n18043), .C2(n18034), .A(
        P3_INSTADDRPOINTER_REG_13__SCAN_IN), .B(n9642), .ZN(n18035) );
  OAI211_X1 U21122 ( .C1(n18037), .C2(n18065), .A(n18036), .B(n18035), .ZN(
        P3_U2849) );
  AOI22_X1 U21123 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n18168), .B1(
        n18174), .B2(P3_REIP_REG_12__SCAN_IN), .ZN(n18046) );
  NOR2_X1 U21124 ( .A1(n18038), .A2(n18049), .ZN(n18039) );
  AOI21_X1 U21125 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n18635), .A(
        n18039), .ZN(n18044) );
  OAI21_X1 U21126 ( .B1(n18041), .B2(n18040), .A(n9931), .ZN(n18042) );
  OAI211_X1 U21127 ( .C1(n18044), .C2(n18043), .A(n18175), .B(n18042), .ZN(
        n18045) );
  OAI211_X1 U21128 ( .C1(n18047), .C2(n18065), .A(n18046), .B(n18045), .ZN(
        P3_U2850) );
  AOI22_X1 U21129 ( .A1(n18174), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n18081), 
        .B2(n18048), .ZN(n18064) );
  INV_X1 U21130 ( .A(n18049), .ZN(n18077) );
  INV_X1 U21131 ( .A(n18050), .ZN(n18056) );
  AOI22_X1 U21132 ( .A1(n18054), .A2(n18053), .B1(n18052), .B2(n18051), .ZN(
        n18055) );
  NAND2_X1 U21133 ( .A1(n18175), .A2(n18055), .ZN(n18074) );
  AOI211_X1 U21134 ( .C1(n18058), .C2(n18057), .A(n18056), .B(n18074), .ZN(
        n18059) );
  OAI221_X1 U21135 ( .B1(n18635), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .C1(
        n18635), .C2(n18077), .A(n18059), .ZN(n18068) );
  OAI22_X1 U21136 ( .A1(n18061), .A2(n18060), .B1(n18635), .B2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n18062) );
  OAI211_X1 U21137 ( .C1(n18068), .C2(n18062), .A(
        P3_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n9642), .ZN(n18063) );
  OAI211_X1 U21138 ( .C1(n18066), .C2(n18065), .A(n18064), .B(n18063), .ZN(
        P3_U2851) );
  NAND2_X1 U21139 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n18081), .ZN(
        n18073) );
  OAI221_X1 U21140 ( .B1(n18068), .B2(n18067), .C1(n18068), .C2(n18080), .A(
        n9642), .ZN(n18071) );
  AOI22_X1 U21141 ( .A1(n18174), .A2(P3_REIP_REG_10__SCAN_IN), .B1(n9743), 
        .B2(n18069), .ZN(n18070) );
  OAI221_X1 U21142 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n18073), 
        .C1(n18072), .C2(n18071), .A(n18070), .ZN(P3_U2852) );
  NAND2_X1 U21143 ( .A1(n18655), .A2(n18092), .ZN(n18076) );
  INV_X1 U21144 ( .A(n18074), .ZN(n18075) );
  OAI211_X1 U21145 ( .C1(n18077), .C2(n18635), .A(n18076), .B(n18075), .ZN(
        n18078) );
  OAI21_X1 U21146 ( .B1(n18079), .B2(n18078), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n18084) );
  AOI22_X1 U21147 ( .A1(n9743), .A2(n18082), .B1(n18081), .B2(n18080), .ZN(
        n18083) );
  OAI221_X1 U21148 ( .B1(n18174), .B2(n18084), .C1(n9642), .C2(n18729), .A(
        n18083), .ZN(P3_U2853) );
  NAND3_X1 U21149 ( .A1(n18142), .A2(n18175), .A3(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18119) );
  INV_X1 U21150 ( .A(n18119), .ZN(n18136) );
  NAND3_X1 U21151 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A3(n18136), .ZN(n18114) );
  NOR2_X1 U21152 ( .A1(n18090), .A2(n18114), .ZN(n18093) );
  INV_X1 U21153 ( .A(n18085), .ZN(n18089) );
  AOI21_X1 U21154 ( .B1(n18153), .B2(n18086), .A(n18129), .ZN(n18088) );
  AOI221_X1 U21155 ( .B1(n18089), .B2(n18088), .C1(n18087), .C2(n18088), .A(
        n18166), .ZN(n18111) );
  AOI21_X1 U21156 ( .B1(n18169), .B2(n18090), .A(n18111), .ZN(n18102) );
  NAND2_X1 U21157 ( .A1(n18102), .A2(n18162), .ZN(n18105) );
  NOR2_X1 U21158 ( .A1(n9642), .A2(n18728), .ZN(n18091) );
  AOI221_X1 U21159 ( .B1(n18093), .B2(n18092), .C1(n18105), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n18091), .ZN(n18098) );
  AOI22_X1 U21160 ( .A1(n18179), .A2(n18096), .B1(n9743), .B2(n18094), .ZN(
        n18097) );
  OAI211_X1 U21161 ( .C1(n18100), .C2(n18099), .A(n18098), .B(n18097), .ZN(
        P3_U2854) );
  INV_X1 U21162 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18725) );
  NOR2_X1 U21163 ( .A1(n9642), .A2(n18725), .ZN(n18104) );
  NOR3_X1 U21164 ( .A1(n18102), .A2(n18101), .A3(n18113), .ZN(n18103) );
  AOI211_X1 U21165 ( .C1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C2(n18105), .A(
        n18104), .B(n18103), .ZN(n18109) );
  AOI22_X1 U21166 ( .A1(n18179), .A2(n18107), .B1(n18164), .B2(n18106), .ZN(
        n18108) );
  NAND2_X1 U21167 ( .A1(n18109), .A2(n18108), .ZN(P3_U2855) );
  INV_X1 U21168 ( .A(n18110), .ZN(n18118) );
  NOR2_X1 U21169 ( .A1(n18168), .A2(n18111), .ZN(n18120) );
  OAI221_X1 U21170 ( .B1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n18114), .C1(
        n18113), .C2(n18120), .A(n18112), .ZN(n18115) );
  AOI21_X1 U21171 ( .B1(n18164), .B2(n18116), .A(n18115), .ZN(n18117) );
  OAI21_X1 U21172 ( .B1(n18141), .B2(n18118), .A(n18117), .ZN(P3_U2856) );
  NOR2_X1 U21173 ( .A1(n9642), .A2(n18722), .ZN(n18124) );
  NOR2_X1 U21174 ( .A1(n18135), .A2(n18119), .ZN(n18122) );
  INV_X1 U21175 ( .A(n18120), .ZN(n18121) );
  MUX2_X1 U21176 ( .A(n18122), .B(n18121), .S(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .Z(n18123) );
  AOI211_X1 U21177 ( .C1(n18125), .C2(n18179), .A(n18124), .B(n18123), .ZN(
        n18126) );
  OAI21_X1 U21178 ( .B1(n18183), .B2(n18127), .A(n18126), .ZN(P3_U2857) );
  AOI22_X1 U21179 ( .A1(n18174), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18164), 
        .B2(n18128), .ZN(n18139) );
  AOI21_X1 U21180 ( .B1(n18131), .B2(n18130), .A(n18129), .ZN(n18149) );
  OAI211_X1 U21181 ( .C1(n18661), .C2(n18132), .A(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .B(n18149), .ZN(n18133) );
  NAND2_X1 U21182 ( .A1(n18175), .A2(n18133), .ZN(n18147) );
  OAI21_X1 U21183 ( .B1(n18134), .B2(n18147), .A(n18162), .ZN(n18137) );
  AOI22_X1 U21184 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18137), .B1(
        n18136), .B2(n18135), .ZN(n18138) );
  OAI211_X1 U21185 ( .C1(n18141), .C2(n18140), .A(n18139), .B(n18138), .ZN(
        P3_U2858) );
  NOR2_X1 U21186 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18142), .ZN(
        n18148) );
  AOI22_X1 U21187 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18168), .B1(
        n18174), .B2(P3_REIP_REG_3__SCAN_IN), .ZN(n18146) );
  AOI22_X1 U21188 ( .A1(n18179), .A2(n18144), .B1(n18164), .B2(n18143), .ZN(
        n18145) );
  OAI211_X1 U21189 ( .C1(n18148), .C2(n18147), .A(n18146), .B(n18145), .ZN(
        P3_U2859) );
  NAND2_X1 U21190 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18150) );
  OAI21_X1 U21191 ( .B1(n18661), .B2(n18150), .A(n18149), .ZN(n18151) );
  AOI22_X1 U21192 ( .A1(n18153), .A2(n18152), .B1(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n18151), .ZN(n18156) );
  NAND3_X1 U21193 ( .A1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n18154), .A3(
        n15627), .ZN(n18155) );
  OAI211_X1 U21194 ( .C1(n18157), .C2(n18630), .A(n18156), .B(n18155), .ZN(
        n18159) );
  AOI22_X1 U21195 ( .A1(n18175), .A2(n18159), .B1(n18164), .B2(n18158), .ZN(
        n18161) );
  OAI211_X1 U21196 ( .C1(n18162), .C2(n15627), .A(n18161), .B(n18160), .ZN(
        P3_U2860) );
  AOI22_X1 U21197 ( .A1(n18179), .A2(n18165), .B1(n18164), .B2(n18163), .ZN(
        n18173) );
  NAND2_X1 U21198 ( .A1(n18174), .A2(P3_REIP_REG_1__SCAN_IN), .ZN(n18172) );
  NOR3_X1 U21199 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n18167), .A3(
        n18166), .ZN(n18178) );
  OAI21_X1 U21200 ( .B1(n18168), .B2(n18178), .A(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18171) );
  OAI211_X1 U21201 ( .C1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .C2(n18655), .A(
        n18169), .B(n18793), .ZN(n18170) );
  NAND4_X1 U21202 ( .A1(n18173), .A2(n18172), .A3(n18171), .A4(n18170), .ZN(
        P3_U2861) );
  AOI211_X1 U21203 ( .C1(n18176), .C2(n18175), .A(n18174), .B(n18810), .ZN(
        n18177) );
  AOI211_X1 U21204 ( .C1(n18179), .C2(n18182), .A(n18178), .B(n18177), .ZN(
        n18181) );
  NAND2_X1 U21205 ( .A1(n18174), .A2(P3_REIP_REG_0__SCAN_IN), .ZN(n18180) );
  OAI211_X1 U21206 ( .C1(n18183), .C2(n18182), .A(n18181), .B(n18180), .ZN(
        P3_U2862) );
  OAI211_X1 U21207 ( .C1(P3_FLUSH_REG_SCAN_IN), .C2(n18184), .A(
        P3_STATE2_REG_2__SCAN_IN), .B(P3_STATE2_REG_1__SCAN_IN), .ZN(n18685)
         );
  OAI21_X1 U21208 ( .B1(n18187), .B2(n18185), .A(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18186) );
  OAI221_X1 U21209 ( .B1(n18187), .B2(n18685), .C1(n18187), .C2(n18470), .A(
        n18186), .ZN(P3_U2863) );
  INV_X1 U21210 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18668) );
  NAND2_X1 U21211 ( .A1(n18193), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18469) );
  INV_X1 U21212 ( .A(n18469), .ZN(n18424) );
  NAND2_X1 U21213 ( .A1(n18544), .A2(n18424), .ZN(n18492) );
  INV_X1 U21214 ( .A(n18492), .ZN(n18471) );
  NAND2_X1 U21215 ( .A1(n18668), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18348) );
  INV_X1 U21216 ( .A(n18348), .ZN(n18375) );
  NOR2_X1 U21217 ( .A1(n18471), .A2(n18375), .ZN(n18189) );
  OAI22_X1 U21218 ( .A1(n18190), .A2(n18668), .B1(n18189), .B2(n18188), .ZN(
        P3_U2866) );
  NOR2_X1 U21219 ( .A1(n18192), .A2(n18191), .ZN(P3_U2867) );
  NAND2_X1 U21220 ( .A1(n18639), .A2(n18638), .ZN(n18306) );
  INV_X1 U21221 ( .A(n18306), .ZN(n18642) );
  NAND2_X1 U21222 ( .A1(n18193), .A2(n18668), .ZN(n18283) );
  INV_X1 U21223 ( .A(n18283), .ZN(n18285) );
  NAND2_X1 U21224 ( .A1(n18642), .A2(n18285), .ZN(n18260) );
  NOR2_X1 U21225 ( .A1(n18195), .A2(n18194), .ZN(n18234) );
  NAND2_X1 U21226 ( .A1(n18234), .A2(n18196), .ZN(n18575) );
  INV_X1 U21227 ( .A(BUF2_REG_24__SCAN_IN), .ZN(n18197) );
  NOR2_X2 U21228 ( .A1(n18197), .A2(n18397), .ZN(n18572) );
  NAND2_X1 U21229 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18201) );
  NOR2_X1 U21230 ( .A1(n18201), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18570) );
  NAND2_X1 U21231 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18570), .ZN(
        n18540) );
  INV_X1 U21232 ( .A(n18540), .ZN(n18612) );
  NOR2_X2 U21233 ( .A1(n18399), .A2(n18198), .ZN(n18566) );
  NOR2_X1 U21234 ( .A1(n18668), .A2(n18373), .ZN(n18569) );
  NAND2_X1 U21235 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18569), .ZN(
        n18622) );
  NAND2_X1 U21236 ( .A1(n18622), .A2(n18260), .ZN(n18200) );
  INV_X1 U21237 ( .A(n18200), .ZN(n18261) );
  NOR2_X1 U21238 ( .A1(n18518), .A2(n18261), .ZN(n18236) );
  AOI22_X1 U21239 ( .A1(n18572), .A2(n18612), .B1(n18566), .B2(n18236), .ZN(
        n18203) );
  NAND2_X1 U21240 ( .A1(n18638), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18445) );
  INV_X1 U21241 ( .A(n18445), .ZN(n18199) );
  NOR2_X1 U21242 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18638), .ZN(
        n18421) );
  NOR2_X1 U21243 ( .A1(n18199), .A2(n18421), .ZN(n18493) );
  NOR2_X1 U21244 ( .A1(n18493), .A2(n18201), .ZN(n18545) );
  AOI21_X1 U21245 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n18399), .ZN(n18542) );
  AOI22_X1 U21246 ( .A1(n18571), .A2(n18545), .B1(n18542), .B2(n18200), .ZN(
        n18238) );
  NOR2_X2 U21247 ( .A1(n18397), .A2(n14995), .ZN(n18567) );
  NOR2_X2 U21248 ( .A1(n18445), .A2(n18201), .ZN(n18541) );
  AOI22_X1 U21249 ( .A1(P3_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n18238), .B1(
        n18567), .B2(n18541), .ZN(n18202) );
  OAI211_X1 U21250 ( .C1(n18260), .C2(n18575), .A(n18203), .B(n18202), .ZN(
        P3_U2868) );
  NAND2_X1 U21251 ( .A1(n18234), .A2(n18204), .ZN(n18581) );
  AND2_X1 U21252 ( .A1(n18495), .A2(BUF2_REG_1__SCAN_IN), .ZN(n18577) );
  NOR2_X2 U21253 ( .A1(n18397), .A2(n19221), .ZN(n18576) );
  AOI22_X1 U21254 ( .A1(n18577), .A2(n18236), .B1(n18576), .B2(n18541), .ZN(
        n18207) );
  INV_X1 U21255 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18205) );
  NOR2_X2 U21256 ( .A1(n18205), .A2(n18397), .ZN(n18578) );
  AOI22_X1 U21257 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n18238), .B1(
        n18578), .B2(n18612), .ZN(n18206) );
  OAI211_X1 U21258 ( .C1(n18260), .C2(n18581), .A(n18207), .B(n18206), .ZN(
        P3_U2869) );
  NAND2_X1 U21259 ( .A1(n18234), .A2(n18208), .ZN(n18587) );
  AND2_X1 U21260 ( .A1(n18571), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18584) );
  NOR2_X2 U21261 ( .A1(n18399), .A2(n18209), .ZN(n18583) );
  AOI22_X1 U21262 ( .A1(n18584), .A2(n18541), .B1(n18583), .B2(n18236), .ZN(
        n18212) );
  INV_X1 U21263 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n18210) );
  NOR2_X2 U21264 ( .A1(n18210), .A2(n18397), .ZN(n18582) );
  AOI22_X1 U21265 ( .A1(P3_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n18238), .B1(
        n18582), .B2(n18612), .ZN(n18211) );
  OAI211_X1 U21266 ( .C1(n18260), .C2(n18587), .A(n18212), .B(n18211), .ZN(
        P3_U2870) );
  NAND2_X1 U21267 ( .A1(n18234), .A2(n18213), .ZN(n18593) );
  NOR2_X2 U21268 ( .A1(n18399), .A2(n18214), .ZN(n18588) );
  AND2_X1 U21269 ( .A1(n18571), .A2(BUF2_REG_19__SCAN_IN), .ZN(n18590) );
  AOI22_X1 U21270 ( .A1(n18588), .A2(n18236), .B1(n18590), .B2(n18541), .ZN(
        n18217) );
  NOR2_X2 U21271 ( .A1(n18215), .A2(n18397), .ZN(n18589) );
  AOI22_X1 U21272 ( .A1(P3_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n18238), .B1(
        n18589), .B2(n18612), .ZN(n18216) );
  OAI211_X1 U21273 ( .C1(n18260), .C2(n18593), .A(n18217), .B(n18216), .ZN(
        P3_U2871) );
  NAND2_X1 U21274 ( .A1(n18234), .A2(n18218), .ZN(n18599) );
  NOR2_X2 U21275 ( .A1(n18219), .A2(n18397), .ZN(n18596) );
  NOR2_X2 U21276 ( .A1(n18399), .A2(n18220), .ZN(n18594) );
  AOI22_X1 U21277 ( .A1(n18596), .A2(n18612), .B1(n18594), .B2(n18236), .ZN(
        n18222) );
  AND2_X1 U21278 ( .A1(n18571), .A2(BUF2_REG_20__SCAN_IN), .ZN(n18595) );
  AOI22_X1 U21279 ( .A1(P3_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n18238), .B1(
        n18595), .B2(n18541), .ZN(n18221) );
  OAI211_X1 U21280 ( .C1(n18260), .C2(n18599), .A(n18222), .B(n18221), .ZN(
        P3_U2872) );
  NAND2_X1 U21281 ( .A1(n18234), .A2(n18223), .ZN(n18605) );
  NOR2_X2 U21282 ( .A1(n18399), .A2(n18224), .ZN(n18601) );
  NOR2_X2 U21283 ( .A1(n18225), .A2(n18397), .ZN(n18600) );
  AOI22_X1 U21284 ( .A1(n18601), .A2(n18236), .B1(n18600), .B2(n18612), .ZN(
        n18227) );
  NOR2_X2 U21285 ( .A1(n18397), .A2(n19237), .ZN(n18602) );
  AOI22_X1 U21286 ( .A1(P3_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n18238), .B1(
        n18602), .B2(n18541), .ZN(n18226) );
  OAI211_X1 U21287 ( .C1(n18260), .C2(n18605), .A(n18227), .B(n18226), .ZN(
        P3_U2873) );
  NAND2_X1 U21288 ( .A1(n18234), .A2(n18228), .ZN(n18611) );
  NOR2_X2 U21289 ( .A1(n18229), .A2(n18397), .ZN(n18607) );
  NOR2_X2 U21290 ( .A1(n18399), .A2(n18230), .ZN(n18606) );
  AOI22_X1 U21291 ( .A1(n18607), .A2(n18612), .B1(n18606), .B2(n18236), .ZN(
        n18232) );
  NOR2_X2 U21292 ( .A1(n18397), .A2(n19243), .ZN(n18608) );
  AOI22_X1 U21293 ( .A1(P3_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n18238), .B1(
        n18608), .B2(n18541), .ZN(n18231) );
  OAI211_X1 U21294 ( .C1(n18260), .C2(n18611), .A(n18232), .B(n18231), .ZN(
        P3_U2874) );
  NAND2_X1 U21295 ( .A1(n18234), .A2(n18233), .ZN(n18621) );
  NOR2_X2 U21296 ( .A1(n18235), .A2(n18399), .ZN(n18615) );
  AND2_X1 U21297 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n18571), .ZN(n18613) );
  AOI22_X1 U21298 ( .A1(n18615), .A2(n18236), .B1(n18613), .B2(n18541), .ZN(
        n18240) );
  NOR2_X2 U21299 ( .A1(n18397), .A2(n18237), .ZN(n18617) );
  AOI22_X1 U21300 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n18238), .B1(
        n18617), .B2(n18612), .ZN(n18239) );
  OAI211_X1 U21301 ( .C1(n18260), .C2(n18621), .A(n18240), .B(n18239), .ZN(
        P3_U2875) );
  NAND2_X1 U21302 ( .A1(n18285), .A2(n18421), .ZN(n18286) );
  INV_X1 U21303 ( .A(n18622), .ZN(n18278) );
  NAND2_X1 U21304 ( .A1(n18639), .A2(n18686), .ZN(n18422) );
  NOR2_X1 U21305 ( .A1(n18283), .A2(n18422), .ZN(n18256) );
  AOI22_X1 U21306 ( .A1(n18278), .A2(n18567), .B1(n18566), .B2(n18256), .ZN(
        n18243) );
  INV_X1 U21307 ( .A(n18470), .ZN(n18241) );
  NOR2_X1 U21308 ( .A1(n18399), .A2(n18241), .ZN(n18568) );
  INV_X1 U21309 ( .A(n18568), .ZN(n18284) );
  NOR2_X1 U21310 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18284), .ZN(
        n18423) );
  AOI22_X1 U21311 ( .A1(n18571), .A2(n18569), .B1(n18285), .B2(n18423), .ZN(
        n18257) );
  AOI22_X1 U21312 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18257), .B1(
        n18572), .B2(n18541), .ZN(n18242) );
  OAI211_X1 U21313 ( .C1(n18286), .C2(n18575), .A(n18243), .B(n18242), .ZN(
        P3_U2876) );
  AOI22_X1 U21314 ( .A1(n18278), .A2(n18576), .B1(n18577), .B2(n18256), .ZN(
        n18245) );
  AOI22_X1 U21315 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18257), .B1(
        n18578), .B2(n18541), .ZN(n18244) );
  OAI211_X1 U21316 ( .C1(n18286), .C2(n18581), .A(n18245), .B(n18244), .ZN(
        P3_U2877) );
  AOI22_X1 U21317 ( .A1(n18583), .A2(n18256), .B1(n18582), .B2(n18541), .ZN(
        n18247) );
  AOI22_X1 U21318 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18257), .B1(
        n18278), .B2(n18584), .ZN(n18246) );
  OAI211_X1 U21319 ( .C1(n18286), .C2(n18587), .A(n18247), .B(n18246), .ZN(
        P3_U2878) );
  AOI22_X1 U21320 ( .A1(n18589), .A2(n18541), .B1(n18588), .B2(n18256), .ZN(
        n18249) );
  AOI22_X1 U21321 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18257), .B1(
        n18278), .B2(n18590), .ZN(n18248) );
  OAI211_X1 U21322 ( .C1(n18286), .C2(n18593), .A(n18249), .B(n18248), .ZN(
        P3_U2879) );
  AOI22_X1 U21323 ( .A1(n18596), .A2(n18541), .B1(n18594), .B2(n18256), .ZN(
        n18251) );
  AOI22_X1 U21324 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18257), .B1(
        n18278), .B2(n18595), .ZN(n18250) );
  OAI211_X1 U21325 ( .C1(n18286), .C2(n18599), .A(n18251), .B(n18250), .ZN(
        P3_U2880) );
  AOI22_X1 U21326 ( .A1(n18601), .A2(n18256), .B1(n18600), .B2(n18541), .ZN(
        n18253) );
  AOI22_X1 U21327 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18257), .B1(
        n18278), .B2(n18602), .ZN(n18252) );
  OAI211_X1 U21328 ( .C1(n18286), .C2(n18605), .A(n18253), .B(n18252), .ZN(
        P3_U2881) );
  AOI22_X1 U21329 ( .A1(n18278), .A2(n18608), .B1(n18606), .B2(n18256), .ZN(
        n18255) );
  AOI22_X1 U21330 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18257), .B1(
        n18607), .B2(n18541), .ZN(n18254) );
  OAI211_X1 U21331 ( .C1(n18286), .C2(n18611), .A(n18255), .B(n18254), .ZN(
        P3_U2882) );
  AOI22_X1 U21332 ( .A1(n18278), .A2(n18613), .B1(n18615), .B2(n18256), .ZN(
        n18259) );
  AOI22_X1 U21333 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18257), .B1(
        n18617), .B2(n18541), .ZN(n18258) );
  OAI211_X1 U21334 ( .C1(n18286), .C2(n18621), .A(n18259), .B(n18258), .ZN(
        P3_U2883) );
  NOR2_X2 U21335 ( .A1(n18445), .A2(n18283), .ZN(n18344) );
  INV_X1 U21336 ( .A(n18344), .ZN(n18282) );
  INV_X1 U21337 ( .A(n18260), .ZN(n18302) );
  AOI21_X1 U21338 ( .B1(n18282), .B2(n18286), .A(n18518), .ZN(n18277) );
  AOI22_X1 U21339 ( .A1(n18302), .A2(n18567), .B1(n18566), .B2(n18277), .ZN(
        n18264) );
  AOI221_X1 U21340 ( .B1(n18261), .B2(n18286), .C1(n18446), .C2(n18286), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18262) );
  OAI21_X1 U21341 ( .B1(n18344), .B2(n18262), .A(n18495), .ZN(n18279) );
  AOI22_X1 U21342 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18279), .B1(
        n18278), .B2(n18572), .ZN(n18263) );
  OAI211_X1 U21343 ( .C1(n18282), .C2(n18575), .A(n18264), .B(n18263), .ZN(
        P3_U2884) );
  AOI22_X1 U21344 ( .A1(n18302), .A2(n18576), .B1(n18277), .B2(n18577), .ZN(
        n18266) );
  AOI22_X1 U21345 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18279), .B1(
        n18278), .B2(n18578), .ZN(n18265) );
  OAI211_X1 U21346 ( .C1(n18282), .C2(n18581), .A(n18266), .B(n18265), .ZN(
        P3_U2885) );
  AOI22_X1 U21347 ( .A1(n18278), .A2(n18582), .B1(n18277), .B2(n18583), .ZN(
        n18268) );
  AOI22_X1 U21348 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18279), .B1(
        n18302), .B2(n18584), .ZN(n18267) );
  OAI211_X1 U21349 ( .C1(n18282), .C2(n18587), .A(n18268), .B(n18267), .ZN(
        P3_U2886) );
  AOI22_X1 U21350 ( .A1(n18302), .A2(n18590), .B1(n18277), .B2(n18588), .ZN(
        n18270) );
  AOI22_X1 U21351 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18279), .B1(
        n18278), .B2(n18589), .ZN(n18269) );
  OAI211_X1 U21352 ( .C1(n18282), .C2(n18593), .A(n18270), .B(n18269), .ZN(
        P3_U2887) );
  AOI22_X1 U21353 ( .A1(n18302), .A2(n18595), .B1(n18277), .B2(n18594), .ZN(
        n18272) );
  AOI22_X1 U21354 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18279), .B1(
        n18278), .B2(n18596), .ZN(n18271) );
  OAI211_X1 U21355 ( .C1(n18282), .C2(n18599), .A(n18272), .B(n18271), .ZN(
        P3_U2888) );
  AOI22_X1 U21356 ( .A1(n18278), .A2(n18600), .B1(n18277), .B2(n18601), .ZN(
        n18274) );
  AOI22_X1 U21357 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18279), .B1(
        n18302), .B2(n18602), .ZN(n18273) );
  OAI211_X1 U21358 ( .C1(n18282), .C2(n18605), .A(n18274), .B(n18273), .ZN(
        P3_U2889) );
  AOI22_X1 U21359 ( .A1(n18278), .A2(n18607), .B1(n18277), .B2(n18606), .ZN(
        n18276) );
  AOI22_X1 U21360 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18279), .B1(
        n18302), .B2(n18608), .ZN(n18275) );
  OAI211_X1 U21361 ( .C1(n18282), .C2(n18611), .A(n18276), .B(n18275), .ZN(
        P3_U2890) );
  AOI22_X1 U21362 ( .A1(n18302), .A2(n18613), .B1(n18277), .B2(n18615), .ZN(
        n18281) );
  AOI22_X1 U21363 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18279), .B1(
        n18278), .B2(n18617), .ZN(n18280) );
  OAI211_X1 U21364 ( .C1(n18282), .C2(n18621), .A(n18281), .B(n18280), .ZN(
        P3_U2891) );
  NOR2_X1 U21365 ( .A1(n18639), .A2(n18283), .ZN(n18328) );
  NAND2_X1 U21366 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18328), .ZN(
        n18350) );
  AOI21_X1 U21367 ( .B1(n18639), .B2(n18446), .A(n18284), .ZN(n18374) );
  NAND2_X1 U21368 ( .A1(n18285), .A2(n18374), .ZN(n18303) );
  AND2_X1 U21369 ( .A1(n18686), .A2(n18328), .ZN(n18301) );
  AOI22_X1 U21370 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18303), .B1(
        n18566), .B2(n18301), .ZN(n18288) );
  INV_X1 U21371 ( .A(n18286), .ZN(n18324) );
  AOI22_X1 U21372 ( .A1(n18572), .A2(n18302), .B1(n18324), .B2(n18567), .ZN(
        n18287) );
  OAI211_X1 U21373 ( .C1(n18575), .C2(n18350), .A(n18288), .B(n18287), .ZN(
        P3_U2892) );
  AOI22_X1 U21374 ( .A1(n18302), .A2(n18578), .B1(n18577), .B2(n18301), .ZN(
        n18290) );
  AOI22_X1 U21375 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18303), .B1(
        n18324), .B2(n18576), .ZN(n18289) );
  OAI211_X1 U21376 ( .C1(n18581), .C2(n18350), .A(n18290), .B(n18289), .ZN(
        P3_U2893) );
  AOI22_X1 U21377 ( .A1(n18324), .A2(n18584), .B1(n18583), .B2(n18301), .ZN(
        n18292) );
  AOI22_X1 U21378 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18303), .B1(
        n18302), .B2(n18582), .ZN(n18291) );
  OAI211_X1 U21379 ( .C1(n18587), .C2(n18350), .A(n18292), .B(n18291), .ZN(
        P3_U2894) );
  AOI22_X1 U21380 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18303), .B1(
        n18588), .B2(n18301), .ZN(n18294) );
  AOI22_X1 U21381 ( .A1(n18324), .A2(n18590), .B1(n18302), .B2(n18589), .ZN(
        n18293) );
  OAI211_X1 U21382 ( .C1(n18593), .C2(n18350), .A(n18294), .B(n18293), .ZN(
        P3_U2895) );
  AOI22_X1 U21383 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18303), .B1(
        n18594), .B2(n18301), .ZN(n18296) );
  AOI22_X1 U21384 ( .A1(n18324), .A2(n18595), .B1(n18302), .B2(n18596), .ZN(
        n18295) );
  OAI211_X1 U21385 ( .C1(n18599), .C2(n18350), .A(n18296), .B(n18295), .ZN(
        P3_U2896) );
  AOI22_X1 U21386 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18303), .B1(
        n18601), .B2(n18301), .ZN(n18298) );
  AOI22_X1 U21387 ( .A1(n18324), .A2(n18602), .B1(n18302), .B2(n18600), .ZN(
        n18297) );
  OAI211_X1 U21388 ( .C1(n18605), .C2(n18350), .A(n18298), .B(n18297), .ZN(
        P3_U2897) );
  AOI22_X1 U21389 ( .A1(n18302), .A2(n18607), .B1(n18606), .B2(n18301), .ZN(
        n18300) );
  AOI22_X1 U21390 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18303), .B1(
        n18324), .B2(n18608), .ZN(n18299) );
  OAI211_X1 U21391 ( .C1(n18611), .C2(n18350), .A(n18300), .B(n18299), .ZN(
        P3_U2898) );
  AOI22_X1 U21392 ( .A1(n18324), .A2(n18613), .B1(n18615), .B2(n18301), .ZN(
        n18305) );
  AOI22_X1 U21393 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18303), .B1(
        n18302), .B2(n18617), .ZN(n18304) );
  OAI211_X1 U21394 ( .C1(n18621), .C2(n18350), .A(n18305), .B(n18304), .ZN(
        P3_U2899) );
  NOR2_X2 U21395 ( .A1(n18306), .A2(n18348), .ZN(n18393) );
  INV_X1 U21396 ( .A(n18393), .ZN(n18349) );
  AOI21_X1 U21397 ( .B1(n18350), .B2(n18349), .A(n18518), .ZN(n18323) );
  AOI22_X1 U21398 ( .A1(n18572), .A2(n18324), .B1(n18566), .B2(n18323), .ZN(
        n18310) );
  NOR2_X1 U21399 ( .A1(n18344), .A2(n18324), .ZN(n18307) );
  AOI221_X1 U21400 ( .B1(n18307), .B2(n18350), .C1(n18446), .C2(n18350), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18308) );
  OAI21_X1 U21401 ( .B1(n18393), .B2(n18308), .A(n18495), .ZN(n18325) );
  AOI22_X1 U21402 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18325), .B1(
        n18344), .B2(n18567), .ZN(n18309) );
  OAI211_X1 U21403 ( .C1(n18575), .C2(n18349), .A(n18310), .B(n18309), .ZN(
        P3_U2900) );
  AOI22_X1 U21404 ( .A1(n18344), .A2(n18576), .B1(n18577), .B2(n18323), .ZN(
        n18312) );
  AOI22_X1 U21405 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18325), .B1(
        n18324), .B2(n18578), .ZN(n18311) );
  OAI211_X1 U21406 ( .C1(n18581), .C2(n18349), .A(n18312), .B(n18311), .ZN(
        P3_U2901) );
  AOI22_X1 U21407 ( .A1(n18324), .A2(n18582), .B1(n18583), .B2(n18323), .ZN(
        n18314) );
  AOI22_X1 U21408 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18325), .B1(
        n18344), .B2(n18584), .ZN(n18313) );
  OAI211_X1 U21409 ( .C1(n18587), .C2(n18349), .A(n18314), .B(n18313), .ZN(
        P3_U2902) );
  AOI22_X1 U21410 ( .A1(n18324), .A2(n18589), .B1(n18588), .B2(n18323), .ZN(
        n18316) );
  AOI22_X1 U21411 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18325), .B1(
        n18344), .B2(n18590), .ZN(n18315) );
  OAI211_X1 U21412 ( .C1(n18593), .C2(n18349), .A(n18316), .B(n18315), .ZN(
        P3_U2903) );
  AOI22_X1 U21413 ( .A1(n18344), .A2(n18595), .B1(n18594), .B2(n18323), .ZN(
        n18318) );
  AOI22_X1 U21414 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18325), .B1(
        n18324), .B2(n18596), .ZN(n18317) );
  OAI211_X1 U21415 ( .C1(n18599), .C2(n18349), .A(n18318), .B(n18317), .ZN(
        P3_U2904) );
  AOI22_X1 U21416 ( .A1(n18324), .A2(n18600), .B1(n18601), .B2(n18323), .ZN(
        n18320) );
  AOI22_X1 U21417 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18325), .B1(
        n18344), .B2(n18602), .ZN(n18319) );
  OAI211_X1 U21418 ( .C1(n18605), .C2(n18349), .A(n18320), .B(n18319), .ZN(
        P3_U2905) );
  AOI22_X1 U21419 ( .A1(n18324), .A2(n18607), .B1(n18606), .B2(n18323), .ZN(
        n18322) );
  AOI22_X1 U21420 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18325), .B1(
        n18344), .B2(n18608), .ZN(n18321) );
  OAI211_X1 U21421 ( .C1(n18611), .C2(n18349), .A(n18322), .B(n18321), .ZN(
        P3_U2906) );
  AOI22_X1 U21422 ( .A1(n18324), .A2(n18617), .B1(n18615), .B2(n18323), .ZN(
        n18327) );
  AOI22_X1 U21423 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18325), .B1(
        n18344), .B2(n18613), .ZN(n18326) );
  OAI211_X1 U21424 ( .C1(n18621), .C2(n18349), .A(n18327), .B(n18326), .ZN(
        P3_U2907) );
  NAND2_X1 U21425 ( .A1(n18421), .A2(n18375), .ZN(n18376) );
  NOR2_X1 U21426 ( .A1(n18348), .A2(n18422), .ZN(n18343) );
  AOI22_X1 U21427 ( .A1(n18572), .A2(n18344), .B1(n18566), .B2(n18343), .ZN(
        n18330) );
  AOI22_X1 U21428 ( .A1(n18571), .A2(n18328), .B1(n18375), .B2(n18423), .ZN(
        n18345) );
  INV_X1 U21429 ( .A(n18350), .ZN(n18368) );
  AOI22_X1 U21430 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18345), .B1(
        n18567), .B2(n18368), .ZN(n18329) );
  OAI211_X1 U21431 ( .C1(n18575), .C2(n18376), .A(n18330), .B(n18329), .ZN(
        P3_U2908) );
  AOI22_X1 U21432 ( .A1(n18577), .A2(n18343), .B1(n18576), .B2(n18368), .ZN(
        n18332) );
  AOI22_X1 U21433 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18345), .B1(
        n18344), .B2(n18578), .ZN(n18331) );
  OAI211_X1 U21434 ( .C1(n18581), .C2(n18376), .A(n18332), .B(n18331), .ZN(
        P3_U2909) );
  AOI22_X1 U21435 ( .A1(n18344), .A2(n18582), .B1(n18583), .B2(n18343), .ZN(
        n18334) );
  AOI22_X1 U21436 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18345), .B1(
        n18584), .B2(n18368), .ZN(n18333) );
  OAI211_X1 U21437 ( .C1(n18587), .C2(n18376), .A(n18334), .B(n18333), .ZN(
        P3_U2910) );
  AOI22_X1 U21438 ( .A1(n18588), .A2(n18343), .B1(n18590), .B2(n18368), .ZN(
        n18336) );
  AOI22_X1 U21439 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18345), .B1(
        n18344), .B2(n18589), .ZN(n18335) );
  OAI211_X1 U21440 ( .C1(n18593), .C2(n18376), .A(n18336), .B(n18335), .ZN(
        P3_U2911) );
  AOI22_X1 U21441 ( .A1(n18344), .A2(n18596), .B1(n18594), .B2(n18343), .ZN(
        n18338) );
  AOI22_X1 U21442 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18345), .B1(
        n18595), .B2(n18368), .ZN(n18337) );
  OAI211_X1 U21443 ( .C1(n18599), .C2(n18376), .A(n18338), .B(n18337), .ZN(
        P3_U2912) );
  AOI22_X1 U21444 ( .A1(n18602), .A2(n18368), .B1(n18601), .B2(n18343), .ZN(
        n18340) );
  AOI22_X1 U21445 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18345), .B1(
        n18344), .B2(n18600), .ZN(n18339) );
  OAI211_X1 U21446 ( .C1(n18605), .C2(n18376), .A(n18340), .B(n18339), .ZN(
        P3_U2913) );
  AOI22_X1 U21447 ( .A1(n18608), .A2(n18368), .B1(n18606), .B2(n18343), .ZN(
        n18342) );
  AOI22_X1 U21448 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18345), .B1(
        n18344), .B2(n18607), .ZN(n18341) );
  OAI211_X1 U21449 ( .C1(n18611), .C2(n18376), .A(n18342), .B(n18341), .ZN(
        P3_U2914) );
  AOI22_X1 U21450 ( .A1(n18615), .A2(n18343), .B1(n18613), .B2(n18368), .ZN(
        n18347) );
  AOI22_X1 U21451 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18345), .B1(
        n18344), .B2(n18617), .ZN(n18346) );
  OAI211_X1 U21452 ( .C1(n18621), .C2(n18376), .A(n18347), .B(n18346), .ZN(
        P3_U2915) );
  NOR2_X2 U21453 ( .A1(n18445), .A2(n18348), .ZN(n18441) );
  INV_X1 U21454 ( .A(n18441), .ZN(n18372) );
  NAND2_X1 U21455 ( .A1(n18376), .A2(n18372), .ZN(n18352) );
  INV_X1 U21456 ( .A(n18352), .ZN(n18398) );
  NOR2_X1 U21457 ( .A1(n18518), .A2(n18398), .ZN(n18367) );
  AOI22_X1 U21458 ( .A1(n18567), .A2(n18393), .B1(n18566), .B2(n18367), .ZN(
        n18354) );
  NAND2_X1 U21459 ( .A1(n18350), .A2(n18349), .ZN(n18351) );
  OAI221_X1 U21460 ( .B1(n18352), .B2(n18544), .C1(n18352), .C2(n18351), .A(
        n18542), .ZN(n18369) );
  AOI22_X1 U21461 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18369), .B1(
        n18572), .B2(n18368), .ZN(n18353) );
  OAI211_X1 U21462 ( .C1(n18575), .C2(n18372), .A(n18354), .B(n18353), .ZN(
        P3_U2916) );
  AOI22_X1 U21463 ( .A1(n18578), .A2(n18368), .B1(n18577), .B2(n18367), .ZN(
        n18356) );
  AOI22_X1 U21464 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18369), .B1(
        n18576), .B2(n18393), .ZN(n18355) );
  OAI211_X1 U21465 ( .C1(n18581), .C2(n18372), .A(n18356), .B(n18355), .ZN(
        P3_U2917) );
  AOI22_X1 U21466 ( .A1(n18583), .A2(n18367), .B1(n18582), .B2(n18368), .ZN(
        n18358) );
  AOI22_X1 U21467 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18369), .B1(
        n18584), .B2(n18393), .ZN(n18357) );
  OAI211_X1 U21468 ( .C1(n18587), .C2(n18372), .A(n18358), .B(n18357), .ZN(
        P3_U2918) );
  AOI22_X1 U21469 ( .A1(n18588), .A2(n18367), .B1(n18590), .B2(n18393), .ZN(
        n18360) );
  AOI22_X1 U21470 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18369), .B1(
        n18589), .B2(n18368), .ZN(n18359) );
  OAI211_X1 U21471 ( .C1(n18593), .C2(n18372), .A(n18360), .B(n18359), .ZN(
        P3_U2919) );
  AOI22_X1 U21472 ( .A1(n18596), .A2(n18368), .B1(n18594), .B2(n18367), .ZN(
        n18362) );
  AOI22_X1 U21473 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18369), .B1(
        n18595), .B2(n18393), .ZN(n18361) );
  OAI211_X1 U21474 ( .C1(n18599), .C2(n18372), .A(n18362), .B(n18361), .ZN(
        P3_U2920) );
  AOI22_X1 U21475 ( .A1(n18602), .A2(n18393), .B1(n18601), .B2(n18367), .ZN(
        n18364) );
  AOI22_X1 U21476 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18369), .B1(
        n18600), .B2(n18368), .ZN(n18363) );
  OAI211_X1 U21477 ( .C1(n18605), .C2(n18372), .A(n18364), .B(n18363), .ZN(
        P3_U2921) );
  AOI22_X1 U21478 ( .A1(n18608), .A2(n18393), .B1(n18606), .B2(n18367), .ZN(
        n18366) );
  AOI22_X1 U21479 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18369), .B1(
        n18607), .B2(n18368), .ZN(n18365) );
  OAI211_X1 U21480 ( .C1(n18611), .C2(n18372), .A(n18366), .B(n18365), .ZN(
        P3_U2922) );
  AOI22_X1 U21481 ( .A1(n18615), .A2(n18367), .B1(n18613), .B2(n18393), .ZN(
        n18371) );
  AOI22_X1 U21482 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18369), .B1(
        n18617), .B2(n18368), .ZN(n18370) );
  OAI211_X1 U21483 ( .C1(n18621), .C2(n18372), .A(n18371), .B(n18370), .ZN(
        P3_U2923) );
  NOR2_X1 U21484 ( .A1(n18373), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18425) );
  NAND2_X1 U21485 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18425), .ZN(
        n18396) );
  AND2_X1 U21486 ( .A1(n18686), .A2(n18425), .ZN(n18391) );
  AOI22_X1 U21487 ( .A1(n18572), .A2(n18393), .B1(n18566), .B2(n18391), .ZN(
        n18378) );
  NAND2_X1 U21488 ( .A1(n18375), .A2(n18374), .ZN(n18392) );
  INV_X1 U21489 ( .A(n18376), .ZN(n18416) );
  AOI22_X1 U21490 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18392), .B1(
        n18567), .B2(n18416), .ZN(n18377) );
  OAI211_X1 U21491 ( .C1(n18575), .C2(n18396), .A(n18378), .B(n18377), .ZN(
        P3_U2924) );
  AOI22_X1 U21492 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18392), .B1(
        n18577), .B2(n18391), .ZN(n18380) );
  AOI22_X1 U21493 ( .A1(n18578), .A2(n18393), .B1(n18576), .B2(n18416), .ZN(
        n18379) );
  OAI211_X1 U21494 ( .C1(n18581), .C2(n18396), .A(n18380), .B(n18379), .ZN(
        P3_U2925) );
  AOI22_X1 U21495 ( .A1(n18583), .A2(n18391), .B1(n18582), .B2(n18393), .ZN(
        n18382) );
  AOI22_X1 U21496 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18392), .B1(
        n18584), .B2(n18416), .ZN(n18381) );
  OAI211_X1 U21497 ( .C1(n18587), .C2(n18396), .A(n18382), .B(n18381), .ZN(
        P3_U2926) );
  AOI22_X1 U21498 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18392), .B1(
        n18588), .B2(n18391), .ZN(n18384) );
  AOI22_X1 U21499 ( .A1(n18589), .A2(n18393), .B1(n18590), .B2(n18416), .ZN(
        n18383) );
  OAI211_X1 U21500 ( .C1(n18593), .C2(n18396), .A(n18384), .B(n18383), .ZN(
        P3_U2927) );
  AOI22_X1 U21501 ( .A1(n18596), .A2(n18393), .B1(n18594), .B2(n18391), .ZN(
        n18386) );
  AOI22_X1 U21502 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18392), .B1(
        n18595), .B2(n18416), .ZN(n18385) );
  OAI211_X1 U21503 ( .C1(n18599), .C2(n18396), .A(n18386), .B(n18385), .ZN(
        P3_U2928) );
  AOI22_X1 U21504 ( .A1(n18601), .A2(n18391), .B1(n18600), .B2(n18393), .ZN(
        n18388) );
  AOI22_X1 U21505 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18392), .B1(
        n18602), .B2(n18416), .ZN(n18387) );
  OAI211_X1 U21506 ( .C1(n18605), .C2(n18396), .A(n18388), .B(n18387), .ZN(
        P3_U2929) );
  AOI22_X1 U21507 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18392), .B1(
        n18606), .B2(n18391), .ZN(n18390) );
  AOI22_X1 U21508 ( .A1(n18608), .A2(n18416), .B1(n18607), .B2(n18393), .ZN(
        n18389) );
  OAI211_X1 U21509 ( .C1(n18611), .C2(n18396), .A(n18390), .B(n18389), .ZN(
        P3_U2930) );
  AOI22_X1 U21510 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18392), .B1(
        n18615), .B2(n18391), .ZN(n18395) );
  AOI22_X1 U21511 ( .A1(n18617), .A2(n18393), .B1(n18613), .B2(n18416), .ZN(
        n18394) );
  OAI211_X1 U21512 ( .C1(n18621), .C2(n18396), .A(n18395), .B(n18394), .ZN(
        P3_U2931) );
  NAND2_X1 U21513 ( .A1(n18642), .A2(n18424), .ZN(n18420) );
  INV_X1 U21514 ( .A(n18420), .ZN(n18489) );
  INV_X1 U21515 ( .A(n18396), .ZN(n18464) );
  NOR2_X1 U21516 ( .A1(n18489), .A2(n18464), .ZN(n18447) );
  NOR2_X1 U21517 ( .A1(n18518), .A2(n18447), .ZN(n18415) );
  AOI22_X1 U21518 ( .A1(n18572), .A2(n18416), .B1(n18566), .B2(n18415), .ZN(
        n18402) );
  OAI22_X1 U21519 ( .A1(n18447), .A2(n18399), .B1(n18398), .B2(n18397), .ZN(
        n18400) );
  OAI21_X1 U21520 ( .B1(n18489), .B2(n18782), .A(n18400), .ZN(n18417) );
  AOI22_X1 U21521 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18417), .B1(
        n18567), .B2(n18441), .ZN(n18401) );
  OAI211_X1 U21522 ( .C1(n18575), .C2(n18420), .A(n18402), .B(n18401), .ZN(
        P3_U2932) );
  AOI22_X1 U21523 ( .A1(n18578), .A2(n18416), .B1(n18577), .B2(n18415), .ZN(
        n18404) );
  AOI22_X1 U21524 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18417), .B1(
        n18576), .B2(n18441), .ZN(n18403) );
  OAI211_X1 U21525 ( .C1(n18581), .C2(n18420), .A(n18404), .B(n18403), .ZN(
        P3_U2933) );
  AOI22_X1 U21526 ( .A1(n18583), .A2(n18415), .B1(n18582), .B2(n18416), .ZN(
        n18406) );
  AOI22_X1 U21527 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18417), .B1(
        n18584), .B2(n18441), .ZN(n18405) );
  OAI211_X1 U21528 ( .C1(n18587), .C2(n18420), .A(n18406), .B(n18405), .ZN(
        P3_U2934) );
  AOI22_X1 U21529 ( .A1(n18589), .A2(n18416), .B1(n18588), .B2(n18415), .ZN(
        n18408) );
  AOI22_X1 U21530 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18417), .B1(
        n18590), .B2(n18441), .ZN(n18407) );
  OAI211_X1 U21531 ( .C1(n18593), .C2(n18420), .A(n18408), .B(n18407), .ZN(
        P3_U2935) );
  AOI22_X1 U21532 ( .A1(n18596), .A2(n18416), .B1(n18594), .B2(n18415), .ZN(
        n18410) );
  AOI22_X1 U21533 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18417), .B1(
        n18595), .B2(n18441), .ZN(n18409) );
  OAI211_X1 U21534 ( .C1(n18599), .C2(n18420), .A(n18410), .B(n18409), .ZN(
        P3_U2936) );
  AOI22_X1 U21535 ( .A1(n18602), .A2(n18441), .B1(n18601), .B2(n18415), .ZN(
        n18412) );
  AOI22_X1 U21536 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18417), .B1(
        n18600), .B2(n18416), .ZN(n18411) );
  OAI211_X1 U21537 ( .C1(n18605), .C2(n18420), .A(n18412), .B(n18411), .ZN(
        P3_U2937) );
  AOI22_X1 U21538 ( .A1(n18608), .A2(n18441), .B1(n18606), .B2(n18415), .ZN(
        n18414) );
  AOI22_X1 U21539 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18417), .B1(
        n18607), .B2(n18416), .ZN(n18413) );
  OAI211_X1 U21540 ( .C1(n18611), .C2(n18420), .A(n18414), .B(n18413), .ZN(
        P3_U2938) );
  AOI22_X1 U21541 ( .A1(n18617), .A2(n18416), .B1(n18615), .B2(n18415), .ZN(
        n18419) );
  AOI22_X1 U21542 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18417), .B1(
        n18613), .B2(n18441), .ZN(n18418) );
  OAI211_X1 U21543 ( .C1(n18621), .C2(n18420), .A(n18419), .B(n18418), .ZN(
        P3_U2939) );
  NAND2_X1 U21544 ( .A1(n18421), .A2(n18424), .ZN(n18472) );
  NOR2_X1 U21545 ( .A1(n18469), .A2(n18422), .ZN(n18440) );
  AOI22_X1 U21546 ( .A1(n18567), .A2(n18464), .B1(n18566), .B2(n18440), .ZN(
        n18427) );
  AOI22_X1 U21547 ( .A1(n18571), .A2(n18425), .B1(n18424), .B2(n18423), .ZN(
        n18442) );
  AOI22_X1 U21548 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18442), .B1(
        n18572), .B2(n18441), .ZN(n18426) );
  OAI211_X1 U21549 ( .C1(n18575), .C2(n18472), .A(n18427), .B(n18426), .ZN(
        P3_U2940) );
  AOI22_X1 U21550 ( .A1(n18577), .A2(n18440), .B1(n18576), .B2(n18464), .ZN(
        n18429) );
  AOI22_X1 U21551 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18442), .B1(
        n18578), .B2(n18441), .ZN(n18428) );
  OAI211_X1 U21552 ( .C1(n18581), .C2(n18472), .A(n18429), .B(n18428), .ZN(
        P3_U2941) );
  AOI22_X1 U21553 ( .A1(n18583), .A2(n18440), .B1(n18582), .B2(n18441), .ZN(
        n18431) );
  AOI22_X1 U21554 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18442), .B1(
        n18584), .B2(n18464), .ZN(n18430) );
  OAI211_X1 U21555 ( .C1(n18587), .C2(n18472), .A(n18431), .B(n18430), .ZN(
        P3_U2942) );
  AOI22_X1 U21556 ( .A1(n18589), .A2(n18441), .B1(n18588), .B2(n18440), .ZN(
        n18433) );
  AOI22_X1 U21557 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18442), .B1(
        n18590), .B2(n18464), .ZN(n18432) );
  OAI211_X1 U21558 ( .C1(n18593), .C2(n18472), .A(n18433), .B(n18432), .ZN(
        P3_U2943) );
  AOI22_X1 U21559 ( .A1(n18595), .A2(n18464), .B1(n18594), .B2(n18440), .ZN(
        n18435) );
  AOI22_X1 U21560 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18442), .B1(
        n18596), .B2(n18441), .ZN(n18434) );
  OAI211_X1 U21561 ( .C1(n18599), .C2(n18472), .A(n18435), .B(n18434), .ZN(
        P3_U2944) );
  AOI22_X1 U21562 ( .A1(n18602), .A2(n18464), .B1(n18601), .B2(n18440), .ZN(
        n18437) );
  AOI22_X1 U21563 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18442), .B1(
        n18600), .B2(n18441), .ZN(n18436) );
  OAI211_X1 U21564 ( .C1(n18605), .C2(n18472), .A(n18437), .B(n18436), .ZN(
        P3_U2945) );
  AOI22_X1 U21565 ( .A1(n18608), .A2(n18464), .B1(n18606), .B2(n18440), .ZN(
        n18439) );
  AOI22_X1 U21566 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18442), .B1(
        n18607), .B2(n18441), .ZN(n18438) );
  OAI211_X1 U21567 ( .C1(n18611), .C2(n18472), .A(n18439), .B(n18438), .ZN(
        P3_U2946) );
  AOI22_X1 U21568 ( .A1(n18615), .A2(n18440), .B1(n18613), .B2(n18464), .ZN(
        n18444) );
  AOI22_X1 U21569 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18442), .B1(
        n18617), .B2(n18441), .ZN(n18443) );
  OAI211_X1 U21570 ( .C1(n18621), .C2(n18472), .A(n18444), .B(n18443), .ZN(
        P3_U2947) );
  NOR2_X2 U21571 ( .A1(n18445), .A2(n18469), .ZN(n18536) );
  INV_X1 U21572 ( .A(n18536), .ZN(n18468) );
  AOI22_X1 U21573 ( .A1(n18567), .A2(n18489), .B1(n18566), .B2(n18463), .ZN(
        n18450) );
  AOI221_X1 U21574 ( .B1(n18447), .B2(n18472), .C1(n18446), .C2(n18472), .A(
        P3_STATE2_REG_3__SCAN_IN), .ZN(n18448) );
  OAI21_X1 U21575 ( .B1(n18536), .B2(n18448), .A(n18495), .ZN(n18465) );
  AOI22_X1 U21576 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18465), .B1(
        n18572), .B2(n18464), .ZN(n18449) );
  OAI211_X1 U21577 ( .C1(n18575), .C2(n18468), .A(n18450), .B(n18449), .ZN(
        P3_U2948) );
  AOI22_X1 U21578 ( .A1(n18577), .A2(n18463), .B1(n18576), .B2(n18489), .ZN(
        n18452) );
  AOI22_X1 U21579 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18465), .B1(
        n18578), .B2(n18464), .ZN(n18451) );
  OAI211_X1 U21580 ( .C1(n18581), .C2(n18468), .A(n18452), .B(n18451), .ZN(
        P3_U2949) );
  AOI22_X1 U21581 ( .A1(n18583), .A2(n18463), .B1(n18582), .B2(n18464), .ZN(
        n18454) );
  AOI22_X1 U21582 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18465), .B1(
        n18584), .B2(n18489), .ZN(n18453) );
  OAI211_X1 U21583 ( .C1(n18587), .C2(n18468), .A(n18454), .B(n18453), .ZN(
        P3_U2950) );
  AOI22_X1 U21584 ( .A1(n18589), .A2(n18464), .B1(n18588), .B2(n18463), .ZN(
        n18456) );
  AOI22_X1 U21585 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18465), .B1(
        n18590), .B2(n18489), .ZN(n18455) );
  OAI211_X1 U21586 ( .C1(n18593), .C2(n18468), .A(n18456), .B(n18455), .ZN(
        P3_U2951) );
  AOI22_X1 U21587 ( .A1(n18595), .A2(n18489), .B1(n18594), .B2(n18463), .ZN(
        n18458) );
  AOI22_X1 U21588 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18465), .B1(
        n18596), .B2(n18464), .ZN(n18457) );
  OAI211_X1 U21589 ( .C1(n18599), .C2(n18468), .A(n18458), .B(n18457), .ZN(
        P3_U2952) );
  AOI22_X1 U21590 ( .A1(n18601), .A2(n18463), .B1(n18600), .B2(n18464), .ZN(
        n18460) );
  AOI22_X1 U21591 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18465), .B1(
        n18602), .B2(n18489), .ZN(n18459) );
  OAI211_X1 U21592 ( .C1(n18605), .C2(n18468), .A(n18460), .B(n18459), .ZN(
        P3_U2953) );
  AOI22_X1 U21593 ( .A1(n18607), .A2(n18464), .B1(n18606), .B2(n18463), .ZN(
        n18462) );
  AOI22_X1 U21594 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18465), .B1(
        n18608), .B2(n18489), .ZN(n18461) );
  OAI211_X1 U21595 ( .C1(n18611), .C2(n18468), .A(n18462), .B(n18461), .ZN(
        P3_U2954) );
  AOI22_X1 U21596 ( .A1(n18615), .A2(n18463), .B1(n18613), .B2(n18489), .ZN(
        n18467) );
  AOI22_X1 U21597 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18465), .B1(
        n18617), .B2(n18464), .ZN(n18466) );
  OAI211_X1 U21598 ( .C1(n18621), .C2(n18468), .A(n18467), .B(n18466), .ZN(
        P3_U2955) );
  NOR2_X1 U21599 ( .A1(n18639), .A2(n18469), .ZN(n18519) );
  NAND2_X1 U21600 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18519), .ZN(
        n18520) );
  OAI211_X1 U21601 ( .C1(n18471), .C2(n18519), .A(n18470), .B(n18495), .ZN(
        n18488) );
  AND2_X1 U21602 ( .A1(n18686), .A2(n18519), .ZN(n18487) );
  AOI22_X1 U21603 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18488), .B1(
        n18566), .B2(n18487), .ZN(n18474) );
  INV_X1 U21604 ( .A(n18472), .ZN(n18512) );
  AOI22_X1 U21605 ( .A1(n18572), .A2(n18489), .B1(n18567), .B2(n18512), .ZN(
        n18473) );
  OAI211_X1 U21606 ( .C1(n18575), .C2(n18520), .A(n18474), .B(n18473), .ZN(
        P3_U2956) );
  AOI22_X1 U21607 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18488), .B1(
        n18577), .B2(n18487), .ZN(n18476) );
  AOI22_X1 U21608 ( .A1(n18578), .A2(n18489), .B1(n18576), .B2(n18512), .ZN(
        n18475) );
  OAI211_X1 U21609 ( .C1(n18581), .C2(n18520), .A(n18476), .B(n18475), .ZN(
        P3_U2957) );
  AOI22_X1 U21610 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18488), .B1(
        n18583), .B2(n18487), .ZN(n18478) );
  AOI22_X1 U21611 ( .A1(n18584), .A2(n18512), .B1(n18582), .B2(n18489), .ZN(
        n18477) );
  OAI211_X1 U21612 ( .C1(n18587), .C2(n18520), .A(n18478), .B(n18477), .ZN(
        P3_U2958) );
  AOI22_X1 U21613 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18488), .B1(
        n18588), .B2(n18487), .ZN(n18480) );
  AOI22_X1 U21614 ( .A1(n18589), .A2(n18489), .B1(n18590), .B2(n18512), .ZN(
        n18479) );
  OAI211_X1 U21615 ( .C1(n18593), .C2(n18520), .A(n18480), .B(n18479), .ZN(
        P3_U2959) );
  AOI22_X1 U21616 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18488), .B1(
        n18594), .B2(n18487), .ZN(n18482) );
  AOI22_X1 U21617 ( .A1(n18596), .A2(n18489), .B1(n18595), .B2(n18512), .ZN(
        n18481) );
  OAI211_X1 U21618 ( .C1(n18599), .C2(n18520), .A(n18482), .B(n18481), .ZN(
        P3_U2960) );
  AOI22_X1 U21619 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18488), .B1(
        n18601), .B2(n18487), .ZN(n18484) );
  AOI22_X1 U21620 ( .A1(n18602), .A2(n18512), .B1(n18600), .B2(n18489), .ZN(
        n18483) );
  OAI211_X1 U21621 ( .C1(n18605), .C2(n18520), .A(n18484), .B(n18483), .ZN(
        P3_U2961) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18488), .B1(
        n18606), .B2(n18487), .ZN(n18486) );
  AOI22_X1 U21623 ( .A1(n18608), .A2(n18512), .B1(n18607), .B2(n18489), .ZN(
        n18485) );
  OAI211_X1 U21624 ( .C1(n18611), .C2(n18520), .A(n18486), .B(n18485), .ZN(
        P3_U2962) );
  AOI22_X1 U21625 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18488), .B1(
        n18615), .B2(n18487), .ZN(n18491) );
  AOI22_X1 U21626 ( .A1(n18617), .A2(n18489), .B1(n18613), .B2(n18512), .ZN(
        n18490) );
  OAI211_X1 U21627 ( .C1(n18621), .C2(n18520), .A(n18491), .B(n18490), .ZN(
        P3_U2963) );
  INV_X1 U21628 ( .A(n18570), .ZN(n18517) );
  NOR2_X2 U21629 ( .A1(n18517), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18616) );
  INV_X1 U21630 ( .A(n18616), .ZN(n18516) );
  NAND2_X1 U21631 ( .A1(n18520), .A2(n18516), .ZN(n18543) );
  INV_X1 U21632 ( .A(n18543), .ZN(n18496) );
  OAI21_X1 U21633 ( .B1(n18493), .B2(n18492), .A(n18496), .ZN(n18494) );
  OAI211_X1 U21634 ( .C1(n18616), .C2(n18782), .A(n18495), .B(n18494), .ZN(
        n18513) );
  NOR2_X1 U21635 ( .A1(n18518), .A2(n18496), .ZN(n18511) );
  AOI22_X1 U21636 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18513), .B1(
        n18566), .B2(n18511), .ZN(n18498) );
  AOI22_X1 U21637 ( .A1(n18572), .A2(n18512), .B1(n18567), .B2(n18536), .ZN(
        n18497) );
  OAI211_X1 U21638 ( .C1(n18575), .C2(n18516), .A(n18498), .B(n18497), .ZN(
        P3_U2964) );
  AOI22_X1 U21639 ( .A1(n18577), .A2(n18511), .B1(n18576), .B2(n18536), .ZN(
        n18500) );
  AOI22_X1 U21640 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18513), .B1(
        n18578), .B2(n18512), .ZN(n18499) );
  OAI211_X1 U21641 ( .C1(n18581), .C2(n18516), .A(n18500), .B(n18499), .ZN(
        P3_U2965) );
  AOI22_X1 U21642 ( .A1(n18583), .A2(n18511), .B1(n18582), .B2(n18512), .ZN(
        n18502) );
  AOI22_X1 U21643 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18513), .B1(
        n18584), .B2(n18536), .ZN(n18501) );
  OAI211_X1 U21644 ( .C1(n18587), .C2(n18516), .A(n18502), .B(n18501), .ZN(
        P3_U2966) );
  AOI22_X1 U21645 ( .A1(n18589), .A2(n18512), .B1(n18588), .B2(n18511), .ZN(
        n18504) );
  AOI22_X1 U21646 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18513), .B1(
        n18590), .B2(n18536), .ZN(n18503) );
  OAI211_X1 U21647 ( .C1(n18593), .C2(n18516), .A(n18504), .B(n18503), .ZN(
        P3_U2967) );
  AOI22_X1 U21648 ( .A1(n18595), .A2(n18536), .B1(n18594), .B2(n18511), .ZN(
        n18506) );
  AOI22_X1 U21649 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18513), .B1(
        n18596), .B2(n18512), .ZN(n18505) );
  OAI211_X1 U21650 ( .C1(n18599), .C2(n18516), .A(n18506), .B(n18505), .ZN(
        P3_U2968) );
  AOI22_X1 U21651 ( .A1(n18601), .A2(n18511), .B1(n18600), .B2(n18512), .ZN(
        n18508) );
  AOI22_X1 U21652 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18513), .B1(
        n18602), .B2(n18536), .ZN(n18507) );
  OAI211_X1 U21653 ( .C1(n18605), .C2(n18516), .A(n18508), .B(n18507), .ZN(
        P3_U2969) );
  AOI22_X1 U21654 ( .A1(n18608), .A2(n18536), .B1(n18606), .B2(n18511), .ZN(
        n18510) );
  AOI22_X1 U21655 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18513), .B1(
        n18607), .B2(n18512), .ZN(n18509) );
  OAI211_X1 U21656 ( .C1(n18611), .C2(n18516), .A(n18510), .B(n18509), .ZN(
        P3_U2970) );
  AOI22_X1 U21657 ( .A1(n18617), .A2(n18512), .B1(n18615), .B2(n18511), .ZN(
        n18515) );
  AOI22_X1 U21658 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18513), .B1(
        n18613), .B2(n18536), .ZN(n18514) );
  OAI211_X1 U21659 ( .C1(n18621), .C2(n18516), .A(n18515), .B(n18514), .ZN(
        P3_U2971) );
  NOR2_X1 U21660 ( .A1(n18518), .A2(n18517), .ZN(n18535) );
  AOI22_X1 U21661 ( .A1(n18572), .A2(n18536), .B1(n18566), .B2(n18535), .ZN(
        n18522) );
  AOI22_X1 U21662 ( .A1(n18571), .A2(n18519), .B1(n18570), .B2(n18568), .ZN(
        n18537) );
  INV_X1 U21663 ( .A(n18520), .ZN(n18561) );
  AOI22_X1 U21664 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18537), .B1(
        n18567), .B2(n18561), .ZN(n18521) );
  OAI211_X1 U21665 ( .C1(n18575), .C2(n18540), .A(n18522), .B(n18521), .ZN(
        P3_U2972) );
  AOI22_X1 U21666 ( .A1(n18578), .A2(n18536), .B1(n18577), .B2(n18535), .ZN(
        n18524) );
  AOI22_X1 U21667 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18537), .B1(
        n18576), .B2(n18561), .ZN(n18523) );
  OAI211_X1 U21668 ( .C1(n18581), .C2(n18540), .A(n18524), .B(n18523), .ZN(
        P3_U2973) );
  AOI22_X1 U21669 ( .A1(n18584), .A2(n18561), .B1(n18583), .B2(n18535), .ZN(
        n18526) );
  AOI22_X1 U21670 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18537), .B1(
        n18582), .B2(n18536), .ZN(n18525) );
  OAI211_X1 U21671 ( .C1(n18587), .C2(n18540), .A(n18526), .B(n18525), .ZN(
        P3_U2974) );
  AOI22_X1 U21672 ( .A1(n18589), .A2(n18536), .B1(n18588), .B2(n18535), .ZN(
        n18528) );
  AOI22_X1 U21673 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18537), .B1(
        n18590), .B2(n18561), .ZN(n18527) );
  OAI211_X1 U21674 ( .C1(n18593), .C2(n18540), .A(n18528), .B(n18527), .ZN(
        P3_U2975) );
  AOI22_X1 U21675 ( .A1(n18595), .A2(n18561), .B1(n18594), .B2(n18535), .ZN(
        n18530) );
  AOI22_X1 U21676 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18537), .B1(
        n18596), .B2(n18536), .ZN(n18529) );
  OAI211_X1 U21677 ( .C1(n18599), .C2(n18540), .A(n18530), .B(n18529), .ZN(
        P3_U2976) );
  AOI22_X1 U21678 ( .A1(n18601), .A2(n18535), .B1(n18600), .B2(n18536), .ZN(
        n18532) );
  AOI22_X1 U21679 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18537), .B1(
        n18602), .B2(n18561), .ZN(n18531) );
  OAI211_X1 U21680 ( .C1(n18605), .C2(n18540), .A(n18532), .B(n18531), .ZN(
        P3_U2977) );
  AOI22_X1 U21681 ( .A1(n18607), .A2(n18536), .B1(n18606), .B2(n18535), .ZN(
        n18534) );
  AOI22_X1 U21682 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18537), .B1(
        n18608), .B2(n18561), .ZN(n18533) );
  OAI211_X1 U21683 ( .C1(n18611), .C2(n18540), .A(n18534), .B(n18533), .ZN(
        P3_U2978) );
  AOI22_X1 U21684 ( .A1(n18615), .A2(n18535), .B1(n18613), .B2(n18561), .ZN(
        n18539) );
  AOI22_X1 U21685 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18537), .B1(
        n18617), .B2(n18536), .ZN(n18538) );
  OAI211_X1 U21686 ( .C1(n18621), .C2(n18540), .A(n18539), .B(n18538), .ZN(
        P3_U2979) );
  INV_X1 U21687 ( .A(n18541), .ZN(n18565) );
  AND2_X1 U21688 ( .A1(n18686), .A2(n18545), .ZN(n18560) );
  AOI22_X1 U21689 ( .A1(n18567), .A2(n18616), .B1(n18566), .B2(n18560), .ZN(
        n18547) );
  OAI221_X1 U21690 ( .B1(n18545), .B2(n18544), .C1(n18545), .C2(n18543), .A(
        n18542), .ZN(n18562) );
  AOI22_X1 U21691 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18562), .B1(
        n18572), .B2(n18561), .ZN(n18546) );
  OAI211_X1 U21692 ( .C1(n18575), .C2(n18565), .A(n18547), .B(n18546), .ZN(
        P3_U2980) );
  AOI22_X1 U21693 ( .A1(n18578), .A2(n18561), .B1(n18577), .B2(n18560), .ZN(
        n18549) );
  AOI22_X1 U21694 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18562), .B1(
        n18576), .B2(n18616), .ZN(n18548) );
  OAI211_X1 U21695 ( .C1(n18581), .C2(n18565), .A(n18549), .B(n18548), .ZN(
        P3_U2981) );
  AOI22_X1 U21696 ( .A1(n18583), .A2(n18560), .B1(n18582), .B2(n18561), .ZN(
        n18551) );
  AOI22_X1 U21697 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18562), .B1(
        n18584), .B2(n18616), .ZN(n18550) );
  OAI211_X1 U21698 ( .C1(n18587), .C2(n18565), .A(n18551), .B(n18550), .ZN(
        P3_U2982) );
  AOI22_X1 U21699 ( .A1(n18588), .A2(n18560), .B1(n18590), .B2(n18616), .ZN(
        n18553) );
  AOI22_X1 U21700 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18562), .B1(
        n18589), .B2(n18561), .ZN(n18552) );
  OAI211_X1 U21701 ( .C1(n18593), .C2(n18565), .A(n18553), .B(n18552), .ZN(
        P3_U2983) );
  AOI22_X1 U21702 ( .A1(n18596), .A2(n18561), .B1(n18594), .B2(n18560), .ZN(
        n18555) );
  AOI22_X1 U21703 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18562), .B1(
        n18595), .B2(n18616), .ZN(n18554) );
  OAI211_X1 U21704 ( .C1(n18599), .C2(n18565), .A(n18555), .B(n18554), .ZN(
        P3_U2984) );
  AOI22_X1 U21705 ( .A1(n18601), .A2(n18560), .B1(n18600), .B2(n18561), .ZN(
        n18557) );
  AOI22_X1 U21706 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18562), .B1(
        n18602), .B2(n18616), .ZN(n18556) );
  OAI211_X1 U21707 ( .C1(n18605), .C2(n18565), .A(n18557), .B(n18556), .ZN(
        P3_U2985) );
  AOI22_X1 U21708 ( .A1(n18608), .A2(n18616), .B1(n18606), .B2(n18560), .ZN(
        n18559) );
  AOI22_X1 U21709 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18562), .B1(
        n18607), .B2(n18561), .ZN(n18558) );
  OAI211_X1 U21710 ( .C1(n18611), .C2(n18565), .A(n18559), .B(n18558), .ZN(
        P3_U2986) );
  AOI22_X1 U21711 ( .A1(n18617), .A2(n18561), .B1(n18615), .B2(n18560), .ZN(
        n18564) );
  AOI22_X1 U21712 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18562), .B1(
        n18613), .B2(n18616), .ZN(n18563) );
  OAI211_X1 U21713 ( .C1(n18621), .C2(n18565), .A(n18564), .B(n18563), .ZN(
        P3_U2987) );
  AND2_X1 U21714 ( .A1(n18686), .A2(n18569), .ZN(n18614) );
  AOI22_X1 U21715 ( .A1(n18567), .A2(n18612), .B1(n18566), .B2(n18614), .ZN(
        n18574) );
  AOI22_X1 U21716 ( .A1(n18571), .A2(n18570), .B1(n18569), .B2(n18568), .ZN(
        n18618) );
  AOI22_X1 U21717 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18618), .B1(
        n18572), .B2(n18616), .ZN(n18573) );
  OAI211_X1 U21718 ( .C1(n18622), .C2(n18575), .A(n18574), .B(n18573), .ZN(
        P3_U2988) );
  AOI22_X1 U21719 ( .A1(n18577), .A2(n18614), .B1(n18576), .B2(n18612), .ZN(
        n18580) );
  AOI22_X1 U21720 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18618), .B1(
        n18578), .B2(n18616), .ZN(n18579) );
  OAI211_X1 U21721 ( .C1(n18622), .C2(n18581), .A(n18580), .B(n18579), .ZN(
        P3_U2989) );
  AOI22_X1 U21722 ( .A1(n18583), .A2(n18614), .B1(n18582), .B2(n18616), .ZN(
        n18586) );
  AOI22_X1 U21723 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18618), .B1(
        n18584), .B2(n18612), .ZN(n18585) );
  OAI211_X1 U21724 ( .C1(n18622), .C2(n18587), .A(n18586), .B(n18585), .ZN(
        P3_U2990) );
  AOI22_X1 U21725 ( .A1(n18589), .A2(n18616), .B1(n18588), .B2(n18614), .ZN(
        n18592) );
  AOI22_X1 U21726 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18618), .B1(
        n18590), .B2(n18612), .ZN(n18591) );
  OAI211_X1 U21727 ( .C1(n18622), .C2(n18593), .A(n18592), .B(n18591), .ZN(
        P3_U2991) );
  AOI22_X1 U21728 ( .A1(n18595), .A2(n18612), .B1(n18594), .B2(n18614), .ZN(
        n18598) );
  AOI22_X1 U21729 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18618), .B1(
        n18596), .B2(n18616), .ZN(n18597) );
  OAI211_X1 U21730 ( .C1(n18622), .C2(n18599), .A(n18598), .B(n18597), .ZN(
        P3_U2992) );
  AOI22_X1 U21731 ( .A1(n18601), .A2(n18614), .B1(n18600), .B2(n18616), .ZN(
        n18604) );
  AOI22_X1 U21732 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18618), .B1(
        n18602), .B2(n18612), .ZN(n18603) );
  OAI211_X1 U21733 ( .C1(n18622), .C2(n18605), .A(n18604), .B(n18603), .ZN(
        P3_U2993) );
  AOI22_X1 U21734 ( .A1(n18607), .A2(n18616), .B1(n18606), .B2(n18614), .ZN(
        n18610) );
  AOI22_X1 U21735 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18618), .B1(
        n18608), .B2(n18612), .ZN(n18609) );
  OAI211_X1 U21736 ( .C1(n18622), .C2(n18611), .A(n18610), .B(n18609), .ZN(
        P3_U2994) );
  AOI22_X1 U21737 ( .A1(n18615), .A2(n18614), .B1(n18613), .B2(n18612), .ZN(
        n18620) );
  AOI22_X1 U21738 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18618), .B1(
        n18617), .B2(n18616), .ZN(n18619) );
  OAI211_X1 U21739 ( .C1(n18622), .C2(n18621), .A(n18620), .B(n18619), .ZN(
        P3_U2995) );
  NAND2_X1 U21740 ( .A1(n18624), .A2(n18623), .ZN(n18625) );
  AOI22_X1 U21741 ( .A1(n18628), .A2(n18627), .B1(n18626), .B2(n18625), .ZN(
        n18629) );
  OAI221_X1 U21742 ( .B1(n18631), .B2(n18661), .C1(n18631), .C2(n18630), .A(
        n18629), .ZN(n18825) );
  AOI21_X1 U21743 ( .B1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n18664), .A(
        n18825), .ZN(n18674) );
  AOI221_X1 U21744 ( .B1(P3_MORE_REG_SCAN_IN), .B2(n18633), .C1(
        P3_FLUSH_REG_SCAN_IN), .C2(n18633), .A(n18632), .ZN(n18673) );
  NAND2_X1 U21745 ( .A1(n18635), .A2(n18634), .ZN(n18637) );
  AOI21_X1 U21746 ( .B1(n18636), .B2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(
        n18655), .ZN(n18660) );
  INV_X1 U21747 ( .A(n18660), .ZN(n18644) );
  AOI22_X1 U21748 ( .A1(n18803), .A2(n18637), .B1(n18806), .B2(n18644), .ZN(
        n18800) );
  AOI22_X1 U21749 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18655), .B1(
        n18637), .B2(n18813), .ZN(n18640) );
  INV_X1 U21750 ( .A(n18640), .ZN(n18808) );
  NOR3_X1 U21751 ( .A1(n18639), .A2(n18638), .A3(n18808), .ZN(n18641) );
  OAI22_X1 U21752 ( .A1(n18800), .A2(n18641), .B1(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n18640), .ZN(n18643) );
  INV_X1 U21753 ( .A(n18664), .ZN(n18650) );
  AOI21_X1 U21754 ( .B1(n18643), .B2(n18650), .A(n18642), .ZN(n18652) );
  OAI211_X1 U21755 ( .C1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n18644), .B(n18659), .ZN(
        n18649) );
  OAI21_X1 U21756 ( .B1(n18647), .B2(n18646), .A(n18645), .ZN(n18653) );
  NAND3_X1 U21757 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n18656), .A3(
        n18653), .ZN(n18648) );
  OAI211_X1 U21758 ( .C1(n18795), .C2(n18661), .A(n18649), .B(n18648), .ZN(
        n18797) );
  AOI22_X1 U21759 ( .A1(n18664), .A2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n18797), .B2(n18650), .ZN(n18666) );
  OR2_X1 U21760 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18666), .ZN(
        n18651) );
  AOI221_X1 U21761 ( .B1(n18652), .B2(n18651), .C1(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .C2(n18666), .A(
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18670) );
  AOI22_X1 U21762 ( .A1(n18659), .A2(n18655), .B1(n18654), .B2(n18653), .ZN(
        n18657) );
  NAND2_X1 U21763 ( .A1(n18799), .A2(n18656), .ZN(n18658) );
  NAND2_X1 U21764 ( .A1(n18657), .A2(n18658), .ZN(n18788) );
  NOR2_X1 U21765 ( .A1(n18664), .A2(n18788), .ZN(n18665) );
  INV_X1 U21766 ( .A(n18658), .ZN(n18662) );
  OAI22_X1 U21767 ( .A1(n18662), .A2(n18661), .B1(n18660), .B2(n18659), .ZN(
        n18785) );
  NAND2_X1 U21768 ( .A1(n18789), .A2(n18785), .ZN(n18663) );
  OAI22_X1 U21769 ( .A1(n18665), .A2(n18789), .B1(n18664), .B2(n18663), .ZN(
        n18669) );
  OAI21_X1 U21770 ( .B1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(n18666), .ZN(n18667) );
  AOI222_X1 U21771 ( .A1(n18670), .A2(n18669), .B1(n18670), .B2(n18668), .C1(
        n18669), .C2(n18667), .ZN(n18672) );
  NAND4_X1 U21772 ( .A1(n18674), .A2(n18673), .A3(n18672), .A4(n18671), .ZN(
        n18683) );
  AOI211_X1 U21773 ( .C1(n18677), .C2(n18676), .A(n18675), .B(n18683), .ZN(
        n18780) );
  AOI21_X1 U21774 ( .B1(n18829), .B2(n18678), .A(n18780), .ZN(n18687) );
  NAND2_X1 U21775 ( .A1(n18829), .A2(n18679), .ZN(n18691) );
  INV_X1 U21776 ( .A(n18691), .ZN(n18680) );
  AOI211_X1 U21777 ( .C1(n18807), .C2(n18837), .A(P3_STATE2_REG_0__SCAN_IN), 
        .B(n18680), .ZN(n18681) );
  AOI211_X1 U21778 ( .C1(n18827), .C2(n18683), .A(n18682), .B(n18681), .ZN(
        n18684) );
  OAI221_X1 U21779 ( .B1(n18779), .B2(n18687), .C1(n18779), .C2(n18685), .A(
        n18684), .ZN(P3_U2996) );
  NOR4_X1 U21780 ( .A1(n18779), .A2(n18792), .A3(n18835), .A4(
        P3_STATE2_REG_2__SCAN_IN), .ZN(n18694) );
  INV_X1 U21781 ( .A(n18694), .ZN(n18690) );
  NAND3_X1 U21782 ( .A1(n18688), .A2(n18687), .A3(n18686), .ZN(n18689) );
  NAND4_X1 U21783 ( .A1(n18692), .A2(n18691), .A3(n18690), .A4(n18689), .ZN(
        P3_U2997) );
  OAI21_X1 U21784 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(
        P3_STATEBS16_REG_SCAN_IN), .A(n18693), .ZN(n18695) );
  AOI21_X1 U21785 ( .B1(n18696), .B2(n18695), .A(n18694), .ZN(P3_U2998) );
  INV_X1 U21786 ( .A(n18778), .ZN(n18775) );
  AND2_X1 U21787 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18775), .ZN(
        P3_U2999) );
  AND2_X1 U21788 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18775), .ZN(
        P3_U3000) );
  AND2_X1 U21789 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18775), .ZN(
        P3_U3001) );
  AND2_X1 U21790 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18775), .ZN(
        P3_U3002) );
  AND2_X1 U21791 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18775), .ZN(
        P3_U3003) );
  AND2_X1 U21792 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18775), .ZN(
        P3_U3004) );
  AND2_X1 U21793 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18775), .ZN(
        P3_U3005) );
  AND2_X1 U21794 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18775), .ZN(
        P3_U3006) );
  AND2_X1 U21795 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18775), .ZN(
        P3_U3007) );
  AND2_X1 U21796 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18775), .ZN(
        P3_U3008) );
  AND2_X1 U21797 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18775), .ZN(
        P3_U3009) );
  AND2_X1 U21798 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18775), .ZN(
        P3_U3010) );
  AND2_X1 U21799 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18775), .ZN(
        P3_U3011) );
  AND2_X1 U21800 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18775), .ZN(
        P3_U3012) );
  AND2_X1 U21801 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18775), .ZN(
        P3_U3013) );
  AND2_X1 U21802 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18775), .ZN(
        P3_U3014) );
  AND2_X1 U21803 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18775), .ZN(
        P3_U3015) );
  AND2_X1 U21804 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18775), .ZN(
        P3_U3016) );
  AND2_X1 U21805 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18775), .ZN(
        P3_U3017) );
  AND2_X1 U21806 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18775), .ZN(
        P3_U3018) );
  AND2_X1 U21807 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18775), .ZN(
        P3_U3019) );
  AND2_X1 U21808 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18775), .ZN(
        P3_U3020) );
  AND2_X1 U21809 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18775), .ZN(P3_U3021) );
  AND2_X1 U21810 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18775), .ZN(P3_U3022) );
  INV_X1 U21811 ( .A(P3_DATAWIDTH_REG_7__SCAN_IN), .ZN(n20817) );
  NOR2_X1 U21812 ( .A1(n20817), .A2(n18778), .ZN(P3_U3023) );
  AND2_X1 U21813 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18775), .ZN(P3_U3024) );
  AND2_X1 U21814 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18775), .ZN(P3_U3025) );
  AND2_X1 U21815 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18775), .ZN(P3_U3026) );
  AND2_X1 U21816 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18775), .ZN(P3_U3027) );
  AND2_X1 U21817 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18775), .ZN(P3_U3028) );
  NAND2_X1 U21818 ( .A1(n18829), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18706) );
  INV_X1 U21819 ( .A(n18706), .ZN(n18704) );
  OAI21_X1 U21820 ( .B1(n18697), .B2(n20687), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18698) );
  AOI22_X1 U21821 ( .A1(n18704), .A2(n18712), .B1(n18842), .B2(n18698), .ZN(
        n18700) );
  NAND3_X1 U21822 ( .A1(NA), .A2(n18710), .A3(n18699), .ZN(n18705) );
  OAI211_X1 U21823 ( .C1(P3_STATE_REG_0__SCAN_IN), .C2(P3_STATE_REG_2__SCAN_IN), .A(n18700), .B(n18705), .ZN(P3_U3029) );
  AOI21_X1 U21824 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(HOLD), .A(
        P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18701) );
  AOI21_X1 U21825 ( .B1(HOLD), .B2(P3_STATE_REG_2__SCAN_IN), .A(n18701), .ZN(
        n18702) );
  AOI22_X1 U21826 ( .A1(n18829), .A2(P3_STATE_REG_1__SCAN_IN), .B1(
        P3_STATE_REG_0__SCAN_IN), .B2(n18702), .ZN(n18703) );
  NAND2_X1 U21827 ( .A1(n18703), .A2(n18832), .ZN(P3_U3030) );
  AOI21_X1 U21828 ( .B1(n18710), .B2(n18705), .A(n18704), .ZN(n18711) );
  NOR2_X1 U21829 ( .A1(n18712), .A2(n20687), .ZN(n18708) );
  OAI22_X1 U21830 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18706), .ZN(n18707) );
  OAI22_X1 U21831 ( .A1(n18708), .A2(n18707), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18709) );
  OAI22_X1 U21832 ( .A1(n18711), .A2(n18712), .B1(n18710), .B2(n18709), .ZN(
        P3_U3031) );
  INV_X1 U21833 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18714) );
  OAI222_X1 U21834 ( .A1(n18714), .A2(n18769), .B1(n18713), .B2(n20776), .C1(
        n18715), .C2(n18765), .ZN(P3_U3032) );
  OAI222_X1 U21835 ( .A1(n18765), .A2(n18717), .B1(n18716), .B2(n20776), .C1(
        n18715), .C2(n18769), .ZN(P3_U3033) );
  OAI222_X1 U21836 ( .A1(n18765), .A2(n18719), .B1(n18718), .B2(n20776), .C1(
        n18717), .C2(n18769), .ZN(P3_U3034) );
  OAI222_X1 U21837 ( .A1(n18765), .A2(n18722), .B1(n18720), .B2(n20776), .C1(
        n18719), .C2(n18769), .ZN(P3_U3035) );
  INV_X1 U21838 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n18723) );
  OAI222_X1 U21839 ( .A1(n18722), .A2(n18769), .B1(n18721), .B2(n20776), .C1(
        n18723), .C2(n18765), .ZN(P3_U3036) );
  OAI222_X1 U21840 ( .A1(n18765), .A2(n18725), .B1(n18724), .B2(n20776), .C1(
        n18723), .C2(n18769), .ZN(P3_U3037) );
  OAI222_X1 U21841 ( .A1(n18765), .A2(n18728), .B1(n18726), .B2(n20776), .C1(
        n18725), .C2(n18769), .ZN(P3_U3038) );
  OAI222_X1 U21842 ( .A1(n18728), .A2(n18769), .B1(n18727), .B2(n20776), .C1(
        n18729), .C2(n18765), .ZN(P3_U3039) );
  OAI222_X1 U21843 ( .A1(n18765), .A2(n18731), .B1(n18730), .B2(n20776), .C1(
        n18729), .C2(n18769), .ZN(P3_U3040) );
  OAI222_X1 U21844 ( .A1(n18765), .A2(n18733), .B1(n18732), .B2(n20776), .C1(
        n18731), .C2(n18769), .ZN(P3_U3041) );
  OAI222_X1 U21845 ( .A1(n18765), .A2(n20954), .B1(n18734), .B2(n20776), .C1(
        n18733), .C2(n18769), .ZN(P3_U3042) );
  INV_X1 U21846 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18736) );
  OAI222_X1 U21847 ( .A1(n18765), .A2(n18736), .B1(n18735), .B2(n20776), .C1(
        n20954), .C2(n18769), .ZN(P3_U3043) );
  OAI222_X1 U21848 ( .A1(n18765), .A2(n20774), .B1(n18737), .B2(n20776), .C1(
        n18736), .C2(n18769), .ZN(P3_U3044) );
  OAI222_X1 U21849 ( .A1(n20773), .A2(n18769), .B1(n18738), .B2(n20776), .C1(
        n18739), .C2(n18765), .ZN(P3_U3046) );
  INV_X1 U21850 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18742) );
  OAI222_X1 U21851 ( .A1(n18765), .A2(n18742), .B1(n18740), .B2(n20776), .C1(
        n18739), .C2(n18769), .ZN(P3_U3047) );
  OAI222_X1 U21852 ( .A1(n18742), .A2(n18769), .B1(n18741), .B2(n20776), .C1(
        n18743), .C2(n18765), .ZN(P3_U3048) );
  OAI222_X1 U21853 ( .A1(n18765), .A2(n18746), .B1(n18744), .B2(n20776), .C1(
        n18743), .C2(n18769), .ZN(P3_U3049) );
  OAI222_X1 U21854 ( .A1(n18746), .A2(n18769), .B1(n18745), .B2(n20776), .C1(
        n18747), .C2(n18765), .ZN(P3_U3050) );
  OAI222_X1 U21855 ( .A1(n18765), .A2(n18750), .B1(n18748), .B2(n20776), .C1(
        n18747), .C2(n18769), .ZN(P3_U3051) );
  OAI222_X1 U21856 ( .A1(n18750), .A2(n18769), .B1(n18749), .B2(n20776), .C1(
        n18751), .C2(n18765), .ZN(P3_U3052) );
  OAI222_X1 U21857 ( .A1(n18765), .A2(n18754), .B1(n18752), .B2(n20776), .C1(
        n18751), .C2(n18769), .ZN(P3_U3053) );
  OAI222_X1 U21858 ( .A1(n18754), .A2(n18769), .B1(n18753), .B2(n20776), .C1(
        n18755), .C2(n18765), .ZN(P3_U3054) );
  OAI222_X1 U21859 ( .A1(n18765), .A2(n18756), .B1(n20938), .B2(n20776), .C1(
        n18755), .C2(n18769), .ZN(P3_U3055) );
  OAI222_X1 U21860 ( .A1(n18765), .A2(n18758), .B1(n18757), .B2(n20776), .C1(
        n18756), .C2(n18769), .ZN(P3_U3056) );
  OAI222_X1 U21861 ( .A1(n18765), .A2(n18759), .B1(n20795), .B2(n20776), .C1(
        n18758), .C2(n18769), .ZN(P3_U3057) );
  OAI222_X1 U21862 ( .A1(n18765), .A2(n18762), .B1(n18760), .B2(n20776), .C1(
        n18759), .C2(n18769), .ZN(P3_U3058) );
  OAI222_X1 U21863 ( .A1(n18762), .A2(n18769), .B1(n18761), .B2(n20776), .C1(
        n18763), .C2(n18765), .ZN(P3_U3059) );
  OAI222_X1 U21864 ( .A1(n18765), .A2(n18768), .B1(n18764), .B2(n20776), .C1(
        n18763), .C2(n18769), .ZN(P3_U3060) );
  OAI222_X1 U21865 ( .A1(n18769), .A2(n18768), .B1(n18767), .B2(n20776), .C1(
        n18766), .C2(n18765), .ZN(P3_U3061) );
  OAI22_X1 U21866 ( .A1(n18842), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n20776), .ZN(n18770) );
  INV_X1 U21867 ( .A(n18770), .ZN(P3_U3274) );
  OAI22_X1 U21868 ( .A1(n18842), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n20776), .ZN(n18771) );
  INV_X1 U21869 ( .A(n18771), .ZN(P3_U3275) );
  OAI22_X1 U21870 ( .A1(n18842), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n20776), .ZN(n18772) );
  INV_X1 U21871 ( .A(n18772), .ZN(P3_U3276) );
  OAI22_X1 U21872 ( .A1(n18842), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n20776), .ZN(n18773) );
  INV_X1 U21873 ( .A(n18773), .ZN(P3_U3277) );
  INV_X1 U21874 ( .A(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18816) );
  INV_X1 U21875 ( .A(n18776), .ZN(n18774) );
  AOI21_X1 U21876 ( .B1(n18775), .B2(n18816), .A(n18774), .ZN(P3_U3280) );
  INV_X1 U21877 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18777) );
  OAI21_X1 U21878 ( .B1(n18778), .B2(n18777), .A(n18776), .ZN(P3_U3281) );
  NOR2_X1 U21879 ( .A1(n18780), .A2(n18779), .ZN(n18783) );
  OAI21_X1 U21880 ( .B1(n18783), .B2(n18782), .A(n18781), .ZN(P3_U3282) );
  INV_X1 U21881 ( .A(n18784), .ZN(n18787) );
  NOR2_X1 U21882 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18844), .ZN(
        n18786) );
  AOI22_X1 U21883 ( .A1(n18807), .A2(n18787), .B1(n18786), .B2(n18785), .ZN(
        n18791) );
  INV_X1 U21884 ( .A(n18844), .ZN(n18809) );
  AOI21_X1 U21885 ( .B1(n18809), .B2(n18788), .A(n18814), .ZN(n18790) );
  OAI22_X1 U21886 ( .A1(n18814), .A2(n18791), .B1(n18790), .B2(n18789), .ZN(
        P3_U3285) );
  NOR2_X1 U21887 ( .A1(n18792), .A2(n18810), .ZN(n18801) );
  OAI22_X1 U21888 ( .A1(n18794), .A2(n18793), .B1(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18802) );
  INV_X1 U21889 ( .A(n18802), .ZN(n18796) );
  AOI222_X1 U21890 ( .A1(n18797), .A2(n18809), .B1(n18801), .B2(n18796), .C1(
        n18807), .C2(n18795), .ZN(n18798) );
  INV_X1 U21891 ( .A(n18814), .ZN(n18811) );
  AOI22_X1 U21892 ( .A1(n18814), .A2(n18799), .B1(n18798), .B2(n18811), .ZN(
        P3_U3288) );
  INV_X1 U21893 ( .A(n18800), .ZN(n18804) );
  AOI222_X1 U21894 ( .A1(n18804), .A2(n18809), .B1(n18807), .B2(n18803), .C1(
        n18802), .C2(n18801), .ZN(n18805) );
  AOI22_X1 U21895 ( .A1(n18814), .A2(n18806), .B1(n18805), .B2(n18811), .ZN(
        P3_U3289) );
  AOI222_X1 U21896 ( .A1(n18810), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18809), 
        .B2(n18808), .C1(n18813), .C2(n18807), .ZN(n18812) );
  AOI22_X1 U21897 ( .A1(n18814), .A2(n18813), .B1(n18812), .B2(n18811), .ZN(
        P3_U3290) );
  NOR3_X1 U21898 ( .A1(n18816), .A2(P3_REIP_REG_0__SCAN_IN), .A3(
        P3_REIP_REG_1__SCAN_IN), .ZN(n18815) );
  AOI221_X1 U21899 ( .B1(n18817), .B2(n18816), .C1(P3_REIP_REG_1__SCAN_IN), 
        .C2(P3_REIP_REG_0__SCAN_IN), .A(n18815), .ZN(n18819) );
  INV_X1 U21900 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18818) );
  INV_X1 U21901 ( .A(n18822), .ZN(n18820) );
  AOI22_X1 U21902 ( .A1(n18822), .A2(n18819), .B1(n18818), .B2(n18820), .ZN(
        P3_U3292) );
  NOR2_X1 U21903 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .ZN(n18821) );
  INV_X1 U21904 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20902) );
  AOI22_X1 U21905 ( .A1(n18822), .A2(n18821), .B1(n20902), .B2(n18820), .ZN(
        P3_U3293) );
  INV_X1 U21906 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18823) );
  AOI22_X1 U21907 ( .A1(n20776), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18823), 
        .B2(n18842), .ZN(P3_U3294) );
  MUX2_X1 U21908 ( .A(P3_MORE_REG_SCAN_IN), .B(n18825), .S(n18824), .Z(
        P3_U3295) );
  OAI22_X1 U21909 ( .A1(n18829), .A2(n18828), .B1(n18827), .B2(n18826), .ZN(
        n18830) );
  NOR2_X1 U21910 ( .A1(n18831), .A2(n18830), .ZN(n18841) );
  AOI21_X1 U21911 ( .B1(n18834), .B2(n18833), .A(n18832), .ZN(n18836) );
  OAI211_X1 U21912 ( .C1(n18845), .C2(n18836), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18835), .ZN(n18838) );
  AOI21_X1 U21913 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18838), .A(n18837), 
        .ZN(n18840) );
  NAND2_X1 U21914 ( .A1(n18841), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18839) );
  OAI21_X1 U21915 ( .B1(n18841), .B2(n18840), .A(n18839), .ZN(P3_U3296) );
  OAI22_X1 U21916 ( .A1(n18842), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n20776), .ZN(n18843) );
  INV_X1 U21917 ( .A(n18843), .ZN(P3_U3297) );
  OAI21_X1 U21918 ( .B1(n18844), .B2(P3_STATE2_REG_2__SCAN_IN), .A(n18846), 
        .ZN(n18849) );
  OAI22_X1 U21919 ( .A1(n18849), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18846), 
        .B2(n18845), .ZN(n18847) );
  INV_X1 U21920 ( .A(n18847), .ZN(P3_U3298) );
  OAI21_X1 U21921 ( .B1(n18849), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n18848), 
        .ZN(n18850) );
  INV_X1 U21922 ( .A(n18850), .ZN(P3_U3299) );
  NAND2_X1 U21923 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19776), .ZN(n19768) );
  NAND2_X1 U21924 ( .A1(n19764), .A2(n19759), .ZN(n19765) );
  OAI21_X1 U21925 ( .B1(n19764), .B2(n19768), .A(n19765), .ZN(n19843) );
  AOI21_X1 U21926 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19843), .ZN(n18851) );
  INV_X1 U21927 ( .A(n18851), .ZN(P2_U2815) );
  INV_X1 U21928 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18854) );
  OAI22_X1 U21929 ( .A1(n19892), .A2(n18854), .B1(n18853), .B2(n18852), .ZN(
        P2_U2816) );
  INV_X1 U21930 ( .A(n19770), .ZN(n18856) );
  AOI22_X1 U21931 ( .A1(P2_D_C_N_REG_SCAN_IN), .A2(n19906), .B1(n18856), .B2(
        n19764), .ZN(n18855) );
  OAI21_X1 U21932 ( .B1(P2_CODEFETCH_REG_SCAN_IN), .B2(n19906), .A(n18855), 
        .ZN(P2_U2817) );
  OAI21_X1 U21933 ( .B1(n18856), .B2(BS16), .A(n19843), .ZN(n19841) );
  OAI21_X1 U21934 ( .B1(n19843), .B2(n19896), .A(n19841), .ZN(P2_U2818) );
  NOR2_X1 U21935 ( .A1(n18858), .A2(n18857), .ZN(n19890) );
  OAI21_X1 U21936 ( .B1(n19890), .B2(n18860), .A(n18859), .ZN(P2_U2819) );
  NOR4_X1 U21937 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(P2_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_23__SCAN_IN), .ZN(n18864) );
  NOR4_X1 U21938 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_17__SCAN_IN), .A3(P2_DATAWIDTH_REG_18__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_19__SCAN_IN), .ZN(n18863) );
  NOR4_X1 U21939 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18862) );
  NOR4_X1 U21940 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18861) );
  NAND4_X1 U21941 ( .A1(n18864), .A2(n18863), .A3(n18862), .A4(n18861), .ZN(
        n18870) );
  NOR4_X1 U21942 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n18868) );
  AOI211_X1 U21943 ( .C1(P2_DATAWIDTH_REG_0__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_1__SCAN_IN), .A(P2_DATAWIDTH_REG_2__SCAN_IN), .B(
        P2_DATAWIDTH_REG_3__SCAN_IN), .ZN(n18867) );
  NOR4_X1 U21944 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_14__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_15__SCAN_IN), .ZN(n18866) );
  NOR4_X1 U21945 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n18865) );
  NAND4_X1 U21946 ( .A1(n18868), .A2(n18867), .A3(n18866), .A4(n18865), .ZN(
        n18869) );
  NOR2_X1 U21947 ( .A1(n18870), .A2(n18869), .ZN(n18879) );
  INV_X1 U21948 ( .A(n18879), .ZN(n18877) );
  NOR2_X1 U21949 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18877), .ZN(n18872) );
  INV_X1 U21950 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20923) );
  AOI22_X1 U21951 ( .A1(n18872), .A2(n14759), .B1(n20923), .B2(n18877), .ZN(
        P2_U2820) );
  OR3_X1 U21952 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18876) );
  INV_X1 U21953 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18871) );
  AOI22_X1 U21954 ( .A1(n18872), .A2(n18876), .B1(n18877), .B2(n18871), .ZN(
        P2_U2821) );
  INV_X1 U21955 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19842) );
  NAND2_X1 U21956 ( .A1(n18872), .A2(n19842), .ZN(n18875) );
  INV_X1 U21957 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n19777) );
  OAI21_X1 U21958 ( .B1(n19777), .B2(n14759), .A(n18879), .ZN(n18873) );
  OAI21_X1 U21959 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18879), .A(n18873), 
        .ZN(n18874) );
  OAI221_X1 U21960 ( .B1(n18875), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18875), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18874), .ZN(P2_U2822) );
  INV_X1 U21961 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18878) );
  OAI221_X1 U21962 ( .B1(n18879), .B2(n18878), .C1(n18877), .C2(n18876), .A(
        n18875), .ZN(P2_U2823) );
  INV_X1 U21963 ( .A(n18880), .ZN(n18884) );
  INV_X1 U21964 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19814) );
  OAI22_X1 U21965 ( .A1(n19104), .A2(n10613), .B1(n19814), .B2(n19110), .ZN(
        n18883) );
  OAI22_X1 U21966 ( .A1(n18881), .A2(n19086), .B1(n19101), .B2(n20917), .ZN(
        n18882) );
  AOI211_X1 U21967 ( .C1(n18884), .C2(n19112), .A(n18883), .B(n18882), .ZN(
        n18888) );
  OAI211_X1 U21968 ( .C1(n18886), .C2(n18890), .A(n19076), .B(n18885), .ZN(
        n18887) );
  OAI211_X1 U21969 ( .C1(n19085), .C2(n18889), .A(n18888), .B(n18887), .ZN(
        P2_U2834) );
  AOI211_X1 U21970 ( .C1(n18892), .C2(n18891), .A(n19116), .B(n18890), .ZN(
        n18895) );
  OAI22_X1 U21971 ( .A1(n19104), .A2(n18893), .B1(n9831), .B2(n19101), .ZN(
        n18894) );
  AOI211_X1 U21972 ( .C1(n19070), .C2(P2_REIP_REG_20__SCAN_IN), .A(n18895), 
        .B(n18894), .ZN(n18902) );
  INV_X1 U21973 ( .A(n18896), .ZN(n19120) );
  OAI22_X1 U21974 ( .A1(n18898), .A2(n19086), .B1(n18897), .B2(n19120), .ZN(
        n18899) );
  AOI21_X1 U21975 ( .B1(n18900), .B2(n19099), .A(n18899), .ZN(n18901) );
  OAI211_X1 U21976 ( .C1(n18903), .C2(n19091), .A(n18902), .B(n18901), .ZN(
        P2_U2835) );
  INV_X1 U21977 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19810) );
  OAI21_X1 U21978 ( .B1(n19810), .B2(n19110), .A(n19089), .ZN(n18907) );
  OAI22_X1 U21979 ( .A1(n18905), .A2(n19086), .B1(n19101), .B2(n18904), .ZN(
        n18906) );
  AOI211_X1 U21980 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n19064), .A(n18907), .B(
        n18906), .ZN(n18914) );
  NOR2_X1 U21981 ( .A1(n13666), .A2(n18908), .ZN(n18910) );
  XOR2_X1 U21982 ( .A(n18910), .B(n18909), .Z(n18911) );
  AOI22_X1 U21983 ( .A1(n18912), .A2(n19112), .B1(n19076), .B2(n18911), .ZN(
        n18913) );
  OAI211_X1 U21984 ( .C1(n18915), .C2(n19085), .A(n18914), .B(n18913), .ZN(
        P2_U2836) );
  NAND2_X1 U21985 ( .A1(n19080), .A2(n18928), .ZN(n18916) );
  XOR2_X1 U21986 ( .A(n18917), .B(n18916), .Z(n18926) );
  INV_X1 U21987 ( .A(n18918), .ZN(n18920) );
  AOI22_X1 U21988 ( .A1(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(n19065), .B1(
        P2_EBX_REG_18__SCAN_IN), .B2(n19064), .ZN(n18919) );
  OAI21_X1 U21989 ( .B1(n18920), .B2(n19086), .A(n18919), .ZN(n18921) );
  AOI211_X1 U21990 ( .C1(P2_REIP_REG_18__SCAN_IN), .C2(n19070), .A(n19069), 
        .B(n18921), .ZN(n18925) );
  AOI22_X1 U21991 ( .A1(n18923), .A2(n19112), .B1(n18922), .B2(n19099), .ZN(
        n18924) );
  OAI211_X1 U21992 ( .C1(n19116), .C2(n18926), .A(n18925), .B(n18924), .ZN(
        P2_U2837) );
  INV_X1 U21993 ( .A(n18927), .ZN(n18933) );
  OAI211_X1 U21994 ( .C1(n18930), .C2(n18940), .A(n18929), .B(n18928), .ZN(
        n18932) );
  AOI22_X1 U21995 ( .A1(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .A2(n19065), .B1(
        P2_EBX_REG_17__SCAN_IN), .B2(n19064), .ZN(n18931) );
  OAI211_X1 U21996 ( .C1(n18933), .C2(n19086), .A(n18932), .B(n18931), .ZN(
        n18934) );
  AOI211_X1 U21997 ( .C1(P2_REIP_REG_17__SCAN_IN), .C2(n19070), .A(n19069), 
        .B(n18934), .ZN(n18939) );
  INV_X1 U21998 ( .A(n18935), .ZN(n18936) );
  AOI22_X1 U21999 ( .A1(n18937), .A2(n19112), .B1(n18936), .B2(n19099), .ZN(
        n18938) );
  OAI211_X1 U22000 ( .C1(n18940), .C2(n19120), .A(n18939), .B(n18938), .ZN(
        P2_U2838) );
  OAI22_X1 U22001 ( .A1(n18942), .A2(n19086), .B1(n19101), .B2(n18941), .ZN(
        n18943) );
  INV_X1 U22002 ( .A(n18943), .ZN(n18944) );
  OAI21_X1 U22003 ( .B1(n19104), .B2(n10610), .A(n18944), .ZN(n18945) );
  AOI211_X1 U22004 ( .C1(P2_REIP_REG_16__SCAN_IN), .C2(n19070), .A(n19069), 
        .B(n18945), .ZN(n18952) );
  NAND2_X1 U22005 ( .A1(n19080), .A2(n18946), .ZN(n18947) );
  XOR2_X1 U22006 ( .A(n18948), .B(n18947), .Z(n18949) );
  AOI22_X1 U22007 ( .A1(n18950), .A2(n19099), .B1(n19076), .B2(n18949), .ZN(
        n18951) );
  OAI211_X1 U22008 ( .C1(n18953), .C2(n19091), .A(n18952), .B(n18951), .ZN(
        P2_U2839) );
  AOI22_X1 U22009 ( .A1(n18954), .A2(n19107), .B1(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n19065), .ZN(n18955) );
  OAI211_X1 U22010 ( .C1(n19803), .C2(n19110), .A(n18955), .B(n19089), .ZN(
        n18956) );
  AOI21_X1 U22011 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(n19064), .A(n18956), .ZN(
        n18964) );
  INV_X1 U22012 ( .A(n18957), .ZN(n18962) );
  NOR2_X1 U22013 ( .A1(n13666), .A2(n18958), .ZN(n18960) );
  XOR2_X1 U22014 ( .A(n18960), .B(n18959), .Z(n18961) );
  AOI22_X1 U22015 ( .A1(n18962), .A2(n19112), .B1(n19076), .B2(n18961), .ZN(
        n18963) );
  OAI211_X1 U22016 ( .C1(n18965), .C2(n19085), .A(n18964), .B(n18963), .ZN(
        P2_U2840) );
  NAND2_X1 U22017 ( .A1(n19080), .A2(n18966), .ZN(n18980) );
  XOR2_X1 U22018 ( .A(n18967), .B(n18980), .Z(n18974) );
  AOI22_X1 U22019 ( .A1(n18968), .A2(n19107), .B1(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n19065), .ZN(n18969) );
  OAI211_X1 U22020 ( .C1(n19801), .C2(n19110), .A(n18969), .B(n19089), .ZN(
        n18970) );
  AOI21_X1 U22021 ( .B1(P2_EBX_REG_14__SCAN_IN), .B2(n19064), .A(n18970), .ZN(
        n18973) );
  AOI22_X1 U22022 ( .A1(n18971), .A2(n19112), .B1(n19126), .B2(n19099), .ZN(
        n18972) );
  OAI211_X1 U22023 ( .C1(n19116), .C2(n18974), .A(n18973), .B(n18972), .ZN(
        P2_U2841) );
  INV_X1 U22024 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n19799) );
  AOI22_X1 U22025 ( .A1(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n19065), .B1(
        P2_EBX_REG_13__SCAN_IN), .B2(n19064), .ZN(n18975) );
  OAI211_X1 U22026 ( .C1(n19799), .C2(n19110), .A(n18975), .B(n19089), .ZN(
        n18978) );
  OAI22_X1 U22027 ( .A1(n18976), .A2(n19086), .B1(n19120), .B2(n18982), .ZN(
        n18977) );
  AOI211_X1 U22028 ( .C1(n18979), .C2(n19112), .A(n18978), .B(n18977), .ZN(
        n18985) );
  INV_X1 U22029 ( .A(n18980), .ZN(n18981) );
  OAI211_X1 U22030 ( .C1(n18983), .C2(n18982), .A(n19076), .B(n18981), .ZN(
        n18984) );
  OAI211_X1 U22031 ( .C1(n19085), .C2(n18986), .A(n18985), .B(n18984), .ZN(
        P2_U2842) );
  NAND2_X1 U22032 ( .A1(n19080), .A2(n18987), .ZN(n19003) );
  XOR2_X1 U22033 ( .A(n18988), .B(n19003), .Z(n18996) );
  AOI22_X1 U22034 ( .A1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(n19065), .B1(
        P2_EBX_REG_12__SCAN_IN), .B2(n19064), .ZN(n18989) );
  OAI21_X1 U22035 ( .B1(n18990), .B2(n19086), .A(n18989), .ZN(n18991) );
  AOI211_X1 U22036 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n19070), .A(n19069), 
        .B(n18991), .ZN(n18995) );
  AOI22_X1 U22037 ( .A1(n18993), .A2(n19112), .B1(n18992), .B2(n19099), .ZN(
        n18994) );
  OAI211_X1 U22038 ( .C1(n19116), .C2(n18996), .A(n18995), .B(n18994), .ZN(
        P2_U2843) );
  AOI22_X1 U22039 ( .A1(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .A2(n19065), .B1(
        P2_EBX_REG_11__SCAN_IN), .B2(n19064), .ZN(n18997) );
  OAI211_X1 U22040 ( .C1(n19795), .C2(n19110), .A(n18997), .B(n19089), .ZN(
        n19001) );
  OAI22_X1 U22041 ( .A1(n18999), .A2(n19085), .B1(n18998), .B2(n19086), .ZN(
        n19000) );
  AOI211_X1 U22042 ( .C1(n19002), .C2(n19112), .A(n19001), .B(n19000), .ZN(
        n19007) );
  INV_X1 U22043 ( .A(n19003), .ZN(n19004) );
  OAI211_X1 U22044 ( .C1(n19005), .C2(n19008), .A(n19076), .B(n19004), .ZN(
        n19006) );
  OAI211_X1 U22045 ( .C1(n19120), .C2(n19008), .A(n19007), .B(n19006), .ZN(
        P2_U2844) );
  OAI21_X1 U22046 ( .B1(n19793), .B2(n19110), .A(n19089), .ZN(n19011) );
  OAI22_X1 U22047 ( .A1(n19009), .A2(n19086), .B1(n19104), .B2(n10598), .ZN(
        n19010) );
  AOI211_X1 U22048 ( .C1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .C2(n19065), .A(
        n19011), .B(n19010), .ZN(n19018) );
  NAND2_X1 U22049 ( .A1(n19080), .A2(n19012), .ZN(n19013) );
  XOR2_X1 U22050 ( .A(n19014), .B(n19013), .Z(n19015) );
  AOI22_X1 U22051 ( .A1(n19016), .A2(n19112), .B1(n19076), .B2(n19015), .ZN(
        n19017) );
  OAI211_X1 U22052 ( .C1(n19019), .C2(n19085), .A(n19018), .B(n19017), .ZN(
        P2_U2845) );
  AOI22_X1 U22053 ( .A1(n19020), .A2(n19107), .B1(
        P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n19065), .ZN(n19021) );
  OAI211_X1 U22054 ( .C1(n19791), .C2(n19110), .A(n19021), .B(n19089), .ZN(
        n19022) );
  AOI21_X1 U22055 ( .B1(P2_EBX_REG_9__SCAN_IN), .B2(n19064), .A(n19022), .ZN(
        n19029) );
  NOR2_X1 U22056 ( .A1(n13666), .A2(n19023), .ZN(n19025) );
  XOR2_X1 U22057 ( .A(n19025), .B(n19024), .Z(n19026) );
  AOI22_X1 U22058 ( .A1(n19027), .A2(n19112), .B1(n19076), .B2(n19026), .ZN(
        n19028) );
  OAI211_X1 U22059 ( .C1(n19030), .C2(n19085), .A(n19029), .B(n19028), .ZN(
        P2_U2846) );
  AOI22_X1 U22060 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n19065), .B1(
        P2_EBX_REG_8__SCAN_IN), .B2(n19064), .ZN(n19031) );
  OAI21_X1 U22061 ( .B1(n19032), .B2(n19086), .A(n19031), .ZN(n19033) );
  AOI211_X1 U22062 ( .C1(P2_REIP_REG_8__SCAN_IN), .C2(n19070), .A(n19069), .B(
        n19033), .ZN(n19039) );
  NAND2_X1 U22063 ( .A1(n19080), .A2(n19034), .ZN(n19035) );
  XNOR2_X1 U22064 ( .A(n19036), .B(n19035), .ZN(n19037) );
  AOI22_X1 U22065 ( .A1(n19076), .A2(n19037), .B1(n19099), .B2(n19129), .ZN(
        n19038) );
  OAI211_X1 U22066 ( .C1(n19091), .C2(n19040), .A(n19039), .B(n19038), .ZN(
        P2_U2847) );
  AOI22_X1 U22067 ( .A1(n19041), .A2(n19107), .B1(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n19065), .ZN(n19042) );
  OAI211_X1 U22068 ( .C1(n19787), .C2(n19110), .A(n19042), .B(n19089), .ZN(
        n19043) );
  AOI21_X1 U22069 ( .B1(P2_EBX_REG_7__SCAN_IN), .B2(n19064), .A(n19043), .ZN(
        n19050) );
  NOR2_X1 U22070 ( .A1(n13666), .A2(n19044), .ZN(n19046) );
  XNOR2_X1 U22071 ( .A(n19046), .B(n19045), .ZN(n19048) );
  AOI22_X1 U22072 ( .A1(n19076), .A2(n19048), .B1(n19112), .B2(n19047), .ZN(
        n19049) );
  OAI211_X1 U22073 ( .C1(n19085), .C2(n19051), .A(n19050), .B(n19049), .ZN(
        P2_U2848) );
  OAI21_X1 U22074 ( .B1(n19786), .B2(n19110), .A(n19089), .ZN(n19055) );
  OAI22_X1 U22075 ( .A1(n19053), .A2(n19086), .B1(n19101), .B2(n19052), .ZN(
        n19054) );
  AOI211_X1 U22076 ( .C1(P2_EBX_REG_6__SCAN_IN), .C2(n19064), .A(n19055), .B(
        n19054), .ZN(n19062) );
  NAND2_X1 U22077 ( .A1(n19080), .A2(n19056), .ZN(n19057) );
  XNOR2_X1 U22078 ( .A(n19058), .B(n19057), .ZN(n19060) );
  AOI22_X1 U22079 ( .A1(n19076), .A2(n19060), .B1(n19112), .B2(n19059), .ZN(
        n19061) );
  OAI211_X1 U22080 ( .C1(n19085), .C2(n19063), .A(n19062), .B(n19061), .ZN(
        P2_U2849) );
  AOI22_X1 U22081 ( .A1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .A2(n19065), .B1(
        P2_EBX_REG_5__SCAN_IN), .B2(n19064), .ZN(n19066) );
  OAI21_X1 U22082 ( .B1(n19067), .B2(n19086), .A(n19066), .ZN(n19068) );
  AOI211_X1 U22083 ( .C1(P2_REIP_REG_5__SCAN_IN), .C2(n19070), .A(n19069), .B(
        n19068), .ZN(n19078) );
  NOR2_X1 U22084 ( .A1(n13666), .A2(n19071), .ZN(n19073) );
  XNOR2_X1 U22085 ( .A(n19073), .B(n19072), .ZN(n19075) );
  AOI22_X1 U22086 ( .A1(n19076), .A2(n19075), .B1(n19112), .B2(n19074), .ZN(
        n19077) );
  OAI211_X1 U22087 ( .C1(n19085), .C2(n19142), .A(n19078), .B(n19077), .ZN(
        P2_U2850) );
  NAND2_X1 U22088 ( .A1(n19080), .A2(n19079), .ZN(n19082) );
  XOR2_X1 U22089 ( .A(n19082), .B(n19081), .Z(n19098) );
  OAI22_X1 U22090 ( .A1(n19104), .A2(n19084), .B1(n19083), .B2(n19101), .ZN(
        n19096) );
  OAI22_X1 U22091 ( .A1(n19087), .A2(n19086), .B1(n19085), .B2(n19144), .ZN(
        n19088) );
  INV_X1 U22092 ( .A(n19088), .ZN(n19090) );
  OAI211_X1 U22093 ( .C1(n19783), .C2(n19110), .A(n19090), .B(n19089), .ZN(
        n19095) );
  OAI22_X1 U22094 ( .A1(n19146), .A2(n19093), .B1(n19092), .B2(n19091), .ZN(
        n19094) );
  NOR3_X1 U22095 ( .A1(n19096), .A2(n19095), .A3(n19094), .ZN(n19097) );
  OAI21_X1 U22096 ( .B1(n19098), .B2(n19116), .A(n19097), .ZN(P2_U2851) );
  NAND2_X1 U22097 ( .A1(n19866), .A2(n19099), .ZN(n19109) );
  INV_X1 U22098 ( .A(n19100), .ZN(n19106) );
  OAI22_X1 U22099 ( .A1(n19104), .A2(n19103), .B1(n19102), .B2(n19101), .ZN(
        n19105) );
  AOI21_X1 U22100 ( .B1(n19107), .B2(n19106), .A(n19105), .ZN(n19108) );
  OAI211_X1 U22101 ( .C1(n19777), .C2(n19110), .A(n19109), .B(n19108), .ZN(
        n19111) );
  AOI21_X1 U22102 ( .B1(n11297), .B2(n19112), .A(n19111), .ZN(n19115) );
  NAND2_X1 U22103 ( .A1(n19870), .A2(n19113), .ZN(n19114) );
  OAI211_X1 U22104 ( .C1(n19117), .C2(n19116), .A(n19115), .B(n19114), .ZN(
        n19118) );
  INV_X1 U22105 ( .A(n19118), .ZN(n19119) );
  OAI21_X1 U22106 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n19120), .A(
        n19119), .ZN(P2_U2854) );
  AOI22_X1 U22107 ( .A1(n19122), .A2(n19163), .B1(n19121), .B2(
        BUF2_REG_31__SCAN_IN), .ZN(n19125) );
  AOI22_X1 U22108 ( .A1(n19123), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19162), .ZN(n19124) );
  NAND2_X1 U22109 ( .A1(n19125), .A2(n19124), .ZN(P2_U2888) );
  INV_X1 U22110 ( .A(n19126), .ZN(n19128) );
  AOI22_X1 U22111 ( .A1(n19134), .A2(n19203), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n19162), .ZN(n19127) );
  OAI21_X1 U22112 ( .B1(n19143), .B2(n19128), .A(n19127), .ZN(P2_U2905) );
  INV_X1 U22113 ( .A(n19129), .ZN(n19132) );
  AOI22_X1 U22114 ( .A1(n19134), .A2(n19130), .B1(P2_EAX_REG_8__SCAN_IN), .B2(
        n19162), .ZN(n19131) );
  OAI21_X1 U22115 ( .B1(n19143), .B2(n19132), .A(n19131), .ZN(P2_U2911) );
  AOI22_X1 U22116 ( .A1(n19134), .A2(n19133), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n19162), .ZN(n19141) );
  INV_X1 U22117 ( .A(n19484), .ZN(n19851) );
  XNOR2_X1 U22118 ( .A(n19484), .B(n19850), .ZN(n19158) );
  NAND2_X1 U22119 ( .A1(n19859), .A2(n19135), .ZN(n19137) );
  NAND2_X1 U22120 ( .A1(n19137), .A2(n19136), .ZN(n19157) );
  NAND2_X1 U22121 ( .A1(n19158), .A2(n19157), .ZN(n19156) );
  OAI21_X1 U22122 ( .B1(n19851), .B2(n19850), .A(n19156), .ZN(n19138) );
  NAND2_X1 U22123 ( .A1(n19138), .A2(n19144), .ZN(n19147) );
  INV_X1 U22124 ( .A(n19146), .ZN(n19139) );
  NAND3_X1 U22125 ( .A1(n19147), .A2(n19139), .A3(n19164), .ZN(n19140) );
  OAI211_X1 U22126 ( .C1(n19143), .C2(n19142), .A(n19141), .B(n19140), .ZN(
        P2_U2914) );
  INV_X1 U22127 ( .A(n19144), .ZN(n19145) );
  AOI22_X1 U22128 ( .A1(n19163), .A2(n19145), .B1(P2_EAX_REG_4__SCAN_IN), .B2(
        n19162), .ZN(n19150) );
  XNOR2_X1 U22129 ( .A(n19147), .B(n19146), .ZN(n19148) );
  NAND2_X1 U22130 ( .A1(n19148), .A2(n19164), .ZN(n19149) );
  OAI211_X1 U22131 ( .C1(n19234), .C2(n19169), .A(n19150), .B(n19149), .ZN(
        P2_U2915) );
  INV_X1 U22132 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19151) );
  OAI22_X1 U22133 ( .A1(n19154), .A2(n19153), .B1(n19152), .B2(n19151), .ZN(
        n19155) );
  INV_X1 U22134 ( .A(n19155), .ZN(n19161) );
  OAI21_X1 U22135 ( .B1(n19158), .B2(n19157), .A(n19156), .ZN(n19159) );
  NAND2_X1 U22136 ( .A1(n19159), .A2(n19164), .ZN(n19160) );
  OAI211_X1 U22137 ( .C1(n19231), .C2(n19169), .A(n19161), .B(n19160), .ZN(
        P2_U2916) );
  AOI22_X1 U22138 ( .A1(n19163), .A2(n19166), .B1(P2_EAX_REG_0__SCAN_IN), .B2(
        n19162), .ZN(n19168) );
  OAI211_X1 U22139 ( .C1(n19877), .C2(n19166), .A(n19165), .B(n19164), .ZN(
        n19167) );
  OAI211_X1 U22140 ( .C1(n19170), .C2(n19169), .A(n19168), .B(n19167), .ZN(
        P2_U2919) );
  NOR2_X1 U22141 ( .A1(n19176), .A2(n19171), .ZN(P2_U2920) );
  INV_X1 U22142 ( .A(n19172), .ZN(n19173) );
  AOI22_X1 U22143 ( .A1(n19173), .A2(P2_EAX_REG_30__SCAN_IN), .B1(
        P2_UWORD_REG_14__SCAN_IN), .B2(n19181), .ZN(n19174) );
  OAI21_X1 U22144 ( .B1(n19176), .B2(n19175), .A(n19174), .ZN(P2_U2921) );
  AOI22_X1 U22145 ( .A1(n19181), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19177) );
  OAI21_X1 U22146 ( .B1(n12787), .B2(n19201), .A(n19177), .ZN(P2_U2936) );
  INV_X1 U22147 ( .A(P2_EAX_REG_14__SCAN_IN), .ZN(n19179) );
  AOI22_X1 U22148 ( .A1(n19181), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_14__SCAN_IN), .ZN(n19178) );
  OAI21_X1 U22149 ( .B1(n19179), .B2(n19201), .A(n19178), .ZN(P2_U2937) );
  AOI22_X1 U22150 ( .A1(n19181), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19180) );
  OAI21_X1 U22151 ( .B1(n12908), .B2(n19201), .A(n19180), .ZN(P2_U2938) );
  AOI22_X1 U22152 ( .A1(n19181), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19182) );
  OAI21_X1 U22153 ( .B1(n12901), .B2(n19201), .A(n19182), .ZN(P2_U2939) );
  AOI22_X1 U22154 ( .A1(n19181), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19183) );
  OAI21_X1 U22155 ( .B1(n12759), .B2(n19201), .A(n19183), .ZN(P2_U2940) );
  AOI22_X1 U22156 ( .A1(n19181), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_10__SCAN_IN), .ZN(n19184) );
  OAI21_X1 U22157 ( .B1(n12755), .B2(n19201), .A(n19184), .ZN(P2_U2941) );
  AOI22_X1 U22158 ( .A1(n19181), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19185) );
  OAI21_X1 U22159 ( .B1(n12914), .B2(n19201), .A(n19185), .ZN(P2_U2942) );
  AOI22_X1 U22160 ( .A1(n19181), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19186) );
  OAI21_X1 U22161 ( .B1(n19187), .B2(n19201), .A(n19186), .ZN(P2_U2943) );
  AOI22_X1 U22162 ( .A1(n19181), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19188) );
  OAI21_X1 U22163 ( .B1(n19189), .B2(n19201), .A(n19188), .ZN(P2_U2944) );
  AOI22_X1 U22164 ( .A1(n19181), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19190) );
  OAI21_X1 U22165 ( .B1(n19191), .B2(n19201), .A(n19190), .ZN(P2_U2945) );
  INV_X1 U22166 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n19193) );
  AOI22_X1 U22167 ( .A1(n19181), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19192) );
  OAI21_X1 U22168 ( .B1(n19193), .B2(n19201), .A(n19192), .ZN(P2_U2946) );
  INV_X1 U22169 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19195) );
  AOI22_X1 U22170 ( .A1(n19181), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19194) );
  OAI21_X1 U22171 ( .B1(n19195), .B2(n19201), .A(n19194), .ZN(P2_U2947) );
  AOI22_X1 U22172 ( .A1(n19181), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19196) );
  OAI21_X1 U22173 ( .B1(n19151), .B2(n19201), .A(n19196), .ZN(P2_U2948) );
  AOI22_X1 U22174 ( .A1(n19181), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19197) );
  OAI21_X1 U22175 ( .B1(n12889), .B2(n19201), .A(n19197), .ZN(P2_U2949) );
  AOI22_X1 U22176 ( .A1(n19181), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19198) );
  OAI21_X1 U22177 ( .B1(n12761), .B2(n19201), .A(n19198), .ZN(P2_U2950) );
  AOI22_X1 U22178 ( .A1(n19181), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19199), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19200) );
  OAI21_X1 U22179 ( .B1(n12892), .B2(n19201), .A(n19200), .ZN(P2_U2951) );
  AOI22_X1 U22180 ( .A1(n19202), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_30__SCAN_IN), .B2(n19206), .ZN(n19205) );
  NAND2_X1 U22181 ( .A1(n19204), .A2(n19203), .ZN(n19207) );
  NAND2_X1 U22182 ( .A1(n19205), .A2(n19207), .ZN(P2_U2966) );
  AOI22_X1 U22183 ( .A1(n19202), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(
        P2_EAX_REG_14__SCAN_IN), .B2(n19206), .ZN(n19208) );
  NAND2_X1 U22184 ( .A1(n19208), .A2(n19207), .ZN(P2_U2981) );
  INV_X1 U22185 ( .A(n19703), .ZN(n19660) );
  NAND2_X1 U22186 ( .A1(n19856), .A2(n19863), .ZN(n19317) );
  NOR2_X1 U22187 ( .A1(n19454), .A2(n19317), .ZN(n19253) );
  AOI22_X1 U22188 ( .A1(n19647), .A2(n19746), .B1(n19694), .B2(n19253), .ZN(
        n19220) );
  NAND2_X1 U22189 ( .A1(n19211), .A2(n19267), .ZN(n19212) );
  AOI21_X1 U22190 ( .B1(n19212), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19650), 
        .ZN(n19216) );
  OAI21_X1 U22191 ( .B1(n19213), .B2(n19691), .A(n19697), .ZN(n19214) );
  AOI21_X1 U22192 ( .B1(n19216), .B2(n19687), .A(n19214), .ZN(n19215) );
  OAI21_X1 U22193 ( .B1(n19215), .B2(n19253), .A(n19695), .ZN(n19256) );
  INV_X1 U22194 ( .A(n19687), .ZN(n19742) );
  OAI21_X1 U22195 ( .B1(n19742), .B2(n19253), .A(n19216), .ZN(n19218) );
  OAI21_X1 U22196 ( .B1(n19213), .B2(n19253), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19217) );
  NAND2_X1 U22197 ( .A1(n19218), .A2(n19217), .ZN(n19255) );
  AOI22_X1 U22198 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n19256), .B1(
        n15506), .B2(n19255), .ZN(n19219) );
  OAI211_X1 U22199 ( .C1(n19660), .C2(n19267), .A(n19220), .B(n19219), .ZN(
        P2_U3048) );
  INV_X1 U22200 ( .A(n19708), .ZN(n19664) );
  AOI22_X1 U22201 ( .A1(BUF1_REG_25__SCAN_IN), .A2(n19250), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n19249), .ZN(n19711) );
  NOR2_X2 U22202 ( .A1(n11518), .A2(n19251), .ZN(n19707) );
  AOI22_X1 U22203 ( .A1(n19661), .A2(n19746), .B1(n19707), .B2(n19253), .ZN(
        n19226) );
  AOI22_X1 U22204 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n19256), .B1(
        n19224), .B2(n19255), .ZN(n19225) );
  OAI211_X1 U22205 ( .C1(n19664), .C2(n19267), .A(n19226), .B(n19225), .ZN(
        P2_U3049) );
  AOI22_X1 U22206 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19250), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19249), .ZN(n19626) );
  AOI22_X1 U22207 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19250), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19249), .ZN(n19716) );
  NOR2_X2 U22208 ( .A1(n10767), .A2(n19251), .ZN(n19712) );
  AOI22_X1 U22209 ( .A1(n19623), .A2(n19746), .B1(n19712), .B2(n19253), .ZN(
        n19230) );
  AOI22_X1 U22210 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n19256), .B1(
        n19228), .B2(n19255), .ZN(n19229) );
  OAI211_X1 U22211 ( .C1(n19626), .C2(n19267), .A(n19230), .B(n19229), .ZN(
        P2_U3050) );
  AOI22_X1 U22212 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19250), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19249), .ZN(n19630) );
  AOI22_X1 U22213 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n19249), .B1(
        BUF1_REG_27__SCAN_IN), .B2(n19250), .ZN(n19722) );
  INV_X1 U22214 ( .A(n19722), .ZN(n19627) );
  NOR2_X2 U22215 ( .A1(n10180), .A2(n19251), .ZN(n19717) );
  AOI22_X1 U22216 ( .A1(n19627), .A2(n19746), .B1(n19717), .B2(n19253), .ZN(
        n19233) );
  NOR2_X2 U22217 ( .A1(n19231), .A2(n19614), .ZN(n19718) );
  AOI22_X1 U22218 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n19256), .B1(
        n19718), .B2(n19255), .ZN(n19232) );
  OAI211_X1 U22219 ( .C1(n19630), .C2(n19267), .A(n19233), .B(n19232), .ZN(
        P2_U3051) );
  AOI22_X1 U22220 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19250), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19249), .ZN(n19634) );
  AOI22_X1 U22221 ( .A1(BUF2_REG_28__SCAN_IN), .A2(n19249), .B1(
        BUF1_REG_28__SCAN_IN), .B2(n19250), .ZN(n19728) );
  INV_X1 U22222 ( .A(n19728), .ZN(n19631) );
  NOR2_X2 U22223 ( .A1(n10200), .A2(n19251), .ZN(n19723) );
  AOI22_X1 U22224 ( .A1(n19631), .A2(n19746), .B1(n19723), .B2(n19253), .ZN(
        n19236) );
  NOR2_X2 U22225 ( .A1(n19234), .A2(n19614), .ZN(n19724) );
  AOI22_X1 U22226 ( .A1(P2_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n19256), .B1(
        n19724), .B2(n19255), .ZN(n19235) );
  OAI211_X1 U22227 ( .C1(n19634), .C2(n19267), .A(n19236), .B(n19235), .ZN(
        P2_U3052) );
  OAI22_X1 U22228 ( .A1(n19238), .A2(n19244), .B1(n19237), .B2(n19242), .ZN(
        n19731) );
  AOI22_X1 U22229 ( .A1(BUF2_REG_29__SCAN_IN), .A2(n19249), .B1(
        BUF1_REG_29__SCAN_IN), .B2(n19250), .ZN(n19734) );
  NOR2_X2 U22230 ( .A1(n11687), .A2(n19251), .ZN(n19729) );
  AOI22_X1 U22231 ( .A1(n19671), .A2(n19746), .B1(n19729), .B2(n19253), .ZN(
        n19241) );
  NOR2_X2 U22232 ( .A1(n19239), .A2(n19614), .ZN(n19730) );
  AOI22_X1 U22233 ( .A1(P2_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n19256), .B1(
        n19730), .B2(n19255), .ZN(n19240) );
  OAI211_X1 U22234 ( .C1(n19674), .C2(n19267), .A(n19241), .B(n19240), .ZN(
        P2_U3053) );
  INV_X1 U22235 ( .A(n19737), .ZN(n19679) );
  AOI22_X1 U22236 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19250), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19249), .ZN(n19740) );
  INV_X1 U22237 ( .A(n19740), .ZN(n19676) );
  NOR2_X2 U22238 ( .A1(n10107), .A2(n19251), .ZN(n19735) );
  AOI22_X1 U22239 ( .A1(n19676), .A2(n19746), .B1(n19735), .B2(n19253), .ZN(
        n19248) );
  NOR2_X2 U22240 ( .A1(n19246), .A2(n19614), .ZN(n19736) );
  AOI22_X1 U22241 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n19256), .B1(
        n19736), .B2(n19255), .ZN(n19247) );
  OAI211_X1 U22242 ( .C1(n19679), .C2(n19267), .A(n19248), .B(n19247), .ZN(
        P2_U3054) );
  AOI22_X1 U22243 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n19250), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n19249), .ZN(n19607) );
  INV_X1 U22244 ( .A(n19751), .ZN(n19602) );
  NOR2_X2 U22245 ( .A1(n19252), .A2(n19251), .ZN(n19741) );
  AOI22_X1 U22246 ( .A1(n19602), .A2(n19746), .B1(n19741), .B2(n19253), .ZN(
        n19258) );
  NOR2_X2 U22247 ( .A1(n19254), .A2(n19614), .ZN(n19743) );
  AOI22_X1 U22248 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n19256), .B1(
        n19743), .B2(n19255), .ZN(n19257) );
  OAI211_X1 U22249 ( .C1(n19607), .C2(n19267), .A(n19258), .B(n19257), .ZN(
        P2_U3055) );
  OR2_X1 U22250 ( .A1(n19317), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19262) );
  NOR3_X2 U22251 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19880), .A3(
        n19317), .ZN(n19282) );
  INV_X1 U22252 ( .A(n19282), .ZN(n19259) );
  NAND2_X1 U22253 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19259), .ZN(n19260) );
  OR2_X1 U22254 ( .A1(n10430), .A2(n19260), .ZN(n19264) );
  INV_X1 U22255 ( .A(n19264), .ZN(n19261) );
  AOI211_X2 U22256 ( .C1(n19262), .C2(n19691), .A(n19752), .B(n19261), .ZN(
        n19283) );
  AOI22_X1 U22257 ( .A1(n19283), .A2(n15506), .B1(n19694), .B2(n19282), .ZN(
        n19269) );
  NAND2_X1 U22258 ( .A1(n19484), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19429) );
  NOR3_X1 U22259 ( .A1(n19485), .A2(n19429), .A3(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n19266) );
  NOR3_X1 U22260 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19874), .A3(
        n19317), .ZN(n19265) );
  OAI211_X1 U22261 ( .C1(n19266), .C2(n19265), .A(n19695), .B(n19264), .ZN(
        n19285) );
  AOI22_X1 U22262 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19285), .B1(
        n19284), .B2(n19647), .ZN(n19268) );
  OAI211_X1 U22263 ( .C1(n19660), .C2(n19316), .A(n19269), .B(n19268), .ZN(
        P2_U3056) );
  AOI22_X1 U22264 ( .A1(n19283), .A2(n19224), .B1(n19707), .B2(n19282), .ZN(
        n19271) );
  AOI22_X1 U22265 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19285), .B1(
        n19284), .B2(n19661), .ZN(n19270) );
  OAI211_X1 U22266 ( .C1(n19664), .C2(n19316), .A(n19271), .B(n19270), .ZN(
        P2_U3057) );
  AOI22_X1 U22267 ( .A1(n19283), .A2(n19228), .B1(n19712), .B2(n19282), .ZN(
        n19273) );
  AOI22_X1 U22268 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19285), .B1(
        n19284), .B2(n19623), .ZN(n19272) );
  OAI211_X1 U22269 ( .C1(n19626), .C2(n19316), .A(n19273), .B(n19272), .ZN(
        P2_U3058) );
  AOI22_X1 U22270 ( .A1(n19283), .A2(n19718), .B1(n19717), .B2(n19282), .ZN(
        n19275) );
  AOI22_X1 U22271 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19285), .B1(
        n19284), .B2(n19627), .ZN(n19274) );
  OAI211_X1 U22272 ( .C1(n19630), .C2(n19316), .A(n19275), .B(n19274), .ZN(
        P2_U3059) );
  AOI22_X1 U22273 ( .A1(n19283), .A2(n19724), .B1(n19723), .B2(n19282), .ZN(
        n19277) );
  AOI22_X1 U22274 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19285), .B1(
        n19284), .B2(n19631), .ZN(n19276) );
  OAI211_X1 U22275 ( .C1(n19634), .C2(n19316), .A(n19277), .B(n19276), .ZN(
        P2_U3060) );
  AOI22_X1 U22276 ( .A1(n19283), .A2(n19730), .B1(n19729), .B2(n19282), .ZN(
        n19279) );
  AOI22_X1 U22277 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19285), .B1(
        n19284), .B2(n19671), .ZN(n19278) );
  OAI211_X1 U22278 ( .C1(n19674), .C2(n19316), .A(n19279), .B(n19278), .ZN(
        P2_U3061) );
  AOI22_X1 U22279 ( .A1(n19283), .A2(n19736), .B1(n19735), .B2(n19282), .ZN(
        n19281) );
  AOI22_X1 U22280 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19285), .B1(
        n19284), .B2(n19676), .ZN(n19280) );
  OAI211_X1 U22281 ( .C1(n19679), .C2(n19316), .A(n19281), .B(n19280), .ZN(
        P2_U3062) );
  AOI22_X1 U22282 ( .A1(n19283), .A2(n19743), .B1(n19741), .B2(n19282), .ZN(
        n19287) );
  AOI22_X1 U22283 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19285), .B1(
        n19284), .B2(n19602), .ZN(n19286) );
  OAI211_X1 U22284 ( .C1(n19607), .C2(n19316), .A(n19287), .B(n19286), .ZN(
        P2_U3063) );
  NOR3_X2 U22285 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19873), .A3(
        n19317), .ZN(n19311) );
  OAI21_X1 U22286 ( .B1(n19288), .B2(n19311), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19291) );
  INV_X1 U22287 ( .A(n19516), .ZN(n19290) );
  INV_X1 U22288 ( .A(n19317), .ZN(n19289) );
  NAND2_X1 U22289 ( .A1(n19290), .A2(n19289), .ZN(n19293) );
  NAND2_X1 U22290 ( .A1(n19291), .A2(n19293), .ZN(n19312) );
  AOI22_X1 U22291 ( .A1(n19312), .A2(n15506), .B1(n19694), .B2(n19311), .ZN(
        n19298) );
  AOI21_X1 U22292 ( .B1(n10435), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19296) );
  INV_X1 U22293 ( .A(n19316), .ZN(n19292) );
  NOR2_X1 U22294 ( .A1(n19337), .A2(n19292), .ZN(n19294) );
  OAI211_X1 U22295 ( .C1(n19294), .C2(n19896), .A(n19844), .B(n19293), .ZN(
        n19295) );
  OAI211_X1 U22296 ( .C1(n19311), .C2(n19296), .A(n19295), .B(n19695), .ZN(
        n19313) );
  AOI22_X1 U22297 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19313), .B1(
        n19337), .B2(n19703), .ZN(n19297) );
  OAI211_X1 U22298 ( .C1(n19706), .C2(n19316), .A(n19298), .B(n19297), .ZN(
        P2_U3064) );
  AOI22_X1 U22299 ( .A1(n19312), .A2(n19224), .B1(n19707), .B2(n19311), .ZN(
        n19300) );
  AOI22_X1 U22300 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19313), .B1(
        n19337), .B2(n19708), .ZN(n19299) );
  OAI211_X1 U22301 ( .C1(n19711), .C2(n19316), .A(n19300), .B(n19299), .ZN(
        P2_U3065) );
  AOI22_X1 U22302 ( .A1(n19312), .A2(n19228), .B1(n19712), .B2(n19311), .ZN(
        n19302) );
  INV_X1 U22303 ( .A(n19626), .ZN(n19713) );
  AOI22_X1 U22304 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19313), .B1(
        n19337), .B2(n19713), .ZN(n19301) );
  OAI211_X1 U22305 ( .C1(n19716), .C2(n19316), .A(n19302), .B(n19301), .ZN(
        P2_U3066) );
  AOI22_X1 U22306 ( .A1(n19312), .A2(n19718), .B1(n19717), .B2(n19311), .ZN(
        n19304) );
  INV_X1 U22307 ( .A(n19630), .ZN(n19719) );
  AOI22_X1 U22308 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19313), .B1(
        n19337), .B2(n19719), .ZN(n19303) );
  OAI211_X1 U22309 ( .C1(n19722), .C2(n19316), .A(n19304), .B(n19303), .ZN(
        P2_U3067) );
  AOI22_X1 U22310 ( .A1(n19312), .A2(n19724), .B1(n19723), .B2(n19311), .ZN(
        n19306) );
  AOI22_X1 U22311 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19313), .B1(
        n19337), .B2(n19725), .ZN(n19305) );
  OAI211_X1 U22312 ( .C1(n19728), .C2(n19316), .A(n19306), .B(n19305), .ZN(
        P2_U3068) );
  AOI22_X1 U22313 ( .A1(n19312), .A2(n19730), .B1(n19729), .B2(n19311), .ZN(
        n19308) );
  AOI22_X1 U22314 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19313), .B1(
        n19337), .B2(n19731), .ZN(n19307) );
  OAI211_X1 U22315 ( .C1(n19734), .C2(n19316), .A(n19308), .B(n19307), .ZN(
        P2_U3069) );
  AOI22_X1 U22316 ( .A1(n19312), .A2(n19736), .B1(n19735), .B2(n19311), .ZN(
        n19310) );
  AOI22_X1 U22317 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19313), .B1(
        n19337), .B2(n19737), .ZN(n19309) );
  OAI211_X1 U22318 ( .C1(n19740), .C2(n19316), .A(n19310), .B(n19309), .ZN(
        P2_U3070) );
  AOI22_X1 U22319 ( .A1(n19312), .A2(n19743), .B1(n19741), .B2(n19311), .ZN(
        n19315) );
  AOI22_X1 U22320 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19313), .B1(
        n19337), .B2(n19745), .ZN(n19314) );
  OAI211_X1 U22321 ( .C1(n19751), .C2(n19316), .A(n19315), .B(n19314), .ZN(
        P2_U3071) );
  INV_X1 U22322 ( .A(n19337), .ZN(n19346) );
  NOR2_X1 U22323 ( .A1(n19544), .A2(n19317), .ZN(n19341) );
  AOI22_X1 U22324 ( .A1(n19703), .A2(n19372), .B1(n19341), .B2(n19694), .ZN(
        n19326) );
  OAI21_X1 U22325 ( .B1(n19429), .B2(n19847), .A(n19844), .ZN(n19324) );
  NOR2_X1 U22326 ( .A1(n19873), .A2(n19317), .ZN(n19321) );
  OAI21_X1 U22327 ( .B1(n10529), .B2(n19691), .A(n19697), .ZN(n19319) );
  INV_X1 U22328 ( .A(n19341), .ZN(n19318) );
  AOI21_X1 U22329 ( .B1(n19319), .B2(n19318), .A(n19614), .ZN(n19320) );
  OAI21_X1 U22330 ( .B1(n19324), .B2(n19321), .A(n19320), .ZN(n19343) );
  INV_X1 U22331 ( .A(n19321), .ZN(n19323) );
  OAI21_X1 U22332 ( .B1(n10529), .B2(n19341), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19322) );
  OAI21_X1 U22333 ( .B1(n19324), .B2(n19323), .A(n19322), .ZN(n19342) );
  AOI22_X1 U22334 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19343), .B1(
        n15506), .B2(n19342), .ZN(n19325) );
  OAI211_X1 U22335 ( .C1(n19706), .C2(n19346), .A(n19326), .B(n19325), .ZN(
        P2_U3072) );
  INV_X1 U22336 ( .A(n19372), .ZN(n19340) );
  AOI22_X1 U22337 ( .A1(n19661), .A2(n19337), .B1(n19341), .B2(n19707), .ZN(
        n19328) );
  AOI22_X1 U22338 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19343), .B1(
        n19224), .B2(n19342), .ZN(n19327) );
  OAI211_X1 U22339 ( .C1(n19664), .C2(n19340), .A(n19328), .B(n19327), .ZN(
        P2_U3073) );
  AOI22_X1 U22340 ( .A1(n19623), .A2(n19337), .B1(n19341), .B2(n19712), .ZN(
        n19330) );
  AOI22_X1 U22341 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19343), .B1(
        n19228), .B2(n19342), .ZN(n19329) );
  OAI211_X1 U22342 ( .C1(n19626), .C2(n19340), .A(n19330), .B(n19329), .ZN(
        P2_U3074) );
  AOI22_X1 U22343 ( .A1(n19719), .A2(n19372), .B1(n19341), .B2(n19717), .ZN(
        n19332) );
  AOI22_X1 U22344 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19343), .B1(
        n19718), .B2(n19342), .ZN(n19331) );
  OAI211_X1 U22345 ( .C1(n19722), .C2(n19346), .A(n19332), .B(n19331), .ZN(
        P2_U3075) );
  AOI22_X1 U22346 ( .A1(n19725), .A2(n19372), .B1(n19341), .B2(n19723), .ZN(
        n19334) );
  AOI22_X1 U22347 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19343), .B1(
        n19724), .B2(n19342), .ZN(n19333) );
  OAI211_X1 U22348 ( .C1(n19728), .C2(n19346), .A(n19334), .B(n19333), .ZN(
        P2_U3076) );
  AOI22_X1 U22349 ( .A1(n19671), .A2(n19337), .B1(n19341), .B2(n19729), .ZN(
        n19336) );
  AOI22_X1 U22350 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19343), .B1(
        n19730), .B2(n19342), .ZN(n19335) );
  OAI211_X1 U22351 ( .C1(n19674), .C2(n19340), .A(n19336), .B(n19335), .ZN(
        P2_U3077) );
  AOI22_X1 U22352 ( .A1(n19676), .A2(n19337), .B1(n19341), .B2(n19735), .ZN(
        n19339) );
  AOI22_X1 U22353 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19343), .B1(
        n19736), .B2(n19342), .ZN(n19338) );
  OAI211_X1 U22354 ( .C1(n19679), .C2(n19340), .A(n19339), .B(n19338), .ZN(
        P2_U3078) );
  AOI22_X1 U22355 ( .A1(n19745), .A2(n19372), .B1(n19341), .B2(n19741), .ZN(
        n19345) );
  AOI22_X1 U22356 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19343), .B1(
        n19743), .B2(n19342), .ZN(n19344) );
  OAI211_X1 U22357 ( .C1(n19751), .C2(n19346), .A(n19345), .B(n19344), .ZN(
        P2_U3079) );
  NOR2_X1 U22358 ( .A1(n19349), .A2(n19348), .ZN(n19580) );
  NAND2_X1 U22359 ( .A1(n19580), .A2(n19856), .ZN(n19354) );
  NOR2_X1 U22360 ( .A1(n19454), .A2(n19426), .ZN(n19370) );
  OAI21_X1 U22361 ( .B1(n19351), .B2(n19370), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19350) );
  OAI21_X1 U22362 ( .B1(n19354), .B2(n19650), .A(n19350), .ZN(n19371) );
  AOI22_X1 U22363 ( .A1(n19371), .A2(n15506), .B1(n19694), .B2(n19370), .ZN(
        n19357) );
  OAI21_X1 U22364 ( .B1(n19372), .B2(n19389), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19353) );
  AOI211_X1 U22365 ( .C1(n19351), .C2(n19697), .A(n19370), .B(n19844), .ZN(
        n19352) );
  AOI211_X1 U22366 ( .C1(n19354), .C2(n19353), .A(n19614), .B(n19352), .ZN(
        n19355) );
  AOI22_X1 U22367 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19373), .B1(
        n19372), .B2(n19647), .ZN(n19356) );
  OAI211_X1 U22368 ( .C1(n19660), .C2(n19405), .A(n19357), .B(n19356), .ZN(
        P2_U3080) );
  AOI22_X1 U22369 ( .A1(n19371), .A2(n19224), .B1(n19707), .B2(n19370), .ZN(
        n19359) );
  AOI22_X1 U22370 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19373), .B1(
        n19372), .B2(n19661), .ZN(n19358) );
  OAI211_X1 U22371 ( .C1(n19664), .C2(n19405), .A(n19359), .B(n19358), .ZN(
        P2_U3081) );
  AOI22_X1 U22372 ( .A1(n19371), .A2(n19228), .B1(n19712), .B2(n19370), .ZN(
        n19361) );
  AOI22_X1 U22373 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19373), .B1(
        n19372), .B2(n19623), .ZN(n19360) );
  OAI211_X1 U22374 ( .C1(n19626), .C2(n19405), .A(n19361), .B(n19360), .ZN(
        P2_U3082) );
  AOI22_X1 U22375 ( .A1(n19371), .A2(n19718), .B1(n19717), .B2(n19370), .ZN(
        n19363) );
  AOI22_X1 U22376 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19373), .B1(
        n19372), .B2(n19627), .ZN(n19362) );
  OAI211_X1 U22377 ( .C1(n19630), .C2(n19405), .A(n19363), .B(n19362), .ZN(
        P2_U3083) );
  AOI22_X1 U22378 ( .A1(n19371), .A2(n19724), .B1(n19723), .B2(n19370), .ZN(
        n19365) );
  AOI22_X1 U22379 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19373), .B1(
        n19372), .B2(n19631), .ZN(n19364) );
  OAI211_X1 U22380 ( .C1(n19634), .C2(n19405), .A(n19365), .B(n19364), .ZN(
        P2_U3084) );
  AOI22_X1 U22381 ( .A1(n19371), .A2(n19730), .B1(n19729), .B2(n19370), .ZN(
        n19367) );
  AOI22_X1 U22382 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19373), .B1(
        n19372), .B2(n19671), .ZN(n19366) );
  OAI211_X1 U22383 ( .C1(n19674), .C2(n19405), .A(n19367), .B(n19366), .ZN(
        P2_U3085) );
  AOI22_X1 U22384 ( .A1(n19371), .A2(n19736), .B1(n19735), .B2(n19370), .ZN(
        n19369) );
  AOI22_X1 U22385 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19373), .B1(
        n19372), .B2(n19676), .ZN(n19368) );
  OAI211_X1 U22386 ( .C1(n19679), .C2(n19405), .A(n19369), .B(n19368), .ZN(
        P2_U3086) );
  AOI22_X1 U22387 ( .A1(n19371), .A2(n19743), .B1(n19741), .B2(n19370), .ZN(
        n19375) );
  AOI22_X1 U22388 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19373), .B1(
        n19372), .B2(n19602), .ZN(n19374) );
  OAI211_X1 U22389 ( .C1(n19607), .C2(n19405), .A(n19375), .B(n19374), .ZN(
        P2_U3087) );
  NAND2_X1 U22390 ( .A1(n19376), .A2(n19873), .ZN(n19383) );
  NOR2_X1 U22391 ( .A1(n19880), .A2(n19383), .ZN(n19400) );
  AOI22_X1 U22392 ( .A1(n19703), .A2(n19414), .B1(n19400), .B2(n19694), .ZN(
        n19386) );
  OAI21_X1 U22393 ( .B1(n19429), .B2(n19608), .A(n19844), .ZN(n19384) );
  INV_X1 U22394 ( .A(n19383), .ZN(n19380) );
  INV_X1 U22395 ( .A(n19381), .ZN(n19378) );
  INV_X1 U22396 ( .A(n19400), .ZN(n19377) );
  OAI211_X1 U22397 ( .C1(n19378), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19377), 
        .B(n19650), .ZN(n19379) );
  OAI211_X1 U22398 ( .C1(n19384), .C2(n19380), .A(n19695), .B(n19379), .ZN(
        n19402) );
  OAI21_X1 U22399 ( .B1(n19381), .B2(n19400), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19382) );
  OAI21_X1 U22400 ( .B1(n19384), .B2(n19383), .A(n19382), .ZN(n19401) );
  AOI22_X1 U22401 ( .A1(P2_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n19402), .B1(
        n15506), .B2(n19401), .ZN(n19385) );
  OAI211_X1 U22402 ( .C1(n19706), .C2(n19405), .A(n19386), .B(n19385), .ZN(
        P2_U3088) );
  AOI22_X1 U22403 ( .A1(n19661), .A2(n19389), .B1(n19707), .B2(n19400), .ZN(
        n19388) );
  AOI22_X1 U22404 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19402), .B1(
        n19224), .B2(n19401), .ZN(n19387) );
  OAI211_X1 U22405 ( .C1(n19664), .C2(n19424), .A(n19388), .B(n19387), .ZN(
        P2_U3089) );
  AOI22_X1 U22406 ( .A1(n19623), .A2(n19389), .B1(n19400), .B2(n19712), .ZN(
        n19391) );
  AOI22_X1 U22407 ( .A1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n19402), .B1(
        n19228), .B2(n19401), .ZN(n19390) );
  OAI211_X1 U22408 ( .C1(n19626), .C2(n19424), .A(n19391), .B(n19390), .ZN(
        P2_U3090) );
  AOI22_X1 U22409 ( .A1(n19719), .A2(n19414), .B1(n19400), .B2(n19717), .ZN(
        n19393) );
  AOI22_X1 U22410 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n19402), .B1(
        n19718), .B2(n19401), .ZN(n19392) );
  OAI211_X1 U22411 ( .C1(n19722), .C2(n19405), .A(n19393), .B(n19392), .ZN(
        P2_U3091) );
  AOI22_X1 U22412 ( .A1(n19725), .A2(n19414), .B1(n19400), .B2(n19723), .ZN(
        n19395) );
  AOI22_X1 U22413 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n19402), .B1(
        n19724), .B2(n19401), .ZN(n19394) );
  OAI211_X1 U22414 ( .C1(n19728), .C2(n19405), .A(n19395), .B(n19394), .ZN(
        P2_U3092) );
  AOI22_X1 U22415 ( .A1(n19731), .A2(n19414), .B1(n19400), .B2(n19729), .ZN(
        n19397) );
  AOI22_X1 U22416 ( .A1(P2_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n19402), .B1(
        n19730), .B2(n19401), .ZN(n19396) );
  OAI211_X1 U22417 ( .C1(n19734), .C2(n19405), .A(n19397), .B(n19396), .ZN(
        P2_U3093) );
  AOI22_X1 U22418 ( .A1(n19737), .A2(n19414), .B1(n19400), .B2(n19735), .ZN(
        n19399) );
  AOI22_X1 U22419 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19402), .B1(
        n19736), .B2(n19401), .ZN(n19398) );
  OAI211_X1 U22420 ( .C1(n19740), .C2(n19405), .A(n19399), .B(n19398), .ZN(
        P2_U3094) );
  AOI22_X1 U22421 ( .A1(n19745), .A2(n19414), .B1(n19400), .B2(n19741), .ZN(
        n19404) );
  AOI22_X1 U22422 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19402), .B1(
        n19743), .B2(n19401), .ZN(n19403) );
  OAI211_X1 U22423 ( .C1(n19751), .C2(n19405), .A(n19404), .B(n19403), .ZN(
        P2_U3095) );
  AOI22_X1 U22424 ( .A1(n19420), .A2(n19224), .B1(n19707), .B2(n19419), .ZN(
        n19407) );
  AOI22_X1 U22425 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19421), .B1(
        n19414), .B2(n19661), .ZN(n19406) );
  OAI211_X1 U22426 ( .C1(n19664), .C2(n19453), .A(n19407), .B(n19406), .ZN(
        P2_U3097) );
  AOI22_X1 U22427 ( .A1(n19420), .A2(n19228), .B1(n19712), .B2(n19419), .ZN(
        n19409) );
  AOI22_X1 U22428 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19421), .B1(
        n19446), .B2(n19713), .ZN(n19408) );
  OAI211_X1 U22429 ( .C1(n19716), .C2(n19424), .A(n19409), .B(n19408), .ZN(
        P2_U3098) );
  AOI22_X1 U22430 ( .A1(n19420), .A2(n19718), .B1(n19717), .B2(n19419), .ZN(
        n19411) );
  AOI22_X1 U22431 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19421), .B1(
        n19446), .B2(n19719), .ZN(n19410) );
  OAI211_X1 U22432 ( .C1(n19722), .C2(n19424), .A(n19411), .B(n19410), .ZN(
        P2_U3099) );
  AOI22_X1 U22433 ( .A1(n19420), .A2(n19724), .B1(n19723), .B2(n19419), .ZN(
        n19413) );
  AOI22_X1 U22434 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19421), .B1(
        n19414), .B2(n19631), .ZN(n19412) );
  OAI211_X1 U22435 ( .C1(n19634), .C2(n19453), .A(n19413), .B(n19412), .ZN(
        P2_U3100) );
  AOI22_X1 U22436 ( .A1(n19420), .A2(n19730), .B1(n19729), .B2(n19419), .ZN(
        n19416) );
  AOI22_X1 U22437 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19421), .B1(
        n19414), .B2(n19671), .ZN(n19415) );
  OAI211_X1 U22438 ( .C1(n19674), .C2(n19453), .A(n19416), .B(n19415), .ZN(
        P2_U3101) );
  AOI22_X1 U22439 ( .A1(n19420), .A2(n19736), .B1(n19735), .B2(n19419), .ZN(
        n19418) );
  AOI22_X1 U22440 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19421), .B1(
        n19446), .B2(n19737), .ZN(n19417) );
  OAI211_X1 U22441 ( .C1(n19740), .C2(n19424), .A(n19418), .B(n19417), .ZN(
        P2_U3102) );
  AOI22_X1 U22442 ( .A1(n19420), .A2(n19743), .B1(n19741), .B2(n19419), .ZN(
        n19423) );
  AOI22_X1 U22443 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19421), .B1(
        n19446), .B2(n19745), .ZN(n19422) );
  OAI211_X1 U22444 ( .C1(n19751), .C2(n19424), .A(n19423), .B(n19422), .ZN(
        P2_U3103) );
  NOR2_X1 U22445 ( .A1(n19690), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19433) );
  INV_X1 U22446 ( .A(n19433), .ZN(n19428) );
  NOR2_X1 U22447 ( .A1(n19544), .A2(n19426), .ZN(n19460) );
  OR2_X1 U22448 ( .A1(n19460), .A2(n19691), .ZN(n19427) );
  NOR2_X1 U22449 ( .A1(n10429), .A2(n19427), .ZN(n19431) );
  AOI211_X2 U22450 ( .C1(n19428), .C2(n19691), .A(n19752), .B(n19431), .ZN(
        n19449) );
  AOI22_X1 U22451 ( .A1(n19449), .A2(n15506), .B1(n19694), .B2(n19460), .ZN(
        n19435) );
  NOR2_X1 U22452 ( .A1(n19429), .A2(n19645), .ZN(n19845) );
  OAI21_X1 U22453 ( .B1(n19460), .B2(n19697), .A(n19695), .ZN(n19430) );
  NOR2_X1 U22454 ( .A1(n19431), .A2(n19430), .ZN(n19432) );
  OAI21_X1 U22455 ( .B1(n19433), .B2(n19845), .A(n19432), .ZN(n19450) );
  AOI22_X1 U22456 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19450), .B1(
        n19446), .B2(n19647), .ZN(n19434) );
  OAI211_X1 U22457 ( .C1(n19660), .C2(n19483), .A(n19435), .B(n19434), .ZN(
        P2_U3104) );
  AOI22_X1 U22458 ( .A1(n19449), .A2(n19224), .B1(n19707), .B2(n19460), .ZN(
        n19437) );
  AOI22_X1 U22459 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19450), .B1(
        n19446), .B2(n19661), .ZN(n19436) );
  OAI211_X1 U22460 ( .C1(n19664), .C2(n19483), .A(n19437), .B(n19436), .ZN(
        P2_U3105) );
  AOI22_X1 U22461 ( .A1(n19449), .A2(n19228), .B1(n19712), .B2(n19460), .ZN(
        n19439) );
  AOI22_X1 U22462 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19450), .B1(
        n19446), .B2(n19623), .ZN(n19438) );
  OAI211_X1 U22463 ( .C1(n19626), .C2(n19483), .A(n19439), .B(n19438), .ZN(
        P2_U3106) );
  AOI22_X1 U22464 ( .A1(n19449), .A2(n19718), .B1(n19717), .B2(n19460), .ZN(
        n19441) );
  AOI22_X1 U22465 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19450), .B1(
        n19446), .B2(n19627), .ZN(n19440) );
  OAI211_X1 U22466 ( .C1(n19630), .C2(n19483), .A(n19441), .B(n19440), .ZN(
        P2_U3107) );
  AOI22_X1 U22467 ( .A1(n19449), .A2(n19724), .B1(n19723), .B2(n19460), .ZN(
        n19443) );
  AOI22_X1 U22468 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19450), .B1(
        n19455), .B2(n19725), .ZN(n19442) );
  OAI211_X1 U22469 ( .C1(n19728), .C2(n19453), .A(n19443), .B(n19442), .ZN(
        P2_U3108) );
  AOI22_X1 U22470 ( .A1(n19449), .A2(n19730), .B1(n19729), .B2(n19460), .ZN(
        n19445) );
  AOI22_X1 U22471 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19450), .B1(
        n19455), .B2(n19731), .ZN(n19444) );
  OAI211_X1 U22472 ( .C1(n19734), .C2(n19453), .A(n19445), .B(n19444), .ZN(
        P2_U3109) );
  AOI22_X1 U22473 ( .A1(n19449), .A2(n19736), .B1(n19735), .B2(n19460), .ZN(
        n19448) );
  AOI22_X1 U22474 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19450), .B1(
        n19446), .B2(n19676), .ZN(n19447) );
  OAI211_X1 U22475 ( .C1(n19679), .C2(n19483), .A(n19448), .B(n19447), .ZN(
        P2_U3110) );
  AOI22_X1 U22476 ( .A1(n19449), .A2(n19743), .B1(n19741), .B2(n19460), .ZN(
        n19452) );
  AOI22_X1 U22477 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19450), .B1(
        n19455), .B2(n19745), .ZN(n19451) );
  OAI211_X1 U22478 ( .C1(n19751), .C2(n19453), .A(n19452), .B(n19451), .ZN(
        P2_U3111) );
  NOR2_X1 U22479 ( .A1(n19856), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n19542) );
  INV_X1 U22480 ( .A(n19542), .ZN(n19545) );
  NOR2_X1 U22481 ( .A1(n19454), .A2(n19545), .ZN(n19478) );
  AOI22_X1 U22482 ( .A1(n19703), .A2(n19506), .B1(n19694), .B2(n19478), .ZN(
        n19465) );
  NOR3_X1 U22483 ( .A1(n19459), .A2(n19478), .A3(n19691), .ZN(n19458) );
  NOR2_X1 U22484 ( .A1(n19506), .A2(n19455), .ZN(n19456) );
  OAI21_X1 U22485 ( .B1(n19456), .B2(n19896), .A(n19844), .ZN(n19463) );
  AOI221_X1 U22486 ( .B1(n19697), .B2(n19463), .C1(n19697), .C2(n19460), .A(
        n19478), .ZN(n19457) );
  OAI21_X1 U22487 ( .B1(n19459), .B2(n19478), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19462) );
  NOR2_X1 U22488 ( .A1(n19478), .A2(n19460), .ZN(n19461) );
  AOI22_X1 U22489 ( .A1(n19463), .A2(n19462), .B1(n19461), .B2(n19691), .ZN(
        n19479) );
  AOI22_X1 U22490 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19480), .B1(
        n15506), .B2(n19479), .ZN(n19464) );
  OAI211_X1 U22491 ( .C1(n19706), .C2(n19483), .A(n19465), .B(n19464), .ZN(
        P2_U3112) );
  AOI22_X1 U22492 ( .A1(n19708), .A2(n19506), .B1(n19707), .B2(n19478), .ZN(
        n19467) );
  AOI22_X1 U22493 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19480), .B1(
        n19224), .B2(n19479), .ZN(n19466) );
  OAI211_X1 U22494 ( .C1(n19711), .C2(n19483), .A(n19467), .B(n19466), .ZN(
        P2_U3113) );
  AOI22_X1 U22495 ( .A1(n19713), .A2(n19506), .B1(n19712), .B2(n19478), .ZN(
        n19469) );
  AOI22_X1 U22496 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19480), .B1(
        n19228), .B2(n19479), .ZN(n19468) );
  OAI211_X1 U22497 ( .C1(n19716), .C2(n19483), .A(n19469), .B(n19468), .ZN(
        P2_U3114) );
  AOI22_X1 U22498 ( .A1(n19719), .A2(n19506), .B1(n19717), .B2(n19478), .ZN(
        n19471) );
  AOI22_X1 U22499 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19480), .B1(
        n19718), .B2(n19479), .ZN(n19470) );
  OAI211_X1 U22500 ( .C1(n19722), .C2(n19483), .A(n19471), .B(n19470), .ZN(
        P2_U3115) );
  AOI22_X1 U22501 ( .A1(n19725), .A2(n19506), .B1(n19723), .B2(n19478), .ZN(
        n19473) );
  AOI22_X1 U22502 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19480), .B1(
        n19724), .B2(n19479), .ZN(n19472) );
  OAI211_X1 U22503 ( .C1(n19728), .C2(n19483), .A(n19473), .B(n19472), .ZN(
        P2_U3116) );
  AOI22_X1 U22504 ( .A1(n19731), .A2(n19506), .B1(n19729), .B2(n19478), .ZN(
        n19475) );
  AOI22_X1 U22505 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19480), .B1(
        n19730), .B2(n19479), .ZN(n19474) );
  OAI211_X1 U22506 ( .C1(n19734), .C2(n19483), .A(n19475), .B(n19474), .ZN(
        P2_U3117) );
  AOI22_X1 U22507 ( .A1(n19737), .A2(n19506), .B1(n19735), .B2(n19478), .ZN(
        n19477) );
  AOI22_X1 U22508 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19480), .B1(
        n19736), .B2(n19479), .ZN(n19476) );
  OAI211_X1 U22509 ( .C1(n19740), .C2(n19483), .A(n19477), .B(n19476), .ZN(
        P2_U3118) );
  AOI22_X1 U22510 ( .A1(n19506), .A2(n19745), .B1(n19741), .B2(n19478), .ZN(
        n19482) );
  AOI22_X1 U22511 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19480), .B1(
        n19743), .B2(n19479), .ZN(n19481) );
  OAI211_X1 U22512 ( .C1(n19751), .C2(n19483), .A(n19482), .B(n19481), .ZN(
        P2_U3119) );
  NOR3_X2 U22513 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19880), .A3(
        n19545), .ZN(n19517) );
  AOI22_X1 U22514 ( .A1(n19703), .A2(n19518), .B1(n19694), .B2(n19517), .ZN(
        n19495) );
  NOR2_X1 U22515 ( .A1(n19484), .A2(n19896), .ZN(n19700) );
  INV_X1 U22516 ( .A(n19700), .ZN(n19486) );
  OAI21_X1 U22517 ( .B1(n19486), .B2(n19485), .A(n19844), .ZN(n19493) );
  NAND2_X1 U22518 ( .A1(n19873), .A2(n19542), .ZN(n19492) );
  INV_X1 U22519 ( .A(n19492), .ZN(n19489) );
  INV_X1 U22520 ( .A(n19517), .ZN(n19487) );
  OAI211_X1 U22521 ( .C1(n10425), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19487), 
        .B(n19650), .ZN(n19488) );
  OAI211_X1 U22522 ( .C1(n19493), .C2(n19489), .A(n19695), .B(n19488), .ZN(
        n19510) );
  OAI21_X1 U22523 ( .B1(n19490), .B2(n19517), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19491) );
  OAI21_X1 U22524 ( .B1(n19493), .B2(n19492), .A(n19491), .ZN(n19509) );
  AOI22_X1 U22525 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19510), .B1(
        n15506), .B2(n19509), .ZN(n19494) );
  OAI211_X1 U22526 ( .C1(n19706), .C2(n19513), .A(n19495), .B(n19494), .ZN(
        P2_U3120) );
  AOI22_X1 U22527 ( .A1(n19708), .A2(n19518), .B1(n19707), .B2(n19517), .ZN(
        n19497) );
  AOI22_X1 U22528 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19510), .B1(
        n19224), .B2(n19509), .ZN(n19496) );
  OAI211_X1 U22529 ( .C1(n19711), .C2(n19513), .A(n19497), .B(n19496), .ZN(
        P2_U3121) );
  AOI22_X1 U22530 ( .A1(n19623), .A2(n19506), .B1(n19712), .B2(n19517), .ZN(
        n19499) );
  AOI22_X1 U22531 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19510), .B1(
        n19228), .B2(n19509), .ZN(n19498) );
  OAI211_X1 U22532 ( .C1(n19626), .C2(n19541), .A(n19499), .B(n19498), .ZN(
        P2_U3122) );
  AOI22_X1 U22533 ( .A1(n19627), .A2(n19506), .B1(n19717), .B2(n19517), .ZN(
        n19501) );
  AOI22_X1 U22534 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19510), .B1(
        n19718), .B2(n19509), .ZN(n19500) );
  OAI211_X1 U22535 ( .C1(n19630), .C2(n19541), .A(n19501), .B(n19500), .ZN(
        P2_U3123) );
  AOI22_X1 U22536 ( .A1(n19725), .A2(n19518), .B1(n19723), .B2(n19517), .ZN(
        n19503) );
  AOI22_X1 U22537 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19510), .B1(
        n19724), .B2(n19509), .ZN(n19502) );
  OAI211_X1 U22538 ( .C1(n19728), .C2(n19513), .A(n19503), .B(n19502), .ZN(
        P2_U3124) );
  AOI22_X1 U22539 ( .A1(n19671), .A2(n19506), .B1(n19729), .B2(n19517), .ZN(
        n19505) );
  AOI22_X1 U22540 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19510), .B1(
        n19730), .B2(n19509), .ZN(n19504) );
  OAI211_X1 U22541 ( .C1(n19674), .C2(n19541), .A(n19505), .B(n19504), .ZN(
        P2_U3125) );
  AOI22_X1 U22542 ( .A1(n19676), .A2(n19506), .B1(n19735), .B2(n19517), .ZN(
        n19508) );
  AOI22_X1 U22543 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19510), .B1(
        n19736), .B2(n19509), .ZN(n19507) );
  OAI211_X1 U22544 ( .C1(n19679), .C2(n19541), .A(n19508), .B(n19507), .ZN(
        P2_U3126) );
  AOI22_X1 U22545 ( .A1(n19518), .A2(n19745), .B1(n19741), .B2(n19517), .ZN(
        n19512) );
  AOI22_X1 U22546 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19510), .B1(
        n19743), .B2(n19509), .ZN(n19511) );
  OAI211_X1 U22547 ( .C1(n19751), .C2(n19513), .A(n19512), .B(n19511), .ZN(
        P2_U3127) );
  INV_X1 U22548 ( .A(n10420), .ZN(n19514) );
  NOR3_X2 U22549 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19873), .A3(
        n19545), .ZN(n19536) );
  OAI21_X1 U22550 ( .B1(n19514), .B2(n19536), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19515) );
  OAI21_X1 U22551 ( .B1(n19545), .B2(n19516), .A(n19515), .ZN(n19537) );
  AOI22_X1 U22552 ( .A1(n19537), .A2(n15506), .B1(n19694), .B2(n19536), .ZN(
        n19523) );
  AOI221_X1 U22553 ( .B1(n19518), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19569), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19517), .ZN(n19519) );
  MUX2_X1 U22554 ( .A(n10420), .B(n19519), .S(n19691), .Z(n19520) );
  NOR2_X1 U22555 ( .A1(n19520), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19521) );
  AOI22_X1 U22556 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19538), .B1(
        n19569), .B2(n19703), .ZN(n19522) );
  OAI211_X1 U22557 ( .C1(n19706), .C2(n19541), .A(n19523), .B(n19522), .ZN(
        P2_U3128) );
  AOI22_X1 U22558 ( .A1(n19537), .A2(n19224), .B1(n19707), .B2(n19536), .ZN(
        n19525) );
  AOI22_X1 U22559 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19538), .B1(
        n19569), .B2(n19708), .ZN(n19524) );
  OAI211_X1 U22560 ( .C1(n19711), .C2(n19541), .A(n19525), .B(n19524), .ZN(
        P2_U3129) );
  AOI22_X1 U22561 ( .A1(n19537), .A2(n19228), .B1(n19712), .B2(n19536), .ZN(
        n19527) );
  AOI22_X1 U22562 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19538), .B1(
        n19569), .B2(n19713), .ZN(n19526) );
  OAI211_X1 U22563 ( .C1(n19716), .C2(n19541), .A(n19527), .B(n19526), .ZN(
        P2_U3130) );
  AOI22_X1 U22564 ( .A1(n19537), .A2(n19718), .B1(n19717), .B2(n19536), .ZN(
        n19529) );
  AOI22_X1 U22565 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19538), .B1(
        n19569), .B2(n19719), .ZN(n19528) );
  OAI211_X1 U22566 ( .C1(n19722), .C2(n19541), .A(n19529), .B(n19528), .ZN(
        P2_U3131) );
  AOI22_X1 U22567 ( .A1(n19537), .A2(n19724), .B1(n19723), .B2(n19536), .ZN(
        n19531) );
  AOI22_X1 U22568 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19538), .B1(
        n19569), .B2(n19725), .ZN(n19530) );
  OAI211_X1 U22569 ( .C1(n19728), .C2(n19541), .A(n19531), .B(n19530), .ZN(
        P2_U3132) );
  AOI22_X1 U22570 ( .A1(n19537), .A2(n19730), .B1(n19729), .B2(n19536), .ZN(
        n19533) );
  AOI22_X1 U22571 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19538), .B1(
        n19569), .B2(n19731), .ZN(n19532) );
  OAI211_X1 U22572 ( .C1(n19734), .C2(n19541), .A(n19533), .B(n19532), .ZN(
        P2_U3133) );
  AOI22_X1 U22573 ( .A1(n19537), .A2(n19736), .B1(n19735), .B2(n19536), .ZN(
        n19535) );
  AOI22_X1 U22574 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19538), .B1(
        n19569), .B2(n19737), .ZN(n19534) );
  OAI211_X1 U22575 ( .C1(n19740), .C2(n19541), .A(n19535), .B(n19534), .ZN(
        P2_U3134) );
  AOI22_X1 U22576 ( .A1(n19537), .A2(n19743), .B1(n19741), .B2(n19536), .ZN(
        n19540) );
  AOI22_X1 U22577 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19538), .B1(
        n19569), .B2(n19745), .ZN(n19539) );
  OAI211_X1 U22578 ( .C1(n19751), .C2(n19541), .A(n19540), .B(n19539), .ZN(
        P2_U3135) );
  NAND2_X1 U22579 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19542), .ZN(
        n19550) );
  INV_X1 U22580 ( .A(n19550), .ZN(n19543) );
  NAND2_X1 U22581 ( .A1(n19543), .A2(n19697), .ZN(n19547) );
  INV_X1 U22582 ( .A(n10062), .ZN(n19546) );
  NOR2_X1 U22583 ( .A1(n19545), .A2(n19544), .ZN(n19567) );
  NOR3_X1 U22584 ( .A1(n19546), .A2(n19567), .A3(n19691), .ZN(n19549) );
  AOI21_X1 U22585 ( .B1(n19691), .B2(n19547), .A(n19549), .ZN(n19568) );
  AOI22_X1 U22586 ( .A1(n19568), .A2(n15506), .B1(n19694), .B2(n19567), .ZN(
        n19554) );
  NAND2_X1 U22587 ( .A1(n19700), .A2(n19548), .ZN(n19551) );
  AOI21_X1 U22588 ( .B1(n19551), .B2(n19550), .A(n19549), .ZN(n19552) );
  OAI211_X1 U22589 ( .C1(n19567), .C2(n19697), .A(n19552), .B(n19695), .ZN(
        n19570) );
  AOI22_X1 U22590 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19570), .B1(
        n19569), .B2(n19647), .ZN(n19553) );
  OAI211_X1 U22591 ( .C1(n19660), .C2(n19573), .A(n19554), .B(n19553), .ZN(
        P2_U3136) );
  AOI22_X1 U22592 ( .A1(n19568), .A2(n19224), .B1(n19707), .B2(n19567), .ZN(
        n19556) );
  AOI22_X1 U22593 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19570), .B1(
        n19569), .B2(n19661), .ZN(n19555) );
  OAI211_X1 U22594 ( .C1(n19664), .C2(n19573), .A(n19556), .B(n19555), .ZN(
        P2_U3137) );
  AOI22_X1 U22595 ( .A1(n19568), .A2(n19228), .B1(n19712), .B2(n19567), .ZN(
        n19558) );
  AOI22_X1 U22596 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19570), .B1(
        n19569), .B2(n19623), .ZN(n19557) );
  OAI211_X1 U22597 ( .C1(n19626), .C2(n19573), .A(n19558), .B(n19557), .ZN(
        P2_U3138) );
  AOI22_X1 U22598 ( .A1(n19568), .A2(n19718), .B1(n19717), .B2(n19567), .ZN(
        n19560) );
  AOI22_X1 U22599 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19570), .B1(
        n19569), .B2(n19627), .ZN(n19559) );
  OAI211_X1 U22600 ( .C1(n19630), .C2(n19573), .A(n19560), .B(n19559), .ZN(
        P2_U3139) );
  AOI22_X1 U22601 ( .A1(n19568), .A2(n19724), .B1(n19723), .B2(n19567), .ZN(
        n19562) );
  AOI22_X1 U22602 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19570), .B1(
        n19569), .B2(n19631), .ZN(n19561) );
  OAI211_X1 U22603 ( .C1(n19634), .C2(n19573), .A(n19562), .B(n19561), .ZN(
        P2_U3140) );
  AOI22_X1 U22604 ( .A1(n19568), .A2(n19730), .B1(n19729), .B2(n19567), .ZN(
        n19564) );
  AOI22_X1 U22605 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19570), .B1(
        n19569), .B2(n19671), .ZN(n19563) );
  OAI211_X1 U22606 ( .C1(n19674), .C2(n19573), .A(n19564), .B(n19563), .ZN(
        P2_U3141) );
  AOI22_X1 U22607 ( .A1(n19568), .A2(n19736), .B1(n19735), .B2(n19567), .ZN(
        n19566) );
  AOI22_X1 U22608 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19570), .B1(
        n19569), .B2(n19676), .ZN(n19565) );
  OAI211_X1 U22609 ( .C1(n19679), .C2(n19573), .A(n19566), .B(n19565), .ZN(
        P2_U3142) );
  AOI22_X1 U22610 ( .A1(n19568), .A2(n19743), .B1(n19741), .B2(n19567), .ZN(
        n19572) );
  AOI22_X1 U22611 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19570), .B1(
        n19569), .B2(n19602), .ZN(n19571) );
  OAI211_X1 U22612 ( .C1(n19607), .C2(n19573), .A(n19572), .B(n19571), .ZN(
        P2_U3143) );
  AOI21_X1 U22613 ( .B1(n19644), .B2(n19573), .A(n19896), .ZN(n19574) );
  AOI21_X1 U22614 ( .B1(n19580), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n19574), .ZN(n19578) );
  NAND3_X1 U22615 ( .A1(n19873), .A2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19611) );
  NOR2_X1 U22616 ( .A1(n19611), .A2(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n19600) );
  INV_X1 U22617 ( .A(n19600), .ZN(n19575) );
  OAI211_X1 U22618 ( .C1(n10422), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19575), 
        .B(n19650), .ZN(n19576) );
  NAND2_X1 U22619 ( .A1(n19576), .A2(n19695), .ZN(n19577) );
  INV_X1 U22620 ( .A(n19604), .ZN(n19589) );
  INV_X1 U22621 ( .A(n19579), .ZN(n19584) );
  INV_X1 U22622 ( .A(n19580), .ZN(n19583) );
  INV_X1 U22623 ( .A(n10422), .ZN(n19581) );
  OAI21_X1 U22624 ( .B1(n19581), .B2(n19600), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19582) );
  OAI21_X1 U22625 ( .B1(n19584), .B2(n19583), .A(n19582), .ZN(n19601) );
  AOI22_X1 U22626 ( .A1(n19601), .A2(n15506), .B1(n19694), .B2(n19600), .ZN(
        n19586) );
  AOI22_X1 U22627 ( .A1(n19603), .A2(n19647), .B1(n19635), .B2(n19703), .ZN(
        n19585) );
  OAI211_X1 U22628 ( .C1(n19589), .C2(n11504), .A(n19586), .B(n19585), .ZN(
        P2_U3144) );
  AOI22_X1 U22629 ( .A1(n19601), .A2(n19224), .B1(n19707), .B2(n19600), .ZN(
        n19588) );
  AOI22_X1 U22630 ( .A1(n19603), .A2(n19661), .B1(n19635), .B2(n19708), .ZN(
        n19587) );
  OAI211_X1 U22631 ( .C1(n19589), .C2(n11347), .A(n19588), .B(n19587), .ZN(
        P2_U3145) );
  AOI22_X1 U22632 ( .A1(n19601), .A2(n19228), .B1(n19712), .B2(n19600), .ZN(
        n19591) );
  AOI22_X1 U22633 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19604), .B1(
        n19603), .B2(n19623), .ZN(n19590) );
  OAI211_X1 U22634 ( .C1(n19626), .C2(n19644), .A(n19591), .B(n19590), .ZN(
        P2_U3146) );
  AOI22_X1 U22635 ( .A1(n19601), .A2(n19718), .B1(n19717), .B2(n19600), .ZN(
        n19593) );
  AOI22_X1 U22636 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19604), .B1(
        n19603), .B2(n19627), .ZN(n19592) );
  OAI211_X1 U22637 ( .C1(n19630), .C2(n19644), .A(n19593), .B(n19592), .ZN(
        P2_U3147) );
  AOI22_X1 U22638 ( .A1(n19601), .A2(n19724), .B1(n19723), .B2(n19600), .ZN(
        n19595) );
  AOI22_X1 U22639 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19604), .B1(
        n19603), .B2(n19631), .ZN(n19594) );
  OAI211_X1 U22640 ( .C1(n19634), .C2(n19644), .A(n19595), .B(n19594), .ZN(
        P2_U3148) );
  AOI22_X1 U22641 ( .A1(n19601), .A2(n19730), .B1(n19729), .B2(n19600), .ZN(
        n19597) );
  AOI22_X1 U22642 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19604), .B1(
        n19603), .B2(n19671), .ZN(n19596) );
  OAI211_X1 U22643 ( .C1(n19674), .C2(n19644), .A(n19597), .B(n19596), .ZN(
        P2_U3149) );
  AOI22_X1 U22644 ( .A1(n19601), .A2(n19736), .B1(n19735), .B2(n19600), .ZN(
        n19599) );
  AOI22_X1 U22645 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19604), .B1(
        n19603), .B2(n19676), .ZN(n19598) );
  OAI211_X1 U22646 ( .C1(n19679), .C2(n19644), .A(n19599), .B(n19598), .ZN(
        P2_U3150) );
  AOI22_X1 U22647 ( .A1(n19601), .A2(n19743), .B1(n19741), .B2(n19600), .ZN(
        n19606) );
  AOI22_X1 U22648 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19604), .B1(
        n19603), .B2(n19602), .ZN(n19605) );
  OAI211_X1 U22649 ( .C1(n19607), .C2(n19644), .A(n19606), .B(n19605), .ZN(
        P2_U3151) );
  INV_X1 U22650 ( .A(n10426), .ZN(n19610) );
  NOR2_X1 U22651 ( .A1(n19880), .A2(n19611), .ZN(n19649) );
  NOR3_X1 U22652 ( .A1(n19610), .A2(n19649), .A3(n19691), .ZN(n19613) );
  INV_X1 U22653 ( .A(n19611), .ZN(n19618) );
  AOI21_X1 U22654 ( .B1(n19697), .B2(n19618), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19612) );
  NOR2_X1 U22655 ( .A1(n19613), .A2(n19612), .ZN(n19640) );
  AOI22_X1 U22656 ( .A1(n19640), .A2(n15506), .B1(n19694), .B2(n19649), .ZN(
        n19620) );
  INV_X1 U22657 ( .A(n19649), .ZN(n19615) );
  AOI211_X1 U22658 ( .C1(P2_STATE2_REG_3__SCAN_IN), .C2(n19615), .A(n19614), 
        .B(n19613), .ZN(n19616) );
  OAI221_X1 U22659 ( .B1(n19618), .B2(n19617), .C1(n19618), .C2(n19700), .A(
        n19616), .ZN(n19641) );
  AOI22_X1 U22660 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19641), .B1(
        n19635), .B2(n19647), .ZN(n19619) );
  OAI211_X1 U22661 ( .C1(n19660), .C2(n19686), .A(n19620), .B(n19619), .ZN(
        P2_U3152) );
  AOI22_X1 U22662 ( .A1(n19640), .A2(n19224), .B1(n19707), .B2(n19649), .ZN(
        n19622) );
  AOI22_X1 U22663 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19641), .B1(
        n19675), .B2(n19708), .ZN(n19621) );
  OAI211_X1 U22664 ( .C1(n19711), .C2(n19644), .A(n19622), .B(n19621), .ZN(
        P2_U3153) );
  AOI22_X1 U22665 ( .A1(n19640), .A2(n19228), .B1(n19712), .B2(n19649), .ZN(
        n19625) );
  AOI22_X1 U22666 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19641), .B1(
        n19635), .B2(n19623), .ZN(n19624) );
  OAI211_X1 U22667 ( .C1(n19626), .C2(n19686), .A(n19625), .B(n19624), .ZN(
        P2_U3154) );
  AOI22_X1 U22668 ( .A1(n19640), .A2(n19718), .B1(n19717), .B2(n19649), .ZN(
        n19629) );
  AOI22_X1 U22669 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19641), .B1(
        n19635), .B2(n19627), .ZN(n19628) );
  OAI211_X1 U22670 ( .C1(n19630), .C2(n19686), .A(n19629), .B(n19628), .ZN(
        P2_U3155) );
  AOI22_X1 U22671 ( .A1(n19640), .A2(n19724), .B1(n19723), .B2(n19649), .ZN(
        n19633) );
  AOI22_X1 U22672 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19641), .B1(
        n19635), .B2(n19631), .ZN(n19632) );
  OAI211_X1 U22673 ( .C1(n19634), .C2(n19686), .A(n19633), .B(n19632), .ZN(
        P2_U3156) );
  AOI22_X1 U22674 ( .A1(n19640), .A2(n19730), .B1(n19729), .B2(n19649), .ZN(
        n19637) );
  AOI22_X1 U22675 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19641), .B1(
        n19635), .B2(n19671), .ZN(n19636) );
  OAI211_X1 U22676 ( .C1(n19674), .C2(n19686), .A(n19637), .B(n19636), .ZN(
        P2_U3157) );
  AOI22_X1 U22677 ( .A1(n19640), .A2(n19736), .B1(n19735), .B2(n19649), .ZN(
        n19639) );
  AOI22_X1 U22678 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19641), .B1(
        n19675), .B2(n19737), .ZN(n19638) );
  OAI211_X1 U22679 ( .C1(n19740), .C2(n19644), .A(n19639), .B(n19638), .ZN(
        P2_U3158) );
  AOI22_X1 U22680 ( .A1(n19640), .A2(n19743), .B1(n19741), .B2(n19649), .ZN(
        n19643) );
  AOI22_X1 U22681 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19641), .B1(
        n19675), .B2(n19745), .ZN(n19642) );
  OAI211_X1 U22682 ( .C1(n19751), .C2(n19644), .A(n19643), .B(n19642), .ZN(
        P2_U3159) );
  NOR3_X2 U22683 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19856), .A3(
        n19690), .ZN(n19680) );
  AOI22_X1 U22684 ( .A1(n19647), .A2(n19675), .B1(n19694), .B2(n19680), .ZN(
        n19659) );
  NOR2_X1 U22685 ( .A1(n19681), .A2(n19675), .ZN(n19648) );
  OAI21_X1 U22686 ( .B1(n19648), .B2(n19896), .A(n19844), .ZN(n19657) );
  NOR2_X1 U22687 ( .A1(n19680), .A2(n19649), .ZN(n19656) );
  INV_X1 U22688 ( .A(n19656), .ZN(n19653) );
  INV_X1 U22689 ( .A(n19680), .ZN(n19651) );
  OAI211_X1 U22690 ( .C1(n10421), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19651), 
        .B(n19650), .ZN(n19652) );
  OAI211_X1 U22691 ( .C1(n19657), .C2(n19653), .A(n19695), .B(n19652), .ZN(
        n19683) );
  OAI21_X1 U22692 ( .B1(n19654), .B2(n19680), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19655) );
  AOI22_X1 U22693 ( .A1(P2_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n19683), .B1(
        n15506), .B2(n19682), .ZN(n19658) );
  OAI211_X1 U22694 ( .C1(n19660), .C2(n19750), .A(n19659), .B(n19658), .ZN(
        P2_U3160) );
  AOI22_X1 U22695 ( .A1(n19661), .A2(n19675), .B1(n19707), .B2(n19680), .ZN(
        n19663) );
  AOI22_X1 U22696 ( .A1(P2_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n19683), .B1(
        n19224), .B2(n19682), .ZN(n19662) );
  OAI211_X1 U22697 ( .C1(n19664), .C2(n19750), .A(n19663), .B(n19662), .ZN(
        P2_U3161) );
  AOI22_X1 U22698 ( .A1(n19713), .A2(n19681), .B1(n19712), .B2(n19680), .ZN(
        n19666) );
  AOI22_X1 U22699 ( .A1(P2_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n19683), .B1(
        n19228), .B2(n19682), .ZN(n19665) );
  OAI211_X1 U22700 ( .C1(n19716), .C2(n19686), .A(n19666), .B(n19665), .ZN(
        P2_U3162) );
  AOI22_X1 U22701 ( .A1(n19719), .A2(n19681), .B1(n19717), .B2(n19680), .ZN(
        n19668) );
  AOI22_X1 U22702 ( .A1(P2_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n19683), .B1(
        n19718), .B2(n19682), .ZN(n19667) );
  OAI211_X1 U22703 ( .C1(n19722), .C2(n19686), .A(n19668), .B(n19667), .ZN(
        P2_U3163) );
  AOI22_X1 U22704 ( .A1(n19725), .A2(n19681), .B1(n19723), .B2(n19680), .ZN(
        n19670) );
  AOI22_X1 U22705 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n19683), .B1(
        n19724), .B2(n19682), .ZN(n19669) );
  OAI211_X1 U22706 ( .C1(n19728), .C2(n19686), .A(n19670), .B(n19669), .ZN(
        P2_U3164) );
  AOI22_X1 U22707 ( .A1(n19671), .A2(n19675), .B1(n19729), .B2(n19680), .ZN(
        n19673) );
  AOI22_X1 U22708 ( .A1(P2_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n19683), .B1(
        n19730), .B2(n19682), .ZN(n19672) );
  OAI211_X1 U22709 ( .C1(n19674), .C2(n19750), .A(n19673), .B(n19672), .ZN(
        P2_U3165) );
  AOI22_X1 U22710 ( .A1(n19676), .A2(n19675), .B1(n19735), .B2(n19680), .ZN(
        n19678) );
  AOI22_X1 U22711 ( .A1(P2_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n19683), .B1(
        n19736), .B2(n19682), .ZN(n19677) );
  OAI211_X1 U22712 ( .C1(n19679), .C2(n19750), .A(n19678), .B(n19677), .ZN(
        P2_U3166) );
  AOI22_X1 U22713 ( .A1(n19681), .A2(n19745), .B1(n19741), .B2(n19680), .ZN(
        n19685) );
  AOI22_X1 U22714 ( .A1(P2_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n19683), .B1(
        n19743), .B2(n19682), .ZN(n19684) );
  OAI211_X1 U22715 ( .C1(n19751), .C2(n19686), .A(n19685), .B(n19684), .ZN(
        P2_U3167) );
  AND2_X1 U22716 ( .A1(n19687), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19688) );
  NAND2_X1 U22717 ( .A1(n19689), .A2(n19688), .ZN(n19696) );
  NOR2_X1 U22718 ( .A1(n19856), .A2(n19690), .ZN(n19702) );
  INV_X1 U22719 ( .A(n19702), .ZN(n19692) );
  OAI21_X1 U22720 ( .B1(n19692), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19691), 
        .ZN(n19693) );
  AND2_X1 U22721 ( .A1(n19696), .A2(n19693), .ZN(n19744) );
  AOI22_X1 U22722 ( .A1(n19744), .A2(n15506), .B1(n19742), .B2(n19694), .ZN(
        n19705) );
  OAI211_X1 U22723 ( .C1(n19742), .C2(n19697), .A(n19696), .B(n19695), .ZN(
        n19698) );
  INV_X1 U22724 ( .A(n19698), .ZN(n19699) );
  OAI221_X1 U22725 ( .B1(n19702), .B2(n19701), .C1(n19702), .C2(n19700), .A(
        n19699), .ZN(n19747) );
  AOI22_X1 U22726 ( .A1(P2_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n19747), .B1(
        n19746), .B2(n19703), .ZN(n19704) );
  OAI211_X1 U22727 ( .C1(n19706), .C2(n19750), .A(n19705), .B(n19704), .ZN(
        P2_U3168) );
  AOI22_X1 U22728 ( .A1(n19744), .A2(n19224), .B1(n19742), .B2(n19707), .ZN(
        n19710) );
  AOI22_X1 U22729 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n19747), .B1(
        n19746), .B2(n19708), .ZN(n19709) );
  OAI211_X1 U22730 ( .C1(n19711), .C2(n19750), .A(n19710), .B(n19709), .ZN(
        P2_U3169) );
  AOI22_X1 U22731 ( .A1(n19744), .A2(n19228), .B1(n19742), .B2(n19712), .ZN(
        n19715) );
  AOI22_X1 U22732 ( .A1(P2_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n19747), .B1(
        n19746), .B2(n19713), .ZN(n19714) );
  OAI211_X1 U22733 ( .C1(n19716), .C2(n19750), .A(n19715), .B(n19714), .ZN(
        P2_U3170) );
  AOI22_X1 U22734 ( .A1(n19744), .A2(n19718), .B1(n19742), .B2(n19717), .ZN(
        n19721) );
  AOI22_X1 U22735 ( .A1(P2_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n19747), .B1(
        n19746), .B2(n19719), .ZN(n19720) );
  OAI211_X1 U22736 ( .C1(n19722), .C2(n19750), .A(n19721), .B(n19720), .ZN(
        P2_U3171) );
  AOI22_X1 U22737 ( .A1(n19744), .A2(n19724), .B1(n19742), .B2(n19723), .ZN(
        n19727) );
  AOI22_X1 U22738 ( .A1(P2_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n19747), .B1(
        n19746), .B2(n19725), .ZN(n19726) );
  OAI211_X1 U22739 ( .C1(n19728), .C2(n19750), .A(n19727), .B(n19726), .ZN(
        P2_U3172) );
  AOI22_X1 U22740 ( .A1(n19744), .A2(n19730), .B1(n19742), .B2(n19729), .ZN(
        n19733) );
  AOI22_X1 U22741 ( .A1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n19747), .B1(
        n19746), .B2(n19731), .ZN(n19732) );
  OAI211_X1 U22742 ( .C1(n19734), .C2(n19750), .A(n19733), .B(n19732), .ZN(
        P2_U3173) );
  AOI22_X1 U22743 ( .A1(n19744), .A2(n19736), .B1(n19742), .B2(n19735), .ZN(
        n19739) );
  AOI22_X1 U22744 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n19747), .B1(
        n19746), .B2(n19737), .ZN(n19738) );
  OAI211_X1 U22745 ( .C1(n19740), .C2(n19750), .A(n19739), .B(n19738), .ZN(
        P2_U3174) );
  AOI22_X1 U22746 ( .A1(n19744), .A2(n19743), .B1(n19742), .B2(n19741), .ZN(
        n19749) );
  AOI22_X1 U22747 ( .A1(P2_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n19747), .B1(
        n19746), .B2(n19745), .ZN(n19748) );
  OAI211_X1 U22748 ( .C1(n19751), .C2(n19750), .A(n19749), .B(n19748), .ZN(
        P2_U3175) );
  OR3_X1 U22749 ( .A1(n19754), .A2(n19753), .A3(n19752), .ZN(n19755) );
  OAI221_X1 U22750 ( .B1(n15828), .B2(n19757), .C1(n15828), .C2(n19756), .A(
        n19755), .ZN(P2_U3177) );
  AND2_X1 U22751 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19758), .ZN(
        P2_U3179) );
  AND2_X1 U22752 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19758), .ZN(
        P2_U3180) );
  AND2_X1 U22753 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19758), .ZN(
        P2_U3181) );
  AND2_X1 U22754 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19758), .ZN(
        P2_U3182) );
  AND2_X1 U22755 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19758), .ZN(
        P2_U3183) );
  AND2_X1 U22756 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19758), .ZN(
        P2_U3184) );
  AND2_X1 U22757 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19758), .ZN(
        P2_U3185) );
  AND2_X1 U22758 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(n19758), .ZN(
        P2_U3186) );
  AND2_X1 U22759 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19758), .ZN(
        P2_U3187) );
  AND2_X1 U22760 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19758), .ZN(
        P2_U3188) );
  AND2_X1 U22761 ( .A1(P2_DATAWIDTH_REG_21__SCAN_IN), .A2(n19758), .ZN(
        P2_U3189) );
  AND2_X1 U22762 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19758), .ZN(
        P2_U3190) );
  AND2_X1 U22763 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19758), .ZN(
        P2_U3191) );
  AND2_X1 U22764 ( .A1(P2_DATAWIDTH_REG_18__SCAN_IN), .A2(n19758), .ZN(
        P2_U3192) );
  AND2_X1 U22765 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19758), .ZN(
        P2_U3193) );
  AND2_X1 U22766 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19758), .ZN(
        P2_U3194) );
  AND2_X1 U22767 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19758), .ZN(
        P2_U3195) );
  AND2_X1 U22768 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19758), .ZN(
        P2_U3196) );
  AND2_X1 U22769 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19758), .ZN(
        P2_U3197) );
  AND2_X1 U22770 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19758), .ZN(
        P2_U3198) );
  AND2_X1 U22771 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19758), .ZN(
        P2_U3199) );
  AND2_X1 U22772 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19758), .ZN(
        P2_U3200) );
  AND2_X1 U22773 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19758), .ZN(P2_U3201) );
  AND2_X1 U22774 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19758), .ZN(P2_U3202) );
  AND2_X1 U22775 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19758), .ZN(P2_U3203) );
  AND2_X1 U22776 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19758), .ZN(P2_U3204) );
  AND2_X1 U22777 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19758), .ZN(P2_U3205) );
  AND2_X1 U22778 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(n19758), .ZN(P2_U3206) );
  AND2_X1 U22779 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19758), .ZN(P2_U3207) );
  AND2_X1 U22780 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19758), .ZN(P2_U3208) );
  INV_X1 U22781 ( .A(NA), .ZN(n20682) );
  OAI21_X1 U22782 ( .B1(n20682), .B2(n19765), .A(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19775) );
  INV_X1 U22783 ( .A(n19775), .ZN(n19762) );
  NOR2_X1 U22784 ( .A1(n19759), .A2(n19898), .ZN(n19769) );
  INV_X1 U22785 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19904) );
  NOR3_X1 U22786 ( .A1(n19769), .A2(n19904), .A3(n19764), .ZN(n19761) );
  OAI211_X1 U22787 ( .C1(HOLD), .C2(n19904), .A(n19906), .B(n19770), .ZN(
        n19760) );
  OAI21_X1 U22788 ( .B1(n19762), .B2(n19761), .A(n19760), .ZN(P2_U3209) );
  NOR2_X1 U22789 ( .A1(n19763), .A2(n19769), .ZN(n19767) );
  NOR2_X1 U22790 ( .A1(HOLD), .A2(n19764), .ZN(n19774) );
  OAI211_X1 U22791 ( .C1(n19774), .C2(n19776), .A(
        P2_REQUESTPENDING_REG_SCAN_IN), .B(n19765), .ZN(n19766) );
  OAI211_X1 U22792 ( .C1(n19768), .C2(n20687), .A(n19767), .B(n19766), .ZN(
        P2_U3210) );
  INV_X1 U22793 ( .A(n19769), .ZN(n19773) );
  OAI22_X1 U22794 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19770), .B1(NA), 
        .B2(n19773), .ZN(n19771) );
  OAI211_X1 U22795 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19771), .ZN(n19772) );
  OAI221_X1 U22796 ( .B1(n19775), .B2(n19774), .C1(n19775), .C2(n19773), .A(
        n19772), .ZN(P2_U3211) );
  INV_X1 U22797 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n19779) );
  OAI222_X1 U22798 ( .A1(n19835), .A2(n19779), .B1(n19778), .B2(n19833), .C1(
        n19777), .C2(n19831), .ZN(P2_U3212) );
  OAI222_X1 U22799 ( .A1(n19835), .A2(n19781), .B1(n19780), .B2(n19833), .C1(
        n19779), .C2(n19831), .ZN(P2_U3213) );
  OAI222_X1 U22800 ( .A1(n19835), .A2(n19783), .B1(n19782), .B2(n19833), .C1(
        n19781), .C2(n19831), .ZN(P2_U3214) );
  OAI222_X1 U22801 ( .A1(n19835), .A2(n13716), .B1(n19784), .B2(n19833), .C1(
        n19783), .C2(n19831), .ZN(P2_U3215) );
  OAI222_X1 U22802 ( .A1(n19835), .A2(n19786), .B1(n19785), .B2(n19833), .C1(
        n13716), .C2(n19831), .ZN(P2_U3216) );
  OAI222_X1 U22803 ( .A1(n19835), .A2(n19787), .B1(n20951), .B2(n19839), .C1(
        n19786), .C2(n19831), .ZN(P2_U3217) );
  INV_X1 U22804 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n19789) );
  OAI222_X1 U22805 ( .A1(n19835), .A2(n19789), .B1(n19788), .B2(n19833), .C1(
        n19787), .C2(n19831), .ZN(P2_U3218) );
  OAI222_X1 U22806 ( .A1(n19835), .A2(n19791), .B1(n19790), .B2(n19833), .C1(
        n19789), .C2(n19831), .ZN(P2_U3219) );
  OAI222_X1 U22807 ( .A1(n19835), .A2(n19793), .B1(n19792), .B2(n19833), .C1(
        n19791), .C2(n19831), .ZN(P2_U3220) );
  OAI222_X1 U22808 ( .A1(n19835), .A2(n19795), .B1(n19794), .B2(n19833), .C1(
        n19793), .C2(n19831), .ZN(P2_U3221) );
  INV_X1 U22809 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n19797) );
  OAI222_X1 U22810 ( .A1(n19835), .A2(n19797), .B1(n19796), .B2(n19839), .C1(
        n19795), .C2(n19831), .ZN(P2_U3222) );
  OAI222_X1 U22811 ( .A1(n19835), .A2(n19799), .B1(n19798), .B2(n19839), .C1(
        n19797), .C2(n19831), .ZN(P2_U3223) );
  OAI222_X1 U22812 ( .A1(n19835), .A2(n19801), .B1(n19800), .B2(n19839), .C1(
        n19799), .C2(n19831), .ZN(P2_U3224) );
  OAI222_X1 U22813 ( .A1(n19835), .A2(n19803), .B1(n19802), .B2(n19839), .C1(
        n19801), .C2(n19831), .ZN(P2_U3225) );
  OAI222_X1 U22814 ( .A1(n19835), .A2(n15142), .B1(n19804), .B2(n19839), .C1(
        n19803), .C2(n19831), .ZN(P2_U3226) );
  INV_X1 U22815 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19806) );
  OAI222_X1 U22816 ( .A1(n19835), .A2(n19806), .B1(n19805), .B2(n19839), .C1(
        n15142), .C2(n19831), .ZN(P2_U3227) );
  INV_X1 U22817 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19808) );
  OAI222_X1 U22818 ( .A1(n19835), .A2(n19808), .B1(n19807), .B2(n19839), .C1(
        n19806), .C2(n19831), .ZN(P2_U3228) );
  OAI222_X1 U22819 ( .A1(n19835), .A2(n19810), .B1(n19809), .B2(n19839), .C1(
        n19808), .C2(n19831), .ZN(P2_U3229) );
  INV_X1 U22820 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19812) );
  OAI222_X1 U22821 ( .A1(n19835), .A2(n19812), .B1(n19811), .B2(n19839), .C1(
        n19810), .C2(n19831), .ZN(P2_U3230) );
  OAI222_X1 U22822 ( .A1(n19835), .A2(n19814), .B1(n19813), .B2(n19839), .C1(
        n19812), .C2(n19831), .ZN(P2_U3231) );
  OAI222_X1 U22823 ( .A1(n19835), .A2(n19816), .B1(n19815), .B2(n19839), .C1(
        n19814), .C2(n19831), .ZN(P2_U3232) );
  OAI222_X1 U22824 ( .A1(n19835), .A2(n19818), .B1(n19817), .B2(n19839), .C1(
        n19816), .C2(n19831), .ZN(P2_U3233) );
  OAI222_X1 U22825 ( .A1(n19835), .A2(n19820), .B1(n19819), .B2(n19833), .C1(
        n19818), .C2(n19831), .ZN(P2_U3234) );
  INV_X1 U22826 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19822) );
  OAI222_X1 U22827 ( .A1(n19835), .A2(n19822), .B1(n19821), .B2(n19833), .C1(
        n19820), .C2(n19831), .ZN(P2_U3235) );
  INV_X1 U22828 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n19824) );
  OAI222_X1 U22829 ( .A1(n19835), .A2(n19824), .B1(n19823), .B2(n19833), .C1(
        n19822), .C2(n19831), .ZN(P2_U3236) );
  INV_X1 U22830 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19827) );
  OAI222_X1 U22831 ( .A1(n19835), .A2(n19827), .B1(n19825), .B2(n19833), .C1(
        n19824), .C2(n19831), .ZN(P2_U3237) );
  OAI222_X1 U22832 ( .A1(n19831), .A2(n19827), .B1(n19826), .B2(n19833), .C1(
        n19828), .C2(n19835), .ZN(P2_U3238) );
  INV_X1 U22833 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n20939) );
  OAI222_X1 U22834 ( .A1(n19835), .A2(n20939), .B1(n19829), .B2(n19833), .C1(
        n19828), .C2(n19831), .ZN(P2_U3239) );
  OAI222_X1 U22835 ( .A1(n19835), .A2(n19832), .B1(n19830), .B2(n19833), .C1(
        n20939), .C2(n19831), .ZN(P2_U3240) );
  OAI222_X1 U22836 ( .A1(n19835), .A2(n16125), .B1(n19834), .B2(n19833), .C1(
        n19832), .C2(n19831), .ZN(P2_U3241) );
  OAI22_X1 U22837 ( .A1(n19906), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19839), .ZN(n19836) );
  INV_X1 U22838 ( .A(n19836), .ZN(P2_U3585) );
  OAI22_X1 U22839 ( .A1(n19906), .A2(P2_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P2_BE_N_REG_2__SCAN_IN), .B2(n19839), .ZN(n19837) );
  INV_X1 U22840 ( .A(n19837), .ZN(P2_U3586) );
  OAI22_X1 U22841 ( .A1(n19906), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19833), .ZN(n19838) );
  INV_X1 U22842 ( .A(n19838), .ZN(P2_U3587) );
  INV_X1 U22843 ( .A(P2_BE_N_REG_0__SCAN_IN), .ZN(n20924) );
  AOI22_X1 U22844 ( .A1(n19839), .A2(n20923), .B1(n20924), .B2(n19906), .ZN(
        P2_U3588) );
  OAI21_X1 U22845 ( .B1(n19843), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19841), 
        .ZN(n19840) );
  INV_X1 U22846 ( .A(n19840), .ZN(P2_U3591) );
  OAI21_X1 U22847 ( .B1(n19843), .B2(n19842), .A(n19841), .ZN(P2_U3592) );
  INV_X1 U22848 ( .A(n19878), .ZN(n19881) );
  NAND2_X1 U22849 ( .A1(n19845), .A2(n19844), .ZN(n19854) );
  INV_X1 U22850 ( .A(n19846), .ZN(n19869) );
  OR2_X1 U22851 ( .A1(n19847), .A2(n19869), .ZN(n19857) );
  NAND3_X1 U22852 ( .A1(n19870), .A2(n19848), .A3(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19849) );
  NAND2_X1 U22853 ( .A1(n19849), .A2(n19876), .ZN(n19858) );
  NAND2_X1 U22854 ( .A1(n19857), .A2(n19858), .ZN(n19852) );
  AOI22_X1 U22855 ( .A1(n19852), .A2(n19851), .B1(P2_STATE2_REG_3__SCAN_IN), 
        .B2(n19850), .ZN(n19853) );
  AND2_X1 U22856 ( .A1(n19854), .A2(n19853), .ZN(n19855) );
  AOI22_X1 U22857 ( .A1(n19881), .A2(n19856), .B1(n19855), .B2(n19878), .ZN(
        P2_U3602) );
  OAI21_X1 U22858 ( .B1(n19859), .B2(n19858), .A(n19857), .ZN(n19860) );
  AOI21_X1 U22859 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19861), .A(n19860), 
        .ZN(n19862) );
  AOI22_X1 U22860 ( .A1(n19881), .A2(n19863), .B1(n19862), .B2(n19878), .ZN(
        P2_U3603) );
  INV_X1 U22861 ( .A(n19864), .ZN(n19865) );
  NAND3_X1 U22862 ( .A1(n19870), .A2(n19876), .A3(n19865), .ZN(n19868) );
  NAND2_X1 U22863 ( .A1(n19866), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19867) );
  OAI211_X1 U22864 ( .C1(n19870), .C2(n19869), .A(n19868), .B(n19867), .ZN(
        n19871) );
  INV_X1 U22865 ( .A(n19871), .ZN(n19872) );
  AOI22_X1 U22866 ( .A1(n19881), .A2(n19873), .B1(n19872), .B2(n19878), .ZN(
        P2_U3604) );
  AOI211_X1 U22867 ( .C1(n19877), .C2(n19876), .A(n19875), .B(n19874), .ZN(
        n19879) );
  AOI22_X1 U22868 ( .A1(n19881), .A2(n19880), .B1(n19879), .B2(n19878), .ZN(
        P2_U3605) );
  INV_X1 U22869 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19882) );
  AOI22_X1 U22870 ( .A1(n19839), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19882), 
        .B2(n19906), .ZN(P2_U3608) );
  INV_X1 U22871 ( .A(n19883), .ZN(n19889) );
  OR3_X1 U22872 ( .A1(n10745), .A2(n19885), .A3(n19884), .ZN(n19886) );
  OAI211_X1 U22873 ( .C1(n19889), .C2(n19888), .A(n19887), .B(n19886), .ZN(
        n19891) );
  MUX2_X1 U22874 ( .A(P2_MORE_REG_SCAN_IN), .B(n19891), .S(n19890), .Z(
        P2_U3609) );
  AOI21_X1 U22875 ( .B1(n19181), .B2(n19898), .A(n19892), .ZN(n19893) );
  OAI21_X1 U22876 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19894), .A(n19893), 
        .ZN(n19905) );
  AOI21_X1 U22877 ( .B1(n19897), .B2(n19896), .A(n19895), .ZN(n19900) );
  OAI211_X1 U22878 ( .C1(n19900), .C2(n19899), .A(P2_STATE2_REG_2__SCAN_IN), 
        .B(n19898), .ZN(n19901) );
  NAND3_X1 U22879 ( .A1(n19905), .A2(n19902), .A3(n19901), .ZN(n19903) );
  OAI21_X1 U22880 ( .B1(n19905), .B2(n19904), .A(n19903), .ZN(P2_U3610) );
  OAI22_X1 U22881 ( .A1(n19906), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19833), .ZN(n19907) );
  INV_X1 U22882 ( .A(n19907), .ZN(P2_U3611) );
  OAI21_X1 U22883 ( .B1(n20674), .B2(P1_STATE_REG_2__SCAN_IN), .A(
        P1_STATE_REG_0__SCAN_IN), .ZN(n19916) );
  NOR2_X1 U22884 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20674), .ZN(n20771) );
  INV_X2 U22885 ( .A(n20771), .ZN(n20732) );
  OAI21_X1 U22886 ( .B1(n19916), .B2(P1_ADS_N_REG_SCAN_IN), .A(n20732), .ZN(
        n19908) );
  INV_X1 U22887 ( .A(n19908), .ZN(P1_U2802) );
  NAND2_X1 U22888 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n19909), .ZN(n19914) );
  INV_X1 U22889 ( .A(n19910), .ZN(n19912) );
  OAI21_X1 U22890 ( .B1(n19912), .B2(n19911), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19913) );
  OAI21_X1 U22891 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n19914), .A(n19913), 
        .ZN(P1_U2803) );
  NOR2_X1 U22892 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19917) );
  OAI21_X1 U22893 ( .B1(n19917), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20732), .ZN(
        n19915) );
  OAI21_X1 U22894 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20732), .A(n19915), 
        .ZN(P1_U2804) );
  NAND2_X1 U22895 ( .A1(n20732), .A2(n19916), .ZN(n20672) );
  INV_X1 U22896 ( .A(n20672), .ZN(n20743) );
  OAI21_X1 U22897 ( .B1(BS16), .B2(n19917), .A(n20743), .ZN(n20741) );
  OAI21_X1 U22898 ( .B1(n20743), .B2(n20761), .A(n20741), .ZN(P1_U2805) );
  OAI21_X1 U22899 ( .B1(n19920), .B2(n19919), .A(n19918), .ZN(P1_U2806) );
  NOR4_X1 U22900 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_19__SCAN_IN), .A3(P1_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_21__SCAN_IN), .ZN(n19924) );
  NOR4_X1 U22901 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_15__SCAN_IN), .A3(P1_DATAWIDTH_REG_16__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_17__SCAN_IN), .ZN(n19923) );
  NOR4_X1 U22902 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_28__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19922) );
  NOR4_X1 U22903 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_23__SCAN_IN), .A3(P1_DATAWIDTH_REG_24__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_25__SCAN_IN), .ZN(n19921) );
  NAND4_X1 U22904 ( .A1(n19924), .A2(n19923), .A3(n19922), .A4(n19921), .ZN(
        n19930) );
  NOR4_X1 U22905 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_2__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_3__SCAN_IN), .ZN(n19928) );
  AOI211_X1 U22906 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_9__SCAN_IN), .B(
        P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n19927) );
  NOR4_X1 U22907 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_10__SCAN_IN), .A3(P1_DATAWIDTH_REG_11__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_12__SCAN_IN), .ZN(n19926) );
  NOR4_X1 U22908 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_5__SCAN_IN), .A3(P1_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_7__SCAN_IN), .ZN(n19925) );
  NAND4_X1 U22909 ( .A1(n19928), .A2(n19927), .A3(n19926), .A4(n19925), .ZN(
        n19929) );
  NOR2_X1 U22910 ( .A1(n19930), .A2(n19929), .ZN(n20757) );
  INV_X1 U22911 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19932) );
  NOR3_X1 U22912 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19933) );
  OAI21_X1 U22913 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19933), .A(n20757), .ZN(
        n19931) );
  OAI21_X1 U22914 ( .B1(n20757), .B2(n19932), .A(n19931), .ZN(P1_U2807) );
  INV_X1 U22915 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20742) );
  AOI21_X1 U22916 ( .B1(n20750), .B2(n20742), .A(n19933), .ZN(n19935) );
  INV_X1 U22917 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19934) );
  INV_X1 U22918 ( .A(n20757), .ZN(n20752) );
  AOI22_X1 U22919 ( .A1(n20757), .A2(n19935), .B1(n19934), .B2(n20752), .ZN(
        P1_U2808) );
  NAND2_X1 U22920 ( .A1(n19937), .A2(n19936), .ZN(n19959) );
  AOI22_X1 U22921 ( .A1(n19938), .A2(n20034), .B1(n20026), .B2(
        P1_EBX_REG_9__SCAN_IN), .ZN(n19939) );
  OAI211_X1 U22922 ( .C1(n20031), .C2(n19940), .A(n19939), .B(n19974), .ZN(
        n19945) );
  OAI22_X1 U22923 ( .A1(n19943), .A2(n19942), .B1(P1_REIP_REG_9__SCAN_IN), 
        .B2(n19941), .ZN(n19944) );
  AOI211_X1 U22924 ( .C1(n19946), .C2(n20014), .A(n19945), .B(n19944), .ZN(
        n19947) );
  OAI21_X1 U22925 ( .B1(n19948), .B2(n19959), .A(n19947), .ZN(P1_U2831) );
  NOR2_X1 U22926 ( .A1(n20017), .A2(n19949), .ZN(n19950) );
  NOR2_X1 U22927 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n19950), .ZN(n19960) );
  AOI22_X1 U22928 ( .A1(n20026), .A2(P1_EBX_REG_8__SCAN_IN), .B1(n20014), .B2(
        n19951), .ZN(n19958) );
  NOR2_X1 U22929 ( .A1(n19952), .A2(n20008), .ZN(n19955) );
  OAI21_X1 U22930 ( .B1(n20031), .B2(n19953), .A(n19974), .ZN(n19954) );
  AOI211_X1 U22931 ( .C1(n19956), .C2(n19978), .A(n19955), .B(n19954), .ZN(
        n19957) );
  OAI211_X1 U22932 ( .C1(n19960), .C2(n19959), .A(n19958), .B(n19957), .ZN(
        P1_U2832) );
  AOI22_X1 U22933 ( .A1(n19961), .A2(n20034), .B1(n20026), .B2(
        P1_EBX_REG_7__SCAN_IN), .ZN(n19970) );
  NOR2_X1 U22934 ( .A1(P1_REIP_REG_7__SCAN_IN), .A2(n20017), .ZN(n19965) );
  INV_X1 U22935 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n19963) );
  OAI22_X1 U22936 ( .A1(n19963), .A2(n20031), .B1(n19962), .B2(n20042), .ZN(
        n19964) );
  AOI21_X1 U22937 ( .B1(n19965), .B2(n19966), .A(n19964), .ZN(n19969) );
  OAI21_X1 U22938 ( .B1(n20017), .B2(n19966), .A(n20029), .ZN(n19981) );
  AOI22_X1 U22939 ( .A1(n19967), .A2(n19978), .B1(P1_REIP_REG_7__SCAN_IN), 
        .B2(n19981), .ZN(n19968) );
  NAND4_X1 U22940 ( .A1(n19970), .A2(n19969), .A3(n19968), .A4(n19974), .ZN(
        P1_U2833) );
  INV_X1 U22941 ( .A(n19971), .ZN(n19972) );
  AOI22_X1 U22942 ( .A1(n20026), .A2(P1_EBX_REG_6__SCAN_IN), .B1(n19972), .B2(
        n20014), .ZN(n19984) );
  NAND2_X1 U22943 ( .A1(n19973), .A2(n20034), .ZN(n19975) );
  OAI211_X1 U22944 ( .C1(n20031), .C2(n19976), .A(n19975), .B(n19974), .ZN(
        n19977) );
  AOI21_X1 U22945 ( .B1(n19979), .B2(n19978), .A(n19977), .ZN(n19983) );
  AOI211_X1 U22946 ( .C1(n20019), .C2(n20004), .A(n20003), .B(n19980), .ZN(
        n19997) );
  OAI21_X1 U22947 ( .B1(P1_REIP_REG_6__SCAN_IN), .B2(n19997), .A(n19981), .ZN(
        n19982) );
  NAND3_X1 U22948 ( .A1(n19984), .A2(n19983), .A3(n19982), .ZN(P1_U2834) );
  INV_X1 U22949 ( .A(n20004), .ZN(n19985) );
  AOI21_X1 U22950 ( .B1(n20019), .B2(n19985), .A(P1_REIP_REG_5__SCAN_IN), .ZN(
        n19996) );
  INV_X1 U22951 ( .A(n19986), .ZN(n19987) );
  AOI22_X1 U22952 ( .A1(n19988), .A2(n20034), .B1(n19987), .B2(n20014), .ZN(
        n19995) );
  AOI21_X1 U22953 ( .B1(n20013), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n20001), .ZN(n19989) );
  OAI21_X1 U22954 ( .B1(n19991), .B2(n19990), .A(n19989), .ZN(n19992) );
  AOI21_X1 U22955 ( .B1(n19993), .B2(n20038), .A(n19992), .ZN(n19994) );
  OAI211_X1 U22956 ( .C1(n19997), .C2(n19996), .A(n19995), .B(n19994), .ZN(
        P1_U2835) );
  INV_X1 U22957 ( .A(n19998), .ZN(n20002) );
  NAND3_X1 U22958 ( .A1(P1_REIP_REG_3__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n19999) );
  NOR3_X1 U22959 ( .A1(n20017), .A2(P1_REIP_REG_4__SCAN_IN), .A3(n19999), .ZN(
        n20000) );
  AOI211_X1 U22960 ( .C1(n20002), .C2(n20028), .A(n20001), .B(n20000), .ZN(
        n20012) );
  AOI21_X1 U22961 ( .B1(n20019), .B2(n20004), .A(n20003), .ZN(n20005) );
  INV_X1 U22962 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20691) );
  NOR2_X1 U22963 ( .A1(n20005), .A2(n20691), .ZN(n20010) );
  INV_X1 U22964 ( .A(n20111), .ZN(n20006) );
  AOI22_X1 U22965 ( .A1(n20026), .A2(P1_EBX_REG_4__SCAN_IN), .B1(n20006), .B2(
        n20014), .ZN(n20007) );
  OAI21_X1 U22966 ( .B1(n20008), .B2(n20136), .A(n20007), .ZN(n20009) );
  AOI211_X1 U22967 ( .C1(n20108), .C2(n20038), .A(n20010), .B(n20009), .ZN(
        n20011) );
  OAI211_X1 U22968 ( .C1(n12031), .C2(n20031), .A(n20012), .B(n20011), .ZN(
        P1_U2836) );
  AOI222_X1 U22969 ( .A1(n20371), .A2(n20028), .B1(n20034), .B2(n20145), .C1(
        n20013), .C2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n20023) );
  INV_X1 U22970 ( .A(n20119), .ZN(n20015) );
  AOI22_X1 U22971 ( .A1(n20026), .A2(P1_EBX_REG_3__SCAN_IN), .B1(n20015), .B2(
        n20014), .ZN(n20022) );
  AND2_X1 U22972 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(P1_REIP_REG_1__SCAN_IN), 
        .ZN(n20016) );
  OAI21_X1 U22973 ( .B1(n20017), .B2(n20016), .A(n20029), .ZN(n20018) );
  AOI22_X1 U22974 ( .A1(n20116), .A2(n20038), .B1(P1_REIP_REG_3__SCAN_IN), 
        .B2(n20018), .ZN(n20021) );
  INV_X1 U22975 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20693) );
  NAND4_X1 U22976 ( .A1(n20019), .A2(P1_REIP_REG_1__SCAN_IN), .A3(
        P1_REIP_REG_2__SCAN_IN), .A4(n20693), .ZN(n20020) );
  NAND4_X1 U22977 ( .A1(n20023), .A2(n20022), .A3(n20021), .A4(n20020), .ZN(
        P1_U2837) );
  INV_X1 U22978 ( .A(n20024), .ZN(n20025) );
  AOI21_X1 U22979 ( .B1(n20026), .B2(P1_EBX_REG_1__SCAN_IN), .A(n20025), .ZN(
        n20041) );
  INV_X1 U22980 ( .A(n20027), .ZN(n20039) );
  INV_X1 U22981 ( .A(n20028), .ZN(n20036) );
  OAI22_X1 U22982 ( .A1(n20031), .A2(n20030), .B1(n20750), .B2(n20029), .ZN(
        n20032) );
  AOI21_X1 U22983 ( .B1(n20034), .B2(n20033), .A(n20032), .ZN(n20035) );
  OAI21_X1 U22984 ( .B1(n20372), .B2(n20036), .A(n20035), .ZN(n20037) );
  AOI21_X1 U22985 ( .B1(n20039), .B2(n20038), .A(n20037), .ZN(n20040) );
  OAI211_X1 U22986 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n20042), .A(
        n20041), .B(n20040), .ZN(P1_U2839) );
  AOI22_X1 U22987 ( .A1(P1_LWORD_REG_15__SCAN_IN), .A2(n20768), .B1(n20064), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n20044) );
  OAI21_X1 U22988 ( .B1(n12986), .B2(n20067), .A(n20044), .ZN(P1_U2921) );
  AOI22_X1 U22989 ( .A1(P1_LWORD_REG_14__SCAN_IN), .A2(n20768), .B1(n20064), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n20045) );
  OAI21_X1 U22990 ( .B1(n13832), .B2(n20067), .A(n20045), .ZN(P1_U2922) );
  AOI22_X1 U22991 ( .A1(P1_LWORD_REG_13__SCAN_IN), .A2(n20768), .B1(n20064), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n20046) );
  OAI21_X1 U22992 ( .B1(n14474), .B2(n20067), .A(n20046), .ZN(P1_U2923) );
  AOI22_X1 U22993 ( .A1(P1_LWORD_REG_12__SCAN_IN), .A2(n20768), .B1(n20064), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n20047) );
  OAI21_X1 U22994 ( .B1(n13801), .B2(n20067), .A(n20047), .ZN(P1_U2924) );
  AOI22_X1 U22995 ( .A1(P1_LWORD_REG_11__SCAN_IN), .A2(n20768), .B1(n20064), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n20048) );
  OAI21_X1 U22996 ( .B1(n20049), .B2(n20067), .A(n20048), .ZN(P1_U2925) );
  AOI22_X1 U22997 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(n20768), .B1(n20064), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n20050) );
  OAI21_X1 U22998 ( .B1(n13665), .B2(n20067), .A(n20050), .ZN(P1_U2926) );
  AOI22_X1 U22999 ( .A1(P1_LWORD_REG_9__SCAN_IN), .A2(n20768), .B1(n20064), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n20051) );
  OAI21_X1 U23000 ( .B1(n13624), .B2(n20067), .A(n20051), .ZN(P1_U2927) );
  AOI22_X1 U23001 ( .A1(P1_LWORD_REG_8__SCAN_IN), .A2(n20768), .B1(n20064), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n20052) );
  OAI21_X1 U23002 ( .B1(n20802), .B2(n20067), .A(n20052), .ZN(P1_U2928) );
  AOI22_X1 U23003 ( .A1(P1_LWORD_REG_7__SCAN_IN), .A2(n20065), .B1(n20064), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n20053) );
  OAI21_X1 U23004 ( .B1(n12085), .B2(n20067), .A(n20053), .ZN(P1_U2929) );
  AOI22_X1 U23005 ( .A1(P1_LWORD_REG_6__SCAN_IN), .A2(n20065), .B1(n20064), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n20054) );
  OAI21_X1 U23006 ( .B1(n13377), .B2(n20067), .A(n20054), .ZN(P1_U2930) );
  AOI22_X1 U23007 ( .A1(P1_LWORD_REG_5__SCAN_IN), .A2(n20065), .B1(n20064), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n20055) );
  OAI21_X1 U23008 ( .B1(n12055), .B2(n20067), .A(n20055), .ZN(P1_U2931) );
  AOI22_X1 U23009 ( .A1(P1_LWORD_REG_4__SCAN_IN), .A2(n20065), .B1(n20064), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n20056) );
  OAI21_X1 U23010 ( .B1(n20057), .B2(n20067), .A(n20056), .ZN(P1_U2932) );
  AOI22_X1 U23011 ( .A1(P1_LWORD_REG_3__SCAN_IN), .A2(n20065), .B1(n20064), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n20058) );
  OAI21_X1 U23012 ( .B1(n20059), .B2(n20067), .A(n20058), .ZN(P1_U2933) );
  AOI22_X1 U23013 ( .A1(P1_LWORD_REG_2__SCAN_IN), .A2(n20065), .B1(n20064), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n20060) );
  OAI21_X1 U23014 ( .B1(n20061), .B2(n20067), .A(n20060), .ZN(P1_U2934) );
  AOI22_X1 U23015 ( .A1(P1_LWORD_REG_1__SCAN_IN), .A2(n20065), .B1(n20064), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n20062) );
  OAI21_X1 U23016 ( .B1(n20063), .B2(n20067), .A(n20062), .ZN(P1_U2935) );
  AOI22_X1 U23017 ( .A1(P1_LWORD_REG_0__SCAN_IN), .A2(n20065), .B1(n20064), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n20066) );
  OAI21_X1 U23018 ( .B1(n20068), .B2(n20067), .A(n20066), .ZN(P1_U2936) );
  AOI22_X1 U23019 ( .A1(n20101), .A2(P1_EAX_REG_24__SCAN_IN), .B1(
        P1_UWORD_REG_8__SCAN_IN), .B2(n20075), .ZN(n20071) );
  INV_X1 U23020 ( .A(n20069), .ZN(n20070) );
  NAND2_X1 U23021 ( .A1(n20088), .A2(n20070), .ZN(n20090) );
  NAND2_X1 U23022 ( .A1(n20071), .A2(n20090), .ZN(P1_U2945) );
  AOI22_X1 U23023 ( .A1(n20101), .A2(P1_EAX_REG_25__SCAN_IN), .B1(
        P1_UWORD_REG_9__SCAN_IN), .B2(n20075), .ZN(n20074) );
  INV_X1 U23024 ( .A(n20072), .ZN(n20073) );
  NAND2_X1 U23025 ( .A1(n20088), .A2(n20073), .ZN(n20092) );
  NAND2_X1 U23026 ( .A1(n20074), .A2(n20092), .ZN(P1_U2946) );
  AOI22_X1 U23027 ( .A1(n20076), .A2(P1_EAX_REG_26__SCAN_IN), .B1(
        P1_UWORD_REG_10__SCAN_IN), .B2(n20075), .ZN(n20079) );
  INV_X1 U23028 ( .A(n20077), .ZN(n20078) );
  NAND2_X1 U23029 ( .A1(n20088), .A2(n20078), .ZN(n20094) );
  NAND2_X1 U23030 ( .A1(n20079), .A2(n20094), .ZN(P1_U2947) );
  AOI22_X1 U23031 ( .A1(n20101), .A2(P1_EAX_REG_28__SCAN_IN), .B1(
        P1_UWORD_REG_12__SCAN_IN), .B2(n20100), .ZN(n20082) );
  INV_X1 U23032 ( .A(n20080), .ZN(n20081) );
  NAND2_X1 U23033 ( .A1(n20088), .A2(n20081), .ZN(n20096) );
  NAND2_X1 U23034 ( .A1(n20082), .A2(n20096), .ZN(P1_U2949) );
  AOI22_X1 U23035 ( .A1(n20101), .A2(P1_EAX_REG_29__SCAN_IN), .B1(
        P1_UWORD_REG_13__SCAN_IN), .B2(n20100), .ZN(n20085) );
  INV_X1 U23036 ( .A(n20083), .ZN(n20084) );
  NAND2_X1 U23037 ( .A1(n20088), .A2(n20084), .ZN(n20098) );
  NAND2_X1 U23038 ( .A1(n20085), .A2(n20098), .ZN(P1_U2950) );
  AOI22_X1 U23039 ( .A1(n20101), .A2(P1_EAX_REG_30__SCAN_IN), .B1(
        P1_UWORD_REG_14__SCAN_IN), .B2(n20100), .ZN(n20089) );
  INV_X1 U23040 ( .A(n20086), .ZN(n20087) );
  NAND2_X1 U23041 ( .A1(n20088), .A2(n20087), .ZN(n20102) );
  NAND2_X1 U23042 ( .A1(n20089), .A2(n20102), .ZN(P1_U2951) );
  AOI22_X1 U23043 ( .A1(n20101), .A2(P1_EAX_REG_8__SCAN_IN), .B1(
        P1_LWORD_REG_8__SCAN_IN), .B2(n20075), .ZN(n20091) );
  NAND2_X1 U23044 ( .A1(n20091), .A2(n20090), .ZN(P1_U2960) );
  AOI22_X1 U23045 ( .A1(n20101), .A2(P1_EAX_REG_9__SCAN_IN), .B1(
        P1_LWORD_REG_9__SCAN_IN), .B2(n20100), .ZN(n20093) );
  NAND2_X1 U23046 ( .A1(n20093), .A2(n20092), .ZN(P1_U2961) );
  AOI22_X1 U23047 ( .A1(n20101), .A2(P1_EAX_REG_10__SCAN_IN), .B1(
        P1_LWORD_REG_10__SCAN_IN), .B2(n20075), .ZN(n20095) );
  NAND2_X1 U23048 ( .A1(n20095), .A2(n20094), .ZN(P1_U2962) );
  AOI22_X1 U23049 ( .A1(n20101), .A2(P1_EAX_REG_12__SCAN_IN), .B1(
        P1_LWORD_REG_12__SCAN_IN), .B2(n20100), .ZN(n20097) );
  NAND2_X1 U23050 ( .A1(n20097), .A2(n20096), .ZN(P1_U2964) );
  AOI22_X1 U23051 ( .A1(n20101), .A2(P1_EAX_REG_13__SCAN_IN), .B1(
        P1_LWORD_REG_13__SCAN_IN), .B2(n20075), .ZN(n20099) );
  NAND2_X1 U23052 ( .A1(n20099), .A2(n20098), .ZN(P1_U2965) );
  AOI22_X1 U23053 ( .A1(n20101), .A2(P1_EAX_REG_14__SCAN_IN), .B1(
        P1_LWORD_REG_14__SCAN_IN), .B2(n20100), .ZN(n20103) );
  NAND2_X1 U23054 ( .A1(n20103), .A2(n20102), .ZN(P1_U2966) );
  AOI22_X1 U23055 ( .A1(n20120), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        n20162), .B2(P1_REIP_REG_4__SCAN_IN), .ZN(n20110) );
  OAI21_X1 U23056 ( .B1(n20106), .B2(n20105), .A(n20104), .ZN(n20107) );
  INV_X1 U23057 ( .A(n20107), .ZN(n20142) );
  AOI22_X1 U23058 ( .A1(n20142), .A2(n12697), .B1(n20125), .B2(n20108), .ZN(
        n20109) );
  OAI211_X1 U23059 ( .C1(n20130), .C2(n20111), .A(n20110), .B(n20109), .ZN(
        P1_U2995) );
  AOI22_X1 U23060 ( .A1(n20120), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B1(
        n20162), .B2(P1_REIP_REG_3__SCAN_IN), .ZN(n20118) );
  OAI21_X1 U23061 ( .B1(n20114), .B2(n20113), .A(n20112), .ZN(n20115) );
  INV_X1 U23062 ( .A(n20115), .ZN(n20147) );
  AOI22_X1 U23063 ( .A1(n20147), .A2(n12697), .B1(n20125), .B2(n20116), .ZN(
        n20117) );
  OAI211_X1 U23064 ( .C1(n20130), .C2(n20119), .A(n20118), .B(n20117), .ZN(
        P1_U2996) );
  AOI22_X1 U23065 ( .A1(n20120), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B1(
        n20162), .B2(P1_REIP_REG_2__SCAN_IN), .ZN(n20128) );
  OAI21_X1 U23066 ( .B1(n20123), .B2(n20122), .A(n20121), .ZN(n20124) );
  INV_X1 U23067 ( .A(n20124), .ZN(n20161) );
  AOI22_X1 U23068 ( .A1(n20126), .A2(n20125), .B1(n20161), .B2(n12697), .ZN(
        n20127) );
  OAI211_X1 U23069 ( .C1(n20130), .C2(n20129), .A(n20128), .B(n20127), .ZN(
        P1_U2997) );
  NOR2_X1 U23070 ( .A1(n20154), .A2(n20131), .ZN(n20156) );
  INV_X1 U23071 ( .A(n20132), .ZN(n20133) );
  OAI21_X1 U23072 ( .B1(n20164), .B2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        n20133), .ZN(n20159) );
  AOI211_X1 U23073 ( .C1(n20152), .C2(n20134), .A(n20156), .B(n20159), .ZN(
        n20151) );
  OAI22_X1 U23074 ( .A1(n20137), .A2(n20136), .B1(n20691), .B2(n20135), .ZN(
        n20141) );
  AOI211_X1 U23075 ( .C1(n20144), .C2(n20150), .A(n20139), .B(n20138), .ZN(
        n20140) );
  AOI211_X1 U23076 ( .C1(n20142), .C2(n20160), .A(n20141), .B(n20140), .ZN(
        n20143) );
  OAI21_X1 U23077 ( .B1(n20151), .B2(n20144), .A(n20143), .ZN(P1_U3027) );
  AOI22_X1 U23078 ( .A1(n20157), .A2(n20145), .B1(n20162), .B2(
        P1_REIP_REG_3__SCAN_IN), .ZN(n20149) );
  AOI22_X1 U23079 ( .A1(n20147), .A2(n20160), .B1(n20150), .B2(n20146), .ZN(
        n20148) );
  OAI211_X1 U23080 ( .C1(n20151), .C2(n20150), .A(n20149), .B(n20148), .ZN(
        P1_U3028) );
  NOR4_X1 U23081 ( .A1(n20154), .A2(n20153), .A3(n20152), .A4(n20165), .ZN(
        n20155) );
  AOI211_X1 U23082 ( .C1(n20158), .C2(n20157), .A(n20156), .B(n20155), .ZN(
        n20169) );
  AOI22_X1 U23083 ( .A1(n20161), .A2(n20160), .B1(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20159), .ZN(n20168) );
  NAND2_X1 U23084 ( .A1(n20162), .A2(P1_REIP_REG_2__SCAN_IN), .ZN(n20167) );
  OR4_X1 U23085 ( .A1(n20165), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A3(
        n20164), .A4(n20163), .ZN(n20166) );
  NAND4_X1 U23086 ( .A1(n20169), .A2(n20168), .A3(n20167), .A4(n20166), .ZN(
        P1_U3029) );
  NOR2_X1 U23087 ( .A1(n12545), .A2(n20170), .ZN(P1_U3032) );
  INV_X1 U23088 ( .A(n20275), .ZN(n20173) );
  NOR3_X1 U23089 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20215) );
  NAND2_X1 U23090 ( .A1(n20553), .A2(n20215), .ZN(n20203) );
  OAI22_X1 U23091 ( .A1(n20204), .A2(n20515), .B1(n20203), .B2(n20503), .ZN(
        n20174) );
  INV_X1 U23092 ( .A(n20174), .ZN(n20184) );
  INV_X1 U23093 ( .A(n20235), .ZN(n20175) );
  OAI21_X1 U23094 ( .B1(n20175), .B2(n20663), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20176) );
  NAND2_X1 U23095 ( .A1(n20176), .A2(n20585), .ZN(n20182) );
  OR2_X1 U23096 ( .A1(n20371), .A2(n20177), .ZN(n20277) );
  INV_X1 U23097 ( .A(n20372), .ZN(n20594) );
  NOR2_X1 U23098 ( .A1(n20277), .A2(n20594), .ZN(n20180) );
  NAND2_X1 U23099 ( .A1(n20435), .A2(n20373), .ZN(n20314) );
  AOI22_X1 U23100 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20314), .B1(
        P1_STATE2_REG_3__SCAN_IN), .B2(n20203), .ZN(n20179) );
  OAI211_X1 U23101 ( .C1(n20182), .C2(n20180), .A(n20433), .B(n20179), .ZN(
        n20207) );
  INV_X1 U23102 ( .A(n20180), .ZN(n20181) );
  OAI22_X1 U23103 ( .A1(n20182), .A2(n20181), .B1(n20436), .B2(n20314), .ZN(
        n20206) );
  AOI22_X1 U23104 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20207), .B1(
        n20592), .B2(n20206), .ZN(n20183) );
  OAI211_X1 U23105 ( .C1(n20604), .C2(n20235), .A(n20184), .B(n20183), .ZN(
        P1_U3033) );
  OAI22_X1 U23106 ( .A1(n20204), .A2(n20520), .B1(n20203), .B2(n20516), .ZN(
        n20185) );
  INV_X1 U23107 ( .A(n20185), .ZN(n20187) );
  AOI22_X1 U23108 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20207), .B1(
        n20606), .B2(n20206), .ZN(n20186) );
  OAI211_X1 U23109 ( .C1(n20610), .C2(n20235), .A(n20187), .B(n20186), .ZN(
        P1_U3034) );
  OAI22_X1 U23110 ( .A1(n20204), .A2(n20651), .B1(n20203), .B2(n20521), .ZN(
        n20188) );
  INV_X1 U23111 ( .A(n20188), .ZN(n20190) );
  AOI22_X1 U23112 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20207), .B1(
        n20647), .B2(n20206), .ZN(n20189) );
  OAI211_X1 U23113 ( .C1(n20614), .C2(n20235), .A(n20190), .B(n20189), .ZN(
        P1_U3035) );
  OAI22_X1 U23114 ( .A1(n20204), .A2(n20529), .B1(n20203), .B2(n20525), .ZN(
        n20191) );
  INV_X1 U23115 ( .A(n20191), .ZN(n20193) );
  AOI22_X1 U23116 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20207), .B1(
        n20616), .B2(n20206), .ZN(n20192) );
  OAI211_X1 U23117 ( .C1(n20620), .C2(n20235), .A(n20193), .B(n20192), .ZN(
        P1_U3036) );
  OAI22_X1 U23118 ( .A1(n20204), .A2(n20657), .B1(n20203), .B2(n20530), .ZN(
        n20194) );
  INV_X1 U23119 ( .A(n20194), .ZN(n20196) );
  AOI22_X1 U23120 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20207), .B1(
        n20653), .B2(n20206), .ZN(n20195) );
  OAI211_X1 U23121 ( .C1(n20624), .C2(n20235), .A(n20196), .B(n20195), .ZN(
        P1_U3037) );
  OAI22_X1 U23122 ( .A1(n20204), .A2(n20538), .B1(n20203), .B2(n20534), .ZN(
        n20197) );
  INV_X1 U23123 ( .A(n20197), .ZN(n20199) );
  AOI22_X1 U23124 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20207), .B1(
        n20626), .B2(n20206), .ZN(n20198) );
  OAI211_X1 U23125 ( .C1(n20630), .C2(n20235), .A(n20199), .B(n20198), .ZN(
        P1_U3038) );
  OAI22_X1 U23126 ( .A1(n20204), .A2(n20543), .B1(n20203), .B2(n20539), .ZN(
        n20200) );
  INV_X1 U23127 ( .A(n20200), .ZN(n20202) );
  AOI22_X1 U23128 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20207), .B1(
        n20632), .B2(n20206), .ZN(n20201) );
  OAI211_X1 U23129 ( .C1(n20636), .C2(n20235), .A(n20202), .B(n20201), .ZN(
        P1_U3039) );
  OAI22_X1 U23130 ( .A1(n20204), .A2(n20668), .B1(n20203), .B2(n20545), .ZN(
        n20205) );
  INV_X1 U23131 ( .A(n20205), .ZN(n20209) );
  AOI22_X1 U23132 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20207), .B1(
        n20661), .B2(n20206), .ZN(n20208) );
  OAI211_X1 U23133 ( .C1(n20644), .C2(n20235), .A(n20209), .B(n20208), .ZN(
        P1_U3040) );
  OR2_X1 U23134 ( .A1(n20277), .A2(n20340), .ZN(n20211) );
  INV_X1 U23135 ( .A(n20215), .ZN(n20212) );
  NOR2_X1 U23136 ( .A1(n20553), .A2(n20212), .ZN(n20230) );
  INV_X1 U23137 ( .A(n20230), .ZN(n20210) );
  AND2_X1 U23138 ( .A1(n20211), .A2(n20210), .ZN(n20213) );
  OAI22_X1 U23139 ( .A1(n20213), .A2(n20556), .B1(n20212), .B2(n20760), .ZN(
        n20231) );
  AOI22_X1 U23140 ( .A1(n20592), .A2(n20231), .B1(n20591), .B2(n20230), .ZN(
        n20217) );
  OAI21_X1 U23141 ( .B1(n20275), .B2(n20761), .A(n20213), .ZN(n20214) );
  OAI221_X1 U23142 ( .B1(n20585), .B2(n20215), .C1(n20556), .C2(n20214), .A(
        n20561), .ZN(n20232) );
  AOI22_X1 U23143 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20232), .B1(
        n20237), .B2(n20404), .ZN(n20216) );
  OAI211_X1 U23144 ( .C1(n20515), .C2(n20235), .A(n20217), .B(n20216), .ZN(
        P1_U3041) );
  AOI22_X1 U23145 ( .A1(n20606), .A2(n20231), .B1(n20605), .B2(n20230), .ZN(
        n20219) );
  AOI22_X1 U23146 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20232), .B1(
        n20237), .B2(n20479), .ZN(n20218) );
  OAI211_X1 U23147 ( .C1(n20520), .C2(n20235), .A(n20219), .B(n20218), .ZN(
        P1_U3042) );
  AOI22_X1 U23148 ( .A1(n20647), .A2(n20231), .B1(n20646), .B2(n20230), .ZN(
        n20221) );
  AOI22_X1 U23149 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20232), .B1(
        n20237), .B2(n20648), .ZN(n20220) );
  OAI211_X1 U23150 ( .C1(n20651), .C2(n20235), .A(n20221), .B(n20220), .ZN(
        P1_U3043) );
  AOI22_X1 U23151 ( .A1(n20616), .A2(n20231), .B1(n20615), .B2(n20230), .ZN(
        n20223) );
  AOI22_X1 U23152 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20232), .B1(
        n20237), .B2(n20411), .ZN(n20222) );
  OAI211_X1 U23153 ( .C1(n20529), .C2(n20235), .A(n20223), .B(n20222), .ZN(
        P1_U3044) );
  AOI22_X1 U23154 ( .A1(n20653), .A2(n20231), .B1(n20652), .B2(n20230), .ZN(
        n20225) );
  AOI22_X1 U23155 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20232), .B1(
        n20237), .B2(n20654), .ZN(n20224) );
  OAI211_X1 U23156 ( .C1(n20657), .C2(n20235), .A(n20225), .B(n20224), .ZN(
        P1_U3045) );
  AOI22_X1 U23157 ( .A1(n20626), .A2(n20231), .B1(n20625), .B2(n20230), .ZN(
        n20227) );
  AOI22_X1 U23158 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20232), .B1(
        n20237), .B2(n20416), .ZN(n20226) );
  OAI211_X1 U23159 ( .C1(n20538), .C2(n20235), .A(n20227), .B(n20226), .ZN(
        P1_U3046) );
  AOI22_X1 U23160 ( .A1(n20632), .A2(n20231), .B1(n20631), .B2(n20230), .ZN(
        n20229) );
  AOI22_X1 U23161 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20232), .B1(
        n20237), .B2(n20419), .ZN(n20228) );
  OAI211_X1 U23162 ( .C1(n20543), .C2(n20235), .A(n20229), .B(n20228), .ZN(
        P1_U3047) );
  AOI22_X1 U23163 ( .A1(n20661), .A2(n20231), .B1(n20658), .B2(n20230), .ZN(
        n20234) );
  AOI22_X1 U23164 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20232), .B1(
        n20237), .B2(n20662), .ZN(n20233) );
  OAI211_X1 U23165 ( .C1(n20668), .C2(n20235), .A(n20234), .B(n20233), .ZN(
        P1_U3048) );
  NAND3_X1 U23166 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n20501), .A3(
        n20502), .ZN(n20281) );
  OR2_X1 U23167 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20281), .ZN(
        n20266) );
  OAI22_X1 U23168 ( .A1(n20267), .A2(n20515), .B1(n20266), .B2(n20503), .ZN(
        n20236) );
  INV_X1 U23169 ( .A(n20236), .ZN(n20247) );
  INV_X1 U23170 ( .A(n20305), .ZN(n20238) );
  OAI21_X1 U23171 ( .B1(n20238), .B2(n20237), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20239) );
  NAND2_X1 U23172 ( .A1(n20239), .A2(n20585), .ZN(n20245) );
  NOR2_X1 U23173 ( .A1(n20277), .A2(n20372), .ZN(n20242) );
  AOI21_X1 U23174 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20266), .A(n20240), 
        .ZN(n20241) );
  OAI211_X1 U23175 ( .C1(n20245), .C2(n20242), .A(n20433), .B(n20241), .ZN(
        n20270) );
  INV_X1 U23176 ( .A(n20242), .ZN(n20244) );
  OAI22_X1 U23177 ( .A1(n20245), .A2(n20244), .B1(n20243), .B2(n20436), .ZN(
        n20269) );
  AOI22_X1 U23178 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20270), .B1(
        n20592), .B2(n20269), .ZN(n20246) );
  OAI211_X1 U23179 ( .C1(n20604), .C2(n20305), .A(n20247), .B(n20246), .ZN(
        P1_U3049) );
  OAI22_X1 U23180 ( .A1(n20305), .A2(n20610), .B1(n20516), .B2(n20266), .ZN(
        n20248) );
  INV_X1 U23181 ( .A(n20248), .ZN(n20250) );
  AOI22_X1 U23182 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20270), .B1(
        n20606), .B2(n20269), .ZN(n20249) );
  OAI211_X1 U23183 ( .C1(n20520), .C2(n20267), .A(n20250), .B(n20249), .ZN(
        P1_U3050) );
  OAI22_X1 U23184 ( .A1(n20267), .A2(n20651), .B1(n20266), .B2(n20521), .ZN(
        n20251) );
  INV_X1 U23185 ( .A(n20251), .ZN(n20253) );
  AOI22_X1 U23186 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20270), .B1(
        n20647), .B2(n20269), .ZN(n20252) );
  OAI211_X1 U23187 ( .C1(n20614), .C2(n20305), .A(n20253), .B(n20252), .ZN(
        P1_U3051) );
  OAI22_X1 U23188 ( .A1(n20305), .A2(n20620), .B1(n20525), .B2(n20266), .ZN(
        n20254) );
  INV_X1 U23189 ( .A(n20254), .ZN(n20256) );
  AOI22_X1 U23190 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20270), .B1(
        n20616), .B2(n20269), .ZN(n20255) );
  OAI211_X1 U23191 ( .C1(n20529), .C2(n20267), .A(n20256), .B(n20255), .ZN(
        P1_U3052) );
  OAI22_X1 U23192 ( .A1(n20267), .A2(n20657), .B1(n20266), .B2(n20530), .ZN(
        n20257) );
  INV_X1 U23193 ( .A(n20257), .ZN(n20259) );
  AOI22_X1 U23194 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20270), .B1(
        n20653), .B2(n20269), .ZN(n20258) );
  OAI211_X1 U23195 ( .C1(n20624), .C2(n20305), .A(n20259), .B(n20258), .ZN(
        P1_U3053) );
  OAI22_X1 U23196 ( .A1(n20305), .A2(n20630), .B1(n20534), .B2(n20266), .ZN(
        n20260) );
  INV_X1 U23197 ( .A(n20260), .ZN(n20262) );
  AOI22_X1 U23198 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20270), .B1(
        n20626), .B2(n20269), .ZN(n20261) );
  OAI211_X1 U23199 ( .C1(n20538), .C2(n20267), .A(n20262), .B(n20261), .ZN(
        P1_U3054) );
  OAI22_X1 U23200 ( .A1(n20267), .A2(n20543), .B1(n20266), .B2(n20539), .ZN(
        n20263) );
  INV_X1 U23201 ( .A(n20263), .ZN(n20265) );
  AOI22_X1 U23202 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20270), .B1(
        n20632), .B2(n20269), .ZN(n20264) );
  OAI211_X1 U23203 ( .C1(n20636), .C2(n20305), .A(n20265), .B(n20264), .ZN(
        P1_U3055) );
  OAI22_X1 U23204 ( .A1(n20267), .A2(n20668), .B1(n20266), .B2(n20545), .ZN(
        n20268) );
  INV_X1 U23205 ( .A(n20268), .ZN(n20272) );
  AOI22_X1 U23206 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20270), .B1(
        n20661), .B2(n20269), .ZN(n20271) );
  OAI211_X1 U23207 ( .C1(n20644), .C2(n20305), .A(n20272), .B(n20271), .ZN(
        P1_U3056) );
  OR2_X1 U23208 ( .A1(n20468), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n20304) );
  OAI22_X1 U23209 ( .A1(n20315), .A2(n20604), .B1(n20503), .B2(n20304), .ZN(
        n20273) );
  INV_X1 U23210 ( .A(n20273), .ZN(n20285) );
  OAI21_X1 U23211 ( .B1(n20275), .B2(n20274), .A(n20585), .ZN(n20283) );
  INV_X1 U23212 ( .A(n20469), .ZN(n20276) );
  OR2_X1 U23213 ( .A1(n20277), .A2(n20276), .ZN(n20278) );
  INV_X1 U23214 ( .A(n20282), .ZN(n20280) );
  NAND2_X1 U23215 ( .A1(n20556), .A2(n20281), .ZN(n20279) );
  OAI211_X1 U23216 ( .C1(n20283), .C2(n20280), .A(n20561), .B(n20279), .ZN(
        n20308) );
  OAI22_X1 U23217 ( .A1(n20283), .A2(n20282), .B1(n20760), .B2(n20281), .ZN(
        n20307) );
  AOI22_X1 U23218 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20308), .B1(
        n20592), .B2(n20307), .ZN(n20284) );
  OAI211_X1 U23219 ( .C1(n20515), .C2(n20305), .A(n20285), .B(n20284), .ZN(
        P1_U3057) );
  OAI22_X1 U23220 ( .A1(n20305), .A2(n20520), .B1(n20304), .B2(n20516), .ZN(
        n20286) );
  INV_X1 U23221 ( .A(n20286), .ZN(n20288) );
  AOI22_X1 U23222 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20308), .B1(
        n20606), .B2(n20307), .ZN(n20287) );
  OAI211_X1 U23223 ( .C1(n20610), .C2(n20315), .A(n20288), .B(n20287), .ZN(
        P1_U3058) );
  OAI22_X1 U23224 ( .A1(n20305), .A2(n20651), .B1(n20304), .B2(n20521), .ZN(
        n20289) );
  INV_X1 U23225 ( .A(n20289), .ZN(n20291) );
  AOI22_X1 U23226 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20308), .B1(
        n20647), .B2(n20307), .ZN(n20290) );
  OAI211_X1 U23227 ( .C1(n20614), .C2(n20315), .A(n20291), .B(n20290), .ZN(
        P1_U3059) );
  OAI22_X1 U23228 ( .A1(n20315), .A2(n20620), .B1(n20525), .B2(n20304), .ZN(
        n20292) );
  INV_X1 U23229 ( .A(n20292), .ZN(n20294) );
  AOI22_X1 U23230 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20308), .B1(
        n20616), .B2(n20307), .ZN(n20293) );
  OAI211_X1 U23231 ( .C1(n20529), .C2(n20305), .A(n20294), .B(n20293), .ZN(
        P1_U3060) );
  OAI22_X1 U23232 ( .A1(n20315), .A2(n20624), .B1(n20530), .B2(n20304), .ZN(
        n20295) );
  INV_X1 U23233 ( .A(n20295), .ZN(n20297) );
  AOI22_X1 U23234 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20308), .B1(
        n20653), .B2(n20307), .ZN(n20296) );
  OAI211_X1 U23235 ( .C1(n20657), .C2(n20305), .A(n20297), .B(n20296), .ZN(
        P1_U3061) );
  OAI22_X1 U23236 ( .A1(n20305), .A2(n20538), .B1(n20304), .B2(n20534), .ZN(
        n20298) );
  INV_X1 U23237 ( .A(n20298), .ZN(n20300) );
  AOI22_X1 U23238 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20308), .B1(
        n20626), .B2(n20307), .ZN(n20299) );
  OAI211_X1 U23239 ( .C1(n20630), .C2(n20315), .A(n20300), .B(n20299), .ZN(
        P1_U3062) );
  OAI22_X1 U23240 ( .A1(n20315), .A2(n20636), .B1(n20539), .B2(n20304), .ZN(
        n20301) );
  INV_X1 U23241 ( .A(n20301), .ZN(n20303) );
  AOI22_X1 U23242 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20308), .B1(
        n20632), .B2(n20307), .ZN(n20302) );
  OAI211_X1 U23243 ( .C1(n20543), .C2(n20305), .A(n20303), .B(n20302), .ZN(
        P1_U3063) );
  OAI22_X1 U23244 ( .A1(n20305), .A2(n20668), .B1(n20304), .B2(n20545), .ZN(
        n20306) );
  INV_X1 U23245 ( .A(n20306), .ZN(n20310) );
  AOI22_X1 U23246 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20308), .B1(
        n20661), .B2(n20307), .ZN(n20309) );
  OAI211_X1 U23247 ( .C1(n20644), .C2(n20315), .A(n20310), .B(n20309), .ZN(
        P1_U3064) );
  INV_X1 U23248 ( .A(n20311), .ZN(n20312) );
  NAND3_X1 U23249 ( .A1(n20341), .A2(n20585), .A3(n20372), .ZN(n20313) );
  OAI21_X1 U23250 ( .B1(n20314), .B2(n20587), .A(n20313), .ZN(n20335) );
  NOR3_X1 U23251 ( .A1(n20502), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20348) );
  INV_X1 U23252 ( .A(n20348), .ZN(n20342) );
  NOR2_X1 U23253 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20342), .ZN(
        n20334) );
  AOI22_X1 U23254 ( .A1(n20592), .A2(n20335), .B1(n20591), .B2(n20334), .ZN(
        n20321) );
  INV_X1 U23255 ( .A(n20369), .ZN(n20316) );
  OAI21_X1 U23256 ( .B1(n20336), .B2(n20316), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20317) );
  OAI21_X1 U23257 ( .B1(n20594), .B2(n20318), .A(n20317), .ZN(n20319) );
  AOI22_X1 U23258 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20337), .B1(
        n20336), .B2(n20601), .ZN(n20320) );
  OAI211_X1 U23259 ( .C1(n20604), .C2(n20369), .A(n20321), .B(n20320), .ZN(
        P1_U3065) );
  AOI22_X1 U23260 ( .A1(n20606), .A2(n20335), .B1(n20605), .B2(n20334), .ZN(
        n20323) );
  AOI22_X1 U23261 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20337), .B1(
        n20336), .B2(n20607), .ZN(n20322) );
  OAI211_X1 U23262 ( .C1(n20610), .C2(n20369), .A(n20323), .B(n20322), .ZN(
        P1_U3066) );
  AOI22_X1 U23263 ( .A1(n20647), .A2(n20335), .B1(n20646), .B2(n20334), .ZN(
        n20325) );
  AOI22_X1 U23264 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20337), .B1(
        n20336), .B2(n20611), .ZN(n20324) );
  OAI211_X1 U23265 ( .C1(n20614), .C2(n20369), .A(n20325), .B(n20324), .ZN(
        P1_U3067) );
  AOI22_X1 U23266 ( .A1(n20616), .A2(n20335), .B1(n20615), .B2(n20334), .ZN(
        n20327) );
  AOI22_X1 U23267 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20337), .B1(
        n20336), .B2(n20617), .ZN(n20326) );
  OAI211_X1 U23268 ( .C1(n20620), .C2(n20369), .A(n20327), .B(n20326), .ZN(
        P1_U3068) );
  AOI22_X1 U23269 ( .A1(n20653), .A2(n20335), .B1(n20652), .B2(n20334), .ZN(
        n20329) );
  AOI22_X1 U23270 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20337), .B1(
        n20336), .B2(n20621), .ZN(n20328) );
  OAI211_X1 U23271 ( .C1(n20624), .C2(n20369), .A(n20329), .B(n20328), .ZN(
        P1_U3069) );
  AOI22_X1 U23272 ( .A1(n20626), .A2(n20335), .B1(n20625), .B2(n20334), .ZN(
        n20331) );
  AOI22_X1 U23273 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20337), .B1(
        n20336), .B2(n20627), .ZN(n20330) );
  OAI211_X1 U23274 ( .C1(n20630), .C2(n20369), .A(n20331), .B(n20330), .ZN(
        P1_U3070) );
  AOI22_X1 U23275 ( .A1(n20632), .A2(n20335), .B1(n20631), .B2(n20334), .ZN(
        n20333) );
  AOI22_X1 U23276 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20337), .B1(
        n20336), .B2(n20633), .ZN(n20332) );
  OAI211_X1 U23277 ( .C1(n20636), .C2(n20369), .A(n20333), .B(n20332), .ZN(
        P1_U3071) );
  AOI22_X1 U23278 ( .A1(n20661), .A2(n20335), .B1(n20658), .B2(n20334), .ZN(
        n20339) );
  AOI22_X1 U23279 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20337), .B1(
        n20336), .B2(n20639), .ZN(n20338) );
  OAI211_X1 U23280 ( .C1(n20644), .C2(n20369), .A(n20339), .B(n20338), .ZN(
        P1_U3072) );
  INV_X1 U23281 ( .A(n20340), .ZN(n20554) );
  NOR2_X1 U23282 ( .A1(n20553), .A2(n20342), .ZN(n20363) );
  AOI21_X1 U23283 ( .B1(n20341), .B2(n20554), .A(n20363), .ZN(n20344) );
  OAI22_X1 U23284 ( .A1(n20344), .A2(n20556), .B1(n20342), .B2(n20760), .ZN(
        n20364) );
  AOI22_X1 U23285 ( .A1(n20592), .A2(n20364), .B1(n20591), .B2(n20363), .ZN(
        n20350) );
  INV_X1 U23286 ( .A(n20343), .ZN(n20346) );
  OAI21_X1 U23287 ( .B1(n20346), .B2(n20345), .A(n20344), .ZN(n20347) );
  OAI211_X1 U23288 ( .C1(n20585), .C2(n20348), .A(n20561), .B(n20347), .ZN(
        n20366) );
  AOI22_X1 U23289 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20366), .B1(
        n20365), .B2(n20404), .ZN(n20349) );
  OAI211_X1 U23290 ( .C1(n20515), .C2(n20369), .A(n20350), .B(n20349), .ZN(
        P1_U3073) );
  AOI22_X1 U23291 ( .A1(n20606), .A2(n20364), .B1(n20605), .B2(n20363), .ZN(
        n20352) );
  AOI22_X1 U23292 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20366), .B1(
        n20365), .B2(n20479), .ZN(n20351) );
  OAI211_X1 U23293 ( .C1(n20520), .C2(n20369), .A(n20352), .B(n20351), .ZN(
        P1_U3074) );
  AOI22_X1 U23294 ( .A1(n20647), .A2(n20364), .B1(n20646), .B2(n20363), .ZN(
        n20354) );
  AOI22_X1 U23295 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20366), .B1(
        n20365), .B2(n20648), .ZN(n20353) );
  OAI211_X1 U23296 ( .C1(n20651), .C2(n20369), .A(n20354), .B(n20353), .ZN(
        P1_U3075) );
  AOI22_X1 U23297 ( .A1(n20616), .A2(n20364), .B1(n20615), .B2(n20363), .ZN(
        n20356) );
  AOI22_X1 U23298 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20366), .B1(
        n20365), .B2(n20411), .ZN(n20355) );
  OAI211_X1 U23299 ( .C1(n20529), .C2(n20369), .A(n20356), .B(n20355), .ZN(
        P1_U3076) );
  AOI22_X1 U23300 ( .A1(n20653), .A2(n20364), .B1(n20652), .B2(n20363), .ZN(
        n20358) );
  AOI22_X1 U23301 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20366), .B1(
        n20365), .B2(n20654), .ZN(n20357) );
  OAI211_X1 U23302 ( .C1(n20657), .C2(n20369), .A(n20358), .B(n20357), .ZN(
        P1_U3077) );
  AOI22_X1 U23303 ( .A1(n20626), .A2(n20364), .B1(n20625), .B2(n20363), .ZN(
        n20360) );
  AOI22_X1 U23304 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20366), .B1(
        n20365), .B2(n20416), .ZN(n20359) );
  OAI211_X1 U23305 ( .C1(n20538), .C2(n20369), .A(n20360), .B(n20359), .ZN(
        P1_U3078) );
  AOI22_X1 U23306 ( .A1(n20632), .A2(n20364), .B1(n20631), .B2(n20363), .ZN(
        n20362) );
  AOI22_X1 U23307 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20366), .B1(
        n20365), .B2(n20419), .ZN(n20361) );
  OAI211_X1 U23308 ( .C1(n20543), .C2(n20369), .A(n20362), .B(n20361), .ZN(
        P1_U3079) );
  AOI22_X1 U23309 ( .A1(n20661), .A2(n20364), .B1(n20658), .B2(n20363), .ZN(
        n20368) );
  AOI22_X1 U23310 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20366), .B1(
        n20365), .B2(n20662), .ZN(n20367) );
  OAI211_X1 U23311 ( .C1(n20668), .C2(n20369), .A(n20368), .B(n20367), .ZN(
        P1_U3080) );
  INV_X1 U23312 ( .A(n20467), .ZN(n20474) );
  AND2_X1 U23313 ( .A1(n13187), .A2(n20371), .ZN(n20470) );
  NOR3_X1 U23314 ( .A1(n20501), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20403) );
  INV_X1 U23315 ( .A(n20403), .ZN(n20400) );
  NOR2_X1 U23316 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20400), .ZN(
        n20394) );
  AOI21_X1 U23317 ( .B1(n20470), .B2(n20372), .A(n20394), .ZN(n20376) );
  INV_X1 U23318 ( .A(n20373), .ZN(n20374) );
  NAND2_X1 U23319 ( .A1(n20374), .A2(n20435), .ZN(n20510) );
  OAI22_X1 U23320 ( .A1(n20376), .A2(n20556), .B1(n20436), .B2(n20510), .ZN(
        n20395) );
  AOI22_X1 U23321 ( .A1(n20592), .A2(n20395), .B1(n20591), .B2(n20394), .ZN(
        n20381) );
  INV_X1 U23322 ( .A(n20428), .ZN(n20375) );
  OAI21_X1 U23323 ( .B1(n20375), .B2(n20396), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20377) );
  NAND2_X1 U23324 ( .A1(n20377), .A2(n20376), .ZN(n20378) );
  AOI22_X1 U23325 ( .A1(n20397), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n20396), .B2(n20601), .ZN(n20380) );
  OAI211_X1 U23326 ( .C1(n20604), .C2(n20428), .A(n20381), .B(n20380), .ZN(
        P1_U3097) );
  AOI22_X1 U23327 ( .A1(n20606), .A2(n20395), .B1(n20605), .B2(n20394), .ZN(
        n20383) );
  AOI22_X1 U23328 ( .A1(n20397), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n20396), .B2(n20607), .ZN(n20382) );
  OAI211_X1 U23329 ( .C1(n20610), .C2(n20428), .A(n20383), .B(n20382), .ZN(
        P1_U3098) );
  AOI22_X1 U23330 ( .A1(n20647), .A2(n20395), .B1(n20646), .B2(n20394), .ZN(
        n20385) );
  AOI22_X1 U23331 ( .A1(n20397), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n20396), .B2(n20611), .ZN(n20384) );
  OAI211_X1 U23332 ( .C1(n20614), .C2(n20428), .A(n20385), .B(n20384), .ZN(
        P1_U3099) );
  AOI22_X1 U23333 ( .A1(n20616), .A2(n20395), .B1(n20615), .B2(n20394), .ZN(
        n20387) );
  AOI22_X1 U23334 ( .A1(n20397), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n20396), .B2(n20617), .ZN(n20386) );
  OAI211_X1 U23335 ( .C1(n20620), .C2(n20428), .A(n20387), .B(n20386), .ZN(
        P1_U3100) );
  AOI22_X1 U23336 ( .A1(n20653), .A2(n20395), .B1(n20652), .B2(n20394), .ZN(
        n20389) );
  AOI22_X1 U23337 ( .A1(n20397), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n20396), .B2(n20621), .ZN(n20388) );
  OAI211_X1 U23338 ( .C1(n20624), .C2(n20428), .A(n20389), .B(n20388), .ZN(
        P1_U3101) );
  AOI22_X1 U23339 ( .A1(n20626), .A2(n20395), .B1(n20625), .B2(n20394), .ZN(
        n20391) );
  AOI22_X1 U23340 ( .A1(n20397), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n20396), .B2(n20627), .ZN(n20390) );
  OAI211_X1 U23341 ( .C1(n20630), .C2(n20428), .A(n20391), .B(n20390), .ZN(
        P1_U3102) );
  AOI22_X1 U23342 ( .A1(n20632), .A2(n20395), .B1(n20631), .B2(n20394), .ZN(
        n20393) );
  AOI22_X1 U23343 ( .A1(n20397), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n20396), .B2(n20633), .ZN(n20392) );
  OAI211_X1 U23344 ( .C1(n20636), .C2(n20428), .A(n20393), .B(n20392), .ZN(
        P1_U3103) );
  AOI22_X1 U23345 ( .A1(n20661), .A2(n20395), .B1(n20658), .B2(n20394), .ZN(
        n20399) );
  AOI22_X1 U23346 ( .A1(n20397), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n20396), .B2(n20639), .ZN(n20398) );
  OAI211_X1 U23347 ( .C1(n20644), .C2(n20428), .A(n20399), .B(n20398), .ZN(
        P1_U3104) );
  NOR2_X1 U23348 ( .A1(n20553), .A2(n20400), .ZN(n20422) );
  AOI21_X1 U23349 ( .B1(n20470), .B2(n20554), .A(n20422), .ZN(n20401) );
  OAI22_X1 U23350 ( .A1(n20401), .A2(n20556), .B1(n20400), .B2(n20760), .ZN(
        n20423) );
  AOI22_X1 U23351 ( .A1(n20592), .A2(n20423), .B1(n20591), .B2(n20422), .ZN(
        n20406) );
  OAI21_X1 U23352 ( .B1(n20467), .B2(n20761), .A(n20401), .ZN(n20402) );
  OAI221_X1 U23353 ( .B1(n20585), .B2(n20403), .C1(n20556), .C2(n20402), .A(
        n20561), .ZN(n20425) );
  AOI22_X1 U23354 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20404), .ZN(n20405) );
  OAI211_X1 U23355 ( .C1(n20515), .C2(n20428), .A(n20406), .B(n20405), .ZN(
        P1_U3105) );
  AOI22_X1 U23356 ( .A1(n20606), .A2(n20423), .B1(n20605), .B2(n20422), .ZN(
        n20408) );
  AOI22_X1 U23357 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20479), .ZN(n20407) );
  OAI211_X1 U23358 ( .C1(n20520), .C2(n20428), .A(n20408), .B(n20407), .ZN(
        P1_U3106) );
  AOI22_X1 U23359 ( .A1(n20647), .A2(n20423), .B1(n20646), .B2(n20422), .ZN(
        n20410) );
  AOI22_X1 U23360 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20648), .ZN(n20409) );
  OAI211_X1 U23361 ( .C1(n20651), .C2(n20428), .A(n20410), .B(n20409), .ZN(
        P1_U3107) );
  AOI22_X1 U23362 ( .A1(n20616), .A2(n20423), .B1(n20615), .B2(n20422), .ZN(
        n20413) );
  AOI22_X1 U23363 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20411), .ZN(n20412) );
  OAI211_X1 U23364 ( .C1(n20529), .C2(n20428), .A(n20413), .B(n20412), .ZN(
        P1_U3108) );
  AOI22_X1 U23365 ( .A1(n20653), .A2(n20423), .B1(n20652), .B2(n20422), .ZN(
        n20415) );
  AOI22_X1 U23366 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20654), .ZN(n20414) );
  OAI211_X1 U23367 ( .C1(n20657), .C2(n20428), .A(n20415), .B(n20414), .ZN(
        P1_U3109) );
  AOI22_X1 U23368 ( .A1(n20626), .A2(n20423), .B1(n20625), .B2(n20422), .ZN(
        n20418) );
  AOI22_X1 U23369 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20416), .ZN(n20417) );
  OAI211_X1 U23370 ( .C1(n20538), .C2(n20428), .A(n20418), .B(n20417), .ZN(
        P1_U3110) );
  AOI22_X1 U23371 ( .A1(n20632), .A2(n20423), .B1(n20631), .B2(n20422), .ZN(
        n20421) );
  AOI22_X1 U23372 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20419), .ZN(n20420) );
  OAI211_X1 U23373 ( .C1(n20543), .C2(n20428), .A(n20421), .B(n20420), .ZN(
        P1_U3111) );
  AOI22_X1 U23374 ( .A1(n20661), .A2(n20423), .B1(n20658), .B2(n20422), .ZN(
        n20427) );
  AOI22_X1 U23375 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20425), .B1(
        n20424), .B2(n20662), .ZN(n20426) );
  OAI211_X1 U23376 ( .C1(n20668), .C2(n20428), .A(n20427), .B(n20426), .ZN(
        P1_U3112) );
  NOR3_X1 U23377 ( .A1(n20501), .A2(n15765), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20475) );
  NAND2_X1 U23378 ( .A1(n20553), .A2(n20475), .ZN(n20459) );
  OAI22_X1 U23379 ( .A1(n20460), .A2(n20515), .B1(n20459), .B2(n20503), .ZN(
        n20430) );
  INV_X1 U23380 ( .A(n20430), .ZN(n20440) );
  NAND2_X1 U23381 ( .A1(n20485), .A2(n20460), .ZN(n20431) );
  AOI21_X1 U23382 ( .B1(n20431), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20556), 
        .ZN(n20434) );
  NAND2_X1 U23383 ( .A1(n20470), .A2(n20594), .ZN(n20437) );
  AOI22_X1 U23384 ( .A1(n20434), .A2(n20437), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20459), .ZN(n20432) );
  OAI21_X1 U23385 ( .B1(n20501), .B2(n20435), .A(P1_STATE2_REG_2__SCAN_IN), 
        .ZN(n20597) );
  NAND3_X1 U23386 ( .A1(n20433), .A2(n20432), .A3(n20597), .ZN(n20463) );
  INV_X1 U23387 ( .A(n20434), .ZN(n20438) );
  OR2_X1 U23388 ( .A1(n20435), .A2(n20501), .ZN(n20588) );
  OAI22_X1 U23389 ( .A1(n20438), .A2(n20437), .B1(n20436), .B2(n20588), .ZN(
        n20462) );
  AOI22_X1 U23390 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20463), .B1(
        n20592), .B2(n20462), .ZN(n20439) );
  OAI211_X1 U23391 ( .C1(n20604), .C2(n20485), .A(n20440), .B(n20439), .ZN(
        P1_U3113) );
  OAI22_X1 U23392 ( .A1(n20460), .A2(n20520), .B1(n20459), .B2(n20516), .ZN(
        n20441) );
  INV_X1 U23393 ( .A(n20441), .ZN(n20443) );
  AOI22_X1 U23394 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20463), .B1(
        n20606), .B2(n20462), .ZN(n20442) );
  OAI211_X1 U23395 ( .C1(n20610), .C2(n20485), .A(n20443), .B(n20442), .ZN(
        P1_U3114) );
  OAI22_X1 U23396 ( .A1(n20485), .A2(n20614), .B1(n20521), .B2(n20459), .ZN(
        n20444) );
  INV_X1 U23397 ( .A(n20444), .ZN(n20446) );
  AOI22_X1 U23398 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20463), .B1(
        n20647), .B2(n20462), .ZN(n20445) );
  OAI211_X1 U23399 ( .C1(n20651), .C2(n20460), .A(n20446), .B(n20445), .ZN(
        P1_U3115) );
  OAI22_X1 U23400 ( .A1(n20460), .A2(n20529), .B1(n20459), .B2(n20525), .ZN(
        n20447) );
  INV_X1 U23401 ( .A(n20447), .ZN(n20449) );
  AOI22_X1 U23402 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20463), .B1(
        n20616), .B2(n20462), .ZN(n20448) );
  OAI211_X1 U23403 ( .C1(n20620), .C2(n20485), .A(n20449), .B(n20448), .ZN(
        P1_U3116) );
  OAI22_X1 U23404 ( .A1(n20460), .A2(n20657), .B1(n20459), .B2(n20530), .ZN(
        n20450) );
  INV_X1 U23405 ( .A(n20450), .ZN(n20452) );
  AOI22_X1 U23406 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20463), .B1(
        n20653), .B2(n20462), .ZN(n20451) );
  OAI211_X1 U23407 ( .C1(n20624), .C2(n20485), .A(n20452), .B(n20451), .ZN(
        P1_U3117) );
  OAI22_X1 U23408 ( .A1(n20460), .A2(n20538), .B1(n20459), .B2(n20534), .ZN(
        n20453) );
  INV_X1 U23409 ( .A(n20453), .ZN(n20455) );
  AOI22_X1 U23410 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20463), .B1(
        n20626), .B2(n20462), .ZN(n20454) );
  OAI211_X1 U23411 ( .C1(n20630), .C2(n20485), .A(n20455), .B(n20454), .ZN(
        P1_U3118) );
  OAI22_X1 U23412 ( .A1(n20460), .A2(n20543), .B1(n20459), .B2(n20539), .ZN(
        n20456) );
  INV_X1 U23413 ( .A(n20456), .ZN(n20458) );
  AOI22_X1 U23414 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20463), .B1(
        n20632), .B2(n20462), .ZN(n20457) );
  OAI211_X1 U23415 ( .C1(n20636), .C2(n20485), .A(n20458), .B(n20457), .ZN(
        P1_U3119) );
  OAI22_X1 U23416 ( .A1(n20460), .A2(n20668), .B1(n20459), .B2(n20545), .ZN(
        n20461) );
  INV_X1 U23417 ( .A(n20461), .ZN(n20465) );
  AOI22_X1 U23418 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20463), .B1(
        n20661), .B2(n20462), .ZN(n20464) );
  OAI211_X1 U23419 ( .C1(n20644), .C2(n20485), .A(n20465), .B(n20464), .ZN(
        P1_U3120) );
  NOR2_X1 U23420 ( .A1(n20468), .A2(n20501), .ZN(n20494) );
  AOI21_X1 U23421 ( .B1(n20470), .B2(n20469), .A(n20494), .ZN(n20472) );
  INV_X1 U23422 ( .A(n20475), .ZN(n20471) );
  OAI22_X1 U23423 ( .A1(n20472), .A2(n20556), .B1(n20471), .B2(n20760), .ZN(
        n20495) );
  AOI22_X1 U23424 ( .A1(n20592), .A2(n20495), .B1(n20591), .B2(n20494), .ZN(
        n20478) );
  AND2_X1 U23425 ( .A1(n20474), .A2(n20473), .ZN(n20476) );
  OAI21_X1 U23426 ( .B1(n20476), .B2(n20475), .A(n20561), .ZN(n20497) );
  AOI22_X1 U23427 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20497), .B1(
        n20496), .B2(n20601), .ZN(n20477) );
  OAI211_X1 U23428 ( .C1(n20604), .C2(n20551), .A(n20478), .B(n20477), .ZN(
        P1_U3121) );
  AOI22_X1 U23429 ( .A1(n20606), .A2(n20495), .B1(n20605), .B2(n20494), .ZN(
        n20481) );
  INV_X1 U23430 ( .A(n20551), .ZN(n20482) );
  AOI22_X1 U23431 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20497), .B1(
        n20482), .B2(n20479), .ZN(n20480) );
  OAI211_X1 U23432 ( .C1(n20520), .C2(n20485), .A(n20481), .B(n20480), .ZN(
        P1_U3122) );
  AOI22_X1 U23433 ( .A1(n20647), .A2(n20495), .B1(n20646), .B2(n20494), .ZN(
        n20484) );
  AOI22_X1 U23434 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20497), .B1(
        n20482), .B2(n20648), .ZN(n20483) );
  OAI211_X1 U23435 ( .C1(n20651), .C2(n20485), .A(n20484), .B(n20483), .ZN(
        P1_U3123) );
  AOI22_X1 U23436 ( .A1(n20616), .A2(n20495), .B1(n20615), .B2(n20494), .ZN(
        n20487) );
  AOI22_X1 U23437 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20497), .B1(
        n20496), .B2(n20617), .ZN(n20486) );
  OAI211_X1 U23438 ( .C1(n20620), .C2(n20551), .A(n20487), .B(n20486), .ZN(
        P1_U3124) );
  AOI22_X1 U23439 ( .A1(n20653), .A2(n20495), .B1(n20652), .B2(n20494), .ZN(
        n20489) );
  AOI22_X1 U23440 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20497), .B1(
        n20496), .B2(n20621), .ZN(n20488) );
  OAI211_X1 U23441 ( .C1(n20624), .C2(n20551), .A(n20489), .B(n20488), .ZN(
        P1_U3125) );
  AOI22_X1 U23442 ( .A1(n20626), .A2(n20495), .B1(n20625), .B2(n20494), .ZN(
        n20491) );
  AOI22_X1 U23443 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20497), .B1(
        n20496), .B2(n20627), .ZN(n20490) );
  OAI211_X1 U23444 ( .C1(n20630), .C2(n20551), .A(n20491), .B(n20490), .ZN(
        P1_U3126) );
  AOI22_X1 U23445 ( .A1(n20632), .A2(n20495), .B1(n20631), .B2(n20494), .ZN(
        n20493) );
  AOI22_X1 U23446 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20497), .B1(
        n20496), .B2(n20633), .ZN(n20492) );
  OAI211_X1 U23447 ( .C1(n20636), .C2(n20551), .A(n20493), .B(n20492), .ZN(
        P1_U3127) );
  AOI22_X1 U23448 ( .A1(n20661), .A2(n20495), .B1(n20658), .B2(n20494), .ZN(
        n20499) );
  AOI22_X1 U23449 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20497), .B1(
        n20496), .B2(n20639), .ZN(n20498) );
  OAI211_X1 U23450 ( .C1(n20644), .C2(n20551), .A(n20499), .B(n20498), .ZN(
        P1_U3128) );
  NOR3_X1 U23451 ( .A1(n20502), .A2(n20501), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20562) );
  NAND2_X1 U23452 ( .A1(n20553), .A2(n20562), .ZN(n20544) );
  OAI22_X1 U23453 ( .A1(n20564), .A2(n20604), .B1(n20503), .B2(n20544), .ZN(
        n20504) );
  INV_X1 U23454 ( .A(n20504), .ZN(n20514) );
  INV_X1 U23455 ( .A(n20510), .ZN(n20508) );
  AOI21_X1 U23456 ( .B1(n20551), .B2(n20564), .A(n20761), .ZN(n20505) );
  NOR2_X1 U23457 ( .A1(n20505), .A2(n20556), .ZN(n20509) );
  OR2_X1 U23458 ( .A1(n20506), .A2(n20594), .ZN(n20511) );
  AOI22_X1 U23459 ( .A1(n20509), .A2(n20511), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20544), .ZN(n20507) );
  OAI211_X1 U23460 ( .C1(n20508), .C2(n20760), .A(n20598), .B(n20507), .ZN(
        n20548) );
  INV_X1 U23461 ( .A(n20509), .ZN(n20512) );
  AOI22_X1 U23462 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20548), .B1(
        n20592), .B2(n20547), .ZN(n20513) );
  OAI211_X1 U23463 ( .C1(n20515), .C2(n20551), .A(n20514), .B(n20513), .ZN(
        P1_U3129) );
  OAI22_X1 U23464 ( .A1(n20564), .A2(n20610), .B1(n20516), .B2(n20544), .ZN(
        n20517) );
  INV_X1 U23465 ( .A(n20517), .ZN(n20519) );
  AOI22_X1 U23466 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20548), .B1(
        n20606), .B2(n20547), .ZN(n20518) );
  OAI211_X1 U23467 ( .C1(n20520), .C2(n20551), .A(n20519), .B(n20518), .ZN(
        P1_U3130) );
  OAI22_X1 U23468 ( .A1(n20564), .A2(n20614), .B1(n20521), .B2(n20544), .ZN(
        n20522) );
  INV_X1 U23469 ( .A(n20522), .ZN(n20524) );
  AOI22_X1 U23470 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20548), .B1(
        n20647), .B2(n20547), .ZN(n20523) );
  OAI211_X1 U23471 ( .C1(n20651), .C2(n20551), .A(n20524), .B(n20523), .ZN(
        P1_U3131) );
  OAI22_X1 U23472 ( .A1(n20564), .A2(n20620), .B1(n20525), .B2(n20544), .ZN(
        n20526) );
  INV_X1 U23473 ( .A(n20526), .ZN(n20528) );
  AOI22_X1 U23474 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20548), .B1(
        n20616), .B2(n20547), .ZN(n20527) );
  OAI211_X1 U23475 ( .C1(n20529), .C2(n20551), .A(n20528), .B(n20527), .ZN(
        P1_U3132) );
  OAI22_X1 U23476 ( .A1(n20564), .A2(n20624), .B1(n20530), .B2(n20544), .ZN(
        n20531) );
  INV_X1 U23477 ( .A(n20531), .ZN(n20533) );
  AOI22_X1 U23478 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20548), .B1(
        n20653), .B2(n20547), .ZN(n20532) );
  OAI211_X1 U23479 ( .C1(n20657), .C2(n20551), .A(n20533), .B(n20532), .ZN(
        P1_U3133) );
  OAI22_X1 U23480 ( .A1(n20564), .A2(n20630), .B1(n20534), .B2(n20544), .ZN(
        n20535) );
  INV_X1 U23481 ( .A(n20535), .ZN(n20537) );
  AOI22_X1 U23482 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20548), .B1(
        n20626), .B2(n20547), .ZN(n20536) );
  OAI211_X1 U23483 ( .C1(n20538), .C2(n20551), .A(n20537), .B(n20536), .ZN(
        P1_U3134) );
  OAI22_X1 U23484 ( .A1(n20564), .A2(n20636), .B1(n20539), .B2(n20544), .ZN(
        n20540) );
  INV_X1 U23485 ( .A(n20540), .ZN(n20542) );
  AOI22_X1 U23486 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20548), .B1(
        n20632), .B2(n20547), .ZN(n20541) );
  OAI211_X1 U23487 ( .C1(n20543), .C2(n20551), .A(n20542), .B(n20541), .ZN(
        P1_U3135) );
  OAI22_X1 U23488 ( .A1(n20564), .A2(n20644), .B1(n20545), .B2(n20544), .ZN(
        n20546) );
  INV_X1 U23489 ( .A(n20546), .ZN(n20550) );
  AOI22_X1 U23490 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20548), .B1(
        n20661), .B2(n20547), .ZN(n20549) );
  OAI211_X1 U23491 ( .C1(n20668), .C2(n20551), .A(n20550), .B(n20549), .ZN(
        P1_U3136) );
  INV_X1 U23492 ( .A(n20562), .ZN(n20555) );
  NOR2_X1 U23493 ( .A1(n20553), .A2(n20555), .ZN(n20579) );
  AOI21_X1 U23494 ( .B1(n20595), .B2(n20554), .A(n20579), .ZN(n20557) );
  OAI22_X1 U23495 ( .A1(n20557), .A2(n20556), .B1(n20555), .B2(n20760), .ZN(
        n20580) );
  AOI22_X1 U23496 ( .A1(n20592), .A2(n20580), .B1(n20591), .B2(n20579), .ZN(
        n20566) );
  INV_X1 U23497 ( .A(n20558), .ZN(n20560) );
  NOR3_X1 U23498 ( .A1(n20560), .A2(n20761), .A3(n20559), .ZN(n20563) );
  OAI21_X1 U23499 ( .B1(n20563), .B2(n20562), .A(n20561), .ZN(n20582) );
  AOI22_X1 U23500 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20582), .B1(
        n20581), .B2(n20601), .ZN(n20565) );
  OAI211_X1 U23501 ( .C1(n20604), .C2(n20600), .A(n20566), .B(n20565), .ZN(
        P1_U3137) );
  AOI22_X1 U23502 ( .A1(n20606), .A2(n20580), .B1(n20605), .B2(n20579), .ZN(
        n20568) );
  AOI22_X1 U23503 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20582), .B1(
        n20581), .B2(n20607), .ZN(n20567) );
  OAI211_X1 U23504 ( .C1(n20610), .C2(n20600), .A(n20568), .B(n20567), .ZN(
        P1_U3138) );
  AOI22_X1 U23505 ( .A1(n20647), .A2(n20580), .B1(n20646), .B2(n20579), .ZN(
        n20570) );
  AOI22_X1 U23506 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20582), .B1(
        n20581), .B2(n20611), .ZN(n20569) );
  OAI211_X1 U23507 ( .C1(n20614), .C2(n20600), .A(n20570), .B(n20569), .ZN(
        P1_U3139) );
  AOI22_X1 U23508 ( .A1(n20616), .A2(n20580), .B1(n20615), .B2(n20579), .ZN(
        n20572) );
  AOI22_X1 U23509 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20582), .B1(
        n20581), .B2(n20617), .ZN(n20571) );
  OAI211_X1 U23510 ( .C1(n20620), .C2(n20600), .A(n20572), .B(n20571), .ZN(
        P1_U3140) );
  AOI22_X1 U23511 ( .A1(n20653), .A2(n20580), .B1(n20652), .B2(n20579), .ZN(
        n20574) );
  AOI22_X1 U23512 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20582), .B1(
        n20581), .B2(n20621), .ZN(n20573) );
  OAI211_X1 U23513 ( .C1(n20624), .C2(n20600), .A(n20574), .B(n20573), .ZN(
        P1_U3141) );
  AOI22_X1 U23514 ( .A1(n20626), .A2(n20580), .B1(n20625), .B2(n20579), .ZN(
        n20576) );
  AOI22_X1 U23515 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20582), .B1(
        n20581), .B2(n20627), .ZN(n20575) );
  OAI211_X1 U23516 ( .C1(n20630), .C2(n20600), .A(n20576), .B(n20575), .ZN(
        P1_U3142) );
  AOI22_X1 U23517 ( .A1(n20632), .A2(n20580), .B1(n20631), .B2(n20579), .ZN(
        n20578) );
  AOI22_X1 U23518 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20582), .B1(
        n20581), .B2(n20633), .ZN(n20577) );
  OAI211_X1 U23519 ( .C1(n20636), .C2(n20600), .A(n20578), .B(n20577), .ZN(
        P1_U3143) );
  AOI22_X1 U23520 ( .A1(n20661), .A2(n20580), .B1(n20658), .B2(n20579), .ZN(
        n20584) );
  AOI22_X1 U23521 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20582), .B1(
        n20581), .B2(n20639), .ZN(n20583) );
  OAI211_X1 U23522 ( .C1(n20644), .C2(n20600), .A(n20584), .B(n20583), .ZN(
        P1_U3144) );
  NAND3_X1 U23523 ( .A1(n20595), .A2(n20594), .A3(n20585), .ZN(n20586) );
  OAI21_X1 U23524 ( .B1(n20588), .B2(n20587), .A(n20586), .ZN(n20638) );
  INV_X1 U23525 ( .A(n20589), .ZN(n20590) );
  NOR2_X1 U23526 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20590), .ZN(
        n20637) );
  AOI22_X1 U23527 ( .A1(n20592), .A2(n20638), .B1(n20591), .B2(n20637), .ZN(
        n20603) );
  AOI21_X1 U23528 ( .B1(n20667), .B2(n20600), .A(n20761), .ZN(n20593) );
  AOI21_X1 U23529 ( .B1(n20595), .B2(n20594), .A(n20593), .ZN(n20596) );
  NOR2_X1 U23530 ( .A1(n20596), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20599) );
  AOI22_X1 U23531 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20641), .B1(
        n20640), .B2(n20601), .ZN(n20602) );
  OAI211_X1 U23532 ( .C1(n20604), .C2(n20667), .A(n20603), .B(n20602), .ZN(
        P1_U3145) );
  AOI22_X1 U23533 ( .A1(n20606), .A2(n20638), .B1(n20605), .B2(n20637), .ZN(
        n20609) );
  AOI22_X1 U23534 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20641), .B1(
        n20640), .B2(n20607), .ZN(n20608) );
  OAI211_X1 U23535 ( .C1(n20610), .C2(n20667), .A(n20609), .B(n20608), .ZN(
        P1_U3146) );
  AOI22_X1 U23536 ( .A1(n20647), .A2(n20638), .B1(n20646), .B2(n20637), .ZN(
        n20613) );
  AOI22_X1 U23537 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20641), .B1(
        n20640), .B2(n20611), .ZN(n20612) );
  OAI211_X1 U23538 ( .C1(n20614), .C2(n20667), .A(n20613), .B(n20612), .ZN(
        P1_U3147) );
  AOI22_X1 U23539 ( .A1(n20616), .A2(n20638), .B1(n20615), .B2(n20637), .ZN(
        n20619) );
  AOI22_X1 U23540 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20641), .B1(
        n20640), .B2(n20617), .ZN(n20618) );
  OAI211_X1 U23541 ( .C1(n20620), .C2(n20667), .A(n20619), .B(n20618), .ZN(
        P1_U3148) );
  AOI22_X1 U23542 ( .A1(n20653), .A2(n20638), .B1(n20652), .B2(n20637), .ZN(
        n20623) );
  AOI22_X1 U23543 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20641), .B1(
        n20640), .B2(n20621), .ZN(n20622) );
  OAI211_X1 U23544 ( .C1(n20624), .C2(n20667), .A(n20623), .B(n20622), .ZN(
        P1_U3149) );
  AOI22_X1 U23545 ( .A1(n20626), .A2(n20638), .B1(n20625), .B2(n20637), .ZN(
        n20629) );
  AOI22_X1 U23546 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20641), .B1(
        n20640), .B2(n20627), .ZN(n20628) );
  OAI211_X1 U23547 ( .C1(n20630), .C2(n20667), .A(n20629), .B(n20628), .ZN(
        P1_U3150) );
  AOI22_X1 U23548 ( .A1(n20632), .A2(n20638), .B1(n20631), .B2(n20637), .ZN(
        n20635) );
  AOI22_X1 U23549 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20641), .B1(
        n20640), .B2(n20633), .ZN(n20634) );
  OAI211_X1 U23550 ( .C1(n20636), .C2(n20667), .A(n20635), .B(n20634), .ZN(
        P1_U3151) );
  AOI22_X1 U23551 ( .A1(n20661), .A2(n20638), .B1(n20658), .B2(n20637), .ZN(
        n20643) );
  AOI22_X1 U23552 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20641), .B1(
        n20640), .B2(n20639), .ZN(n20642) );
  OAI211_X1 U23553 ( .C1(n20644), .C2(n20667), .A(n20643), .B(n20642), .ZN(
        P1_U3152) );
  INV_X1 U23554 ( .A(n20645), .ZN(n20660) );
  AOI22_X1 U23555 ( .A1(n20647), .A2(n20660), .B1(n20659), .B2(n20646), .ZN(
        n20650) );
  AOI22_X1 U23556 ( .A1(n20664), .A2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n20663), .B2(n20648), .ZN(n20649) );
  OAI211_X1 U23557 ( .C1(n20651), .C2(n20667), .A(n20650), .B(n20649), .ZN(
        P1_U3155) );
  AOI22_X1 U23558 ( .A1(n20653), .A2(n20660), .B1(n20659), .B2(n20652), .ZN(
        n20656) );
  AOI22_X1 U23559 ( .A1(n20664), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n20663), .B2(n20654), .ZN(n20655) );
  OAI211_X1 U23560 ( .C1(n20657), .C2(n20667), .A(n20656), .B(n20655), .ZN(
        P1_U3157) );
  AOI22_X1 U23561 ( .A1(n20661), .A2(n20660), .B1(n20659), .B2(n20658), .ZN(
        n20666) );
  AOI22_X1 U23562 ( .A1(n20664), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n20663), .B2(n20662), .ZN(n20665) );
  OAI211_X1 U23563 ( .C1(n20668), .C2(n20667), .A(n20666), .B(n20665), .ZN(
        P1_U3160) );
  NOR2_X1 U23564 ( .A1(n9755), .A2(n20669), .ZN(n20671) );
  OAI21_X1 U23565 ( .B1(n20671), .B2(n20760), .A(n20670), .ZN(P1_U3163) );
  AND2_X1 U23566 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20672), .ZN(
        P1_U3164) );
  AND2_X1 U23567 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20672), .ZN(
        P1_U3165) );
  INV_X1 U23568 ( .A(P1_DATAWIDTH_REG_29__SCAN_IN), .ZN(n20945) );
  NOR2_X1 U23569 ( .A1(n20743), .A2(n20945), .ZN(P1_U3166) );
  AND2_X1 U23570 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20672), .ZN(
        P1_U3167) );
  AND2_X1 U23571 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20672), .ZN(
        P1_U3168) );
  INV_X1 U23572 ( .A(P1_DATAWIDTH_REG_26__SCAN_IN), .ZN(n20813) );
  NOR2_X1 U23573 ( .A1(n20743), .A2(n20813), .ZN(P1_U3169) );
  AND2_X1 U23574 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20672), .ZN(
        P1_U3170) );
  AND2_X1 U23575 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20672), .ZN(
        P1_U3171) );
  AND2_X1 U23576 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20672), .ZN(
        P1_U3172) );
  AND2_X1 U23577 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20672), .ZN(
        P1_U3173) );
  AND2_X1 U23578 ( .A1(P1_DATAWIDTH_REG_21__SCAN_IN), .A2(n20672), .ZN(
        P1_U3174) );
  AND2_X1 U23579 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20672), .ZN(
        P1_U3175) );
  AND2_X1 U23580 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20672), .ZN(
        P1_U3176) );
  AND2_X1 U23581 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20672), .ZN(
        P1_U3177) );
  AND2_X1 U23582 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20672), .ZN(
        P1_U3178) );
  AND2_X1 U23583 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20672), .ZN(
        P1_U3179) );
  AND2_X1 U23584 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20672), .ZN(
        P1_U3180) );
  AND2_X1 U23585 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20672), .ZN(
        P1_U3181) );
  INV_X1 U23586 ( .A(P1_DATAWIDTH_REG_13__SCAN_IN), .ZN(n20921) );
  NOR2_X1 U23587 ( .A1(n20743), .A2(n20921), .ZN(P1_U3182) );
  AND2_X1 U23588 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20672), .ZN(
        P1_U3183) );
  AND2_X1 U23589 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20672), .ZN(
        P1_U3184) );
  AND2_X1 U23590 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20672), .ZN(
        P1_U3185) );
  AND2_X1 U23591 ( .A1(n20672), .A2(P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(P1_U3186) );
  AND2_X1 U23592 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20672), .ZN(P1_U3187) );
  AND2_X1 U23593 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20672), .ZN(P1_U3188) );
  AND2_X1 U23594 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20672), .ZN(P1_U3189) );
  AND2_X1 U23595 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20672), .ZN(P1_U3190) );
  AND2_X1 U23596 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20672), .ZN(P1_U3191) );
  AND2_X1 U23597 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20672), .ZN(P1_U3192) );
  AND2_X1 U23598 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20672), .ZN(P1_U3193) );
  NAND2_X1 U23599 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20673), .ZN(n20681) );
  INV_X1 U23600 ( .A(n20681), .ZN(n20678) );
  INV_X1 U23601 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20680) );
  OAI22_X1 U23602 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20682), .B1(n20674), 
        .B2(n20687), .ZN(n20675) );
  NOR3_X1 U23603 ( .A1(n20676), .A2(n20680), .A3(n20675), .ZN(n20677) );
  OAI22_X1 U23604 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20678), .B1(n20771), 
        .B2(n20677), .ZN(P1_U3194) );
  OAI211_X1 U23605 ( .C1(NA), .C2(n20767), .A(P1_STATE_REG_1__SCAN_IN), .B(
        n20688), .ZN(n20679) );
  OAI211_X1 U23606 ( .C1(P1_STATE_REG_2__SCAN_IN), .C2(n20680), .A(
        P1_STATE_REG_0__SCAN_IN), .B(n20679), .ZN(n20686) );
  OAI211_X1 U23607 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n20682), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20681), .ZN(n20685) );
  NAND4_X1 U23608 ( .A1(P1_REQUESTPENDING_REG_SCAN_IN), .A2(
        P1_STATE_REG_0__SCAN_IN), .A3(n20683), .A4(n20682), .ZN(n20684) );
  OAI211_X1 U23609 ( .C1(n20687), .C2(n20686), .A(n20685), .B(n20684), .ZN(
        P1_U3196) );
  OR2_X1 U23610 ( .A1(n20732), .A2(P1_STATE_REG_2__SCAN_IN), .ZN(n20734) );
  OR2_X1 U23611 ( .A1(n20688), .A2(n20732), .ZN(n20729) );
  AOI222_X1 U23612 ( .A1(n20727), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_0__SCAN_IN), .B2(n20732), .C1(P1_REIP_REG_1__SCAN_IN), 
        .C2(n20731), .ZN(n20689) );
  INV_X1 U23613 ( .A(n20689), .ZN(P1_U3197) );
  AOI222_X1 U23614 ( .A1(n20731), .A2(P1_REIP_REG_2__SCAN_IN), .B1(
        P1_ADDRESS_REG_1__SCAN_IN), .B2(n20732), .C1(P1_REIP_REG_3__SCAN_IN), 
        .C2(n20727), .ZN(n20690) );
  INV_X1 U23615 ( .A(n20690), .ZN(P1_U3198) );
  OAI222_X1 U23616 ( .A1(n20729), .A2(n20693), .B1(n20692), .B2(n20771), .C1(
        n20691), .C2(n20734), .ZN(P1_U3199) );
  AOI222_X1 U23617 ( .A1(n20731), .A2(P1_REIP_REG_4__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20732), .C1(P1_REIP_REG_5__SCAN_IN), 
        .C2(n20727), .ZN(n20694) );
  INV_X1 U23618 ( .A(n20694), .ZN(P1_U3200) );
  AOI222_X1 U23619 ( .A1(n20731), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20732), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20727), .ZN(n20695) );
  INV_X1 U23620 ( .A(n20695), .ZN(P1_U3201) );
  AOI22_X1 U23621 ( .A1(P1_ADDRESS_REG_5__SCAN_IN), .A2(n20732), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20727), .ZN(n20696) );
  OAI21_X1 U23622 ( .B1(n20697), .B2(n20729), .A(n20696), .ZN(P1_U3202) );
  AOI22_X1 U23623 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20732), .B1(
        P1_REIP_REG_7__SCAN_IN), .B2(n20731), .ZN(n20698) );
  OAI21_X1 U23624 ( .B1(n20699), .B2(n20734), .A(n20698), .ZN(P1_U3203) );
  AOI222_X1 U23625 ( .A1(n20727), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_7__SCAN_IN), .B2(n20732), .C1(P1_REIP_REG_8__SCAN_IN), 
        .C2(n20731), .ZN(n20700) );
  INV_X1 U23626 ( .A(n20700), .ZN(P1_U3204) );
  AOI222_X1 U23627 ( .A1(n20731), .A2(P1_REIP_REG_9__SCAN_IN), .B1(
        P1_ADDRESS_REG_8__SCAN_IN), .B2(n20732), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20727), .ZN(n20701) );
  INV_X1 U23628 ( .A(n20701), .ZN(P1_U3205) );
  AOI222_X1 U23629 ( .A1(n20727), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20732), .C1(P1_REIP_REG_10__SCAN_IN), 
        .C2(n20731), .ZN(n20702) );
  INV_X1 U23630 ( .A(n20702), .ZN(P1_U3206) );
  AOI222_X1 U23631 ( .A1(n20731), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20732), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20727), .ZN(n20703) );
  INV_X1 U23632 ( .A(n20703), .ZN(P1_U3207) );
  AOI222_X1 U23633 ( .A1(n20731), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20732), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20727), .ZN(n20704) );
  INV_X1 U23634 ( .A(n20704), .ZN(P1_U3208) );
  AOI222_X1 U23635 ( .A1(n20731), .A2(P1_REIP_REG_13__SCAN_IN), .B1(
        P1_ADDRESS_REG_12__SCAN_IN), .B2(n20732), .C1(P1_REIP_REG_14__SCAN_IN), 
        .C2(n20727), .ZN(n20705) );
  INV_X1 U23636 ( .A(n20705), .ZN(P1_U3209) );
  AOI222_X1 U23637 ( .A1(n20731), .A2(P1_REIP_REG_14__SCAN_IN), .B1(
        P1_ADDRESS_REG_13__SCAN_IN), .B2(n20732), .C1(P1_REIP_REG_15__SCAN_IN), 
        .C2(n20727), .ZN(n20706) );
  INV_X1 U23638 ( .A(n20706), .ZN(P1_U3210) );
  AOI222_X1 U23639 ( .A1(n20731), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20732), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20727), .ZN(n20707) );
  INV_X1 U23640 ( .A(n20707), .ZN(P1_U3211) );
  AOI22_X1 U23641 ( .A1(P1_ADDRESS_REG_15__SCAN_IN), .A2(n20732), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20727), .ZN(n20708) );
  OAI21_X1 U23642 ( .B1(n14588), .B2(n20729), .A(n20708), .ZN(P1_U3212) );
  INV_X1 U23643 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20711) );
  AOI22_X1 U23644 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(n20732), .B1(
        P1_REIP_REG_17__SCAN_IN), .B2(n20731), .ZN(n20709) );
  OAI21_X1 U23645 ( .B1(n20711), .B2(n20734), .A(n20709), .ZN(P1_U3213) );
  AOI22_X1 U23646 ( .A1(P1_ADDRESS_REG_17__SCAN_IN), .A2(n20732), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20727), .ZN(n20710) );
  OAI21_X1 U23647 ( .B1(n20711), .B2(n20729), .A(n20710), .ZN(P1_U3214) );
  AOI22_X1 U23648 ( .A1(P1_ADDRESS_REG_18__SCAN_IN), .A2(n20732), .B1(
        P1_REIP_REG_19__SCAN_IN), .B2(n20731), .ZN(n20712) );
  OAI21_X1 U23649 ( .B1(n20713), .B2(n20734), .A(n20712), .ZN(P1_U3215) );
  AOI222_X1 U23650 ( .A1(n20731), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20732), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20727), .ZN(n20714) );
  INV_X1 U23651 ( .A(n20714), .ZN(P1_U3216) );
  AOI22_X1 U23652 ( .A1(P1_ADDRESS_REG_20__SCAN_IN), .A2(n20732), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(n20727), .ZN(n20715) );
  OAI21_X1 U23653 ( .B1(n20716), .B2(n20729), .A(n20715), .ZN(P1_U3217) );
  AOI22_X1 U23654 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20732), .B1(
        P1_REIP_REG_22__SCAN_IN), .B2(n20731), .ZN(n20717) );
  OAI21_X1 U23655 ( .B1(n20718), .B2(n20734), .A(n20717), .ZN(P1_U3218) );
  AOI222_X1 U23656 ( .A1(n20731), .A2(P1_REIP_REG_23__SCAN_IN), .B1(
        P1_ADDRESS_REG_22__SCAN_IN), .B2(n20732), .C1(P1_REIP_REG_24__SCAN_IN), 
        .C2(n20727), .ZN(n20719) );
  INV_X1 U23657 ( .A(n20719), .ZN(P1_U3219) );
  AOI222_X1 U23658 ( .A1(n20731), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20732), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20727), .ZN(n20720) );
  INV_X1 U23659 ( .A(n20720), .ZN(P1_U3220) );
  AOI22_X1 U23660 ( .A1(P1_ADDRESS_REG_24__SCAN_IN), .A2(n20732), .B1(
        P1_REIP_REG_26__SCAN_IN), .B2(n20727), .ZN(n20721) );
  OAI21_X1 U23661 ( .B1(n20722), .B2(n20729), .A(n20721), .ZN(P1_U3221) );
  AOI22_X1 U23662 ( .A1(P1_ADDRESS_REG_25__SCAN_IN), .A2(n20732), .B1(
        P1_REIP_REG_26__SCAN_IN), .B2(n20731), .ZN(n20723) );
  OAI21_X1 U23663 ( .B1(n20724), .B2(n20734), .A(n20723), .ZN(P1_U3222) );
  AOI222_X1 U23664 ( .A1(n20731), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20732), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20727), .ZN(n20725) );
  INV_X1 U23665 ( .A(n20725), .ZN(P1_U3223) );
  AOI222_X1 U23666 ( .A1(n20731), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20732), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20727), .ZN(n20726) );
  INV_X1 U23667 ( .A(n20726), .ZN(P1_U3224) );
  AOI22_X1 U23668 ( .A1(P1_ADDRESS_REG_28__SCAN_IN), .A2(n20732), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(n20727), .ZN(n20728) );
  OAI21_X1 U23669 ( .B1(n20730), .B2(n20729), .A(n20728), .ZN(P1_U3225) );
  AOI22_X1 U23670 ( .A1(P1_ADDRESS_REG_29__SCAN_IN), .A2(n20732), .B1(
        P1_REIP_REG_30__SCAN_IN), .B2(n20731), .ZN(n20733) );
  OAI21_X1 U23671 ( .B1(n20735), .B2(n20734), .A(n20733), .ZN(P1_U3226) );
  OAI22_X1 U23672 ( .A1(n20732), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20771), .ZN(n20736) );
  INV_X1 U23673 ( .A(n20736), .ZN(P1_U3458) );
  OAI22_X1 U23674 ( .A1(n20732), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20771), .ZN(n20737) );
  INV_X1 U23675 ( .A(n20737), .ZN(P1_U3459) );
  OAI22_X1 U23676 ( .A1(n20732), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20771), .ZN(n20738) );
  INV_X1 U23677 ( .A(n20738), .ZN(P1_U3460) );
  OAI22_X1 U23678 ( .A1(n20732), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20771), .ZN(n20739) );
  INV_X1 U23679 ( .A(n20739), .ZN(P1_U3461) );
  OAI21_X1 U23680 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20743), .A(n20741), 
        .ZN(n20740) );
  INV_X1 U23681 ( .A(n20740), .ZN(P1_U3464) );
  OAI21_X1 U23682 ( .B1(n20743), .B2(n20742), .A(n20741), .ZN(P1_U3465) );
  OAI22_X1 U23683 ( .A1(n20747), .A2(n20746), .B1(n20745), .B2(n20744), .ZN(
        n20749) );
  MUX2_X1 U23684 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20749), .S(
        n20748), .Z(P1_U3469) );
  AOI21_X1 U23685 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20751) );
  AOI22_X1 U23686 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20751), .B2(n20750), .ZN(n20754) );
  INV_X1 U23687 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20753) );
  AOI22_X1 U23688 ( .A1(n20757), .A2(n20754), .B1(n20753), .B2(n20752), .ZN(
        P1_U3481) );
  INV_X1 U23689 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20756) );
  OAI21_X1 U23690 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20757), .ZN(n20755) );
  OAI21_X1 U23691 ( .B1(n20757), .B2(n20756), .A(n20755), .ZN(P1_U3482) );
  AOI22_X1 U23692 ( .A1(n20771), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20758), 
        .B2(n20732), .ZN(P1_U3483) );
  AOI211_X1 U23693 ( .C1(n20762), .C2(n20761), .A(n20760), .B(n20759), .ZN(
        n20764) );
  OAI21_X1 U23694 ( .B1(n20764), .B2(n9755), .A(n20763), .ZN(n20770) );
  AOI211_X1 U23695 ( .C1(n20768), .C2(n20767), .A(n20766), .B(n20765), .ZN(
        n20769) );
  MUX2_X1 U23696 ( .A(n20770), .B(P1_REQUESTPENDING_REG_SCAN_IN), .S(n20769), 
        .Z(P1_U3485) );
  OAI22_X1 U23697 ( .A1(n20732), .A2(P1_MEMORYFETCH_REG_SCAN_IN), .B1(
        P1_M_IO_N_REG_SCAN_IN), .B2(n20771), .ZN(n20772) );
  INV_X1 U23698 ( .A(n20772), .ZN(P1_U3486) );
  OAI222_X1 U23699 ( .A1(n20776), .A2(n20775), .B1(n18769), .B2(n20774), .C1(
        n20773), .C2(n18765), .ZN(n20969) );
  AOI22_X1 U23700 ( .A1(n20778), .A2(keyinput97), .B1(n20933), .B2(keyinput127), .ZN(n20777) );
  OAI221_X1 U23701 ( .B1(n20778), .B2(keyinput97), .C1(n20933), .C2(
        keyinput127), .A(n20777), .ZN(n20789) );
  INV_X1 U23702 ( .A(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n20780) );
  AOI22_X1 U23703 ( .A1(n20939), .A2(keyinput76), .B1(keyinput90), .B2(n20780), 
        .ZN(n20779) );
  OAI221_X1 U23704 ( .B1(n20939), .B2(keyinput76), .C1(n20780), .C2(keyinput90), .A(n20779), .ZN(n20788) );
  INV_X1 U23705 ( .A(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n20783) );
  INV_X1 U23706 ( .A(P2_BE_N_REG_2__SCAN_IN), .ZN(n20782) );
  AOI22_X1 U23707 ( .A1(n20783), .A2(keyinput64), .B1(keyinput89), .B2(n20782), 
        .ZN(n20781) );
  OAI221_X1 U23708 ( .B1(n20783), .B2(keyinput64), .C1(n20782), .C2(keyinput89), .A(n20781), .ZN(n20787) );
  INV_X1 U23709 ( .A(P3_DATAO_REG_17__SCAN_IN), .ZN(n20785) );
  AOI22_X1 U23710 ( .A1(n20785), .A2(keyinput110), .B1(n10392), .B2(keyinput69), .ZN(n20784) );
  OAI221_X1 U23711 ( .B1(n20785), .B2(keyinput110), .C1(n10392), .C2(
        keyinput69), .A(n20784), .ZN(n20786) );
  NOR4_X1 U23712 ( .A1(n20789), .A2(n20788), .A3(n20787), .A4(n20786), .ZN(
        n20826) );
  AOI22_X1 U23713 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(keyinput72), 
        .B1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B2(keyinput99), .ZN(n20790) );
  OAI221_X1 U23714 ( .B1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(keyinput72), 
        .C1(P2_INSTQUEUE_REG_15__5__SCAN_IN), .C2(keyinput99), .A(n20790), 
        .ZN(n20800) );
  AOI22_X1 U23715 ( .A1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(keyinput114), 
        .B1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .B2(keyinput105), .ZN(n20791) );
  OAI221_X1 U23716 ( .B1(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(keyinput114), 
        .C1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .C2(keyinput105), .A(n20791), 
        .ZN(n20799) );
  AOI22_X1 U23717 ( .A1(n20793), .A2(keyinput96), .B1(n12761), .B2(keyinput75), 
        .ZN(n20792) );
  OAI221_X1 U23718 ( .B1(n20793), .B2(keyinput96), .C1(n12761), .C2(keyinput75), .A(n20792), .ZN(n20798) );
  AOI22_X1 U23719 ( .A1(n20796), .A2(keyinput81), .B1(keyinput68), .B2(n20795), 
        .ZN(n20794) );
  OAI221_X1 U23720 ( .B1(n20796), .B2(keyinput81), .C1(n20795), .C2(keyinput68), .A(n20794), .ZN(n20797) );
  NOR4_X1 U23721 ( .A1(n20800), .A2(n20799), .A3(n20798), .A4(n20797), .ZN(
        n20825) );
  INV_X1 U23722 ( .A(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n20803) );
  AOI22_X1 U23723 ( .A1(n20803), .A2(keyinput73), .B1(keyinput100), .B2(n20802), .ZN(n20801) );
  OAI221_X1 U23724 ( .B1(n20803), .B2(keyinput73), .C1(n20802), .C2(
        keyinput100), .A(n20801), .ZN(n20811) );
  AOI22_X1 U23725 ( .A1(n20805), .A2(keyinput78), .B1(keyinput79), .B2(n20900), 
        .ZN(n20804) );
  OAI221_X1 U23726 ( .B1(n20805), .B2(keyinput78), .C1(n20900), .C2(keyinput79), .A(n20804), .ZN(n20810) );
  AOI22_X1 U23727 ( .A1(n20948), .A2(keyinput83), .B1(keyinput118), .B2(n20945), .ZN(n20806) );
  OAI221_X1 U23728 ( .B1(n20948), .B2(keyinput83), .C1(n20945), .C2(
        keyinput118), .A(n20806), .ZN(n20809) );
  AOI22_X1 U23729 ( .A1(n20921), .A2(keyinput71), .B1(n20930), .B2(keyinput126), .ZN(n20807) );
  OAI221_X1 U23730 ( .B1(n20921), .B2(keyinput71), .C1(n20930), .C2(
        keyinput126), .A(n20807), .ZN(n20808) );
  NOR4_X1 U23731 ( .A1(n20811), .A2(n20810), .A3(n20809), .A4(n20808), .ZN(
        n20824) );
  INV_X1 U23732 ( .A(P1_LWORD_REG_10__SCAN_IN), .ZN(n20920) );
  AOI22_X1 U23733 ( .A1(n20813), .A2(keyinput65), .B1(n20920), .B2(keyinput94), 
        .ZN(n20812) );
  OAI221_X1 U23734 ( .B1(n20813), .B2(keyinput65), .C1(n20920), .C2(keyinput94), .A(n20812), .ZN(n20822) );
  AOI22_X1 U23735 ( .A1(n20815), .A2(keyinput120), .B1(n11347), .B2(keyinput80), .ZN(n20814) );
  OAI221_X1 U23736 ( .B1(n20815), .B2(keyinput120), .C1(n11347), .C2(
        keyinput80), .A(n20814), .ZN(n20821) );
  AOI22_X1 U23737 ( .A1(n20817), .A2(keyinput95), .B1(n13539), .B2(keyinput121), .ZN(n20816) );
  OAI221_X1 U23738 ( .B1(n20817), .B2(keyinput95), .C1(n13539), .C2(
        keyinput121), .A(n20816), .ZN(n20820) );
  AOI22_X1 U23739 ( .A1(n20931), .A2(keyinput98), .B1(n20946), .B2(keyinput85), 
        .ZN(n20818) );
  OAI221_X1 U23740 ( .B1(n20931), .B2(keyinput98), .C1(n20946), .C2(keyinput85), .A(n20818), .ZN(n20819) );
  NOR4_X1 U23741 ( .A1(n20822), .A2(n20821), .A3(n20820), .A4(n20819), .ZN(
        n20823) );
  AND4_X1 U23742 ( .A1(n20826), .A2(n20825), .A3(n20824), .A4(n20823), .ZN(
        n20967) );
  OAI22_X1 U23743 ( .A1(P2_EAX_REG_25__SCAN_IN), .A2(keyinput86), .B1(
        P1_INSTQUEUE_REG_10__0__SCAN_IN), .B2(keyinput117), .ZN(n20827) );
  AOI221_X1 U23744 ( .B1(P2_EAX_REG_25__SCAN_IN), .B2(keyinput86), .C1(
        keyinput117), .C2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A(n20827), .ZN(
        n20834) );
  OAI22_X1 U23745 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(keyinput122), 
        .B1(keyinput115), .B2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n20828)
         );
  AOI221_X1 U23746 ( .B1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(keyinput122), 
        .C1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(keyinput115), .A(n20828), 
        .ZN(n20833) );
  OAI22_X1 U23747 ( .A1(P1_EAX_REG_17__SCAN_IN), .A2(keyinput66), .B1(
        P3_REIP_REG_12__SCAN_IN), .B2(keyinput67), .ZN(n20829) );
  AOI221_X1 U23748 ( .B1(P1_EAX_REG_17__SCAN_IN), .B2(keyinput66), .C1(
        keyinput67), .C2(P3_REIP_REG_12__SCAN_IN), .A(n20829), .ZN(n20832) );
  OAI22_X1 U23749 ( .A1(P3_EAX_REG_29__SCAN_IN), .A2(keyinput107), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(keyinput101), .ZN(n20830) );
  AOI221_X1 U23750 ( .B1(P3_EAX_REG_29__SCAN_IN), .B2(keyinput107), .C1(
        keyinput101), .C2(P2_DATAO_REG_16__SCAN_IN), .A(n20830), .ZN(n20831)
         );
  NAND4_X1 U23751 ( .A1(n20834), .A2(n20833), .A3(n20832), .A4(n20831), .ZN(
        n20862) );
  OAI22_X1 U23752 ( .A1(DATAI_19_), .A2(keyinput74), .B1(
        P3_DATAO_REG_8__SCAN_IN), .B2(keyinput92), .ZN(n20835) );
  AOI221_X1 U23753 ( .B1(DATAI_19_), .B2(keyinput74), .C1(keyinput92), .C2(
        P3_DATAO_REG_8__SCAN_IN), .A(n20835), .ZN(n20842) );
  OAI22_X1 U23754 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(keyinput111), .B1(
        P3_BYTEENABLE_REG_0__SCAN_IN), .B2(keyinput108), .ZN(n20836) );
  AOI221_X1 U23755 ( .B1(P1_ADDRESS_REG_9__SCAN_IN), .B2(keyinput111), .C1(
        keyinput108), .C2(P3_BYTEENABLE_REG_0__SCAN_IN), .A(n20836), .ZN(
        n20841) );
  OAI22_X1 U23756 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(keyinput84), 
        .B1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B2(keyinput77), .ZN(n20837) );
  AOI221_X1 U23757 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(keyinput84), 
        .C1(keyinput77), .C2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A(n20837), 
        .ZN(n20840) );
  OAI22_X1 U23758 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(keyinput70), .B1(
        keyinput112), .B2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n20838) );
  AOI221_X1 U23759 ( .B1(P2_EAX_REG_10__SCAN_IN), .B2(keyinput70), .C1(
        P3_PHYADDRPOINTER_REG_27__SCAN_IN), .C2(keyinput112), .A(n20838), .ZN(
        n20839) );
  NAND4_X1 U23760 ( .A1(n20842), .A2(n20841), .A3(n20840), .A4(n20839), .ZN(
        n20861) );
  OAI22_X1 U23761 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(keyinput119), .B1(
        P2_DATAO_REG_14__SCAN_IN), .B2(keyinput104), .ZN(n20843) );
  AOI221_X1 U23762 ( .B1(P3_EAX_REG_24__SCAN_IN), .B2(keyinput119), .C1(
        keyinput104), .C2(P2_DATAO_REG_14__SCAN_IN), .A(n20843), .ZN(n20850)
         );
  OAI22_X1 U23763 ( .A1(BUF2_REG_3__SCAN_IN), .A2(keyinput82), .B1(keyinput113), .B2(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20844) );
  AOI221_X1 U23764 ( .B1(BUF2_REG_3__SCAN_IN), .B2(keyinput82), .C1(
        P2_BYTEENABLE_REG_0__SCAN_IN), .C2(keyinput113), .A(n20844), .ZN(
        n20849) );
  OAI22_X1 U23765 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(keyinput102), 
        .B1(P2_EAX_REG_20__SCAN_IN), .B2(keyinput116), .ZN(n20845) );
  AOI221_X1 U23766 ( .B1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(keyinput102), 
        .C1(keyinput116), .C2(P2_EAX_REG_20__SCAN_IN), .A(n20845), .ZN(n20848)
         );
  OAI22_X1 U23767 ( .A1(P2_ADDRESS_REG_5__SCAN_IN), .A2(keyinput106), .B1(
        keyinput103), .B2(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n20846) );
  AOI221_X1 U23768 ( .B1(P2_ADDRESS_REG_5__SCAN_IN), .B2(keyinput106), .C1(
        P1_BYTEENABLE_REG_3__SCAN_IN), .C2(keyinput103), .A(n20846), .ZN(
        n20847) );
  NAND4_X1 U23769 ( .A1(n20850), .A2(n20849), .A3(n20848), .A4(n20847), .ZN(
        n20860) );
  OAI22_X1 U23770 ( .A1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .A2(keyinput123), 
        .B1(keyinput88), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n20851) );
  AOI221_X1 U23771 ( .B1(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B2(keyinput123), 
        .C1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .C2(keyinput88), .A(n20851), 
        .ZN(n20858) );
  OAI22_X1 U23772 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(keyinput125), 
        .B1(keyinput109), .B2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n20852)
         );
  AOI221_X1 U23773 ( .B1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B2(keyinput125), 
        .C1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(keyinput109), .A(n20852), 
        .ZN(n20857) );
  OAI22_X1 U23774 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(keyinput93), .B1(
        keyinput124), .B2(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n20853) );
  AOI221_X1 U23775 ( .B1(P2_BE_N_REG_0__SCAN_IN), .B2(keyinput93), .C1(
        P3_ADDRESS_REG_23__SCAN_IN), .C2(keyinput124), .A(n20853), .ZN(n20856)
         );
  OAI22_X1 U23776 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(keyinput91), .B1(
        keyinput87), .B2(P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n20854) );
  AOI221_X1 U23777 ( .B1(P1_DATAO_REG_4__SCAN_IN), .B2(keyinput91), .C1(
        P1_DATAWIDTH_REG_9__SCAN_IN), .C2(keyinput87), .A(n20854), .ZN(n20855)
         );
  NAND4_X1 U23778 ( .A1(n20858), .A2(n20857), .A3(n20856), .A4(n20855), .ZN(
        n20859) );
  NOR4_X1 U23779 ( .A1(n20862), .A2(n20861), .A3(n20860), .A4(n20859), .ZN(
        n20966) );
  AOI22_X1 U23780 ( .A1(P3_DATAO_REG_8__SCAN_IN), .A2(keyinput28), .B1(
        P3_INSTQUEUE_REG_14__6__SCAN_IN), .B2(keyinput13), .ZN(n20863) );
  OAI221_X1 U23781 ( .B1(P3_DATAO_REG_8__SCAN_IN), .B2(keyinput28), .C1(
        P3_INSTQUEUE_REG_14__6__SCAN_IN), .C2(keyinput13), .A(n20863), .ZN(
        n20870) );
  AOI22_X1 U23782 ( .A1(BUF1_REG_5__SCAN_IN), .A2(keyinput32), .B1(
        P1_EAX_REG_8__SCAN_IN), .B2(keyinput36), .ZN(n20864) );
  OAI221_X1 U23783 ( .B1(BUF1_REG_5__SCAN_IN), .B2(keyinput32), .C1(
        P1_EAX_REG_8__SCAN_IN), .C2(keyinput36), .A(n20864), .ZN(n20869) );
  AOI22_X1 U23784 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(keyinput58), .B1(
        P2_INSTQUEUE_REG_5__2__SCAN_IN), .B2(keyinput5), .ZN(n20865) );
  OAI221_X1 U23785 ( .B1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(keyinput58), 
        .C1(P2_INSTQUEUE_REG_5__2__SCAN_IN), .C2(keyinput5), .A(n20865), .ZN(
        n20868) );
  AOI22_X1 U23786 ( .A1(P3_ADDRESS_REG_25__SCAN_IN), .A2(keyinput4), .B1(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(keyinput57), .ZN(n20866) );
  OAI221_X1 U23787 ( .B1(P3_ADDRESS_REG_25__SCAN_IN), .B2(keyinput4), .C1(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(keyinput57), .A(n20866), .ZN(
        n20867) );
  NOR4_X1 U23788 ( .A1(n20870), .A2(n20869), .A3(n20868), .A4(n20867), .ZN(
        n20898) );
  AOI22_X1 U23789 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(keyinput31), .B1(
        P2_INSTQUEUE_REG_12__1__SCAN_IN), .B2(keyinput16), .ZN(n20871) );
  OAI221_X1 U23790 ( .B1(P3_DATAWIDTH_REG_7__SCAN_IN), .B2(keyinput31), .C1(
        P2_INSTQUEUE_REG_12__1__SCAN_IN), .C2(keyinput16), .A(n20871), .ZN(
        n20878) );
  AOI22_X1 U23791 ( .A1(P1_DATAWIDTH_REG_9__SCAN_IN), .A2(keyinput23), .B1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .B2(keyinput38), .ZN(n20872) );
  OAI221_X1 U23792 ( .B1(P1_DATAWIDTH_REG_9__SCAN_IN), .B2(keyinput23), .C1(
        P2_PHYADDRPOINTER_REG_31__SCAN_IN), .C2(keyinput38), .A(n20872), .ZN(
        n20877) );
  AOI22_X1 U23793 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(keyinput25), .B1(
        P1_INSTQUEUE_REG_14__3__SCAN_IN), .B2(keyinput0), .ZN(n20873) );
  OAI221_X1 U23794 ( .B1(P2_BE_N_REG_2__SCAN_IN), .B2(keyinput25), .C1(
        P1_INSTQUEUE_REG_14__3__SCAN_IN), .C2(keyinput0), .A(n20873), .ZN(
        n20876) );
  AOI22_X1 U23795 ( .A1(BUF2_REG_3__SCAN_IN), .A2(keyinput18), .B1(
        P1_INSTQUEUE_REG_4__1__SCAN_IN), .B2(keyinput26), .ZN(n20874) );
  OAI221_X1 U23796 ( .B1(BUF2_REG_3__SCAN_IN), .B2(keyinput18), .C1(
        P1_INSTQUEUE_REG_4__1__SCAN_IN), .C2(keyinput26), .A(n20874), .ZN(
        n20875) );
  NOR4_X1 U23797 ( .A1(n20878), .A2(n20877), .A3(n20876), .A4(n20875), .ZN(
        n20897) );
  AOI22_X1 U23798 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(keyinput45), 
        .B1(P2_EAX_REG_10__SCAN_IN), .B2(keyinput6), .ZN(n20879) );
  OAI221_X1 U23799 ( .B1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(keyinput45), 
        .C1(P2_EAX_REG_10__SCAN_IN), .C2(keyinput6), .A(n20879), .ZN(n20886)
         );
  AOI22_X1 U23800 ( .A1(P1_BYTEENABLE_REG_3__SCAN_IN), .A2(keyinput39), .B1(
        P3_DATAO_REG_17__SCAN_IN), .B2(keyinput46), .ZN(n20880) );
  OAI221_X1 U23801 ( .B1(P1_BYTEENABLE_REG_3__SCAN_IN), .B2(keyinput39), .C1(
        P3_DATAO_REG_17__SCAN_IN), .C2(keyinput46), .A(n20880), .ZN(n20885) );
  AOI22_X1 U23802 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(keyinput20), 
        .B1(P2_EAX_REG_1__SCAN_IN), .B2(keyinput11), .ZN(n20881) );
  OAI221_X1 U23803 ( .B1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(keyinput20), 
        .C1(P2_EAX_REG_1__SCAN_IN), .C2(keyinput11), .A(n20881), .ZN(n20884)
         );
  AOI22_X1 U23804 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(keyinput9), .B1(
        P2_INSTQUEUE_REG_12__4__SCAN_IN), .B2(keyinput41), .ZN(n20882) );
  OAI221_X1 U23805 ( .B1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(keyinput9), .C1(
        P2_INSTQUEUE_REG_12__4__SCAN_IN), .C2(keyinput41), .A(n20882), .ZN(
        n20883) );
  NOR4_X1 U23806 ( .A1(n20886), .A2(n20885), .A3(n20884), .A4(n20883), .ZN(
        n20896) );
  AOI22_X1 U23807 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(keyinput53), 
        .B1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(keyinput17), .ZN(n20887)
         );
  OAI221_X1 U23808 ( .B1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B2(keyinput53), 
        .C1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(keyinput17), .A(n20887), 
        .ZN(n20894) );
  AOI22_X1 U23809 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(keyinput33), .B1(DATAI_19_), .B2(keyinput10), .ZN(n20888) );
  OAI221_X1 U23810 ( .B1(P3_EAX_REG_8__SCAN_IN), .B2(keyinput33), .C1(
        DATAI_19_), .C2(keyinput10), .A(n20888), .ZN(n20893) );
  AOI22_X1 U23811 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(keyinput55), .B1(
        P2_EAX_REG_25__SCAN_IN), .B2(keyinput22), .ZN(n20889) );
  OAI221_X1 U23812 ( .B1(P3_EAX_REG_24__SCAN_IN), .B2(keyinput55), .C1(
        P2_EAX_REG_25__SCAN_IN), .C2(keyinput22), .A(n20889), .ZN(n20892) );
  AOI22_X1 U23813 ( .A1(P1_ADDRESS_REG_9__SCAN_IN), .A2(keyinput47), .B1(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .B2(keyinput8), .ZN(n20890) );
  OAI221_X1 U23814 ( .B1(P1_ADDRESS_REG_9__SCAN_IN), .B2(keyinput47), .C1(
        P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(keyinput8), .A(n20890), .ZN(
        n20891) );
  NOR4_X1 U23815 ( .A1(n20894), .A2(n20893), .A3(n20892), .A4(n20891), .ZN(
        n20895) );
  NAND4_X1 U23816 ( .A1(n20898), .A2(n20897), .A3(n20896), .A4(n20895), .ZN(
        n20965) );
  AOI22_X1 U23817 ( .A1(n20901), .A2(keyinput2), .B1(keyinput15), .B2(n20900), 
        .ZN(n20899) );
  OAI221_X1 U23818 ( .B1(n20901), .B2(keyinput2), .C1(n20900), .C2(keyinput15), 
        .A(n20899), .ZN(n20906) );
  XNOR2_X1 U23819 ( .A(n20902), .B(keyinput44), .ZN(n20905) );
  XNOR2_X1 U23820 ( .A(n20903), .B(keyinput51), .ZN(n20904) );
  OR3_X1 U23821 ( .A1(n20906), .A2(n20905), .A3(n20904), .ZN(n20915) );
  AOI22_X1 U23822 ( .A1(n20909), .A2(keyinput35), .B1(keyinput24), .B2(n20908), 
        .ZN(n20907) );
  OAI221_X1 U23823 ( .B1(n20909), .B2(keyinput35), .C1(n20908), .C2(keyinput24), .A(n20907), .ZN(n20914) );
  AOI22_X1 U23824 ( .A1(n20912), .A2(keyinput48), .B1(n20911), .B2(keyinput52), 
        .ZN(n20910) );
  OAI221_X1 U23825 ( .B1(n20912), .B2(keyinput48), .C1(n20911), .C2(keyinput52), .A(n20910), .ZN(n20913) );
  NOR3_X1 U23826 ( .A1(n20915), .A2(n20914), .A3(n20913), .ZN(n20963) );
  AOI22_X1 U23827 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(keyinput14), .B1(
        n20917), .B2(keyinput50), .ZN(n20916) );
  OAI221_X1 U23828 ( .B1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B2(keyinput14), 
        .C1(n20917), .C2(keyinput50), .A(n20916), .ZN(n20928) );
  AOI22_X1 U23829 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(keyinput1), .B1(
        BUF1_REG_2__SCAN_IN), .B2(keyinput56), .ZN(n20918) );
  OAI221_X1 U23830 ( .B1(P1_DATAWIDTH_REG_26__SCAN_IN), .B2(keyinput1), .C1(
        BUF1_REG_2__SCAN_IN), .C2(keyinput56), .A(n20918), .ZN(n20927) );
  AOI22_X1 U23831 ( .A1(n20921), .A2(keyinput7), .B1(n20920), .B2(keyinput30), 
        .ZN(n20919) );
  OAI221_X1 U23832 ( .B1(n20921), .B2(keyinput7), .C1(n20920), .C2(keyinput30), 
        .A(n20919), .ZN(n20926) );
  AOI22_X1 U23833 ( .A1(n20924), .A2(keyinput29), .B1(keyinput49), .B2(n20923), 
        .ZN(n20922) );
  OAI221_X1 U23834 ( .B1(n20924), .B2(keyinput29), .C1(n20923), .C2(keyinput49), .A(n20922), .ZN(n20925) );
  NOR4_X1 U23835 ( .A1(n20928), .A2(n20927), .A3(n20926), .A4(n20925), .ZN(
        n20962) );
  AOI22_X1 U23836 ( .A1(n20931), .A2(keyinput34), .B1(n20930), .B2(keyinput62), 
        .ZN(n20929) );
  OAI221_X1 U23837 ( .B1(n20931), .B2(keyinput34), .C1(n20930), .C2(keyinput62), .A(n20929), .ZN(n20943) );
  AOI22_X1 U23838 ( .A1(n20933), .A2(keyinput63), .B1(n10300), .B2(keyinput59), 
        .ZN(n20932) );
  OAI221_X1 U23839 ( .B1(n20933), .B2(keyinput63), .C1(n10300), .C2(keyinput59), .A(n20932), .ZN(n20942) );
  AOI22_X1 U23840 ( .A1(n20936), .A2(keyinput37), .B1(n20935), .B2(keyinput43), 
        .ZN(n20934) );
  OAI221_X1 U23841 ( .B1(n20936), .B2(keyinput37), .C1(n20935), .C2(keyinput43), .A(n20934), .ZN(n20941) );
  AOI22_X1 U23842 ( .A1(n20939), .A2(keyinput12), .B1(keyinput60), .B2(n20938), 
        .ZN(n20937) );
  OAI221_X1 U23843 ( .B1(n20939), .B2(keyinput12), .C1(n20938), .C2(keyinput60), .A(n20937), .ZN(n20940) );
  NOR4_X1 U23844 ( .A1(n20943), .A2(n20942), .A3(n20941), .A4(n20940), .ZN(
        n20961) );
  AOI22_X1 U23845 ( .A1(n20946), .A2(keyinput21), .B1(keyinput54), .B2(n20945), 
        .ZN(n20944) );
  OAI221_X1 U23846 ( .B1(n20946), .B2(keyinput21), .C1(n20945), .C2(keyinput54), .A(n20944), .ZN(n20959) );
  AOI22_X1 U23847 ( .A1(n20949), .A2(keyinput40), .B1(n20948), .B2(keyinput19), 
        .ZN(n20947) );
  OAI221_X1 U23848 ( .B1(n20949), .B2(keyinput40), .C1(n20948), .C2(keyinput19), .A(n20947), .ZN(n20958) );
  INV_X1 U23849 ( .A(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n20952) );
  AOI22_X1 U23850 ( .A1(n20952), .A2(keyinput61), .B1(n20951), .B2(keyinput42), 
        .ZN(n20950) );
  OAI221_X1 U23851 ( .B1(n20952), .B2(keyinput61), .C1(n20951), .C2(keyinput42), .A(n20950), .ZN(n20957) );
  AOI22_X1 U23852 ( .A1(n20955), .A2(keyinput27), .B1(n20954), .B2(keyinput3), 
        .ZN(n20953) );
  OAI221_X1 U23853 ( .B1(n20955), .B2(keyinput27), .C1(n20954), .C2(keyinput3), 
        .A(n20953), .ZN(n20956) );
  NOR4_X1 U23854 ( .A1(n20959), .A2(n20958), .A3(n20957), .A4(n20956), .ZN(
        n20960) );
  NAND4_X1 U23855 ( .A1(n20963), .A2(n20962), .A3(n20961), .A4(n20960), .ZN(
        n20964) );
  AOI211_X1 U23856 ( .C1(n20967), .C2(n20966), .A(n20965), .B(n20964), .ZN(
        n20968) );
  XOR2_X1 U23857 ( .A(n20969), .B(n20968), .Z(P3_U3045) );
  CLKBUF_X1 U11092 ( .A(n9628), .Z(n12515) );
  INV_X1 U11086 ( .A(n11518), .ZN(n14806) );
  XNOR2_X1 U14915 ( .A(n12039), .B(n10057), .ZN(n12631) );
  CLKBUF_X2 U12326 ( .A(n10934), .Z(n10671) );
  INV_X1 U11142 ( .A(n10671), .ZN(n11687) );
  BUF_X2 U11087 ( .A(n13892), .Z(n17175) );
  CLKBUF_X1 U11089 ( .A(n11846), .Z(n13169) );
  CLKBUF_X1 U11279 ( .A(n14026), .Z(n17145) );
  CLKBUF_X1 U11427 ( .A(n10836), .Z(n11250) );
  CLKBUF_X1 U11471 ( .A(n10217), .Z(n11192) );
  CLKBUF_X1 U11968 ( .A(n14241), .Z(n14242) );
  CLKBUF_X1 U12127 ( .A(n15035), .Z(n15038) );
  CLKBUF_X2 U12253 ( .A(n17229), .Z(n9654) );
  CLKBUF_X1 U12354 ( .A(n16497), .Z(n16503) );
  INV_X2 U12705 ( .A(n18828), .ZN(n18679) );
  AND2_X2 U13072 ( .A1(n13739), .A2(n14201), .ZN(n13762) );
endmodule

