

module b14_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043, keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, 
        keyinput5, keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, 
        keyinput11, keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, 
        keyinput17, keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, 
        keyinput23, keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, 
        keyinput29, keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, 
        keyinput35, keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, 
        keyinput41, keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, 
        keyinput47, keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, 
        keyinput53, keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, 
        keyinput59, keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, 
        keyinput65, keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, 
        keyinput71, keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, 
        keyinput77, keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, 
        keyinput83, keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, 
        keyinput89, keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, 
        keyinput95, keyinput96, keyinput97, keyinput98, keyinput99, 
        keyinput100, keyinput101, keyinput102, keyinput103, keyinput104, 
        keyinput105, keyinput106, keyinput107, keyinput108, keyinput109, 
        keyinput110, keyinput111, keyinput112, keyinput113, keyinput114, 
        keyinput115, keyinput116, keyinput117, keyinput118, keyinput119, 
        keyinput120, keyinput121, keyinput122, keyinput123, keyinput124, 
        keyinput125, keyinput126, keyinput127 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN, keyinput0, keyinput1, keyinput2, keyinput3,
         keyinput4, keyinput5, keyinput6, keyinput7, keyinput8, keyinput9,
         keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019;

  XNOR2_X1 U2384 ( .A(n3686), .B(n4883), .ZN(n3674) );
  NAND2_X1 U2386 ( .A1(n2841), .A2(IR_REG_31__SCAN_IN), .ZN(n2842) );
  NAND2_X1 U2387 ( .A1(n4879), .A2(n4339), .ZN(n3334) );
  NOR2_X1 U2388 ( .A1(n3598), .A2(n3597), .ZN(n3596) );
  INV_X1 U2389 ( .A(n3720), .ZN(n3391) );
  INV_X1 U2390 ( .A(n4688), .ZN(n2309) );
  INV_X1 U2391 ( .A(n2863), .ZN(n2865) );
  INV_X1 U2392 ( .A(n4391), .ZN(n4418) );
  INV_X1 U2393 ( .A(n4881), .ZN(n4339) );
  INV_X1 U2394 ( .A(n3628), .ZN(n3634) );
  AND2_X2 U2395 ( .A1(n2783), .A2(n2782), .ZN(n4369) );
  XNOR2_X1 U2396 ( .A(n3209), .B(n4885), .ZN(n3211) );
  OAI21_X1 U2397 ( .B1(n4423), .B2(n2832), .A(n2756), .ZN(n4399) );
  NAND4_X1 U2398 ( .A1(n2578), .A2(n2577), .A3(n2576), .A4(n2575), .ZN(n4282)
         );
  XNOR2_X2 U2399 ( .A(n3188), .B(n3186), .ZN(n3187) );
  NAND2_X2 U2400 ( .A1(n4297), .A2(n3173), .ZN(n3188) );
  XNOR2_X2 U2401 ( .A(n3194), .B(n3186), .ZN(n3193) );
  NAND3_X2 U2402 ( .A1(n2293), .A2(n2292), .A3(n3178), .ZN(n3194) );
  NOR2_X2 U2403 ( .A1(n4491), .A2(n4476), .ZN(n4475) );
  AND2_X2 U2404 ( .A1(n3746), .A2(n3935), .ZN(n2457) );
  NOR2_X2 U2405 ( .A1(n2668), .A2(n3019), .ZN(n2677) );
  NAND2_X2 U2406 ( .A1(n2224), .A2(IR_REG_31__SCAN_IN), .ZN(n2518) );
  XNOR2_X2 U2407 ( .A(n2842), .B(n2843), .ZN(n2863) );
  XNOR2_X2 U2408 ( .A(n3191), .B(n4896), .ZN(n4890) );
  NAND2_X2 U2409 ( .A1(n3190), .A2(n3189), .ZN(n3191) );
  XNOR2_X2 U2410 ( .A(n4325), .B(n3704), .ZN(n3706) );
  XNOR2_X2 U2411 ( .A(n3174), .B(REG2_REG_2__SCAN_IN), .ZN(n4293) );
  NAND2_X1 U2412 ( .A1(n4928), .A2(n4929), .ZN(n4927) );
  NAND2_X1 U2413 ( .A1(n3695), .A2(n2190), .ZN(n4316) );
  AND2_X1 U2414 ( .A1(n4419), .A2(n4720), .ZN(n4382) );
  INV_X2 U2415 ( .A(n3841), .ZN(n3871) );
  NAND4_X1 U2416 ( .A1(n2549), .A2(n2548), .A3(n2547), .A4(n2546), .ZN(n4284)
         );
  NOR2_X2 U2417 ( .A1(n4023), .A2(n3553), .ZN(n2308) );
  NAND2_X2 U2418 ( .A1(n2868), .A2(n4264), .ZN(n3408) );
  INV_X1 U2419 ( .A(n3262), .ZN(n2511) );
  INV_X4 U2421 ( .A(n2903), .ZN(n2482) );
  INV_X1 U2422 ( .A(n4886), .ZN(n3186) );
  NOR2_X1 U2423 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2470)
         );
  NAND2_X2 U2424 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2317)
         );
  AND2_X1 U2425 ( .A1(n2322), .A2(n2321), .ZN(n2214) );
  CLKBUF_X1 U2426 ( .A(n3972), .Z(n3976) );
  NAND2_X1 U2427 ( .A1(n4931), .A2(n4932), .ZN(n4930) );
  NAND2_X1 U2428 ( .A1(n4927), .A2(n2227), .ZN(n4940) );
  AND2_X1 U2429 ( .A1(n4719), .A2(n2254), .ZN(n4817) );
  NAND2_X1 U2430 ( .A1(n2404), .A2(n2406), .ZN(n4365) );
  OR2_X1 U2431 ( .A1(n4411), .A2(n2821), .ZN(n2410) );
  OR2_X1 U2432 ( .A1(n4411), .A2(n2409), .ZN(n2404) );
  NAND2_X1 U2433 ( .A1(n2258), .A2(n4196), .ZN(n4411) );
  OAI21_X1 U2434 ( .B1(n4481), .B2(n4216), .A(n4174), .ZN(n4468) );
  XNOR2_X1 U2435 ( .A(n4316), .B(n3704), .ZN(n3697) );
  NAND2_X1 U2436 ( .A1(n2250), .A2(n2249), .ZN(n4501) );
  NAND2_X1 U2437 ( .A1(n3690), .A2(n3689), .ZN(n3695) );
  NAND2_X1 U2438 ( .A1(n3688), .A2(n3687), .ZN(n3690) );
  NAND2_X1 U2439 ( .A1(n3674), .A2(REG1_REG_12__SCAN_IN), .ZN(n3688) );
  NAND2_X1 U2440 ( .A1(n4547), .A2(n2729), .ZN(n4548) );
  NAND2_X1 U2441 ( .A1(n2775), .A2(n2774), .ZN(n4400) );
  NAND2_X1 U2442 ( .A1(n2245), .A2(n2242), .ZN(n4611) );
  OR2_X1 U2443 ( .A1(n2427), .A2(n2246), .ZN(n2245) );
  AND2_X1 U2444 ( .A1(n2148), .A2(n2243), .ZN(n2242) );
  NAND2_X1 U2445 ( .A1(n3443), .A2(n2220), .ZN(n4305) );
  NOR2_X1 U2446 ( .A1(n2805), .A2(n2429), .ZN(n2428) );
  AOI21_X1 U2447 ( .B1(n3577), .B2(n4151), .A(n3576), .ZN(n3496) );
  NAND2_X1 U2448 ( .A1(n2247), .A2(n2244), .ZN(n2243) );
  OAI21_X1 U2449 ( .B1(n3545), .B2(n2239), .A(n2236), .ZN(n3577) );
  OR2_X1 U2450 ( .A1(n2804), .A2(n2810), .ZN(n2805) );
  AND2_X1 U2451 ( .A1(n4661), .A2(n3652), .ZN(n3663) );
  NAND2_X1 U2452 ( .A1(n3388), .A2(n4130), .ZN(n3545) );
  OR2_X1 U2453 ( .A1(n2607), .A2(n3615), .ZN(n2608) );
  AND2_X1 U2454 ( .A1(n4653), .A2(n4208), .ZN(n2806) );
  XNOR2_X1 U2455 ( .A(n3564), .B(n3841), .ZN(n3926) );
  INV_X2 U2456 ( .A(n4957), .ZN(n2142) );
  AND2_X1 U2457 ( .A1(n2731), .A2(REG3_REG_19__SCAN_IN), .ZN(n2733) );
  AOI21_X1 U2458 ( .B1(n2238), .B2(n2240), .A(n2237), .ZN(n2236) );
  NAND2_X1 U2459 ( .A1(n4131), .A2(n4128), .ZN(n4220) );
  NOR2_X1 U2460 ( .A1(n2376), .A2(n2631), .ZN(n2371) );
  INV_X1 U2462 ( .A(n4142), .ZN(n2429) );
  OR2_X1 U2463 ( .A1(n3322), .A2(n3348), .ZN(n4131) );
  NAND2_X1 U2464 ( .A1(n3308), .A2(n3369), .ZN(n3737) );
  NAND4_X1 U2465 ( .A1(n2590), .A2(n2589), .A3(n2588), .A4(n2587), .ZN(n4283)
         );
  NAND4_X2 U2466 ( .A1(n2515), .A2(n2514), .A3(n2513), .A4(n2512), .ZN(n3712)
         );
  AND2_X1 U2467 ( .A1(n2530), .A2(n2529), .ZN(n3321) );
  NAND4_X1 U2468 ( .A1(n2617), .A2(n2616), .A3(n2615), .A4(n2614), .ZN(n4280)
         );
  NAND4_X2 U2469 ( .A1(n2569), .A2(n2568), .A3(n2567), .A4(n2566), .ZN(n4281)
         );
  OAI21_X1 U2470 ( .B1(n2144), .B2(n2521), .A(n2520), .ZN(n3720) );
  AND2_X2 U2471 ( .A1(n3724), .A2(n2903), .ZN(n2778) );
  NAND2_X1 U2472 ( .A1(n2785), .A2(IR_REG_31__SCAN_IN), .ZN(n2786) );
  BUF_X4 U2473 ( .A(n4186), .Z(n2144) );
  NAND3_X1 U2474 ( .A1(n2300), .A2(n2299), .A3(n2158), .ZN(n4186) );
  NAND2_X1 U2475 ( .A1(n2791), .A2(IR_REG_31__SCAN_IN), .ZN(n2792) );
  XNOR2_X1 U2476 ( .A(n2790), .B(IR_REG_21__SCAN_IN), .ZN(n4264) );
  XNOR2_X1 U2477 ( .A(n2849), .B(IR_REG_26__SCAN_IN), .ZN(n4878) );
  NAND2_X1 U2478 ( .A1(n2225), .A2(IR_REG_31__SCAN_IN), .ZN(n2784) );
  OR2_X1 U2479 ( .A1(n2839), .A2(IR_REG_21__SCAN_IN), .ZN(n2791) );
  NAND2_X1 U2480 ( .A1(n2256), .A2(IR_REG_31__SCAN_IN), .ZN(n2480) );
  INV_X1 U2481 ( .A(n2591), .ZN(n2349) );
  NAND4_X1 U2482 ( .A1(n2473), .A2(n2472), .A3(n2471), .A4(n2470), .ZN(n2474)
         );
  INV_X1 U2483 ( .A(IR_REG_3__SCAN_IN), .ZN(n2558) );
  NOR2_X1 U2484 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2471)
         );
  NOR2_X1 U2485 ( .A1(IR_REG_5__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2473)
         );
  INV_X1 U2486 ( .A(IR_REG_2__SCAN_IN), .ZN(n2517) );
  NOR2_X1 U2487 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_9__SCAN_IN), .ZN(n2472)
         );
  INV_X1 U2488 ( .A(IR_REG_23__SCAN_IN), .ZN(n2867) );
  INV_X1 U2489 ( .A(IR_REG_4__SCAN_IN), .ZN(n2561) );
  NOR2_X1 U2490 ( .A1(IR_REG_13__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2345)
         );
  NOR2_X1 U2491 ( .A1(IR_REG_19__SCAN_IN), .A2(IR_REG_20__SCAN_IN), .ZN(n2348)
         );
  NOR2_X1 U2492 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2347)
         );
  NOR2_X1 U2493 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2346)
         );
  XNOR2_X2 U2494 ( .A(n3198), .B(n4896), .ZN(n4893) );
  NAND2_X2 U2495 ( .A1(n3196), .A2(n3195), .ZN(n3198) );
  NAND2_X1 U2496 ( .A1(n4921), .A2(n4920), .ZN(n4919) );
  XNOR2_X1 U2497 ( .A(n4331), .B(n2700), .ZN(n4921) );
  XNOR2_X2 U2498 ( .A(n3680), .B(n3685), .ZN(n3679) );
  NAND2_X2 U2499 ( .A1(n3670), .A2(n3669), .ZN(n3680) );
  OAI21_X2 U2500 ( .B1(n4047), .B2(n4048), .A(n4049), .ZN(n3907) );
  NAND2_X1 U2501 ( .A1(n3174), .A2(REG1_REG_2__SCAN_IN), .ZN(n2228) );
  OR2_X1 U2502 ( .A1(n3174), .A2(REG1_REG_2__SCAN_IN), .ZN(n2203) );
  AND2_X4 U2503 ( .A1(n3724), .A2(n2482), .ZN(n2572) );
  INV_X2 U2504 ( .A(n2481), .ZN(n3724) );
  INV_X2 U2505 ( .A(n3755), .ZN(n3874) );
  OR2_X1 U2506 ( .A1(n4400), .A2(n4384), .ZN(n4185) );
  INV_X1 U2507 ( .A(n4074), .ZN(n2451) );
  INV_X1 U2508 ( .A(n2778), .ZN(n2832) );
  AOI21_X1 U2509 ( .B1(n2396), .B2(n2757), .A(n2168), .ZN(n2394) );
  OR2_X1 U2510 ( .A1(n3712), .A2(n3391), .ZN(n2539) );
  AND2_X1 U2511 ( .A1(n4879), .A2(n4264), .ZN(n3167) );
  AND2_X1 U2512 ( .A1(n2788), .A2(n2180), .ZN(n2291) );
  INV_X1 U2513 ( .A(IR_REG_15__SCAN_IN), .ZN(n2686) );
  AOI22_X1 U2514 ( .A1(n3745), .A2(n3933), .B1(n3744), .B2(n3743), .ZN(n3746)
         );
  XNOR2_X1 U2515 ( .A(n3445), .B(n3436), .ZN(n3301) );
  NAND2_X1 U2516 ( .A1(n2338), .A2(n2337), .ZN(n2336) );
  INV_X1 U2517 ( .A(n4904), .ZN(n2337) );
  NAND2_X1 U2518 ( .A1(n4919), .A2(n4332), .ZN(n4931) );
  AND2_X1 U2519 ( .A1(n4948), .A2(n2327), .ZN(n2326) );
  AND2_X1 U2520 ( .A1(n2333), .A2(n2328), .ZN(n2327) );
  AND2_X1 U2521 ( .A1(n2392), .A2(n2173), .ZN(n2391) );
  NAND2_X1 U2522 ( .A1(n2394), .A2(n2160), .ZN(n2393) );
  AND2_X1 U2523 ( .A1(n4202), .A2(n4254), .ZN(n4402) );
  AOI21_X1 U2524 ( .B1(n2362), .B2(n2364), .A(n2366), .ZN(n2360) );
  INV_X1 U2525 ( .A(n4678), .ZN(n4563) );
  OAI22_X1 U2526 ( .A1(n3543), .A2(n2551), .B1(n3553), .B2(n4284), .ZN(n3454)
         );
  OR2_X1 U2527 ( .A1(n3454), .A2(n4199), .ZN(n3498) );
  NAND2_X1 U2528 ( .A1(n2793), .A2(n4339), .ZN(n3574) );
  AND3_X1 U2529 ( .A1(n2873), .A2(n2872), .A3(n2871), .ZN(n2879) );
  INV_X1 U2530 ( .A(n4369), .ZN(n4392) );
  OR2_X1 U2531 ( .A1(n4386), .A2(n2832), .ZN(n2775) );
  NAND2_X1 U2532 ( .A1(n2763), .A2(n2762), .ZN(n4391) );
  INV_X1 U2533 ( .A(n4455), .ZN(n4415) );
  XNOR2_X1 U2534 ( .A(n3419), .B(n3841), .ZN(n3466) );
  NAND2_X1 U2535 ( .A1(n3951), .A2(n3950), .ZN(n2460) );
  NAND2_X1 U2536 ( .A1(n3466), .A2(n3467), .ZN(n2446) );
  INV_X1 U2537 ( .A(n4433), .ZN(n2233) );
  NOR2_X1 U2538 ( .A1(n4448), .A2(n2235), .ZN(n2234) );
  NAND2_X1 U2539 ( .A1(n4303), .A2(n2184), .ZN(n3521) );
  INV_X1 U2540 ( .A(n2823), .ZN(n2408) );
  OAI21_X1 U2541 ( .B1(n4469), .B2(n2356), .A(n2749), .ZN(n2355) );
  NAND2_X1 U2542 ( .A1(n4473), .A2(n4451), .ZN(n2357) );
  INV_X1 U2543 ( .A(n2424), .ZN(n2423) );
  AOI21_X1 U2544 ( .B1(n4216), .B2(n4174), .A(n2425), .ZN(n2424) );
  NOR2_X1 U2545 ( .A1(n2165), .A2(n2422), .ZN(n2421) );
  NOR2_X1 U2546 ( .A1(n2423), .A2(n4174), .ZN(n2422) );
  INV_X1 U2547 ( .A(n2363), .ZN(n2362) );
  OAI21_X1 U2548 ( .B1(n2159), .B2(n2364), .A(n2367), .ZN(n2363) );
  OR2_X1 U2549 ( .A1(n4484), .A2(n4745), .ZN(n2367) );
  INV_X1 U2550 ( .A(n4235), .ZN(n2249) );
  INV_X1 U2551 ( .A(n4560), .ZN(n2250) );
  NOR2_X1 U2552 ( .A1(n2248), .A2(n2403), .ZN(n2247) );
  OR2_X1 U2553 ( .A1(n3858), .A2(n4224), .ZN(n2386) );
  INV_X1 U2554 ( .A(n4136), .ZN(n2241) );
  INV_X1 U2555 ( .A(n4221), .ZN(n2238) );
  INV_X1 U2556 ( .A(n4140), .ZN(n2237) );
  OR2_X1 U2557 ( .A1(n2789), .A2(n2416), .ZN(n2415) );
  AND2_X1 U2558 ( .A1(n2305), .A2(IR_REG_31__SCAN_IN), .ZN(n2304) );
  INV_X1 U2559 ( .A(IR_REG_27__SCAN_IN), .ZN(n2305) );
  NOR2_X1 U2560 ( .A1(n4435), .A2(n4451), .ZN(n2310) );
  NAND2_X1 U2561 ( .A1(n2377), .A2(n2379), .ZN(n4547) );
  AOI21_X1 U2562 ( .B1(n2381), .B2(n2380), .A(n2166), .ZN(n2379) );
  AND2_X1 U2563 ( .A1(n4594), .A2(n4561), .ZN(n2316) );
  AND2_X1 U2564 ( .A1(n2476), .A2(n2418), .ZN(n2417) );
  INV_X1 U2565 ( .A(IR_REG_26__SCAN_IN), .ZN(n2418) );
  AND2_X1 U2566 ( .A1(n2291), .A2(n2176), .ZN(n2289) );
  OR3_X1 U2567 ( .A1(n2714), .A2(IR_REG_16__SCAN_IN), .A3(n2713), .ZN(n2725)
         );
  OAI21_X1 U2568 ( .B1(n3561), .B2(n3560), .A(n3559), .ZN(n3748) );
  XNOR2_X1 U2569 ( .A(n3467), .B(n2259), .ZN(n2260) );
  INV_X1 U2570 ( .A(n3466), .ZN(n2259) );
  NAND2_X1 U2571 ( .A1(n3917), .A2(n3819), .ZN(n4008) );
  NOR2_X2 U2572 ( .A1(n2743), .A2(n3920), .ZN(n2744) );
  NAND2_X1 U2573 ( .A1(n2733), .A2(REG3_REG_20__SCAN_IN), .ZN(n2504) );
  OAI21_X1 U2574 ( .B1(n3943), .B2(n3942), .A(n3795), .ZN(n4037) );
  OR2_X1 U2575 ( .A1(n3794), .A2(n3793), .ZN(n3795) );
  NAND2_X1 U2576 ( .A1(n2461), .A2(n2460), .ZN(n2288) );
  AOI21_X1 U2577 ( .B1(n2457), .B2(n3747), .A(n2169), .ZN(n2454) );
  INV_X1 U2578 ( .A(n3749), .ZN(n2456) );
  OR2_X1 U2579 ( .A1(n3907), .A2(n3903), .ZN(n3984) );
  NAND2_X1 U2580 ( .A1(n4008), .A2(n4011), .ZN(n3825) );
  NAND2_X1 U2581 ( .A1(n2279), .A2(n2282), .ZN(n3824) );
  AOI21_X1 U2582 ( .B1(n2287), .B2(n3814), .A(n2283), .ZN(n2282) );
  AOI21_X1 U2583 ( .B1(n3276), .B2(n3270), .A(n3269), .ZN(n3176) );
  INV_X1 U2584 ( .A(n4888), .ZN(n4287) );
  NAND2_X1 U2585 ( .A1(n2318), .A2(n2167), .ZN(n3445) );
  NAND2_X1 U2586 ( .A1(n3297), .A2(n2319), .ZN(n2318) );
  NAND2_X1 U2587 ( .A1(n3301), .A2(REG1_REG_8__SCAN_IN), .ZN(n3443) );
  XNOR2_X1 U2588 ( .A(n3521), .B(n3526), .ZN(n3447) );
  NAND2_X1 U2589 ( .A1(n3529), .A2(n3528), .ZN(n3531) );
  NAND2_X1 U2590 ( .A1(n4318), .A2(n4317), .ZN(n2338) );
  OR2_X1 U2591 ( .A1(n4333), .A2(REG2_REG_17__SCAN_IN), .ZN(n2230) );
  INV_X1 U2592 ( .A(n4476), .ZN(n4465) );
  NAND2_X1 U2593 ( .A1(n4464), .A2(n4469), .ZN(n4463) );
  AND2_X1 U2594 ( .A1(n2495), .A2(n2494), .ZN(n4487) );
  NAND2_X1 U2595 ( .A1(n2146), .A2(n2161), .ZN(n2365) );
  NOR2_X1 U2596 ( .A1(n2383), .A2(n2667), .ZN(n2382) );
  INV_X1 U2597 ( .A(n2705), .ZN(n2383) );
  AND3_X1 U2598 ( .A1(n2696), .A2(n2695), .A3(n2694), .ZN(n4609) );
  INV_X1 U2599 ( .A(n2402), .ZN(n2401) );
  OAI21_X1 U2600 ( .B1(n4164), .B2(n2403), .A(n4161), .ZN(n2402) );
  NAND2_X1 U2601 ( .A1(n4629), .A2(n2247), .ZN(n2400) );
  CLKBUF_X1 U2602 ( .A(n4625), .Z(n4626) );
  NAND2_X1 U2603 ( .A1(n2427), .A2(n4165), .ZN(n4629) );
  INV_X1 U2604 ( .A(n3593), .ZN(n3597) );
  OR2_X1 U2605 ( .A1(n4989), .A2(n4264), .ZN(n3341) );
  AND2_X1 U2606 ( .A1(n4137), .A2(n4140), .ZN(n4199) );
  AND2_X1 U2607 ( .A1(n3283), .A2(n2539), .ZN(n2540) );
  AND2_X1 U2608 ( .A1(n4136), .A2(n4133), .ZN(n4221) );
  NAND2_X1 U2609 ( .A1(n3545), .A2(n4221), .ZN(n3544) );
  NAND2_X1 U2610 ( .A1(n3369), .A2(n4978), .ZN(n3403) );
  NAND2_X1 U2611 ( .A1(n2794), .A2(n4125), .ZN(n3329) );
  NAND2_X1 U2612 ( .A1(n2315), .A2(n2314), .ZN(n2313) );
  AOI21_X1 U2613 ( .B1(n4368), .B2(n4525), .A(n2430), .ZN(n4711) );
  OAI22_X1 U2614 ( .A1(n4369), .A2(n4659), .B1(n4371), .B2(n4370), .ZN(n2430)
         );
  INV_X1 U2615 ( .A(n4384), .ZN(n4714) );
  OR2_X1 U2616 ( .A1(n3329), .A2(n2868), .ZN(n4795) );
  INV_X1 U2617 ( .A(n4795), .ZN(n4768) );
  OR2_X1 U2618 ( .A1(n4951), .A2(n4879), .ZN(n4989) );
  NAND2_X1 U2619 ( .A1(n2850), .A2(n4878), .ZN(n3326) );
  NAND2_X1 U2620 ( .A1(n2844), .A2(IR_REG_31__SCAN_IN), .ZN(n2866) );
  XNOR2_X1 U2621 ( .A(n2866), .B(n2867), .ZN(n3368) );
  AND2_X1 U2622 ( .A1(n2688), .A2(n2697), .ZN(n4330) );
  CLKBUF_X1 U2623 ( .A(n3748), .Z(n3928) );
  NAND2_X1 U2624 ( .A1(n4019), .A2(n2211), .ZN(n4020) );
  AND2_X1 U2625 ( .A1(n4021), .A2(n4018), .ZN(n2211) );
  NAND2_X1 U2626 ( .A1(n3365), .A2(n2217), .ZN(n3717) );
  OR2_X1 U2627 ( .A1(n3362), .A2(n3361), .ZN(n2217) );
  NAND2_X1 U2628 ( .A1(n4305), .A2(n4304), .ZN(n4303) );
  NAND2_X1 U2629 ( .A1(n3697), .A2(REG1_REG_14__SCAN_IN), .ZN(n4318) );
  NAND2_X1 U2630 ( .A1(n4916), .A2(n4321), .ZN(n4928) );
  NAND2_X1 U2631 ( .A1(n3225), .A2(n4888), .ZN(n4949) );
  OR2_X1 U2632 ( .A1(n4940), .A2(n2323), .ZN(n2322) );
  NAND2_X1 U2633 ( .A1(n4935), .A2(n2325), .ZN(n2323) );
  NAND2_X1 U2634 ( .A1(n2331), .A2(n2329), .ZN(n2325) );
  OR2_X1 U2635 ( .A1(n4939), .A2(n2332), .ZN(n2331) );
  AOI21_X1 U2636 ( .B1(n4940), .B2(n2154), .A(n2193), .ZN(n2321) );
  AND2_X1 U2637 ( .A1(n4948), .A2(n2328), .ZN(n2226) );
  OAI21_X1 U2638 ( .B1(n4410), .B2(n2393), .A(n2391), .ZN(n4357) );
  NAND2_X1 U2639 ( .A1(n2390), .A2(n2394), .ZN(n4381) );
  NAND2_X1 U2640 ( .A1(n2405), .A2(n2411), .ZN(n4389) );
  NAND2_X1 U2641 ( .A1(n2410), .A2(n2823), .ZN(n2413) );
  OAI21_X1 U2642 ( .B1(n4411), .B2(n4396), .A(n4397), .ZN(n4398) );
  OR2_X1 U2643 ( .A1(n3403), .A2(n3341), .ZN(n4643) );
  INV_X1 U2644 ( .A(n2382), .ZN(n2380) );
  INV_X1 U2645 ( .A(n3420), .ZN(n3870) );
  INV_X1 U2646 ( .A(n3821), .ZN(n2283) );
  NOR2_X1 U2647 ( .A1(n2284), .A2(n2281), .ZN(n2280) );
  INV_X1 U2648 ( .A(n2460), .ZN(n2281) );
  INV_X1 U2649 ( .A(n3814), .ZN(n2284) );
  INV_X1 U2650 ( .A(REG3_REG_12__SCAN_IN), .ZN(n2659) );
  INV_X1 U2651 ( .A(REG3_REG_7__SCAN_IN), .ZN(n2563) );
  OR2_X1 U2652 ( .A1(n3299), .A2(n3298), .ZN(n2319) );
  NAND2_X1 U2653 ( .A1(n4418), .A2(n2207), .ZN(n4202) );
  NAND2_X1 U2654 ( .A1(n2421), .A2(n2423), .ZN(n2419) );
  INV_X1 U2655 ( .A(n2365), .ZN(n2364) );
  INV_X1 U2656 ( .A(n4165), .ZN(n2244) );
  INV_X1 U2657 ( .A(n2247), .ZN(n2246) );
  INV_X1 U2658 ( .A(n4200), .ZN(n2403) );
  NAND2_X1 U2659 ( .A1(n2209), .A2(n2208), .ZN(n2668) );
  NOR2_X1 U2660 ( .A1(n2659), .A2(n2993), .ZN(n2208) );
  INV_X1 U2661 ( .A(n2660), .ZN(n2209) );
  OR2_X1 U2662 ( .A1(n3646), .A2(n2654), .ZN(n2658) );
  NAND2_X1 U2663 ( .A1(n3643), .A2(n2811), .ZN(n2427) );
  INV_X1 U2664 ( .A(n4712), .ZN(n2314) );
  INV_X1 U2665 ( .A(n3326), .ZN(n2861) );
  NOR2_X1 U2666 ( .A1(IR_REG_15__SCAN_IN), .A2(IR_REG_14__SCAN_IN), .ZN(n2741)
         );
  NOR2_X1 U2667 ( .A1(IR_REG_17__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .ZN(n2740)
         );
  INV_X1 U2668 ( .A(IR_REG_9__SCAN_IN), .ZN(n2628) );
  NOR2_X2 U2669 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2516)
         );
  INV_X1 U2670 ( .A(IR_REG_19__SCAN_IN), .ZN(n2925) );
  INV_X1 U2671 ( .A(REG3_REG_13__SCAN_IN), .ZN(n2993) );
  INV_X1 U2672 ( .A(IR_REG_6__SCAN_IN), .ZN(n2570) );
  INV_X1 U2673 ( .A(REG3_REG_14__SCAN_IN), .ZN(n3019) );
  AND2_X1 U2674 ( .A1(n3918), .A2(n3919), .ZN(n3814) );
  NOR2_X1 U2675 ( .A1(n2621), .A2(n3042), .ZN(n2634) );
  XNOR2_X1 U2676 ( .A(n3354), .B(n3841), .ZN(n3423) );
  INV_X1 U2677 ( .A(n4400), .ZN(n3887) );
  INV_X1 U2678 ( .A(n3321), .ZN(n3348) );
  INV_X1 U2679 ( .A(REG3_REG_21__SCAN_IN), .ZN(n3954) );
  INV_X1 U2680 ( .A(n3826), .ZN(n3873) );
  XNOR2_X1 U2681 ( .A(n3740), .B(n3871), .ZN(n3933) );
  AOI21_X1 U2682 ( .B1(n2266), .B2(n2268), .A(n2265), .ZN(n2264) );
  INV_X1 U2683 ( .A(n2450), .ZN(n2268) );
  AND3_X2 U2684 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .A3(
        REG3_REG_5__SCAN_IN), .ZN(n2583) );
  NAND2_X1 U2685 ( .A1(n2446), .A2(n2447), .ZN(n2444) );
  INV_X1 U2686 ( .A(n2446), .ZN(n2442) );
  AND2_X1 U2687 ( .A1(n2677), .A2(REG3_REG_15__SCAN_IN), .ZN(n2689) );
  OR2_X1 U2688 ( .A1(n3874), .A2(n3336), .ZN(n3344) );
  AND2_X1 U2689 ( .A1(n4229), .A2(n2231), .ZN(n4266) );
  NOR2_X1 U2690 ( .A1(n4366), .A2(n2232), .ZN(n2231) );
  NAND2_X1 U2691 ( .A1(n2234), .A2(n2233), .ZN(n2232) );
  NAND2_X1 U2692 ( .A1(n2572), .A2(REG2_REG_7__SCAN_IN), .ZN(n2569) );
  OR2_X1 U2693 ( .A1(n3524), .A2(n4799), .ZN(n2342) );
  NAND2_X1 U2694 ( .A1(n3522), .A2(n2340), .ZN(n2339) );
  INV_X1 U2695 ( .A(n3524), .ZN(n2340) );
  NAND2_X1 U2696 ( .A1(n4330), .A2(REG1_REG_15__SCAN_IN), .ZN(n2335) );
  AND2_X1 U2697 ( .A1(n3183), .A2(n3181), .ZN(n3225) );
  INV_X1 U2698 ( .A(n4322), .ZN(n2332) );
  AOI21_X1 U2699 ( .B1(n4939), .B2(n2188), .A(n2330), .ZN(n2329) );
  AND2_X1 U2700 ( .A1(n2334), .A2(n4322), .ZN(n2330) );
  INV_X1 U2701 ( .A(n2329), .ZN(n2324) );
  AND2_X1 U2702 ( .A1(n4334), .A2(REG2_REG_18__SCAN_IN), .ZN(n2333) );
  INV_X1 U2703 ( .A(n4336), .ZN(n2328) );
  AOI21_X1 U2704 ( .B1(n2411), .B2(n2408), .A(n2407), .ZN(n2406) );
  INV_X1 U2705 ( .A(n4185), .ZN(n2407) );
  NAND2_X1 U2706 ( .A1(n2206), .A2(n4254), .ZN(n2823) );
  INV_X1 U2707 ( .A(n4251), .ZN(n2206) );
  NAND2_X1 U2708 ( .A1(n4411), .A2(n2823), .ZN(n2405) );
  AND2_X1 U2709 ( .A1(n2412), .A2(n4390), .ZN(n2411) );
  NAND2_X1 U2710 ( .A1(n2821), .A2(n2823), .ZN(n2412) );
  NAND2_X1 U2711 ( .A1(n2357), .A2(n2358), .ZN(n2353) );
  INV_X1 U2712 ( .A(n2357), .ZN(n2352) );
  INV_X1 U2713 ( .A(n2355), .ZN(n2354) );
  INV_X1 U2714 ( .A(n4440), .ZN(n4435) );
  OAI21_X1 U2715 ( .B1(n4481), .B2(n2423), .A(n2421), .ZN(n4431) );
  AND2_X1 U2716 ( .A1(n2487), .A2(n2486), .ZN(n4455) );
  AND2_X1 U2717 ( .A1(n4521), .A2(n4522), .ZN(n4551) );
  NAND2_X1 U2718 ( .A1(n2689), .A2(REG3_REG_16__SCAN_IN), .ZN(n2707) );
  NAND2_X1 U2719 ( .A1(n4586), .A2(n4234), .ZN(n4560) );
  AND2_X1 U2720 ( .A1(n4237), .A2(n4234), .ZN(n4600) );
  NAND2_X1 U2721 ( .A1(n2384), .A2(n2386), .ZN(n4596) );
  NAND2_X1 U2722 ( .A1(n2385), .A2(n2387), .ZN(n2384) );
  NAND2_X1 U2723 ( .A1(n2814), .A2(n4164), .ZN(n4233) );
  NAND2_X1 U2724 ( .A1(n4629), .A2(n4160), .ZN(n2814) );
  AND2_X1 U2725 ( .A1(n4161), .A2(n4147), .ZN(n4200) );
  NAND2_X1 U2726 ( .A1(n2223), .A2(REG3_REG_9__SCAN_IN), .ZN(n2621) );
  INV_X1 U2727 ( .A(n2611), .ZN(n2223) );
  AND2_X1 U2728 ( .A1(n4672), .A2(n4674), .ZN(n4210) );
  NAND2_X1 U2729 ( .A1(n2799), .A2(n4142), .ZN(n3622) );
  INV_X1 U2730 ( .A(n2240), .ZN(n2239) );
  NOR2_X1 U2731 ( .A1(n2797), .A2(n2241), .ZN(n2240) );
  NAND2_X1 U2732 ( .A1(n2307), .A2(n2308), .ZN(n3583) );
  NOR2_X1 U2733 ( .A1(n3552), .A2(n3553), .ZN(n3551) );
  NAND2_X1 U2734 ( .A1(n2414), .A2(n2304), .ZN(n2300) );
  OAI211_X1 U2735 ( .C1(n2417), .C2(n2416), .A(n2415), .B(IR_REG_28__SCAN_IN), 
        .ZN(n2299) );
  NAND2_X1 U2736 ( .A1(n2302), .A2(n2301), .ZN(n3315) );
  NAND2_X1 U2737 ( .A1(n2143), .A2(DATAI_0_), .ZN(n2301) );
  OR2_X1 U2738 ( .A1(n2143), .A2(n2303), .ZN(n2302) );
  INV_X1 U2739 ( .A(n3895), .ZN(n4358) );
  NAND2_X1 U2740 ( .A1(n4382), .A2(n4342), .ZN(n4374) );
  NOR2_X1 U2741 ( .A1(n4374), .A2(n4350), .ZN(n4349) );
  AND2_X1 U2742 ( .A1(n4475), .A2(n2194), .ZN(n4419) );
  NAND2_X1 U2743 ( .A1(n4475), .A2(n2310), .ZN(n4439) );
  NAND2_X1 U2744 ( .A1(n4475), .A2(n4457), .ZN(n4456) );
  OR2_X1 U2745 ( .A1(n4511), .A2(n4483), .ZN(n4491) );
  INV_X1 U2746 ( .A(n4745), .ZN(n4512) );
  AND2_X1 U2747 ( .A1(n4588), .A2(n2185), .ZN(n4533) );
  AND2_X1 U2748 ( .A1(n4620), .A2(n2875), .ZN(n4588) );
  NAND2_X1 U2749 ( .A1(n4588), .A2(n2316), .ZN(n4571) );
  NAND2_X1 U2750 ( .A1(n4588), .A2(n4594), .ZN(n4589) );
  NOR2_X1 U2751 ( .A1(n4642), .A2(n3910), .ZN(n4620) );
  OR2_X1 U2752 ( .A1(n4640), .A2(n4639), .ZN(n4642) );
  INV_X1 U2753 ( .A(n3965), .ZN(n4784) );
  AND2_X1 U2754 ( .A1(n3596), .A2(n2178), .ZN(n4661) );
  NAND2_X1 U2755 ( .A1(n3596), .A2(n2145), .ZN(n4691) );
  NAND2_X1 U2756 ( .A1(n3596), .A2(n3634), .ZN(n4689) );
  AND2_X1 U2757 ( .A1(n3348), .A2(n3855), .ZN(n3393) );
  INV_X1 U2758 ( .A(IR_REG_29__SCAN_IN), .ZN(n2478) );
  AND2_X1 U2759 ( .A1(n2162), .A2(n2834), .ZN(n2463) );
  INV_X1 U2760 ( .A(n2474), .ZN(n2351) );
  NAND2_X1 U2761 ( .A1(n2290), .A2(IR_REG_31__SCAN_IN), .ZN(n2846) );
  XNOR2_X1 U2762 ( .A(n2715), .B(IR_REG_17__SCAN_IN), .ZN(n4333) );
  INV_X1 U2763 ( .A(IR_REG_13__SCAN_IN), .ZN(n2674) );
  INV_X1 U2764 ( .A(IR_REG_11__SCAN_IN), .ZN(n2649) );
  OR3_X1 U2765 ( .A1(n2618), .A2(IR_REG_8__SCAN_IN), .A3(IR_REG_7__SCAN_IN), 
        .ZN(n2627) );
  INV_X1 U2766 ( .A(IR_REG_7__SCAN_IN), .ZN(n2911) );
  CLKBUF_X1 U2767 ( .A(IR_REG_0__SCAN_IN), .Z(n2222) );
  OAI211_X1 U2768 ( .C1(n4020), .C2(n2438), .A(n2439), .B(n2437), .ZN(n3489)
         );
  NAND2_X1 U2769 ( .A1(n2189), .A2(n2445), .ZN(n2439) );
  NAND2_X1 U2770 ( .A1(n2171), .A2(n2441), .ZN(n2437) );
  NAND2_X1 U2771 ( .A1(n2441), .A2(n2445), .ZN(n2438) );
  NAND2_X1 U2772 ( .A1(n3489), .A2(n3488), .ZN(n3559) );
  INV_X1 U2773 ( .A(n4116), .ZN(n4065) );
  AOI21_X1 U2774 ( .B1(n2277), .B2(n2274), .A(n2273), .ZN(n2272) );
  INV_X1 U2775 ( .A(n4100), .ZN(n2273) );
  NAND2_X1 U2776 ( .A1(n4060), .A2(n3814), .ZN(n3917) );
  NAND2_X1 U2777 ( .A1(n2457), .A2(n2453), .ZN(n3934) );
  OR2_X1 U2778 ( .A1(n3928), .A2(n3747), .ZN(n2453) );
  AND2_X1 U2779 ( .A1(n2777), .A2(n2156), .ZN(n3894) );
  INV_X1 U2780 ( .A(n2432), .ZN(n2431) );
  INV_X1 U2781 ( .A(n3355), .ZN(n2436) );
  AOI22_X1 U2782 ( .A1(n3851), .A2(n3849), .B1(n3319), .B2(n3871), .ZN(n3356)
         );
  INV_X1 U2783 ( .A(n2461), .ZN(n3953) );
  NAND2_X1 U2784 ( .A1(n2450), .A2(n2269), .ZN(n3962) );
  NAND2_X1 U2785 ( .A1(n3928), .A2(n2448), .ZN(n2269) );
  OR2_X1 U2786 ( .A1(n2768), .A2(n2752), .ZN(n4423) );
  AND3_X1 U2787 ( .A1(n2712), .A2(n2711), .A3(n2710), .ZN(n4584) );
  NAND2_X1 U2788 ( .A1(n4020), .A2(n2447), .ZN(n3468) );
  INV_X1 U2789 ( .A(n2260), .ZN(n2261) );
  INV_X1 U2790 ( .A(n3427), .ZN(n3422) );
  INV_X1 U2791 ( .A(n3315), .ZN(n3855) );
  INV_X1 U2792 ( .A(n4117), .ZN(n4064) );
  INV_X1 U2793 ( .A(n4067), .ZN(n4115) );
  CLKBUF_X1 U2794 ( .A(n4047), .Z(n4052) );
  AOI21_X1 U2795 ( .B1(n4458), .B2(n2778), .A(n2748), .ZN(n4068) );
  INV_X1 U2796 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4066) );
  NOR2_X1 U2797 ( .A1(n2285), .A2(n2458), .ZN(n4061) );
  INV_X1 U2798 ( .A(n2288), .ZN(n2285) );
  NAND2_X1 U2799 ( .A1(n2457), .A2(n3928), .ZN(n2455) );
  NAND2_X1 U2800 ( .A1(n2199), .A2(n2200), .ZN(n4090) );
  OR2_X1 U2801 ( .A1(n3780), .A2(n3781), .ZN(n2200) );
  NAND2_X1 U2802 ( .A1(n2440), .A2(n2441), .ZN(n3484) );
  NAND2_X1 U2803 ( .A1(n4020), .A2(n2443), .ZN(n2440) );
  INV_X1 U2804 ( .A(n2444), .ZN(n2443) );
  NAND2_X1 U2805 ( .A1(n3342), .A2(n4643), .ZN(n4117) );
  NAND2_X1 U2806 ( .A1(n2276), .A2(n2275), .ZN(n4098) );
  NAND2_X1 U2807 ( .A1(n2278), .A2(n2274), .ZN(n2275) );
  NAND2_X1 U2808 ( .A1(n3346), .A2(n3330), .ZN(n4108) );
  INV_X1 U2809 ( .A(n4108), .ZN(n4122) );
  INV_X1 U2810 ( .A(n4487), .ZN(n4452) );
  OR2_X1 U2811 ( .A1(n4490), .A2(n2832), .ZN(n2502) );
  NAND2_X1 U2812 ( .A1(n2509), .A2(n2508), .ZN(n4484) );
  NAND2_X1 U2813 ( .A1(n2738), .A2(n2737), .ZN(n4545) );
  OAI21_X1 U2814 ( .B1(n4555), .B2(n2832), .A(n2724), .ZN(n4564) );
  INV_X1 U2815 ( .A(n4584), .ZN(n4091) );
  INV_X1 U2816 ( .A(n4609), .ZN(n4277) );
  NAND2_X1 U2817 ( .A1(n2778), .A2(n3508), .ZN(n2578) );
  NAND4_X1 U2818 ( .A1(n2557), .A2(n2556), .A3(n2555), .A4(n2554), .ZN(n3578)
         );
  NAND2_X1 U2819 ( .A1(n2778), .A2(REG3_REG_2__SCAN_IN), .ZN(n2513) );
  OR2_X1 U2820 ( .A1(n3369), .A2(n2885), .ZN(n4285) );
  XNOR2_X1 U2821 ( .A(n3175), .B(REG1_REG_1__SCAN_IN), .ZN(n3267) );
  NAND2_X1 U2822 ( .A1(n2295), .A2(n3177), .ZN(n4294) );
  AND2_X1 U2823 ( .A1(n3191), .A2(n3197), .ZN(n2229) );
  NAND2_X1 U2824 ( .A1(n3217), .A2(n3216), .ZN(n3221) );
  NAND2_X1 U2825 ( .A1(n2221), .A2(n3436), .ZN(n2220) );
  INV_X1 U2826 ( .A(n3445), .ZN(n2221) );
  OR2_X1 U2827 ( .A1(n3447), .A2(n4799), .ZN(n2344) );
  INV_X1 U2828 ( .A(n3522), .ZN(n2343) );
  NAND2_X1 U2829 ( .A1(n2341), .A2(n2339), .ZN(n3672) );
  AND2_X1 U2830 ( .A1(n4328), .A2(n4327), .ZN(n2216) );
  INV_X1 U2831 ( .A(n2338), .ZN(n4905) );
  INV_X1 U2832 ( .A(n2336), .ZN(n4903) );
  INV_X1 U2833 ( .A(n4939), .ZN(n2219) );
  AND2_X1 U2834 ( .A1(n3225), .A2(n4270), .ZN(n4948) );
  AOI21_X1 U2835 ( .B1(n2391), .B2(n2393), .A(n4204), .ZN(n2388) );
  NAND2_X1 U2836 ( .A1(n4711), .A2(n2182), .ZN(n4378) );
  NAND2_X1 U2837 ( .A1(n4463), .A2(n2358), .ZN(n4447) );
  NAND2_X1 U2838 ( .A1(n2361), .A2(n2365), .ZN(n4509) );
  NAND2_X1 U2839 ( .A1(n4548), .A2(n2159), .ZN(n2361) );
  NAND2_X1 U2840 ( .A1(n2378), .A2(n2381), .ZN(n4568) );
  NAND2_X1 U2841 ( .A1(n2385), .A2(n2382), .ZN(n2378) );
  INV_X1 U2842 ( .A(n4763), .ZN(n4594) );
  NAND2_X1 U2843 ( .A1(n2400), .A2(n2401), .ZN(n4607) );
  AND2_X1 U2844 ( .A1(n2373), .A2(n2609), .ZN(n4671) );
  AND2_X1 U2845 ( .A1(n2608), .A2(n2157), .ZN(n2373) );
  NAND2_X1 U2846 ( .A1(n4957), .A2(n3575), .ZN(n4697) );
  NAND2_X1 U2847 ( .A1(n3544), .A2(n4136), .ZN(n3452) );
  INV_X1 U2848 ( .A(n4572), .ZN(n4693) );
  INV_X1 U2849 ( .A(n4619), .ZN(n4666) );
  INV_X1 U2850 ( .A(n4643), .ZN(n4953) );
  OR2_X1 U2851 ( .A1(n3405), .A2(n3404), .ZN(n3406) );
  INV_X1 U2852 ( .A(REG1_REG_10__SCAN_IN), .ZN(n4799) );
  NAND2_X1 U2853 ( .A1(n4711), .A2(n2204), .ZN(n4815) );
  INV_X1 U2854 ( .A(n2205), .ZN(n2204) );
  OAI21_X1 U2855 ( .B1(n4709), .B2(n5000), .A(n2311), .ZN(n2205) );
  INV_X1 U2856 ( .A(n2312), .ZN(n2311) );
  OAI21_X1 U2857 ( .B1(n3902), .B2(n5002), .A(n2838), .ZN(n2880) );
  NAND2_X1 U2858 ( .A1(n2213), .A2(n5007), .ZN(n2212) );
  INV_X1 U2859 ( .A(n4718), .ZN(n2213) );
  AOI21_X1 U2860 ( .B1(n4721), .B2(n5007), .A(n2255), .ZN(n2254) );
  NOR2_X1 U2861 ( .A1(n4795), .A2(n4720), .ZN(n2255) );
  INV_X1 U2862 ( .A(n3407), .ZN(n2874) );
  NAND2_X1 U2863 ( .A1(n3326), .A2(n3338), .ZN(n4975) );
  AND2_X1 U2864 ( .A1(n2476), .A2(n2162), .ZN(n2462) );
  NAND2_X1 U2865 ( .A1(n2414), .A2(IR_REG_31__SCAN_IN), .ZN(n2895) );
  INV_X1 U2866 ( .A(n2868), .ZN(n4880) );
  INV_X1 U2867 ( .A(n4334), .ZN(n4980) );
  INV_X1 U2868 ( .A(IR_REG_16__SCAN_IN), .ZN(n2698) );
  XNOR2_X1 U2869 ( .A(n2650), .B(n2649), .ZN(n3671) );
  NAND2_X1 U2870 ( .A1(n2298), .A2(n2153), .ZN(n2320) );
  OAI21_X1 U2871 ( .B1(n4817), .B2(n5017), .A(n2251), .ZN(U3544) );
  AND2_X1 U2872 ( .A1(n2253), .A2(n2252), .ZN(n2251) );
  OR2_X1 U2873 ( .A1(n5019), .A2(n4722), .ZN(n2252) );
  OR2_X1 U2874 ( .A1(n4820), .A2(n4801), .ZN(n2253) );
  AND2_X1 U2875 ( .A1(n2457), .A2(n2449), .ZN(n2448) );
  INV_X1 U2876 ( .A(n2448), .ZN(n2267) );
  INV_X1 U2877 ( .A(n3582), .ZN(n2306) );
  AND2_X1 U2878 ( .A1(n3634), .A2(n2309), .ZN(n2145) );
  OR2_X1 U2879 ( .A1(n4545), .A2(n4527), .ZN(n2146) );
  AND2_X1 U2880 ( .A1(n3754), .A2(n3753), .ZN(n2147) );
  AND2_X1 U2881 ( .A1(n2401), .A2(n2399), .ZN(n2148) );
  NAND2_X1 U2882 ( .A1(n2175), .A2(n2386), .ZN(n2149) );
  NAND2_X1 U2883 ( .A1(n3807), .A2(n3806), .ZN(n2459) );
  AND2_X1 U2884 ( .A1(n2316), .A2(n4552), .ZN(n2150) );
  NAND2_X1 U2885 ( .A1(n2307), .A2(n2195), .ZN(n2151) );
  XNOR2_X1 U2886 ( .A(n3841), .B(n3756), .ZN(n2152) );
  AND2_X1 U2887 ( .A1(n4948), .A2(n2198), .ZN(n2153) );
  AND2_X1 U2888 ( .A1(n4935), .A2(n2192), .ZN(n2154) );
  NOR2_X1 U2889 ( .A1(n4944), .A2(n2196), .ZN(n2155) );
  OR2_X1 U2890 ( .A1(n2776), .A2(n3079), .ZN(n2156) );
  INV_X1 U2891 ( .A(n3737), .ZN(n3755) );
  OR2_X1 U2892 ( .A1(n4681), .A2(n3628), .ZN(n2157) );
  NAND4_X1 U2893 ( .A1(n2538), .A2(n2537), .A3(n2536), .A4(n2535), .ZN(n3313)
         );
  NAND2_X1 U2894 ( .A1(n2834), .A2(IR_REG_27__SCAN_IN), .ZN(n2158) );
  AND2_X1 U2895 ( .A1(n2146), .A2(n2730), .ZN(n2159) );
  INV_X1 U2896 ( .A(n4204), .ZN(n4356) );
  AND2_X1 U2897 ( .A1(n4362), .A2(n4364), .ZN(n4204) );
  OR2_X1 U2898 ( .A1(n4400), .A2(n4714), .ZN(n2160) );
  INV_X1 U2899 ( .A(IR_REG_31__SCAN_IN), .ZN(n2416) );
  AND2_X1 U2900 ( .A1(n4545), .A2(n4527), .ZN(n2161) );
  NOR2_X1 U2901 ( .A1(IR_REG_27__SCAN_IN), .A2(IR_REG_26__SCAN_IN), .ZN(n2162)
         );
  OR2_X1 U2902 ( .A1(n3262), .A2(n3129), .ZN(n2163) );
  AND3_X1 U2903 ( .A1(n3775), .A2(n3774), .A3(n3776), .ZN(n2164) );
  INV_X1 U2904 ( .A(n2376), .ZN(n2375) );
  OAI22_X1 U2905 ( .A1(n2157), .A2(n2620), .B1(n4280), .B2(n4688), .ZN(n2376)
         );
  NAND2_X1 U2906 ( .A1(n4198), .A2(n2820), .ZN(n2165) );
  NAND2_X1 U2907 ( .A1(n2389), .A2(n2388), .ZN(n4713) );
  AND2_X1 U2908 ( .A1(n4584), .A2(n4561), .ZN(n2166) );
  INV_X1 U2909 ( .A(n3483), .ZN(n2445) );
  OR2_X1 U2910 ( .A1(n3300), .A2(REG1_REG_7__SCAN_IN), .ZN(n2167) );
  INV_X1 U2911 ( .A(REG3_REG_9__SCAN_IN), .ZN(n2610) );
  INV_X1 U2912 ( .A(n2358), .ZN(n2356) );
  OR2_X1 U2913 ( .A1(n4487), .A2(n4465), .ZN(n2358) );
  NOR2_X1 U2914 ( .A1(n4391), .A2(n2207), .ZN(n2168) );
  INV_X1 U2915 ( .A(n2398), .ZN(n2397) );
  NOR2_X1 U2916 ( .A1(n4438), .A2(n4421), .ZN(n2398) );
  INV_X1 U2917 ( .A(IR_REG_21__SCAN_IN), .ZN(n3096) );
  INV_X1 U2918 ( .A(n2287), .ZN(n2286) );
  NAND2_X1 U2919 ( .A1(n4062), .A2(n2459), .ZN(n2287) );
  NOR2_X1 U2920 ( .A1(n4530), .A2(n4512), .ZN(n2366) );
  AND2_X1 U2921 ( .A1(n3741), .A2(n2456), .ZN(n2169) );
  AND3_X1 U2922 ( .A1(n3888), .A2(n3889), .A3(n4122), .ZN(n2170) );
  AND2_X1 U2923 ( .A1(n2444), .A2(n2445), .ZN(n2171) );
  AND2_X1 U2924 ( .A1(n2306), .A2(n2798), .ZN(n2172) );
  INV_X1 U2925 ( .A(n2620), .ZN(n2374) );
  OR2_X1 U2926 ( .A1(n3887), .A2(n4384), .ZN(n2173) );
  AND3_X1 U2927 ( .A1(n2739), .A2(n2740), .A3(n2741), .ZN(n2174) );
  NOR2_X1 U2928 ( .A1(n4595), .A2(n2704), .ZN(n2175) );
  AND2_X1 U2929 ( .A1(n2843), .A2(n2867), .ZN(n2176) );
  INV_X1 U2930 ( .A(n2396), .ZN(n2395) );
  NOR2_X1 U2931 ( .A1(n2764), .A2(n2398), .ZN(n2396) );
  AND2_X1 U2932 ( .A1(n2419), .A2(n4245), .ZN(n2177) );
  AND2_X1 U2933 ( .A1(n2145), .A2(n4794), .ZN(n2178) );
  AND2_X1 U2934 ( .A1(n2172), .A2(n2308), .ZN(n2179) );
  NAND2_X1 U2935 ( .A1(n2149), .A2(n2705), .ZN(n2381) );
  AND2_X1 U2936 ( .A1(n3096), .A2(n2840), .ZN(n2180) );
  INV_X1 U2937 ( .A(IR_REG_28__SCAN_IN), .ZN(n2834) );
  AND2_X1 U2938 ( .A1(n2278), .A2(n4099), .ZN(n2277) );
  OR2_X1 U2939 ( .A1(n2267), .A2(n3960), .ZN(n2181) );
  INV_X1 U2940 ( .A(n4626), .ZN(n2385) );
  INV_X1 U2941 ( .A(n4720), .ZN(n2207) );
  INV_X1 U2942 ( .A(n4244), .ZN(n2425) );
  INV_X1 U2943 ( .A(n4216), .ZN(n2426) );
  NAND2_X1 U2944 ( .A1(n4548), .A2(n2730), .ZN(n4531) );
  NAND2_X1 U2945 ( .A1(n2454), .A2(n2455), .ZN(n4073) );
  INV_X1 U2946 ( .A(n3973), .ZN(n2274) );
  INV_X1 U2947 ( .A(n4160), .ZN(n2248) );
  OR2_X1 U2948 ( .A1(n2156), .A2(n4643), .ZN(n2182) );
  INV_X1 U2949 ( .A(n4552), .ZN(n4092) );
  AND2_X1 U2950 ( .A1(n4588), .A2(n2150), .ZN(n2183) );
  OR2_X1 U2951 ( .A1(n4306), .A2(n3446), .ZN(n2184) );
  INV_X1 U2952 ( .A(n2459), .ZN(n2458) );
  INV_X1 U2953 ( .A(n4561), .ZN(n4569) );
  AND2_X1 U2954 ( .A1(n2150), .A2(n4535), .ZN(n2185) );
  AND2_X1 U2955 ( .A1(n2344), .A2(n2343), .ZN(n2186) );
  NAND2_X1 U2956 ( .A1(n3673), .A2(REG1_REG_11__SCAN_IN), .ZN(n2187) );
  XNOR2_X1 U2957 ( .A(n2699), .B(n2698), .ZN(n4983) );
  AND2_X2 U2958 ( .A1(n2879), .A2(n3407), .ZN(n5019) );
  AND2_X2 U2959 ( .A1(n2874), .A2(n2879), .ZN(n5013) );
  OR2_X1 U2960 ( .A1(n2260), .A2(n2442), .ZN(n2441) );
  NOR2_X1 U2961 ( .A1(n2334), .A2(n4322), .ZN(n2188) );
  INV_X1 U2962 ( .A(n4615), .ZN(n2399) );
  NAND2_X1 U2963 ( .A1(n2431), .A2(n2433), .ZN(n3357) );
  AND2_X1 U2964 ( .A1(n3574), .A2(n4989), .ZN(n5002) );
  INV_X1 U2965 ( .A(n5002), .ZN(n5007) );
  NOR2_X1 U2966 ( .A1(n3473), .A2(n3472), .ZN(n2189) );
  NAND2_X1 U2967 ( .A1(n2789), .A2(n2462), .ZN(n2833) );
  OR2_X1 U2968 ( .A1(n3696), .A2(n4782), .ZN(n2190) );
  AND2_X1 U2969 ( .A1(n4330), .A2(REG2_REG_15__SCAN_IN), .ZN(n2191) );
  INV_X1 U2970 ( .A(n2147), .ZN(n2449) );
  OR2_X1 U2971 ( .A1(n2324), .A2(n2188), .ZN(n2192) );
  OR2_X1 U2972 ( .A1(n4340), .A2(n2326), .ZN(n2193) );
  AND2_X1 U2973 ( .A1(n2310), .A2(n4421), .ZN(n2194) );
  AND2_X1 U2974 ( .A1(n2308), .A2(n2306), .ZN(n2195) );
  NOR2_X1 U2975 ( .A1(n4949), .A2(n4980), .ZN(n2196) );
  INV_X1 U2976 ( .A(n2222), .ZN(n2303) );
  INV_X1 U2977 ( .A(IR_REG_30__SCAN_IN), .ZN(n3867) );
  INV_X1 U2978 ( .A(IR_REG_20__SCAN_IN), .ZN(n2924) );
  AND2_X1 U2979 ( .A1(n3176), .A2(n3177), .ZN(n2197) );
  NOR2_X1 U2980 ( .A1(n2333), .A2(n2328), .ZN(n2198) );
  XNOR2_X1 U2981 ( .A(n4940), .B(n2219), .ZN(n2218) );
  NAND3_X1 U2982 ( .A1(n3985), .A2(n3984), .A3(n2164), .ZN(n2199) );
  NAND2_X1 U2983 ( .A1(n2201), .A2(n2181), .ZN(n2263) );
  NOR2_X2 U2984 ( .A1(n2452), .A2(n2451), .ZN(n2450) );
  INV_X1 U2985 ( .A(n2266), .ZN(n2201) );
  AOI21_X2 U2986 ( .B1(n2450), .B2(n2267), .A(n2152), .ZN(n2266) );
  NOR2_X1 U2987 ( .A1(n2454), .A2(n2147), .ZN(n2452) );
  AOI21_X1 U2988 ( .B1(n3907), .B2(n3903), .A(n3904), .ZN(n3764) );
  NAND3_X1 U2989 ( .A1(n2202), .A2(n2296), .A3(n2155), .ZN(U3258) );
  NAND2_X1 U2990 ( .A1(n2218), .A2(n4935), .ZN(n2202) );
  NAND2_X1 U2991 ( .A1(n2228), .A2(n2203), .ZN(n4299) );
  NAND2_X1 U2992 ( .A1(n4580), .A2(n4600), .ZN(n4586) );
  NAND2_X1 U2993 ( .A1(n2420), .A2(n2177), .ZN(n2258) );
  NOR2_X1 U2994 ( .A1(n2803), .A2(n4652), .ZN(n2808) );
  OAI21_X2 U2995 ( .B1(n4501), .B2(n4172), .A(n4175), .ZN(n4481) );
  NAND2_X1 U2996 ( .A1(n3366), .A2(n3367), .ZN(n4019) );
  AOI21_X1 U2997 ( .B1(n3356), .B2(n2433), .A(n2432), .ZN(n3718) );
  INV_X4 U2998 ( .A(n3737), .ZN(n3760) );
  OAI211_X1 U2999 ( .C1(n3884), .C2(n3893), .A(n2210), .B(n3892), .ZN(U3217)
         );
  NAND2_X1 U3000 ( .A1(n3884), .A2(n2170), .ZN(n2210) );
  AND2_X4 U3001 ( .A1(n3826), .A2(n5000), .ZN(n3420) );
  NAND3_X1 U3002 ( .A1(n4717), .A2(n4716), .A3(n2212), .ZN(n4816) );
  OAI211_X1 U3003 ( .C1(n2315), .C2(n2465), .A(n2313), .B(n4710), .ZN(n2312)
         );
  INV_X1 U3004 ( .A(n4713), .ZN(n2315) );
  OAI21_X2 U3005 ( .B1(n4435), .B2(n4415), .A(n2750), .ZN(n4410) );
  NAND2_X1 U3006 ( .A1(n4410), .A2(n2391), .ZN(n2389) );
  AOI21_X1 U3007 ( .B1(n4466), .B2(n4492), .A(n2742), .ZN(n4464) );
  NAND2_X1 U3008 ( .A1(n4298), .A2(n4299), .ZN(n4297) );
  NAND2_X1 U3009 ( .A1(n4945), .A2(n2226), .ZN(n2215) );
  NAND2_X1 U3010 ( .A1(n2262), .A2(n2264), .ZN(n4047) );
  NAND2_X1 U3011 ( .A1(n4037), .A2(n4038), .ZN(n4036) );
  XNOR2_X2 U3012 ( .A(n3437), .B(n3444), .ZN(n3435) );
  NAND3_X1 U3013 ( .A1(n2215), .A2(n2320), .A3(n2214), .ZN(U3259) );
  INV_X1 U3014 ( .A(n2516), .ZN(n2224) );
  NOR2_X2 U3015 ( .A1(n4326), .A2(n2216), .ZN(n4909) );
  NOR2_X2 U3016 ( .A1(n3706), .A2(n3707), .ZN(n4326) );
  AOI21_X2 U3017 ( .B1(n4090), .B2(n4086), .A(n4088), .ZN(n3943) );
  NAND2_X2 U3018 ( .A1(n4918), .A2(n4917), .ZN(n4916) );
  NAND2_X1 U3019 ( .A1(n3267), .A2(n3268), .ZN(n3172) );
  NAND2_X1 U3020 ( .A1(n3881), .A2(n3880), .ZN(n3884) );
  INV_X1 U3021 ( .A(n2411), .ZN(n2409) );
  XNOR2_X2 U3022 ( .A(n3215), .B(n3204), .ZN(n3214) );
  XNOR2_X2 U3023 ( .A(n3527), .B(n3442), .ZN(n3525) );
  NOR2_X2 U3024 ( .A1(n4909), .A2(n4910), .ZN(n4908) );
  INV_X1 U3025 ( .A(n2298), .ZN(n4945) );
  NOR2_X2 U3026 ( .A1(n2787), .A2(n2257), .ZN(n2476) );
  NAND4_X1 U3027 ( .A1(n2348), .A2(n2347), .A3(n2345), .A4(n2346), .ZN(n2787)
         );
  NAND2_X1 U3028 ( .A1(n2789), .A2(n2174), .ZN(n2225) );
  NAND2_X1 U3029 ( .A1(n2271), .A2(n2277), .ZN(n3881) );
  AOI22_X1 U3030 ( .A1(n3755), .A2(n3322), .B1(n3826), .B2(n3321), .ZN(n3320)
         );
  NAND2_X1 U3031 ( .A1(n2436), .A2(n2434), .ZN(n2433) );
  NAND2_X2 U3032 ( .A1(n4309), .A2(n3440), .ZN(n3527) );
  NAND2_X2 U3033 ( .A1(n3237), .A2(n3202), .ZN(n3215) );
  NAND2_X2 U3034 ( .A1(n3296), .A2(n3295), .ZN(n3437) );
  NAND2_X1 U3035 ( .A1(n4930), .A2(n2230), .ZN(n4946) );
  NAND2_X1 U3036 ( .A1(n2294), .A2(n4293), .ZN(n2292) );
  AND2_X2 U3037 ( .A1(n4036), .A2(n4040), .ZN(n2461) );
  NAND2_X1 U3038 ( .A1(n2263), .A2(n3748), .ZN(n2262) );
  NAND2_X1 U3039 ( .A1(n3972), .A2(n3973), .ZN(n2271) );
  OR2_X1 U3040 ( .A1(n4333), .A2(REG1_REG_17__SCAN_IN), .ZN(n2227) );
  AOI21_X2 U3041 ( .B1(n4890), .B2(REG1_REG_4__SCAN_IN), .A(n2229), .ZN(n3236)
         );
  NOR2_X2 U3042 ( .A1(n2571), .A2(n2563), .ZN(n2595) );
  NAND3_X1 U3043 ( .A1(n4230), .A2(n4228), .A3(n4488), .ZN(n2235) );
  NAND3_X1 U3044 ( .A1(n2350), .A2(n2349), .A3(n2476), .ZN(n2256) );
  NAND4_X1 U3045 ( .A1(n2475), .A2(n3096), .A3(n2843), .A4(n2867), .ZN(n2257)
         );
  XNOR2_X1 U3046 ( .A(n3468), .B(n2261), .ZN(n3433) );
  AOI21_X1 U3047 ( .B1(n2450), .B2(n2152), .A(n3960), .ZN(n2265) );
  NAND3_X1 U3048 ( .A1(n3825), .A2(n4009), .A3(n2277), .ZN(n2270) );
  NAND2_X1 U3049 ( .A1(n3825), .A2(n4009), .ZN(n3972) );
  NAND2_X1 U3050 ( .A1(n2270), .A2(n2272), .ZN(n3843) );
  NAND3_X1 U3051 ( .A1(n3825), .A2(n4009), .A3(n2278), .ZN(n2276) );
  INV_X1 U3052 ( .A(n3974), .ZN(n2278) );
  NAND2_X1 U3053 ( .A1(n2461), .A2(n2280), .ZN(n2279) );
  NAND2_X2 U3054 ( .A1(n2288), .A2(n2286), .ZN(n4060) );
  NAND2_X1 U3055 ( .A1(n2289), .A2(n2789), .ZN(n2290) );
  NAND2_X1 U3056 ( .A1(n2789), .A2(n2291), .ZN(n2844) );
  NAND2_X1 U3057 ( .A1(n2789), .A2(n2788), .ZN(n2839) );
  INV_X1 U3058 ( .A(n3176), .ZN(n2295) );
  NAND2_X1 U3059 ( .A1(n3176), .A2(n4293), .ZN(n2293) );
  INV_X1 U3060 ( .A(n3177), .ZN(n2294) );
  OAI21_X2 U3061 ( .B1(n3702), .B2(n3701), .A(n3703), .ZN(n4325) );
  NAND2_X2 U3062 ( .A1(n3682), .A2(n3681), .ZN(n3702) );
  NOR2_X2 U3063 ( .A1(n4908), .A2(n2191), .ZN(n4331) );
  NAND3_X1 U3064 ( .A1(n2298), .A2(n4948), .A3(n2297), .ZN(n2296) );
  NAND2_X1 U3065 ( .A1(n4946), .A2(n4947), .ZN(n2297) );
  OR2_X2 U3066 ( .A1(n4946), .A2(n4947), .ZN(n2298) );
  INV_X1 U3067 ( .A(n3552), .ZN(n2307) );
  NAND2_X1 U3068 ( .A1(n2307), .A2(n2179), .ZN(n3598) );
  XNOR2_X2 U3069 ( .A(n2317), .B(n2527), .ZN(n3175) );
  AND2_X1 U3070 ( .A1(n4334), .A2(REG1_REG_18__SCAN_IN), .ZN(n2334) );
  XNOR2_X2 U3071 ( .A(n4320), .B(n2700), .ZN(n4918) );
  AND2_X2 U3072 ( .A1(n2336), .A2(n2335), .ZN(n4320) );
  AND3_X2 U3073 ( .A1(n2341), .A2(n2339), .A3(n2187), .ZN(n3686) );
  OR2_X2 U3074 ( .A1(n3447), .A2(n2342), .ZN(n2341) );
  INV_X1 U3075 ( .A(n2344), .ZN(n3523) );
  NOR2_X4 U3076 ( .A1(n2591), .A2(n2474), .ZN(n2789) );
  XNOR2_X2 U3077 ( .A(n2518), .B(n2517), .ZN(n3174) );
  NAND2_X1 U3078 ( .A1(n3866), .A2(IR_REG_31__SCAN_IN), .ZN(n2479) );
  NAND4_X1 U3079 ( .A1(n2349), .A2(n2350), .A3(n2478), .A4(n2476), .ZN(n3866)
         );
  AND2_X2 U3080 ( .A1(n2463), .A2(n2351), .ZN(n2350) );
  OAI22_X1 U3081 ( .A1(n4464), .A2(n2353), .B1(n2354), .B2(n2352), .ZN(n4429)
         );
  NAND2_X1 U3082 ( .A1(n4429), .A2(n2468), .ZN(n2750) );
  NAND2_X1 U3083 ( .A1(n4548), .A2(n2362), .ZN(n2359) );
  NAND2_X1 U3084 ( .A1(n2359), .A2(n2360), .ZN(n4489) );
  INV_X1 U3085 ( .A(n2608), .ZN(n2368) );
  NAND3_X1 U3086 ( .A1(n2372), .A2(n2371), .A3(n2370), .ZN(n2633) );
  NAND2_X1 U3087 ( .A1(n2368), .A2(n2374), .ZN(n2370) );
  NAND2_X1 U3088 ( .A1(n2369), .A2(n2374), .ZN(n2372) );
  INV_X1 U3089 ( .A(n2609), .ZN(n2369) );
  NAND3_X1 U3090 ( .A1(n2372), .A2(n2375), .A3(n2370), .ZN(n4651) );
  NAND2_X1 U3091 ( .A1(n4625), .A2(n2381), .ZN(n2377) );
  INV_X1 U3092 ( .A(n2667), .ZN(n2387) );
  OAI21_X1 U3093 ( .B1(n4410), .B2(n2757), .A(n2397), .ZN(n4403) );
  NAND2_X1 U3094 ( .A1(n4410), .A2(n2396), .ZN(n2390) );
  NAND3_X1 U3095 ( .A1(n2394), .A2(n2395), .A3(n2160), .ZN(n2392) );
  NAND2_X1 U3096 ( .A1(n2417), .A2(n2789), .ZN(n2414) );
  NAND2_X1 U3097 ( .A1(n2789), .A2(n2476), .ZN(n2848) );
  NAND2_X1 U3098 ( .A1(n4481), .A2(n2421), .ZN(n2420) );
  NAND2_X1 U3099 ( .A1(n2428), .A2(n2799), .ZN(n3643) );
  INV_X1 U3100 ( .A(n2435), .ZN(n2434) );
  XNOR2_X1 U3101 ( .A(n3320), .B(n3841), .ZN(n2435) );
  AND2_X1 U3102 ( .A1(n2435), .A2(n3355), .ZN(n2432) );
  OR2_X1 U3103 ( .A1(n3426), .A2(n3427), .ZN(n2447) );
  AND2_X1 U3104 ( .A1(n3313), .A2(n3315), .ZN(n3283) );
  NAND2_X1 U3105 ( .A1(n2880), .A2(n5013), .ZN(n2878) );
  AOI22_X2 U3106 ( .A1(n3211), .A2(REG1_REG_6__SCAN_IN), .B1(n4885), .B2(n3210), .ZN(n3297) );
  NAND2_X1 U3107 ( .A1(n2511), .A2(REG1_REG_2__SCAN_IN), .ZN(n2512) );
  INV_X1 U3108 ( .A(n2533), .ZN(n2542) );
  AND2_X1 U3109 ( .A1(n2144), .A2(DATAI_28_), .ZN(n3895) );
  NAND2_X1 U3110 ( .A1(n2144), .A2(n2519), .ZN(n2520) );
  AND2_X1 U3111 ( .A1(n2144), .A2(DATAI_21_), .ZN(n4483) );
  AND2_X1 U3112 ( .A1(n2144), .A2(DATAI_22_), .ZN(n4476) );
  NAND2_X1 U3113 ( .A1(n4220), .A2(n2540), .ZN(n2541) );
  NAND2_X1 U3114 ( .A1(n2778), .A2(REG3_REG_1__SCAN_IN), .ZN(n2526) );
  AND2_X1 U3115 ( .A1(n2877), .A2(n2876), .ZN(n2464) );
  OR3_X1 U3116 ( .A1(n4705), .A2(n4704), .A3(n5002), .ZN(n2465) );
  AND2_X1 U3117 ( .A1(n4681), .A2(n3628), .ZN(n2466) );
  AND2_X1 U3118 ( .A1(n4632), .A2(n3965), .ZN(n2467) );
  INV_X1 U3119 ( .A(n3174), .ZN(n2521) );
  AND2_X1 U3120 ( .A1(n3167), .A2(n4287), .ZN(n4682) );
  NAND2_X1 U3121 ( .A1(n2825), .A2(n2824), .ZN(n4525) );
  INV_X1 U3122 ( .A(n4525), .ZN(n4684) );
  OR2_X1 U3123 ( .A1(n4455), .A2(n4440), .ZN(n2468) );
  INV_X1 U3124 ( .A(IR_REG_22__SCAN_IN), .ZN(n2840) );
  OR2_X1 U3125 ( .A1(n3259), .A2(n4818), .ZN(n2759) );
  INV_X1 U3126 ( .A(REG3_REG_17__SCAN_IN), .ZN(n2706) );
  NAND2_X1 U3127 ( .A1(n2143), .A2(n2528), .ZN(n2529) );
  INV_X1 U3128 ( .A(n4769), .ZN(n2875) );
  OR2_X1 U3129 ( .A1(n2714), .A2(IR_REG_14__SCAN_IN), .ZN(n2685) );
  AND2_X1 U3130 ( .A1(n3821), .A2(n3822), .ZN(n3819) );
  INV_X1 U3131 ( .A(REG3_REG_18__SCAN_IN), .ZN(n2717) );
  AND2_X1 U3132 ( .A1(n3201), .A2(REG1_REG_5__SCAN_IN), .ZN(n3192) );
  NAND2_X1 U3133 ( .A1(n4316), .A2(n4327), .ZN(n4317) );
  INV_X1 U3134 ( .A(n4774), .ZN(n3910) );
  NAND2_X1 U3135 ( .A1(n2542), .A2(n2541), .ZN(n3543) );
  INV_X1 U3136 ( .A(IR_REG_25__SCAN_IN), .ZN(n2845) );
  INV_X1 U3137 ( .A(REG3_REG_23__SCAN_IN), .ZN(n3920) );
  INV_X1 U3138 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3042) );
  INV_X1 U3139 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3079) );
  NAND2_X1 U3140 ( .A1(n2511), .A2(REG1_REG_0__SCAN_IN), .ZN(n2536) );
  AND2_X1 U3141 ( .A1(n3521), .A2(n3526), .ZN(n3522) );
  AOI21_X1 U3142 ( .B1(n4942), .B2(ADDR_REG_18__SCAN_IN), .A(n4941), .ZN(n4943) );
  AND2_X1 U3143 ( .A1(n4203), .A2(n4397), .ZN(n4412) );
  INV_X1 U3144 ( .A(n4505), .ZN(n4466) );
  AND2_X1 U3145 ( .A1(n4519), .A2(n4518), .ZN(n4567) );
  NAND2_X1 U3146 ( .A1(n2800), .A2(n4144), .ZN(n3610) );
  AND2_X1 U3147 ( .A1(n4130), .A2(n4134), .ZN(n4223) );
  AND2_X1 U31480 ( .A1(n2144), .A2(DATAI_25_), .ZN(n4414) );
  INV_X1 U31490 ( .A(n4682), .ZN(n4659) );
  OR2_X1 U3150 ( .A1(n4287), .A2(n3328), .ZN(n4678) );
  AND2_X1 U3151 ( .A1(n3346), .A2(n3345), .ZN(n4116) );
  INV_X1 U3152 ( .A(n4120), .ZN(n4102) );
  AND2_X1 U3153 ( .A1(n3407), .A2(n3327), .ZN(n3346) );
  INV_X1 U3154 ( .A(n4068), .ZN(n4473) );
  INV_X1 U3155 ( .A(n4943), .ZN(n4944) );
  AND2_X1 U3156 ( .A1(n3225), .A2(n4289), .ZN(n4935) );
  AND2_X1 U3157 ( .A1(n4185), .A2(n4182), .ZN(n4390) );
  AND2_X1 U3158 ( .A1(n2144), .A2(DATAI_20_), .ZN(n4745) );
  AND2_X1 U3159 ( .A1(n4209), .A2(n4208), .ZN(n4656) );
  INV_X1 U3160 ( .A(n4697), .ZN(n4577) );
  AND2_X1 U3161 ( .A1(n4139), .A2(n4151), .ZN(n4212) );
  INV_X1 U3162 ( .A(REG1_REG_13__SCAN_IN), .ZN(n4782) );
  AND2_X1 U3163 ( .A1(n2851), .A2(n3161), .ZN(n3407) );
  INV_X1 U3164 ( .A(n4414), .ZN(n4421) );
  INV_X1 U3165 ( .A(n3731), .ZN(n4794) );
  INV_X1 U3166 ( .A(n5000), .ZN(n4994) );
  INV_X1 U3167 ( .A(n3403), .ZN(n3338) );
  AND2_X1 U3168 ( .A1(n3183), .A2(n3182), .ZN(n4942) );
  AND2_X1 U3169 ( .A1(n3373), .A2(n3372), .ZN(n4120) );
  AND4_X1 U3170 ( .A1(n4106), .A2(n4105), .A3(n4104), .A4(n4103), .ZN(n4107)
         );
  OAI21_X1 U3171 ( .B1(n2156), .B2(n2832), .A(n2831), .ZN(n4276) );
  NAND2_X1 U3172 ( .A1(n2502), .A2(n2501), .ZN(n4505) );
  INV_X1 U3173 ( .A(n4948), .ZN(n3705) );
  INV_X1 U3174 ( .A(n4935), .ZN(n4938) );
  OR2_X1 U3175 ( .A1(n4554), .A2(n5000), .ZN(n4572) );
  INV_X1 U3176 ( .A(n2882), .ZN(n2883) );
  NAND2_X1 U3177 ( .A1(n5019), .A2(n4994), .ZN(n4801) );
  INV_X1 U3178 ( .A(n5019), .ZN(n5017) );
  NAND2_X1 U3179 ( .A1(n5013), .A2(n4994), .ZN(n4872) );
  INV_X1 U3180 ( .A(n5013), .ZN(n5012) );
  INV_X1 U3181 ( .A(n4975), .ZN(n4977) );
  INV_X1 U3182 ( .A(D_REG_0__SCAN_IN), .ZN(n3163) );
  AND2_X1 U3183 ( .A1(n3368), .A2(STATE_REG_SCAN_IN), .ZN(n4978) );
  INV_X1 U3184 ( .A(n4333), .ZN(n4981) );
  INV_X2 U3185 ( .A(n4285), .ZN(U4043) );
  NAND2_X1 U3186 ( .A1(n2878), .A2(n2464), .ZN(U3514) );
  NAND2_X1 U3187 ( .A1(n2516), .A2(n2517), .ZN(n2550) );
  NAND2_X1 U3188 ( .A1(n2558), .A2(n2561), .ZN(n2469) );
  OR2_X2 U3189 ( .A1(n2550), .A2(n2469), .ZN(n2591) );
  NOR2_X1 U3190 ( .A1(IR_REG_22__SCAN_IN), .A2(IR_REG_25__SCAN_IN), .ZN(n2475)
         );
  INV_X2 U3191 ( .A(IR_REG_24__SCAN_IN), .ZN(n2843) );
  NAND2_X1 U3192 ( .A1(n2144), .A2(DATAI_24_), .ZN(n4440) );
  NAND2_X1 U3193 ( .A1(n2583), .A2(REG3_REG_6__SCAN_IN), .ZN(n2571) );
  NAND2_X1 U3194 ( .A1(n2595), .A2(REG3_REG_8__SCAN_IN), .ZN(n2611) );
  NAND2_X1 U3195 ( .A1(n2634), .A2(REG3_REG_11__SCAN_IN), .ZN(n2660) );
  OR2_X2 U3196 ( .A1(n2707), .A2(n2706), .ZN(n2718) );
  NOR2_X2 U3197 ( .A1(n2718), .A2(n2717), .ZN(n2731) );
  OR2_X2 U3198 ( .A1(n2504), .A2(n3954), .ZN(n2497) );
  OR2_X2 U3199 ( .A1(n2497), .A2(n4066), .ZN(n2743) );
  AND2_X2 U3200 ( .A1(n2744), .A2(REG3_REG_24__SCAN_IN), .ZN(n2751) );
  NOR2_X1 U3201 ( .A1(n2744), .A2(REG3_REG_24__SCAN_IN), .ZN(n2477) );
  NOR2_X1 U3202 ( .A1(n2751), .A2(n2477), .ZN(n4442) );
  XNOR2_X2 U3203 ( .A(n2479), .B(n3867), .ZN(n2481) );
  XNOR2_X2 U3204 ( .A(n2480), .B(IR_REG_29__SCAN_IN), .ZN(n2903) );
  NAND2_X1 U3205 ( .A1(n4442), .A2(n2778), .ZN(n2487) );
  NAND2_X4 U3206 ( .A1(n2481), .A2(n2903), .ZN(n3262) );
  INV_X1 U3207 ( .A(REG1_REG_24__SCAN_IN), .ZN(n4729) );
  NAND2_X1 U3208 ( .A1(n2572), .A2(REG2_REG_24__SCAN_IN), .ZN(n2484) );
  NAND2_X4 U3209 ( .A1(n2482), .A2(n2481), .ZN(n3259) );
  INV_X1 U32100 ( .A(REG0_REG_24__SCAN_IN), .ZN(n4826) );
  OR2_X1 U32110 ( .A1(n3259), .A2(n4826), .ZN(n2483) );
  OAI211_X1 U32120 ( .C1(n3262), .C2(n4729), .A(n2484), .B(n2483), .ZN(n2485)
         );
  INV_X1 U32130 ( .A(n2485), .ZN(n2486) );
  NAND2_X1 U32140 ( .A1(n2497), .A2(n4066), .ZN(n2488) );
  AND2_X1 U32150 ( .A1(n2743), .A2(n2488), .ZN(n4474) );
  NAND2_X1 U32160 ( .A1(n4474), .A2(n2778), .ZN(n2495) );
  INV_X1 U32170 ( .A(REG1_REG_22__SCAN_IN), .ZN(n2492) );
  NAND2_X1 U32180 ( .A1(n2572), .A2(REG2_REG_22__SCAN_IN), .ZN(n2491) );
  INV_X1 U32190 ( .A(REG0_REG_22__SCAN_IN), .ZN(n2489) );
  OR2_X1 U32200 ( .A1(n3259), .A2(n2489), .ZN(n2490) );
  OAI211_X1 U32210 ( .C1(n3262), .C2(n2492), .A(n2491), .B(n2490), .ZN(n2493)
         );
  INV_X1 U32220 ( .A(n2493), .ZN(n2494) );
  NAND2_X1 U32230 ( .A1(n2504), .A2(n3954), .ZN(n2496) );
  NAND2_X1 U32240 ( .A1(n2497), .A2(n2496), .ZN(n4490) );
  INV_X1 U32250 ( .A(REG1_REG_21__SCAN_IN), .ZN(n4742) );
  NAND2_X1 U32260 ( .A1(n2572), .A2(REG2_REG_21__SCAN_IN), .ZN(n2499) );
  INV_X1 U32270 ( .A(REG0_REG_21__SCAN_IN), .ZN(n4835) );
  OR2_X1 U32280 ( .A1(n3259), .A2(n4835), .ZN(n2498) );
  OAI211_X1 U32290 ( .C1(n3262), .C2(n4742), .A(n2499), .B(n2498), .ZN(n2500)
         );
  INV_X1 U32300 ( .A(n2500), .ZN(n2501) );
  INV_X1 U32310 ( .A(n4483), .ZN(n4492) );
  OR2_X1 U32320 ( .A1(n2733), .A2(REG3_REG_20__SCAN_IN), .ZN(n2503) );
  NAND2_X1 U32330 ( .A1(n2504), .A2(n2503), .ZN(n4510) );
  OR2_X1 U32340 ( .A1(n4510), .A2(n2832), .ZN(n2509) );
  INV_X1 U32350 ( .A(REG1_REG_20__SCAN_IN), .ZN(n4750) );
  NAND2_X1 U32360 ( .A1(n2572), .A2(REG2_REG_20__SCAN_IN), .ZN(n2506) );
  INV_X1 U32370 ( .A(REG0_REG_20__SCAN_IN), .ZN(n4839) );
  OR2_X1 U32380 ( .A1(n3259), .A2(n4839), .ZN(n2505) );
  OAI211_X1 U32390 ( .C1(n3262), .C2(n4750), .A(n2506), .B(n2505), .ZN(n2507)
         );
  INV_X1 U32400 ( .A(n2507), .ZN(n2508) );
  INV_X1 U32410 ( .A(n4484), .ZN(n4530) );
  INV_X1 U32420 ( .A(REG0_REG_2__SCAN_IN), .ZN(n2510) );
  OR2_X1 U32430 ( .A1(n3259), .A2(n2510), .ZN(n2515) );
  NAND2_X1 U32440 ( .A1(n2572), .A2(REG2_REG_2__SCAN_IN), .ZN(n2514) );
  INV_X1 U32450 ( .A(DATAI_2_), .ZN(n2519) );
  INV_X1 U32460 ( .A(n2539), .ZN(n2532) );
  INV_X1 U32470 ( .A(REG0_REG_1__SCAN_IN), .ZN(n2522) );
  OR2_X1 U32480 ( .A1(n3259), .A2(n2522), .ZN(n2525) );
  NAND2_X1 U32490 ( .A1(n2511), .A2(REG1_REG_1__SCAN_IN), .ZN(n2524) );
  NAND2_X1 U32500 ( .A1(n2572), .A2(REG2_REG_1__SCAN_IN), .ZN(n2523) );
  NAND4_X2 U32510 ( .A1(n2526), .A2(n2525), .A3(n2524), .A4(n2523), .ZN(n3322)
         );
  INV_X1 U32520 ( .A(IR_REG_1__SCAN_IN), .ZN(n2527) );
  INV_X1 U32530 ( .A(n3175), .ZN(n3170) );
  INV_X1 U32540 ( .A(n3170), .ZN(n3276) );
  NAND2_X1 U32550 ( .A1(n2653), .A2(n3276), .ZN(n2530) );
  INV_X1 U32560 ( .A(DATAI_1_), .ZN(n2528) );
  NAND2_X1 U32570 ( .A1(n3322), .A2(n3321), .ZN(n3380) );
  OR2_X1 U32580 ( .A1(n3712), .A2(n3720), .ZN(n4130) );
  NAND2_X1 U32590 ( .A1(n4130), .A2(n3391), .ZN(n2531) );
  OAI21_X1 U32600 ( .B1(n2532), .B2(n3380), .A(n2531), .ZN(n2533) );
  NAND2_X1 U32610 ( .A1(n3322), .A2(n3348), .ZN(n4128) );
  NAND2_X1 U32620 ( .A1(n2778), .A2(REG3_REG_0__SCAN_IN), .ZN(n2538) );
  INV_X1 U32630 ( .A(REG0_REG_0__SCAN_IN), .ZN(n2534) );
  OR2_X1 U32640 ( .A1(n3259), .A2(n2534), .ZN(n2537) );
  NAND2_X1 U32650 ( .A1(n2572), .A2(REG2_REG_0__SCAN_IN), .ZN(n2535) );
  INV_X1 U32660 ( .A(REG3_REG_3__SCAN_IN), .ZN(n2543) );
  NAND2_X1 U32670 ( .A1(n2778), .A2(n2543), .ZN(n2549) );
  NAND2_X1 U32680 ( .A1(n2572), .A2(REG2_REG_3__SCAN_IN), .ZN(n2548) );
  INV_X1 U32690 ( .A(REG0_REG_3__SCAN_IN), .ZN(n2544) );
  OR2_X1 U32700 ( .A1(n3259), .A2(n2544), .ZN(n2547) );
  INV_X1 U32710 ( .A(REG1_REG_3__SCAN_IN), .ZN(n2545) );
  OR2_X1 U32720 ( .A1(n3262), .A2(n2545), .ZN(n2546) );
  NAND2_X1 U32730 ( .A1(n2550), .A2(IR_REG_31__SCAN_IN), .ZN(n2559) );
  XNOR2_X1 U32740 ( .A(n2559), .B(IR_REG_3__SCAN_IN), .ZN(n4886) );
  MUX2_X1 U32750 ( .A(n4886), .B(DATAI_3_), .S(n2144), .Z(n3553) );
  AND2_X1 U32760 ( .A1(n4284), .A2(n3553), .ZN(n2551) );
  INV_X1 U32770 ( .A(REG3_REG_4__SCAN_IN), .ZN(n2552) );
  XNOR2_X1 U32780 ( .A(n2552), .B(REG3_REG_3__SCAN_IN), .ZN(n3461) );
  NAND2_X1 U32790 ( .A1(n2778), .A2(n3461), .ZN(n2557) );
  NAND2_X1 U32800 ( .A1(n2572), .A2(REG2_REG_4__SCAN_IN), .ZN(n2556) );
  INV_X1 U32810 ( .A(REG1_REG_4__SCAN_IN), .ZN(n4889) );
  OR2_X1 U32820 ( .A1(n3262), .A2(n4889), .ZN(n2555) );
  INV_X1 U32830 ( .A(REG0_REG_4__SCAN_IN), .ZN(n2553) );
  OR2_X1 U32840 ( .A1(n3259), .A2(n2553), .ZN(n2554) );
  NAND2_X1 U32850 ( .A1(n2559), .A2(n2558), .ZN(n2560) );
  NAND2_X1 U32860 ( .A1(n2560), .A2(IR_REG_31__SCAN_IN), .ZN(n2562) );
  XNOR2_X1 U32870 ( .A(n2562), .B(n2561), .ZN(n4896) );
  INV_X1 U32880 ( .A(DATAI_4_), .ZN(n2886) );
  MUX2_X1 U32890 ( .A(n4896), .B(n2886), .S(n2144), .Z(n3460) );
  OR2_X1 U32900 ( .A1(n3578), .A2(n3460), .ZN(n4137) );
  NAND2_X1 U32910 ( .A1(n3578), .A2(n3460), .ZN(n4140) );
  INV_X1 U32920 ( .A(n3460), .ZN(n4023) );
  NAND2_X1 U32930 ( .A1(n3578), .A2(n4023), .ZN(n3497) );
  AND2_X1 U32940 ( .A1(n2571), .A2(n2563), .ZN(n2564) );
  NOR2_X1 U32950 ( .A1(n2595), .A2(n2564), .ZN(n3482) );
  NAND2_X1 U32960 ( .A1(n2778), .A2(n3482), .ZN(n2568) );
  INV_X1 U32970 ( .A(REG1_REG_7__SCAN_IN), .ZN(n3298) );
  OR2_X1 U32980 ( .A1(n3262), .A2(n3298), .ZN(n2567) );
  INV_X1 U32990 ( .A(REG0_REG_7__SCAN_IN), .ZN(n2565) );
  OR2_X1 U33000 ( .A1(n3259), .A2(n2565), .ZN(n2566) );
  NOR2_X1 U33010 ( .A1(n2591), .A2(IR_REG_5__SCAN_IN), .ZN(n2579) );
  NAND2_X1 U33020 ( .A1(n2579), .A2(n2570), .ZN(n2618) );
  NAND2_X1 U33030 ( .A1(n2618), .A2(IR_REG_31__SCAN_IN), .ZN(n2601) );
  XNOR2_X1 U33040 ( .A(n2601), .B(n2911), .ZN(n3299) );
  INV_X1 U33050 ( .A(DATAI_7_), .ZN(n2893) );
  MUX2_X1 U33060 ( .A(n3299), .B(n2893), .S(n2144), .Z(n3593) );
  OR2_X1 U33070 ( .A1(n4281), .A2(n3593), .ZN(n2800) );
  NAND2_X1 U33080 ( .A1(n4281), .A2(n3593), .ZN(n4144) );
  OAI21_X1 U33090 ( .B1(n2583), .B2(REG3_REG_6__SCAN_IN), .A(n2571), .ZN(n3478) );
  INV_X1 U33100 ( .A(n3478), .ZN(n3508) );
  NAND2_X1 U33110 ( .A1(n2572), .A2(REG2_REG_6__SCAN_IN), .ZN(n2577) );
  INV_X1 U33120 ( .A(REG1_REG_6__SCAN_IN), .ZN(n2573) );
  OR2_X1 U33130 ( .A1(n3262), .A2(n2573), .ZN(n2576) );
  INV_X1 U33140 ( .A(REG0_REG_6__SCAN_IN), .ZN(n2574) );
  OR2_X1 U33150 ( .A1(n3259), .A2(n2574), .ZN(n2575) );
  INV_X1 U33160 ( .A(n2579), .ZN(n2580) );
  NAND2_X1 U33170 ( .A1(n2580), .A2(IR_REG_31__SCAN_IN), .ZN(n2581) );
  XNOR2_X1 U33180 ( .A(n2581), .B(IR_REG_6__SCAN_IN), .ZN(n4885) );
  MUX2_X1 U33190 ( .A(n4885), .B(DATAI_6_), .S(n2144), .Z(n3605) );
  OR2_X1 U33200 ( .A1(n4282), .A2(n3605), .ZN(n2582) );
  NAND2_X1 U33210 ( .A1(n3610), .A2(n2582), .ZN(n2606) );
  AOI21_X1 U33220 ( .B1(REG3_REG_3__SCAN_IN), .B2(REG3_REG_4__SCAN_IN), .A(
        REG3_REG_5__SCAN_IN), .ZN(n2584) );
  NOR2_X1 U33230 ( .A1(n2584), .A2(n2583), .ZN(n3428) );
  NAND2_X1 U33240 ( .A1(n2778), .A2(n3428), .ZN(n2590) );
  NAND2_X1 U33250 ( .A1(n2572), .A2(REG2_REG_5__SCAN_IN), .ZN(n2589) );
  INV_X1 U33260 ( .A(REG0_REG_5__SCAN_IN), .ZN(n2585) );
  OR2_X1 U33270 ( .A1(n3259), .A2(n2585), .ZN(n2588) );
  INV_X1 U33280 ( .A(REG1_REG_5__SCAN_IN), .ZN(n2586) );
  OR2_X1 U33290 ( .A1(n3262), .A2(n2586), .ZN(n2587) );
  NAND2_X1 U33300 ( .A1(n2591), .A2(IR_REG_31__SCAN_IN), .ZN(n2592) );
  XNOR2_X1 U33310 ( .A(n2592), .B(IR_REG_5__SCAN_IN), .ZN(n3201) );
  MUX2_X1 U33320 ( .A(n3201), .B(DATAI_5_), .S(n2144), .Z(n3582) );
  NAND2_X1 U33330 ( .A1(n4283), .A2(n3582), .ZN(n3501) );
  NAND3_X1 U33340 ( .A1(n3610), .A2(n3605), .A3(n4282), .ZN(n2594) );
  NAND2_X1 U33350 ( .A1(n4281), .A2(n3597), .ZN(n2593) );
  OAI211_X1 U33360 ( .C1(n2606), .C2(n3501), .A(n2594), .B(n2593), .ZN(n3617)
         );
  OR2_X1 U33370 ( .A1(n2595), .A2(REG3_REG_8__SCAN_IN), .ZN(n2596) );
  AND2_X1 U33380 ( .A1(n2611), .A2(n2596), .ZN(n3629) );
  NAND2_X1 U33390 ( .A1(n2778), .A2(n3629), .ZN(n2600) );
  NAND2_X1 U33400 ( .A1(n2572), .A2(REG2_REG_8__SCAN_IN), .ZN(n2599) );
  INV_X1 U33410 ( .A(REG0_REG_8__SCAN_IN), .ZN(n2597) );
  OR2_X1 U33420 ( .A1(n3259), .A2(n2597), .ZN(n2598) );
  INV_X1 U33430 ( .A(REG1_REG_8__SCAN_IN), .ZN(n3129) );
  NAND4_X1 U33440 ( .A1(n2600), .A2(n2599), .A3(n2598), .A4(n2163), .ZN(n4681)
         );
  NAND2_X1 U33450 ( .A1(n2601), .A2(n2911), .ZN(n2602) );
  NAND2_X1 U33460 ( .A1(n2602), .A2(IR_REG_31__SCAN_IN), .ZN(n2603) );
  XNOR2_X1 U33470 ( .A(n2603), .B(IR_REG_8__SCAN_IN), .ZN(n3436) );
  MUX2_X1 U33480 ( .A(n3436), .B(DATAI_8_), .S(n2144), .Z(n3628) );
  NOR2_X1 U33490 ( .A1(n3617), .A2(n2466), .ZN(n2605) );
  AND2_X1 U33500 ( .A1(n3497), .A2(n2605), .ZN(n2604) );
  NAND2_X1 U33510 ( .A1(n3498), .A2(n2604), .ZN(n2609) );
  INV_X1 U33520 ( .A(n2605), .ZN(n2607) );
  NOR2_X1 U3353 ( .A1(n4283), .A2(n3582), .ZN(n3499) );
  NOR2_X1 U33540 ( .A1(n2606), .A2(n3499), .ZN(n3615) );
  NAND2_X1 U3355 ( .A1(n2611), .A2(n2610), .ZN(n2612) );
  AND2_X1 U3356 ( .A1(n2621), .A2(n2612), .ZN(n4692) );
  NAND2_X1 U3357 ( .A1(n2778), .A2(n4692), .ZN(n2617) );
  NAND2_X1 U3358 ( .A1(n2572), .A2(REG2_REG_9__SCAN_IN), .ZN(n2616) );
  INV_X1 U3359 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3446) );
  OR2_X1 U3360 ( .A1(n3262), .A2(n3446), .ZN(n2615) );
  INV_X1 U3361 ( .A(REG0_REG_9__SCAN_IN), .ZN(n2613) );
  OR2_X1 U3362 ( .A1(n3259), .A2(n2613), .ZN(n2614) );
  NAND2_X1 U3363 ( .A1(n2627), .A2(IR_REG_31__SCAN_IN), .ZN(n2619) );
  XNOR2_X1 U3364 ( .A(n2619), .B(IR_REG_9__SCAN_IN), .ZN(n4884) );
  MUX2_X1 U3365 ( .A(n4884), .B(DATAI_9_), .S(n2144), .Z(n4688) );
  AND2_X1 U3366 ( .A1(n4280), .A2(n4688), .ZN(n2620) );
  AND2_X1 U3367 ( .A1(n2621), .A2(n3042), .ZN(n2622) );
  OR2_X1 U3368 ( .A1(n2634), .A2(n2622), .ZN(n3941) );
  INV_X1 U3369 ( .A(n3941), .ZN(n4664) );
  NAND2_X1 U3370 ( .A1(n2778), .A2(n4664), .ZN(n2626) );
  NAND2_X1 U3371 ( .A1(n2572), .A2(REG2_REG_10__SCAN_IN), .ZN(n2625) );
  INV_X1 U3372 ( .A(REG0_REG_10__SCAN_IN), .ZN(n4870) );
  OR2_X1 U3373 ( .A1(n3259), .A2(n4870), .ZN(n2624) );
  OR2_X1 U3374 ( .A1(n3262), .A2(n4799), .ZN(n2623) );
  NAND4_X1 U3375 ( .A1(n2626), .A2(n2625), .A3(n2624), .A4(n2623), .ZN(n4078)
         );
  INV_X1 U3376 ( .A(n2627), .ZN(n2629) );
  NAND2_X1 U3377 ( .A1(n2629), .A2(n2628), .ZN(n2640) );
  NAND2_X1 U3378 ( .A1(n2640), .A2(IR_REG_31__SCAN_IN), .ZN(n2630) );
  XNOR2_X1 U3379 ( .A(n2630), .B(IR_REG_10__SCAN_IN), .ZN(n3526) );
  MUX2_X1 U3380 ( .A(n3526), .B(DATAI_10_), .S(n2144), .Z(n3731) );
  NOR2_X1 U3381 ( .A1(n4078), .A2(n3731), .ZN(n2631) );
  NAND2_X1 U3382 ( .A1(n4078), .A2(n3731), .ZN(n2632) );
  NAND2_X1 U3383 ( .A1(n2633), .A2(n2632), .ZN(n3646) );
  OR2_X1 U3384 ( .A1(n2634), .A2(REG3_REG_11__SCAN_IN), .ZN(n2635) );
  AND2_X1 U3385 ( .A1(n2660), .A2(n2635), .ZN(n4076) );
  NAND2_X1 U3386 ( .A1(n2778), .A2(n4076), .ZN(n2639) );
  NAND2_X1 U3387 ( .A1(n2572), .A2(REG2_REG_11__SCAN_IN), .ZN(n2638) );
  INV_X1 U3388 ( .A(REG0_REG_11__SCAN_IN), .ZN(n4866) );
  OR2_X1 U3389 ( .A1(n3259), .A2(n4866), .ZN(n2637) );
  INV_X1 U3390 ( .A(REG1_REG_11__SCAN_IN), .ZN(n4792) );
  OR2_X1 U3391 ( .A1(n3262), .A2(n4792), .ZN(n2636) );
  NAND4_X1 U3392 ( .A1(n2639), .A2(n2638), .A3(n2637), .A4(n2636), .ZN(n4279)
         );
  INV_X1 U3393 ( .A(n2640), .ZN(n2642) );
  INV_X1 U3394 ( .A(IR_REG_10__SCAN_IN), .ZN(n2641) );
  NAND2_X1 U3395 ( .A1(n2642), .A2(n2641), .ZN(n2643) );
  NAND2_X1 U3396 ( .A1(n2643), .A2(IR_REG_31__SCAN_IN), .ZN(n2650) );
  INV_X1 U3397 ( .A(DATAI_11_), .ZN(n2644) );
  MUX2_X1 U3398 ( .A(n3671), .B(n2644), .S(n2144), .Z(n3652) );
  OR2_X1 U3399 ( .A1(n4279), .A2(n3652), .ZN(n4165) );
  NAND2_X1 U3400 ( .A1(n4279), .A2(n3652), .ZN(n4159) );
  AND2_X1 U3401 ( .A1(n4165), .A2(n4159), .ZN(n3645) );
  XNOR2_X1 U3402 ( .A(n2660), .B(REG3_REG_12__SCAN_IN), .ZN(n3963) );
  NAND2_X1 U3403 ( .A1(n2778), .A2(n3963), .ZN(n2648) );
  NAND2_X1 U3404 ( .A1(n2572), .A2(REG2_REG_12__SCAN_IN), .ZN(n2647) );
  INV_X1 U3405 ( .A(REG1_REG_12__SCAN_IN), .ZN(n4788) );
  OR2_X1 U3406 ( .A1(n3262), .A2(n4788), .ZN(n2646) );
  INV_X1 U3407 ( .A(REG0_REG_12__SCAN_IN), .ZN(n4862) );
  OR2_X1 U3408 ( .A1(n3259), .A2(n4862), .ZN(n2645) );
  NAND4_X1 U3409 ( .A1(n2648), .A2(n2647), .A3(n2646), .A4(n2645), .ZN(n4632)
         );
  NAND2_X1 U3410 ( .A1(n2650), .A2(n2649), .ZN(n2651) );
  NAND2_X1 U3411 ( .A1(n2651), .A2(IR_REG_31__SCAN_IN), .ZN(n2652) );
  XNOR2_X1 U3412 ( .A(n2652), .B(IR_REG_12__SCAN_IN), .ZN(n4883) );
  INV_X1 U3413 ( .A(n2143), .ZN(n2653) );
  MUX2_X1 U3414 ( .A(DATAI_12_), .B(n4883), .S(n2653), .Z(n3965) );
  OR2_X1 U3415 ( .A1(n3645), .A2(n2467), .ZN(n2654) );
  INV_X1 U3416 ( .A(n3652), .ZN(n4079) );
  OR2_X1 U3417 ( .A1(n4279), .A2(n4079), .ZN(n3660) );
  OR2_X1 U3418 ( .A1(n4632), .A2(n3965), .ZN(n2655) );
  AND2_X1 U3419 ( .A1(n3660), .A2(n2655), .ZN(n2656) );
  OR2_X1 U3420 ( .A1(n2467), .A2(n2656), .ZN(n2657) );
  NAND2_X1 U3421 ( .A1(n2658), .A2(n2657), .ZN(n4625) );
  OAI21_X1 U3422 ( .B1(n2660), .B2(n2659), .A(n2993), .ZN(n2661) );
  AND2_X1 U3423 ( .A1(n2661), .A2(n2668), .ZN(n4053) );
  NAND2_X1 U3424 ( .A1(n2778), .A2(n4053), .ZN(n2665) );
  NAND2_X1 U3425 ( .A1(n2572), .A2(REG2_REG_13__SCAN_IN), .ZN(n2664) );
  OR2_X1 U3426 ( .A1(n3262), .A2(n4782), .ZN(n2663) );
  INV_X1 U3427 ( .A(REG0_REG_13__SCAN_IN), .ZN(n4858) );
  OR2_X1 U3428 ( .A1(n3259), .A2(n4858), .ZN(n2662) );
  NAND4_X1 U3429 ( .A1(n2665), .A2(n2664), .A3(n2663), .A4(n2662), .ZN(n4278)
         );
  OR2_X1 U3430 ( .A1(n2789), .A2(n2416), .ZN(n2666) );
  XNOR2_X1 U3431 ( .A(n2666), .B(IR_REG_13__SCAN_IN), .ZN(n4882) );
  MUX2_X1 U3432 ( .A(n4882), .B(DATAI_13_), .S(n2144), .Z(n4639) );
  NOR2_X1 U3433 ( .A1(n4278), .A2(n4639), .ZN(n2667) );
  INV_X1 U3434 ( .A(n4278), .ZN(n3858) );
  INV_X1 U3435 ( .A(n4639), .ZN(n4224) );
  AND2_X1 U3436 ( .A1(n2668), .A2(n3019), .ZN(n2669) );
  NOR2_X1 U3437 ( .A1(n2677), .A2(n2669), .ZN(n3908) );
  NAND2_X1 U3438 ( .A1(n2778), .A2(n3908), .ZN(n2673) );
  NAND2_X1 U3439 ( .A1(n2572), .A2(REG2_REG_14__SCAN_IN), .ZN(n2672) );
  INV_X1 U3440 ( .A(REG0_REG_14__SCAN_IN), .ZN(n4854) );
  OR2_X1 U3441 ( .A1(n3259), .A2(n4854), .ZN(n2671) );
  INV_X1 U3442 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4778) );
  OR2_X1 U3443 ( .A1(n3262), .A2(n4778), .ZN(n2670) );
  NAND4_X1 U3444 ( .A1(n2673), .A2(n2672), .A3(n2671), .A4(n2670), .ZN(n4608)
         );
  NAND2_X1 U3445 ( .A1(n2789), .A2(n2674), .ZN(n2714) );
  NAND2_X1 U3446 ( .A1(n2714), .A2(IR_REG_31__SCAN_IN), .ZN(n2676) );
  INV_X1 U3447 ( .A(IR_REG_14__SCAN_IN), .ZN(n2675) );
  XNOR2_X1 U3448 ( .A(n2676), .B(n2675), .ZN(n3704) );
  INV_X1 U3449 ( .A(DATAI_14_), .ZN(n2948) );
  MUX2_X1 U3450 ( .A(n3704), .B(n2948), .S(n2144), .Z(n4774) );
  OR2_X1 U3451 ( .A1(n4608), .A2(n4774), .ZN(n4161) );
  NAND2_X1 U3452 ( .A1(n4608), .A2(n4774), .ZN(n4147) );
  NOR2_X1 U3453 ( .A1(n2677), .A2(REG3_REG_15__SCAN_IN), .ZN(n2678) );
  OR2_X1 U3454 ( .A1(n2689), .A2(n2678), .ZN(n4617) );
  INV_X1 U3455 ( .A(n4617), .ZN(n2679) );
  NAND2_X1 U3456 ( .A1(n2679), .A2(n2778), .ZN(n2684) );
  INV_X1 U3457 ( .A(REG1_REG_15__SCAN_IN), .ZN(n4319) );
  OR2_X1 U34580 ( .A1(n3262), .A2(n4319), .ZN(n2683) );
  INV_X1 U34590 ( .A(REG0_REG_15__SCAN_IN), .ZN(n2680) );
  OR2_X1 U3460 ( .A1(n3259), .A2(n2680), .ZN(n2682) );
  NAND2_X1 U3461 ( .A1(n2572), .A2(REG2_REG_15__SCAN_IN), .ZN(n2681) );
  NAND4_X1 U3462 ( .A1(n2684), .A2(n2683), .A3(n2682), .A4(n2681), .ZN(n3990)
         );
  NAND2_X1 U3463 ( .A1(n2685), .A2(IR_REG_31__SCAN_IN), .ZN(n2687) );
  OR2_X1 U3464 ( .A1(n2687), .A2(n2686), .ZN(n2688) );
  NAND2_X1 U3465 ( .A1(n2687), .A2(n2686), .ZN(n2697) );
  MUX2_X1 U3466 ( .A(n4330), .B(DATAI_15_), .S(n2144), .Z(n4769) );
  AND2_X1 U34670 ( .A1(n3990), .A2(n4769), .ZN(n2701) );
  OR2_X1 U3468 ( .A1(n4200), .A2(n2701), .ZN(n4595) );
  OR2_X1 U34690 ( .A1(n2689), .A2(REG3_REG_16__SCAN_IN), .ZN(n2690) );
  AND2_X1 U3470 ( .A1(n2707), .A2(n2690), .ZN(n4592) );
  NAND2_X1 U34710 ( .A1(n4592), .A2(n2778), .ZN(n2696) );
  INV_X1 U3472 ( .A(REG1_REG_16__SCAN_IN), .ZN(n4917) );
  OR2_X1 U34730 ( .A1(n3262), .A2(n4917), .ZN(n2693) );
  INV_X1 U3474 ( .A(REG0_REG_16__SCAN_IN), .ZN(n2691) );
  OR2_X1 U34750 ( .A1(n3259), .A2(n2691), .ZN(n2692) );
  AND2_X1 U3476 ( .A1(n2693), .A2(n2692), .ZN(n2695) );
  NAND2_X1 U34770 ( .A1(n2572), .A2(REG2_REG_16__SCAN_IN), .ZN(n2694) );
  NAND2_X1 U3478 ( .A1(n2697), .A2(IR_REG_31__SCAN_IN), .ZN(n2699) );
  INV_X1 U34790 ( .A(n4983), .ZN(n2700) );
  MUX2_X1 U3480 ( .A(n2700), .B(DATAI_16_), .S(n2144), .Z(n4763) );
  AND2_X1 U34810 ( .A1(n4277), .A2(n4763), .ZN(n2704) );
  NAND2_X1 U3482 ( .A1(n4609), .A2(n4763), .ZN(n4237) );
  NAND2_X1 U34830 ( .A1(n4277), .A2(n4594), .ZN(n4234) );
  INV_X1 U3484 ( .A(n4600), .ZN(n4581) );
  OR2_X1 U34850 ( .A1(n4608), .A2(n3910), .ZN(n4613) );
  OR2_X1 U3486 ( .A1(n2701), .A2(n4613), .ZN(n2703) );
  OR2_X1 U34870 ( .A1(n3990), .A2(n4769), .ZN(n2702) );
  AND2_X1 U3488 ( .A1(n2703), .A2(n2702), .ZN(n4598) );
  AND2_X1 U34890 ( .A1(n4581), .A2(n4598), .ZN(n4597) );
  OR2_X1 U3490 ( .A1(n2704), .A2(n4597), .ZN(n2705) );
  NAND2_X1 U34910 ( .A1(n2707), .A2(n2706), .ZN(n2708) );
  NAND2_X1 U3492 ( .A1(n2718), .A2(n2708), .ZN(n4573) );
  OR2_X1 U34930 ( .A1(n4573), .A2(n2832), .ZN(n2712) );
  INV_X1 U3494 ( .A(REG1_REG_17__SCAN_IN), .ZN(n4761) );
  INV_X1 U34950 ( .A(REG0_REG_17__SCAN_IN), .ZN(n4848) );
  OAI22_X1 U3496 ( .A1(n3262), .A2(n4761), .B1(n3259), .B2(n4848), .ZN(n2709)
         );
  INV_X1 U34970 ( .A(n2709), .ZN(n2711) );
  NAND2_X1 U3498 ( .A1(n2572), .A2(REG2_REG_17__SCAN_IN), .ZN(n2710) );
  INV_X1 U34990 ( .A(n2741), .ZN(n2713) );
  NAND2_X1 U3500 ( .A1(n2725), .A2(IR_REG_31__SCAN_IN), .ZN(n2715) );
  INV_X1 U35010 ( .A(DATAI_17_), .ZN(n2716) );
  MUX2_X1 U3502 ( .A(n4981), .B(n2716), .S(n2144), .Z(n4561) );
  NAND2_X1 U35030 ( .A1(n4091), .A2(n4569), .ZN(n4546) );
  AND2_X1 U3504 ( .A1(n2718), .A2(n2717), .ZN(n2719) );
  OR2_X1 U35050 ( .A1(n2719), .A2(n2731), .ZN(n4555) );
  INV_X1 U35060 ( .A(REG1_REG_18__SCAN_IN), .ZN(n4315) );
  NAND2_X1 U35070 ( .A1(n2572), .A2(REG2_REG_18__SCAN_IN), .ZN(n2722) );
  INV_X1 U35080 ( .A(REG0_REG_18__SCAN_IN), .ZN(n2720) );
  OR2_X1 U35090 ( .A1(n3259), .A2(n2720), .ZN(n2721) );
  OAI211_X1 U35100 ( .C1(n3262), .C2(n4315), .A(n2722), .B(n2721), .ZN(n2723)
         );
  INV_X1 U35110 ( .A(n2723), .ZN(n2724) );
  OAI21_X1 U35120 ( .B1(n2725), .B2(IR_REG_17__SCAN_IN), .A(IR_REG_31__SCAN_IN), .ZN(n2726) );
  XNOR2_X1 U35130 ( .A(n2726), .B(IR_REG_18__SCAN_IN), .ZN(n4334) );
  INV_X1 U35140 ( .A(DATAI_18_), .ZN(n2727) );
  MUX2_X1 U35150 ( .A(n4980), .B(n2727), .S(n2144), .Z(n4552) );
  OR2_X1 U35160 ( .A1(n4564), .A2(n4552), .ZN(n4521) );
  NAND2_X1 U35170 ( .A1(n4564), .A2(n4552), .ZN(n4522) );
  INV_X1 U35180 ( .A(n4551), .ZN(n2728) );
  AND2_X1 U35190 ( .A1(n4546), .A2(n2728), .ZN(n2729) );
  OR2_X1 U35200 ( .A1(n4564), .A2(n4092), .ZN(n2730) );
  NOR2_X1 U35210 ( .A1(n2731), .A2(REG3_REG_19__SCAN_IN), .ZN(n2732) );
  OR2_X1 U35220 ( .A1(n2733), .A2(n2732), .ZN(n4536) );
  OR2_X1 U35230 ( .A1(n4536), .A2(n2832), .ZN(n2738) );
  INV_X1 U35240 ( .A(REG1_REG_19__SCAN_IN), .ZN(n4754) );
  NAND2_X1 U35250 ( .A1(n2572), .A2(REG2_REG_19__SCAN_IN), .ZN(n2735) );
  INV_X1 U35260 ( .A(REG0_REG_19__SCAN_IN), .ZN(n4843) );
  OR2_X1 U35270 ( .A1(n3259), .A2(n4843), .ZN(n2734) );
  OAI211_X1 U35280 ( .C1(n3262), .C2(n4754), .A(n2735), .B(n2734), .ZN(n2736)
         );
  INV_X1 U35290 ( .A(n2736), .ZN(n2737) );
  NOR2_X1 U35300 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_16__SCAN_IN), .ZN(n2739) );
  XNOR2_X2 U35310 ( .A(n2784), .B(IR_REG_19__SCAN_IN), .ZN(n4881) );
  MUX2_X1 U35320 ( .A(n4881), .B(DATAI_19_), .S(n2144), .Z(n4527) );
  AOI21_X1 U35330 ( .B1(n4483), .B2(n4505), .A(n4489), .ZN(n2742) );
  NAND2_X1 U35340 ( .A1(n4487), .A2(n4476), .ZN(n4244) );
  NAND2_X1 U35350 ( .A1(n4452), .A2(n4465), .ZN(n2820) );
  NAND2_X1 U35360 ( .A1(n4244), .A2(n2820), .ZN(n4469) );
  AND2_X1 U35370 ( .A1(n2743), .A2(n3920), .ZN(n2745) );
  NOR2_X1 U35380 ( .A1(n2745), .A2(n2744), .ZN(n4458) );
  INV_X1 U35390 ( .A(REG1_REG_23__SCAN_IN), .ZN(n4733) );
  NAND2_X1 U35400 ( .A1(n2572), .A2(REG2_REG_23__SCAN_IN), .ZN(n2747) );
  INV_X1 U35410 ( .A(REG0_REG_23__SCAN_IN), .ZN(n4830) );
  OR2_X1 U35420 ( .A1(n3259), .A2(n4830), .ZN(n2746) );
  OAI211_X1 U35430 ( .C1(n3262), .C2(n4733), .A(n2747), .B(n2746), .ZN(n2748)
         );
  NAND2_X1 U35440 ( .A1(n2144), .A2(DATAI_23_), .ZN(n4457) );
  NAND2_X1 U35450 ( .A1(n4068), .A2(n4457), .ZN(n2749) );
  INV_X1 U35460 ( .A(n4457), .ZN(n4451) );
  AND2_X2 U35470 ( .A1(n2751), .A2(REG3_REG_25__SCAN_IN), .ZN(n2768) );
  NOR2_X1 U35480 ( .A1(n2751), .A2(REG3_REG_25__SCAN_IN), .ZN(n2752) );
  INV_X1 U35490 ( .A(REG1_REG_25__SCAN_IN), .ZN(n4725) );
  NAND2_X1 U35500 ( .A1(n2572), .A2(REG2_REG_25__SCAN_IN), .ZN(n2754) );
  INV_X1 U35510 ( .A(REG0_REG_25__SCAN_IN), .ZN(n4822) );
  OR2_X1 U35520 ( .A1(n3259), .A2(n4822), .ZN(n2753) );
  OAI211_X1 U35530 ( .C1(n3262), .C2(n4725), .A(n2754), .B(n2753), .ZN(n2755)
         );
  INV_X1 U35540 ( .A(n2755), .ZN(n2756) );
  NOR2_X1 U35550 ( .A1(n4399), .A2(n4414), .ZN(n2757) );
  INV_X1 U35560 ( .A(n4399), .ZN(n4438) );
  INV_X1 U35570 ( .A(REG3_REG_26__SCAN_IN), .ZN(n2758) );
  XNOR2_X1 U35580 ( .A(n2768), .B(n2758), .ZN(n4407) );
  NAND2_X1 U35590 ( .A1(n4407), .A2(n2778), .ZN(n2763) );
  INV_X1 U35600 ( .A(REG1_REG_26__SCAN_IN), .ZN(n4722) );
  NAND2_X1 U35610 ( .A1(n2572), .A2(REG2_REG_26__SCAN_IN), .ZN(n2760) );
  INV_X1 U35620 ( .A(REG0_REG_26__SCAN_IN), .ZN(n4818) );
  OAI211_X1 U35630 ( .C1(n3262), .C2(n4722), .A(n2760), .B(n2759), .ZN(n2761)
         );
  INV_X1 U35640 ( .A(n2761), .ZN(n2762) );
  NAND2_X1 U35650 ( .A1(n2144), .A2(DATAI_26_), .ZN(n4720) );
  NOR2_X1 U35660 ( .A1(n4418), .A2(n4720), .ZN(n2764) );
  NAND2_X1 U35670 ( .A1(n2768), .A2(REG3_REG_26__SCAN_IN), .ZN(n2766) );
  INV_X1 U35680 ( .A(REG3_REG_27__SCAN_IN), .ZN(n2765) );
  NAND2_X1 U35690 ( .A1(n2766), .A2(n2765), .ZN(n2769) );
  AND2_X1 U35700 ( .A1(REG3_REG_27__SCAN_IN), .A2(REG3_REG_26__SCAN_IN), .ZN(
        n2767) );
  NAND2_X1 U35710 ( .A1(n2768), .A2(n2767), .ZN(n2776) );
  NAND2_X1 U35720 ( .A1(n2769), .A2(n2776), .ZN(n4386) );
  INV_X1 U35730 ( .A(REG1_REG_27__SCAN_IN), .ZN(n2772) );
  NAND2_X1 U35740 ( .A1(n2572), .A2(REG2_REG_27__SCAN_IN), .ZN(n2771) );
  INV_X1 U35750 ( .A(REG0_REG_27__SCAN_IN), .ZN(n3080) );
  OR2_X1 U35760 ( .A1(n3259), .A2(n3080), .ZN(n2770) );
  OAI211_X1 U35770 ( .C1(n3262), .C2(n2772), .A(n2771), .B(n2770), .ZN(n2773)
         );
  INV_X1 U35780 ( .A(n2773), .ZN(n2774) );
  NAND2_X1 U35790 ( .A1(n2144), .A2(DATAI_27_), .ZN(n4384) );
  NAND2_X1 U35800 ( .A1(n2776), .A2(n3079), .ZN(n2777) );
  NAND2_X1 U35810 ( .A1(n3894), .A2(n2778), .ZN(n2783) );
  INV_X1 U3582 ( .A(REG1_REG_28__SCAN_IN), .ZN(n3033) );
  NAND2_X1 U3583 ( .A1(n2572), .A2(REG2_REG_28__SCAN_IN), .ZN(n2780) );
  INV_X1 U3584 ( .A(REG0_REG_28__SCAN_IN), .ZN(n3032) );
  OR2_X1 U3585 ( .A1(n3259), .A2(n3032), .ZN(n2779) );
  OAI211_X1 U3586 ( .C1(n3033), .C2(n3262), .A(n2780), .B(n2779), .ZN(n2781)
         );
  INV_X1 U3587 ( .A(n2781), .ZN(n2782) );
  NAND2_X1 U3588 ( .A1(n4369), .A2(n3895), .ZN(n4362) );
  NAND2_X1 U3589 ( .A1(n4392), .A2(n4358), .ZN(n4364) );
  XNOR2_X1 U3590 ( .A(n4357), .B(n4356), .ZN(n3902) );
  NAND2_X1 U3591 ( .A1(n2784), .A2(n2925), .ZN(n2785) );
  XNOR2_X2 U3592 ( .A(n2786), .B(n2924), .ZN(n2868) );
  INV_X1 U3593 ( .A(n2787), .ZN(n2788) );
  NAND2_X1 U3594 ( .A1(n2839), .A2(IR_REG_31__SCAN_IN), .ZN(n2790) );
  XNOR2_X2 U3595 ( .A(n2792), .B(IR_REG_22__SCAN_IN), .ZN(n4879) );
  XNOR2_X1 U3596 ( .A(n3408), .B(n4879), .ZN(n2793) );
  NAND2_X1 U3597 ( .A1(n2868), .A2(n4881), .ZN(n4951) );
  INV_X1 U3598 ( .A(n4879), .ZN(n2794) );
  INV_X1 U3599 ( .A(n4264), .ZN(n4125) );
  INV_X1 U3600 ( .A(n4220), .ZN(n3284) );
  OR2_X1 U3601 ( .A1(n3313), .A2(n3855), .ZN(n4126) );
  INV_X1 U3602 ( .A(n4126), .ZN(n3285) );
  NAND2_X1 U3603 ( .A1(n3284), .A2(n3285), .ZN(n3386) );
  NAND2_X1 U3604 ( .A1(n3386), .A2(n4131), .ZN(n2795) );
  NAND2_X1 U3605 ( .A1(n3712), .A2(n3720), .ZN(n4134) );
  NAND2_X1 U3606 ( .A1(n2795), .A2(n4223), .ZN(n3388) );
  INV_X1 U3607 ( .A(n3553), .ZN(n2796) );
  OR2_X1 U3608 ( .A1(n4284), .A2(n2796), .ZN(n4136) );
  NAND2_X1 U3609 ( .A1(n4284), .A2(n2796), .ZN(n4133) );
  INV_X1 U3610 ( .A(n4137), .ZN(n2797) );
  OR2_X1 U3611 ( .A1(n4283), .A2(n2306), .ZN(n4151) );
  AND2_X1 U3612 ( .A1(n4283), .A2(n2306), .ZN(n3576) );
  INV_X1 U3613 ( .A(n3605), .ZN(n2798) );
  NAND2_X1 U3614 ( .A1(n4282), .A2(n2798), .ZN(n4152) );
  NAND2_X1 U3615 ( .A1(n3496), .A2(n4152), .ZN(n2799) );
  OR2_X1 U3616 ( .A1(n4282), .A2(n2798), .ZN(n4142) );
  INV_X1 U3617 ( .A(n2800), .ZN(n3621) );
  OR2_X1 U3618 ( .A1(n4280), .A2(n2309), .ZN(n4217) );
  INV_X1 U3619 ( .A(n4217), .ZN(n2802) );
  NAND2_X1 U3620 ( .A1(n4681), .A2(n3634), .ZN(n4674) );
  AND2_X1 U3621 ( .A1(n4280), .A2(n2309), .ZN(n4149) );
  INV_X1 U3622 ( .A(n4149), .ZN(n4218) );
  AND2_X1 U3623 ( .A1(n4218), .A2(n4674), .ZN(n2801) );
  OR2_X1 U3624 ( .A1(n2802), .A2(n2801), .ZN(n4653) );
  NAND2_X1 U3625 ( .A1(n4078), .A2(n4794), .ZN(n4208) );
  INV_X1 U3626 ( .A(n2806), .ZN(n2803) );
  OR2_X1 U3627 ( .A1(n4681), .A2(n3634), .ZN(n4672) );
  AND2_X1 U3628 ( .A1(n4672), .A2(n4217), .ZN(n4652) );
  OR2_X1 U3629 ( .A1(n3621), .A2(n2808), .ZN(n2804) );
  OR2_X1 U3630 ( .A1(n4078), .A2(n4794), .ZN(n4209) );
  INV_X1 U3631 ( .A(n4209), .ZN(n2810) );
  AND2_X1 U3632 ( .A1(n4144), .A2(n2806), .ZN(n2807) );
  OR2_X1 U3633 ( .A1(n2808), .A2(n2807), .ZN(n2809) );
  OR2_X1 U3634 ( .A1(n2810), .A2(n2809), .ZN(n3642) );
  AND2_X1 U3635 ( .A1(n3642), .A2(n4159), .ZN(n2811) );
  NAND2_X1 U3636 ( .A1(n4632), .A2(n4784), .ZN(n4627) );
  NAND2_X1 U3637 ( .A1(n4278), .A2(n4224), .ZN(n2812) );
  AND2_X1 U3638 ( .A1(n4627), .A2(n2812), .ZN(n4160) );
  NOR2_X1 U3639 ( .A1(n4632), .A2(n4784), .ZN(n4628) );
  NOR2_X1 U3640 ( .A1(n4278), .A2(n4224), .ZN(n2813) );
  AOI21_X1 U3641 ( .B1(n4160), .B2(n4628), .A(n2813), .ZN(n4164) );
  OR2_X1 U3642 ( .A1(n3990), .A2(n2875), .ZN(n4162) );
  NAND2_X1 U3643 ( .A1(n3990), .A2(n2875), .ZN(n4148) );
  NAND2_X1 U3644 ( .A1(n4162), .A2(n4148), .ZN(n4615) );
  NAND2_X1 U3645 ( .A1(n4611), .A2(n4148), .ZN(n4580) );
  INV_X1 U3646 ( .A(n4527), .ZN(n4535) );
  NAND2_X1 U3647 ( .A1(n4545), .A2(n4535), .ZN(n2815) );
  AND2_X1 U3648 ( .A1(n2815), .A2(n4522), .ZN(n2816) );
  NAND2_X1 U3649 ( .A1(n4091), .A2(n4561), .ZN(n4518) );
  NAND2_X1 U3650 ( .A1(n2816), .A2(n4518), .ZN(n4235) );
  AND2_X1 U3651 ( .A1(n4484), .A2(n4512), .ZN(n4172) );
  INV_X1 U3652 ( .A(n2816), .ZN(n2818) );
  NAND2_X1 U3653 ( .A1(n4584), .A2(n4569), .ZN(n4519) );
  AND2_X1 U3654 ( .A1(n4521), .A2(n4519), .ZN(n2817) );
  OAI22_X1 U3655 ( .A1(n2818), .A2(n2817), .B1(n4535), .B2(n4545), .ZN(n4499)
         );
  NOR2_X1 U3656 ( .A1(n4484), .A2(n4512), .ZN(n2819) );
  OR2_X1 U3657 ( .A1(n4499), .A2(n2819), .ZN(n4240) );
  INV_X1 U3658 ( .A(n4172), .ZN(n4239) );
  NAND2_X1 U3659 ( .A1(n4240), .A2(n4239), .ZN(n4175) );
  AND2_X1 U3660 ( .A1(n4466), .A2(n4483), .ZN(n4216) );
  NAND2_X1 U3661 ( .A1(n4505), .A2(n4492), .ZN(n4174) );
  NAND2_X1 U3662 ( .A1(n4473), .A2(n4457), .ZN(n4198) );
  OR2_X1 U3663 ( .A1(n4415), .A2(n4440), .ZN(n4197) );
  OR2_X1 U3664 ( .A1(n4473), .A2(n4457), .ZN(n4430) );
  AND2_X1 U3665 ( .A1(n4197), .A2(n4430), .ZN(n4245) );
  NAND2_X1 U3666 ( .A1(n4415), .A2(n4440), .ZN(n4196) );
  AND2_X1 U3667 ( .A1(n4399), .A2(n4421), .ZN(n4396) );
  NAND2_X1 U3668 ( .A1(n4391), .A2(n4720), .ZN(n4254) );
  INV_X1 U3669 ( .A(n4254), .ZN(n2822) );
  OR2_X1 U3670 ( .A1(n4396), .A2(n2822), .ZN(n2821) );
  OR2_X1 U3671 ( .A1(n4399), .A2(n4421), .ZN(n4397) );
  AND2_X1 U3672 ( .A1(n4202), .A2(n4397), .ZN(n4251) );
  NAND2_X1 U3673 ( .A1(n4400), .A2(n4384), .ZN(n4182) );
  XNOR2_X1 U3674 ( .A(n4365), .B(n4204), .ZN(n2826) );
  NAND2_X1 U3675 ( .A1(n4880), .A2(n4264), .ZN(n2825) );
  NAND2_X1 U3676 ( .A1(n4879), .A2(n4881), .ZN(n2824) );
  NAND2_X1 U3677 ( .A1(n2826), .A2(n4525), .ZN(n2837) );
  INV_X1 U3678 ( .A(REG1_REG_29__SCAN_IN), .ZN(n2829) );
  NAND2_X1 U3679 ( .A1(n2572), .A2(REG2_REG_29__SCAN_IN), .ZN(n2828) );
  INV_X1 U3680 ( .A(REG0_REG_29__SCAN_IN), .ZN(n3060) );
  OR2_X1 U3681 ( .A1(n3259), .A2(n3060), .ZN(n2827) );
  OAI211_X1 U3682 ( .C1(n3262), .C2(n2829), .A(n2828), .B(n2827), .ZN(n2830)
         );
  INV_X1 U3683 ( .A(n2830), .ZN(n2831) );
  NAND2_X1 U3684 ( .A1(n2833), .A2(IR_REG_31__SCAN_IN), .ZN(n2835) );
  XNOR2_X1 U3685 ( .A(n2835), .B(n2834), .ZN(n4888) );
  INV_X1 U3686 ( .A(n3167), .ZN(n3328) );
  AOI22_X1 U3687 ( .A1(n4276), .A2(n4563), .B1(n4400), .B2(n4682), .ZN(n2836)
         );
  NAND2_X1 U3688 ( .A1(n2837), .A2(n2836), .ZN(n3900) );
  AOI21_X1 U3689 ( .B1(n3895), .B2(n4768), .A(n3900), .ZN(n2838) );
  NAND2_X1 U3690 ( .A1(n2866), .A2(n2867), .ZN(n2841) );
  XNOR2_X1 U3691 ( .A(n2846), .B(n2845), .ZN(n2864) );
  NAND2_X1 U3692 ( .A1(n2863), .A2(n2864), .ZN(n2847) );
  MUX2_X1 U3693 ( .A(n2863), .B(n2847), .S(B_REG_SCAN_IN), .Z(n2850) );
  NAND2_X1 U3694 ( .A1(n2848), .A2(IR_REG_31__SCAN_IN), .ZN(n2849) );
  NAND2_X1 U3695 ( .A1(n2861), .A2(n3163), .ZN(n2851) );
  INV_X1 U3696 ( .A(n4878), .ZN(n2862) );
  NAND2_X1 U3697 ( .A1(n2863), .A2(n2862), .ZN(n3161) );
  NOR4_X1 U3698 ( .A1(D_REG_7__SCAN_IN), .A2(D_REG_9__SCAN_IN), .A3(
        D_REG_10__SCAN_IN), .A4(D_REG_15__SCAN_IN), .ZN(n2855) );
  NOR4_X1 U3699 ( .A1(D_REG_8__SCAN_IN), .A2(D_REG_3__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_6__SCAN_IN), .ZN(n2854) );
  INV_X1 U3700 ( .A(D_REG_19__SCAN_IN), .ZN(n4968) );
  INV_X1 U3701 ( .A(D_REG_31__SCAN_IN), .ZN(n4959) );
  INV_X1 U3702 ( .A(D_REG_23__SCAN_IN), .ZN(n4965) );
  INV_X1 U3703 ( .A(D_REG_25__SCAN_IN), .ZN(n4964) );
  NAND4_X1 U3704 ( .A1(n4968), .A2(n4959), .A3(n4965), .A4(n4964), .ZN(n2852)
         );
  NOR2_X1 U3705 ( .A1(D_REG_20__SCAN_IN), .A2(n2852), .ZN(n2909) );
  NOR4_X1 U3706 ( .A1(D_REG_22__SCAN_IN), .A2(D_REG_16__SCAN_IN), .A3(
        D_REG_12__SCAN_IN), .A4(D_REG_13__SCAN_IN), .ZN(n2853) );
  AND4_X1 U3707 ( .A1(n2855), .A2(n2854), .A3(n2909), .A4(n2853), .ZN(n2860)
         );
  NOR4_X1 U3708 ( .A1(D_REG_24__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_2__SCAN_IN), .A4(D_REG_11__SCAN_IN), .ZN(n2858) );
  NOR4_X1 U3709 ( .A1(D_REG_17__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        D_REG_30__SCAN_IN), .A4(D_REG_4__SCAN_IN), .ZN(n2857) );
  NOR4_X1 U3710 ( .A1(D_REG_18__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_28__SCAN_IN), .A4(D_REG_26__SCAN_IN), .ZN(n2856) );
  INV_X1 U3711 ( .A(D_REG_21__SCAN_IN), .ZN(n4966) );
  AND4_X1 U3712 ( .A1(n2858), .A2(n2857), .A3(n2856), .A4(n4966), .ZN(n2859)
         );
  NAND2_X1 U3713 ( .A1(n2860), .A2(n2859), .ZN(n3323) );
  NAND2_X1 U3714 ( .A1(n2861), .A2(n3323), .ZN(n2873) );
  NAND2_X1 U3715 ( .A1(n2864), .A2(n2862), .ZN(n3324) );
  OAI21_X1 U3716 ( .B1(n3326), .B2(D_REG_1__SCAN_IN), .A(n3324), .ZN(n2872) );
  INV_X1 U3717 ( .A(n2864), .ZN(n2897) );
  NAND3_X2 U3718 ( .A1(n2865), .A2(n4878), .A3(n2897), .ZN(n3369) );
  NAND2_X1 U3719 ( .A1(n2868), .A2(n4339), .ZN(n2869) );
  NAND2_X1 U3720 ( .A1(n3167), .A2(n2869), .ZN(n3401) );
  NAND2_X1 U3721 ( .A1(n3341), .A2(n3401), .ZN(n2870) );
  NOR2_X1 U3722 ( .A1(n3403), .A2(n2870), .ZN(n2871) );
  NAND2_X1 U3723 ( .A1(n3393), .A2(n3720), .ZN(n3552) );
  NAND2_X1 U3724 ( .A1(n3663), .A2(n4784), .ZN(n4640) );
  NAND2_X1 U3725 ( .A1(n4533), .A2(n4512), .ZN(n4511) );
  AND2_X1 U3726 ( .A1(n4382), .A2(n4384), .ZN(n4383) );
  NOR2_X1 U3727 ( .A1(n4714), .A2(n3895), .ZN(n4341) );
  NAND2_X1 U3728 ( .A1(n4382), .A2(n4341), .ZN(n4372) );
  OAI21_X1 U3729 ( .B1(n4383), .B2(n4358), .A(n4372), .ZN(n3898) );
  OR2_X1 U3731 ( .A1(n3898), .A2(n4872), .ZN(n2877) );
  NAND2_X1 U3732 ( .A1(n5012), .A2(REG0_REG_28__SCAN_IN), .ZN(n2876) );
  NAND2_X1 U3733 ( .A1(n2880), .A2(n5019), .ZN(n2884) );
  OR2_X1 U3734 ( .A1(n5019), .A2(n3033), .ZN(n2881) );
  OAI21_X1 U3735 ( .B1(n3898), .B2(n4801), .A(n2881), .ZN(n2882) );
  NAND2_X1 U3736 ( .A1(n2884), .A2(n2883), .ZN(U3546) );
  INV_X1 U3737 ( .A(n4978), .ZN(n2885) );
  INV_X2 U3738 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  MUX2_X1 U3739 ( .A(n2886), .B(n4896), .S(STATE_REG_SCAN_IN), .Z(n2887) );
  INV_X1 U3740 ( .A(n2887), .ZN(U3348) );
  INV_X1 U3741 ( .A(n3201), .ZN(n3243) );
  INV_X1 U3742 ( .A(DATAI_5_), .ZN(n2888) );
  MUX2_X1 U3743 ( .A(n3243), .B(n2888), .S(U3149), .Z(n2889) );
  INV_X1 U3744 ( .A(n2889), .ZN(U3347) );
  INV_X1 U3745 ( .A(DATAI_21_), .ZN(n2891) );
  NAND2_X1 U3746 ( .A1(n4264), .A2(STATE_REG_SCAN_IN), .ZN(n2890) );
  OAI21_X1 U3747 ( .B1(STATE_REG_SCAN_IN), .B2(n2891), .A(n2890), .ZN(U3331)
         );
  MUX2_X1 U3748 ( .A(n2948), .B(n3704), .S(STATE_REG_SCAN_IN), .Z(n2892) );
  INV_X1 U3749 ( .A(n2892), .ZN(U3338) );
  MUX2_X1 U3750 ( .A(n2893), .B(n3299), .S(STATE_REG_SCAN_IN), .Z(n2894) );
  INV_X1 U3751 ( .A(n2894), .ZN(U3345) );
  INV_X1 U3752 ( .A(DATAI_27_), .ZN(n3090) );
  XNOR2_X1 U3753 ( .A(n2895), .B(IR_REG_27__SCAN_IN), .ZN(n4343) );
  NAND2_X1 U3754 ( .A1(n4343), .A2(STATE_REG_SCAN_IN), .ZN(n2896) );
  OAI21_X1 U3755 ( .B1(STATE_REG_SCAN_IN), .B2(n3090), .A(n2896), .ZN(U3325)
         );
  INV_X1 U3756 ( .A(DATAI_25_), .ZN(n3068) );
  NAND2_X1 U3757 ( .A1(n2897), .A2(STATE_REG_SCAN_IN), .ZN(n2898) );
  OAI21_X1 U3758 ( .B1(STATE_REG_SCAN_IN), .B2(n3068), .A(n2898), .ZN(U3327)
         );
  INV_X1 U3759 ( .A(DATAI_8_), .ZN(n2899) );
  INV_X1 U3760 ( .A(n3436), .ZN(n3444) );
  MUX2_X1 U3761 ( .A(n2899), .B(n3444), .S(STATE_REG_SCAN_IN), .Z(n2900) );
  INV_X1 U3762 ( .A(n2900), .ZN(U3344) );
  INV_X1 U3763 ( .A(DATAI_24_), .ZN(n2901) );
  MUX2_X1 U3764 ( .A(n2863), .B(n2901), .S(U3149), .Z(n2902) );
  INV_X1 U3765 ( .A(n2902), .ZN(U3328) );
  INV_X1 U3766 ( .A(DATAI_29_), .ZN(n2905) );
  NAND2_X1 U3767 ( .A1(n2903), .A2(STATE_REG_SCAN_IN), .ZN(n2904) );
  OAI21_X1 U3768 ( .B1(STATE_REG_SCAN_IN), .B2(n2905), .A(n2904), .ZN(U3323)
         );
  MUX2_X1 U3769 ( .A(n2644), .B(n3671), .S(STATE_REG_SCAN_IN), .Z(n2906) );
  INV_X1 U3770 ( .A(n2906), .ZN(U3341) );
  INV_X1 U3771 ( .A(DATAI_10_), .ZN(n2907) );
  INV_X1 U3772 ( .A(n3526), .ZN(n3442) );
  MUX2_X1 U3773 ( .A(n2907), .B(n3442), .S(STATE_REG_SCAN_IN), .Z(n2908) );
  INV_X1 U3774 ( .A(n2908), .ZN(U3342) );
  INV_X1 U3775 ( .A(DATAO_REG_31__SCAN_IN), .ZN(n3258) );
  NAND4_X1 U3776 ( .A1(IR_REG_29__SCAN_IN), .A2(n2909), .A3(
        DATAO_REG_2__SCAN_IN), .A4(n3258), .ZN(n2944) );
  INV_X1 U3777 ( .A(REG3_REG_15__SCAN_IN), .ZN(n3024) );
  NAND4_X1 U3778 ( .A1(REG0_REG_3__SCAN_IN), .A2(ADDR_REG_4__SCAN_IN), .A3(
        n3024), .A4(n3019), .ZN(n2910) );
  NOR3_X1 U3779 ( .A1(REG1_REG_9__SCAN_IN), .A2(ADDR_REG_16__SCAN_IN), .A3(
        n2910), .ZN(n2917) );
  INV_X1 U3780 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4012) );
  INV_X1 U3781 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4920) );
  INV_X1 U3782 ( .A(ADDR_REG_0__SCAN_IN), .ZN(n3013) );
  NAND4_X1 U3783 ( .A1(ADDR_REG_1__SCAN_IN), .A2(n4012), .A3(n4920), .A4(n3013), .ZN(n2915) );
  INV_X1 U3784 ( .A(ADDR_REG_3__SCAN_IN), .ZN(n3008) );
  NAND4_X1 U3785 ( .A1(DATAI_20_), .A2(REG3_REG_25__SCAN_IN), .A3(
        ADDR_REG_19__SCAN_IN), .A4(n3008), .ZN(n2914) );
  NAND4_X1 U3786 ( .A1(D_REG_8__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        REG1_REG_28__SCAN_IN), .A4(n3032), .ZN(n2913) );
  NAND4_X1 U3787 ( .A1(n2911), .A2(IR_REG_8__SCAN_IN), .A3(IR_REG_5__SCAN_IN), 
        .A4(D_REG_30__SCAN_IN), .ZN(n2912) );
  NOR4_X1 U3788 ( .A1(n2915), .A2(n2914), .A3(n2913), .A4(n2912), .ZN(n2916)
         );
  NAND4_X1 U3789 ( .A1(IR_REG_3__SCAN_IN), .A2(DATAI_2_), .A3(n2917), .A4(
        n2916), .ZN(n2943) );
  INV_X1 U3790 ( .A(REG2_REG_21__SCAN_IN), .ZN(n3141) );
  INV_X1 U3791 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n3264) );
  NAND4_X1 U3792 ( .A1(ADDR_REG_14__SCAN_IN), .A2(ADDR_REG_11__SCAN_IN), .A3(
        n3141), .A4(n3264), .ZN(n2922) );
  INV_X1 U3793 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n3253) );
  NAND4_X1 U3794 ( .A1(REG1_REG_14__SCAN_IN), .A2(n2510), .A3(n3129), .A4(
        n3253), .ZN(n2918) );
  NOR2_X1 U3795 ( .A1(REG3_REG_6__SCAN_IN), .A2(n2918), .ZN(n2919) );
  INV_X1 U3796 ( .A(REG2_REG_30__SCAN_IN), .ZN(n4355) );
  NAND4_X1 U3797 ( .A1(n2919), .A2(REG2_REG_3__SCAN_IN), .A3(D_REG_11__SCAN_IN), .A4(n4355), .ZN(n2921) );
  NAND4_X1 U3798 ( .A1(IR_REG_17__SCAN_IN), .A2(REG2_REG_20__SCAN_IN), .A3(
        REG0_REG_14__SCAN_IN), .A4(DATAO_REG_12__SCAN_IN), .ZN(n2920) );
  NOR3_X1 U3799 ( .A1(n2922), .A2(n2921), .A3(n2920), .ZN(n2941) );
  AND4_X1 U3800 ( .A1(D_REG_1__SCAN_IN), .A2(D_REG_2__SCAN_IN), .A3(
        REG2_REG_11__SCAN_IN), .A4(DATAI_26_), .ZN(n2928) );
  INV_X1 U3801 ( .A(REG3_REG_19__SCAN_IN), .ZN(n3118) );
  AND4_X1 U3802 ( .A1(REG1_REG_11__SCAN_IN), .A2(DATAI_7_), .A3(DATAI_1_), 
        .A4(n3118), .ZN(n2923) );
  AND4_X1 U3803 ( .A1(n2925), .A2(n2924), .A3(DATAI_17_), .A4(n2923), .ZN(
        n2927) );
  INV_X1 U3804 ( .A(DATAO_REG_15__SCAN_IN), .ZN(n3266) );
  AND2_X1 U3805 ( .A1(REG2_REG_5__SCAN_IN), .A2(D_REG_0__SCAN_IN), .ZN(n2926)
         );
  AND4_X1 U3806 ( .A1(n2928), .A2(n2927), .A3(n3266), .A4(n2926), .ZN(n2940)
         );
  NAND4_X1 U3807 ( .A1(D_REG_28__SCAN_IN), .A2(D_REG_26__SCAN_IN), .A3(
        D_REG_17__SCAN_IN), .A4(REG0_REG_1__SCAN_IN), .ZN(n2932) );
  NAND4_X1 U3808 ( .A1(ADDR_REG_7__SCAN_IN), .A2(n2570), .A3(n4830), .A4(n4733), .ZN(n2931) );
  NAND4_X1 U3809 ( .A1(REG3_REG_5__SCAN_IN), .A2(REG2_REG_26__SCAN_IN), .A3(
        DATAO_REG_10__SCAN_IN), .A4(n3867), .ZN(n2930) );
  NAND4_X1 U3810 ( .A1(REG3_REG_13__SCAN_IN), .A2(D_REG_29__SCAN_IN), .A3(
        DATAO_REG_4__SCAN_IN), .A4(n4866), .ZN(n2929) );
  NOR4_X1 U3811 ( .A1(n2932), .A2(n2931), .A3(n2930), .A4(n2929), .ZN(n2939)
         );
  NAND4_X1 U3812 ( .A1(D_REG_14__SCAN_IN), .A2(REG3_REG_20__SCAN_IN), .A3(
        REG0_REG_0__SCAN_IN), .A4(n2641), .ZN(n2937) );
  INV_X1 U3813 ( .A(ADDR_REG_8__SCAN_IN), .ZN(n2935) );
  INV_X1 U3814 ( .A(DATAI_31_), .ZN(n3868) );
  INV_X1 U3815 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n3280) );
  NAND4_X1 U3816 ( .A1(REG2_REG_31__SCAN_IN), .A2(REG2_REG_18__SCAN_IN), .A3(
        n3868), .A4(n3280), .ZN(n2934) );
  INV_X1 U3817 ( .A(DATAO_REG_27__SCAN_IN), .ZN(n3495) );
  NAND4_X1 U3818 ( .A1(REG3_REG_23__SCAN_IN), .A2(IR_REG_13__SCAN_IN), .A3(
        REG0_REG_31__SCAN_IN), .A4(n3495), .ZN(n2933) );
  OR4_X1 U3819 ( .A1(n2935), .A2(IR_REG_9__SCAN_IN), .A3(n2934), .A4(n2933), 
        .ZN(n2936) );
  NOR4_X1 U3820 ( .A1(n2937), .A2(n2936), .A3(DATAI_22_), .A4(n4799), .ZN(
        n2938) );
  NAND4_X1 U3821 ( .A1(n2941), .A2(n2940), .A3(n2939), .A4(n2938), .ZN(n2942)
         );
  NOR4_X1 U3822 ( .A1(REG3_REG_10__SCAN_IN), .A2(n2944), .A3(n2943), .A4(n2942), .ZN(n2960) );
  INV_X1 U3823 ( .A(D_REG_18__SCAN_IN), .ZN(n4969) );
  NOR4_X1 U3824 ( .A1(ADDR_REG_5__SCAN_IN), .A2(n3060), .A3(n4969), .A4(n2585), 
        .ZN(n2958) );
  INV_X1 U3825 ( .A(IR_REG_12__SCAN_IN), .ZN(n3092) );
  INV_X1 U3826 ( .A(REG2_REG_25__SCAN_IN), .ZN(n3056) );
  NOR4_X1 U3827 ( .A1(IR_REG_24__SCAN_IN), .A2(n3092), .A3(n3056), .A4(n4835), 
        .ZN(n2957) );
  INV_X1 U3828 ( .A(DATAI_3_), .ZN(n2946) );
  INV_X1 U3829 ( .A(REG2_REG_2__SCAN_IN), .ZN(n2945) );
  NOR4_X1 U3830 ( .A1(n2946), .A2(n2945), .A3(REG0_REG_18__SCAN_IN), .A4(
        ADDR_REG_6__SCAN_IN), .ZN(n2956) );
  INV_X1 U3831 ( .A(DATAI_12_), .ZN(n2947) );
  NAND4_X1 U3832 ( .A1(n2948), .A2(n2947), .A3(DATAI_4_), .A4(DATAI_6_), .ZN(
        n2954) );
  INV_X1 U3833 ( .A(DATAO_REG_23__SCAN_IN), .ZN(n3400) );
  NAND4_X1 U3834 ( .A1(REG3_REG_11__SCAN_IN), .A2(ADDR_REG_10__SCAN_IN), .A3(
        n2543), .A4(n3400), .ZN(n2950) );
  NAND4_X1 U3835 ( .A1(REG1_REG_26__SCAN_IN), .A2(IR_REG_28__SCAN_IN), .A3(
        n3068), .A4(n2586), .ZN(n2949) );
  NOR2_X1 U3836 ( .A1(n2950), .A2(n2949), .ZN(n2952) );
  NOR4_X1 U3837 ( .A1(IR_REG_21__SCAN_IN), .A2(n2222), .A3(
        REG0_REG_13__SCAN_IN), .A4(n3090), .ZN(n2951) );
  NAND4_X1 U3838 ( .A1(IR_REG_25__SCAN_IN), .A2(n2952), .A3(n2951), .A4(
        REG3_REG_9__SCAN_IN), .ZN(n2953) );
  NOR4_X1 U3839 ( .A1(n2954), .A2(n2953), .A3(n3079), .A4(REG0_REG_27__SCAN_IN), .ZN(n2955) );
  AND4_X1 U3840 ( .A1(n2958), .A2(n2957), .A3(n2956), .A4(n2955), .ZN(n2959)
         );
  AOI21_X1 U3841 ( .B1(n2960), .B2(n2959), .A(DATAO_REG_19__SCAN_IN), .ZN(
        n3158) );
  AOI22_X1 U3842 ( .A1(n3495), .A2(keyinput35), .B1(n2935), .B2(keyinput55), 
        .ZN(n2961) );
  OAI221_X1 U3843 ( .B1(n3495), .B2(keyinput35), .C1(n2935), .C2(keyinput55), 
        .A(n2961), .ZN(n2970) );
  INV_X1 U3844 ( .A(D_REG_14__SCAN_IN), .ZN(n4971) );
  INV_X1 U3845 ( .A(REG3_REG_20__SCAN_IN), .ZN(n2963) );
  AOI22_X1 U3846 ( .A1(n4971), .A2(keyinput29), .B1(keyinput95), .B2(n2963), 
        .ZN(n2962) );
  OAI221_X1 U3847 ( .B1(n4971), .B2(keyinput29), .C1(n2963), .C2(keyinput95), 
        .A(n2962), .ZN(n2969) );
  INV_X1 U3848 ( .A(REG0_REG_31__SCAN_IN), .ZN(n3254) );
  AOI22_X1 U3849 ( .A1(n3920), .A2(keyinput67), .B1(keyinput43), .B2(n3254), 
        .ZN(n2964) );
  OAI221_X1 U3850 ( .B1(n3920), .B2(keyinput67), .C1(n3254), .C2(keyinput43), 
        .A(n2964), .ZN(n2968) );
  XOR2_X1 U3851 ( .A(n2641), .B(keyinput59), .Z(n2966) );
  XNOR2_X1 U3852 ( .A(IR_REG_13__SCAN_IN), .B(keyinput79), .ZN(n2965) );
  NAND2_X1 U3853 ( .A1(n2966), .A2(n2965), .ZN(n2967) );
  NOR4_X1 U3854 ( .A1(n2970), .A2(n2969), .A3(n2968), .A4(n2967), .ZN(n3004)
         );
  INV_X1 U3855 ( .A(ADDR_REG_7__SCAN_IN), .ZN(n2972) );
  AOI22_X1 U3856 ( .A1(n3868), .A2(keyinput87), .B1(keyinput91), .B2(n2972), 
        .ZN(n2971) );
  OAI221_X1 U3857 ( .B1(n3868), .B2(keyinput87), .C1(n2972), .C2(keyinput91), 
        .A(n2971), .ZN(n2982) );
  INV_X1 U3858 ( .A(REG2_REG_18__SCAN_IN), .ZN(n2974) );
  AOI22_X1 U3859 ( .A1(n3280), .A2(keyinput103), .B1(n2974), .B2(keyinput75), 
        .ZN(n2973) );
  OAI221_X1 U3860 ( .B1(n3280), .B2(keyinput103), .C1(n2974), .C2(keyinput75), 
        .A(n2973), .ZN(n2981) );
  INV_X1 U3861 ( .A(REG2_REG_31__SCAN_IN), .ZN(n2976) );
  AOI22_X1 U3862 ( .A1(n4799), .A2(keyinput123), .B1(keyinput107), .B2(n2976), 
        .ZN(n2975) );
  OAI221_X1 U3863 ( .B1(n4799), .B2(keyinput123), .C1(n2976), .C2(keyinput107), 
        .A(n2975), .ZN(n2980) );
  XNOR2_X1 U3864 ( .A(IR_REG_9__SCAN_IN), .B(keyinput51), .ZN(n2978) );
  XNOR2_X1 U3865 ( .A(DATAI_22_), .B(keyinput115), .ZN(n2977) );
  NAND2_X1 U3866 ( .A1(n2978), .A2(n2977), .ZN(n2979) );
  NOR4_X1 U3867 ( .A1(n2982), .A2(n2981), .A3(n2980), .A4(n2979), .ZN(n3003)
         );
  AOI22_X1 U3868 ( .A1(n2570), .A2(keyinput111), .B1(keyinput127), .B2(n4830), 
        .ZN(n2983) );
  OAI221_X1 U3869 ( .B1(n2570), .B2(keyinput111), .C1(n4830), .C2(keyinput127), 
        .A(n2983), .ZN(n2990) );
  INV_X1 U3870 ( .A(D_REG_20__SCAN_IN), .ZN(n4967) );
  AOI22_X1 U3871 ( .A1(n4967), .A2(keyinput119), .B1(keyinput63), .B2(n4733), 
        .ZN(n2984) );
  OAI221_X1 U3872 ( .B1(n4967), .B2(keyinput119), .C1(n4733), .C2(keyinput63), 
        .A(n2984), .ZN(n2989) );
  INV_X1 U3873 ( .A(D_REG_28__SCAN_IN), .ZN(n4962) );
  AOI22_X1 U3874 ( .A1(n2522), .A2(keyinput31), .B1(n4962), .B2(keyinput83), 
        .ZN(n2985) );
  OAI221_X1 U3875 ( .B1(n2522), .B2(keyinput31), .C1(n4962), .C2(keyinput83), 
        .A(n2985), .ZN(n2988) );
  INV_X1 U3876 ( .A(D_REG_26__SCAN_IN), .ZN(n4963) );
  INV_X1 U3877 ( .A(D_REG_17__SCAN_IN), .ZN(n4970) );
  AOI22_X1 U3878 ( .A1(n4963), .A2(keyinput3), .B1(keyinput99), .B2(n4970), 
        .ZN(n2986) );
  OAI221_X1 U3879 ( .B1(n4963), .B2(keyinput3), .C1(n4970), .C2(keyinput99), 
        .A(n2986), .ZN(n2987) );
  NOR4_X1 U3880 ( .A1(n2990), .A2(n2989), .A3(n2988), .A4(n2987), .ZN(n3002)
         );
  INV_X1 U3881 ( .A(D_REG_29__SCAN_IN), .ZN(n4961) );
  AOI22_X1 U3882 ( .A1(n4961), .A2(keyinput71), .B1(keyinput19), .B2(n4866), 
        .ZN(n2991) );
  OAI221_X1 U3883 ( .B1(n4961), .B2(keyinput71), .C1(n4866), .C2(keyinput19), 
        .A(n2991), .ZN(n3000) );
  INV_X1 U3884 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n3247) );
  AOI22_X1 U3885 ( .A1(n3247), .A2(keyinput27), .B1(n2993), .B2(keyinput39), 
        .ZN(n2992) );
  OAI221_X1 U3886 ( .B1(n3247), .B2(keyinput27), .C1(n2993), .C2(keyinput39), 
        .A(n2992), .ZN(n2999) );
  INV_X1 U3887 ( .A(REG2_REG_26__SCAN_IN), .ZN(n2995) );
  AOI22_X1 U3888 ( .A1(n3867), .A2(keyinput47), .B1(keyinput7), .B2(n2995), 
        .ZN(n2994) );
  OAI221_X1 U3889 ( .B1(n3867), .B2(keyinput47), .C1(n2995), .C2(keyinput7), 
        .A(n2994), .ZN(n2998) );
  INV_X1 U3890 ( .A(REG3_REG_5__SCAN_IN), .ZN(n3240) );
  INV_X1 U3891 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n3251) );
  AOI22_X1 U3892 ( .A1(n3240), .A2(keyinput15), .B1(keyinput11), .B2(n3251), 
        .ZN(n2996) );
  OAI221_X1 U3893 ( .B1(n3240), .B2(keyinput15), .C1(n3251), .C2(keyinput11), 
        .A(n2996), .ZN(n2997) );
  NOR4_X1 U3894 ( .A1(n3000), .A2(n2999), .A3(n2998), .A4(n2997), .ZN(n3001)
         );
  NAND4_X1 U3895 ( .A1(n3004), .A2(n3003), .A3(n3002), .A4(n3001), .ZN(n3156)
         );
  INV_X1 U3896 ( .A(DATAI_20_), .ZN(n3006) );
  INV_X1 U3897 ( .A(REG3_REG_25__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U3898 ( .A1(n3006), .A2(keyinput23), .B1(n3977), .B2(keyinput52), 
        .ZN(n3005) );
  OAI221_X1 U3899 ( .B1(n3006), .B2(keyinput23), .C1(n3977), .C2(keyinput52), 
        .A(n3005), .ZN(n3017) );
  INV_X1 U3900 ( .A(ADDR_REG_19__SCAN_IN), .ZN(n3009) );
  AOI22_X1 U3901 ( .A1(n3009), .A2(keyinput60), .B1(keyinput80), .B2(n3008), 
        .ZN(n3007) );
  OAI221_X1 U3902 ( .B1(n3009), .B2(keyinput60), .C1(n3008), .C2(keyinput80), 
        .A(n3007), .ZN(n3016) );
  AOI22_X1 U3903 ( .A1(n4012), .A2(keyinput46), .B1(keyinput73), .B2(n4920), 
        .ZN(n3010) );
  OAI221_X1 U3904 ( .B1(n4012), .B2(keyinput46), .C1(n4920), .C2(keyinput73), 
        .A(n3010), .ZN(n3015) );
  INV_X1 U3905 ( .A(ADDR_REG_1__SCAN_IN), .ZN(n3012) );
  AOI22_X1 U3906 ( .A1(n3013), .A2(keyinput78), .B1(keyinput72), .B2(n3012), 
        .ZN(n3011) );
  OAI221_X1 U3907 ( .B1(n3013), .B2(keyinput78), .C1(n3012), .C2(keyinput72), 
        .A(n3011), .ZN(n3014) );
  NOR4_X1 U3908 ( .A1(n3017), .A2(n3016), .A3(n3015), .A4(n3014), .ZN(n3054)
         );
  INV_X1 U3909 ( .A(ADDR_REG_4__SCAN_IN), .ZN(n3020) );
  AOI22_X1 U3910 ( .A1(n3020), .A2(keyinput58), .B1(n3019), .B2(keyinput42), 
        .ZN(n3018) );
  OAI221_X1 U3911 ( .B1(n3020), .B2(keyinput58), .C1(n3019), .C2(keyinput42), 
        .A(n3018), .ZN(n3029) );
  INV_X1 U3912 ( .A(ADDR_REG_16__SCAN_IN), .ZN(n3022) );
  AOI22_X1 U3913 ( .A1(n3022), .A2(keyinput64), .B1(n3446), .B2(keyinput53), 
        .ZN(n3021) );
  OAI221_X1 U3914 ( .B1(n3022), .B2(keyinput64), .C1(n3446), .C2(keyinput53), 
        .A(n3021), .ZN(n3028) );
  AOI22_X1 U3915 ( .A1(n3024), .A2(keyinput68), .B1(keyinput85), .B2(n2544), 
        .ZN(n3023) );
  OAI221_X1 U3916 ( .B1(n3024), .B2(keyinput68), .C1(n2544), .C2(keyinput85), 
        .A(n3023), .ZN(n3027) );
  AOI22_X1 U3917 ( .A1(n2519), .A2(keyinput45), .B1(n2558), .B2(keyinput69), 
        .ZN(n3025) );
  OAI221_X1 U3918 ( .B1(n2519), .B2(keyinput45), .C1(n2558), .C2(keyinput69), 
        .A(n3025), .ZN(n3026) );
  NOR4_X1 U3919 ( .A1(n3029), .A2(n3028), .A3(n3027), .A4(n3026), .ZN(n3053)
         );
  INV_X1 U3920 ( .A(D_REG_4__SCAN_IN), .ZN(n4974) );
  INV_X1 U3921 ( .A(D_REG_8__SCAN_IN), .ZN(n4973) );
  AOI22_X1 U3922 ( .A1(n4974), .A2(keyinput56), .B1(keyinput44), .B2(n4973), 
        .ZN(n3030) );
  OAI221_X1 U3923 ( .B1(n4974), .B2(keyinput56), .C1(n4973), .C2(keyinput44), 
        .A(n3030), .ZN(n3040) );
  AOI22_X1 U3924 ( .A1(n3033), .A2(keyinput65), .B1(n3032), .B2(keyinput70), 
        .ZN(n3031) );
  OAI221_X1 U3925 ( .B1(n3033), .B2(keyinput65), .C1(n3032), .C2(keyinput70), 
        .A(n3031), .ZN(n3039) );
  INV_X1 U3926 ( .A(D_REG_30__SCAN_IN), .ZN(n4960) );
  XOR2_X1 U3927 ( .A(n4960), .B(keyinput61), .Z(n3037) );
  XNOR2_X1 U3928 ( .A(IR_REG_5__SCAN_IN), .B(keyinput66), .ZN(n3036) );
  XNOR2_X1 U3929 ( .A(IR_REG_7__SCAN_IN), .B(keyinput76), .ZN(n3035) );
  XNOR2_X1 U3930 ( .A(IR_REG_8__SCAN_IN), .B(keyinput50), .ZN(n3034) );
  NAND4_X1 U3931 ( .A1(n3037), .A2(n3036), .A3(n3035), .A4(n3034), .ZN(n3038)
         );
  NOR3_X1 U3932 ( .A1(n3040), .A2(n3039), .A3(n3038), .ZN(n3052) );
  AOI22_X1 U3933 ( .A1(n3266), .A2(keyinput57), .B1(n3163), .B2(keyinput54), 
        .ZN(n3041) );
  OAI221_X1 U3934 ( .B1(n3266), .B2(keyinput57), .C1(n3163), .C2(keyinput54), 
        .A(n3041), .ZN(n3045) );
  XNOR2_X1 U3935 ( .A(n3042), .B(keyinput74), .ZN(n3044) );
  INV_X1 U3936 ( .A(DATAO_REG_2__SCAN_IN), .ZN(n3714) );
  XNOR2_X1 U3937 ( .A(n3714), .B(keyinput81), .ZN(n3043) );
  OR3_X1 U3938 ( .A1(n3045), .A2(n3044), .A3(n3043), .ZN(n3050) );
  AOI22_X1 U3939 ( .A1(n3258), .A2(keyinput49), .B1(n4959), .B2(keyinput62), 
        .ZN(n3046) );
  OAI221_X1 U3940 ( .B1(n3258), .B2(keyinput49), .C1(n4959), .C2(keyinput62), 
        .A(n3046), .ZN(n3049) );
  AOI22_X1 U3941 ( .A1(n2478), .A2(keyinput77), .B1(n4968), .B2(keyinput82), 
        .ZN(n3047) );
  OAI221_X1 U3942 ( .B1(n2478), .B2(keyinput77), .C1(n4968), .C2(keyinput82), 
        .A(n3047), .ZN(n3048) );
  NOR3_X1 U3943 ( .A1(n3050), .A2(n3049), .A3(n3048), .ZN(n3051) );
  NAND4_X1 U3944 ( .A1(n3054), .A2(n3053), .A3(n3052), .A4(n3051), .ZN(n3155)
         );
  AOI22_X1 U3945 ( .A1(n4964), .A2(keyinput9), .B1(keyinput6), .B2(n3056), 
        .ZN(n3055) );
  OAI221_X1 U3946 ( .B1(n4964), .B2(keyinput9), .C1(n3056), .C2(keyinput6), 
        .A(n3055), .ZN(n3066) );
  INV_X1 U3947 ( .A(ADDR_REG_5__SCAN_IN), .ZN(n3058) );
  AOI22_X1 U3948 ( .A1(n4969), .A2(keyinput5), .B1(keyinput0), .B2(n3058), 
        .ZN(n3057) );
  OAI221_X1 U3949 ( .B1(n4969), .B2(keyinput5), .C1(n3058), .C2(keyinput0), 
        .A(n3057), .ZN(n3065) );
  AOI22_X1 U3950 ( .A1(n2585), .A2(keyinput1), .B1(n3060), .B2(keyinput8), 
        .ZN(n3059) );
  OAI221_X1 U3951 ( .B1(n2585), .B2(keyinput1), .C1(n3060), .C2(keyinput8), 
        .A(n3059), .ZN(n3064) );
  XNOR2_X1 U3952 ( .A(REG2_REG_2__SCAN_IN), .B(keyinput2), .ZN(n3062) );
  XNOR2_X1 U3953 ( .A(REG0_REG_18__SCAN_IN), .B(keyinput17), .ZN(n3061) );
  NAND2_X1 U3954 ( .A1(n3062), .A2(n3061), .ZN(n3063) );
  NOR4_X1 U3955 ( .A1(n3066), .A2(n3065), .A3(n3064), .A4(n3063), .ZN(n3104)
         );
  AOI22_X1 U3956 ( .A1(n2586), .A2(keyinput14), .B1(n3068), .B2(keyinput10), 
        .ZN(n3067) );
  OAI221_X1 U3957 ( .B1(n2586), .B2(keyinput14), .C1(n3068), .C2(keyinput10), 
        .A(n3067), .ZN(n3077) );
  INV_X1 U3958 ( .A(ADDR_REG_10__SCAN_IN), .ZN(n3070) );
  AOI22_X1 U3959 ( .A1(n2924), .A2(keyinput126), .B1(keyinput12), .B2(n3070), 
        .ZN(n3069) );
  OAI221_X1 U3960 ( .B1(n2924), .B2(keyinput126), .C1(n3070), .C2(keyinput12), 
        .A(n3069), .ZN(n3076) );
  XNOR2_X1 U3961 ( .A(IR_REG_25__SCAN_IN), .B(keyinput18), .ZN(n3074) );
  XNOR2_X1 U3962 ( .A(IR_REG_28__SCAN_IN), .B(keyinput21), .ZN(n3073) );
  XNOR2_X1 U3963 ( .A(REG1_REG_26__SCAN_IN), .B(keyinput13), .ZN(n3072) );
  XNOR2_X1 U3964 ( .A(keyinput16), .B(REG3_REG_9__SCAN_IN), .ZN(n3071) );
  NAND4_X1 U3965 ( .A1(n3074), .A2(n3073), .A3(n3072), .A4(n3071), .ZN(n3075)
         );
  NOR3_X1 U3966 ( .A1(n3077), .A2(n3076), .A3(n3075), .ZN(n3103) );
  AOI22_X1 U3967 ( .A1(n2948), .A2(keyinput38), .B1(n3079), .B2(keyinput24), 
        .ZN(n3078) );
  OAI221_X1 U3968 ( .B1(n2948), .B2(keyinput38), .C1(n3079), .C2(keyinput24), 
        .A(n3078), .ZN(n3088) );
  XNOR2_X1 U3969 ( .A(n3080), .B(keyinput20), .ZN(n3087) );
  XNOR2_X1 U3970 ( .A(DATAI_6_), .B(keyinput25), .ZN(n3084) );
  XNOR2_X1 U3971 ( .A(DATAI_12_), .B(keyinput22), .ZN(n3083) );
  XNOR2_X1 U3972 ( .A(DATAI_3_), .B(keyinput30), .ZN(n3082) );
  XNOR2_X1 U3973 ( .A(DATAI_4_), .B(keyinput28), .ZN(n3081) );
  NAND4_X1 U3974 ( .A1(n3084), .A2(n3083), .A3(n3082), .A4(n3081), .ZN(n3086)
         );
  XNOR2_X1 U3975 ( .A(keyinput26), .B(n2534), .ZN(n3085) );
  NOR4_X1 U3976 ( .A1(n3088), .A2(n3087), .A3(n3086), .A4(n3085), .ZN(n3102)
         );
  AOI22_X1 U3977 ( .A1(n4835), .A2(keyinput34), .B1(n3090), .B2(keyinput32), 
        .ZN(n3089) );
  OAI221_X1 U3978 ( .B1(n4835), .B2(keyinput34), .C1(n3090), .C2(keyinput32), 
        .A(n3089), .ZN(n3100) );
  AOI22_X1 U3979 ( .A1(n2843), .A2(keyinput4), .B1(keyinput37), .B2(n3092), 
        .ZN(n3091) );
  OAI221_X1 U3980 ( .B1(n2843), .B2(keyinput4), .C1(n3092), .C2(keyinput37), 
        .A(n3091), .ZN(n3099) );
  INV_X1 U3981 ( .A(ADDR_REG_6__SCAN_IN), .ZN(n3094) );
  AOI22_X1 U3982 ( .A1(n4858), .A2(keyinput41), .B1(keyinput36), .B2(n3094), 
        .ZN(n3093) );
  OAI221_X1 U3983 ( .B1(n4858), .B2(keyinput41), .C1(n3094), .C2(keyinput36), 
        .A(n3093), .ZN(n3098) );
  AOI22_X1 U3984 ( .A1(n3096), .A2(keyinput33), .B1(keyinput40), .B2(n2303), 
        .ZN(n3095) );
  OAI221_X1 U3985 ( .B1(n3096), .B2(keyinput33), .C1(n2303), .C2(keyinput40), 
        .A(n3095), .ZN(n3097) );
  NOR4_X1 U3986 ( .A1(n3100), .A2(n3099), .A3(n3098), .A4(n3097), .ZN(n3101)
         );
  NAND4_X1 U3987 ( .A1(n3104), .A2(n3103), .A3(n3102), .A4(n3101), .ZN(n3154)
         );
  INV_X1 U3988 ( .A(D_REG_1__SCAN_IN), .ZN(n3165) );
  INV_X1 U3989 ( .A(DATAI_26_), .ZN(n3106) );
  AOI22_X1 U3990 ( .A1(n3165), .A2(keyinput92), .B1(keyinput96), .B2(n3106), 
        .ZN(n3105) );
  OAI221_X1 U3991 ( .B1(n3165), .B2(keyinput92), .C1(n3106), .C2(keyinput96), 
        .A(n3105), .ZN(n3116) );
  INV_X1 U3992 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3109) );
  INV_X1 U3993 ( .A(REG2_REG_20__SCAN_IN), .ZN(n3108) );
  AOI22_X1 U3994 ( .A1(n3109), .A2(keyinput97), .B1(n3108), .B2(keyinput98), 
        .ZN(n3107) );
  OAI221_X1 U3995 ( .B1(n3109), .B2(keyinput97), .C1(n3108), .C2(keyinput98), 
        .A(n3107), .ZN(n3115) );
  INV_X1 U3996 ( .A(DATAO_REG_12__SCAN_IN), .ZN(n3249) );
  AOI22_X1 U3997 ( .A1(n3249), .A2(keyinput100), .B1(n4854), .B2(keyinput104), 
        .ZN(n3110) );
  OAI221_X1 U3998 ( .B1(n3249), .B2(keyinput100), .C1(n4854), .C2(keyinput104), 
        .A(n3110), .ZN(n3114) );
  XOR2_X1 U3999 ( .A(n2925), .B(keyinput102), .Z(n3112) );
  XNOR2_X1 U4000 ( .A(IR_REG_17__SCAN_IN), .B(keyinput101), .ZN(n3111) );
  NAND2_X1 U4001 ( .A1(n3112), .A2(n3111), .ZN(n3113) );
  NOR4_X1 U4002 ( .A1(n3116), .A2(n3115), .A3(n3114), .A4(n3113), .ZN(n3152)
         );
  INV_X1 U4003 ( .A(D_REG_2__SCAN_IN), .ZN(n4976) );
  AOI22_X1 U4004 ( .A1(n3118), .A2(keyinput93), .B1(n4976), .B2(keyinput94), 
        .ZN(n3117) );
  OAI221_X1 U4005 ( .B1(n3118), .B2(keyinput93), .C1(n4976), .C2(keyinput94), 
        .A(n3117), .ZN(n3126) );
  INV_X1 U4006 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3586) );
  AOI22_X1 U4007 ( .A1(n2716), .A2(keyinput86), .B1(keyinput84), .B2(n3586), 
        .ZN(n3119) );
  OAI221_X1 U4008 ( .B1(n2716), .B2(keyinput86), .C1(n3586), .C2(keyinput84), 
        .A(n3119), .ZN(n3125) );
  INV_X1 U4009 ( .A(DATAO_REG_19__SCAN_IN), .ZN(n3278) );
  AOI22_X1 U4010 ( .A1(keyinput89), .A2(n4792), .B1(keyinput48), .B2(n3278), 
        .ZN(n3120) );
  OAI21_X1 U4011 ( .B1(n4792), .B2(keyinput89), .A(n3120), .ZN(n3124) );
  XOR2_X1 U4012 ( .A(n2528), .B(keyinput90), .Z(n3122) );
  XNOR2_X1 U4013 ( .A(DATAI_7_), .B(keyinput88), .ZN(n3121) );
  NAND2_X1 U4014 ( .A1(n3122), .A2(n3121), .ZN(n3123) );
  NOR4_X1 U4015 ( .A1(n3126), .A2(n3125), .A3(n3124), .A4(n3123), .ZN(n3151)
         );
  AOI22_X1 U4016 ( .A1(n4778), .A2(keyinput116), .B1(keyinput121), .B2(n2510), 
        .ZN(n3127) );
  OAI221_X1 U4017 ( .B1(n4778), .B2(keyinput116), .C1(n2510), .C2(keyinput121), 
        .A(n3127), .ZN(n3136) );
  AOI22_X1 U4018 ( .A1(n3264), .A2(keyinput114), .B1(n3129), .B2(keyinput118), 
        .ZN(n3128) );
  OAI221_X1 U4019 ( .B1(n3264), .B2(keyinput114), .C1(n3129), .C2(keyinput118), 
        .A(n3128), .ZN(n3135) );
  INV_X1 U4020 ( .A(REG3_REG_11__SCAN_IN), .ZN(n3131) );
  AOI22_X1 U4021 ( .A1(n3400), .A2(keyinput122), .B1(n3131), .B2(keyinput124), 
        .ZN(n3130) );
  OAI221_X1 U4022 ( .B1(n3400), .B2(keyinput122), .C1(n3131), .C2(keyinput124), 
        .A(n3130), .ZN(n3134) );
  AOI22_X1 U4023 ( .A1(n3253), .A2(keyinput120), .B1(n2543), .B2(keyinput125), 
        .ZN(n3132) );
  OAI221_X1 U4024 ( .B1(n3253), .B2(keyinput120), .C1(n2543), .C2(keyinput125), 
        .A(n3132), .ZN(n3133) );
  NOR4_X1 U4025 ( .A1(n3136), .A2(n3135), .A3(n3134), .A4(n3133), .ZN(n3150)
         );
  INV_X1 U4026 ( .A(ADDR_REG_14__SCAN_IN), .ZN(n3699) );
  INV_X1 U4027 ( .A(ADDR_REG_11__SCAN_IN), .ZN(n3138) );
  AOI22_X1 U4028 ( .A1(n3699), .A2(keyinput113), .B1(keyinput117), .B2(n3138), 
        .ZN(n3137) );
  OAI221_X1 U4029 ( .B1(n3699), .B2(keyinput113), .C1(n3138), .C2(keyinput117), 
        .A(n3137), .ZN(n3148) );
  INV_X1 U4030 ( .A(D_REG_11__SCAN_IN), .ZN(n4972) );
  AOI22_X1 U4031 ( .A1(n4972), .A2(keyinput105), .B1(keyinput106), .B2(n4965), 
        .ZN(n3139) );
  OAI221_X1 U4032 ( .B1(n4972), .B2(keyinput105), .C1(n4965), .C2(keyinput106), 
        .A(n3139), .ZN(n3147) );
  AOI22_X1 U4033 ( .A1(n4355), .A2(keyinput110), .B1(n3141), .B2(keyinput112), 
        .ZN(n3140) );
  OAI221_X1 U4034 ( .B1(n4355), .B2(keyinput110), .C1(n3141), .C2(keyinput112), 
        .A(n3140), .ZN(n3146) );
  INV_X1 U4035 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3142) );
  XOR2_X1 U4036 ( .A(n3142), .B(keyinput108), .Z(n3144) );
  XNOR2_X1 U4037 ( .A(REG3_REG_6__SCAN_IN), .B(keyinput109), .ZN(n3143) );
  NAND2_X1 U4038 ( .A1(n3144), .A2(n3143), .ZN(n3145) );
  NOR4_X1 U4039 ( .A1(n3148), .A2(n3147), .A3(n3146), .A4(n3145), .ZN(n3149)
         );
  NAND4_X1 U4040 ( .A1(n3152), .A2(n3151), .A3(n3150), .A4(n3149), .ZN(n3153)
         );
  NOR4_X1 U4041 ( .A1(n3156), .A2(n3155), .A3(n3154), .A4(n3153), .ZN(n3157)
         );
  OAI21_X1 U4042 ( .B1(n3158), .B2(keyinput48), .A(n3157), .ZN(n3160) );
  MUX2_X1 U40430 ( .A(n3170), .B(DATAI_1_), .S(U3149), .Z(n3159) );
  XNOR2_X1 U4044 ( .A(n3160), .B(n3159), .ZN(U3351) );
  INV_X1 U4045 ( .A(n3161), .ZN(n3162) );
  AOI22_X1 U4046 ( .A1(n4975), .A2(n3163), .B1(n3162), .B2(n4978), .ZN(U3458)
         );
  INV_X1 U4047 ( .A(n3324), .ZN(n3164) );
  AOI22_X1 U4048 ( .A1(n4975), .A2(n3165), .B1(n3164), .B2(n4978), .ZN(U3459)
         );
  INV_X1 U4049 ( .A(n3368), .ZN(n3166) );
  NAND2_X1 U4050 ( .A1(n3166), .A2(STATE_REG_SCAN_IN), .ZN(n4274) );
  NAND2_X1 U4051 ( .A1(n3403), .A2(n4274), .ZN(n3183) );
  NAND2_X1 U4052 ( .A1(n3167), .A2(n3368), .ZN(n3168) );
  AND2_X1 U4053 ( .A1(n3168), .A2(n2144), .ZN(n3181) );
  INV_X1 U4054 ( .A(n4343), .ZN(n4289) );
  INV_X1 U4055 ( .A(REG1_REG_2__SCAN_IN), .ZN(n3169) );
  AND2_X1 U4056 ( .A1(n2222), .A2(REG1_REG_0__SCAN_IN), .ZN(n3268) );
  NAND2_X1 U4057 ( .A1(n3170), .A2(REG1_REG_1__SCAN_IN), .ZN(n3171) );
  NAND2_X1 U4058 ( .A1(n3172), .A2(n3171), .ZN(n4298) );
  NAND2_X1 U4059 ( .A1(n2521), .A2(REG1_REG_2__SCAN_IN), .ZN(n3173) );
  XOR2_X1 U4060 ( .A(n3187), .B(REG1_REG_3__SCAN_IN), .Z(n3180) );
  AND2_X1 U4061 ( .A1(n4287), .A2(n4343), .ZN(n4270) );
  INV_X1 U4062 ( .A(REG2_REG_1__SCAN_IN), .ZN(n3270) );
  NAND2_X1 U4063 ( .A1(n2222), .A2(REG2_REG_0__SCAN_IN), .ZN(n3269) );
  OR2_X1 U4064 ( .A1(n3175), .A2(n3270), .ZN(n3177) );
  NAND2_X1 U4065 ( .A1(n2521), .A2(REG2_REG_2__SCAN_IN), .ZN(n3178) );
  XOR2_X1 U4066 ( .A(n3193), .B(REG2_REG_3__SCAN_IN), .Z(n3179) );
  AOI22_X1 U4067 ( .A1(n4935), .A2(n3180), .B1(n4948), .B2(n3179), .ZN(n3185)
         );
  INV_X1 U4068 ( .A(n3181), .ZN(n3182) );
  NOR2_X1 U4069 ( .A1(STATE_REG_SCAN_IN), .A2(n2543), .ZN(n3374) );
  AOI21_X1 U4070 ( .B1(n4942), .B2(ADDR_REG_3__SCAN_IN), .A(n3374), .ZN(n3184)
         );
  OAI211_X1 U4071 ( .C1(n3186), .C2(n4949), .A(n3185), .B(n3184), .ZN(U3243)
         );
  NAND2_X1 U4072 ( .A1(n3187), .A2(REG1_REG_3__SCAN_IN), .ZN(n3190) );
  NAND2_X1 U4073 ( .A1(n3188), .A2(n4886), .ZN(n3189) );
  INV_X1 U4074 ( .A(n4896), .ZN(n3197) );
  MUX2_X1 U4075 ( .A(n2586), .B(REG1_REG_5__SCAN_IN), .S(n3201), .Z(n3235) );
  NOR2_X2 U4076 ( .A1(n3236), .A2(n3235), .ZN(n3234) );
  NOR2_X2 U4077 ( .A1(n3234), .A2(n3192), .ZN(n3209) );
  XNOR2_X1 U4078 ( .A(n3211), .B(REG1_REG_6__SCAN_IN), .ZN(n3208) );
  NAND2_X1 U4079 ( .A1(n3193), .A2(REG2_REG_3__SCAN_IN), .ZN(n3196) );
  NAND2_X1 U4080 ( .A1(n3194), .A2(n4886), .ZN(n3195) );
  NAND2_X1 U4081 ( .A1(n4893), .A2(REG2_REG_4__SCAN_IN), .ZN(n3200) );
  NAND2_X1 U4082 ( .A1(n3198), .A2(n3197), .ZN(n3199) );
  NAND2_X1 U4083 ( .A1(n3200), .A2(n3199), .ZN(n3238) );
  MUX2_X1 U4084 ( .A(REG2_REG_5__SCAN_IN), .B(n3586), .S(n3201), .Z(n3239) );
  NAND2_X1 U4085 ( .A1(n3238), .A2(n3239), .ZN(n3237) );
  NAND2_X1 U4086 ( .A1(n3201), .A2(REG2_REG_5__SCAN_IN), .ZN(n3202) );
  INV_X1 U4087 ( .A(n4885), .ZN(n3204) );
  XOR2_X1 U4088 ( .A(n3214), .B(REG2_REG_6__SCAN_IN), .Z(n3206) );
  AND2_X1 U4089 ( .A1(U3149), .A2(REG3_REG_6__SCAN_IN), .ZN(n3475) );
  AOI21_X1 U4090 ( .B1(n4942), .B2(ADDR_REG_6__SCAN_IN), .A(n3475), .ZN(n3203)
         );
  OAI21_X1 U4091 ( .B1(n4949), .B2(n3204), .A(n3203), .ZN(n3205) );
  AOI21_X1 U4092 ( .B1(n3206), .B2(n4948), .A(n3205), .ZN(n3207) );
  OAI21_X1 U4093 ( .B1(n3208), .B2(n4938), .A(n3207), .ZN(U3246) );
  INV_X1 U4094 ( .A(n3209), .ZN(n3210) );
  MUX2_X1 U4095 ( .A(REG1_REG_7__SCAN_IN), .B(n3298), .S(n3299), .Z(n3212) );
  XNOR2_X1 U4096 ( .A(n3297), .B(n3212), .ZN(n3224) );
  AND2_X1 U4097 ( .A1(REG3_REG_7__SCAN_IN), .A2(U3149), .ZN(n3491) );
  NOR2_X1 U4098 ( .A1(n4949), .A2(n3299), .ZN(n3213) );
  AOI211_X1 U4099 ( .C1(n4942), .C2(ADDR_REG_7__SCAN_IN), .A(n3491), .B(n3213), 
        .ZN(n3223) );
  NAND2_X1 U4100 ( .A1(n3214), .A2(REG2_REG_6__SCAN_IN), .ZN(n3217) );
  NAND2_X1 U4101 ( .A1(n3215), .A2(n4885), .ZN(n3216) );
  INV_X1 U4102 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3601) );
  MUX2_X1 U4103 ( .A(REG2_REG_7__SCAN_IN), .B(n3601), .S(n3299), .Z(n3218) );
  INV_X1 U4104 ( .A(n3218), .ZN(n3220) );
  MUX2_X1 U4105 ( .A(n3601), .B(REG2_REG_7__SCAN_IN), .S(n3299), .Z(n3219) );
  NAND2_X1 U4106 ( .A1(n3221), .A2(n3219), .ZN(n3296) );
  OAI211_X1 U4107 ( .C1(n3221), .C2(n3220), .A(n3296), .B(n4948), .ZN(n3222)
         );
  OAI211_X1 U4108 ( .C1(n3224), .C2(n4938), .A(n3223), .B(n3222), .ZN(U3247)
         );
  INV_X1 U4109 ( .A(n3225), .ZN(n3230) );
  INV_X1 U4110 ( .A(REG2_REG_0__SCAN_IN), .ZN(n3226) );
  AOI21_X1 U4111 ( .B1(n4343), .B2(n3226), .A(n4888), .ZN(n4292) );
  OAI21_X1 U4112 ( .B1(REG1_REG_0__SCAN_IN), .B2(n4343), .A(n4292), .ZN(n3227)
         );
  MUX2_X1 U4113 ( .A(n3227), .B(n4292), .S(n2222), .Z(n3229) );
  INV_X1 U4114 ( .A(REG3_REG_0__SCAN_IN), .ZN(n3228) );
  OAI22_X1 U4115 ( .A1(n3230), .A2(n3229), .B1(STATE_REG_SCAN_IN), .B2(n3228), 
        .ZN(n3232) );
  NOR3_X1 U4116 ( .A1(n4938), .A2(REG1_REG_0__SCAN_IN), .A3(n2303), .ZN(n3231)
         );
  AOI211_X1 U4117 ( .C1(n4942), .C2(ADDR_REG_0__SCAN_IN), .A(n3232), .B(n3231), 
        .ZN(n3233) );
  INV_X1 U4118 ( .A(n3233), .ZN(U3240) );
  NOR2_X1 U4119 ( .A1(n4942), .A2(U4043), .ZN(U3148) );
  AOI211_X1 U4120 ( .C1(n3236), .C2(n3235), .A(n3234), .B(n4938), .ZN(n3245)
         );
  OAI211_X1 U4121 ( .C1(n3239), .C2(n3238), .A(n4948), .B(n3237), .ZN(n3242)
         );
  NOR2_X1 U4122 ( .A1(STATE_REG_SCAN_IN), .A2(n3240), .ZN(n3429) );
  AOI21_X1 U4123 ( .B1(n4942), .B2(ADDR_REG_5__SCAN_IN), .A(n3429), .ZN(n3241)
         );
  OAI211_X1 U4124 ( .C1(n4949), .C2(n3243), .A(n3242), .B(n3241), .ZN(n3244)
         );
  OR2_X1 U4125 ( .A1(n3245), .A2(n3244), .ZN(U3245) );
  NAND2_X1 U4126 ( .A1(n3578), .A2(U4043), .ZN(n3246) );
  OAI21_X1 U4127 ( .B1(U4043), .B2(n3247), .A(n3246), .ZN(U3554) );
  NAND2_X1 U4128 ( .A1(n4632), .A2(U4043), .ZN(n3248) );
  OAI21_X1 U4129 ( .B1(U4043), .B2(n3249), .A(n3248), .ZN(U3562) );
  NAND2_X1 U4130 ( .A1(n4078), .A2(U4043), .ZN(n3250) );
  OAI21_X1 U4131 ( .B1(U4043), .B2(n3251), .A(n3250), .ZN(U3560) );
  NAND2_X1 U4132 ( .A1(n4091), .A2(U4043), .ZN(n3252) );
  OAI21_X1 U4133 ( .B1(U4043), .B2(n3253), .A(n3252), .ZN(U3567) );
  INV_X1 U4134 ( .A(REG1_REG_31__SCAN_IN), .ZN(n4698) );
  NAND2_X1 U4135 ( .A1(n2572), .A2(REG2_REG_31__SCAN_IN), .ZN(n3256) );
  OR2_X1 U4136 ( .A1(n3259), .A2(n3254), .ZN(n3255) );
  OAI211_X1 U4137 ( .C1(n3262), .C2(n4698), .A(n3256), .B(n3255), .ZN(n4345)
         );
  NAND2_X1 U4138 ( .A1(n4345), .A2(U4043), .ZN(n3257) );
  OAI21_X1 U4139 ( .B1(U4043), .B2(n3258), .A(n3257), .ZN(U3581) );
  INV_X1 U4140 ( .A(REG1_REG_30__SCAN_IN), .ZN(n4703) );
  NAND2_X1 U4141 ( .A1(n2572), .A2(REG2_REG_30__SCAN_IN), .ZN(n3261) );
  INV_X1 U4142 ( .A(REG0_REG_30__SCAN_IN), .ZN(n4814) );
  OR2_X1 U4143 ( .A1(n3259), .A2(n4814), .ZN(n3260) );
  OAI211_X1 U4144 ( .C1(n3262), .C2(n4703), .A(n3261), .B(n3260), .ZN(n4360)
         );
  NAND2_X1 U4145 ( .A1(n4360), .A2(U4043), .ZN(n3263) );
  OAI21_X1 U4146 ( .B1(U4043), .B2(n3264), .A(n3263), .ZN(U3580) );
  NAND2_X1 U4147 ( .A1(n3990), .A2(U4043), .ZN(n3265) );
  OAI21_X1 U4148 ( .B1(U4043), .B2(n3266), .A(n3265), .ZN(U3565) );
  XOR2_X1 U4149 ( .A(n3267), .B(n3268), .Z(n3273) );
  INV_X1 U4150 ( .A(n3269), .ZN(n4290) );
  MUX2_X1 U4151 ( .A(REG2_REG_1__SCAN_IN), .B(n3270), .S(n3276), .Z(n3271) );
  AOI211_X1 U4152 ( .C1(n3269), .C2(n3271), .A(n2197), .B(n3705), .ZN(n3272)
         );
  AOI21_X1 U4153 ( .B1(n4935), .B2(n3273), .A(n3272), .ZN(n3275) );
  AOI22_X1 U4154 ( .A1(n4942), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3274) );
  OAI211_X1 U4155 ( .C1(n3276), .C2(n4949), .A(n3275), .B(n3274), .ZN(U3241)
         );
  NAND2_X1 U4156 ( .A1(n4545), .A2(U4043), .ZN(n3277) );
  OAI21_X1 U4157 ( .B1(U4043), .B2(n3278), .A(n3277), .ZN(U3569) );
  NAND2_X1 U4158 ( .A1(n4484), .A2(U4043), .ZN(n3279) );
  OAI21_X1 U4159 ( .B1(U4043), .B2(n3280), .A(n3279), .ZN(U3570) );
  INV_X1 U4160 ( .A(n4989), .ZN(n4998) );
  NAND2_X1 U4161 ( .A1(n3313), .A2(n3855), .ZN(n4127) );
  NAND2_X1 U4162 ( .A1(n4126), .A2(n4127), .ZN(n4954) );
  NOR2_X1 U4163 ( .A1(n3855), .A2(n3329), .ZN(n4952) );
  INV_X1 U4164 ( .A(n3322), .ZN(n3384) );
  INV_X1 U4165 ( .A(n3574), .ZN(n4636) );
  OAI21_X1 U4166 ( .B1(n4636), .B2(n4525), .A(n4954), .ZN(n3281) );
  OAI21_X1 U4167 ( .B1(n3384), .B2(n4678), .A(n3281), .ZN(n4950) );
  AOI211_X1 U4168 ( .C1(n4998), .C2(n4954), .A(n4952), .B(n4950), .ZN(n4987)
         );
  NAND2_X1 U4169 ( .A1(n5017), .A2(REG1_REG_0__SCAN_IN), .ZN(n3282) );
  OAI21_X1 U4170 ( .B1(n4987), .B2(n5017), .A(n3282), .ZN(U3518) );
  NAND2_X1 U4171 ( .A1(n4220), .A2(n3283), .ZN(n3381) );
  OAI21_X1 U4172 ( .B1(n4220), .B2(n3283), .A(n3381), .ZN(n3410) );
  OAI21_X1 U4173 ( .B1(n3284), .B2(n3285), .A(n3386), .ZN(n3289) );
  NAND2_X1 U4174 ( .A1(n3313), .A2(n4682), .ZN(n3287) );
  NAND2_X1 U4175 ( .A1(n3712), .A2(n4563), .ZN(n3286) );
  OAI211_X1 U4176 ( .C1(n4795), .C2(n3348), .A(n3287), .B(n3286), .ZN(n3288)
         );
  AOI21_X1 U4177 ( .B1(n3289), .B2(n4525), .A(n3288), .ZN(n3290) );
  OAI21_X1 U4178 ( .B1(n3574), .B2(n3410), .A(n3290), .ZN(n3411) );
  INV_X1 U4179 ( .A(n3393), .ZN(n3292) );
  NAND2_X1 U4180 ( .A1(n3321), .A2(n3315), .ZN(n3291) );
  NAND2_X1 U4181 ( .A1(n3292), .A2(n3291), .ZN(n3416) );
  OAI22_X1 U4182 ( .A1(n3410), .A2(n4989), .B1(n5000), .B2(n3416), .ZN(n3293)
         );
  NOR2_X1 U4183 ( .A1(n3411), .A2(n3293), .ZN(n4988) );
  NAND2_X1 U4184 ( .A1(n5017), .A2(REG1_REG_1__SCAN_IN), .ZN(n3294) );
  OAI21_X1 U4185 ( .B1(n4988), .B2(n5017), .A(n3294), .ZN(U3519) );
  OR2_X1 U4186 ( .A1(n3299), .A2(n3601), .ZN(n3295) );
  XOR2_X1 U4187 ( .A(n3435), .B(REG2_REG_8__SCAN_IN), .Z(n3306) );
  INV_X1 U4188 ( .A(n3299), .ZN(n3300) );
  OAI211_X1 U4189 ( .C1(n3301), .C2(REG1_REG_8__SCAN_IN), .A(n3443), .B(n4935), 
        .ZN(n3304) );
  NAND2_X1 U4190 ( .A1(REG3_REG_8__SCAN_IN), .A2(U3149), .ZN(n3568) );
  INV_X1 U4191 ( .A(n3568), .ZN(n3302) );
  AOI21_X1 U4192 ( .B1(n4942), .B2(ADDR_REG_8__SCAN_IN), .A(n3302), .ZN(n3303)
         );
  OAI211_X1 U4193 ( .C1(n4949), .C2(n3444), .A(n3304), .B(n3303), .ZN(n3305)
         );
  AOI21_X1 U4194 ( .B1(n4948), .B2(n3306), .A(n3305), .ZN(n3307) );
  INV_X1 U4195 ( .A(n3307), .ZN(U3248) );
  INV_X1 U4196 ( .A(n3408), .ZN(n3308) );
  NAND2_X1 U4197 ( .A1(n3313), .A2(n3760), .ZN(n3310) );
  AND2_X4 U4198 ( .A1(n3408), .A2(n3369), .ZN(n3826) );
  NAND2_X1 U4199 ( .A1(n3826), .A2(n3315), .ZN(n3309) );
  NAND2_X1 U4200 ( .A1(n3310), .A2(n3309), .ZN(n3318) );
  INV_X1 U4201 ( .A(REG1_REG_0__SCAN_IN), .ZN(n3311) );
  NOR2_X1 U4202 ( .A1(n3369), .A2(n3311), .ZN(n3312) );
  OR2_X1 U4203 ( .A1(n3318), .A2(n3312), .ZN(n3851) );
  NAND2_X1 U4204 ( .A1(n3420), .A2(n3313), .ZN(n3317) );
  INV_X1 U4205 ( .A(n3369), .ZN(n3314) );
  AOI22_X1 U4206 ( .A1(n3760), .A2(n3315), .B1(n3314), .B2(n2222), .ZN(n3316)
         );
  NAND2_X1 U4207 ( .A1(n3317), .A2(n3316), .ZN(n3849) );
  INV_X1 U4208 ( .A(n3318), .ZN(n3319) );
  NAND2_X4 U4209 ( .A1(n3408), .A2(n3334), .ZN(n3841) );
  AOI22_X1 U4210 ( .A1(n3420), .A2(n3322), .B1(n3321), .B2(n3760), .ZN(n3355)
         );
  XNOR2_X1 U4211 ( .A(n3356), .B(n3357), .ZN(n3351) );
  NOR2_X1 U4212 ( .A1(n3323), .A2(n3165), .ZN(n3325) );
  OAI21_X1 U4213 ( .B1(n3326), .B2(n3325), .A(n3324), .ZN(n3405) );
  INV_X1 U4214 ( .A(n3405), .ZN(n3327) );
  OAI211_X1 U4215 ( .C1(n3329), .C2(n4339), .A(n3328), .B(n4795), .ZN(n3331)
         );
  NOR2_X1 U4216 ( .A1(n3403), .A2(n3331), .ZN(n3330) );
  INV_X1 U4217 ( .A(n3346), .ZN(n3337) );
  NAND2_X1 U4218 ( .A1(n3331), .A2(n4795), .ZN(n3332) );
  NAND2_X1 U4219 ( .A1(n3337), .A2(n3332), .ZN(n3333) );
  NAND2_X1 U4220 ( .A1(n3333), .A2(n3401), .ZN(n3371) );
  INV_X1 U4221 ( .A(n3371), .ZN(n3339) );
  INV_X1 U4222 ( .A(n3334), .ZN(n3335) );
  NAND2_X1 U4223 ( .A1(n4978), .A2(n3335), .ZN(n3336) );
  INV_X1 U4224 ( .A(n3344), .ZN(n4271) );
  NAND2_X1 U4225 ( .A1(n3337), .A2(n4271), .ZN(n3372) );
  NAND3_X1 U4226 ( .A1(n3339), .A2(n3338), .A3(n3372), .ZN(n3852) );
  NOR2_X1 U4227 ( .A1(n3403), .A2(n4795), .ZN(n3340) );
  NAND2_X1 U4228 ( .A1(n3346), .A2(n3340), .ZN(n3342) );
  NOR2_X1 U4229 ( .A1(n3344), .A2(n4287), .ZN(n3343) );
  NAND2_X1 U4230 ( .A1(n3346), .A2(n3343), .ZN(n4067) );
  NOR2_X1 U4231 ( .A1(n3344), .A2(n4888), .ZN(n3345) );
  AOI22_X1 U4232 ( .A1(n4115), .A2(n3712), .B1(n4116), .B2(n3313), .ZN(n3347)
         );
  OAI21_X1 U4233 ( .B1(n4064), .B2(n3348), .A(n3347), .ZN(n3349) );
  AOI21_X1 U4234 ( .B1(REG3_REG_1__SCAN_IN), .B2(n3852), .A(n3349), .ZN(n3350)
         );
  OAI21_X1 U4235 ( .B1(n3351), .B2(n4108), .A(n3350), .ZN(U3219) );
  NAND2_X1 U4236 ( .A1(n4284), .A2(n3760), .ZN(n3353) );
  NAND2_X1 U4237 ( .A1(n3826), .A2(n3553), .ZN(n3352) );
  NAND2_X1 U4238 ( .A1(n3353), .A2(n3352), .ZN(n3354) );
  AOI22_X1 U4239 ( .A1(n3420), .A2(n4284), .B1(n3760), .B2(n3553), .ZN(n3424)
         );
  XNOR2_X1 U4240 ( .A(n3423), .B(n3424), .ZN(n3367) );
  INV_X1 U4241 ( .A(n3718), .ZN(n3364) );
  NAND2_X1 U4242 ( .A1(n3712), .A2(n3760), .ZN(n3359) );
  NAND2_X1 U4243 ( .A1(n3391), .A2(n3826), .ZN(n3358) );
  NAND2_X1 U4244 ( .A1(n3359), .A2(n3358), .ZN(n3360) );
  XNOR2_X1 U4245 ( .A(n3360), .B(n3871), .ZN(n3362) );
  AOI22_X1 U4246 ( .A1(n3420), .A2(n3712), .B1(n3391), .B2(n3760), .ZN(n3361)
         );
  NAND2_X1 U4247 ( .A1(n3362), .A2(n3361), .ZN(n3365) );
  INV_X1 U4248 ( .A(n3717), .ZN(n3363) );
  NAND2_X1 U4249 ( .A1(n3364), .A2(n3363), .ZN(n3715) );
  NAND2_X1 U4250 ( .A1(n3715), .A2(n3365), .ZN(n3366) );
  OAI21_X1 U4251 ( .B1(n3367), .B2(n3366), .A(n4019), .ZN(n3378) );
  NAND2_X1 U4252 ( .A1(n3369), .A2(n3368), .ZN(n3370) );
  OAI21_X1 U4253 ( .B1(n3371), .B2(n3370), .A(STATE_REG_SCAN_IN), .ZN(n3373)
         );
  AOI21_X1 U4254 ( .B1(n4115), .B2(n3578), .A(n3374), .ZN(n3376) );
  AOI22_X1 U4255 ( .A1(n3553), .A2(n4117), .B1(n4116), .B2(n3712), .ZN(n3375)
         );
  OAI211_X1 U4256 ( .C1(n4120), .C2(REG3_REG_3__SCAN_IN), .A(n3376), .B(n3375), 
        .ZN(n3377) );
  AOI21_X1 U4257 ( .B1(n3378), .B2(n4122), .A(n3377), .ZN(n3379) );
  INV_X1 U4258 ( .A(n3379), .ZN(U3215) );
  NAND2_X1 U4259 ( .A1(n3381), .A2(n3380), .ZN(n3382) );
  XNOR2_X1 U4260 ( .A(n3382), .B(n4223), .ZN(n3540) );
  INV_X1 U4261 ( .A(n4284), .ZN(n3383) );
  OAI22_X1 U4262 ( .A1(n3384), .A2(n4659), .B1(n3383), .B2(n4678), .ZN(n3390)
         );
  INV_X1 U4263 ( .A(n4223), .ZN(n3385) );
  NAND3_X1 U4264 ( .A1(n3386), .A2(n3385), .A3(n4131), .ZN(n3387) );
  AOI21_X1 U4265 ( .B1(n3388), .B2(n3387), .A(n4684), .ZN(n3389) );
  AOI211_X1 U4266 ( .C1(n3540), .C2(n4636), .A(n3390), .B(n3389), .ZN(n3542)
         );
  AOI22_X1 U4267 ( .A1(n3540), .A2(n4998), .B1(n3391), .B2(n4768), .ZN(n3392)
         );
  NAND2_X1 U4268 ( .A1(n3542), .A2(n3392), .ZN(n3397) );
  OAI21_X1 U4269 ( .B1(n3393), .B2(n3720), .A(n3552), .ZN(n3536) );
  OAI22_X1 U4270 ( .A1(n4872), .A2(n3536), .B1(n5013), .B2(n2510), .ZN(n3394)
         );
  AOI21_X1 U4271 ( .B1(n3397), .B2(n5013), .A(n3394), .ZN(n3395) );
  INV_X1 U4272 ( .A(n3395), .ZN(U3471) );
  OAI22_X1 U4273 ( .A1(n4801), .A2(n3536), .B1(n5019), .B2(n3169), .ZN(n3396)
         );
  AOI21_X1 U4274 ( .B1(n3397), .B2(n5019), .A(n3396), .ZN(n3398) );
  INV_X1 U4275 ( .A(n3398), .ZN(U3520) );
  NAND2_X1 U4276 ( .A1(n4473), .A2(U4043), .ZN(n3399) );
  OAI21_X1 U4277 ( .B1(U4043), .B2(n3400), .A(n3399), .ZN(U3573) );
  INV_X1 U4278 ( .A(n3401), .ZN(n3402) );
  OR2_X1 U4279 ( .A1(n3403), .A2(n3402), .ZN(n3404) );
  OAI21_X4 U4280 ( .B1(n3407), .B2(n3406), .A(n4643), .ZN(n4957) );
  NAND2_X1 U4281 ( .A1(n4957), .A2(n4339), .ZN(n4554) );
  OR2_X1 U4282 ( .A1(n3408), .A2(n4339), .ZN(n3573) );
  INV_X1 U4283 ( .A(n3573), .ZN(n3409) );
  NAND2_X1 U4284 ( .A1(n4957), .A2(n3409), .ZN(n4649) );
  INV_X1 U4285 ( .A(n4649), .ZN(n4955) );
  INV_X1 U4286 ( .A(n3410), .ZN(n3414) );
  AOI22_X1 U4287 ( .A1(n3411), .A2(n4957), .B1(REG3_REG_1__SCAN_IN), .B2(n4953), .ZN(n3412) );
  OAI21_X1 U4288 ( .B1(n3270), .B2(n4957), .A(n3412), .ZN(n3413) );
  AOI21_X1 U4289 ( .B1(n4955), .B2(n3414), .A(n3413), .ZN(n3415) );
  OAI21_X1 U4290 ( .B1(n4572), .B2(n3416), .A(n3415), .ZN(U3289) );
  NAND2_X1 U4291 ( .A1(n4283), .A2(n3760), .ZN(n3418) );
  NAND2_X1 U4292 ( .A1(n3826), .A2(n3582), .ZN(n3417) );
  NAND2_X1 U4293 ( .A1(n3418), .A2(n3417), .ZN(n3419) );
  AOI22_X1 U4294 ( .A1(n3831), .A2(n4283), .B1(n3582), .B2(n3760), .ZN(n3465)
         );
  AOI22_X1 U4295 ( .A1(n3420), .A2(n3578), .B1(n4023), .B2(n3760), .ZN(n3427)
         );
  AOI22_X1 U4296 ( .A1(n3578), .A2(n3760), .B1(n4023), .B2(n3826), .ZN(n3421)
         );
  XNOR2_X1 U4297 ( .A(n3421), .B(n3841), .ZN(n3426) );
  XNOR2_X1 U4298 ( .A(n3426), .B(n3422), .ZN(n4021) );
  INV_X1 U4299 ( .A(n3423), .ZN(n3425) );
  NAND2_X1 U4300 ( .A1(n3425), .A2(n3424), .ZN(n4018) );
  INV_X1 U4301 ( .A(n3428), .ZN(n3585) );
  AOI21_X1 U4302 ( .B1(n4115), .B2(n4282), .A(n3429), .ZN(n3431) );
  AOI22_X1 U4303 ( .A1(n3582), .A2(n4117), .B1(n4116), .B2(n3578), .ZN(n3430)
         );
  OAI211_X1 U4304 ( .C1(n4120), .C2(n3585), .A(n3431), .B(n3430), .ZN(n3432)
         );
  AOI21_X1 U4305 ( .B1(n3433), .B2(n4122), .A(n3432), .ZN(n3434) );
  INV_X1 U4306 ( .A(n3434), .ZN(U3224) );
  NAND2_X1 U4307 ( .A1(n3435), .A2(REG2_REG_8__SCAN_IN), .ZN(n3439) );
  NAND2_X1 U4308 ( .A1(n3437), .A2(n3436), .ZN(n3438) );
  NAND2_X1 U4309 ( .A1(n3439), .A2(n3438), .ZN(n4311) );
  INV_X1 U4310 ( .A(REG2_REG_9__SCAN_IN), .ZN(n4687) );
  MUX2_X1 U4311 ( .A(REG2_REG_9__SCAN_IN), .B(n4687), .S(n4884), .Z(n4310) );
  NAND2_X1 U4312 ( .A1(n4311), .A2(n4310), .ZN(n4309) );
  NAND2_X1 U4313 ( .A1(n4884), .A2(REG2_REG_9__SCAN_IN), .ZN(n3440) );
  XOR2_X1 U4314 ( .A(n3525), .B(REG2_REG_10__SCAN_IN), .Z(n3450) );
  AND2_X1 U4315 ( .A1(U3149), .A2(REG3_REG_10__SCAN_IN), .ZN(n3938) );
  AOI21_X1 U4316 ( .B1(n4942), .B2(ADDR_REG_10__SCAN_IN), .A(n3938), .ZN(n3441) );
  OAI21_X1 U4317 ( .B1(n4949), .B2(n3442), .A(n3441), .ZN(n3449) );
  INV_X1 U4318 ( .A(n4884), .ZN(n4306) );
  XOR2_X1 U4319 ( .A(REG1_REG_9__SCAN_IN), .B(n4884), .Z(n4304) );
  AOI211_X1 U4320 ( .C1(n3447), .C2(n4799), .A(n4938), .B(n3523), .ZN(n3448)
         );
  AOI211_X1 U4321 ( .C1(n4948), .C2(n3450), .A(n3449), .B(n3448), .ZN(n3451)
         );
  INV_X1 U4322 ( .A(n3451), .ZN(U3250) );
  XOR2_X1 U4323 ( .A(n4199), .B(n3452), .Z(n3459) );
  INV_X1 U4324 ( .A(n3498), .ZN(n3453) );
  AOI21_X1 U4325 ( .B1(n4199), .B2(n3454), .A(n3453), .ZN(n4999) );
  INV_X1 U4326 ( .A(n4283), .ZN(n3456) );
  AOI22_X1 U4327 ( .A1(n4284), .A2(n4682), .B1(n4023), .B2(n4768), .ZN(n3455)
         );
  OAI21_X1 U4328 ( .B1(n3456), .B2(n4678), .A(n3455), .ZN(n3457) );
  AOI21_X1 U4329 ( .B1(n4999), .B2(n4636), .A(n3457), .ZN(n3458) );
  OAI21_X1 U4330 ( .B1(n4684), .B2(n3459), .A(n3458), .ZN(n4996) );
  OAI211_X1 U4331 ( .C1(n3551), .C2(n3460), .A(n3583), .B(n4994), .ZN(n4995)
         );
  INV_X1 U4332 ( .A(n3461), .ZN(n4024) );
  OAI22_X1 U4333 ( .A1(n4995), .A2(n4881), .B1(n4643), .B2(n4024), .ZN(n3462)
         );
  OAI21_X1 U4334 ( .B1(n4996), .B2(n3462), .A(n4957), .ZN(n3464) );
  AOI22_X1 U4335 ( .A1(n4999), .A2(n4955), .B1(REG2_REG_4__SCAN_IN), .B2(n2142), .ZN(n3463) );
  NAND2_X1 U4336 ( .A1(n3464), .A2(n3463), .ZN(U3286) );
  INV_X1 U4337 ( .A(n3465), .ZN(n3467) );
  NAND2_X1 U4338 ( .A1(n4282), .A2(n3760), .ZN(n3470) );
  NAND2_X1 U4339 ( .A1(n3826), .A2(n3605), .ZN(n3469) );
  NAND2_X1 U4340 ( .A1(n3470), .A2(n3469), .ZN(n3471) );
  XNOR2_X1 U4341 ( .A(n3471), .B(n3871), .ZN(n3473) );
  AOI22_X1 U4342 ( .A1(n3831), .A2(n4282), .B1(n3605), .B2(n3796), .ZN(n3472)
         );
  AND2_X1 U4343 ( .A1(n3473), .A2(n3472), .ZN(n3483) );
  NOR2_X1 U4344 ( .A1(n2189), .A2(n3483), .ZN(n3474) );
  XNOR2_X1 U4345 ( .A(n3484), .B(n3474), .ZN(n3480) );
  AOI21_X1 U4346 ( .B1(n4115), .B2(n4281), .A(n3475), .ZN(n3477) );
  AOI22_X1 U4347 ( .A1(n3605), .A2(n4117), .B1(n4116), .B2(n4283), .ZN(n3476)
         );
  OAI211_X1 U4348 ( .C1(n4120), .C2(n3478), .A(n3477), .B(n3476), .ZN(n3479)
         );
  AOI21_X1 U4349 ( .B1(n3480), .B2(n4122), .A(n3479), .ZN(n3481) );
  INV_X1 U4350 ( .A(n3481), .ZN(U3236) );
  INV_X1 U4351 ( .A(n3482), .ZN(n3600) );
  NAND2_X1 U4352 ( .A1(n4281), .A2(n3760), .ZN(n3486) );
  NAND2_X1 U4353 ( .A1(n3826), .A2(n3597), .ZN(n3485) );
  NAND2_X1 U4354 ( .A1(n3486), .A2(n3485), .ZN(n3487) );
  XNOR2_X1 U4355 ( .A(n3487), .B(n3841), .ZN(n3558) );
  AOI22_X1 U4356 ( .A1(n3420), .A2(n4281), .B1(n3597), .B2(n3796), .ZN(n3561)
         );
  XNOR2_X1 U4357 ( .A(n3558), .B(n3561), .ZN(n3488) );
  OAI211_X1 U4358 ( .C1(n3489), .C2(n3488), .A(n3559), .B(n4122), .ZN(n3493)
         );
  INV_X1 U4359 ( .A(n4282), .ZN(n3608) );
  OAI22_X1 U4360 ( .A1(n4064), .A2(n3593), .B1(n4065), .B2(n3608), .ZN(n3490)
         );
  AOI211_X1 U4361 ( .C1(n4115), .C2(n4681), .A(n3491), .B(n3490), .ZN(n3492)
         );
  OAI211_X1 U4362 ( .C1(n4120), .C2(n3600), .A(n3493), .B(n3492), .ZN(U3210)
         );
  NAND2_X1 U4363 ( .A1(n4400), .A2(U4043), .ZN(n3494) );
  OAI21_X1 U4364 ( .B1(U4043), .B2(n3495), .A(n3494), .ZN(U3577) );
  NAND2_X1 U4365 ( .A1(n4142), .A2(n4152), .ZN(n4219) );
  XOR2_X1 U4366 ( .A(n4219), .B(n3496), .Z(n3506) );
  NAND2_X1 U4367 ( .A1(n3498), .A2(n3497), .ZN(n3616) );
  INV_X1 U4368 ( .A(n3499), .ZN(n3500) );
  NAND2_X1 U4369 ( .A1(n3616), .A2(n3500), .ZN(n3502) );
  NAND2_X1 U4370 ( .A1(n3502), .A2(n3501), .ZN(n3606) );
  XNOR2_X1 U4371 ( .A(n3606), .B(n4219), .ZN(n3514) );
  AOI22_X1 U4372 ( .A1(n4283), .A2(n4682), .B1(n4768), .B2(n3605), .ZN(n3504)
         );
  NAND2_X1 U4373 ( .A1(n4281), .A2(n4563), .ZN(n3503) );
  OAI211_X1 U4374 ( .C1(n3514), .C2(n3574), .A(n3504), .B(n3503), .ZN(n3505)
         );
  AOI21_X1 U4375 ( .B1(n4525), .B2(n3506), .A(n3505), .ZN(n3513) );
  INV_X1 U4376 ( .A(n3514), .ZN(n3511) );
  NAND2_X1 U4377 ( .A1(n2151), .A2(n3605), .ZN(n3507) );
  NAND2_X1 U4378 ( .A1(n3598), .A2(n3507), .ZN(n3517) );
  AOI22_X1 U4379 ( .A1(n2142), .A2(REG2_REG_6__SCAN_IN), .B1(n3508), .B2(n4953), .ZN(n3509) );
  OAI21_X1 U4380 ( .B1(n4572), .B2(n3517), .A(n3509), .ZN(n3510) );
  AOI21_X1 U4381 ( .B1(n3511), .B2(n4955), .A(n3510), .ZN(n3512) );
  OAI21_X1 U4382 ( .B1(n3513), .B2(n2142), .A(n3512), .ZN(U3284) );
  OAI21_X1 U4383 ( .B1(n4989), .B2(n3514), .A(n3513), .ZN(n3519) );
  OAI22_X1 U4384 ( .A1(n3517), .A2(n4801), .B1(n5019), .B2(n2573), .ZN(n3515)
         );
  AOI21_X1 U4385 ( .B1(n3519), .B2(n5019), .A(n3515), .ZN(n3516) );
  INV_X1 U4386 ( .A(n3516), .ZN(U3524) );
  OAI22_X1 U4387 ( .A1(n3517), .A2(n4872), .B1(n5013), .B2(n2574), .ZN(n3518)
         );
  AOI21_X1 U4388 ( .B1(n3519), .B2(n5013), .A(n3518), .ZN(n3520) );
  INV_X1 U4389 ( .A(n3520), .ZN(U3479) );
  XOR2_X1 U4390 ( .A(REG1_REG_11__SCAN_IN), .B(n3671), .Z(n3524) );
  AOI211_X1 U4391 ( .C1(n2186), .C2(n3524), .A(n4938), .B(n3672), .ZN(n3535)
         );
  NAND2_X1 U4392 ( .A1(n3525), .A2(REG2_REG_10__SCAN_IN), .ZN(n3529) );
  NAND2_X1 U4393 ( .A1(n3527), .A2(n3526), .ZN(n3528) );
  MUX2_X1 U4394 ( .A(n3109), .B(REG2_REG_11__SCAN_IN), .S(n3671), .Z(n3530) );
  NAND2_X1 U4395 ( .A1(n3531), .A2(n3530), .ZN(n3670) );
  OAI211_X1 U4396 ( .C1(n3531), .C2(n3530), .A(n3670), .B(n4948), .ZN(n3533)
         );
  AND2_X1 U4397 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n4077) );
  AOI21_X1 U4398 ( .B1(n4942), .B2(ADDR_REG_11__SCAN_IN), .A(n4077), .ZN(n3532) );
  OAI211_X1 U4399 ( .C1(n4949), .C2(n3671), .A(n3533), .B(n3532), .ZN(n3534)
         );
  OR2_X1 U4400 ( .A1(n3535), .A2(n3534), .ZN(U3251) );
  NOR2_X1 U4401 ( .A1(n4572), .A2(n3536), .ZN(n3539) );
  AND2_X1 U4402 ( .A1(n4957), .A2(n4768), .ZN(n4619) );
  AOI22_X1 U4403 ( .A1(n2142), .A2(REG2_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(n4953), .ZN(n3537) );
  OAI21_X1 U4404 ( .B1(n4666), .B2(n3720), .A(n3537), .ZN(n3538) );
  AOI211_X1 U4405 ( .C1(n3540), .C2(n4955), .A(n3539), .B(n3538), .ZN(n3541)
         );
  OAI21_X1 U4406 ( .B1(n2142), .B2(n3542), .A(n3541), .ZN(U3288) );
  XOR2_X1 U4407 ( .A(n4221), .B(n3543), .Z(n4990) );
  OAI21_X1 U4408 ( .B1(n4221), .B2(n3545), .A(n3544), .ZN(n3549) );
  INV_X1 U4409 ( .A(n3578), .ZN(n3547) );
  AOI22_X1 U4410 ( .A1(n3712), .A2(n4682), .B1(n3553), .B2(n4768), .ZN(n3546)
         );
  OAI21_X1 U4411 ( .B1(n3547), .B2(n4678), .A(n3546), .ZN(n3548) );
  AOI21_X1 U4412 ( .B1(n3549), .B2(n4525), .A(n3548), .ZN(n3550) );
  OAI21_X1 U4413 ( .B1(n4990), .B2(n3574), .A(n3550), .ZN(n4991) );
  INV_X1 U4414 ( .A(n4991), .ZN(n3557) );
  AOI21_X1 U4415 ( .B1(n3553), .B2(n3552), .A(n3551), .ZN(n4993) );
  AOI22_X1 U4416 ( .A1(n2142), .A2(REG2_REG_3__SCAN_IN), .B1(n4953), .B2(n2543), .ZN(n3554) );
  OAI21_X1 U4417 ( .B1(n4990), .B2(n4649), .A(n3554), .ZN(n3555) );
  AOI21_X1 U4418 ( .B1(n4693), .B2(n4993), .A(n3555), .ZN(n3556) );
  OAI21_X1 U4419 ( .B1(n3557), .B2(n2142), .A(n3556), .ZN(U3287) );
  INV_X1 U4420 ( .A(n3558), .ZN(n3560) );
  NAND2_X1 U4421 ( .A1(n4681), .A2(n3755), .ZN(n3563) );
  NAND2_X1 U4422 ( .A1(n3826), .A2(n3628), .ZN(n3562) );
  NAND2_X1 U4423 ( .A1(n3563), .A2(n3562), .ZN(n3564) );
  NAND2_X1 U4424 ( .A1(n3420), .A2(n4681), .ZN(n3566) );
  NAND2_X1 U4425 ( .A1(n3760), .A2(n3628), .ZN(n3565) );
  NAND2_X1 U4426 ( .A1(n3566), .A2(n3565), .ZN(n3927) );
  INV_X1 U4427 ( .A(n3927), .ZN(n3930) );
  XNOR2_X1 U4428 ( .A(n3926), .B(n3930), .ZN(n3567) );
  XNOR2_X1 U4429 ( .A(n3928), .B(n3567), .ZN(n3572) );
  INV_X1 U4430 ( .A(n4280), .ZN(n4658) );
  AOI22_X1 U4431 ( .A1(n3628), .A2(n4117), .B1(n4116), .B2(n4281), .ZN(n3569)
         );
  OAI211_X1 U4432 ( .C1(n4658), .C2(n4067), .A(n3569), .B(n3568), .ZN(n3570)
         );
  AOI21_X1 U4433 ( .B1(n3629), .B2(n4102), .A(n3570), .ZN(n3571) );
  OAI21_X1 U4434 ( .B1(n3572), .B2(n4108), .A(n3571), .ZN(U3218) );
  NAND2_X1 U4435 ( .A1(n3574), .A2(n3573), .ZN(n3575) );
  INV_X1 U4436 ( .A(n3576), .ZN(n4139) );
  XOR2_X1 U4437 ( .A(n4212), .B(n3616), .Z(n5003) );
  XNOR2_X1 U4438 ( .A(n3577), .B(n4212), .ZN(n3581) );
  AOI22_X1 U4439 ( .A1(n3578), .A2(n4682), .B1(n4768), .B2(n3582), .ZN(n3580)
         );
  NAND2_X1 U4440 ( .A1(n4282), .A2(n4563), .ZN(n3579) );
  OAI211_X1 U4441 ( .C1(n3581), .C2(n4684), .A(n3580), .B(n3579), .ZN(n5004)
         );
  NAND2_X1 U4442 ( .A1(n5004), .A2(n4957), .ZN(n3590) );
  NAND2_X1 U4443 ( .A1(n3583), .A2(n3582), .ZN(n3584) );
  NAND2_X1 U4444 ( .A1(n2151), .A2(n3584), .ZN(n5001) );
  INV_X1 U4445 ( .A(n5001), .ZN(n3588) );
  OAI22_X1 U4446 ( .A1(n4957), .A2(n3586), .B1(n3585), .B2(n4643), .ZN(n3587)
         );
  AOI21_X1 U4447 ( .B1(n4693), .B2(n3588), .A(n3587), .ZN(n3589) );
  OAI211_X1 U4448 ( .C1(n4697), .C2(n5003), .A(n3590), .B(n3589), .ZN(U3285)
         );
  INV_X1 U4449 ( .A(n3610), .ZN(n4222) );
  XNOR2_X1 U4450 ( .A(n3622), .B(n4222), .ZN(n3595) );
  NAND2_X1 U4451 ( .A1(n4681), .A2(n4563), .ZN(n3592) );
  NAND2_X1 U4452 ( .A1(n4282), .A2(n4682), .ZN(n3591) );
  OAI211_X1 U4453 ( .C1(n4795), .C2(n3593), .A(n3592), .B(n3591), .ZN(n3594)
         );
  AOI21_X1 U4454 ( .B1(n3595), .B2(n4525), .A(n3594), .ZN(n5011) );
  INV_X1 U4455 ( .A(n3596), .ZN(n3627) );
  AOI21_X1 U4456 ( .B1(n3598), .B2(n3597), .A(n5000), .ZN(n3599) );
  NAND2_X1 U4457 ( .A1(n3627), .A2(n3599), .ZN(n5010) );
  INV_X1 U4458 ( .A(n5010), .ZN(n3604) );
  INV_X1 U4459 ( .A(n4554), .ZN(n3603) );
  OAI22_X1 U4460 ( .A1(n4957), .A2(n3601), .B1(n3600), .B2(n4643), .ZN(n3602)
         );
  AOI21_X1 U4461 ( .B1(n3604), .B2(n3603), .A(n3602), .ZN(n3614) );
  INV_X1 U4462 ( .A(n3606), .ZN(n3609) );
  AOI21_X1 U4463 ( .B1(n3606), .B2(n4282), .A(n3605), .ZN(n3607) );
  AOI21_X1 U4464 ( .B1(n3609), .B2(n3608), .A(n3607), .ZN(n3611) );
  NAND2_X1 U4465 ( .A1(n3611), .A2(n3610), .ZN(n5008) );
  INV_X1 U4466 ( .A(n3611), .ZN(n3612) );
  NAND2_X1 U4467 ( .A1(n3612), .A2(n4222), .ZN(n5006) );
  NAND3_X1 U4468 ( .A1(n5008), .A2(n4577), .A3(n5006), .ZN(n3613) );
  OAI211_X1 U4469 ( .C1(n5011), .C2(n2142), .A(n3614), .B(n3613), .ZN(U3283)
         );
  NAND2_X1 U4470 ( .A1(n3616), .A2(n3615), .ZN(n3619) );
  INV_X1 U4471 ( .A(n3617), .ZN(n3618) );
  NAND2_X1 U4472 ( .A1(n3619), .A2(n3618), .ZN(n3620) );
  XOR2_X1 U4473 ( .A(n4210), .B(n3620), .Z(n3635) );
  INV_X1 U4474 ( .A(n4281), .ZN(n3625) );
  OR2_X1 U4475 ( .A1(n3622), .A2(n3621), .ZN(n3623) );
  NAND2_X1 U4476 ( .A1(n3623), .A2(n4144), .ZN(n4673) );
  XNOR2_X1 U4477 ( .A(n4673), .B(n4210), .ZN(n3624) );
  OAI222_X1 U4478 ( .A1(n4678), .A2(n4658), .B1(n4659), .B2(n3625), .C1(n4684), 
        .C2(n3624), .ZN(n3637) );
  NAND2_X1 U4479 ( .A1(n3637), .A2(n4957), .ZN(n3633) );
  INV_X1 U4480 ( .A(n4689), .ZN(n3626) );
  AOI21_X1 U4481 ( .B1(n3628), .B2(n3627), .A(n3626), .ZN(n3639) );
  AOI22_X1 U4482 ( .A1(n2142), .A2(REG2_REG_8__SCAN_IN), .B1(n3629), .B2(n4953), .ZN(n3630) );
  OAI21_X1 U4483 ( .B1(n4666), .B2(n3634), .A(n3630), .ZN(n3631) );
  AOI21_X1 U4484 ( .B1(n3639), .B2(n4693), .A(n3631), .ZN(n3632) );
  OAI211_X1 U4485 ( .C1(n4697), .C2(n3635), .A(n3633), .B(n3632), .ZN(U3282)
         );
  OAI22_X1 U4486 ( .A1(n3635), .A2(n5002), .B1(n4795), .B2(n3634), .ZN(n3636)
         );
  NOR2_X1 U4487 ( .A1(n3637), .A2(n3636), .ZN(n3641) );
  INV_X1 U4488 ( .A(n4801), .ZN(n4804) );
  AOI22_X1 U4489 ( .A1(n3639), .A2(n4804), .B1(REG1_REG_8__SCAN_IN), .B2(n5017), .ZN(n3638) );
  OAI21_X1 U4490 ( .B1(n3641), .B2(n5017), .A(n3638), .ZN(U3526) );
  INV_X1 U4491 ( .A(n4872), .ZN(n4874) );
  AOI22_X1 U4492 ( .A1(n3639), .A2(n4874), .B1(REG0_REG_8__SCAN_IN), .B2(n5012), .ZN(n3640) );
  OAI21_X1 U4493 ( .B1(n3641), .B2(n5012), .A(n3640), .ZN(U3483) );
  AND2_X1 U4494 ( .A1(n3643), .A2(n3642), .ZN(n3644) );
  INV_X1 U4495 ( .A(n3645), .ZN(n4201) );
  XNOR2_X1 U4496 ( .A(n3644), .B(n4201), .ZN(n3651) );
  INV_X1 U4497 ( .A(n3646), .ZN(n3647) );
  OR2_X1 U4498 ( .A1(n3646), .A2(n3645), .ZN(n3661) );
  OAI21_X1 U4499 ( .B1(n3647), .B2(n4201), .A(n3661), .ZN(n4791) );
  AOI22_X1 U4500 ( .A1(n4563), .A2(n4632), .B1(n4078), .B2(n4682), .ZN(n3648)
         );
  OAI21_X1 U4501 ( .B1(n3652), .B2(n4795), .A(n3648), .ZN(n3649) );
  AOI21_X1 U4502 ( .B1(n4791), .B2(n4636), .A(n3649), .ZN(n3650) );
  OAI21_X1 U4503 ( .B1(n3651), .B2(n4684), .A(n3650), .ZN(n4790) );
  INV_X1 U4504 ( .A(n4790), .ZN(n3657) );
  NOR2_X1 U4505 ( .A1(n4661), .A2(n3652), .ZN(n3653) );
  OR2_X1 U4506 ( .A1(n3663), .A2(n3653), .ZN(n4868) );
  AOI22_X1 U4507 ( .A1(n2142), .A2(REG2_REG_11__SCAN_IN), .B1(n4076), .B2(
        n4953), .ZN(n3654) );
  OAI21_X1 U4508 ( .B1(n4868), .B2(n4572), .A(n3654), .ZN(n3655) );
  AOI21_X1 U4509 ( .B1(n4791), .B2(n4955), .A(n3655), .ZN(n3656) );
  OAI21_X1 U4510 ( .B1(n3657), .B2(n2142), .A(n3656), .ZN(U3279) );
  INV_X1 U4511 ( .A(n4279), .ZN(n4660) );
  INV_X1 U4512 ( .A(n4627), .ZN(n3658) );
  OR2_X1 U4513 ( .A1(n4628), .A2(n3658), .ZN(n4225) );
  XNOR2_X1 U4514 ( .A(n4629), .B(n4225), .ZN(n3659) );
  OAI222_X1 U4515 ( .A1(n4678), .A2(n3858), .B1(n4659), .B2(n4660), .C1(n3659), 
        .C2(n4684), .ZN(n4785) );
  INV_X1 U4516 ( .A(n4785), .ZN(n3668) );
  NAND2_X1 U4517 ( .A1(n3661), .A2(n3660), .ZN(n3662) );
  XNOR2_X1 U4518 ( .A(n3662), .B(n4225), .ZN(n4787) );
  OAI21_X1 U4519 ( .B1(n3663), .B2(n4784), .A(n4640), .ZN(n4864) );
  AOI22_X1 U4520 ( .A1(n2142), .A2(REG2_REG_12__SCAN_IN), .B1(n3963), .B2(
        n4953), .ZN(n3665) );
  NAND2_X1 U4521 ( .A1(n4619), .A2(n3965), .ZN(n3664) );
  OAI211_X1 U4522 ( .C1(n4864), .C2(n4572), .A(n3665), .B(n3664), .ZN(n3666)
         );
  AOI21_X1 U4523 ( .B1(n4787), .B2(n4577), .A(n3666), .ZN(n3667) );
  OAI21_X1 U4524 ( .B1(n3668), .B2(n2142), .A(n3667), .ZN(U3278) );
  OR2_X1 U4525 ( .A1(n3671), .A2(n3109), .ZN(n3669) );
  INV_X1 U4526 ( .A(n4883), .ZN(n3685) );
  XNOR2_X1 U4527 ( .A(n3679), .B(REG2_REG_12__SCAN_IN), .ZN(n3678) );
  INV_X1 U4528 ( .A(n3671), .ZN(n3673) );
  OAI211_X1 U4529 ( .C1(n3674), .C2(REG1_REG_12__SCAN_IN), .A(n3688), .B(n4935), .ZN(n3677) );
  AND2_X1 U4530 ( .A1(U3149), .A2(REG3_REG_12__SCAN_IN), .ZN(n3964) );
  NOR2_X1 U4531 ( .A1(n4949), .A2(n3685), .ZN(n3675) );
  AOI211_X1 U4532 ( .C1(n4942), .C2(ADDR_REG_12__SCAN_IN), .A(n3964), .B(n3675), .ZN(n3676) );
  OAI211_X1 U4533 ( .C1(n3678), .C2(n3705), .A(n3677), .B(n3676), .ZN(U3252)
         );
  NAND2_X1 U4534 ( .A1(n3679), .A2(REG2_REG_12__SCAN_IN), .ZN(n3682) );
  NAND2_X1 U4535 ( .A1(n3680), .A2(n4883), .ZN(n3681) );
  INV_X1 U4536 ( .A(REG2_REG_13__SCAN_IN), .ZN(n3683) );
  INV_X1 U4537 ( .A(n4882), .ZN(n3696) );
  AND2_X1 U4538 ( .A1(n4882), .A2(REG2_REG_13__SCAN_IN), .ZN(n3701) );
  AOI21_X1 U4539 ( .B1(n3683), .B2(n3696), .A(n3701), .ZN(n3684) );
  XNOR2_X1 U4540 ( .A(n3702), .B(n3684), .ZN(n3694) );
  OR2_X1 U4541 ( .A1(n3686), .A2(n3685), .ZN(n3687) );
  XNOR2_X1 U4542 ( .A(n4882), .B(n4782), .ZN(n3689) );
  OAI211_X1 U4543 ( .C1(n3690), .C2(n3689), .A(n3695), .B(n4935), .ZN(n3693)
         );
  AND2_X1 U4544 ( .A1(U3149), .A2(REG3_REG_13__SCAN_IN), .ZN(n4054) );
  NOR2_X1 U4545 ( .A1(n4949), .A2(n3696), .ZN(n3691) );
  AOI211_X1 U4546 ( .C1(n4942), .C2(ADDR_REG_13__SCAN_IN), .A(n4054), .B(n3691), .ZN(n3692) );
  OAI211_X1 U4547 ( .C1(n3694), .C2(n3705), .A(n3693), .B(n3692), .ZN(U3253)
         );
  OAI211_X1 U4548 ( .C1(n3697), .C2(REG1_REG_14__SCAN_IN), .A(n4318), .B(n4935), .ZN(n3711) );
  INV_X1 U4549 ( .A(n4949), .ZN(n4296) );
  INV_X1 U4550 ( .A(n3704), .ZN(n4327) );
  INV_X1 U4551 ( .A(n4942), .ZN(n3700) );
  AND2_X1 U4552 ( .A1(U3149), .A2(REG3_REG_14__SCAN_IN), .ZN(n3909) );
  INV_X1 U4553 ( .A(n3909), .ZN(n3698) );
  OAI21_X1 U4554 ( .B1(n3700), .B2(n3699), .A(n3698), .ZN(n3709) );
  INV_X1 U4555 ( .A(REG2_REG_14__SCAN_IN), .ZN(n3707) );
  OR2_X1 U4556 ( .A1(n4882), .A2(REG2_REG_13__SCAN_IN), .ZN(n3703) );
  AOI211_X1 U4557 ( .C1(n3707), .C2(n3706), .A(n3705), .B(n4326), .ZN(n3708)
         );
  AOI211_X1 U4558 ( .C1(n4296), .C2(n4327), .A(n3709), .B(n3708), .ZN(n3710)
         );
  NAND2_X1 U4559 ( .A1(n3711), .A2(n3710), .ZN(U3254) );
  NAND2_X1 U4560 ( .A1(n3712), .A2(U4043), .ZN(n3713) );
  OAI21_X1 U4561 ( .B1(U4043), .B2(n3714), .A(n3713), .ZN(U3552) );
  INV_X1 U4562 ( .A(n3715), .ZN(n3716) );
  AOI21_X1 U4563 ( .B1(n3718), .B2(n3717), .A(n3716), .ZN(n3723) );
  AOI22_X1 U4564 ( .A1(n4115), .A2(n4284), .B1(n4116), .B2(n3322), .ZN(n3719)
         );
  OAI21_X1 U4565 ( .B1(n4064), .B2(n3720), .A(n3719), .ZN(n3721) );
  AOI21_X1 U4566 ( .B1(REG3_REG_2__SCAN_IN), .B2(n3852), .A(n3721), .ZN(n3722)
         );
  OAI21_X1 U4567 ( .B1(n3723), .B2(n4108), .A(n3722), .ZN(U3234) );
  INV_X1 U4568 ( .A(DATAI_30_), .ZN(n3726) );
  NAND2_X1 U4569 ( .A1(n3724), .A2(STATE_REG_SCAN_IN), .ZN(n3725) );
  OAI21_X1 U4570 ( .B1(STATE_REG_SCAN_IN), .B2(n3726), .A(n3725), .ZN(U3322)
         );
  NAND2_X1 U4571 ( .A1(n4505), .A2(n3796), .ZN(n3728) );
  NAND2_X1 U4572 ( .A1(n3826), .A2(n4483), .ZN(n3727) );
  NAND2_X1 U4573 ( .A1(n3728), .A2(n3727), .ZN(n3729) );
  XNOR2_X1 U4574 ( .A(n3729), .B(n3871), .ZN(n3951) );
  INV_X1 U4575 ( .A(n3951), .ZN(n3807) );
  NOR2_X1 U4576 ( .A1(n3874), .A2(n4492), .ZN(n3730) );
  AOI21_X1 U4577 ( .B1(n4505), .B2(n3831), .A(n3730), .ZN(n3950) );
  INV_X1 U4578 ( .A(n3950), .ZN(n3806) );
  AOI22_X1 U4579 ( .A1(n3420), .A2(n4078), .B1(n3760), .B2(n3731), .ZN(n3749)
         );
  NAND2_X1 U4580 ( .A1(n4078), .A2(n3760), .ZN(n3733) );
  NAND2_X1 U4581 ( .A1(n3826), .A2(n3731), .ZN(n3732) );
  NAND2_X1 U4582 ( .A1(n3733), .A2(n3732), .ZN(n3734) );
  XNOR2_X1 U4583 ( .A(n3734), .B(n3841), .ZN(n3741) );
  NAND2_X1 U4584 ( .A1(n3420), .A2(n4280), .ZN(n3736) );
  NAND2_X1 U4585 ( .A1(n3760), .A2(n4688), .ZN(n3735) );
  NAND2_X1 U4586 ( .A1(n3736), .A2(n3735), .ZN(n3742) );
  INV_X1 U4587 ( .A(n3742), .ZN(n3932) );
  NAND2_X1 U4588 ( .A1(n4280), .A2(n3760), .ZN(n3739) );
  NAND2_X1 U4589 ( .A1(n3826), .A2(n4688), .ZN(n3738) );
  NAND2_X1 U4590 ( .A1(n3739), .A2(n3738), .ZN(n3740) );
  INV_X1 U4591 ( .A(n3926), .ZN(n3744) );
  OAI22_X1 U4592 ( .A1(n3932), .A2(n3933), .B1(n3744), .B2(n3930), .ZN(n3747)
         );
  XNOR2_X1 U4593 ( .A(n3741), .B(n3749), .ZN(n3935) );
  OAI21_X1 U4594 ( .B1(n3926), .B2(n3927), .A(n3742), .ZN(n3745) );
  NOR2_X1 U4595 ( .A1(n3742), .A2(n3927), .ZN(n3743) );
  NAND2_X1 U4596 ( .A1(n4279), .A2(n3796), .ZN(n3751) );
  NAND2_X1 U4597 ( .A1(n4079), .A2(n3826), .ZN(n3750) );
  NAND2_X1 U4598 ( .A1(n3751), .A2(n3750), .ZN(n3752) );
  XNOR2_X1 U4599 ( .A(n3752), .B(n3871), .ZN(n3754) );
  AOI22_X1 U4600 ( .A1(n3831), .A2(n4279), .B1(n3796), .B2(n4079), .ZN(n3753)
         );
  OR2_X1 U4601 ( .A1(n3754), .A2(n3753), .ZN(n4074) );
  AOI22_X1 U4602 ( .A1(n4632), .A2(n3755), .B1(n3965), .B2(n3826), .ZN(n3756)
         );
  AOI22_X1 U4603 ( .A1(n3831), .A2(n4632), .B1(n3965), .B2(n3760), .ZN(n3960)
         );
  NAND2_X1 U4604 ( .A1(n4278), .A2(n3760), .ZN(n3758) );
  NAND2_X1 U4605 ( .A1(n3826), .A2(n4639), .ZN(n3757) );
  NAND2_X1 U4606 ( .A1(n3758), .A2(n3757), .ZN(n3759) );
  XNOR2_X1 U4607 ( .A(n3759), .B(n3871), .ZN(n3762) );
  AOI22_X1 U4608 ( .A1(n3831), .A2(n4278), .B1(n4639), .B2(n3760), .ZN(n3761)
         );
  NOR2_X1 U4609 ( .A1(n3762), .A2(n3761), .ZN(n4048) );
  NAND2_X1 U4610 ( .A1(n3762), .A2(n3761), .ZN(n4049) );
  AOI22_X1 U4611 ( .A1(n4608), .A2(n3796), .B1(n3910), .B2(n3826), .ZN(n3763)
         );
  XNOR2_X1 U4612 ( .A(n3763), .B(n3841), .ZN(n3903) );
  AOI22_X1 U4613 ( .A1(n3831), .A2(n4608), .B1(n3910), .B2(n3760), .ZN(n3904)
         );
  INV_X1 U4614 ( .A(n3764), .ZN(n3985) );
  NAND2_X1 U4615 ( .A1(n3990), .A2(n3796), .ZN(n3766) );
  NAND2_X1 U4616 ( .A1(n3826), .A2(n4769), .ZN(n3765) );
  NAND2_X1 U4617 ( .A1(n3766), .A2(n3765), .ZN(n3767) );
  XNOR2_X1 U4618 ( .A(n3767), .B(n3841), .ZN(n3986) );
  NAND2_X1 U4619 ( .A1(n3990), .A2(n3831), .ZN(n3769) );
  NAND2_X1 U4620 ( .A1(n3796), .A2(n4769), .ZN(n3768) );
  NAND2_X1 U4621 ( .A1(n3769), .A2(n3768), .ZN(n3983) );
  NAND2_X1 U4622 ( .A1(n3986), .A2(n3983), .ZN(n3775) );
  OAI22_X1 U4623 ( .A1(n4609), .A2(n3874), .B1(n3873), .B2(n4594), .ZN(n3770)
         );
  XNOR2_X1 U4624 ( .A(n3770), .B(n3841), .ZN(n3997) );
  OR2_X1 U4625 ( .A1(n4609), .A2(n3870), .ZN(n3772) );
  NAND2_X1 U4626 ( .A1(n3796), .A2(n4763), .ZN(n3771) );
  NAND2_X1 U4627 ( .A1(n3772), .A2(n3771), .ZN(n3998) );
  NAND2_X1 U4628 ( .A1(n3997), .A2(n3998), .ZN(n3774) );
  OAI22_X1 U4629 ( .A1(n4584), .A2(n3874), .B1(n4561), .B2(n3873), .ZN(n3773)
         );
  XNOR2_X1 U4630 ( .A(n3773), .B(n3841), .ZN(n3999) );
  OAI22_X1 U4631 ( .A1(n4584), .A2(n3870), .B1(n4561), .B2(n3874), .ZN(n4000)
         );
  NAND2_X1 U4632 ( .A1(n3999), .A2(n4000), .ZN(n3776) );
  INV_X1 U4633 ( .A(n3776), .ZN(n3781) );
  INV_X1 U4634 ( .A(n3997), .ZN(n3988) );
  OAI21_X1 U4635 ( .B1(n3986), .B2(n3983), .A(n3998), .ZN(n3779) );
  NOR3_X1 U4636 ( .A1(n3986), .A2(n3998), .A3(n3983), .ZN(n3778) );
  NOR2_X1 U4637 ( .A1(n3999), .A2(n4000), .ZN(n3777) );
  AOI211_X1 U4638 ( .C1(n3988), .C2(n3779), .A(n3778), .B(n3777), .ZN(n3780)
         );
  NAND2_X1 U4639 ( .A1(n4564), .A2(n3760), .ZN(n3783) );
  NAND2_X1 U4640 ( .A1(n3826), .A2(n4092), .ZN(n3782) );
  NAND2_X1 U4641 ( .A1(n3783), .A2(n3782), .ZN(n3784) );
  XNOR2_X1 U4642 ( .A(n3784), .B(n3841), .ZN(n3788) );
  NAND2_X1 U4643 ( .A1(n4564), .A2(n3831), .ZN(n3786) );
  NAND2_X1 U4644 ( .A1(n3796), .A2(n4092), .ZN(n3785) );
  NAND2_X1 U4645 ( .A1(n3786), .A2(n3785), .ZN(n3787) );
  NAND2_X1 U4646 ( .A1(n3788), .A2(n3787), .ZN(n4086) );
  NOR2_X1 U4647 ( .A1(n3788), .A2(n3787), .ZN(n4088) );
  NAND2_X1 U4648 ( .A1(n4545), .A2(n3760), .ZN(n3790) );
  NAND2_X1 U4649 ( .A1(n3826), .A2(n4527), .ZN(n3789) );
  NAND2_X1 U4650 ( .A1(n3790), .A2(n3789), .ZN(n3791) );
  XNOR2_X1 U4651 ( .A(n3791), .B(n3841), .ZN(n3794) );
  AOI22_X1 U4652 ( .A1(n4545), .A2(n3831), .B1(n4527), .B2(n3760), .ZN(n3792)
         );
  XOR2_X1 U4653 ( .A(n3794), .B(n3792), .Z(n3942) );
  INV_X1 U4654 ( .A(n3792), .ZN(n3793) );
  NAND2_X1 U4655 ( .A1(n4484), .A2(n3796), .ZN(n3798) );
  NAND2_X1 U4656 ( .A1(n3826), .A2(n4745), .ZN(n3797) );
  NAND2_X1 U4657 ( .A1(n3798), .A2(n3797), .ZN(n3799) );
  XNOR2_X1 U4658 ( .A(n3799), .B(n3841), .ZN(n3802) );
  NAND2_X1 U4659 ( .A1(n4484), .A2(n3831), .ZN(n3801) );
  NAND2_X1 U4660 ( .A1(n3760), .A2(n4745), .ZN(n3800) );
  NAND2_X1 U4661 ( .A1(n3801), .A2(n3800), .ZN(n3803) );
  NAND2_X1 U4662 ( .A1(n3802), .A2(n3803), .ZN(n4038) );
  INV_X1 U4663 ( .A(n3802), .ZN(n3805) );
  INV_X1 U4664 ( .A(n3803), .ZN(n3804) );
  NAND2_X1 U4665 ( .A1(n3805), .A2(n3804), .ZN(n4040) );
  OAI22_X1 U4666 ( .A1(n4487), .A2(n3870), .B1(n4465), .B2(n3874), .ZN(n3812)
         );
  OAI22_X1 U4667 ( .A1(n4487), .A2(n3874), .B1(n4465), .B2(n3873), .ZN(n3808)
         );
  XNOR2_X1 U4668 ( .A(n3808), .B(n3841), .ZN(n3813) );
  XOR2_X1 U4669 ( .A(n3812), .B(n3813), .Z(n4062) );
  OAI22_X1 U4670 ( .A1(n4068), .A2(n3874), .B1(n4457), .B2(n3873), .ZN(n3809)
         );
  XNOR2_X1 U4671 ( .A(n3809), .B(n3871), .ZN(n3815) );
  OR2_X1 U4672 ( .A1(n4068), .A2(n3870), .ZN(n3811) );
  NAND2_X1 U4673 ( .A1(n3755), .A2(n4451), .ZN(n3810) );
  NAND2_X1 U4674 ( .A1(n3811), .A2(n3810), .ZN(n3816) );
  XNOR2_X1 U4675 ( .A(n3815), .B(n3816), .ZN(n3918) );
  OR2_X1 U4676 ( .A1(n3813), .A2(n3812), .ZN(n3919) );
  INV_X1 U4677 ( .A(n3815), .ZN(n3817) );
  NAND2_X1 U4678 ( .A1(n3817), .A2(n3816), .ZN(n3821) );
  NOR2_X1 U4679 ( .A1(n3874), .A2(n4440), .ZN(n3818) );
  AOI21_X1 U4680 ( .B1(n4415), .B2(n3420), .A(n3818), .ZN(n3822) );
  OAI22_X1 U4681 ( .A1(n4455), .A2(n3874), .B1(n4440), .B2(n3873), .ZN(n3820)
         );
  XNOR2_X1 U4682 ( .A(n3820), .B(n3841), .ZN(n4011) );
  INV_X1 U4683 ( .A(n3822), .ZN(n3823) );
  NAND2_X1 U4684 ( .A1(n3824), .A2(n3823), .ZN(n4009) );
  NAND2_X1 U4685 ( .A1(n4399), .A2(n3796), .ZN(n3828) );
  NAND2_X1 U4686 ( .A1(n3826), .A2(n4414), .ZN(n3827) );
  NAND2_X1 U4687 ( .A1(n3828), .A2(n3827), .ZN(n3829) );
  XNOR2_X1 U4688 ( .A(n3829), .B(n3871), .ZN(n3833) );
  NOR2_X1 U4689 ( .A1(n3874), .A2(n4421), .ZN(n3830) );
  AOI21_X1 U4690 ( .B1(n4399), .B2(n3831), .A(n3830), .ZN(n3832) );
  NAND2_X1 U4691 ( .A1(n3833), .A2(n3832), .ZN(n3973) );
  NOR2_X1 U4692 ( .A1(n3833), .A2(n3832), .ZN(n3974) );
  OAI22_X1 U4693 ( .A1(n4418), .A2(n3874), .B1(n3873), .B2(n4720), .ZN(n3834)
         );
  XNOR2_X1 U4694 ( .A(n3834), .B(n3841), .ZN(n3837) );
  OR2_X1 U4695 ( .A1(n4418), .A2(n3870), .ZN(n3836) );
  NAND2_X1 U4696 ( .A1(n3796), .A2(n2207), .ZN(n3835) );
  NAND2_X1 U4697 ( .A1(n3836), .A2(n3835), .ZN(n3838) );
  NAND2_X1 U4698 ( .A1(n3837), .A2(n3838), .ZN(n4099) );
  INV_X1 U4699 ( .A(n3837), .ZN(n3840) );
  INV_X1 U4700 ( .A(n3838), .ZN(n3839) );
  NAND2_X1 U4701 ( .A1(n3840), .A2(n3839), .ZN(n4100) );
  OAI22_X1 U4702 ( .A1(n3887), .A2(n3874), .B1(n3873), .B2(n4384), .ZN(n3842)
         );
  XNOR2_X1 U4703 ( .A(n3842), .B(n3841), .ZN(n3883) );
  OAI22_X1 U4704 ( .A1(n3887), .A2(n3870), .B1(n3874), .B2(n4384), .ZN(n3882)
         );
  XNOR2_X1 U4705 ( .A(n3883), .B(n3882), .ZN(n3878) );
  XNOR2_X1 U4706 ( .A(n3843), .B(n3878), .ZN(n3848) );
  NOR2_X1 U4707 ( .A1(n4386), .A2(n4120), .ZN(n3846) );
  AOI22_X1 U4708 ( .A1(n4117), .A2(n4714), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n3844) );
  OAI21_X1 U4709 ( .B1(n4369), .B2(n4067), .A(n3844), .ZN(n3845) );
  AOI211_X1 U4710 ( .C1(n4116), .C2(n4391), .A(n3846), .B(n3845), .ZN(n3847)
         );
  OAI21_X1 U4711 ( .B1(n3848), .B2(n4108), .A(n3847), .ZN(U3211) );
  INV_X1 U4712 ( .A(n3849), .ZN(n3850) );
  XNOR2_X1 U4713 ( .A(n3851), .B(n3850), .ZN(n4286) );
  AOI22_X1 U4714 ( .A1(n4286), .A2(n4122), .B1(n4115), .B2(n3322), .ZN(n3854)
         );
  NAND2_X1 U4715 ( .A1(n3852), .A2(REG3_REG_0__SCAN_IN), .ZN(n3853) );
  OAI211_X1 U4716 ( .C1(n4064), .C2(n3855), .A(n3854), .B(n3853), .ZN(U3229)
         );
  OR2_X1 U4717 ( .A1(n4596), .A2(n4200), .ZN(n4614) );
  INV_X1 U4718 ( .A(n4614), .ZN(n3856) );
  AOI21_X1 U4719 ( .B1(n4200), .B2(n4596), .A(n3856), .ZN(n4775) );
  INV_X1 U4720 ( .A(n3990), .ZN(n4583) );
  XOR2_X1 U4721 ( .A(n4233), .B(n4200), .Z(n3857) );
  OAI222_X1 U4722 ( .A1(n4659), .A2(n3858), .B1(n4678), .B2(n4583), .C1(n3857), 
        .C2(n4684), .ZN(n4777) );
  NAND2_X1 U4723 ( .A1(n4777), .A2(n4957), .ZN(n3865) );
  INV_X1 U4724 ( .A(n4642), .ZN(n3860) );
  INV_X1 U4725 ( .A(n4620), .ZN(n3859) );
  OAI21_X1 U4726 ( .B1(n3860), .B2(n4774), .A(n3859), .ZN(n4856) );
  INV_X1 U4727 ( .A(n4856), .ZN(n3863) );
  AOI22_X1 U4728 ( .A1(n2142), .A2(REG2_REG_14__SCAN_IN), .B1(n3908), .B2(
        n4953), .ZN(n3861) );
  OAI21_X1 U4729 ( .B1(n4666), .B2(n4774), .A(n3861), .ZN(n3862) );
  AOI21_X1 U4730 ( .B1(n3863), .B2(n4693), .A(n3862), .ZN(n3864) );
  OAI211_X1 U4731 ( .C1(n4697), .C2(n4775), .A(n3865), .B(n3864), .ZN(U3276)
         );
  NAND3_X1 U4732 ( .A1(n3867), .A2(IR_REG_31__SCAN_IN), .A3(STATE_REG_SCAN_IN), 
        .ZN(n3869) );
  OAI22_X1 U4733 ( .A1(n3866), .A2(n3869), .B1(STATE_REG_SCAN_IN), .B2(n3868), 
        .ZN(U3321) );
  OAI22_X1 U4734 ( .A1(n4369), .A2(n3870), .B1(n4358), .B2(n3874), .ZN(n3872)
         );
  XNOR2_X1 U4735 ( .A(n3872), .B(n3871), .ZN(n3876) );
  OAI22_X1 U4736 ( .A1(n4369), .A2(n3874), .B1(n4358), .B2(n3873), .ZN(n3875)
         );
  XNOR2_X1 U4737 ( .A(n3876), .B(n3875), .ZN(n3889) );
  INV_X1 U4738 ( .A(n3889), .ZN(n3877) );
  NAND2_X1 U4739 ( .A1(n3877), .A2(n4122), .ZN(n3893) );
  INV_X1 U4740 ( .A(n3878), .ZN(n3879) );
  AND2_X1 U4741 ( .A1(n4100), .A2(n3879), .ZN(n3880) );
  NAND2_X1 U4742 ( .A1(n3883), .A2(n3882), .ZN(n3888) );
  AOI22_X1 U4743 ( .A1(n4117), .A2(n3895), .B1(REG3_REG_28__SCAN_IN), .B2(
        U3149), .ZN(n3886) );
  NAND2_X1 U4744 ( .A1(n4276), .A2(n4115), .ZN(n3885) );
  OAI211_X1 U4745 ( .C1(n3887), .C2(n4065), .A(n3886), .B(n3885), .ZN(n3891)
         );
  NOR3_X1 U4746 ( .A1(n3889), .A2(n4108), .A3(n3888), .ZN(n3890) );
  AOI211_X1 U4747 ( .C1(n3894), .C2(n4102), .A(n3891), .B(n3890), .ZN(n3892)
         );
  AOI22_X1 U4748 ( .A1(n3894), .A2(n4953), .B1(REG2_REG_28__SCAN_IN), .B2(
        n2142), .ZN(n3897) );
  NAND2_X1 U4749 ( .A1(n4619), .A2(n3895), .ZN(n3896) );
  OAI211_X1 U4750 ( .C1(n3898), .C2(n4572), .A(n3897), .B(n3896), .ZN(n3899)
         );
  AOI21_X1 U4751 ( .B1(n3900), .B2(n4957), .A(n3899), .ZN(n3901) );
  OAI21_X1 U4752 ( .B1(n3902), .B2(n4697), .A(n3901), .ZN(U3262) );
  INV_X1 U4753 ( .A(n3903), .ZN(n3905) );
  XNOR2_X1 U4754 ( .A(n3905), .B(n3904), .ZN(n3906) );
  XNOR2_X1 U4755 ( .A(n3907), .B(n3906), .ZN(n3915) );
  INV_X1 U4756 ( .A(n3908), .ZN(n3913) );
  AOI21_X1 U4757 ( .B1(n4116), .B2(n4278), .A(n3909), .ZN(n3912) );
  AOI22_X1 U4758 ( .A1(n4115), .A2(n3990), .B1(n4117), .B2(n3910), .ZN(n3911)
         );
  OAI211_X1 U4759 ( .C1(n4120), .C2(n3913), .A(n3912), .B(n3911), .ZN(n3914)
         );
  AOI21_X1 U4760 ( .B1(n3915), .B2(n4122), .A(n3914), .ZN(n3916) );
  INV_X1 U4761 ( .A(n3916), .ZN(U3212) );
  NAND2_X1 U4762 ( .A1(n3917), .A2(n4122), .ZN(n3925) );
  AOI21_X1 U4763 ( .B1(n4060), .B2(n3919), .A(n3918), .ZN(n3924) );
  OAI22_X1 U4764 ( .A1(n4487), .A2(n4065), .B1(STATE_REG_SCAN_IN), .B2(n3920), 
        .ZN(n3922) );
  OAI22_X1 U4765 ( .A1(n4455), .A2(n4067), .B1(n4064), .B2(n4457), .ZN(n3921)
         );
  AOI211_X1 U4766 ( .C1(n4458), .C2(n4102), .A(n3922), .B(n3921), .ZN(n3923)
         );
  OAI21_X1 U4767 ( .B1(n3925), .B2(n3924), .A(n3923), .ZN(U3213) );
  INV_X1 U4768 ( .A(n3928), .ZN(n3931) );
  OAI21_X1 U4769 ( .B1(n3928), .B2(n3927), .A(n3926), .ZN(n3929) );
  OAI21_X1 U4770 ( .B1(n3931), .B2(n3930), .A(n3929), .ZN(n4030) );
  XNOR2_X1 U4771 ( .A(n3933), .B(n3932), .ZN(n4031) );
  NOR2_X1 U4772 ( .A1(n4030), .A2(n4031), .ZN(n4029) );
  AOI21_X1 U4773 ( .B1(n3933), .B2(n3932), .A(n4029), .ZN(n3936) );
  OAI211_X1 U4774 ( .C1(n3936), .C2(n3935), .A(n4122), .B(n3934), .ZN(n3940)
         );
  OAI22_X1 U4775 ( .A1(n4064), .A2(n4794), .B1(n4660), .B2(n4067), .ZN(n3937)
         );
  AOI211_X1 U4776 ( .C1(n4116), .C2(n4280), .A(n3938), .B(n3937), .ZN(n3939)
         );
  OAI211_X1 U4777 ( .C1(n4120), .C2(n3941), .A(n3940), .B(n3939), .ZN(U3214)
         );
  XNOR2_X1 U4778 ( .A(n3943), .B(n3942), .ZN(n3948) );
  NAND2_X1 U4779 ( .A1(U3149), .A2(REG3_REG_19__SCAN_IN), .ZN(n4338) );
  INV_X1 U4780 ( .A(n4338), .ZN(n3944) );
  AOI21_X1 U4781 ( .B1(n4115), .B2(n4484), .A(n3944), .ZN(n3946) );
  AOI22_X1 U4782 ( .A1(n4527), .A2(n4117), .B1(n4116), .B2(n4564), .ZN(n3945)
         );
  OAI211_X1 U4783 ( .C1(n4120), .C2(n4536), .A(n3946), .B(n3945), .ZN(n3947)
         );
  AOI21_X1 U4784 ( .B1(n3948), .B2(n4122), .A(n3947), .ZN(n3949) );
  INV_X1 U4785 ( .A(n3949), .ZN(U3216) );
  XNOR2_X1 U4786 ( .A(n3951), .B(n3950), .ZN(n3952) );
  XNOR2_X1 U4787 ( .A(n3953), .B(n3952), .ZN(n3959) );
  INV_X1 U4788 ( .A(n4490), .ZN(n3957) );
  OAI22_X1 U4789 ( .A1(n4530), .A2(n4065), .B1(n4064), .B2(n4492), .ZN(n3956)
         );
  OAI22_X1 U4790 ( .A1(n4487), .A2(n4067), .B1(STATE_REG_SCAN_IN), .B2(n3954), 
        .ZN(n3955) );
  AOI211_X1 U4791 ( .C1(n3957), .C2(n4102), .A(n3956), .B(n3955), .ZN(n3958)
         );
  OAI21_X1 U4792 ( .B1(n3959), .B2(n4108), .A(n3958), .ZN(U3220) );
  XNOR2_X1 U4793 ( .A(n2152), .B(n3960), .ZN(n3961) );
  XNOR2_X1 U4794 ( .A(n3962), .B(n3961), .ZN(n3970) );
  INV_X1 U4795 ( .A(n3963), .ZN(n3968) );
  AOI21_X1 U4796 ( .B1(n4116), .B2(n4279), .A(n3964), .ZN(n3967) );
  AOI22_X1 U4797 ( .A1(n4115), .A2(n4278), .B1(n4117), .B2(n3965), .ZN(n3966)
         );
  OAI211_X1 U4798 ( .C1(n4120), .C2(n3968), .A(n3967), .B(n3966), .ZN(n3969)
         );
  AOI21_X1 U4799 ( .B1(n3970), .B2(n4122), .A(n3969), .ZN(n3971) );
  INV_X1 U4800 ( .A(n3971), .ZN(U3221) );
  NOR2_X1 U4801 ( .A1(n3974), .A2(n2274), .ZN(n3975) );
  XNOR2_X1 U4802 ( .A(n3976), .B(n3975), .ZN(n3982) );
  OAI22_X1 U4803 ( .A1(n4455), .A2(n4065), .B1(STATE_REG_SCAN_IN), .B2(n3977), 
        .ZN(n3978) );
  AOI21_X1 U4804 ( .B1(n4414), .B2(n4117), .A(n3978), .ZN(n3979) );
  OAI21_X1 U4805 ( .B1(n4120), .B2(n4423), .A(n3979), .ZN(n3980) );
  AOI21_X1 U4806 ( .B1(n4115), .B2(n4391), .A(n3980), .ZN(n3981) );
  OAI21_X1 U4807 ( .B1(n3982), .B2(n4108), .A(n3981), .ZN(U3222) );
  INV_X1 U4808 ( .A(n3983), .ZN(n4113) );
  NAND2_X1 U4809 ( .A1(n3985), .A2(n3984), .ZN(n3987) );
  NAND2_X1 U4810 ( .A1(n3987), .A2(n3986), .ZN(n4110) );
  NOR2_X1 U4811 ( .A1(n3987), .A2(n3986), .ZN(n4112) );
  AOI21_X1 U4812 ( .B1(n4113), .B2(n4110), .A(n4112), .ZN(n3989) );
  XNOR2_X1 U4813 ( .A(n3988), .B(n3998), .ZN(n3995) );
  XNOR2_X1 U4814 ( .A(n3989), .B(n3995), .ZN(n3994) );
  AOI22_X1 U4815 ( .A1(n4763), .A2(n4117), .B1(n4116), .B2(n3990), .ZN(n3991)
         );
  NAND2_X1 U4816 ( .A1(U3149), .A2(REG3_REG_16__SCAN_IN), .ZN(n4914) );
  OAI211_X1 U4817 ( .C1(n4584), .C2(n4067), .A(n3991), .B(n4914), .ZN(n3992)
         );
  AOI21_X1 U4818 ( .B1(n4592), .B2(n4102), .A(n3992), .ZN(n3993) );
  OAI21_X1 U4819 ( .B1(n3994), .B2(n4108), .A(n3993), .ZN(U3223) );
  OAI211_X1 U4820 ( .C1(n4112), .C2(n4113), .A(n3995), .B(n4110), .ZN(n3996)
         );
  OAI21_X1 U4821 ( .B1(n3998), .B2(n3997), .A(n3996), .ZN(n4002) );
  XOR2_X1 U4822 ( .A(n4000), .B(n3999), .Z(n4001) );
  XNOR2_X1 U4823 ( .A(n4002), .B(n4001), .ZN(n4006) );
  AND2_X1 U4824 ( .A1(U3149), .A2(REG3_REG_17__SCAN_IN), .ZN(n4926) );
  AOI21_X1 U4825 ( .B1(n4116), .B2(n4277), .A(n4926), .ZN(n4004) );
  AOI22_X1 U4826 ( .A1(n4115), .A2(n4564), .B1(n4117), .B2(n4569), .ZN(n4003)
         );
  OAI211_X1 U4827 ( .C1(n4120), .C2(n4573), .A(n4004), .B(n4003), .ZN(n4005)
         );
  AOI21_X1 U4828 ( .B1(n4006), .B2(n4122), .A(n4005), .ZN(n4007) );
  INV_X1 U4829 ( .A(n4007), .ZN(U3225) );
  NAND2_X1 U4830 ( .A1(n4009), .A2(n4008), .ZN(n4010) );
  XOR2_X1 U4831 ( .A(n4011), .B(n4010), .Z(n4017) );
  OAI22_X1 U4832 ( .A1(n4068), .A2(n4065), .B1(STATE_REG_SCAN_IN), .B2(n4012), 
        .ZN(n4013) );
  AOI21_X1 U4833 ( .B1(n4435), .B2(n4117), .A(n4013), .ZN(n4014) );
  OAI21_X1 U4834 ( .B1(n4438), .B2(n4067), .A(n4014), .ZN(n4015) );
  AOI21_X1 U4835 ( .B1(n4442), .B2(n4102), .A(n4015), .ZN(n4016) );
  OAI21_X1 U4836 ( .B1(n4017), .B2(n4108), .A(n4016), .ZN(U3226) );
  AND2_X1 U4837 ( .A1(n4019), .A2(n4018), .ZN(n4022) );
  OAI211_X1 U4838 ( .C1(n4022), .C2(n4021), .A(n4122), .B(n4020), .ZN(n4028)
         );
  AND2_X1 U4839 ( .A1(U3149), .A2(REG3_REG_4__SCAN_IN), .ZN(n4895) );
  AOI21_X1 U4840 ( .B1(n4115), .B2(n4283), .A(n4895), .ZN(n4027) );
  AOI22_X1 U4841 ( .A1(n4023), .A2(n4117), .B1(n4116), .B2(n4284), .ZN(n4026)
         );
  OR2_X1 U4842 ( .A1(n4120), .A2(n4024), .ZN(n4025) );
  NAND4_X1 U4843 ( .A1(n4028), .A2(n4027), .A3(n4026), .A4(n4025), .ZN(U3227)
         );
  AOI21_X1 U4844 ( .B1(n4031), .B2(n4030), .A(n4029), .ZN(n4035) );
  NOR2_X1 U4845 ( .A1(STATE_REG_SCAN_IN), .A2(n2610), .ZN(n4308) );
  INV_X1 U4846 ( .A(n4078), .ZN(n4679) );
  OAI22_X1 U4847 ( .A1(n4064), .A2(n2309), .B1(n4679), .B2(n4067), .ZN(n4032)
         );
  AOI211_X1 U4848 ( .C1(n4116), .C2(n4681), .A(n4308), .B(n4032), .ZN(n4034)
         );
  NAND2_X1 U4849 ( .A1(n4102), .A2(n4692), .ZN(n4033) );
  OAI211_X1 U4850 ( .C1(n4035), .C2(n4108), .A(n4034), .B(n4033), .ZN(U3228)
         );
  INV_X1 U4851 ( .A(n4036), .ZN(n4041) );
  AOI21_X1 U4852 ( .B1(n4040), .B2(n4038), .A(n4037), .ZN(n4039) );
  AOI21_X1 U4853 ( .B1(n4041), .B2(n4040), .A(n4039), .ZN(n4046) );
  AOI22_X1 U4854 ( .A1(n4505), .A2(n4115), .B1(REG3_REG_20__SCAN_IN), .B2(
        U3149), .ZN(n4043) );
  AOI22_X1 U4855 ( .A1(n4745), .A2(n4117), .B1(n4116), .B2(n4545), .ZN(n4042)
         );
  OAI211_X1 U4856 ( .C1(n4120), .C2(n4510), .A(n4043), .B(n4042), .ZN(n4044)
         );
  INV_X1 U4857 ( .A(n4044), .ZN(n4045) );
  OAI21_X1 U4858 ( .B1(n4046), .B2(n4108), .A(n4045), .ZN(U3230) );
  INV_X1 U4859 ( .A(n4048), .ZN(n4050) );
  NAND2_X1 U4860 ( .A1(n4050), .A2(n4049), .ZN(n4051) );
  XNOR2_X1 U4861 ( .A(n4052), .B(n4051), .ZN(n4058) );
  INV_X1 U4862 ( .A(n4053), .ZN(n4644) );
  AOI21_X1 U4863 ( .B1(n4116), .B2(n4632), .A(n4054), .ZN(n4056) );
  AOI22_X1 U4864 ( .A1(n4115), .A2(n4608), .B1(n4117), .B2(n4639), .ZN(n4055)
         );
  OAI211_X1 U4865 ( .C1(n4120), .C2(n4644), .A(n4056), .B(n4055), .ZN(n4057)
         );
  AOI21_X1 U4866 ( .B1(n4058), .B2(n4122), .A(n4057), .ZN(n4059) );
  INV_X1 U4867 ( .A(n4059), .ZN(U3231) );
  OAI21_X1 U4868 ( .B1(n4062), .B2(n4061), .A(n4060), .ZN(n4063) );
  NAND2_X1 U4869 ( .A1(n4063), .A2(n4122), .ZN(n4072) );
  OAI22_X1 U4870 ( .A1(n4466), .A2(n4065), .B1(n4064), .B2(n4465), .ZN(n4070)
         );
  OAI22_X1 U4871 ( .A1(n4068), .A2(n4067), .B1(STATE_REG_SCAN_IN), .B2(n4066), 
        .ZN(n4069) );
  AOI211_X1 U4872 ( .C1(n4474), .C2(n4102), .A(n4070), .B(n4069), .ZN(n4071)
         );
  NAND2_X1 U4873 ( .A1(n4072), .A2(n4071), .ZN(U3232) );
  NAND2_X1 U4874 ( .A1(n2449), .A2(n4074), .ZN(n4075) );
  XNOR2_X1 U4875 ( .A(n4073), .B(n4075), .ZN(n4084) );
  INV_X1 U4876 ( .A(n4076), .ZN(n4082) );
  AOI21_X1 U4877 ( .B1(n4116), .B2(n4078), .A(n4077), .ZN(n4081) );
  AOI22_X1 U4878 ( .A1(n4115), .A2(n4632), .B1(n4117), .B2(n4079), .ZN(n4080)
         );
  OAI211_X1 U4879 ( .C1(n4120), .C2(n4082), .A(n4081), .B(n4080), .ZN(n4083)
         );
  AOI21_X1 U4880 ( .B1(n4084), .B2(n4122), .A(n4083), .ZN(n4085) );
  INV_X1 U4881 ( .A(n4085), .ZN(U3233) );
  INV_X1 U4882 ( .A(n4086), .ZN(n4087) );
  NOR2_X1 U4883 ( .A1(n4088), .A2(n4087), .ZN(n4089) );
  XNOR2_X1 U4884 ( .A(n4090), .B(n4089), .ZN(n4096) );
  AND2_X1 U4885 ( .A1(U3149), .A2(REG3_REG_18__SCAN_IN), .ZN(n4941) );
  AOI21_X1 U4886 ( .B1(n4116), .B2(n4091), .A(n4941), .ZN(n4094) );
  AOI22_X1 U4887 ( .A1(n4115), .A2(n4545), .B1(n4117), .B2(n4092), .ZN(n4093)
         );
  OAI211_X1 U4888 ( .C1(n4120), .C2(n4555), .A(n4094), .B(n4093), .ZN(n4095)
         );
  AOI21_X1 U4889 ( .B1(n4096), .B2(n4122), .A(n4095), .ZN(n4097) );
  INV_X1 U4890 ( .A(n4097), .ZN(U3235) );
  NAND2_X1 U4891 ( .A1(n4100), .A2(n4099), .ZN(n4101) );
  XNOR2_X1 U4892 ( .A(n4098), .B(n4101), .ZN(n4109) );
  NAND2_X1 U4893 ( .A1(n4400), .A2(n4115), .ZN(n4106) );
  AOI22_X1 U4894 ( .A1(n4117), .A2(n2207), .B1(REG3_REG_26__SCAN_IN), .B2(
        U3149), .ZN(n4105) );
  NAND2_X1 U4895 ( .A1(n4407), .A2(n4102), .ZN(n4104) );
  NAND2_X1 U4896 ( .A1(n4399), .A2(n4116), .ZN(n4103) );
  OAI21_X1 U4897 ( .B1(n4109), .B2(n4108), .A(n4107), .ZN(U3237) );
  INV_X1 U4898 ( .A(n4110), .ZN(n4111) );
  NOR2_X1 U4899 ( .A1(n4112), .A2(n4111), .ZN(n4114) );
  XNOR2_X1 U4900 ( .A(n4114), .B(n4113), .ZN(n4123) );
  AND2_X1 U4901 ( .A1(U3149), .A2(REG3_REG_15__SCAN_IN), .ZN(n4907) );
  AOI21_X1 U4902 ( .B1(n4115), .B2(n4277), .A(n4907), .ZN(n4119) );
  AOI22_X1 U4903 ( .A1(n4769), .A2(n4117), .B1(n4116), .B2(n4608), .ZN(n4118)
         );
  OAI211_X1 U4904 ( .C1(n4120), .C2(n4617), .A(n4119), .B(n4118), .ZN(n4121)
         );
  AOI21_X1 U4905 ( .B1(n4123), .B2(n4122), .A(n4121), .ZN(n4124) );
  INV_X1 U4906 ( .A(n4124), .ZN(U3238) );
  NAND2_X1 U4907 ( .A1(n4126), .A2(n4125), .ZN(n4129) );
  NAND3_X1 U4908 ( .A1(n4129), .A2(n4128), .A3(n4127), .ZN(n4132) );
  NAND3_X1 U4909 ( .A1(n4132), .A2(n4131), .A3(n4130), .ZN(n4135) );
  NAND3_X1 U4910 ( .A1(n4135), .A2(n4134), .A3(n4133), .ZN(n4138) );
  NAND3_X1 U4911 ( .A1(n4138), .A2(n4137), .A3(n4136), .ZN(n4141) );
  NAND4_X1 U4912 ( .A1(n4141), .A2(n4140), .A3(n4152), .A4(n4139), .ZN(n4143)
         );
  NAND3_X1 U4913 ( .A1(n4143), .A2(n4222), .A3(n4142), .ZN(n4145) );
  AND2_X1 U4914 ( .A1(n4144), .A2(n4674), .ZN(n4154) );
  NAND2_X1 U4915 ( .A1(n4145), .A2(n4154), .ZN(n4146) );
  NAND3_X1 U4916 ( .A1(n4146), .A2(n4217), .A3(n4672), .ZN(n4158) );
  NAND2_X1 U4917 ( .A1(n4148), .A2(n4147), .ZN(n4150) );
  NOR2_X1 U4918 ( .A1(n4150), .A2(n4149), .ZN(n4157) );
  NAND2_X1 U4919 ( .A1(n4150), .A2(n4162), .ZN(n4231) );
  INV_X1 U4920 ( .A(n4151), .ZN(n4153) );
  NAND4_X1 U4921 ( .A1(n4154), .A2(n4218), .A3(n4153), .A4(n4152), .ZN(n4155)
         );
  NAND2_X1 U4922 ( .A1(n4155), .A2(n4209), .ZN(n4156) );
  AOI22_X1 U4923 ( .A1(n4158), .A2(n4157), .B1(n4231), .B2(n4156), .ZN(n4169)
         );
  NAND3_X1 U4924 ( .A1(n4160), .A2(n4159), .A3(n4208), .ZN(n4168) );
  NAND2_X1 U4925 ( .A1(n4162), .A2(n4161), .ZN(n4232) );
  INV_X1 U4926 ( .A(n4232), .ZN(n4163) );
  OAI211_X1 U4927 ( .C1(n4165), .C2(n2248), .A(n4164), .B(n4163), .ZN(n4166)
         );
  NAND2_X1 U4928 ( .A1(n4166), .A2(n4231), .ZN(n4167) );
  OAI21_X1 U4929 ( .B1(n4169), .B2(n4168), .A(n4167), .ZN(n4171) );
  INV_X1 U4930 ( .A(n4237), .ZN(n4170) );
  AOI21_X1 U4931 ( .B1(n4171), .B2(n4234), .A(n4170), .ZN(n4173) );
  OR3_X1 U4932 ( .A1(n4173), .A2(n4172), .A3(n4235), .ZN(n4176) );
  INV_X1 U4933 ( .A(n4174), .ZN(n4242) );
  AOI21_X1 U4934 ( .B1(n4176), .B2(n4175), .A(n4242), .ZN(n4180) );
  NAND3_X1 U4935 ( .A1(n4245), .A2(n4244), .A3(n2426), .ZN(n4179) );
  INV_X1 U4936 ( .A(n4396), .ZN(n4203) );
  NAND2_X1 U4937 ( .A1(n4245), .A2(n2165), .ZN(n4177) );
  NAND3_X1 U4938 ( .A1(n4203), .A2(n4196), .A3(n4177), .ZN(n4252) );
  INV_X1 U4939 ( .A(n4252), .ZN(n4178) );
  OAI21_X1 U4940 ( .B1(n4180), .B2(n4179), .A(n4178), .ZN(n4184) );
  AND2_X1 U4941 ( .A1(n2144), .A2(DATAI_29_), .ZN(n4375) );
  INV_X1 U4942 ( .A(n4375), .ZN(n4706) );
  INV_X1 U4943 ( .A(n4364), .ZN(n4181) );
  AOI21_X1 U4944 ( .B1(n4276), .B2(n4706), .A(n4181), .ZN(n4255) );
  NAND3_X1 U4945 ( .A1(n4255), .A2(n4254), .A3(n4182), .ZN(n4183) );
  AOI21_X1 U4946 ( .B1(n4251), .B2(n4184), .A(n4183), .ZN(n4190) );
  NAND2_X1 U4947 ( .A1(n4362), .A2(n4185), .ZN(n4249) );
  OR2_X1 U4948 ( .A1(n4276), .A2(n4706), .ZN(n4188) );
  NAND2_X1 U4949 ( .A1(n2144), .A2(DATAI_31_), .ZN(n4346) );
  NAND2_X1 U4950 ( .A1(n4345), .A2(n4346), .ZN(n4193) );
  AND2_X1 U4951 ( .A1(n2144), .A2(DATAI_30_), .ZN(n4350) );
  INV_X1 U4952 ( .A(n4350), .ZN(n4191) );
  OR2_X1 U4953 ( .A1(n4360), .A2(n4191), .ZN(n4187) );
  AND2_X1 U4954 ( .A1(n4193), .A2(n4187), .ZN(n4206) );
  NAND2_X1 U4955 ( .A1(n4188), .A2(n4206), .ZN(n4248) );
  AOI21_X1 U4956 ( .B1(n4255), .B2(n4249), .A(n4248), .ZN(n4257) );
  INV_X1 U4957 ( .A(n4257), .ZN(n4189) );
  NOR2_X1 U4958 ( .A1(n4190), .A2(n4189), .ZN(n4195) );
  NAND2_X1 U4959 ( .A1(n4360), .A2(n4191), .ZN(n4261) );
  OR2_X1 U4960 ( .A1(n4345), .A2(n4346), .ZN(n4192) );
  AND2_X1 U4961 ( .A1(n4261), .A2(n4192), .ZN(n4211) );
  INV_X1 U4962 ( .A(n4211), .ZN(n4194) );
  OAI21_X1 U4963 ( .B1(n4195), .B2(n4194), .A(n4193), .ZN(n4268) );
  XNOR2_X1 U4964 ( .A(n4276), .B(n4375), .ZN(n4704) );
  INV_X1 U4965 ( .A(n4704), .ZN(n4366) );
  NAND2_X1 U4966 ( .A1(n4197), .A2(n4196), .ZN(n4433) );
  NAND2_X1 U4967 ( .A1(n4430), .A2(n4198), .ZN(n4448) );
  XNOR2_X1 U4968 ( .A(n4484), .B(n4512), .ZN(n4502) );
  NOR2_X1 U4969 ( .A1(n4469), .A2(n4502), .ZN(n4230) );
  NAND3_X1 U4970 ( .A1(n4551), .A2(n4200), .A3(n4199), .ZN(n4215) );
  XNOR2_X1 U4971 ( .A(n4545), .B(n4535), .ZN(n4532) );
  NOR2_X1 U4972 ( .A1(n4201), .A2(n4954), .ZN(n4207) );
  AND4_X1 U4973 ( .A1(n4204), .A2(n4390), .A3(n4402), .A4(n4412), .ZN(n4205)
         );
  NAND4_X1 U4974 ( .A1(n4207), .A2(n4600), .A3(n4206), .A4(n4205), .ZN(n4214)
         );
  NAND4_X1 U4975 ( .A1(n4212), .A2(n4211), .A3(n4210), .A4(n4656), .ZN(n4213)
         );
  NOR4_X1 U4976 ( .A1(n4215), .A2(n4532), .A3(n4214), .A4(n4213), .ZN(n4229)
         );
  NOR2_X1 U4977 ( .A1(n4216), .A2(n4242), .ZN(n4488) );
  NAND2_X1 U4978 ( .A1(n4218), .A2(n4217), .ZN(n4677) );
  OR4_X1 U4979 ( .A1(n4220), .A2(n4615), .A3(n4677), .A4(n4219), .ZN(n4227) );
  NAND4_X1 U4980 ( .A1(n4567), .A2(n4223), .A3(n4222), .A4(n4221), .ZN(n4226)
         );
  XNOR2_X1 U4981 ( .A(n4278), .B(n4224), .ZN(n4631) );
  NOR4_X1 U4982 ( .A1(n4227), .A2(n4226), .A3(n4631), .A4(n4225), .ZN(n4228)
         );
  OAI21_X1 U4983 ( .B1(n4233), .B2(n4232), .A(n4231), .ZN(n4238) );
  INV_X1 U4984 ( .A(n4234), .ZN(n4236) );
  AOI211_X1 U4985 ( .C1(n4238), .C2(n4237), .A(n4236), .B(n4235), .ZN(n4241)
         );
  OAI21_X1 U4986 ( .B1(n4241), .B2(n4240), .A(n4239), .ZN(n4243) );
  AOI21_X1 U4987 ( .B1(n4243), .B2(n2426), .A(n4242), .ZN(n4247) );
  INV_X1 U4988 ( .A(n4245), .ZN(n4246) );
  NOR3_X1 U4989 ( .A1(n4247), .A2(n2425), .A3(n4246), .ZN(n4253) );
  NOR2_X1 U4990 ( .A1(n4249), .A2(n4248), .ZN(n4250) );
  OAI211_X1 U4991 ( .C1(n4253), .C2(n4252), .A(n4251), .B(n4250), .ZN(n4260)
         );
  NAND3_X1 U4992 ( .A1(n4255), .A2(n4390), .A3(n4254), .ZN(n4256) );
  NAND2_X1 U4993 ( .A1(n4257), .A2(n4256), .ZN(n4259) );
  INV_X1 U4994 ( .A(n4345), .ZN(n4258) );
  AOI22_X1 U4995 ( .A1(n4260), .A2(n4259), .B1(n4258), .B2(n4350), .ZN(n4263)
         );
  AOI21_X1 U4996 ( .B1(n4261), .B2(n4345), .A(n4346), .ZN(n4262) );
  NOR2_X1 U4997 ( .A1(n4263), .A2(n4262), .ZN(n4265) );
  MUX2_X1 U4998 ( .A(n4266), .B(n4265), .S(n4264), .Z(n4267) );
  MUX2_X1 U4999 ( .A(n4268), .B(n4267), .S(n4880), .Z(n4269) );
  XNOR2_X1 U5000 ( .A(n4269), .B(n4881), .ZN(n4275) );
  NAND2_X1 U5001 ( .A1(n4271), .A2(n4270), .ZN(n4272) );
  OAI211_X1 U5002 ( .C1(n4879), .C2(n4274), .A(n4272), .B(B_REG_SCAN_IN), .ZN(
        n4273) );
  OAI21_X1 U5003 ( .B1(n4275), .B2(n4274), .A(n4273), .ZN(U3239) );
  MUX2_X1 U5004 ( .A(n4276), .B(DATAO_REG_29__SCAN_IN), .S(n4285), .Z(U3579)
         );
  MUX2_X1 U5005 ( .A(DATAO_REG_28__SCAN_IN), .B(n4392), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U5006 ( .A(n4391), .B(DATAO_REG_26__SCAN_IN), .S(n4285), .Z(U3576)
         );
  MUX2_X1 U5007 ( .A(n4399), .B(DATAO_REG_25__SCAN_IN), .S(n4285), .Z(U3575)
         );
  MUX2_X1 U5008 ( .A(n4415), .B(DATAO_REG_24__SCAN_IN), .S(n4285), .Z(U3574)
         );
  MUX2_X1 U5009 ( .A(n4452), .B(DATAO_REG_22__SCAN_IN), .S(n4285), .Z(U3572)
         );
  MUX2_X1 U5010 ( .A(n4505), .B(DATAO_REG_21__SCAN_IN), .S(n4285), .Z(U3571)
         );
  MUX2_X1 U5011 ( .A(n4564), .B(DATAO_REG_18__SCAN_IN), .S(n4285), .Z(U3568)
         );
  MUX2_X1 U5012 ( .A(DATAO_REG_16__SCAN_IN), .B(n4277), .S(U4043), .Z(U3566)
         );
  MUX2_X1 U5013 ( .A(n4608), .B(DATAO_REG_14__SCAN_IN), .S(n4285), .Z(U3564)
         );
  MUX2_X1 U5014 ( .A(n4278), .B(DATAO_REG_13__SCAN_IN), .S(n4285), .Z(U3563)
         );
  MUX2_X1 U5015 ( .A(n4279), .B(DATAO_REG_11__SCAN_IN), .S(n4285), .Z(U3561)
         );
  MUX2_X1 U5016 ( .A(n4280), .B(DATAO_REG_9__SCAN_IN), .S(n4285), .Z(U3559) );
  MUX2_X1 U5017 ( .A(n4681), .B(DATAO_REG_8__SCAN_IN), .S(n4285), .Z(U3558) );
  MUX2_X1 U5018 ( .A(n4281), .B(DATAO_REG_7__SCAN_IN), .S(n4285), .Z(U3557) );
  MUX2_X1 U5019 ( .A(n4282), .B(DATAO_REG_6__SCAN_IN), .S(n4285), .Z(U3556) );
  MUX2_X1 U5020 ( .A(n4283), .B(DATAO_REG_5__SCAN_IN), .S(n4285), .Z(U3555) );
  MUX2_X1 U5021 ( .A(n4284), .B(DATAO_REG_3__SCAN_IN), .S(n4285), .Z(U3553) );
  MUX2_X1 U5022 ( .A(n3322), .B(DATAO_REG_1__SCAN_IN), .S(n4285), .Z(U3551) );
  MUX2_X1 U5023 ( .A(n3313), .B(DATAO_REG_0__SCAN_IN), .S(n4285), .Z(U3550) );
  NAND2_X1 U5024 ( .A1(n4286), .A2(n4289), .ZN(n4288) );
  OAI211_X1 U5025 ( .C1(n4290), .C2(n4289), .A(n4288), .B(n4287), .ZN(n4291)
         );
  OAI211_X1 U5026 ( .C1(n2222), .C2(n4292), .A(n4291), .B(U4043), .ZN(n4901)
         );
  AOI22_X1 U5027 ( .A1(ADDR_REG_2__SCAN_IN), .A2(n4942), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n4302) );
  XOR2_X1 U5028 ( .A(n4293), .B(n4294), .Z(n4295) );
  AOI22_X1 U5029 ( .A1(n4296), .A2(n2521), .B1(n4948), .B2(n4295), .ZN(n4301)
         );
  OAI211_X1 U5030 ( .C1(n4299), .C2(n4298), .A(n4935), .B(n4297), .ZN(n4300)
         );
  NAND4_X1 U5031 ( .A1(n4901), .A2(n4302), .A3(n4301), .A4(n4300), .ZN(U3242)
         );
  OAI211_X1 U5032 ( .C1(n4305), .C2(n4304), .A(n4303), .B(n4935), .ZN(n4314)
         );
  NOR2_X1 U5033 ( .A1(n4949), .A2(n4306), .ZN(n4307) );
  AOI211_X1 U5034 ( .C1(n4942), .C2(ADDR_REG_9__SCAN_IN), .A(n4308), .B(n4307), 
        .ZN(n4313) );
  OAI211_X1 U5035 ( .C1(n4311), .C2(n4310), .A(n4309), .B(n4948), .ZN(n4312)
         );
  NAND3_X1 U5036 ( .A1(n4314), .A2(n4313), .A3(n4312), .ZN(U3249) );
  AOI22_X1 U5037 ( .A1(REG1_REG_18__SCAN_IN), .A2(n4980), .B1(n4334), .B2(
        n4315), .ZN(n4939) );
  AOI22_X1 U5038 ( .A1(n4333), .A2(REG1_REG_17__SCAN_IN), .B1(n4761), .B2(
        n4981), .ZN(n4929) );
  INV_X1 U5039 ( .A(n4330), .ZN(n4985) );
  AOI22_X1 U5040 ( .A1(REG1_REG_15__SCAN_IN), .A2(n4985), .B1(n4330), .B2(
        n4319), .ZN(n4904) );
  NAND2_X1 U5041 ( .A1(n4320), .A2(n4983), .ZN(n4321) );
  XNOR2_X1 U5042 ( .A(n4881), .B(REG1_REG_19__SCAN_IN), .ZN(n4322) );
  NAND2_X1 U5043 ( .A1(REG2_REG_18__SCAN_IN), .A2(n4334), .ZN(n4323) );
  OAI21_X1 U5044 ( .B1(REG2_REG_18__SCAN_IN), .B2(n4334), .A(n4323), .ZN(n4947) );
  NOR2_X1 U5045 ( .A1(n4333), .A2(REG2_REG_17__SCAN_IN), .ZN(n4324) );
  AOI21_X1 U5046 ( .B1(REG2_REG_17__SCAN_IN), .B2(n4333), .A(n4324), .ZN(n4932) );
  INV_X1 U5047 ( .A(n4325), .ZN(n4328) );
  INV_X1 U5048 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4329) );
  AOI22_X1 U5049 ( .A1(REG2_REG_15__SCAN_IN), .A2(n4985), .B1(n4330), .B2(
        n4329), .ZN(n4910) );
  NAND2_X1 U5050 ( .A1(n4331), .A2(n4983), .ZN(n4332) );
  INV_X1 U5051 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4335) );
  MUX2_X1 U5052 ( .A(REG2_REG_19__SCAN_IN), .B(n4335), .S(n4881), .Z(n4336) );
  NAND2_X1 U5053 ( .A1(n4942), .A2(ADDR_REG_19__SCAN_IN), .ZN(n4337) );
  OAI211_X1 U5054 ( .C1(n4949), .C2(n4339), .A(n4338), .B(n4337), .ZN(n4340)
         );
  AND2_X1 U5055 ( .A1(n4706), .A2(n4341), .ZN(n4342) );
  XNOR2_X1 U5056 ( .A(n4349), .B(n4346), .ZN(n4809) );
  AND2_X1 U5057 ( .A1(n4343), .A2(B_REG_SCAN_IN), .ZN(n4344) );
  NOR2_X1 U5058 ( .A1(n4678), .A2(n4344), .ZN(n4361) );
  NAND2_X1 U5059 ( .A1(n4345), .A2(n4361), .ZN(n4352) );
  OAI21_X1 U5060 ( .B1(n4346), .B2(n4795), .A(n4352), .ZN(n4806) );
  NAND2_X1 U5061 ( .A1(n4957), .A2(n4806), .ZN(n4348) );
  NAND2_X1 U5062 ( .A1(n2142), .A2(REG2_REG_31__SCAN_IN), .ZN(n4347) );
  OAI211_X1 U5063 ( .C1(n4809), .C2(n4572), .A(n4348), .B(n4347), .ZN(U3260)
         );
  AOI21_X1 U5064 ( .B1(n4350), .B2(n4374), .A(n4349), .ZN(n4810) );
  NAND2_X1 U5065 ( .A1(n4810), .A2(n4693), .ZN(n4354) );
  NAND2_X1 U5066 ( .A1(n4768), .A2(n4350), .ZN(n4351) );
  NAND2_X1 U5067 ( .A1(n4352), .A2(n4351), .ZN(n4811) );
  NAND2_X1 U5068 ( .A1(n4957), .A2(n4811), .ZN(n4353) );
  OAI211_X1 U5069 ( .C1(n4957), .C2(n4355), .A(n4354), .B(n4353), .ZN(U3261)
         );
  NOR2_X1 U5070 ( .A1(n4369), .A2(n4358), .ZN(n4705) );
  INV_X1 U5071 ( .A(n4705), .ZN(n4707) );
  NAND2_X1 U5072 ( .A1(n4713), .A2(n4707), .ZN(n4359) );
  XNOR2_X1 U5073 ( .A(n4359), .B(n4366), .ZN(n4380) );
  INV_X1 U5074 ( .A(n4360), .ZN(n4371) );
  INV_X1 U5075 ( .A(n4361), .ZN(n4370) );
  INV_X1 U5076 ( .A(n4362), .ZN(n4363) );
  AOI21_X1 U5077 ( .B1(n4365), .B2(n4364), .A(n4363), .ZN(n4367) );
  XNOR2_X1 U5078 ( .A(n4367), .B(n4366), .ZN(n4368) );
  NAND2_X1 U5079 ( .A1(n4372), .A2(n4375), .ZN(n4373) );
  NAND2_X1 U5080 ( .A1(n4374), .A2(n4373), .ZN(n4709) );
  AOI22_X1 U5081 ( .A1(n4619), .A2(n4375), .B1(n2142), .B2(
        REG2_REG_29__SCAN_IN), .ZN(n4376) );
  OAI21_X1 U5082 ( .B1(n4709), .B2(n4572), .A(n4376), .ZN(n4377) );
  AOI21_X1 U5083 ( .B1(n4378), .B2(n4957), .A(n4377), .ZN(n4379) );
  OAI21_X1 U5084 ( .B1(n4380), .B2(n4697), .A(n4379), .ZN(U3354) );
  XNOR2_X1 U5085 ( .A(n4381), .B(n4390), .ZN(n4718) );
  INV_X1 U5086 ( .A(n4382), .ZN(n4404) );
  AOI21_X1 U5087 ( .B1(n4714), .B2(n4404), .A(n4383), .ZN(n4715) );
  NOR2_X1 U5088 ( .A1(n4666), .A2(n4384), .ZN(n4388) );
  INV_X1 U5089 ( .A(REG2_REG_27__SCAN_IN), .ZN(n4385) );
  OAI22_X1 U5090 ( .A1(n4386), .A2(n4643), .B1(n4385), .B2(n4957), .ZN(n4387)
         );
  AOI211_X1 U5091 ( .C1(n4715), .C2(n4693), .A(n4388), .B(n4387), .ZN(n4395)
         );
  OAI21_X1 U5092 ( .B1(n2413), .B2(n4390), .A(n4389), .ZN(n4393) );
  AOI222_X1 U5093 ( .A1(n4525), .A2(n4393), .B1(n4392), .B2(n4563), .C1(n4391), 
        .C2(n4682), .ZN(n4717) );
  OR2_X1 U5094 ( .A1(n4717), .A2(n2142), .ZN(n4394) );
  OAI211_X1 U5095 ( .C1(n4718), .C2(n4697), .A(n4395), .B(n4394), .ZN(U3263)
         );
  XNOR2_X1 U5096 ( .A(n4398), .B(n4402), .ZN(n4401) );
  AOI222_X1 U5097 ( .A1(n4525), .A2(n4401), .B1(n4400), .B2(n4563), .C1(n4399), 
        .C2(n4682), .ZN(n4719) );
  XNOR2_X1 U5098 ( .A(n4403), .B(n4402), .ZN(n4721) );
  NAND2_X1 U5099 ( .A1(n4721), .A2(n4577), .ZN(n4409) );
  OAI22_X1 U5100 ( .A1(n4666), .A2(n4720), .B1(n2995), .B2(n4957), .ZN(n4406)
         );
  OAI21_X1 U5101 ( .B1(n4419), .B2(n4720), .A(n4404), .ZN(n4820) );
  NOR2_X1 U5102 ( .A1(n4820), .A2(n4572), .ZN(n4405) );
  AOI211_X1 U5103 ( .C1(n4953), .C2(n4407), .A(n4406), .B(n4405), .ZN(n4408)
         );
  OAI211_X1 U5104 ( .C1(n4719), .C2(n2142), .A(n4409), .B(n4408), .ZN(U3264)
         );
  XOR2_X1 U5105 ( .A(n4412), .B(n4410), .Z(n4724) );
  INV_X1 U5106 ( .A(n4724), .ZN(n4428) );
  XOR2_X1 U5107 ( .A(n4412), .B(n4411), .Z(n4413) );
  NAND2_X1 U5108 ( .A1(n4413), .A2(n4525), .ZN(n4417) );
  AOI22_X1 U5109 ( .A1(n4415), .A2(n4682), .B1(n4414), .B2(n4768), .ZN(n4416)
         );
  OAI211_X1 U5110 ( .C1(n4418), .C2(n4678), .A(n4417), .B(n4416), .ZN(n4723)
         );
  INV_X1 U5111 ( .A(n4439), .ZN(n4422) );
  INV_X1 U5112 ( .A(n4419), .ZN(n4420) );
  OAI21_X1 U5113 ( .B1(n4422), .B2(n4421), .A(n4420), .ZN(n4824) );
  INV_X1 U5114 ( .A(n4423), .ZN(n4424) );
  AOI22_X1 U5115 ( .A1(n4424), .A2(n4953), .B1(REG2_REG_25__SCAN_IN), .B2(
        n2142), .ZN(n4425) );
  OAI21_X1 U5116 ( .B1(n4824), .B2(n4572), .A(n4425), .ZN(n4426) );
  AOI21_X1 U5117 ( .B1(n4723), .B2(n4957), .A(n4426), .ZN(n4427) );
  OAI21_X1 U5118 ( .B1(n4428), .B2(n4697), .A(n4427), .ZN(U3265) );
  XNOR2_X1 U5119 ( .A(n4429), .B(n4433), .ZN(n4728) );
  INV_X1 U5120 ( .A(n4728), .ZN(n4446) );
  NAND2_X1 U5121 ( .A1(n4431), .A2(n4430), .ZN(n4432) );
  XOR2_X1 U5122 ( .A(n4433), .B(n4432), .Z(n4434) );
  NAND2_X1 U5123 ( .A1(n4434), .A2(n4525), .ZN(n4437) );
  AOI22_X1 U5124 ( .A1(n4473), .A2(n4682), .B1(n4435), .B2(n4768), .ZN(n4436)
         );
  OAI211_X1 U5125 ( .C1(n4438), .C2(n4678), .A(n4437), .B(n4436), .ZN(n4727)
         );
  INV_X1 U5126 ( .A(n4456), .ZN(n4441) );
  OAI21_X1 U5127 ( .B1(n4441), .B2(n4440), .A(n4439), .ZN(n4828) );
  AOI22_X1 U5128 ( .A1(n4442), .A2(n4953), .B1(REG2_REG_24__SCAN_IN), .B2(
        n2142), .ZN(n4443) );
  OAI21_X1 U5129 ( .B1(n4828), .B2(n4572), .A(n4443), .ZN(n4444) );
  AOI21_X1 U5130 ( .B1(n4727), .B2(n4957), .A(n4444), .ZN(n4445) );
  OAI21_X1 U5131 ( .B1(n4446), .B2(n4697), .A(n4445), .ZN(U3266) );
  XOR2_X1 U5132 ( .A(n4448), .B(n4447), .Z(n4732) );
  INV_X1 U5133 ( .A(n4732), .ZN(n4462) );
  NOR2_X1 U5134 ( .A1(n4468), .A2(n4469), .ZN(n4467) );
  NOR2_X1 U5135 ( .A1(n4467), .A2(n2425), .ZN(n4449) );
  XNOR2_X1 U5136 ( .A(n4449), .B(n4448), .ZN(n4450) );
  NAND2_X1 U5137 ( .A1(n4450), .A2(n4525), .ZN(n4454) );
  AOI22_X1 U5138 ( .A1(n4452), .A2(n4682), .B1(n4768), .B2(n4451), .ZN(n4453)
         );
  OAI211_X1 U5139 ( .C1(n4455), .C2(n4678), .A(n4454), .B(n4453), .ZN(n4731)
         );
  OAI21_X1 U5140 ( .B1(n4475), .B2(n4457), .A(n4456), .ZN(n4832) );
  AOI22_X1 U5141 ( .A1(n4458), .A2(n4953), .B1(REG2_REG_23__SCAN_IN), .B2(
        n2142), .ZN(n4459) );
  OAI21_X1 U5142 ( .B1(n4832), .B2(n4572), .A(n4459), .ZN(n4460) );
  AOI21_X1 U5143 ( .B1(n4731), .B2(n4957), .A(n4460), .ZN(n4461) );
  OAI21_X1 U5144 ( .B1(n4462), .B2(n4697), .A(n4461), .ZN(U3267) );
  OAI21_X1 U5145 ( .B1(n4464), .B2(n4469), .A(n4463), .ZN(n4739) );
  OAI22_X1 U5146 ( .A1(n4466), .A2(n4659), .B1(n4465), .B2(n4795), .ZN(n4472)
         );
  AOI21_X1 U5147 ( .B1(n4469), .B2(n4468), .A(n4467), .ZN(n4470) );
  NOR2_X1 U5148 ( .A1(n4470), .A2(n4684), .ZN(n4471) );
  AOI211_X1 U5149 ( .C1(n4563), .C2(n4473), .A(n4472), .B(n4471), .ZN(n4738)
         );
  AOI22_X1 U5150 ( .A1(n4474), .A2(n4953), .B1(n2142), .B2(
        REG2_REG_22__SCAN_IN), .ZN(n4478) );
  INV_X1 U5151 ( .A(n4475), .ZN(n4736) );
  NAND2_X1 U5152 ( .A1(n4491), .A2(n4476), .ZN(n4735) );
  NAND3_X1 U5153 ( .A1(n4736), .A2(n4693), .A3(n4735), .ZN(n4477) );
  OAI211_X1 U5154 ( .C1(n4738), .C2(n2142), .A(n4478), .B(n4477), .ZN(n4479)
         );
  INV_X1 U5155 ( .A(n4479), .ZN(n4480) );
  OAI21_X1 U5156 ( .B1(n4697), .B2(n4739), .A(n4480), .ZN(U3268) );
  XNOR2_X1 U5157 ( .A(n4481), .B(n4488), .ZN(n4482) );
  NAND2_X1 U5158 ( .A1(n4482), .A2(n4525), .ZN(n4486) );
  AOI22_X1 U5159 ( .A1(n4484), .A2(n4682), .B1(n4483), .B2(n4768), .ZN(n4485)
         );
  OAI211_X1 U5160 ( .C1(n4487), .C2(n4678), .A(n4486), .B(n4485), .ZN(n4740)
         );
  INV_X1 U5161 ( .A(n4740), .ZN(n4498) );
  XNOR2_X1 U5162 ( .A(n4489), .B(n4488), .ZN(n4741) );
  NAND2_X1 U5163 ( .A1(n4741), .A2(n4577), .ZN(n4497) );
  NOR2_X1 U5164 ( .A1(n4490), .A2(n4643), .ZN(n4495) );
  INV_X1 U5165 ( .A(n4511), .ZN(n4493) );
  OAI21_X1 U5166 ( .B1(n4493), .B2(n4492), .A(n4491), .ZN(n4837) );
  NOR2_X1 U5167 ( .A1(n4837), .A2(n4572), .ZN(n4494) );
  AOI211_X1 U5168 ( .C1(n2142), .C2(REG2_REG_21__SCAN_IN), .A(n4495), .B(n4494), .ZN(n4496) );
  OAI211_X1 U5169 ( .C1(n2142), .C2(n4498), .A(n4497), .B(n4496), .ZN(U3269)
         );
  INV_X1 U5170 ( .A(n4499), .ZN(n4500) );
  NAND2_X1 U5171 ( .A1(n4501), .A2(n4500), .ZN(n4503) );
  INV_X1 U5172 ( .A(n4502), .ZN(n4508) );
  XNOR2_X1 U5173 ( .A(n4503), .B(n4508), .ZN(n4504) );
  NAND2_X1 U5174 ( .A1(n4504), .A2(n4525), .ZN(n4507) );
  AOI22_X1 U5175 ( .A1(n4505), .A2(n4563), .B1(n4682), .B2(n4545), .ZN(n4506)
         );
  NAND2_X1 U5176 ( .A1(n4507), .A2(n4506), .ZN(n4747) );
  INV_X1 U5177 ( .A(n4747), .ZN(n4517) );
  XNOR2_X1 U5178 ( .A(n4509), .B(n4508), .ZN(n4744) );
  NAND2_X1 U5179 ( .A1(n4744), .A2(n4577), .ZN(n4516) );
  OAI22_X1 U5180 ( .A1(n4957), .A2(n3108), .B1(n4510), .B2(n4643), .ZN(n4514)
         );
  OAI21_X1 U5181 ( .B1(n4533), .B2(n4512), .A(n4511), .ZN(n4841) );
  NOR2_X1 U5182 ( .A1(n4841), .A2(n4572), .ZN(n4513) );
  AOI211_X1 U5183 ( .C1(n4619), .C2(n4745), .A(n4514), .B(n4513), .ZN(n4515)
         );
  OAI211_X1 U5184 ( .C1(n2142), .C2(n4517), .A(n4516), .B(n4515), .ZN(U3270)
         );
  INV_X1 U5185 ( .A(n4518), .ZN(n4520) );
  OAI21_X1 U5186 ( .B1(n4560), .B2(n4520), .A(n4519), .ZN(n4541) );
  INV_X1 U5187 ( .A(n4521), .ZN(n4523) );
  OAI21_X1 U5188 ( .B1(n4541), .B2(n4523), .A(n4522), .ZN(n4524) );
  XNOR2_X1 U5189 ( .A(n4524), .B(n4532), .ZN(n4526) );
  NAND2_X1 U5190 ( .A1(n4526), .A2(n4525), .ZN(n4529) );
  AOI22_X1 U5191 ( .A1(n4564), .A2(n4682), .B1(n4768), .B2(n4527), .ZN(n4528)
         );
  OAI211_X1 U5192 ( .C1(n4530), .C2(n4678), .A(n4529), .B(n4528), .ZN(n4752)
         );
  INV_X1 U5193 ( .A(n4752), .ZN(n4540) );
  XNOR2_X1 U5194 ( .A(n4531), .B(n4532), .ZN(n4753) );
  INV_X1 U5195 ( .A(n4533), .ZN(n4534) );
  OAI21_X1 U5196 ( .B1(n2183), .B2(n4535), .A(n4534), .ZN(n4845) );
  NOR2_X1 U5197 ( .A1(n4845), .A2(n4572), .ZN(n4538) );
  OAI22_X1 U5198 ( .A1(n4957), .A2(n4335), .B1(n4536), .B2(n4643), .ZN(n4537)
         );
  AOI211_X1 U5199 ( .C1(n4753), .C2(n4577), .A(n4538), .B(n4537), .ZN(n4539)
         );
  OAI21_X1 U5200 ( .B1(n4540), .B2(n2142), .A(n4539), .ZN(U3271) );
  OAI22_X1 U5201 ( .A1(n4584), .A2(n4659), .B1(n4552), .B2(n4795), .ZN(n4544)
         );
  XOR2_X1 U5202 ( .A(n4551), .B(n4541), .Z(n4542) );
  NOR2_X1 U5203 ( .A1(n4542), .A2(n4684), .ZN(n4543) );
  AOI211_X1 U5204 ( .C1(n4563), .C2(n4545), .A(n4544), .B(n4543), .ZN(n4757)
         );
  NAND2_X1 U5205 ( .A1(n4547), .A2(n4546), .ZN(n4550) );
  INV_X1 U5206 ( .A(n4548), .ZN(n4549) );
  AOI21_X1 U5207 ( .B1(n4551), .B2(n4550), .A(n4549), .ZN(n4758) );
  INV_X1 U5208 ( .A(n4758), .ZN(n4558) );
  XNOR2_X1 U5209 ( .A(n4571), .B(n4552), .ZN(n4553) );
  NAND2_X1 U5210 ( .A1(n4553), .A2(n4994), .ZN(n4756) );
  NOR2_X1 U5211 ( .A1(n4756), .A2(n4554), .ZN(n4557) );
  OAI22_X1 U5212 ( .A1(n4957), .A2(n2974), .B1(n4555), .B2(n4643), .ZN(n4556)
         );
  AOI211_X1 U5213 ( .C1(n4558), .C2(n4577), .A(n4557), .B(n4556), .ZN(n4559)
         );
  OAI21_X1 U5214 ( .B1(n4757), .B2(n2142), .A(n4559), .ZN(U3272) );
  XNOR2_X1 U5215 ( .A(n4560), .B(n4567), .ZN(n4566) );
  OAI22_X1 U5216 ( .A1(n4609), .A2(n4659), .B1(n4795), .B2(n4561), .ZN(n4562)
         );
  AOI21_X1 U5217 ( .B1(n4564), .B2(n4563), .A(n4562), .ZN(n4565) );
  OAI21_X1 U5218 ( .B1(n4566), .B2(n4684), .A(n4565), .ZN(n4759) );
  INV_X1 U5219 ( .A(n4759), .ZN(n4579) );
  XNOR2_X1 U5220 ( .A(n4568), .B(n4567), .ZN(n4760) );
  NAND2_X1 U5221 ( .A1(n4589), .A2(n4569), .ZN(n4570) );
  NAND2_X1 U5222 ( .A1(n4571), .A2(n4570), .ZN(n4850) );
  NOR2_X1 U5223 ( .A1(n4850), .A2(n4572), .ZN(n4576) );
  INV_X1 U5224 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4574) );
  OAI22_X1 U5225 ( .A1(n4957), .A2(n4574), .B1(n4573), .B2(n4643), .ZN(n4575)
         );
  AOI211_X1 U5226 ( .C1(n4760), .C2(n4577), .A(n4576), .B(n4575), .ZN(n4578)
         );
  OAI21_X1 U5227 ( .B1(n4579), .B2(n2142), .A(n4578), .ZN(U3273) );
  INV_X1 U5228 ( .A(n4580), .ZN(n4582) );
  AOI21_X1 U5229 ( .B1(n4582), .B2(n4581), .A(n4684), .ZN(n4587) );
  OAI22_X1 U5230 ( .A1(n4584), .A2(n4678), .B1(n4583), .B2(n4659), .ZN(n4585)
         );
  AOI21_X1 U5231 ( .B1(n4587), .B2(n4586), .A(n4585), .ZN(n4766) );
  INV_X1 U5232 ( .A(n4588), .ZN(n4591) );
  INV_X1 U5233 ( .A(n4589), .ZN(n4590) );
  AOI21_X1 U5234 ( .B1(n4763), .B2(n4591), .A(n4590), .ZN(n4764) );
  AOI22_X1 U5235 ( .A1(n2142), .A2(REG2_REG_16__SCAN_IN), .B1(n4592), .B2(
        n4953), .ZN(n4593) );
  OAI21_X1 U5236 ( .B1(n4666), .B2(n4594), .A(n4593), .ZN(n4605) );
  OR2_X1 U5237 ( .A1(n4596), .A2(n4595), .ZN(n4599) );
  NAND2_X1 U5238 ( .A1(n4599), .A2(n4597), .ZN(n4603) );
  NAND2_X1 U5239 ( .A1(n4599), .A2(n4598), .ZN(n4601) );
  NAND2_X1 U5240 ( .A1(n4601), .A2(n4600), .ZN(n4602) );
  NAND2_X1 U5241 ( .A1(n4603), .A2(n4602), .ZN(n4767) );
  NOR2_X1 U5242 ( .A1(n4767), .A2(n4697), .ZN(n4604) );
  AOI211_X1 U5243 ( .C1(n4764), .C2(n4693), .A(n4605), .B(n4604), .ZN(n4606)
         );
  OAI21_X1 U5244 ( .B1(n2142), .B2(n4766), .A(n4606), .ZN(U3274) );
  AOI21_X1 U5245 ( .B1(n4607), .B2(n4615), .A(n4684), .ZN(n4612) );
  INV_X1 U5246 ( .A(n4608), .ZN(n4634) );
  OAI22_X1 U5247 ( .A1(n4609), .A2(n4678), .B1(n4634), .B2(n4659), .ZN(n4610)
         );
  AOI21_X1 U5248 ( .B1(n4612), .B2(n4611), .A(n4610), .ZN(n4772) );
  NAND2_X1 U5249 ( .A1(n4614), .A2(n4613), .ZN(n4616) );
  XNOR2_X1 U5250 ( .A(n4616), .B(n2399), .ZN(n4773) );
  OAI22_X1 U5251 ( .A1(n4957), .A2(n4329), .B1(n4617), .B2(n4643), .ZN(n4618)
         );
  AOI21_X1 U5252 ( .B1(n4769), .B2(n4619), .A(n4618), .ZN(n4622) );
  XNOR2_X1 U5253 ( .A(n4620), .B(n4769), .ZN(n4770) );
  NAND2_X1 U5254 ( .A1(n4770), .A2(n4693), .ZN(n4621) );
  OAI211_X1 U5255 ( .C1(n4773), .C2(n4697), .A(n4622), .B(n4621), .ZN(n4623)
         );
  INV_X1 U5256 ( .A(n4623), .ZN(n4624) );
  OAI21_X1 U5257 ( .B1(n4772), .B2(n2142), .A(n4624), .ZN(U3275) );
  XNOR2_X1 U5258 ( .A(n4626), .B(n4631), .ZN(n4781) );
  INV_X1 U5259 ( .A(n4781), .ZN(n4650) );
  OAI21_X1 U5260 ( .B1(n4629), .B2(n4628), .A(n4627), .ZN(n4630) );
  XOR2_X1 U5261 ( .A(n4631), .B(n4630), .Z(n4638) );
  AOI22_X1 U5262 ( .A1(n4632), .A2(n4682), .B1(n4639), .B2(n4768), .ZN(n4633)
         );
  OAI21_X1 U5263 ( .B1(n4634), .B2(n4678), .A(n4633), .ZN(n4635) );
  AOI21_X1 U5264 ( .B1(n4781), .B2(n4636), .A(n4635), .ZN(n4637) );
  OAI21_X1 U5265 ( .B1(n4638), .B2(n4684), .A(n4637), .ZN(n4780) );
  NAND2_X1 U5266 ( .A1(n4780), .A2(n4957), .ZN(n4648) );
  NAND2_X1 U5267 ( .A1(n4640), .A2(n4639), .ZN(n4641) );
  NAND2_X1 U5268 ( .A1(n4642), .A2(n4641), .ZN(n4860) );
  INV_X1 U5269 ( .A(n4860), .ZN(n4646) );
  OAI22_X1 U5270 ( .A1(n4957), .A2(n3683), .B1(n4644), .B2(n4643), .ZN(n4645)
         );
  AOI21_X1 U5271 ( .B1(n4646), .B2(n4693), .A(n4645), .ZN(n4647) );
  OAI211_X1 U5272 ( .C1(n4650), .C2(n4649), .A(n4648), .B(n4647), .ZN(U3277)
         );
  XNOR2_X1 U5273 ( .A(n4651), .B(n4656), .ZN(n4796) );
  NAND2_X1 U5274 ( .A1(n4673), .A2(n4652), .ZN(n4654) );
  AND2_X1 U5275 ( .A1(n4654), .A2(n4653), .ZN(n4655) );
  XOR2_X1 U5276 ( .A(n4656), .B(n4655), .Z(n4657) );
  OAI222_X1 U5277 ( .A1(n4678), .A2(n4660), .B1(n4659), .B2(n4658), .C1(n4657), 
        .C2(n4684), .ZN(n4798) );
  NAND2_X1 U5278 ( .A1(n4798), .A2(n4957), .ZN(n4670) );
  INV_X1 U5279 ( .A(n4691), .ZN(n4663) );
  INV_X1 U5280 ( .A(n4661), .ZN(n4662) );
  OAI21_X1 U5281 ( .B1(n4663), .B2(n4794), .A(n4662), .ZN(n4873) );
  INV_X1 U5282 ( .A(n4873), .ZN(n4668) );
  AOI22_X1 U5283 ( .A1(n2142), .A2(REG2_REG_10__SCAN_IN), .B1(n4664), .B2(
        n4953), .ZN(n4665) );
  OAI21_X1 U5284 ( .B1(n4666), .B2(n4794), .A(n4665), .ZN(n4667) );
  AOI21_X1 U5285 ( .B1(n4668), .B2(n4693), .A(n4667), .ZN(n4669) );
  OAI211_X1 U5286 ( .C1(n4697), .C2(n4796), .A(n4670), .B(n4669), .ZN(U3280)
         );
  XOR2_X1 U5287 ( .A(n4671), .B(n4677), .Z(n4803) );
  INV_X1 U5288 ( .A(n4803), .ZN(n4696) );
  NAND2_X1 U5289 ( .A1(n4673), .A2(n4672), .ZN(n4675) );
  NAND2_X1 U5290 ( .A1(n4675), .A2(n4674), .ZN(n4676) );
  XOR2_X1 U5291 ( .A(n4677), .B(n4676), .Z(n4685) );
  OAI22_X1 U5292 ( .A1(n4679), .A2(n4678), .B1(n4795), .B2(n2309), .ZN(n4680)
         );
  AOI21_X1 U5293 ( .B1(n4682), .B2(n4681), .A(n4680), .ZN(n4683) );
  OAI21_X1 U5294 ( .B1(n4685), .B2(n4684), .A(n4683), .ZN(n4802) );
  INV_X1 U5295 ( .A(n4802), .ZN(n4686) );
  MUX2_X1 U5296 ( .A(n4687), .B(n4686), .S(n4957), .Z(n4695) );
  NAND2_X1 U5297 ( .A1(n4689), .A2(n4688), .ZN(n4690) );
  AND2_X1 U5298 ( .A1(n4691), .A2(n4690), .ZN(n4875) );
  AOI22_X1 U5299 ( .A1(n4875), .A2(n4693), .B1(n4692), .B2(n4953), .ZN(n4694)
         );
  OAI211_X1 U5300 ( .C1(n4697), .C2(n4696), .A(n4695), .B(n4694), .ZN(U3281)
         );
  NOR2_X1 U5301 ( .A1(n5019), .A2(n4698), .ZN(n4699) );
  AOI21_X1 U5302 ( .B1(n5019), .B2(n4806), .A(n4699), .ZN(n4700) );
  OAI21_X1 U5303 ( .B1(n4809), .B2(n4801), .A(n4700), .ZN(U3549) );
  NAND2_X1 U5304 ( .A1(n4810), .A2(n4804), .ZN(n4702) );
  NAND2_X1 U5305 ( .A1(n5019), .A2(n4811), .ZN(n4701) );
  OAI211_X1 U5306 ( .C1(n5019), .C2(n4703), .A(n4702), .B(n4701), .ZN(U3548)
         );
  NAND2_X1 U5307 ( .A1(n4704), .A2(n5007), .ZN(n4712) );
  OAI22_X1 U5308 ( .A1(n4712), .A2(n4707), .B1(n4795), .B2(n4706), .ZN(n4708)
         );
  INV_X1 U5309 ( .A(n4708), .ZN(n4710) );
  MUX2_X1 U5310 ( .A(REG1_REG_29__SCAN_IN), .B(n4815), .S(n5019), .Z(U3547) );
  AOI22_X1 U5311 ( .A1(n4715), .A2(n4994), .B1(n4714), .B2(n4768), .ZN(n4716)
         );
  MUX2_X1 U5312 ( .A(REG1_REG_27__SCAN_IN), .B(n4816), .S(n5019), .Z(U3545) );
  AOI21_X1 U5313 ( .B1(n4724), .B2(n5007), .A(n4723), .ZN(n4821) );
  MUX2_X1 U5314 ( .A(n4725), .B(n4821), .S(n5019), .Z(n4726) );
  OAI21_X1 U5315 ( .B1(n4801), .B2(n4824), .A(n4726), .ZN(U3543) );
  AOI21_X1 U5316 ( .B1(n4728), .B2(n5007), .A(n4727), .ZN(n4825) );
  MUX2_X1 U5317 ( .A(n4729), .B(n4825), .S(n5019), .Z(n4730) );
  OAI21_X1 U5318 ( .B1(n4801), .B2(n4828), .A(n4730), .ZN(U3542) );
  AOI21_X1 U5319 ( .B1(n4732), .B2(n5007), .A(n4731), .ZN(n4829) );
  MUX2_X1 U5320 ( .A(n4733), .B(n4829), .S(n5019), .Z(n4734) );
  OAI21_X1 U5321 ( .B1(n4801), .B2(n4832), .A(n4734), .ZN(U3541) );
  NAND3_X1 U5322 ( .A1(n4736), .A2(n4994), .A3(n4735), .ZN(n4737) );
  OAI211_X1 U5323 ( .C1(n5002), .C2(n4739), .A(n4738), .B(n4737), .ZN(n4833)
         );
  MUX2_X1 U5324 ( .A(REG1_REG_22__SCAN_IN), .B(n4833), .S(n5019), .Z(U3540) );
  AOI21_X1 U5325 ( .B1(n4741), .B2(n5007), .A(n4740), .ZN(n4834) );
  MUX2_X1 U5326 ( .A(n4742), .B(n4834), .S(n5019), .Z(n4743) );
  OAI21_X1 U5327 ( .B1(n4801), .B2(n4837), .A(n4743), .ZN(U3539) );
  NAND2_X1 U5328 ( .A1(n4744), .A2(n5007), .ZN(n4749) );
  AND2_X1 U5329 ( .A1(n4768), .A2(n4745), .ZN(n4746) );
  NOR2_X1 U5330 ( .A1(n4747), .A2(n4746), .ZN(n4748) );
  AND2_X1 U5331 ( .A1(n4749), .A2(n4748), .ZN(n4838) );
  MUX2_X1 U5332 ( .A(n4750), .B(n4838), .S(n5019), .Z(n4751) );
  OAI21_X1 U5333 ( .B1(n4801), .B2(n4841), .A(n4751), .ZN(U3538) );
  AOI21_X1 U5334 ( .B1(n5007), .B2(n4753), .A(n4752), .ZN(n4842) );
  MUX2_X1 U5335 ( .A(n4754), .B(n4842), .S(n5019), .Z(n4755) );
  OAI21_X1 U5336 ( .B1(n4801), .B2(n4845), .A(n4755), .ZN(U3537) );
  OAI211_X1 U5337 ( .C1(n5002), .C2(n4758), .A(n4757), .B(n4756), .ZN(n4846)
         );
  MUX2_X1 U5338 ( .A(REG1_REG_18__SCAN_IN), .B(n4846), .S(n5019), .Z(U3536) );
  AOI21_X1 U5339 ( .B1(n4760), .B2(n5007), .A(n4759), .ZN(n4847) );
  MUX2_X1 U5340 ( .A(n4761), .B(n4847), .S(n5019), .Z(n4762) );
  OAI21_X1 U5341 ( .B1(n4801), .B2(n4850), .A(n4762), .ZN(U3535) );
  AOI22_X1 U5342 ( .A1(n4764), .A2(n4994), .B1(n4763), .B2(n4768), .ZN(n4765)
         );
  OAI211_X1 U5343 ( .C1(n5002), .C2(n4767), .A(n4766), .B(n4765), .ZN(n4851)
         );
  MUX2_X1 U5344 ( .A(REG1_REG_16__SCAN_IN), .B(n4851), .S(n5019), .Z(U3534) );
  AOI22_X1 U5345 ( .A1(n4770), .A2(n4994), .B1(n4769), .B2(n4768), .ZN(n4771)
         );
  OAI211_X1 U5346 ( .C1(n5002), .C2(n4773), .A(n4772), .B(n4771), .ZN(n4852)
         );
  MUX2_X1 U5347 ( .A(REG1_REG_15__SCAN_IN), .B(n4852), .S(n5019), .Z(U3533) );
  OAI22_X1 U5348 ( .A1(n4775), .A2(n5002), .B1(n4795), .B2(n4774), .ZN(n4776)
         );
  NOR2_X1 U5349 ( .A1(n4777), .A2(n4776), .ZN(n4853) );
  MUX2_X1 U5350 ( .A(n4778), .B(n4853), .S(n5019), .Z(n4779) );
  OAI21_X1 U5351 ( .B1(n4801), .B2(n4856), .A(n4779), .ZN(U3532) );
  AOI21_X1 U5352 ( .B1(n4998), .B2(n4781), .A(n4780), .ZN(n4857) );
  MUX2_X1 U5353 ( .A(n4782), .B(n4857), .S(n5019), .Z(n4783) );
  OAI21_X1 U5354 ( .B1(n4801), .B2(n4860), .A(n4783), .ZN(U3531) );
  NOR2_X1 U5355 ( .A1(n4784), .A2(n4795), .ZN(n4786) );
  AOI211_X1 U5356 ( .C1(n5007), .C2(n4787), .A(n4786), .B(n4785), .ZN(n4861)
         );
  MUX2_X1 U5357 ( .A(n4788), .B(n4861), .S(n5019), .Z(n4789) );
  OAI21_X1 U5358 ( .B1(n4801), .B2(n4864), .A(n4789), .ZN(U3530) );
  AOI21_X1 U5359 ( .B1(n4998), .B2(n4791), .A(n4790), .ZN(n4865) );
  MUX2_X1 U5360 ( .A(n4792), .B(n4865), .S(n5019), .Z(n4793) );
  OAI21_X1 U5361 ( .B1(n4801), .B2(n4868), .A(n4793), .ZN(U3529) );
  OAI22_X1 U5362 ( .A1(n4796), .A2(n5002), .B1(n4795), .B2(n4794), .ZN(n4797)
         );
  NOR2_X1 U5363 ( .A1(n4798), .A2(n4797), .ZN(n4869) );
  MUX2_X1 U5364 ( .A(n4799), .B(n4869), .S(n5019), .Z(n4800) );
  OAI21_X1 U5365 ( .B1(n4801), .B2(n4873), .A(n4800), .ZN(U3528) );
  AOI21_X1 U5366 ( .B1(n4803), .B2(n5007), .A(n4802), .ZN(n4877) );
  AOI22_X1 U5367 ( .A1(n4875), .A2(n4804), .B1(REG1_REG_9__SCAN_IN), .B2(n5017), .ZN(n4805) );
  OAI21_X1 U5368 ( .B1(n4877), .B2(n5017), .A(n4805), .ZN(U3527) );
  NAND2_X1 U5369 ( .A1(n5013), .A2(n4806), .ZN(n4808) );
  NAND2_X1 U5370 ( .A1(n5012), .A2(REG0_REG_31__SCAN_IN), .ZN(n4807) );
  OAI211_X1 U5371 ( .C1(n4809), .C2(n4872), .A(n4808), .B(n4807), .ZN(U3517)
         );
  NAND2_X1 U5372 ( .A1(n4810), .A2(n4874), .ZN(n4813) );
  NAND2_X1 U5373 ( .A1(n5013), .A2(n4811), .ZN(n4812) );
  OAI211_X1 U5374 ( .C1(n5013), .C2(n4814), .A(n4813), .B(n4812), .ZN(U3516)
         );
  MUX2_X1 U5375 ( .A(REG0_REG_29__SCAN_IN), .B(n4815), .S(n5013), .Z(U3515) );
  MUX2_X1 U5376 ( .A(REG0_REG_27__SCAN_IN), .B(n4816), .S(n5013), .Z(U3513) );
  MUX2_X1 U5377 ( .A(n4818), .B(n4817), .S(n5013), .Z(n4819) );
  OAI21_X1 U5378 ( .B1(n4820), .B2(n4872), .A(n4819), .ZN(U3512) );
  MUX2_X1 U5379 ( .A(n4822), .B(n4821), .S(n5013), .Z(n4823) );
  OAI21_X1 U5380 ( .B1(n4824), .B2(n4872), .A(n4823), .ZN(U3511) );
  MUX2_X1 U5381 ( .A(n4826), .B(n4825), .S(n5013), .Z(n4827) );
  OAI21_X1 U5382 ( .B1(n4828), .B2(n4872), .A(n4827), .ZN(U3510) );
  MUX2_X1 U5383 ( .A(n4830), .B(n4829), .S(n5013), .Z(n4831) );
  OAI21_X1 U5384 ( .B1(n4832), .B2(n4872), .A(n4831), .ZN(U3509) );
  MUX2_X1 U5385 ( .A(REG0_REG_22__SCAN_IN), .B(n4833), .S(n5013), .Z(U3508) );
  MUX2_X1 U5386 ( .A(n4835), .B(n4834), .S(n5013), .Z(n4836) );
  OAI21_X1 U5387 ( .B1(n4837), .B2(n4872), .A(n4836), .ZN(U3507) );
  MUX2_X1 U5388 ( .A(n4839), .B(n4838), .S(n5013), .Z(n4840) );
  OAI21_X1 U5389 ( .B1(n4841), .B2(n4872), .A(n4840), .ZN(U3506) );
  MUX2_X1 U5390 ( .A(n4843), .B(n4842), .S(n5013), .Z(n4844) );
  OAI21_X1 U5391 ( .B1(n4845), .B2(n4872), .A(n4844), .ZN(U3505) );
  MUX2_X1 U5392 ( .A(REG0_REG_18__SCAN_IN), .B(n4846), .S(n5013), .Z(U3503) );
  MUX2_X1 U5393 ( .A(n4848), .B(n4847), .S(n5013), .Z(n4849) );
  OAI21_X1 U5394 ( .B1(n4850), .B2(n4872), .A(n4849), .ZN(U3501) );
  MUX2_X1 U5395 ( .A(REG0_REG_16__SCAN_IN), .B(n4851), .S(n5013), .Z(U3499) );
  MUX2_X1 U5396 ( .A(REG0_REG_15__SCAN_IN), .B(n4852), .S(n5013), .Z(U3497) );
  MUX2_X1 U5397 ( .A(n4854), .B(n4853), .S(n5013), .Z(n4855) );
  OAI21_X1 U5398 ( .B1(n4856), .B2(n4872), .A(n4855), .ZN(U3495) );
  MUX2_X1 U5399 ( .A(n4858), .B(n4857), .S(n5013), .Z(n4859) );
  OAI21_X1 U5400 ( .B1(n4860), .B2(n4872), .A(n4859), .ZN(U3493) );
  MUX2_X1 U5401 ( .A(n4862), .B(n4861), .S(n5013), .Z(n4863) );
  OAI21_X1 U5402 ( .B1(n4864), .B2(n4872), .A(n4863), .ZN(U3491) );
  MUX2_X1 U5403 ( .A(n4866), .B(n4865), .S(n5013), .Z(n4867) );
  OAI21_X1 U5404 ( .B1(n4868), .B2(n4872), .A(n4867), .ZN(U3489) );
  MUX2_X1 U5405 ( .A(n4870), .B(n4869), .S(n5013), .Z(n4871) );
  OAI21_X1 U5406 ( .B1(n4873), .B2(n4872), .A(n4871), .ZN(U3487) );
  AOI22_X1 U5407 ( .A1(n4875), .A2(n4874), .B1(REG0_REG_9__SCAN_IN), .B2(n5012), .ZN(n4876) );
  OAI21_X1 U5408 ( .B1(n4877), .B2(n5012), .A(n4876), .ZN(U3485) );
  MUX2_X1 U5409 ( .A(DATAI_26_), .B(n4878), .S(STATE_REG_SCAN_IN), .Z(U3326)
         );
  MUX2_X1 U5410 ( .A(DATAI_22_), .B(n4879), .S(STATE_REG_SCAN_IN), .Z(U3330)
         );
  MUX2_X1 U5411 ( .A(DATAI_20_), .B(n4880), .S(STATE_REG_SCAN_IN), .Z(U3332)
         );
  MUX2_X1 U5412 ( .A(DATAI_19_), .B(n4881), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U5413 ( .A(n4882), .B(DATAI_13_), .S(U3149), .Z(U3339) );
  MUX2_X1 U5414 ( .A(DATAI_12_), .B(n4883), .S(STATE_REG_SCAN_IN), .Z(U3340)
         );
  MUX2_X1 U5415 ( .A(n4884), .B(DATAI_9_), .S(U3149), .Z(U3343) );
  MUX2_X1 U5416 ( .A(DATAI_6_), .B(n4885), .S(STATE_REG_SCAN_IN), .Z(U3346) );
  MUX2_X1 U5417 ( .A(DATAI_3_), .B(n4886), .S(STATE_REG_SCAN_IN), .Z(U3349) );
  MUX2_X1 U5418 ( .A(n2521), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  INV_X1 U5419 ( .A(DATAI_28_), .ZN(n4887) );
  AOI22_X1 U5420 ( .A1(STATE_REG_SCAN_IN), .A2(n4888), .B1(n4887), .B2(U3149), 
        .ZN(U3324) );
  XNOR2_X1 U5421 ( .A(n4890), .B(n4889), .ZN(n4891) );
  NAND2_X1 U5422 ( .A1(n4935), .A2(n4891), .ZN(n4900) );
  INV_X1 U5423 ( .A(REG2_REG_4__SCAN_IN), .ZN(n4892) );
  XNOR2_X1 U5424 ( .A(n4893), .B(n4892), .ZN(n4894) );
  NAND2_X1 U5425 ( .A1(n4948), .A2(n4894), .ZN(n4899) );
  AOI21_X1 U5426 ( .B1(n4942), .B2(ADDR_REG_4__SCAN_IN), .A(n4895), .ZN(n4898)
         );
  OR2_X1 U5427 ( .A1(n4949), .A2(n4896), .ZN(n4897) );
  AND4_X1 U5428 ( .A1(n4900), .A2(n4899), .A3(n4898), .A4(n4897), .ZN(n4902)
         );
  NAND2_X1 U5429 ( .A1(n4902), .A2(n4901), .ZN(U3244) );
  AOI211_X1 U5430 ( .C1(n4905), .C2(n4904), .A(n4903), .B(n4938), .ZN(n4906)
         );
  AOI211_X1 U5431 ( .C1(n4942), .C2(ADDR_REG_15__SCAN_IN), .A(n4907), .B(n4906), .ZN(n4913) );
  AOI21_X1 U5432 ( .B1(n4910), .B2(n4909), .A(n4908), .ZN(n4911) );
  NAND2_X1 U5433 ( .A1(n4948), .A2(n4911), .ZN(n4912) );
  OAI211_X1 U5434 ( .C1(n4949), .C2(n4985), .A(n4913), .B(n4912), .ZN(U3255)
         );
  INV_X1 U5435 ( .A(n4914), .ZN(n4915) );
  AOI21_X1 U5436 ( .B1(n4942), .B2(ADDR_REG_16__SCAN_IN), .A(n4915), .ZN(n4925) );
  OAI21_X1 U5437 ( .B1(n4918), .B2(n4917), .A(n4916), .ZN(n4923) );
  OAI21_X1 U5438 ( .B1(n4921), .B2(n4920), .A(n4919), .ZN(n4922) );
  AOI22_X1 U5439 ( .A1(n4935), .A2(n4923), .B1(n4948), .B2(n4922), .ZN(n4924)
         );
  OAI211_X1 U5440 ( .C1(n4983), .C2(n4949), .A(n4925), .B(n4924), .ZN(U3256)
         );
  AOI21_X1 U5441 ( .B1(n4942), .B2(ADDR_REG_17__SCAN_IN), .A(n4926), .ZN(n4937) );
  OAI21_X1 U5442 ( .B1(n4929), .B2(n4928), .A(n4927), .ZN(n4934) );
  OAI21_X1 U5443 ( .B1(n4932), .B2(n4931), .A(n4930), .ZN(n4933) );
  AOI22_X1 U5444 ( .A1(n4935), .A2(n4934), .B1(n4948), .B2(n4933), .ZN(n4936)
         );
  OAI211_X1 U5445 ( .C1(n4981), .C2(n4949), .A(n4937), .B(n4936), .ZN(U3257)
         );
  AOI21_X1 U5446 ( .B1(n4952), .B2(n4951), .A(n4950), .ZN(n4958) );
  AOI22_X1 U5447 ( .A1(n4955), .A2(n4954), .B1(REG3_REG_0__SCAN_IN), .B2(n4953), .ZN(n4956) );
  OAI221_X1 U5448 ( .B1(n2142), .B2(n4958), .C1(n4957), .C2(n3226), .A(n4956), 
        .ZN(U3290) );
  NOR2_X1 U5449 ( .A1(n4977), .A2(n4959), .ZN(U3291) );
  NOR2_X1 U5450 ( .A1(n4977), .A2(n4960), .ZN(U3292) );
  NOR2_X1 U5451 ( .A1(n4977), .A2(n4961), .ZN(U3293) );
  NOR2_X1 U5452 ( .A1(n4977), .A2(n4962), .ZN(U3294) );
  AND2_X1 U5453 ( .A1(D_REG_27__SCAN_IN), .A2(n4975), .ZN(U3295) );
  NOR2_X1 U5454 ( .A1(n4977), .A2(n4963), .ZN(U3296) );
  NOR2_X1 U5455 ( .A1(n4977), .A2(n4964), .ZN(U3297) );
  AND2_X1 U5456 ( .A1(D_REG_24__SCAN_IN), .A2(n4975), .ZN(U3298) );
  NOR2_X1 U5457 ( .A1(n4977), .A2(n4965), .ZN(U3299) );
  AND2_X1 U5458 ( .A1(D_REG_22__SCAN_IN), .A2(n4975), .ZN(U3300) );
  NOR2_X1 U5459 ( .A1(n4977), .A2(n4966), .ZN(U3301) );
  NOR2_X1 U5460 ( .A1(n4977), .A2(n4967), .ZN(U3302) );
  NOR2_X1 U5461 ( .A1(n4977), .A2(n4968), .ZN(U3303) );
  NOR2_X1 U5462 ( .A1(n4977), .A2(n4969), .ZN(U3304) );
  NOR2_X1 U5463 ( .A1(n4977), .A2(n4970), .ZN(U3305) );
  AND2_X1 U5464 ( .A1(D_REG_16__SCAN_IN), .A2(n4975), .ZN(U3306) );
  AND2_X1 U5465 ( .A1(D_REG_15__SCAN_IN), .A2(n4975), .ZN(U3307) );
  NOR2_X1 U5466 ( .A1(n4977), .A2(n4971), .ZN(U3308) );
  AND2_X1 U5467 ( .A1(D_REG_13__SCAN_IN), .A2(n4975), .ZN(U3309) );
  AND2_X1 U5468 ( .A1(D_REG_12__SCAN_IN), .A2(n4975), .ZN(U3310) );
  NOR2_X1 U5469 ( .A1(n4977), .A2(n4972), .ZN(U3311) );
  AND2_X1 U5470 ( .A1(D_REG_10__SCAN_IN), .A2(n4975), .ZN(U3312) );
  AND2_X1 U5471 ( .A1(D_REG_9__SCAN_IN), .A2(n4975), .ZN(U3313) );
  NOR2_X1 U5472 ( .A1(n4977), .A2(n4973), .ZN(U3314) );
  AND2_X1 U5473 ( .A1(D_REG_7__SCAN_IN), .A2(n4975), .ZN(U3315) );
  AND2_X1 U5474 ( .A1(D_REG_6__SCAN_IN), .A2(n4975), .ZN(U3316) );
  AND2_X1 U5475 ( .A1(D_REG_5__SCAN_IN), .A2(n4975), .ZN(U3317) );
  NOR2_X1 U5476 ( .A1(n4977), .A2(n4974), .ZN(U3318) );
  AND2_X1 U5477 ( .A1(D_REG_3__SCAN_IN), .A2(n4975), .ZN(U3319) );
  NOR2_X1 U5478 ( .A1(n4977), .A2(n4976), .ZN(U3320) );
  INV_X1 U5479 ( .A(DATAI_23_), .ZN(n4979) );
  AOI21_X1 U5480 ( .B1(U3149), .B2(n4979), .A(n4978), .ZN(U3329) );
  AOI22_X1 U5481 ( .A1(STATE_REG_SCAN_IN), .A2(n4980), .B1(n2727), .B2(U3149), 
        .ZN(U3334) );
  AOI22_X1 U5482 ( .A1(STATE_REG_SCAN_IN), .A2(n4981), .B1(n2716), .B2(U3149), 
        .ZN(U3335) );
  INV_X1 U5483 ( .A(DATAI_16_), .ZN(n4982) );
  AOI22_X1 U5484 ( .A1(STATE_REG_SCAN_IN), .A2(n4983), .B1(n4982), .B2(U3149), 
        .ZN(U3336) );
  INV_X1 U5485 ( .A(DATAI_15_), .ZN(n4984) );
  AOI22_X1 U5486 ( .A1(STATE_REG_SCAN_IN), .A2(n4985), .B1(n4984), .B2(U3149), 
        .ZN(U3337) );
  INV_X1 U5487 ( .A(DATAI_0_), .ZN(n4986) );
  AOI22_X1 U5488 ( .A1(STATE_REG_SCAN_IN), .A2(n2303), .B1(n4986), .B2(U3149), 
        .ZN(U3352) );
  AOI22_X1 U5489 ( .A1(n5013), .A2(n4987), .B1(n2534), .B2(n5012), .ZN(U3467)
         );
  AOI22_X1 U5490 ( .A1(n5013), .A2(n4988), .B1(n2522), .B2(n5012), .ZN(U3469)
         );
  NOR2_X1 U5491 ( .A1(n4990), .A2(n4989), .ZN(n4992) );
  AOI211_X1 U5492 ( .C1(n4994), .C2(n4993), .A(n4992), .B(n4991), .ZN(n5014)
         );
  AOI22_X1 U5493 ( .A1(n5013), .A2(n5014), .B1(n2544), .B2(n5012), .ZN(U3473)
         );
  INV_X1 U5494 ( .A(n4995), .ZN(n4997) );
  AOI211_X1 U5495 ( .C1(n4999), .C2(n4998), .A(n4997), .B(n4996), .ZN(n5015)
         );
  AOI22_X1 U5496 ( .A1(n5013), .A2(n5015), .B1(n2553), .B2(n5012), .ZN(U3475)
         );
  OAI22_X1 U5497 ( .A1(n5003), .A2(n5002), .B1(n5001), .B2(n5000), .ZN(n5005)
         );
  NOR2_X1 U5498 ( .A1(n5005), .A2(n5004), .ZN(n5016) );
  AOI22_X1 U5499 ( .A1(n5013), .A2(n5016), .B1(n2585), .B2(n5012), .ZN(U3477)
         );
  NAND3_X1 U5500 ( .A1(n5008), .A2(n5007), .A3(n5006), .ZN(n5009) );
  AND3_X1 U5501 ( .A1(n5011), .A2(n5010), .A3(n5009), .ZN(n5018) );
  AOI22_X1 U5502 ( .A1(n5013), .A2(n5018), .B1(n2565), .B2(n5012), .ZN(U3481)
         );
  AOI22_X1 U5503 ( .A1(n5019), .A2(n5014), .B1(n2545), .B2(n5017), .ZN(U3521)
         );
  AOI22_X1 U5504 ( .A1(n5019), .A2(n5015), .B1(n4889), .B2(n5017), .ZN(U3522)
         );
  AOI22_X1 U5505 ( .A1(n5019), .A2(n5016), .B1(n2586), .B2(n5017), .ZN(U3523)
         );
  AOI22_X1 U5506 ( .A1(n5019), .A2(n5018), .B1(n3298), .B2(n5017), .ZN(U3525)
         );
  OR2_X1 U3730 ( .A1(n3329), .A2(n4880), .ZN(n5000) );
  INV_X2 U2385 ( .A(n3874), .ZN(n3796) );
  CLKBUF_X2 U2420 ( .A(n3420), .Z(n3831) );
  CLKBUF_X1 U2461 ( .A(n4186), .Z(n2143) );
endmodule

