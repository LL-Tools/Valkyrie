

module b17_C_AntiSAT_k_256_2 ( P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, 
        DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_, DATAI_25_, 
        DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_, DATAI_19_, 
        DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_, DATAI_13_, 
        DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_, DATAI_7_, 
        DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_, DATAI_0_, 
        HOLD, NA, BS16, READY1, READY2, P1_READREQUEST_REG_SCAN_IN, 
        P1_ADS_N_REG_SCAN_IN, P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, 
        P1_D_C_N_REG_SCAN_IN, P1_REQUESTPENDING_REG_SCAN_IN, 
        P1_STATEBS16_REG_SCAN_IN, P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, 
        P1_W_R_N_REG_SCAN_IN, P1_BYTEENABLE_REG_0__SCAN_IN, 
        P1_BYTEENABLE_REG_1__SCAN_IN, P1_BYTEENABLE_REG_2__SCAN_IN, 
        P1_BYTEENABLE_REG_3__SCAN_IN, P1_REIP_REG_31__SCAN_IN, 
        P1_REIP_REG_30__SCAN_IN, P1_REIP_REG_29__SCAN_IN, 
        P1_REIP_REG_28__SCAN_IN, P1_REIP_REG_27__SCAN_IN, 
        P1_REIP_REG_26__SCAN_IN, P1_REIP_REG_25__SCAN_IN, 
        P1_REIP_REG_24__SCAN_IN, P1_REIP_REG_23__SCAN_IN, 
        P1_REIP_REG_22__SCAN_IN, P1_REIP_REG_21__SCAN_IN, 
        P1_REIP_REG_20__SCAN_IN, P1_REIP_REG_19__SCAN_IN, 
        P1_REIP_REG_18__SCAN_IN, P1_REIP_REG_17__SCAN_IN, 
        P1_REIP_REG_16__SCAN_IN, P1_REIP_REG_15__SCAN_IN, 
        P1_REIP_REG_14__SCAN_IN, P1_REIP_REG_13__SCAN_IN, 
        P1_REIP_REG_12__SCAN_IN, P1_REIP_REG_11__SCAN_IN, 
        P1_REIP_REG_10__SCAN_IN, P1_REIP_REG_9__SCAN_IN, 
        P1_REIP_REG_8__SCAN_IN, P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN, 
        P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN, P1_REIP_REG_3__SCAN_IN, 
        P1_REIP_REG_2__SCAN_IN, P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN, 
        P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN, P1_EBX_REG_29__SCAN_IN, 
        P1_EBX_REG_28__SCAN_IN, P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN, 
        P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN, P1_EBX_REG_23__SCAN_IN, 
        P1_EBX_REG_22__SCAN_IN, P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN, 
        P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN, P1_EBX_REG_17__SCAN_IN, 
        P1_EBX_REG_16__SCAN_IN, P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN, 
        P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN, P1_EBX_REG_11__SCAN_IN, 
        P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN, P1_EBX_REG_8__SCAN_IN, 
        P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN, P1_EBX_REG_5__SCAN_IN, 
        P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN, P1_EBX_REG_2__SCAN_IN, 
        P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN, P1_EAX_REG_31__SCAN_IN, 
        P1_EAX_REG_30__SCAN_IN, P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN, 
        P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN, P1_EAX_REG_25__SCAN_IN, 
        P1_EAX_REG_24__SCAN_IN, P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN, 
        P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN, P1_EAX_REG_19__SCAN_IN, 
        P1_EAX_REG_18__SCAN_IN, P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN, 
        P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN, P1_EAX_REG_13__SCAN_IN, 
        P1_EAX_REG_12__SCAN_IN, P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, 
        P1_EAX_REG_9__SCAN_IN, P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, 
        P1_EAX_REG_6__SCAN_IN, P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, 
        P1_EAX_REG_3__SCAN_IN, P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, 
        P1_EAX_REG_0__SCAN_IN, P1_DATAO_REG_31__SCAN_IN, 
        P1_DATAO_REG_30__SCAN_IN, P1_DATAO_REG_29__SCAN_IN, 
        P1_DATAO_REG_28__SCAN_IN, P1_DATAO_REG_27__SCAN_IN, 
        P1_DATAO_REG_26__SCAN_IN, P1_DATAO_REG_25__SCAN_IN, 
        P1_DATAO_REG_24__SCAN_IN, P1_DATAO_REG_23__SCAN_IN, 
        P1_DATAO_REG_22__SCAN_IN, P1_DATAO_REG_21__SCAN_IN, 
        P1_DATAO_REG_20__SCAN_IN, P1_DATAO_REG_19__SCAN_IN, 
        P1_DATAO_REG_18__SCAN_IN, P1_DATAO_REG_17__SCAN_IN, 
        P1_DATAO_REG_16__SCAN_IN, P1_DATAO_REG_15__SCAN_IN, 
        P1_DATAO_REG_14__SCAN_IN, P1_DATAO_REG_13__SCAN_IN, 
        P1_DATAO_REG_12__SCAN_IN, P1_DATAO_REG_11__SCAN_IN, 
        P1_DATAO_REG_10__SCAN_IN, P1_DATAO_REG_9__SCAN_IN, 
        P1_DATAO_REG_8__SCAN_IN, P1_DATAO_REG_7__SCAN_IN, 
        P1_DATAO_REG_6__SCAN_IN, P1_DATAO_REG_5__SCAN_IN, 
        P1_DATAO_REG_4__SCAN_IN, P1_DATAO_REG_3__SCAN_IN, 
        P1_DATAO_REG_2__SCAN_IN, P1_DATAO_REG_1__SCAN_IN, 
        P1_DATAO_REG_0__SCAN_IN, P1_UWORD_REG_0__SCAN_IN, 
        P1_UWORD_REG_1__SCAN_IN, P1_UWORD_REG_2__SCAN_IN, 
        P1_UWORD_REG_3__SCAN_IN, P1_UWORD_REG_4__SCAN_IN, 
        P1_UWORD_REG_5__SCAN_IN, P1_UWORD_REG_6__SCAN_IN, 
        P1_UWORD_REG_7__SCAN_IN, P1_UWORD_REG_8__SCAN_IN, 
        P1_UWORD_REG_9__SCAN_IN, P1_UWORD_REG_10__SCAN_IN, 
        P1_UWORD_REG_11__SCAN_IN, P1_UWORD_REG_12__SCAN_IN, 
        P1_UWORD_REG_13__SCAN_IN, P1_UWORD_REG_14__SCAN_IN, 
        P1_LWORD_REG_0__SCAN_IN, P1_LWORD_REG_1__SCAN_IN, 
        P1_LWORD_REG_2__SCAN_IN, P1_LWORD_REG_3__SCAN_IN, 
        P1_LWORD_REG_4__SCAN_IN, P1_LWORD_REG_5__SCAN_IN, 
        P1_LWORD_REG_6__SCAN_IN, P1_LWORD_REG_7__SCAN_IN, 
        P1_LWORD_REG_8__SCAN_IN, P1_LWORD_REG_9__SCAN_IN, 
        P1_LWORD_REG_10__SCAN_IN, P1_LWORD_REG_11__SCAN_IN, 
        P1_LWORD_REG_12__SCAN_IN, P1_LWORD_REG_13__SCAN_IN, 
        P1_LWORD_REG_14__SCAN_IN, P1_LWORD_REG_15__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_31__SCAN_IN, P1_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_29__SCAN_IN, P1_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_27__SCAN_IN, P1_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_25__SCAN_IN, P1_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_23__SCAN_IN, P1_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_21__SCAN_IN, P1_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_19__SCAN_IN, P1_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_17__SCAN_IN, P1_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_13__SCAN_IN, P1_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_11__SCAN_IN, P1_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_9__SCAN_IN, P1_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_7__SCAN_IN, P1_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_5__SCAN_IN, P1_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_3__SCAN_IN, P1_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P1_PHYADDRPOINTER_REG_1__SCAN_IN, P1_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_31__SCAN_IN, P1_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_29__SCAN_IN, P1_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_27__SCAN_IN, P1_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_25__SCAN_IN, P1_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_23__SCAN_IN, P1_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_21__SCAN_IN, P1_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_19__SCAN_IN, P1_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_17__SCAN_IN, P1_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_15__SCAN_IN, P1_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_13__SCAN_IN, P1_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_11__SCAN_IN, P1_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_9__SCAN_IN, P1_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_7__SCAN_IN, P1_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_5__SCAN_IN, P1_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_3__SCAN_IN, P1_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P1_INSTADDRPOINTER_REG_1__SCAN_IN, P1_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P1_INSTQUEUE_REG_0__0__SCAN_IN, P1_INSTQUEUE_REG_0__1__SCAN_IN, 
        P1_INSTQUEUE_REG_0__2__SCAN_IN, P1_INSTQUEUE_REG_0__3__SCAN_IN, 
        P1_INSTQUEUE_REG_0__4__SCAN_IN, P1_INSTQUEUE_REG_0__5__SCAN_IN, 
        P1_INSTQUEUE_REG_0__6__SCAN_IN, P1_INSTQUEUE_REG_0__7__SCAN_IN, 
        P1_INSTQUEUE_REG_1__0__SCAN_IN, P1_INSTQUEUE_REG_1__1__SCAN_IN, 
        P1_INSTQUEUE_REG_1__2__SCAN_IN, P1_INSTQUEUE_REG_1__3__SCAN_IN, 
        P1_INSTQUEUE_REG_1__4__SCAN_IN, P1_INSTQUEUE_REG_1__5__SCAN_IN, 
        P1_INSTQUEUE_REG_1__6__SCAN_IN, P1_INSTQUEUE_REG_1__7__SCAN_IN, 
        P1_INSTQUEUE_REG_2__0__SCAN_IN, P1_INSTQUEUE_REG_2__1__SCAN_IN, 
        P1_INSTQUEUE_REG_2__2__SCAN_IN, P1_INSTQUEUE_REG_2__3__SCAN_IN, 
        P1_INSTQUEUE_REG_2__4__SCAN_IN, P1_INSTQUEUE_REG_2__5__SCAN_IN, 
        P1_INSTQUEUE_REG_2__6__SCAN_IN, P1_INSTQUEUE_REG_2__7__SCAN_IN, 
        P1_INSTQUEUE_REG_3__0__SCAN_IN, P1_INSTQUEUE_REG_3__1__SCAN_IN, 
        P1_INSTQUEUE_REG_3__2__SCAN_IN, P1_INSTQUEUE_REG_3__3__SCAN_IN, 
        P1_INSTQUEUE_REG_3__4__SCAN_IN, P1_INSTQUEUE_REG_3__5__SCAN_IN, 
        P1_INSTQUEUE_REG_3__6__SCAN_IN, P1_INSTQUEUE_REG_3__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__0__SCAN_IN, BUF1_REG_0__SCAN_IN, 
        BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN, BUF1_REG_3__SCAN_IN, 
        BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN, BUF1_REG_6__SCAN_IN, 
        BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN, BUF1_REG_9__SCAN_IN, 
        BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN, BUF1_REG_12__SCAN_IN, 
        BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN, BUF1_REG_15__SCAN_IN, 
        BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN, BUF1_REG_18__SCAN_IN, 
        BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN, BUF1_REG_21__SCAN_IN, 
        BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN, BUF1_REG_24__SCAN_IN, 
        BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN, BUF1_REG_27__SCAN_IN, 
        BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN, BUF1_REG_30__SCAN_IN, 
        BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN, BUF2_REG_1__SCAN_IN, 
        BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN, BUF2_REG_4__SCAN_IN, 
        BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN, BUF2_REG_7__SCAN_IN, 
        BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN, BUF2_REG_10__SCAN_IN, 
        BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN, BUF2_REG_13__SCAN_IN, 
        BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN, BUF2_REG_16__SCAN_IN, 
        BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN, BUF2_REG_19__SCAN_IN, 
        BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN, BUF2_REG_22__SCAN_IN, 
        BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN, BUF2_REG_25__SCAN_IN, 
        BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN, BUF2_REG_28__SCAN_IN, 
        BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN, BUF2_REG_31__SCAN_IN, 
        READY12_REG_SCAN_IN, READY21_REG_SCAN_IN, READY22_REG_SCAN_IN, 
        READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN, P3_BE_N_REG_2__SCAN_IN, 
        P3_BE_N_REG_1__SCAN_IN, P3_BE_N_REG_0__SCAN_IN, 
        P3_ADDRESS_REG_29__SCAN_IN, P3_ADDRESS_REG_28__SCAN_IN, 
        P3_ADDRESS_REG_27__SCAN_IN, P3_ADDRESS_REG_26__SCAN_IN, 
        P3_ADDRESS_REG_25__SCAN_IN, P3_ADDRESS_REG_24__SCAN_IN, 
        P3_ADDRESS_REG_23__SCAN_IN, P3_ADDRESS_REG_22__SCAN_IN, 
        P3_ADDRESS_REG_21__SCAN_IN, P3_ADDRESS_REG_20__SCAN_IN, 
        P3_ADDRESS_REG_19__SCAN_IN, P3_ADDRESS_REG_18__SCAN_IN, 
        P3_ADDRESS_REG_17__SCAN_IN, P3_ADDRESS_REG_16__SCAN_IN, 
        P3_ADDRESS_REG_15__SCAN_IN, P3_ADDRESS_REG_14__SCAN_IN, 
        P3_ADDRESS_REG_13__SCAN_IN, P3_ADDRESS_REG_12__SCAN_IN, 
        P3_ADDRESS_REG_11__SCAN_IN, P3_ADDRESS_REG_10__SCAN_IN, 
        P3_ADDRESS_REG_9__SCAN_IN, P3_ADDRESS_REG_8__SCAN_IN, 
        P3_ADDRESS_REG_7__SCAN_IN, P3_ADDRESS_REG_6__SCAN_IN, 
        P3_ADDRESS_REG_5__SCAN_IN, P3_ADDRESS_REG_4__SCAN_IN, 
        P3_ADDRESS_REG_3__SCAN_IN, P3_ADDRESS_REG_2__SCAN_IN, 
        P3_ADDRESS_REG_1__SCAN_IN, P3_ADDRESS_REG_0__SCAN_IN, 
        P3_STATE_REG_2__SCAN_IN, P3_STATE_REG_1__SCAN_IN, 
        P3_STATE_REG_0__SCAN_IN, P3_DATAWIDTH_REG_0__SCAN_IN, 
        P3_DATAWIDTH_REG_1__SCAN_IN, P3_DATAWIDTH_REG_2__SCAN_IN, 
        P3_DATAWIDTH_REG_3__SCAN_IN, P3_DATAWIDTH_REG_4__SCAN_IN, 
        P3_DATAWIDTH_REG_5__SCAN_IN, P3_DATAWIDTH_REG_6__SCAN_IN, 
        P3_DATAWIDTH_REG_7__SCAN_IN, P3_DATAWIDTH_REG_8__SCAN_IN, 
        P3_DATAWIDTH_REG_9__SCAN_IN, P3_DATAWIDTH_REG_10__SCAN_IN, 
        P3_DATAWIDTH_REG_11__SCAN_IN, P3_DATAWIDTH_REG_12__SCAN_IN, 
        P3_DATAWIDTH_REG_13__SCAN_IN, P3_DATAWIDTH_REG_14__SCAN_IN, 
        P3_DATAWIDTH_REG_15__SCAN_IN, P3_DATAWIDTH_REG_16__SCAN_IN, 
        P3_DATAWIDTH_REG_17__SCAN_IN, P3_DATAWIDTH_REG_18__SCAN_IN, 
        P3_DATAWIDTH_REG_19__SCAN_IN, P3_DATAWIDTH_REG_20__SCAN_IN, 
        P3_DATAWIDTH_REG_21__SCAN_IN, P3_DATAWIDTH_REG_22__SCAN_IN, 
        P3_DATAWIDTH_REG_23__SCAN_IN, P3_DATAWIDTH_REG_24__SCAN_IN, 
        P3_DATAWIDTH_REG_25__SCAN_IN, P3_DATAWIDTH_REG_26__SCAN_IN, 
        P3_DATAWIDTH_REG_27__SCAN_IN, P3_DATAWIDTH_REG_28__SCAN_IN, 
        P3_DATAWIDTH_REG_29__SCAN_IN, P3_DATAWIDTH_REG_30__SCAN_IN, 
        P3_DATAWIDTH_REG_31__SCAN_IN, P3_STATE2_REG_3__SCAN_IN, 
        P3_STATE2_REG_2__SCAN_IN, P3_STATE2_REG_1__SCAN_IN, 
        P3_STATE2_REG_0__SCAN_IN, P3_INSTQUEUE_REG_15__7__SCAN_IN, 
        P3_INSTQUEUE_REG_15__6__SCAN_IN, P3_INSTQUEUE_REG_15__5__SCAN_IN, 
        P3_INSTQUEUE_REG_15__4__SCAN_IN, P3_INSTQUEUE_REG_15__3__SCAN_IN, 
        P3_INSTQUEUE_REG_15__2__SCAN_IN, P3_INSTQUEUE_REG_15__1__SCAN_IN, 
        P3_INSTQUEUE_REG_15__0__SCAN_IN, P3_INSTQUEUE_REG_14__7__SCAN_IN, 
        P3_INSTQUEUE_REG_14__6__SCAN_IN, P3_INSTQUEUE_REG_14__5__SCAN_IN, 
        P3_INSTQUEUE_REG_14__4__SCAN_IN, P3_INSTQUEUE_REG_14__3__SCAN_IN, 
        P3_INSTQUEUE_REG_14__2__SCAN_IN, P3_INSTQUEUE_REG_14__1__SCAN_IN, 
        P3_INSTQUEUE_REG_14__0__SCAN_IN, P3_INSTQUEUE_REG_13__7__SCAN_IN, 
        P3_INSTQUEUE_REG_13__6__SCAN_IN, P3_INSTQUEUE_REG_13__5__SCAN_IN, 
        P3_INSTQUEUE_REG_13__4__SCAN_IN, P3_INSTQUEUE_REG_13__3__SCAN_IN, 
        P3_INSTQUEUE_REG_13__2__SCAN_IN, P3_INSTQUEUE_REG_13__1__SCAN_IN, 
        P3_INSTQUEUE_REG_13__0__SCAN_IN, P3_INSTQUEUE_REG_12__7__SCAN_IN, 
        P3_INSTQUEUE_REG_12__6__SCAN_IN, P3_INSTQUEUE_REG_12__5__SCAN_IN, 
        P3_INSTQUEUE_REG_12__4__SCAN_IN, P3_INSTQUEUE_REG_12__3__SCAN_IN, 
        P3_INSTQUEUE_REG_12__2__SCAN_IN, P3_INSTQUEUE_REG_12__1__SCAN_IN, 
        P3_INSTQUEUE_REG_12__0__SCAN_IN, P3_INSTQUEUE_REG_11__7__SCAN_IN, 
        P3_INSTQUEUE_REG_11__6__SCAN_IN, P3_INSTQUEUE_REG_11__5__SCAN_IN, 
        P3_INSTQUEUE_REG_11__4__SCAN_IN, P3_INSTQUEUE_REG_11__3__SCAN_IN, 
        P3_INSTQUEUE_REG_11__2__SCAN_IN, P3_INSTQUEUE_REG_11__1__SCAN_IN, 
        P3_INSTQUEUE_REG_11__0__SCAN_IN, P3_INSTQUEUE_REG_10__7__SCAN_IN, 
        P3_INSTQUEUE_REG_10__6__SCAN_IN, P3_INSTQUEUE_REG_10__5__SCAN_IN, 
        P3_INSTQUEUE_REG_10__4__SCAN_IN, P3_INSTQUEUE_REG_10__3__SCAN_IN, 
        P3_INSTQUEUE_REG_10__2__SCAN_IN, P3_INSTQUEUE_REG_10__1__SCAN_IN, 
        P3_INSTQUEUE_REG_10__0__SCAN_IN, P3_INSTQUEUE_REG_9__7__SCAN_IN, 
        P3_INSTQUEUE_REG_9__6__SCAN_IN, P3_INSTQUEUE_REG_9__5__SCAN_IN, 
        P3_INSTQUEUE_REG_9__4__SCAN_IN, P3_INSTQUEUE_REG_9__3__SCAN_IN, 
        P3_INSTQUEUE_REG_9__2__SCAN_IN, P3_INSTQUEUE_REG_9__1__SCAN_IN, 
        P3_INSTQUEUE_REG_9__0__SCAN_IN, P3_INSTQUEUE_REG_8__7__SCAN_IN, 
        P3_INSTQUEUE_REG_8__6__SCAN_IN, P3_INSTQUEUE_REG_8__5__SCAN_IN, 
        P3_INSTQUEUE_REG_8__4__SCAN_IN, P3_INSTQUEUE_REG_8__3__SCAN_IN, 
        P3_INSTQUEUE_REG_8__2__SCAN_IN, P3_INSTQUEUE_REG_8__1__SCAN_IN, 
        P3_INSTQUEUE_REG_8__0__SCAN_IN, P3_INSTQUEUE_REG_7__7__SCAN_IN, 
        P3_INSTQUEUE_REG_7__6__SCAN_IN, P3_INSTQUEUE_REG_7__5__SCAN_IN, 
        P3_INSTQUEUE_REG_7__4__SCAN_IN, P3_INSTQUEUE_REG_7__3__SCAN_IN, 
        P3_INSTQUEUE_REG_7__2__SCAN_IN, P3_INSTQUEUE_REG_7__1__SCAN_IN, 
        P3_INSTQUEUE_REG_7__0__SCAN_IN, P3_INSTQUEUE_REG_6__7__SCAN_IN, 
        P3_INSTQUEUE_REG_6__6__SCAN_IN, P3_INSTQUEUE_REG_6__5__SCAN_IN, 
        P3_INSTQUEUE_REG_6__4__SCAN_IN, P3_INSTQUEUE_REG_6__3__SCAN_IN, 
        P3_INSTQUEUE_REG_6__2__SCAN_IN, P3_INSTQUEUE_REG_6__1__SCAN_IN, 
        P3_INSTQUEUE_REG_6__0__SCAN_IN, P3_INSTQUEUE_REG_5__7__SCAN_IN, 
        P3_INSTQUEUE_REG_5__6__SCAN_IN, P3_INSTQUEUE_REG_5__5__SCAN_IN, 
        P3_INSTQUEUE_REG_5__4__SCAN_IN, P3_INSTQUEUE_REG_5__3__SCAN_IN, 
        P3_INSTQUEUE_REG_5__2__SCAN_IN, P3_INSTQUEUE_REG_5__1__SCAN_IN, 
        P3_INSTQUEUE_REG_5__0__SCAN_IN, P3_INSTQUEUE_REG_4__7__SCAN_IN, 
        P3_INSTQUEUE_REG_4__6__SCAN_IN, P3_INSTQUEUE_REG_4__5__SCAN_IN, 
        P3_INSTQUEUE_REG_4__4__SCAN_IN, P3_INSTQUEUE_REG_4__3__SCAN_IN, 
        P3_INSTQUEUE_REG_4__2__SCAN_IN, P3_INSTQUEUE_REG_4__1__SCAN_IN, 
        P3_INSTQUEUE_REG_4__0__SCAN_IN, P3_INSTQUEUE_REG_3__7__SCAN_IN, 
        P3_INSTQUEUE_REG_3__6__SCAN_IN, P3_INSTQUEUE_REG_3__5__SCAN_IN, 
        P3_INSTQUEUE_REG_3__4__SCAN_IN, P3_INSTQUEUE_REG_3__3__SCAN_IN, 
        P3_INSTQUEUE_REG_3__2__SCAN_IN, P3_INSTQUEUE_REG_3__1__SCAN_IN, 
        P3_INSTQUEUE_REG_3__0__SCAN_IN, P3_INSTQUEUE_REG_2__7__SCAN_IN, 
        P3_INSTQUEUE_REG_2__6__SCAN_IN, P3_INSTQUEUE_REG_2__5__SCAN_IN, 
        P3_INSTQUEUE_REG_2__4__SCAN_IN, P3_INSTQUEUE_REG_2__3__SCAN_IN, 
        P3_INSTQUEUE_REG_2__2__SCAN_IN, P3_INSTQUEUE_REG_2__1__SCAN_IN, 
        P3_INSTQUEUE_REG_2__0__SCAN_IN, P3_INSTQUEUE_REG_1__7__SCAN_IN, 
        P3_INSTQUEUE_REG_1__6__SCAN_IN, P3_INSTQUEUE_REG_1__5__SCAN_IN, 
        P3_INSTQUEUE_REG_1__4__SCAN_IN, P3_INSTQUEUE_REG_1__3__SCAN_IN, 
        P3_INSTQUEUE_REG_1__2__SCAN_IN, P3_INSTQUEUE_REG_1__1__SCAN_IN, 
        P3_INSTQUEUE_REG_1__0__SCAN_IN, P3_INSTQUEUE_REG_0__7__SCAN_IN, 
        P3_INSTQUEUE_REG_0__6__SCAN_IN, P3_INSTQUEUE_REG_0__5__SCAN_IN, 
        P3_INSTQUEUE_REG_0__4__SCAN_IN, P3_INSTQUEUE_REG_0__3__SCAN_IN, 
        P3_INSTQUEUE_REG_0__2__SCAN_IN, P3_INSTQUEUE_REG_0__1__SCAN_IN, 
        P3_INSTQUEUE_REG_0__0__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_11__SCAN_IN, P3_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_13__SCAN_IN, P3_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_15__SCAN_IN, P3_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_17__SCAN_IN, P3_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_19__SCAN_IN, P3_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_21__SCAN_IN, P3_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_23__SCAN_IN, P3_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_25__SCAN_IN, P3_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_27__SCAN_IN, P3_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_29__SCAN_IN, P3_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN, 
        P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN, 
        P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN, 
        P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN, 
        P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN, 
        P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN, 
        P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN, 
        P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN, 
        P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN, 
        P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN, 
        P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN, 
        P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN, 
        P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN, 
        P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN, 
        P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN, 
        P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN, 
        P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN, 
        P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN, 
        P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN, 
        P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN, 
        P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN, 
        P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN, 
        P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN, 
        P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN, 
        P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN, 
        P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN, 
        P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN, 
        P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN, 
        P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN, 
        P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN, 
        P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN, 
        P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN, 
        P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN, 
        P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN, 
        P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN, 
        P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN, 
        P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN, P3_EAX_REG_14__SCAN_IN, 
        P3_EAX_REG_15__SCAN_IN, P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN, 
        P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN, P3_EAX_REG_20__SCAN_IN, 
        P3_EAX_REG_21__SCAN_IN, P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN, 
        P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN, P3_EAX_REG_26__SCAN_IN, 
        P3_EAX_REG_27__SCAN_IN, P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN, 
        P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN, 
        P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN, 
        P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN, 
        P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN, 
        P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN, P3_EBX_REG_12__SCAN_IN, 
        P3_EBX_REG_13__SCAN_IN, P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN, 
        P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN, P3_EBX_REG_18__SCAN_IN, 
        P3_EBX_REG_19__SCAN_IN, P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN, 
        P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN, P3_EBX_REG_24__SCAN_IN, 
        P3_EBX_REG_25__SCAN_IN, P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN, 
        P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN, P3_EBX_REG_30__SCAN_IN, 
        P3_EBX_REG_31__SCAN_IN, P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN, 
        P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN, P3_REIP_REG_4__SCAN_IN, 
        P3_REIP_REG_5__SCAN_IN, P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN, 
        P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN, 
        P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN, 
        P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN, 
        P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN, 
        P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN, 
        P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN, 
        P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN, 
        P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN, 
        P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN, 
        P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN, 
        P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN, 
        P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN, 
        P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN, 
        P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN, 
        P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN, 
        P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN, 
        P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN, 
        P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN, 
        P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN, 
        P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN, P2_BE_N_REG_0__SCAN_IN, 
        P2_ADDRESS_REG_29__SCAN_IN, P2_ADDRESS_REG_28__SCAN_IN, 
        P2_ADDRESS_REG_27__SCAN_IN, P2_ADDRESS_REG_26__SCAN_IN, 
        P2_ADDRESS_REG_25__SCAN_IN, P2_ADDRESS_REG_24__SCAN_IN, 
        P2_ADDRESS_REG_23__SCAN_IN, P2_ADDRESS_REG_22__SCAN_IN, 
        P2_ADDRESS_REG_21__SCAN_IN, P2_ADDRESS_REG_20__SCAN_IN, 
        P2_ADDRESS_REG_19__SCAN_IN, P2_ADDRESS_REG_18__SCAN_IN, 
        P2_ADDRESS_REG_17__SCAN_IN, P2_ADDRESS_REG_16__SCAN_IN, 
        P2_ADDRESS_REG_15__SCAN_IN, P2_ADDRESS_REG_14__SCAN_IN, 
        P2_ADDRESS_REG_13__SCAN_IN, P2_ADDRESS_REG_12__SCAN_IN, 
        P2_ADDRESS_REG_11__SCAN_IN, P2_ADDRESS_REG_10__SCAN_IN, 
        P2_ADDRESS_REG_9__SCAN_IN, P2_ADDRESS_REG_8__SCAN_IN, 
        P2_ADDRESS_REG_7__SCAN_IN, P2_ADDRESS_REG_6__SCAN_IN, 
        P2_ADDRESS_REG_5__SCAN_IN, P2_ADDRESS_REG_4__SCAN_IN, 
        P2_ADDRESS_REG_3__SCAN_IN, P2_ADDRESS_REG_2__SCAN_IN, 
        P2_ADDRESS_REG_1__SCAN_IN, P2_ADDRESS_REG_0__SCAN_IN, 
        P2_STATE_REG_2__SCAN_IN, P2_STATE_REG_1__SCAN_IN, 
        P2_STATE_REG_0__SCAN_IN, P2_DATAWIDTH_REG_0__SCAN_IN, 
        P2_DATAWIDTH_REG_1__SCAN_IN, P2_DATAWIDTH_REG_2__SCAN_IN, 
        P2_DATAWIDTH_REG_3__SCAN_IN, P2_DATAWIDTH_REG_4__SCAN_IN, 
        P2_DATAWIDTH_REG_5__SCAN_IN, P2_DATAWIDTH_REG_6__SCAN_IN, 
        P2_DATAWIDTH_REG_7__SCAN_IN, P2_DATAWIDTH_REG_8__SCAN_IN, 
        P2_DATAWIDTH_REG_9__SCAN_IN, P2_DATAWIDTH_REG_10__SCAN_IN, 
        P2_DATAWIDTH_REG_11__SCAN_IN, P2_DATAWIDTH_REG_12__SCAN_IN, 
        P2_DATAWIDTH_REG_13__SCAN_IN, P2_DATAWIDTH_REG_14__SCAN_IN, 
        P2_DATAWIDTH_REG_15__SCAN_IN, P2_DATAWIDTH_REG_16__SCAN_IN, 
        P2_DATAWIDTH_REG_17__SCAN_IN, P2_DATAWIDTH_REG_18__SCAN_IN, 
        P2_DATAWIDTH_REG_19__SCAN_IN, P2_DATAWIDTH_REG_20__SCAN_IN, 
        P2_DATAWIDTH_REG_21__SCAN_IN, P2_DATAWIDTH_REG_22__SCAN_IN, 
        P2_DATAWIDTH_REG_23__SCAN_IN, P2_DATAWIDTH_REG_24__SCAN_IN, 
        P2_DATAWIDTH_REG_25__SCAN_IN, P2_DATAWIDTH_REG_26__SCAN_IN, 
        P2_DATAWIDTH_REG_27__SCAN_IN, P2_DATAWIDTH_REG_28__SCAN_IN, 
        P2_DATAWIDTH_REG_29__SCAN_IN, P2_DATAWIDTH_REG_30__SCAN_IN, 
        P2_DATAWIDTH_REG_31__SCAN_IN, P2_STATE2_REG_3__SCAN_IN, 
        P2_STATE2_REG_2__SCAN_IN, P2_STATE2_REG_1__SCAN_IN, 
        P2_STATE2_REG_0__SCAN_IN, P2_INSTQUEUE_REG_15__7__SCAN_IN, 
        P2_INSTQUEUE_REG_15__6__SCAN_IN, P2_INSTQUEUE_REG_15__5__SCAN_IN, 
        P2_INSTQUEUE_REG_15__4__SCAN_IN, P2_INSTQUEUE_REG_15__3__SCAN_IN, 
        P2_INSTQUEUE_REG_15__2__SCAN_IN, P2_INSTQUEUE_REG_15__1__SCAN_IN, 
        P2_INSTQUEUE_REG_15__0__SCAN_IN, P2_INSTQUEUE_REG_14__7__SCAN_IN, 
        P2_INSTQUEUE_REG_14__6__SCAN_IN, P2_INSTQUEUE_REG_14__5__SCAN_IN, 
        P2_INSTQUEUE_REG_14__4__SCAN_IN, P2_INSTQUEUE_REG_14__3__SCAN_IN, 
        P2_INSTQUEUE_REG_14__2__SCAN_IN, P2_INSTQUEUE_REG_14__1__SCAN_IN, 
        P2_INSTQUEUE_REG_14__0__SCAN_IN, P2_INSTQUEUE_REG_13__7__SCAN_IN, 
        P2_INSTQUEUE_REG_13__6__SCAN_IN, P2_INSTQUEUE_REG_13__5__SCAN_IN, 
        P2_INSTQUEUE_REG_13__4__SCAN_IN, P2_INSTQUEUE_REG_13__3__SCAN_IN, 
        P2_INSTQUEUE_REG_13__2__SCAN_IN, P2_INSTQUEUE_REG_13__1__SCAN_IN, 
        P2_INSTQUEUE_REG_13__0__SCAN_IN, P2_INSTQUEUE_REG_12__7__SCAN_IN, 
        P2_INSTQUEUE_REG_12__6__SCAN_IN, P2_INSTQUEUE_REG_12__5__SCAN_IN, 
        P2_INSTQUEUE_REG_12__4__SCAN_IN, P2_INSTQUEUE_REG_12__3__SCAN_IN, 
        P2_INSTQUEUE_REG_12__2__SCAN_IN, P2_INSTQUEUE_REG_12__1__SCAN_IN, 
        P2_INSTQUEUE_REG_12__0__SCAN_IN, P2_INSTQUEUE_REG_11__7__SCAN_IN, 
        P2_INSTQUEUE_REG_11__6__SCAN_IN, P2_INSTQUEUE_REG_11__5__SCAN_IN, 
        P2_INSTQUEUE_REG_11__4__SCAN_IN, P2_INSTQUEUE_REG_11__3__SCAN_IN, 
        P2_INSTQUEUE_REG_11__2__SCAN_IN, P2_INSTQUEUE_REG_11__1__SCAN_IN, 
        P2_INSTQUEUE_REG_11__0__SCAN_IN, P2_INSTQUEUE_REG_10__7__SCAN_IN, 
        P2_INSTQUEUE_REG_10__6__SCAN_IN, P2_INSTQUEUE_REG_10__5__SCAN_IN, 
        P2_INSTQUEUE_REG_10__4__SCAN_IN, P2_INSTQUEUE_REG_10__3__SCAN_IN, 
        P2_INSTQUEUE_REG_10__2__SCAN_IN, P2_INSTQUEUE_REG_10__1__SCAN_IN, 
        P2_INSTQUEUE_REG_10__0__SCAN_IN, P2_INSTQUEUE_REG_9__7__SCAN_IN, 
        P2_INSTQUEUE_REG_9__6__SCAN_IN, P2_INSTQUEUE_REG_9__5__SCAN_IN, 
        P2_INSTQUEUE_REG_9__4__SCAN_IN, P2_INSTQUEUE_REG_9__3__SCAN_IN, 
        P2_INSTQUEUE_REG_9__2__SCAN_IN, P2_INSTQUEUE_REG_9__1__SCAN_IN, 
        P2_INSTQUEUE_REG_9__0__SCAN_IN, P2_INSTQUEUE_REG_8__7__SCAN_IN, 
        P2_INSTQUEUE_REG_8__6__SCAN_IN, P2_INSTQUEUE_REG_8__5__SCAN_IN, 
        P2_INSTQUEUE_REG_8__4__SCAN_IN, P2_INSTQUEUE_REG_8__3__SCAN_IN, 
        P2_INSTQUEUE_REG_8__2__SCAN_IN, P2_INSTQUEUE_REG_8__1__SCAN_IN, 
        P2_INSTQUEUE_REG_8__0__SCAN_IN, P2_INSTQUEUE_REG_7__7__SCAN_IN, 
        P2_INSTQUEUE_REG_7__6__SCAN_IN, P2_INSTQUEUE_REG_7__5__SCAN_IN, 
        P2_INSTQUEUE_REG_7__4__SCAN_IN, P2_INSTQUEUE_REG_7__3__SCAN_IN, 
        P2_INSTQUEUE_REG_7__2__SCAN_IN, P2_INSTQUEUE_REG_7__1__SCAN_IN, 
        P2_INSTQUEUE_REG_7__0__SCAN_IN, P2_INSTQUEUE_REG_6__7__SCAN_IN, 
        P2_INSTQUEUE_REG_6__6__SCAN_IN, P2_INSTQUEUE_REG_6__5__SCAN_IN, 
        P2_INSTQUEUE_REG_6__4__SCAN_IN, P2_INSTQUEUE_REG_6__3__SCAN_IN, 
        P2_INSTQUEUE_REG_6__2__SCAN_IN, P2_INSTQUEUE_REG_6__1__SCAN_IN, 
        P2_INSTQUEUE_REG_6__0__SCAN_IN, P2_INSTQUEUE_REG_5__7__SCAN_IN, 
        P2_INSTQUEUE_REG_5__6__SCAN_IN, P2_INSTQUEUE_REG_5__5__SCAN_IN, 
        P2_INSTQUEUE_REG_5__4__SCAN_IN, P2_INSTQUEUE_REG_5__3__SCAN_IN, 
        P2_INSTQUEUE_REG_5__2__SCAN_IN, P2_INSTQUEUE_REG_5__1__SCAN_IN, 
        P2_INSTQUEUE_REG_5__0__SCAN_IN, P2_INSTQUEUE_REG_4__7__SCAN_IN, 
        P2_INSTQUEUE_REG_4__6__SCAN_IN, P2_INSTQUEUE_REG_4__5__SCAN_IN, 
        P2_INSTQUEUE_REG_4__4__SCAN_IN, P2_INSTQUEUE_REG_4__3__SCAN_IN, 
        P2_INSTQUEUE_REG_4__2__SCAN_IN, P2_INSTQUEUE_REG_4__1__SCAN_IN, 
        P2_INSTQUEUE_REG_4__0__SCAN_IN, P2_INSTQUEUE_REG_3__7__SCAN_IN, 
        P2_INSTQUEUE_REG_3__6__SCAN_IN, P2_INSTQUEUE_REG_3__5__SCAN_IN, 
        P2_INSTQUEUE_REG_3__4__SCAN_IN, P2_INSTQUEUE_REG_3__3__SCAN_IN, 
        P2_INSTQUEUE_REG_3__2__SCAN_IN, P2_INSTQUEUE_REG_3__1__SCAN_IN, 
        P2_INSTQUEUE_REG_3__0__SCAN_IN, P2_INSTQUEUE_REG_2__7__SCAN_IN, 
        P2_INSTQUEUE_REG_2__6__SCAN_IN, P2_INSTQUEUE_REG_2__5__SCAN_IN, 
        P2_INSTQUEUE_REG_2__4__SCAN_IN, P2_INSTQUEUE_REG_2__3__SCAN_IN, 
        P2_INSTQUEUE_REG_2__2__SCAN_IN, P2_INSTQUEUE_REG_2__1__SCAN_IN, 
        P2_INSTQUEUE_REG_2__0__SCAN_IN, P2_INSTQUEUE_REG_1__7__SCAN_IN, 
        P2_INSTQUEUE_REG_1__6__SCAN_IN, P2_INSTQUEUE_REG_1__5__SCAN_IN, 
        P2_INSTQUEUE_REG_1__4__SCAN_IN, P2_INSTQUEUE_REG_1__3__SCAN_IN, 
        P2_INSTQUEUE_REG_1__2__SCAN_IN, P2_INSTQUEUE_REG_1__1__SCAN_IN, 
        P2_INSTQUEUE_REG_1__0__SCAN_IN, P2_INSTQUEUE_REG_0__7__SCAN_IN, 
        P2_INSTQUEUE_REG_0__6__SCAN_IN, P2_INSTQUEUE_REG_0__5__SCAN_IN, 
        P2_INSTQUEUE_REG_0__4__SCAN_IN, P2_INSTQUEUE_REG_0__3__SCAN_IN, 
        P2_INSTQUEUE_REG_0__2__SCAN_IN, P2_INSTQUEUE_REG_0__1__SCAN_IN, 
        P2_INSTQUEUE_REG_0__0__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN, 
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN, P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN, P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN, 
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_11__SCAN_IN, P2_INSTADDRPOINTER_REG_12__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_13__SCAN_IN, P2_INSTADDRPOINTER_REG_14__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_15__SCAN_IN, P2_INSTADDRPOINTER_REG_16__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_17__SCAN_IN, P2_INSTADDRPOINTER_REG_18__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_19__SCAN_IN, P2_INSTADDRPOINTER_REG_20__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_21__SCAN_IN, P2_INSTADDRPOINTER_REG_22__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_23__SCAN_IN, P2_INSTADDRPOINTER_REG_24__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_25__SCAN_IN, P2_INSTADDRPOINTER_REG_26__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_27__SCAN_IN, P2_INSTADDRPOINTER_REG_28__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_29__SCAN_IN, P2_INSTADDRPOINTER_REG_30__SCAN_IN, 
        P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN, 
        P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN, 
        P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN, 
        P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN, 
        P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN, 
        P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN, 
        P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN, 
        P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN, 
        P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN, 
        P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN, 
        P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN, 
        P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN, 
        P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN, 
        P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN, 
        P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN, 
        P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN, 
        P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN, 
        P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN, 
        P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN, 
        P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN, 
        P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN, 
        P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN, 
        P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN, 
        P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN, P2_EAX_REG_14__SCAN_IN, 
        P2_EAX_REG_15__SCAN_IN, P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN, 
        P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN, P2_EAX_REG_20__SCAN_IN, 
        P2_EAX_REG_21__SCAN_IN, P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN, 
        P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN, P2_EAX_REG_26__SCAN_IN, 
        P2_EAX_REG_27__SCAN_IN, P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN, 
        P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN, 
        P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN, 
        P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN, 
        P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN, 
        P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN, P2_EBX_REG_12__SCAN_IN, 
        P2_EBX_REG_13__SCAN_IN, P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN, 
        P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN, P2_EBX_REG_18__SCAN_IN, 
        P2_EBX_REG_19__SCAN_IN, P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN, 
        P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN, P2_EBX_REG_24__SCAN_IN, 
        P2_EBX_REG_25__SCAN_IN, P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN, 
        P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN, P2_EBX_REG_30__SCAN_IN, 
        P2_EBX_REG_31__SCAN_IN, P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN, 
        P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN, P2_REIP_REG_4__SCAN_IN, 
        P2_REIP_REG_5__SCAN_IN, P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN, 
        P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN, 
        P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN, 
        P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN, 
        P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN, 
        P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN, 
        P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN, 
        P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN, 
        P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN, 
        P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN, 
        P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN, 
        P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN, 
        P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN, 
        P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN, 
        P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN, 
        P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN, 
        P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN, 
        P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN, 
        P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN, 
        P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN, 
        P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN, P1_BE_N_REG_0__SCAN_IN, 
        P1_ADDRESS_REG_29__SCAN_IN, P1_ADDRESS_REG_28__SCAN_IN, 
        P1_ADDRESS_REG_27__SCAN_IN, P1_ADDRESS_REG_26__SCAN_IN, 
        P1_ADDRESS_REG_25__SCAN_IN, P1_ADDRESS_REG_24__SCAN_IN, 
        P1_ADDRESS_REG_23__SCAN_IN, P1_ADDRESS_REG_22__SCAN_IN, 
        P1_ADDRESS_REG_21__SCAN_IN, P1_ADDRESS_REG_20__SCAN_IN, 
        P1_ADDRESS_REG_19__SCAN_IN, P1_ADDRESS_REG_18__SCAN_IN, 
        P1_ADDRESS_REG_17__SCAN_IN, P1_ADDRESS_REG_16__SCAN_IN, 
        P1_ADDRESS_REG_15__SCAN_IN, P1_ADDRESS_REG_14__SCAN_IN, 
        P1_ADDRESS_REG_13__SCAN_IN, P1_ADDRESS_REG_12__SCAN_IN, 
        P1_ADDRESS_REG_11__SCAN_IN, P1_ADDRESS_REG_10__SCAN_IN, 
        P1_ADDRESS_REG_9__SCAN_IN, P1_ADDRESS_REG_8__SCAN_IN, 
        P1_ADDRESS_REG_7__SCAN_IN, P1_ADDRESS_REG_6__SCAN_IN, 
        P1_ADDRESS_REG_5__SCAN_IN, P1_ADDRESS_REG_4__SCAN_IN, 
        P1_ADDRESS_REG_3__SCAN_IN, P1_ADDRESS_REG_2__SCAN_IN, 
        P1_ADDRESS_REG_1__SCAN_IN, P1_ADDRESS_REG_0__SCAN_IN, 
        P1_STATE_REG_2__SCAN_IN, P1_STATE_REG_1__SCAN_IN, 
        P1_STATE_REG_0__SCAN_IN, P1_DATAWIDTH_REG_0__SCAN_IN, 
        P1_DATAWIDTH_REG_1__SCAN_IN, P1_DATAWIDTH_REG_2__SCAN_IN, 
        P1_DATAWIDTH_REG_3__SCAN_IN, P1_DATAWIDTH_REG_4__SCAN_IN, 
        P1_DATAWIDTH_REG_5__SCAN_IN, P1_DATAWIDTH_REG_6__SCAN_IN, 
        P1_DATAWIDTH_REG_7__SCAN_IN, P1_DATAWIDTH_REG_8__SCAN_IN, 
        P1_DATAWIDTH_REG_9__SCAN_IN, P1_DATAWIDTH_REG_10__SCAN_IN, 
        P1_DATAWIDTH_REG_11__SCAN_IN, P1_DATAWIDTH_REG_12__SCAN_IN, 
        P1_DATAWIDTH_REG_13__SCAN_IN, P1_DATAWIDTH_REG_14__SCAN_IN, 
        P1_DATAWIDTH_REG_15__SCAN_IN, P1_DATAWIDTH_REG_16__SCAN_IN, 
        P1_DATAWIDTH_REG_17__SCAN_IN, P1_DATAWIDTH_REG_18__SCAN_IN, 
        P1_DATAWIDTH_REG_19__SCAN_IN, P1_DATAWIDTH_REG_20__SCAN_IN, 
        P1_DATAWIDTH_REG_21__SCAN_IN, P1_DATAWIDTH_REG_22__SCAN_IN, 
        P1_DATAWIDTH_REG_23__SCAN_IN, P1_DATAWIDTH_REG_24__SCAN_IN, 
        P1_DATAWIDTH_REG_25__SCAN_IN, P1_DATAWIDTH_REG_26__SCAN_IN, 
        P1_DATAWIDTH_REG_27__SCAN_IN, P1_DATAWIDTH_REG_28__SCAN_IN, 
        P1_DATAWIDTH_REG_29__SCAN_IN, P1_DATAWIDTH_REG_30__SCAN_IN, 
        P1_DATAWIDTH_REG_31__SCAN_IN, P1_STATE2_REG_3__SCAN_IN, 
        P1_STATE2_REG_2__SCAN_IN, P1_STATE2_REG_1__SCAN_IN, 
        P1_STATE2_REG_0__SCAN_IN, P1_INSTQUEUE_REG_15__7__SCAN_IN, 
        P1_INSTQUEUE_REG_15__6__SCAN_IN, P1_INSTQUEUE_REG_15__5__SCAN_IN, 
        P1_INSTQUEUE_REG_15__4__SCAN_IN, P1_INSTQUEUE_REG_15__3__SCAN_IN, 
        P1_INSTQUEUE_REG_15__2__SCAN_IN, P1_INSTQUEUE_REG_15__1__SCAN_IN, 
        P1_INSTQUEUE_REG_15__0__SCAN_IN, P1_INSTQUEUE_REG_14__7__SCAN_IN, 
        P1_INSTQUEUE_REG_14__6__SCAN_IN, P1_INSTQUEUE_REG_14__5__SCAN_IN, 
        P1_INSTQUEUE_REG_14__4__SCAN_IN, P1_INSTQUEUE_REG_14__3__SCAN_IN, 
        P1_INSTQUEUE_REG_14__2__SCAN_IN, P1_INSTQUEUE_REG_14__1__SCAN_IN, 
        P1_INSTQUEUE_REG_14__0__SCAN_IN, P1_INSTQUEUE_REG_13__7__SCAN_IN, 
        P1_INSTQUEUE_REG_13__6__SCAN_IN, P1_INSTQUEUE_REG_13__5__SCAN_IN, 
        P1_INSTQUEUE_REG_13__4__SCAN_IN, P1_INSTQUEUE_REG_13__3__SCAN_IN, 
        P1_INSTQUEUE_REG_13__2__SCAN_IN, P1_INSTQUEUE_REG_13__1__SCAN_IN, 
        P1_INSTQUEUE_REG_13__0__SCAN_IN, P1_INSTQUEUE_REG_12__7__SCAN_IN, 
        P1_INSTQUEUE_REG_12__6__SCAN_IN, P1_INSTQUEUE_REG_12__5__SCAN_IN, 
        P1_INSTQUEUE_REG_12__4__SCAN_IN, P1_INSTQUEUE_REG_12__3__SCAN_IN, 
        P1_INSTQUEUE_REG_12__2__SCAN_IN, P1_INSTQUEUE_REG_12__1__SCAN_IN, 
        P1_INSTQUEUE_REG_12__0__SCAN_IN, P1_INSTQUEUE_REG_11__7__SCAN_IN, 
        P1_INSTQUEUE_REG_11__6__SCAN_IN, P1_INSTQUEUE_REG_11__5__SCAN_IN, 
        P1_INSTQUEUE_REG_11__4__SCAN_IN, P1_INSTQUEUE_REG_11__3__SCAN_IN, 
        P1_INSTQUEUE_REG_11__2__SCAN_IN, P1_INSTQUEUE_REG_11__1__SCAN_IN, 
        P1_INSTQUEUE_REG_11__0__SCAN_IN, P1_INSTQUEUE_REG_10__7__SCAN_IN, 
        P1_INSTQUEUE_REG_10__6__SCAN_IN, P1_INSTQUEUE_REG_10__5__SCAN_IN, 
        P1_INSTQUEUE_REG_10__4__SCAN_IN, P1_INSTQUEUE_REG_10__3__SCAN_IN, 
        P1_INSTQUEUE_REG_10__2__SCAN_IN, P1_INSTQUEUE_REG_10__1__SCAN_IN, 
        P1_INSTQUEUE_REG_10__0__SCAN_IN, P1_INSTQUEUE_REG_9__7__SCAN_IN, 
        P1_INSTQUEUE_REG_9__6__SCAN_IN, P1_INSTQUEUE_REG_9__5__SCAN_IN, 
        P1_INSTQUEUE_REG_9__4__SCAN_IN, P1_INSTQUEUE_REG_9__3__SCAN_IN, 
        P1_INSTQUEUE_REG_9__2__SCAN_IN, P1_INSTQUEUE_REG_9__1__SCAN_IN, 
        P1_INSTQUEUE_REG_9__0__SCAN_IN, P1_INSTQUEUE_REG_8__7__SCAN_IN, 
        P1_INSTQUEUE_REG_8__6__SCAN_IN, P1_INSTQUEUE_REG_8__5__SCAN_IN, 
        P1_INSTQUEUE_REG_8__4__SCAN_IN, P1_INSTQUEUE_REG_8__3__SCAN_IN, 
        P1_INSTQUEUE_REG_8__2__SCAN_IN, P1_INSTQUEUE_REG_8__1__SCAN_IN, 
        P1_INSTQUEUE_REG_8__0__SCAN_IN, P1_INSTQUEUE_REG_7__7__SCAN_IN, 
        P1_INSTQUEUE_REG_7__6__SCAN_IN, P1_INSTQUEUE_REG_7__5__SCAN_IN, 
        P1_INSTQUEUE_REG_7__4__SCAN_IN, P1_INSTQUEUE_REG_7__3__SCAN_IN, 
        P1_INSTQUEUE_REG_7__2__SCAN_IN, P1_INSTQUEUE_REG_7__1__SCAN_IN, 
        P1_INSTQUEUE_REG_7__0__SCAN_IN, P1_INSTQUEUE_REG_6__7__SCAN_IN, 
        P1_INSTQUEUE_REG_6__6__SCAN_IN, P1_INSTQUEUE_REG_6__5__SCAN_IN, 
        P1_INSTQUEUE_REG_6__4__SCAN_IN, P1_INSTQUEUE_REG_6__3__SCAN_IN, 
        P1_INSTQUEUE_REG_6__2__SCAN_IN, P1_INSTQUEUE_REG_6__1__SCAN_IN, 
        P1_INSTQUEUE_REG_6__0__SCAN_IN, P1_INSTQUEUE_REG_5__7__SCAN_IN, 
        P1_INSTQUEUE_REG_5__6__SCAN_IN, P1_INSTQUEUE_REG_5__5__SCAN_IN, 
        P1_INSTQUEUE_REG_5__4__SCAN_IN, P1_INSTQUEUE_REG_5__3__SCAN_IN, 
        P1_INSTQUEUE_REG_5__2__SCAN_IN, P1_INSTQUEUE_REG_5__1__SCAN_IN, 
        P1_INSTQUEUE_REG_5__0__SCAN_IN, P1_INSTQUEUE_REG_4__7__SCAN_IN, 
        P1_INSTQUEUE_REG_4__6__SCAN_IN, P1_INSTQUEUE_REG_4__5__SCAN_IN, 
        P1_INSTQUEUE_REG_4__4__SCAN_IN, P1_INSTQUEUE_REG_4__3__SCAN_IN, 
        P1_INSTQUEUE_REG_4__2__SCAN_IN, P1_INSTQUEUE_REG_4__1__SCAN_IN, 
        keyinput0, keyinput1, keyinput2, keyinput3, keyinput4, keyinput5, 
        keyinput6, keyinput7, keyinput8, keyinput9, keyinput10, keyinput11, 
        keyinput12, keyinput13, keyinput14, keyinput15, keyinput16, keyinput17, 
        keyinput18, keyinput19, keyinput20, keyinput21, keyinput22, keyinput23, 
        keyinput24, keyinput25, keyinput26, keyinput27, keyinput28, keyinput29, 
        keyinput30, keyinput31, keyinput32, keyinput33, keyinput34, keyinput35, 
        keyinput36, keyinput37, keyinput38, keyinput39, keyinput40, keyinput41, 
        keyinput42, keyinput43, keyinput44, keyinput45, keyinput46, keyinput47, 
        keyinput48, keyinput49, keyinput50, keyinput51, keyinput52, keyinput53, 
        keyinput54, keyinput55, keyinput56, keyinput57, keyinput58, keyinput59, 
        keyinput60, keyinput61, keyinput62, keyinput63, keyinput64, keyinput65, 
        keyinput66, keyinput67, keyinput68, keyinput69, keyinput70, keyinput71, 
        keyinput72, keyinput73, keyinput74, keyinput75, keyinput76, keyinput77, 
        keyinput78, keyinput79, keyinput80, keyinput81, keyinput82, keyinput83, 
        keyinput84, keyinput85, keyinput86, keyinput87, keyinput88, keyinput89, 
        keyinput90, keyinput91, keyinput92, keyinput93, keyinput94, keyinput95, 
        keyinput96, keyinput97, keyinput98, keyinput99, keyinput100, 
        keyinput101, keyinput102, keyinput103, keyinput104, keyinput105, 
        keyinput106, keyinput107, keyinput108, keyinput109, keyinput110, 
        keyinput111, keyinput112, keyinput113, keyinput114, keyinput115, 
        keyinput116, keyinput117, keyinput118, keyinput119, keyinput120, 
        keyinput121, keyinput122, keyinput123, keyinput124, keyinput125, 
        keyinput126, keyinput127, keyinput128, keyinput129, keyinput130, 
        keyinput131, keyinput132, keyinput133, keyinput134, keyinput135, 
        keyinput136, keyinput137, keyinput138, keyinput139, keyinput140, 
        keyinput141, keyinput142, keyinput143, keyinput144, keyinput145, 
        keyinput146, keyinput147, keyinput148, keyinput149, keyinput150, 
        keyinput151, keyinput152, keyinput153, keyinput154, keyinput155, 
        keyinput156, keyinput157, keyinput158, keyinput159, keyinput160, 
        keyinput161, keyinput162, keyinput163, keyinput164, keyinput165, 
        keyinput166, keyinput167, keyinput168, keyinput169, keyinput170, 
        keyinput171, keyinput172, keyinput173, keyinput174, keyinput175, 
        keyinput176, keyinput177, keyinput178, keyinput179, keyinput180, 
        keyinput181, keyinput182, keyinput183, keyinput184, keyinput185, 
        keyinput186, keyinput187, keyinput188, keyinput189, keyinput190, 
        keyinput191, keyinput192, keyinput193, keyinput194, keyinput195, 
        keyinput196, keyinput197, keyinput198, keyinput199, keyinput200, 
        keyinput201, keyinput202, keyinput203, keyinput204, keyinput205, 
        keyinput206, keyinput207, keyinput208, keyinput209, keyinput210, 
        keyinput211, keyinput212, keyinput213, keyinput214, keyinput215, 
        keyinput216, keyinput217, keyinput218, keyinput219, keyinput220, 
        keyinput221, keyinput222, keyinput223, keyinput224, keyinput225, 
        keyinput226, keyinput227, keyinput228, keyinput229, keyinput230, 
        keyinput231, keyinput232, keyinput233, keyinput234, keyinput235, 
        keyinput236, keyinput237, keyinput238, keyinput239, keyinput240, 
        keyinput241, keyinput242, keyinput243, keyinput244, keyinput245, 
        keyinput246, keyinput247, keyinput248, keyinput249, keyinput250, 
        keyinput251, keyinput252, keyinput253, keyinput254, keyinput255, U355, 
        U356, U357, U358, U359, U360, U361, U362, U363, U364, U366, U367, U368, 
        U369, U370, U371, U372, U373, U374, U375, U347, U348, U349, U350, U351, 
        U352, U353, U354, U365, U376, U247, U246, U245, U244, U243, U242, U241, 
        U240, U239, U238, U237, U236, U235, U234, U233, U232, U231, U230, U229, 
        U228, U227, U226, U225, U224, U223, U222, U221, U220, U219, U218, U217, 
        U216, U251, U252, U253, U254, U255, U256, U257, U258, U259, U260, U261, 
        U262, U263, U264, U265, U266, U267, U268, U269, U270, U271, U272, U273, 
        U274, U275, U276, U277, U278, U279, U280, U281, U282, U212, U215, U213, 
        U214, P3_U3274, P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, 
        P3_U3059, P3_U3058, P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, 
        P3_U3052, P3_U3051, P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, 
        P3_U3045, P3_U3044, P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, 
        P3_U3038, P3_U3037, P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, 
        P3_U3031, P3_U3030, P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, 
        P3_U3026, P3_U3025, P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, 
        P3_U3019, P3_U3018, P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, 
        P3_U3012, P3_U3011, P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, 
        P3_U3005, P3_U3004, P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, 
        P3_U3282, P3_U2998, P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, 
        P3_U2992, P3_U2991, P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, 
        P3_U2985, P3_U2984, P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, 
        P3_U2978, P3_U2977, P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, 
        P3_U2971, P3_U2970, P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, 
        P3_U2964, P3_U2963, P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, 
        P3_U2957, P3_U2956, P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, 
        P3_U2950, P3_U2949, P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, 
        P3_U2943, P3_U2942, P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, 
        P3_U2936, P3_U2935, P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, 
        P3_U2929, P3_U2928, P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, 
        P3_U2922, P3_U2921, P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, 
        P3_U2915, P3_U2914, P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, 
        P3_U2908, P3_U2907, P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, 
        P3_U2901, P3_U2900, P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, 
        P3_U2894, P3_U2893, P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, 
        P3_U2887, P3_U2886, P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, 
        P3_U2880, P3_U2879, P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, 
        P3_U2873, P3_U2872, P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, 
        P3_U3285, P3_U3288, P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, 
        P3_U2864, P3_U2863, P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, 
        P3_U2857, P3_U2856, P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, 
        P3_U2850, P3_U2849, P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, 
        P3_U2843, P3_U2842, P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, 
        P3_U2836, P3_U2835, P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, 
        P3_U2829, P3_U2828, P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, 
        P3_U2822, P3_U2821, P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, 
        P3_U2815, P3_U2814, P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, 
        P3_U2808, P3_U2807, P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, 
        P3_U2801, P3_U2800, P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, 
        P3_U2794, P3_U2793, P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, 
        P3_U2787, P3_U2786, P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, 
        P3_U2780, P3_U2779, P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, 
        P3_U2773, P3_U2772, P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, 
        P3_U2766, P3_U2765, P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, 
        P3_U2759, P3_U2758, P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, 
        P3_U2752, P3_U2751, P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, 
        P3_U2745, P3_U2744, P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, 
        P3_U2738, P3_U2737, P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, 
        P3_U2731, P3_U2730, P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, 
        P3_U2724, P3_U2723, P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, 
        P3_U2717, P3_U2716, P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, 
        P3_U2710, P3_U2709, P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, 
        P3_U2703, P3_U2702, P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, 
        P3_U2696, P3_U2695, P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, 
        P3_U2689, P3_U2688, P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, 
        P3_U2682, P3_U2681, P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, 
        P3_U2675, P3_U2674, P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, 
        P3_U2668, P3_U2667, P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, 
        P3_U2661, P3_U2660, P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, 
        P3_U2654, P3_U2653, P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, 
        P3_U2647, P3_U2646, P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, 
        P3_U2640, P3_U2639, P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, 
        P3_U3295, P3_U2636, P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, 
        P3_U3298, P3_U3299, P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, 
        P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, 
        P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, 
        P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, 
        P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, 
        P2_U3212, P2_U3211, P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, 
        P2_U3207, P2_U3206, P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, 
        P2_U3200, P2_U3199, P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, 
        P2_U3193, P2_U3192, P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, 
        P2_U3186, P2_U3185, P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, 
        P2_U3179, P2_U3593, P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, 
        P2_U3173, P2_U3172, P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, 
        P2_U3166, P2_U3165, P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, 
        P2_U3159, P2_U3158, P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, 
        P2_U3152, P2_U3151, P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, 
        P2_U3145, P2_U3144, P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, 
        P2_U3138, P2_U3137, P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, 
        P2_U3131, P2_U3130, P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, 
        P2_U3124, P2_U3123, P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, 
        P2_U3117, P2_U3116, P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, 
        P2_U3110, P2_U3109, P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, 
        P2_U3103, P2_U3102, P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, 
        P2_U3096, P2_U3095, P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, 
        P2_U3089, P2_U3088, P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, 
        P2_U3082, P2_U3081, P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, 
        P2_U3075, P2_U3074, P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, 
        P2_U3068, P2_U3067, P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, 
        P2_U3061, P2_U3060, P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, 
        P2_U3054, P2_U3053, P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, 
        P2_U3595, P2_U3596, P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, 
        P2_U3603, P2_U3604, P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, 
        P2_U3042, P2_U3041, P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, 
        P2_U3035, P2_U3034, P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, 
        P2_U3028, P2_U3027, P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, 
        P2_U3021, P2_U3020, P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, 
        P2_U3014, P2_U3013, P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, 
        P2_U3007, P2_U3006, P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, 
        P2_U3000, P2_U2999, P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, 
        P2_U2993, P2_U2992, P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, 
        P2_U2986, P2_U2985, P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, 
        P2_U2979, P2_U2978, P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, 
        P2_U2972, P2_U2971, P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, 
        P2_U2965, P2_U2964, P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, 
        P2_U2958, P2_U2957, P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, 
        P2_U2951, P2_U2950, P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, 
        P2_U2944, P2_U2943, P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, 
        P2_U2937, P2_U2936, P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, 
        P2_U2930, P2_U2929, P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, 
        P2_U2923, P2_U2922, P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, 
        P2_U2916, P2_U2915, P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, 
        P2_U2909, P2_U2908, P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, 
        P2_U2902, P2_U2901, P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, 
        P2_U2895, P2_U2894, P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, 
        P2_U2888, P2_U2887, P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, 
        P2_U2881, P2_U2880, P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, 
        P2_U2874, P2_U2873, P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, 
        P2_U2867, P2_U2866, P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, 
        P2_U2860, P2_U2859, P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, 
        P2_U2853, P2_U2852, P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, 
        P2_U2846, P2_U2845, P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, 
        P2_U2839, P2_U2838, P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, 
        P2_U2832, P2_U2831, P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, 
        P2_U2825, P2_U2824, P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, 
        P2_U2819, P2_U3609, P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, 
        P2_U2815, P2_U3612, P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, 
        P1_U3226, P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, 
        P1_U3219, P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, 
        P1_U3212, P1_U3211, P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, 
        P1_U3205, P1_U3204, P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, 
        P1_U3198, P1_U3197, P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, 
        P1_U3193, P1_U3192, P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, 
        P1_U3186, P1_U3185, P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, 
        P1_U3179, P1_U3178, P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, 
        P1_U3172, P1_U3171, P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, 
        P1_U3165, P1_U3164, P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, 
        P1_U3159, P1_U3158, P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, 
        P1_U3152, P1_U3151, P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, 
        P1_U3145, P1_U3144, P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, 
        P1_U3138, P1_U3137, P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, 
        P1_U3131, P1_U3130, P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, 
        P1_U3124, P1_U3123, P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, 
        P1_U3117, P1_U3116, P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, 
        P1_U3110, P1_U3109, P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, 
        P1_U3103, P1_U3102, P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, 
        P1_U3096, P1_U3095, P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, 
        P1_U3089, P1_U3088, P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, 
        P1_U3082, P1_U3081, P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, 
        P1_U3075, P1_U3074, P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, 
        P1_U3068, P1_U3067, P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, 
        P1_U3061, P1_U3060, P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, 
        P1_U3054, P1_U3053, P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, 
        P1_U3047, P1_U3046, P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, 
        P1_U3040, P1_U3039, P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, 
        P1_U3033, P1_U3468, P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, 
        P1_U3475, P1_U3476, P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, 
        P1_U3028, P1_U3027, P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, 
        P1_U3021, P1_U3020, P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, 
        P1_U3014, P1_U3013, P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, 
        P1_U3007, P1_U3006, P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, 
        P1_U3000, P1_U2999, P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, 
        P1_U2993, P1_U2992, P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, 
        P1_U2986, P1_U2985, P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, 
        P1_U2979, P1_U2978, P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, 
        P1_U2972, P1_U2971, P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, 
        P1_U2965, P1_U2964, P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, 
        P1_U2958, P1_U2957, P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, 
        P1_U2951, P1_U2950, P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, 
        P1_U2944, P1_U2943, P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, 
        P1_U2937, P1_U2936, P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, 
        P1_U2930, P1_U2929, P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, 
        P1_U2923, P1_U2922, P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, 
        P1_U2916, P1_U2915, P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, 
        P1_U2909, P1_U2908, P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, 
        P1_U2902, P1_U2901, P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, 
        P1_U2895, P1_U2894, P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, 
        P1_U2888, P1_U2887, P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, 
        P1_U2881, P1_U2880, P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, 
        P1_U2874, P1_U2873, P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, 
        P1_U2867, P1_U2866, P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, 
        P1_U2860, P1_U2859, P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, 
        P1_U2853, P1_U2852, P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, 
        P1_U2846, P1_U2845, P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, 
        P1_U2839, P1_U2838, P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, 
        P1_U2832, P1_U2831, P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, 
        P1_U2825, P1_U2824, P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, 
        P1_U2818, P1_U2817, P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, 
        P1_U2811, P1_U2810, P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, 
        P1_U3483, P1_U2806, P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, 
        P1_U2803, P1_U2802, P1_U3487, P1_U2801 );
  input P1_MEMORYFETCH_REG_SCAN_IN, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_,
         DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_,
         DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_,
         DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_,
         DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_,
         DATAI_2_, DATAI_1_, DATAI_0_, HOLD, NA, BS16, READY1, READY2,
         P1_READREQUEST_REG_SCAN_IN, P1_ADS_N_REG_SCAN_IN,
         P1_CODEFETCH_REG_SCAN_IN, P1_M_IO_N_REG_SCAN_IN, P1_D_C_N_REG_SCAN_IN,
         P1_REQUESTPENDING_REG_SCAN_IN, P1_STATEBS16_REG_SCAN_IN,
         P1_MORE_REG_SCAN_IN, P1_FLUSH_REG_SCAN_IN, P1_W_R_N_REG_SCAN_IN,
         P1_BYTEENABLE_REG_0__SCAN_IN, P1_BYTEENABLE_REG_1__SCAN_IN,
         P1_BYTEENABLE_REG_2__SCAN_IN, P1_BYTEENABLE_REG_3__SCAN_IN,
         P1_REIP_REG_31__SCAN_IN, P1_REIP_REG_30__SCAN_IN,
         P1_REIP_REG_29__SCAN_IN, P1_REIP_REG_28__SCAN_IN,
         P1_REIP_REG_27__SCAN_IN, P1_REIP_REG_26__SCAN_IN,
         P1_REIP_REG_25__SCAN_IN, P1_REIP_REG_24__SCAN_IN,
         P1_REIP_REG_23__SCAN_IN, P1_REIP_REG_22__SCAN_IN,
         P1_REIP_REG_21__SCAN_IN, P1_REIP_REG_20__SCAN_IN,
         P1_REIP_REG_19__SCAN_IN, P1_REIP_REG_18__SCAN_IN,
         P1_REIP_REG_17__SCAN_IN, P1_REIP_REG_16__SCAN_IN,
         P1_REIP_REG_15__SCAN_IN, P1_REIP_REG_14__SCAN_IN,
         P1_REIP_REG_13__SCAN_IN, P1_REIP_REG_12__SCAN_IN,
         P1_REIP_REG_11__SCAN_IN, P1_REIP_REG_10__SCAN_IN,
         P1_REIP_REG_9__SCAN_IN, P1_REIP_REG_8__SCAN_IN,
         P1_REIP_REG_7__SCAN_IN, P1_REIP_REG_6__SCAN_IN,
         P1_REIP_REG_5__SCAN_IN, P1_REIP_REG_4__SCAN_IN,
         P1_REIP_REG_3__SCAN_IN, P1_REIP_REG_2__SCAN_IN,
         P1_REIP_REG_1__SCAN_IN, P1_REIP_REG_0__SCAN_IN,
         P1_EBX_REG_31__SCAN_IN, P1_EBX_REG_30__SCAN_IN,
         P1_EBX_REG_29__SCAN_IN, P1_EBX_REG_28__SCAN_IN,
         P1_EBX_REG_27__SCAN_IN, P1_EBX_REG_26__SCAN_IN,
         P1_EBX_REG_25__SCAN_IN, P1_EBX_REG_24__SCAN_IN,
         P1_EBX_REG_23__SCAN_IN, P1_EBX_REG_22__SCAN_IN,
         P1_EBX_REG_21__SCAN_IN, P1_EBX_REG_20__SCAN_IN,
         P1_EBX_REG_19__SCAN_IN, P1_EBX_REG_18__SCAN_IN,
         P1_EBX_REG_17__SCAN_IN, P1_EBX_REG_16__SCAN_IN,
         P1_EBX_REG_15__SCAN_IN, P1_EBX_REG_14__SCAN_IN,
         P1_EBX_REG_13__SCAN_IN, P1_EBX_REG_12__SCAN_IN,
         P1_EBX_REG_11__SCAN_IN, P1_EBX_REG_10__SCAN_IN, P1_EBX_REG_9__SCAN_IN,
         P1_EBX_REG_8__SCAN_IN, P1_EBX_REG_7__SCAN_IN, P1_EBX_REG_6__SCAN_IN,
         P1_EBX_REG_5__SCAN_IN, P1_EBX_REG_4__SCAN_IN, P1_EBX_REG_3__SCAN_IN,
         P1_EBX_REG_2__SCAN_IN, P1_EBX_REG_1__SCAN_IN, P1_EBX_REG_0__SCAN_IN,
         P1_EAX_REG_31__SCAN_IN, P1_EAX_REG_30__SCAN_IN,
         P1_EAX_REG_29__SCAN_IN, P1_EAX_REG_28__SCAN_IN,
         P1_EAX_REG_27__SCAN_IN, P1_EAX_REG_26__SCAN_IN,
         P1_EAX_REG_25__SCAN_IN, P1_EAX_REG_24__SCAN_IN,
         P1_EAX_REG_23__SCAN_IN, P1_EAX_REG_22__SCAN_IN,
         P1_EAX_REG_21__SCAN_IN, P1_EAX_REG_20__SCAN_IN,
         P1_EAX_REG_19__SCAN_IN, P1_EAX_REG_18__SCAN_IN,
         P1_EAX_REG_17__SCAN_IN, P1_EAX_REG_16__SCAN_IN,
         P1_EAX_REG_15__SCAN_IN, P1_EAX_REG_14__SCAN_IN,
         P1_EAX_REG_13__SCAN_IN, P1_EAX_REG_12__SCAN_IN,
         P1_EAX_REG_11__SCAN_IN, P1_EAX_REG_10__SCAN_IN, P1_EAX_REG_9__SCAN_IN,
         P1_EAX_REG_8__SCAN_IN, P1_EAX_REG_7__SCAN_IN, P1_EAX_REG_6__SCAN_IN,
         P1_EAX_REG_5__SCAN_IN, P1_EAX_REG_4__SCAN_IN, P1_EAX_REG_3__SCAN_IN,
         P1_EAX_REG_2__SCAN_IN, P1_EAX_REG_1__SCAN_IN, P1_EAX_REG_0__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_UWORD_REG_0__SCAN_IN, P1_UWORD_REG_1__SCAN_IN,
         P1_UWORD_REG_2__SCAN_IN, P1_UWORD_REG_3__SCAN_IN,
         P1_UWORD_REG_4__SCAN_IN, P1_UWORD_REG_5__SCAN_IN,
         P1_UWORD_REG_6__SCAN_IN, P1_UWORD_REG_7__SCAN_IN,
         P1_UWORD_REG_8__SCAN_IN, P1_UWORD_REG_9__SCAN_IN,
         P1_UWORD_REG_10__SCAN_IN, P1_UWORD_REG_11__SCAN_IN,
         P1_UWORD_REG_12__SCAN_IN, P1_UWORD_REG_13__SCAN_IN,
         P1_UWORD_REG_14__SCAN_IN, P1_LWORD_REG_0__SCAN_IN,
         P1_LWORD_REG_1__SCAN_IN, P1_LWORD_REG_2__SCAN_IN,
         P1_LWORD_REG_3__SCAN_IN, P1_LWORD_REG_4__SCAN_IN,
         P1_LWORD_REG_5__SCAN_IN, P1_LWORD_REG_6__SCAN_IN,
         P1_LWORD_REG_7__SCAN_IN, P1_LWORD_REG_8__SCAN_IN,
         P1_LWORD_REG_9__SCAN_IN, P1_LWORD_REG_10__SCAN_IN,
         P1_LWORD_REG_11__SCAN_IN, P1_LWORD_REG_12__SCAN_IN,
         P1_LWORD_REG_13__SCAN_IN, P1_LWORD_REG_14__SCAN_IN,
         P1_LWORD_REG_15__SCAN_IN, P1_PHYADDRPOINTER_REG_31__SCAN_IN,
         P1_PHYADDRPOINTER_REG_30__SCAN_IN, P1_PHYADDRPOINTER_REG_29__SCAN_IN,
         P1_PHYADDRPOINTER_REG_28__SCAN_IN, P1_PHYADDRPOINTER_REG_27__SCAN_IN,
         P1_PHYADDRPOINTER_REG_26__SCAN_IN, P1_PHYADDRPOINTER_REG_25__SCAN_IN,
         P1_PHYADDRPOINTER_REG_24__SCAN_IN, P1_PHYADDRPOINTER_REG_23__SCAN_IN,
         P1_PHYADDRPOINTER_REG_22__SCAN_IN, P1_PHYADDRPOINTER_REG_21__SCAN_IN,
         P1_PHYADDRPOINTER_REG_20__SCAN_IN, P1_PHYADDRPOINTER_REG_19__SCAN_IN,
         P1_PHYADDRPOINTER_REG_18__SCAN_IN, P1_PHYADDRPOINTER_REG_17__SCAN_IN,
         P1_PHYADDRPOINTER_REG_16__SCAN_IN, P1_PHYADDRPOINTER_REG_15__SCAN_IN,
         P1_PHYADDRPOINTER_REG_14__SCAN_IN, P1_PHYADDRPOINTER_REG_13__SCAN_IN,
         P1_PHYADDRPOINTER_REG_12__SCAN_IN, P1_PHYADDRPOINTER_REG_11__SCAN_IN,
         P1_PHYADDRPOINTER_REG_10__SCAN_IN, P1_PHYADDRPOINTER_REG_9__SCAN_IN,
         P1_PHYADDRPOINTER_REG_8__SCAN_IN, P1_PHYADDRPOINTER_REG_7__SCAN_IN,
         P1_PHYADDRPOINTER_REG_6__SCAN_IN, P1_PHYADDRPOINTER_REG_5__SCAN_IN,
         P1_PHYADDRPOINTER_REG_4__SCAN_IN, P1_PHYADDRPOINTER_REG_3__SCAN_IN,
         P1_PHYADDRPOINTER_REG_2__SCAN_IN, P1_PHYADDRPOINTER_REG_1__SCAN_IN,
         P1_PHYADDRPOINTER_REG_0__SCAN_IN, P1_INSTADDRPOINTER_REG_31__SCAN_IN,
         P1_INSTADDRPOINTER_REG_30__SCAN_IN,
         P1_INSTADDRPOINTER_REG_29__SCAN_IN,
         P1_INSTADDRPOINTER_REG_28__SCAN_IN,
         P1_INSTADDRPOINTER_REG_27__SCAN_IN,
         P1_INSTADDRPOINTER_REG_26__SCAN_IN,
         P1_INSTADDRPOINTER_REG_25__SCAN_IN,
         P1_INSTADDRPOINTER_REG_24__SCAN_IN,
         P1_INSTADDRPOINTER_REG_23__SCAN_IN,
         P1_INSTADDRPOINTER_REG_22__SCAN_IN,
         P1_INSTADDRPOINTER_REG_21__SCAN_IN,
         P1_INSTADDRPOINTER_REG_20__SCAN_IN,
         P1_INSTADDRPOINTER_REG_19__SCAN_IN,
         P1_INSTADDRPOINTER_REG_18__SCAN_IN,
         P1_INSTADDRPOINTER_REG_17__SCAN_IN,
         P1_INSTADDRPOINTER_REG_16__SCAN_IN,
         P1_INSTADDRPOINTER_REG_15__SCAN_IN,
         P1_INSTADDRPOINTER_REG_14__SCAN_IN,
         P1_INSTADDRPOINTER_REG_13__SCAN_IN,
         P1_INSTADDRPOINTER_REG_12__SCAN_IN,
         P1_INSTADDRPOINTER_REG_11__SCAN_IN,
         P1_INSTADDRPOINTER_REG_10__SCAN_IN, P1_INSTADDRPOINTER_REG_9__SCAN_IN,
         P1_INSTADDRPOINTER_REG_8__SCAN_IN, P1_INSTADDRPOINTER_REG_7__SCAN_IN,
         P1_INSTADDRPOINTER_REG_6__SCAN_IN, P1_INSTADDRPOINTER_REG_5__SCAN_IN,
         P1_INSTADDRPOINTER_REG_4__SCAN_IN, P1_INSTADDRPOINTER_REG_3__SCAN_IN,
         P1_INSTADDRPOINTER_REG_2__SCAN_IN, P1_INSTADDRPOINTER_REG_1__SCAN_IN,
         P1_INSTADDRPOINTER_REG_0__SCAN_IN, P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN, P1_INSTQUEUE_REG_0__0__SCAN_IN,
         P1_INSTQUEUE_REG_0__1__SCAN_IN, P1_INSTQUEUE_REG_0__2__SCAN_IN,
         P1_INSTQUEUE_REG_0__3__SCAN_IN, P1_INSTQUEUE_REG_0__4__SCAN_IN,
         P1_INSTQUEUE_REG_0__5__SCAN_IN, P1_INSTQUEUE_REG_0__6__SCAN_IN,
         P1_INSTQUEUE_REG_0__7__SCAN_IN, P1_INSTQUEUE_REG_1__0__SCAN_IN,
         P1_INSTQUEUE_REG_1__1__SCAN_IN, P1_INSTQUEUE_REG_1__2__SCAN_IN,
         P1_INSTQUEUE_REG_1__3__SCAN_IN, P1_INSTQUEUE_REG_1__4__SCAN_IN,
         P1_INSTQUEUE_REG_1__5__SCAN_IN, P1_INSTQUEUE_REG_1__6__SCAN_IN,
         P1_INSTQUEUE_REG_1__7__SCAN_IN, P1_INSTQUEUE_REG_2__0__SCAN_IN,
         P1_INSTQUEUE_REG_2__1__SCAN_IN, P1_INSTQUEUE_REG_2__2__SCAN_IN,
         P1_INSTQUEUE_REG_2__3__SCAN_IN, P1_INSTQUEUE_REG_2__4__SCAN_IN,
         P1_INSTQUEUE_REG_2__5__SCAN_IN, P1_INSTQUEUE_REG_2__6__SCAN_IN,
         P1_INSTQUEUE_REG_2__7__SCAN_IN, P1_INSTQUEUE_REG_3__0__SCAN_IN,
         P1_INSTQUEUE_REG_3__1__SCAN_IN, P1_INSTQUEUE_REG_3__2__SCAN_IN,
         P1_INSTQUEUE_REG_3__3__SCAN_IN, P1_INSTQUEUE_REG_3__4__SCAN_IN,
         P1_INSTQUEUE_REG_3__5__SCAN_IN, P1_INSTQUEUE_REG_3__6__SCAN_IN,
         P1_INSTQUEUE_REG_3__7__SCAN_IN, P1_INSTQUEUE_REG_4__0__SCAN_IN,
         BUF1_REG_0__SCAN_IN, BUF1_REG_1__SCAN_IN, BUF1_REG_2__SCAN_IN,
         BUF1_REG_3__SCAN_IN, BUF1_REG_4__SCAN_IN, BUF1_REG_5__SCAN_IN,
         BUF1_REG_6__SCAN_IN, BUF1_REG_7__SCAN_IN, BUF1_REG_8__SCAN_IN,
         BUF1_REG_9__SCAN_IN, BUF1_REG_10__SCAN_IN, BUF1_REG_11__SCAN_IN,
         BUF1_REG_12__SCAN_IN, BUF1_REG_13__SCAN_IN, BUF1_REG_14__SCAN_IN,
         BUF1_REG_15__SCAN_IN, BUF1_REG_16__SCAN_IN, BUF1_REG_17__SCAN_IN,
         BUF1_REG_18__SCAN_IN, BUF1_REG_19__SCAN_IN, BUF1_REG_20__SCAN_IN,
         BUF1_REG_21__SCAN_IN, BUF1_REG_22__SCAN_IN, BUF1_REG_23__SCAN_IN,
         BUF1_REG_24__SCAN_IN, BUF1_REG_25__SCAN_IN, BUF1_REG_26__SCAN_IN,
         BUF1_REG_27__SCAN_IN, BUF1_REG_28__SCAN_IN, BUF1_REG_29__SCAN_IN,
         BUF1_REG_30__SCAN_IN, BUF1_REG_31__SCAN_IN, BUF2_REG_0__SCAN_IN,
         BUF2_REG_1__SCAN_IN, BUF2_REG_2__SCAN_IN, BUF2_REG_3__SCAN_IN,
         BUF2_REG_4__SCAN_IN, BUF2_REG_5__SCAN_IN, BUF2_REG_6__SCAN_IN,
         BUF2_REG_7__SCAN_IN, BUF2_REG_8__SCAN_IN, BUF2_REG_9__SCAN_IN,
         BUF2_REG_10__SCAN_IN, BUF2_REG_11__SCAN_IN, BUF2_REG_12__SCAN_IN,
         BUF2_REG_13__SCAN_IN, BUF2_REG_14__SCAN_IN, BUF2_REG_15__SCAN_IN,
         BUF2_REG_16__SCAN_IN, BUF2_REG_17__SCAN_IN, BUF2_REG_18__SCAN_IN,
         BUF2_REG_19__SCAN_IN, BUF2_REG_20__SCAN_IN, BUF2_REG_21__SCAN_IN,
         BUF2_REG_22__SCAN_IN, BUF2_REG_23__SCAN_IN, BUF2_REG_24__SCAN_IN,
         BUF2_REG_25__SCAN_IN, BUF2_REG_26__SCAN_IN, BUF2_REG_27__SCAN_IN,
         BUF2_REG_28__SCAN_IN, BUF2_REG_29__SCAN_IN, BUF2_REG_30__SCAN_IN,
         BUF2_REG_31__SCAN_IN, READY12_REG_SCAN_IN, READY21_REG_SCAN_IN,
         READY22_REG_SCAN_IN, READY11_REG_SCAN_IN, P3_BE_N_REG_3__SCAN_IN,
         P3_BE_N_REG_2__SCAN_IN, P3_BE_N_REG_1__SCAN_IN,
         P3_BE_N_REG_0__SCAN_IN, P3_ADDRESS_REG_29__SCAN_IN,
         P3_ADDRESS_REG_28__SCAN_IN, P3_ADDRESS_REG_27__SCAN_IN,
         P3_ADDRESS_REG_26__SCAN_IN, P3_ADDRESS_REG_25__SCAN_IN,
         P3_ADDRESS_REG_24__SCAN_IN, P3_ADDRESS_REG_23__SCAN_IN,
         P3_ADDRESS_REG_22__SCAN_IN, P3_ADDRESS_REG_21__SCAN_IN,
         P3_ADDRESS_REG_20__SCAN_IN, P3_ADDRESS_REG_19__SCAN_IN,
         P3_ADDRESS_REG_18__SCAN_IN, P3_ADDRESS_REG_17__SCAN_IN,
         P3_ADDRESS_REG_16__SCAN_IN, P3_ADDRESS_REG_15__SCAN_IN,
         P3_ADDRESS_REG_14__SCAN_IN, P3_ADDRESS_REG_13__SCAN_IN,
         P3_ADDRESS_REG_12__SCAN_IN, P3_ADDRESS_REG_11__SCAN_IN,
         P3_ADDRESS_REG_10__SCAN_IN, P3_ADDRESS_REG_9__SCAN_IN,
         P3_ADDRESS_REG_8__SCAN_IN, P3_ADDRESS_REG_7__SCAN_IN,
         P3_ADDRESS_REG_6__SCAN_IN, P3_ADDRESS_REG_5__SCAN_IN,
         P3_ADDRESS_REG_4__SCAN_IN, P3_ADDRESS_REG_3__SCAN_IN,
         P3_ADDRESS_REG_2__SCAN_IN, P3_ADDRESS_REG_1__SCAN_IN,
         P3_ADDRESS_REG_0__SCAN_IN, P3_STATE_REG_2__SCAN_IN,
         P3_STATE_REG_1__SCAN_IN, P3_STATE_REG_0__SCAN_IN,
         P3_DATAWIDTH_REG_0__SCAN_IN, P3_DATAWIDTH_REG_1__SCAN_IN,
         P3_DATAWIDTH_REG_2__SCAN_IN, P3_DATAWIDTH_REG_3__SCAN_IN,
         P3_DATAWIDTH_REG_4__SCAN_IN, P3_DATAWIDTH_REG_5__SCAN_IN,
         P3_DATAWIDTH_REG_6__SCAN_IN, P3_DATAWIDTH_REG_7__SCAN_IN,
         P3_DATAWIDTH_REG_8__SCAN_IN, P3_DATAWIDTH_REG_9__SCAN_IN,
         P3_DATAWIDTH_REG_10__SCAN_IN, P3_DATAWIDTH_REG_11__SCAN_IN,
         P3_DATAWIDTH_REG_12__SCAN_IN, P3_DATAWIDTH_REG_13__SCAN_IN,
         P3_DATAWIDTH_REG_14__SCAN_IN, P3_DATAWIDTH_REG_15__SCAN_IN,
         P3_DATAWIDTH_REG_16__SCAN_IN, P3_DATAWIDTH_REG_17__SCAN_IN,
         P3_DATAWIDTH_REG_18__SCAN_IN, P3_DATAWIDTH_REG_19__SCAN_IN,
         P3_DATAWIDTH_REG_20__SCAN_IN, P3_DATAWIDTH_REG_21__SCAN_IN,
         P3_DATAWIDTH_REG_22__SCAN_IN, P3_DATAWIDTH_REG_23__SCAN_IN,
         P3_DATAWIDTH_REG_24__SCAN_IN, P3_DATAWIDTH_REG_25__SCAN_IN,
         P3_DATAWIDTH_REG_26__SCAN_IN, P3_DATAWIDTH_REG_27__SCAN_IN,
         P3_DATAWIDTH_REG_28__SCAN_IN, P3_DATAWIDTH_REG_29__SCAN_IN,
         P3_DATAWIDTH_REG_30__SCAN_IN, P3_DATAWIDTH_REG_31__SCAN_IN,
         P3_STATE2_REG_3__SCAN_IN, P3_STATE2_REG_2__SCAN_IN,
         P3_STATE2_REG_1__SCAN_IN, P3_STATE2_REG_0__SCAN_IN,
         P3_INSTQUEUE_REG_15__7__SCAN_IN, P3_INSTQUEUE_REG_15__6__SCAN_IN,
         P3_INSTQUEUE_REG_15__5__SCAN_IN, P3_INSTQUEUE_REG_15__4__SCAN_IN,
         P3_INSTQUEUE_REG_15__3__SCAN_IN, P3_INSTQUEUE_REG_15__2__SCAN_IN,
         P3_INSTQUEUE_REG_15__1__SCAN_IN, P3_INSTQUEUE_REG_15__0__SCAN_IN,
         P3_INSTQUEUE_REG_14__7__SCAN_IN, P3_INSTQUEUE_REG_14__6__SCAN_IN,
         P3_INSTQUEUE_REG_14__5__SCAN_IN, P3_INSTQUEUE_REG_14__4__SCAN_IN,
         P3_INSTQUEUE_REG_14__3__SCAN_IN, P3_INSTQUEUE_REG_14__2__SCAN_IN,
         P3_INSTQUEUE_REG_14__1__SCAN_IN, P3_INSTQUEUE_REG_14__0__SCAN_IN,
         P3_INSTQUEUE_REG_13__7__SCAN_IN, P3_INSTQUEUE_REG_13__6__SCAN_IN,
         P3_INSTQUEUE_REG_13__5__SCAN_IN, P3_INSTQUEUE_REG_13__4__SCAN_IN,
         P3_INSTQUEUE_REG_13__3__SCAN_IN, P3_INSTQUEUE_REG_13__2__SCAN_IN,
         P3_INSTQUEUE_REG_13__1__SCAN_IN, P3_INSTQUEUE_REG_13__0__SCAN_IN,
         P3_INSTQUEUE_REG_12__7__SCAN_IN, P3_INSTQUEUE_REG_12__6__SCAN_IN,
         P3_INSTQUEUE_REG_12__5__SCAN_IN, P3_INSTQUEUE_REG_12__4__SCAN_IN,
         P3_INSTQUEUE_REG_12__3__SCAN_IN, P3_INSTQUEUE_REG_12__2__SCAN_IN,
         P3_INSTQUEUE_REG_12__1__SCAN_IN, P3_INSTQUEUE_REG_12__0__SCAN_IN,
         P3_INSTQUEUE_REG_11__7__SCAN_IN, P3_INSTQUEUE_REG_11__6__SCAN_IN,
         P3_INSTQUEUE_REG_11__5__SCAN_IN, P3_INSTQUEUE_REG_11__4__SCAN_IN,
         P3_INSTQUEUE_REG_11__3__SCAN_IN, P3_INSTQUEUE_REG_11__2__SCAN_IN,
         P3_INSTQUEUE_REG_11__1__SCAN_IN, P3_INSTQUEUE_REG_11__0__SCAN_IN,
         P3_INSTQUEUE_REG_10__7__SCAN_IN, P3_INSTQUEUE_REG_10__6__SCAN_IN,
         P3_INSTQUEUE_REG_10__5__SCAN_IN, P3_INSTQUEUE_REG_10__4__SCAN_IN,
         P3_INSTQUEUE_REG_10__3__SCAN_IN, P3_INSTQUEUE_REG_10__2__SCAN_IN,
         P3_INSTQUEUE_REG_10__1__SCAN_IN, P3_INSTQUEUE_REG_10__0__SCAN_IN,
         P3_INSTQUEUE_REG_9__7__SCAN_IN, P3_INSTQUEUE_REG_9__6__SCAN_IN,
         P3_INSTQUEUE_REG_9__5__SCAN_IN, P3_INSTQUEUE_REG_9__4__SCAN_IN,
         P3_INSTQUEUE_REG_9__3__SCAN_IN, P3_INSTQUEUE_REG_9__2__SCAN_IN,
         P3_INSTQUEUE_REG_9__1__SCAN_IN, P3_INSTQUEUE_REG_9__0__SCAN_IN,
         P3_INSTQUEUE_REG_8__7__SCAN_IN, P3_INSTQUEUE_REG_8__6__SCAN_IN,
         P3_INSTQUEUE_REG_8__5__SCAN_IN, P3_INSTQUEUE_REG_8__4__SCAN_IN,
         P3_INSTQUEUE_REG_8__3__SCAN_IN, P3_INSTQUEUE_REG_8__2__SCAN_IN,
         P3_INSTQUEUE_REG_8__1__SCAN_IN, P3_INSTQUEUE_REG_8__0__SCAN_IN,
         P3_INSTQUEUE_REG_7__7__SCAN_IN, P3_INSTQUEUE_REG_7__6__SCAN_IN,
         P3_INSTQUEUE_REG_7__5__SCAN_IN, P3_INSTQUEUE_REG_7__4__SCAN_IN,
         P3_INSTQUEUE_REG_7__3__SCAN_IN, P3_INSTQUEUE_REG_7__2__SCAN_IN,
         P3_INSTQUEUE_REG_7__1__SCAN_IN, P3_INSTQUEUE_REG_7__0__SCAN_IN,
         P3_INSTQUEUE_REG_6__7__SCAN_IN, P3_INSTQUEUE_REG_6__6__SCAN_IN,
         P3_INSTQUEUE_REG_6__5__SCAN_IN, P3_INSTQUEUE_REG_6__4__SCAN_IN,
         P3_INSTQUEUE_REG_6__3__SCAN_IN, P3_INSTQUEUE_REG_6__2__SCAN_IN,
         P3_INSTQUEUE_REG_6__1__SCAN_IN, P3_INSTQUEUE_REG_6__0__SCAN_IN,
         P3_INSTQUEUE_REG_5__7__SCAN_IN, P3_INSTQUEUE_REG_5__6__SCAN_IN,
         P3_INSTQUEUE_REG_5__5__SCAN_IN, P3_INSTQUEUE_REG_5__4__SCAN_IN,
         P3_INSTQUEUE_REG_5__3__SCAN_IN, P3_INSTQUEUE_REG_5__2__SCAN_IN,
         P3_INSTQUEUE_REG_5__1__SCAN_IN, P3_INSTQUEUE_REG_5__0__SCAN_IN,
         P3_INSTQUEUE_REG_4__7__SCAN_IN, P3_INSTQUEUE_REG_4__6__SCAN_IN,
         P3_INSTQUEUE_REG_4__5__SCAN_IN, P3_INSTQUEUE_REG_4__4__SCAN_IN,
         P3_INSTQUEUE_REG_4__3__SCAN_IN, P3_INSTQUEUE_REG_4__2__SCAN_IN,
         P3_INSTQUEUE_REG_4__1__SCAN_IN, P3_INSTQUEUE_REG_4__0__SCAN_IN,
         P3_INSTQUEUE_REG_3__7__SCAN_IN, P3_INSTQUEUE_REG_3__6__SCAN_IN,
         P3_INSTQUEUE_REG_3__5__SCAN_IN, P3_INSTQUEUE_REG_3__4__SCAN_IN,
         P3_INSTQUEUE_REG_3__3__SCAN_IN, P3_INSTQUEUE_REG_3__2__SCAN_IN,
         P3_INSTQUEUE_REG_3__1__SCAN_IN, P3_INSTQUEUE_REG_3__0__SCAN_IN,
         P3_INSTQUEUE_REG_2__7__SCAN_IN, P3_INSTQUEUE_REG_2__6__SCAN_IN,
         P3_INSTQUEUE_REG_2__5__SCAN_IN, P3_INSTQUEUE_REG_2__4__SCAN_IN,
         P3_INSTQUEUE_REG_2__3__SCAN_IN, P3_INSTQUEUE_REG_2__2__SCAN_IN,
         P3_INSTQUEUE_REG_2__1__SCAN_IN, P3_INSTQUEUE_REG_2__0__SCAN_IN,
         P3_INSTQUEUE_REG_1__7__SCAN_IN, P3_INSTQUEUE_REG_1__6__SCAN_IN,
         P3_INSTQUEUE_REG_1__5__SCAN_IN, P3_INSTQUEUE_REG_1__4__SCAN_IN,
         P3_INSTQUEUE_REG_1__3__SCAN_IN, P3_INSTQUEUE_REG_1__2__SCAN_IN,
         P3_INSTQUEUE_REG_1__1__SCAN_IN, P3_INSTQUEUE_REG_1__0__SCAN_IN,
         P3_INSTQUEUE_REG_0__7__SCAN_IN, P3_INSTQUEUE_REG_0__6__SCAN_IN,
         P3_INSTQUEUE_REG_0__5__SCAN_IN, P3_INSTQUEUE_REG_0__4__SCAN_IN,
         P3_INSTQUEUE_REG_0__3__SCAN_IN, P3_INSTQUEUE_REG_0__2__SCAN_IN,
         P3_INSTQUEUE_REG_0__1__SCAN_IN, P3_INSTQUEUE_REG_0__0__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P3_INSTADDRPOINTER_REG_0__SCAN_IN,
         P3_INSTADDRPOINTER_REG_1__SCAN_IN, P3_INSTADDRPOINTER_REG_2__SCAN_IN,
         P3_INSTADDRPOINTER_REG_3__SCAN_IN, P3_INSTADDRPOINTER_REG_4__SCAN_IN,
         P3_INSTADDRPOINTER_REG_5__SCAN_IN, P3_INSTADDRPOINTER_REG_6__SCAN_IN,
         P3_INSTADDRPOINTER_REG_7__SCAN_IN, P3_INSTADDRPOINTER_REG_8__SCAN_IN,
         P3_INSTADDRPOINTER_REG_9__SCAN_IN, P3_INSTADDRPOINTER_REG_10__SCAN_IN,
         P3_INSTADDRPOINTER_REG_11__SCAN_IN,
         P3_INSTADDRPOINTER_REG_12__SCAN_IN,
         P3_INSTADDRPOINTER_REG_13__SCAN_IN,
         P3_INSTADDRPOINTER_REG_14__SCAN_IN,
         P3_INSTADDRPOINTER_REG_15__SCAN_IN,
         P3_INSTADDRPOINTER_REG_16__SCAN_IN,
         P3_INSTADDRPOINTER_REG_17__SCAN_IN,
         P3_INSTADDRPOINTER_REG_18__SCAN_IN,
         P3_INSTADDRPOINTER_REG_19__SCAN_IN,
         P3_INSTADDRPOINTER_REG_20__SCAN_IN,
         P3_INSTADDRPOINTER_REG_21__SCAN_IN,
         P3_INSTADDRPOINTER_REG_22__SCAN_IN,
         P3_INSTADDRPOINTER_REG_23__SCAN_IN,
         P3_INSTADDRPOINTER_REG_24__SCAN_IN,
         P3_INSTADDRPOINTER_REG_25__SCAN_IN,
         P3_INSTADDRPOINTER_REG_26__SCAN_IN,
         P3_INSTADDRPOINTER_REG_27__SCAN_IN,
         P3_INSTADDRPOINTER_REG_28__SCAN_IN,
         P3_INSTADDRPOINTER_REG_29__SCAN_IN,
         P3_INSTADDRPOINTER_REG_30__SCAN_IN,
         P3_INSTADDRPOINTER_REG_31__SCAN_IN, P3_PHYADDRPOINTER_REG_0__SCAN_IN,
         P3_PHYADDRPOINTER_REG_1__SCAN_IN, P3_PHYADDRPOINTER_REG_2__SCAN_IN,
         P3_PHYADDRPOINTER_REG_3__SCAN_IN, P3_PHYADDRPOINTER_REG_4__SCAN_IN,
         P3_PHYADDRPOINTER_REG_5__SCAN_IN, P3_PHYADDRPOINTER_REG_6__SCAN_IN,
         P3_PHYADDRPOINTER_REG_7__SCAN_IN, P3_PHYADDRPOINTER_REG_8__SCAN_IN,
         P3_PHYADDRPOINTER_REG_9__SCAN_IN, P3_PHYADDRPOINTER_REG_10__SCAN_IN,
         P3_PHYADDRPOINTER_REG_11__SCAN_IN, P3_PHYADDRPOINTER_REG_12__SCAN_IN,
         P3_PHYADDRPOINTER_REG_13__SCAN_IN, P3_PHYADDRPOINTER_REG_14__SCAN_IN,
         P3_PHYADDRPOINTER_REG_15__SCAN_IN, P3_PHYADDRPOINTER_REG_16__SCAN_IN,
         P3_PHYADDRPOINTER_REG_17__SCAN_IN, P3_PHYADDRPOINTER_REG_18__SCAN_IN,
         P3_PHYADDRPOINTER_REG_19__SCAN_IN, P3_PHYADDRPOINTER_REG_20__SCAN_IN,
         P3_PHYADDRPOINTER_REG_21__SCAN_IN, P3_PHYADDRPOINTER_REG_22__SCAN_IN,
         P3_PHYADDRPOINTER_REG_23__SCAN_IN, P3_PHYADDRPOINTER_REG_24__SCAN_IN,
         P3_PHYADDRPOINTER_REG_25__SCAN_IN, P3_PHYADDRPOINTER_REG_26__SCAN_IN,
         P3_PHYADDRPOINTER_REG_27__SCAN_IN, P3_PHYADDRPOINTER_REG_28__SCAN_IN,
         P3_PHYADDRPOINTER_REG_29__SCAN_IN, P3_PHYADDRPOINTER_REG_30__SCAN_IN,
         P3_PHYADDRPOINTER_REG_31__SCAN_IN, P3_LWORD_REG_15__SCAN_IN,
         P3_LWORD_REG_14__SCAN_IN, P3_LWORD_REG_13__SCAN_IN,
         P3_LWORD_REG_12__SCAN_IN, P3_LWORD_REG_11__SCAN_IN,
         P3_LWORD_REG_10__SCAN_IN, P3_LWORD_REG_9__SCAN_IN,
         P3_LWORD_REG_8__SCAN_IN, P3_LWORD_REG_7__SCAN_IN,
         P3_LWORD_REG_6__SCAN_IN, P3_LWORD_REG_5__SCAN_IN,
         P3_LWORD_REG_4__SCAN_IN, P3_LWORD_REG_3__SCAN_IN,
         P3_LWORD_REG_2__SCAN_IN, P3_LWORD_REG_1__SCAN_IN,
         P3_LWORD_REG_0__SCAN_IN, P3_UWORD_REG_14__SCAN_IN,
         P3_UWORD_REG_13__SCAN_IN, P3_UWORD_REG_12__SCAN_IN,
         P3_UWORD_REG_11__SCAN_IN, P3_UWORD_REG_10__SCAN_IN,
         P3_UWORD_REG_9__SCAN_IN, P3_UWORD_REG_8__SCAN_IN,
         P3_UWORD_REG_7__SCAN_IN, P3_UWORD_REG_6__SCAN_IN,
         P3_UWORD_REG_5__SCAN_IN, P3_UWORD_REG_4__SCAN_IN,
         P3_UWORD_REG_3__SCAN_IN, P3_UWORD_REG_2__SCAN_IN,
         P3_UWORD_REG_1__SCAN_IN, P3_UWORD_REG_0__SCAN_IN,
         P3_DATAO_REG_0__SCAN_IN, P3_DATAO_REG_1__SCAN_IN,
         P3_DATAO_REG_2__SCAN_IN, P3_DATAO_REG_3__SCAN_IN,
         P3_DATAO_REG_4__SCAN_IN, P3_DATAO_REG_5__SCAN_IN,
         P3_DATAO_REG_6__SCAN_IN, P3_DATAO_REG_7__SCAN_IN,
         P3_DATAO_REG_8__SCAN_IN, P3_DATAO_REG_9__SCAN_IN,
         P3_DATAO_REG_10__SCAN_IN, P3_DATAO_REG_11__SCAN_IN,
         P3_DATAO_REG_12__SCAN_IN, P3_DATAO_REG_13__SCAN_IN,
         P3_DATAO_REG_14__SCAN_IN, P3_DATAO_REG_15__SCAN_IN,
         P3_DATAO_REG_16__SCAN_IN, P3_DATAO_REG_17__SCAN_IN,
         P3_DATAO_REG_18__SCAN_IN, P3_DATAO_REG_19__SCAN_IN,
         P3_DATAO_REG_20__SCAN_IN, P3_DATAO_REG_21__SCAN_IN,
         P3_DATAO_REG_22__SCAN_IN, P3_DATAO_REG_23__SCAN_IN,
         P3_DATAO_REG_24__SCAN_IN, P3_DATAO_REG_25__SCAN_IN,
         P3_DATAO_REG_26__SCAN_IN, P3_DATAO_REG_27__SCAN_IN,
         P3_DATAO_REG_28__SCAN_IN, P3_DATAO_REG_29__SCAN_IN,
         P3_DATAO_REG_30__SCAN_IN, P3_DATAO_REG_31__SCAN_IN,
         P3_EAX_REG_0__SCAN_IN, P3_EAX_REG_1__SCAN_IN, P3_EAX_REG_2__SCAN_IN,
         P3_EAX_REG_3__SCAN_IN, P3_EAX_REG_4__SCAN_IN, P3_EAX_REG_5__SCAN_IN,
         P3_EAX_REG_6__SCAN_IN, P3_EAX_REG_7__SCAN_IN, P3_EAX_REG_8__SCAN_IN,
         P3_EAX_REG_9__SCAN_IN, P3_EAX_REG_10__SCAN_IN, P3_EAX_REG_11__SCAN_IN,
         P3_EAX_REG_12__SCAN_IN, P3_EAX_REG_13__SCAN_IN,
         P3_EAX_REG_14__SCAN_IN, P3_EAX_REG_15__SCAN_IN,
         P3_EAX_REG_16__SCAN_IN, P3_EAX_REG_17__SCAN_IN,
         P3_EAX_REG_18__SCAN_IN, P3_EAX_REG_19__SCAN_IN,
         P3_EAX_REG_20__SCAN_IN, P3_EAX_REG_21__SCAN_IN,
         P3_EAX_REG_22__SCAN_IN, P3_EAX_REG_23__SCAN_IN,
         P3_EAX_REG_24__SCAN_IN, P3_EAX_REG_25__SCAN_IN,
         P3_EAX_REG_26__SCAN_IN, P3_EAX_REG_27__SCAN_IN,
         P3_EAX_REG_28__SCAN_IN, P3_EAX_REG_29__SCAN_IN,
         P3_EAX_REG_30__SCAN_IN, P3_EAX_REG_31__SCAN_IN, P3_EBX_REG_0__SCAN_IN,
         P3_EBX_REG_1__SCAN_IN, P3_EBX_REG_2__SCAN_IN, P3_EBX_REG_3__SCAN_IN,
         P3_EBX_REG_4__SCAN_IN, P3_EBX_REG_5__SCAN_IN, P3_EBX_REG_6__SCAN_IN,
         P3_EBX_REG_7__SCAN_IN, P3_EBX_REG_8__SCAN_IN, P3_EBX_REG_9__SCAN_IN,
         P3_EBX_REG_10__SCAN_IN, P3_EBX_REG_11__SCAN_IN,
         P3_EBX_REG_12__SCAN_IN, P3_EBX_REG_13__SCAN_IN,
         P3_EBX_REG_14__SCAN_IN, P3_EBX_REG_15__SCAN_IN,
         P3_EBX_REG_16__SCAN_IN, P3_EBX_REG_17__SCAN_IN,
         P3_EBX_REG_18__SCAN_IN, P3_EBX_REG_19__SCAN_IN,
         P3_EBX_REG_20__SCAN_IN, P3_EBX_REG_21__SCAN_IN,
         P3_EBX_REG_22__SCAN_IN, P3_EBX_REG_23__SCAN_IN,
         P3_EBX_REG_24__SCAN_IN, P3_EBX_REG_25__SCAN_IN,
         P3_EBX_REG_26__SCAN_IN, P3_EBX_REG_27__SCAN_IN,
         P3_EBX_REG_28__SCAN_IN, P3_EBX_REG_29__SCAN_IN,
         P3_EBX_REG_30__SCAN_IN, P3_EBX_REG_31__SCAN_IN,
         P3_REIP_REG_0__SCAN_IN, P3_REIP_REG_1__SCAN_IN,
         P3_REIP_REG_2__SCAN_IN, P3_REIP_REG_3__SCAN_IN,
         P3_REIP_REG_4__SCAN_IN, P3_REIP_REG_5__SCAN_IN,
         P3_REIP_REG_6__SCAN_IN, P3_REIP_REG_7__SCAN_IN,
         P3_REIP_REG_8__SCAN_IN, P3_REIP_REG_9__SCAN_IN,
         P3_REIP_REG_10__SCAN_IN, P3_REIP_REG_11__SCAN_IN,
         P3_REIP_REG_12__SCAN_IN, P3_REIP_REG_13__SCAN_IN,
         P3_REIP_REG_14__SCAN_IN, P3_REIP_REG_15__SCAN_IN,
         P3_REIP_REG_16__SCAN_IN, P3_REIP_REG_17__SCAN_IN,
         P3_REIP_REG_18__SCAN_IN, P3_REIP_REG_19__SCAN_IN,
         P3_REIP_REG_20__SCAN_IN, P3_REIP_REG_21__SCAN_IN,
         P3_REIP_REG_22__SCAN_IN, P3_REIP_REG_23__SCAN_IN,
         P3_REIP_REG_24__SCAN_IN, P3_REIP_REG_25__SCAN_IN,
         P3_REIP_REG_26__SCAN_IN, P3_REIP_REG_27__SCAN_IN,
         P3_REIP_REG_28__SCAN_IN, P3_REIP_REG_29__SCAN_IN,
         P3_REIP_REG_30__SCAN_IN, P3_REIP_REG_31__SCAN_IN,
         P3_BYTEENABLE_REG_3__SCAN_IN, P3_BYTEENABLE_REG_2__SCAN_IN,
         P3_BYTEENABLE_REG_1__SCAN_IN, P3_BYTEENABLE_REG_0__SCAN_IN,
         P3_W_R_N_REG_SCAN_IN, P3_FLUSH_REG_SCAN_IN, P3_MORE_REG_SCAN_IN,
         P3_STATEBS16_REG_SCAN_IN, P3_REQUESTPENDING_REG_SCAN_IN,
         P3_D_C_N_REG_SCAN_IN, P3_M_IO_N_REG_SCAN_IN, P3_CODEFETCH_REG_SCAN_IN,
         P3_ADS_N_REG_SCAN_IN, P3_READREQUEST_REG_SCAN_IN,
         P3_MEMORYFETCH_REG_SCAN_IN, P2_BE_N_REG_3__SCAN_IN,
         P2_BE_N_REG_2__SCAN_IN, P2_BE_N_REG_1__SCAN_IN,
         P2_BE_N_REG_0__SCAN_IN, P2_ADDRESS_REG_29__SCAN_IN,
         P2_ADDRESS_REG_28__SCAN_IN, P2_ADDRESS_REG_27__SCAN_IN,
         P2_ADDRESS_REG_26__SCAN_IN, P2_ADDRESS_REG_25__SCAN_IN,
         P2_ADDRESS_REG_24__SCAN_IN, P2_ADDRESS_REG_23__SCAN_IN,
         P2_ADDRESS_REG_22__SCAN_IN, P2_ADDRESS_REG_21__SCAN_IN,
         P2_ADDRESS_REG_20__SCAN_IN, P2_ADDRESS_REG_19__SCAN_IN,
         P2_ADDRESS_REG_18__SCAN_IN, P2_ADDRESS_REG_17__SCAN_IN,
         P2_ADDRESS_REG_16__SCAN_IN, P2_ADDRESS_REG_15__SCAN_IN,
         P2_ADDRESS_REG_14__SCAN_IN, P2_ADDRESS_REG_13__SCAN_IN,
         P2_ADDRESS_REG_12__SCAN_IN, P2_ADDRESS_REG_11__SCAN_IN,
         P2_ADDRESS_REG_10__SCAN_IN, P2_ADDRESS_REG_9__SCAN_IN,
         P2_ADDRESS_REG_8__SCAN_IN, P2_ADDRESS_REG_7__SCAN_IN,
         P2_ADDRESS_REG_6__SCAN_IN, P2_ADDRESS_REG_5__SCAN_IN,
         P2_ADDRESS_REG_4__SCAN_IN, P2_ADDRESS_REG_3__SCAN_IN,
         P2_ADDRESS_REG_2__SCAN_IN, P2_ADDRESS_REG_1__SCAN_IN,
         P2_ADDRESS_REG_0__SCAN_IN, P2_STATE_REG_2__SCAN_IN,
         P2_STATE_REG_1__SCAN_IN, P2_STATE_REG_0__SCAN_IN,
         P2_DATAWIDTH_REG_0__SCAN_IN, P2_DATAWIDTH_REG_1__SCAN_IN,
         P2_DATAWIDTH_REG_2__SCAN_IN, P2_DATAWIDTH_REG_3__SCAN_IN,
         P2_DATAWIDTH_REG_4__SCAN_IN, P2_DATAWIDTH_REG_5__SCAN_IN,
         P2_DATAWIDTH_REG_6__SCAN_IN, P2_DATAWIDTH_REG_7__SCAN_IN,
         P2_DATAWIDTH_REG_8__SCAN_IN, P2_DATAWIDTH_REG_9__SCAN_IN,
         P2_DATAWIDTH_REG_10__SCAN_IN, P2_DATAWIDTH_REG_11__SCAN_IN,
         P2_DATAWIDTH_REG_12__SCAN_IN, P2_DATAWIDTH_REG_13__SCAN_IN,
         P2_DATAWIDTH_REG_14__SCAN_IN, P2_DATAWIDTH_REG_15__SCAN_IN,
         P2_DATAWIDTH_REG_16__SCAN_IN, P2_DATAWIDTH_REG_17__SCAN_IN,
         P2_DATAWIDTH_REG_18__SCAN_IN, P2_DATAWIDTH_REG_19__SCAN_IN,
         P2_DATAWIDTH_REG_20__SCAN_IN, P2_DATAWIDTH_REG_21__SCAN_IN,
         P2_DATAWIDTH_REG_22__SCAN_IN, P2_DATAWIDTH_REG_23__SCAN_IN,
         P2_DATAWIDTH_REG_24__SCAN_IN, P2_DATAWIDTH_REG_25__SCAN_IN,
         P2_DATAWIDTH_REG_26__SCAN_IN, P2_DATAWIDTH_REG_27__SCAN_IN,
         P2_DATAWIDTH_REG_28__SCAN_IN, P2_DATAWIDTH_REG_29__SCAN_IN,
         P2_DATAWIDTH_REG_30__SCAN_IN, P2_DATAWIDTH_REG_31__SCAN_IN,
         P2_STATE2_REG_3__SCAN_IN, P2_STATE2_REG_2__SCAN_IN,
         P2_STATE2_REG_1__SCAN_IN, P2_STATE2_REG_0__SCAN_IN,
         P2_INSTQUEUE_REG_15__7__SCAN_IN, P2_INSTQUEUE_REG_15__6__SCAN_IN,
         P2_INSTQUEUE_REG_15__5__SCAN_IN, P2_INSTQUEUE_REG_15__4__SCAN_IN,
         P2_INSTQUEUE_REG_15__3__SCAN_IN, P2_INSTQUEUE_REG_15__2__SCAN_IN,
         P2_INSTQUEUE_REG_15__1__SCAN_IN, P2_INSTQUEUE_REG_15__0__SCAN_IN,
         P2_INSTQUEUE_REG_14__7__SCAN_IN, P2_INSTQUEUE_REG_14__6__SCAN_IN,
         P2_INSTQUEUE_REG_14__5__SCAN_IN, P2_INSTQUEUE_REG_14__4__SCAN_IN,
         P2_INSTQUEUE_REG_14__3__SCAN_IN, P2_INSTQUEUE_REG_14__2__SCAN_IN,
         P2_INSTQUEUE_REG_14__1__SCAN_IN, P2_INSTQUEUE_REG_14__0__SCAN_IN,
         P2_INSTQUEUE_REG_13__7__SCAN_IN, P2_INSTQUEUE_REG_13__6__SCAN_IN,
         P2_INSTQUEUE_REG_13__5__SCAN_IN, P2_INSTQUEUE_REG_13__4__SCAN_IN,
         P2_INSTQUEUE_REG_13__3__SCAN_IN, P2_INSTQUEUE_REG_13__2__SCAN_IN,
         P2_INSTQUEUE_REG_13__1__SCAN_IN, P2_INSTQUEUE_REG_13__0__SCAN_IN,
         P2_INSTQUEUE_REG_12__7__SCAN_IN, P2_INSTQUEUE_REG_12__6__SCAN_IN,
         P2_INSTQUEUE_REG_12__5__SCAN_IN, P2_INSTQUEUE_REG_12__4__SCAN_IN,
         P2_INSTQUEUE_REG_12__3__SCAN_IN, P2_INSTQUEUE_REG_12__2__SCAN_IN,
         P2_INSTQUEUE_REG_12__1__SCAN_IN, P2_INSTQUEUE_REG_12__0__SCAN_IN,
         P2_INSTQUEUE_REG_11__7__SCAN_IN, P2_INSTQUEUE_REG_11__6__SCAN_IN,
         P2_INSTQUEUE_REG_11__5__SCAN_IN, P2_INSTQUEUE_REG_11__4__SCAN_IN,
         P2_INSTQUEUE_REG_11__3__SCAN_IN, P2_INSTQUEUE_REG_11__2__SCAN_IN,
         P2_INSTQUEUE_REG_11__1__SCAN_IN, P2_INSTQUEUE_REG_11__0__SCAN_IN,
         P2_INSTQUEUE_REG_10__7__SCAN_IN, P2_INSTQUEUE_REG_10__6__SCAN_IN,
         P2_INSTQUEUE_REG_10__5__SCAN_IN, P2_INSTQUEUE_REG_10__4__SCAN_IN,
         P2_INSTQUEUE_REG_10__3__SCAN_IN, P2_INSTQUEUE_REG_10__2__SCAN_IN,
         P2_INSTQUEUE_REG_10__1__SCAN_IN, P2_INSTQUEUE_REG_10__0__SCAN_IN,
         P2_INSTQUEUE_REG_9__7__SCAN_IN, P2_INSTQUEUE_REG_9__6__SCAN_IN,
         P2_INSTQUEUE_REG_9__5__SCAN_IN, P2_INSTQUEUE_REG_9__4__SCAN_IN,
         P2_INSTQUEUE_REG_9__3__SCAN_IN, P2_INSTQUEUE_REG_9__2__SCAN_IN,
         P2_INSTQUEUE_REG_9__1__SCAN_IN, P2_INSTQUEUE_REG_9__0__SCAN_IN,
         P2_INSTQUEUE_REG_8__7__SCAN_IN, P2_INSTQUEUE_REG_8__6__SCAN_IN,
         P2_INSTQUEUE_REG_8__5__SCAN_IN, P2_INSTQUEUE_REG_8__4__SCAN_IN,
         P2_INSTQUEUE_REG_8__3__SCAN_IN, P2_INSTQUEUE_REG_8__2__SCAN_IN,
         P2_INSTQUEUE_REG_8__1__SCAN_IN, P2_INSTQUEUE_REG_8__0__SCAN_IN,
         P2_INSTQUEUE_REG_7__7__SCAN_IN, P2_INSTQUEUE_REG_7__6__SCAN_IN,
         P2_INSTQUEUE_REG_7__5__SCAN_IN, P2_INSTQUEUE_REG_7__4__SCAN_IN,
         P2_INSTQUEUE_REG_7__3__SCAN_IN, P2_INSTQUEUE_REG_7__2__SCAN_IN,
         P2_INSTQUEUE_REG_7__1__SCAN_IN, P2_INSTQUEUE_REG_7__0__SCAN_IN,
         P2_INSTQUEUE_REG_6__7__SCAN_IN, P2_INSTQUEUE_REG_6__6__SCAN_IN,
         P2_INSTQUEUE_REG_6__5__SCAN_IN, P2_INSTQUEUE_REG_6__4__SCAN_IN,
         P2_INSTQUEUE_REG_6__3__SCAN_IN, P2_INSTQUEUE_REG_6__2__SCAN_IN,
         P2_INSTQUEUE_REG_6__1__SCAN_IN, P2_INSTQUEUE_REG_6__0__SCAN_IN,
         P2_INSTQUEUE_REG_5__7__SCAN_IN, P2_INSTQUEUE_REG_5__6__SCAN_IN,
         P2_INSTQUEUE_REG_5__5__SCAN_IN, P2_INSTQUEUE_REG_5__4__SCAN_IN,
         P2_INSTQUEUE_REG_5__3__SCAN_IN, P2_INSTQUEUE_REG_5__2__SCAN_IN,
         P2_INSTQUEUE_REG_5__1__SCAN_IN, P2_INSTQUEUE_REG_5__0__SCAN_IN,
         P2_INSTQUEUE_REG_4__7__SCAN_IN, P2_INSTQUEUE_REG_4__6__SCAN_IN,
         P2_INSTQUEUE_REG_4__5__SCAN_IN, P2_INSTQUEUE_REG_4__4__SCAN_IN,
         P2_INSTQUEUE_REG_4__3__SCAN_IN, P2_INSTQUEUE_REG_4__2__SCAN_IN,
         P2_INSTQUEUE_REG_4__1__SCAN_IN, P2_INSTQUEUE_REG_4__0__SCAN_IN,
         P2_INSTQUEUE_REG_3__7__SCAN_IN, P2_INSTQUEUE_REG_3__6__SCAN_IN,
         P2_INSTQUEUE_REG_3__5__SCAN_IN, P2_INSTQUEUE_REG_3__4__SCAN_IN,
         P2_INSTQUEUE_REG_3__3__SCAN_IN, P2_INSTQUEUE_REG_3__2__SCAN_IN,
         P2_INSTQUEUE_REG_3__1__SCAN_IN, P2_INSTQUEUE_REG_3__0__SCAN_IN,
         P2_INSTQUEUE_REG_2__7__SCAN_IN, P2_INSTQUEUE_REG_2__6__SCAN_IN,
         P2_INSTQUEUE_REG_2__5__SCAN_IN, P2_INSTQUEUE_REG_2__4__SCAN_IN,
         P2_INSTQUEUE_REG_2__3__SCAN_IN, P2_INSTQUEUE_REG_2__2__SCAN_IN,
         P2_INSTQUEUE_REG_2__1__SCAN_IN, P2_INSTQUEUE_REG_2__0__SCAN_IN,
         P2_INSTQUEUE_REG_1__7__SCAN_IN, P2_INSTQUEUE_REG_1__6__SCAN_IN,
         P2_INSTQUEUE_REG_1__5__SCAN_IN, P2_INSTQUEUE_REG_1__4__SCAN_IN,
         P2_INSTQUEUE_REG_1__3__SCAN_IN, P2_INSTQUEUE_REG_1__2__SCAN_IN,
         P2_INSTQUEUE_REG_1__1__SCAN_IN, P2_INSTQUEUE_REG_1__0__SCAN_IN,
         P2_INSTQUEUE_REG_0__7__SCAN_IN, P2_INSTQUEUE_REG_0__6__SCAN_IN,
         P2_INSTQUEUE_REG_0__5__SCAN_IN, P2_INSTQUEUE_REG_0__4__SCAN_IN,
         P2_INSTQUEUE_REG_0__3__SCAN_IN, P2_INSTQUEUE_REG_0__2__SCAN_IN,
         P2_INSTQUEUE_REG_0__1__SCAN_IN, P2_INSTQUEUE_REG_0__0__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN,
         P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN, P2_INSTADDRPOINTER_REG_0__SCAN_IN,
         P2_INSTADDRPOINTER_REG_1__SCAN_IN, P2_INSTADDRPOINTER_REG_2__SCAN_IN,
         P2_INSTADDRPOINTER_REG_3__SCAN_IN, P2_INSTADDRPOINTER_REG_4__SCAN_IN,
         P2_INSTADDRPOINTER_REG_5__SCAN_IN, P2_INSTADDRPOINTER_REG_6__SCAN_IN,
         P2_INSTADDRPOINTER_REG_7__SCAN_IN, P2_INSTADDRPOINTER_REG_8__SCAN_IN,
         P2_INSTADDRPOINTER_REG_9__SCAN_IN, P2_INSTADDRPOINTER_REG_10__SCAN_IN,
         P2_INSTADDRPOINTER_REG_11__SCAN_IN,
         P2_INSTADDRPOINTER_REG_12__SCAN_IN,
         P2_INSTADDRPOINTER_REG_13__SCAN_IN,
         P2_INSTADDRPOINTER_REG_14__SCAN_IN,
         P2_INSTADDRPOINTER_REG_15__SCAN_IN,
         P2_INSTADDRPOINTER_REG_16__SCAN_IN,
         P2_INSTADDRPOINTER_REG_17__SCAN_IN,
         P2_INSTADDRPOINTER_REG_18__SCAN_IN,
         P2_INSTADDRPOINTER_REG_19__SCAN_IN,
         P2_INSTADDRPOINTER_REG_20__SCAN_IN,
         P2_INSTADDRPOINTER_REG_21__SCAN_IN,
         P2_INSTADDRPOINTER_REG_22__SCAN_IN,
         P2_INSTADDRPOINTER_REG_23__SCAN_IN,
         P2_INSTADDRPOINTER_REG_24__SCAN_IN,
         P2_INSTADDRPOINTER_REG_25__SCAN_IN,
         P2_INSTADDRPOINTER_REG_26__SCAN_IN,
         P2_INSTADDRPOINTER_REG_27__SCAN_IN,
         P2_INSTADDRPOINTER_REG_28__SCAN_IN,
         P2_INSTADDRPOINTER_REG_29__SCAN_IN,
         P2_INSTADDRPOINTER_REG_30__SCAN_IN,
         P2_INSTADDRPOINTER_REG_31__SCAN_IN, P2_PHYADDRPOINTER_REG_0__SCAN_IN,
         P2_PHYADDRPOINTER_REG_1__SCAN_IN, P2_PHYADDRPOINTER_REG_2__SCAN_IN,
         P2_PHYADDRPOINTER_REG_3__SCAN_IN, P2_PHYADDRPOINTER_REG_4__SCAN_IN,
         P2_PHYADDRPOINTER_REG_5__SCAN_IN, P2_PHYADDRPOINTER_REG_6__SCAN_IN,
         P2_PHYADDRPOINTER_REG_7__SCAN_IN, P2_PHYADDRPOINTER_REG_8__SCAN_IN,
         P2_PHYADDRPOINTER_REG_9__SCAN_IN, P2_PHYADDRPOINTER_REG_10__SCAN_IN,
         P2_PHYADDRPOINTER_REG_11__SCAN_IN, P2_PHYADDRPOINTER_REG_12__SCAN_IN,
         P2_PHYADDRPOINTER_REG_13__SCAN_IN, P2_PHYADDRPOINTER_REG_14__SCAN_IN,
         P2_PHYADDRPOINTER_REG_15__SCAN_IN, P2_PHYADDRPOINTER_REG_16__SCAN_IN,
         P2_PHYADDRPOINTER_REG_17__SCAN_IN, P2_PHYADDRPOINTER_REG_18__SCAN_IN,
         P2_PHYADDRPOINTER_REG_19__SCAN_IN, P2_PHYADDRPOINTER_REG_20__SCAN_IN,
         P2_PHYADDRPOINTER_REG_21__SCAN_IN, P2_PHYADDRPOINTER_REG_22__SCAN_IN,
         P2_PHYADDRPOINTER_REG_23__SCAN_IN, P2_PHYADDRPOINTER_REG_24__SCAN_IN,
         P2_PHYADDRPOINTER_REG_25__SCAN_IN, P2_PHYADDRPOINTER_REG_26__SCAN_IN,
         P2_PHYADDRPOINTER_REG_27__SCAN_IN, P2_PHYADDRPOINTER_REG_28__SCAN_IN,
         P2_PHYADDRPOINTER_REG_29__SCAN_IN, P2_PHYADDRPOINTER_REG_30__SCAN_IN,
         P2_PHYADDRPOINTER_REG_31__SCAN_IN, P2_LWORD_REG_15__SCAN_IN,
         P2_LWORD_REG_14__SCAN_IN, P2_LWORD_REG_13__SCAN_IN,
         P2_LWORD_REG_12__SCAN_IN, P2_LWORD_REG_11__SCAN_IN,
         P2_LWORD_REG_10__SCAN_IN, P2_LWORD_REG_9__SCAN_IN,
         P2_LWORD_REG_8__SCAN_IN, P2_LWORD_REG_7__SCAN_IN,
         P2_LWORD_REG_6__SCAN_IN, P2_LWORD_REG_5__SCAN_IN,
         P2_LWORD_REG_4__SCAN_IN, P2_LWORD_REG_3__SCAN_IN,
         P2_LWORD_REG_2__SCAN_IN, P2_LWORD_REG_1__SCAN_IN,
         P2_LWORD_REG_0__SCAN_IN, P2_UWORD_REG_14__SCAN_IN,
         P2_UWORD_REG_13__SCAN_IN, P2_UWORD_REG_12__SCAN_IN,
         P2_UWORD_REG_11__SCAN_IN, P2_UWORD_REG_10__SCAN_IN,
         P2_UWORD_REG_9__SCAN_IN, P2_UWORD_REG_8__SCAN_IN,
         P2_UWORD_REG_7__SCAN_IN, P2_UWORD_REG_6__SCAN_IN,
         P2_UWORD_REG_5__SCAN_IN, P2_UWORD_REG_4__SCAN_IN,
         P2_UWORD_REG_3__SCAN_IN, P2_UWORD_REG_2__SCAN_IN,
         P2_UWORD_REG_1__SCAN_IN, P2_UWORD_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_EAX_REG_0__SCAN_IN, P2_EAX_REG_1__SCAN_IN, P2_EAX_REG_2__SCAN_IN,
         P2_EAX_REG_3__SCAN_IN, P2_EAX_REG_4__SCAN_IN, P2_EAX_REG_5__SCAN_IN,
         P2_EAX_REG_6__SCAN_IN, P2_EAX_REG_7__SCAN_IN, P2_EAX_REG_8__SCAN_IN,
         P2_EAX_REG_9__SCAN_IN, P2_EAX_REG_10__SCAN_IN, P2_EAX_REG_11__SCAN_IN,
         P2_EAX_REG_12__SCAN_IN, P2_EAX_REG_13__SCAN_IN,
         P2_EAX_REG_14__SCAN_IN, P2_EAX_REG_15__SCAN_IN,
         P2_EAX_REG_16__SCAN_IN, P2_EAX_REG_17__SCAN_IN,
         P2_EAX_REG_18__SCAN_IN, P2_EAX_REG_19__SCAN_IN,
         P2_EAX_REG_20__SCAN_IN, P2_EAX_REG_21__SCAN_IN,
         P2_EAX_REG_22__SCAN_IN, P2_EAX_REG_23__SCAN_IN,
         P2_EAX_REG_24__SCAN_IN, P2_EAX_REG_25__SCAN_IN,
         P2_EAX_REG_26__SCAN_IN, P2_EAX_REG_27__SCAN_IN,
         P2_EAX_REG_28__SCAN_IN, P2_EAX_REG_29__SCAN_IN,
         P2_EAX_REG_30__SCAN_IN, P2_EAX_REG_31__SCAN_IN, P2_EBX_REG_0__SCAN_IN,
         P2_EBX_REG_1__SCAN_IN, P2_EBX_REG_2__SCAN_IN, P2_EBX_REG_3__SCAN_IN,
         P2_EBX_REG_4__SCAN_IN, P2_EBX_REG_5__SCAN_IN, P2_EBX_REG_6__SCAN_IN,
         P2_EBX_REG_7__SCAN_IN, P2_EBX_REG_8__SCAN_IN, P2_EBX_REG_9__SCAN_IN,
         P2_EBX_REG_10__SCAN_IN, P2_EBX_REG_11__SCAN_IN,
         P2_EBX_REG_12__SCAN_IN, P2_EBX_REG_13__SCAN_IN,
         P2_EBX_REG_14__SCAN_IN, P2_EBX_REG_15__SCAN_IN,
         P2_EBX_REG_16__SCAN_IN, P2_EBX_REG_17__SCAN_IN,
         P2_EBX_REG_18__SCAN_IN, P2_EBX_REG_19__SCAN_IN,
         P2_EBX_REG_20__SCAN_IN, P2_EBX_REG_21__SCAN_IN,
         P2_EBX_REG_22__SCAN_IN, P2_EBX_REG_23__SCAN_IN,
         P2_EBX_REG_24__SCAN_IN, P2_EBX_REG_25__SCAN_IN,
         P2_EBX_REG_26__SCAN_IN, P2_EBX_REG_27__SCAN_IN,
         P2_EBX_REG_28__SCAN_IN, P2_EBX_REG_29__SCAN_IN,
         P2_EBX_REG_30__SCAN_IN, P2_EBX_REG_31__SCAN_IN,
         P2_REIP_REG_0__SCAN_IN, P2_REIP_REG_1__SCAN_IN,
         P2_REIP_REG_2__SCAN_IN, P2_REIP_REG_3__SCAN_IN,
         P2_REIP_REG_4__SCAN_IN, P2_REIP_REG_5__SCAN_IN,
         P2_REIP_REG_6__SCAN_IN, P2_REIP_REG_7__SCAN_IN,
         P2_REIP_REG_8__SCAN_IN, P2_REIP_REG_9__SCAN_IN,
         P2_REIP_REG_10__SCAN_IN, P2_REIP_REG_11__SCAN_IN,
         P2_REIP_REG_12__SCAN_IN, P2_REIP_REG_13__SCAN_IN,
         P2_REIP_REG_14__SCAN_IN, P2_REIP_REG_15__SCAN_IN,
         P2_REIP_REG_16__SCAN_IN, P2_REIP_REG_17__SCAN_IN,
         P2_REIP_REG_18__SCAN_IN, P2_REIP_REG_19__SCAN_IN,
         P2_REIP_REG_20__SCAN_IN, P2_REIP_REG_21__SCAN_IN,
         P2_REIP_REG_22__SCAN_IN, P2_REIP_REG_23__SCAN_IN,
         P2_REIP_REG_24__SCAN_IN, P2_REIP_REG_25__SCAN_IN,
         P2_REIP_REG_26__SCAN_IN, P2_REIP_REG_27__SCAN_IN,
         P2_REIP_REG_28__SCAN_IN, P2_REIP_REG_29__SCAN_IN,
         P2_REIP_REG_30__SCAN_IN, P2_REIP_REG_31__SCAN_IN,
         P2_BYTEENABLE_REG_3__SCAN_IN, P2_BYTEENABLE_REG_2__SCAN_IN,
         P2_BYTEENABLE_REG_1__SCAN_IN, P2_BYTEENABLE_REG_0__SCAN_IN,
         P2_W_R_N_REG_SCAN_IN, P2_FLUSH_REG_SCAN_IN, P2_MORE_REG_SCAN_IN,
         P2_STATEBS16_REG_SCAN_IN, P2_REQUESTPENDING_REG_SCAN_IN,
         P2_D_C_N_REG_SCAN_IN, P2_M_IO_N_REG_SCAN_IN, P2_CODEFETCH_REG_SCAN_IN,
         P2_ADS_N_REG_SCAN_IN, P2_READREQUEST_REG_SCAN_IN,
         P2_MEMORYFETCH_REG_SCAN_IN, P1_BE_N_REG_3__SCAN_IN,
         P1_BE_N_REG_2__SCAN_IN, P1_BE_N_REG_1__SCAN_IN,
         P1_BE_N_REG_0__SCAN_IN, P1_ADDRESS_REG_29__SCAN_IN,
         P1_ADDRESS_REG_28__SCAN_IN, P1_ADDRESS_REG_27__SCAN_IN,
         P1_ADDRESS_REG_26__SCAN_IN, P1_ADDRESS_REG_25__SCAN_IN,
         P1_ADDRESS_REG_24__SCAN_IN, P1_ADDRESS_REG_23__SCAN_IN,
         P1_ADDRESS_REG_22__SCAN_IN, P1_ADDRESS_REG_21__SCAN_IN,
         P1_ADDRESS_REG_20__SCAN_IN, P1_ADDRESS_REG_19__SCAN_IN,
         P1_ADDRESS_REG_18__SCAN_IN, P1_ADDRESS_REG_17__SCAN_IN,
         P1_ADDRESS_REG_16__SCAN_IN, P1_ADDRESS_REG_15__SCAN_IN,
         P1_ADDRESS_REG_14__SCAN_IN, P1_ADDRESS_REG_13__SCAN_IN,
         P1_ADDRESS_REG_12__SCAN_IN, P1_ADDRESS_REG_11__SCAN_IN,
         P1_ADDRESS_REG_10__SCAN_IN, P1_ADDRESS_REG_9__SCAN_IN,
         P1_ADDRESS_REG_8__SCAN_IN, P1_ADDRESS_REG_7__SCAN_IN,
         P1_ADDRESS_REG_6__SCAN_IN, P1_ADDRESS_REG_5__SCAN_IN,
         P1_ADDRESS_REG_4__SCAN_IN, P1_ADDRESS_REG_3__SCAN_IN,
         P1_ADDRESS_REG_2__SCAN_IN, P1_ADDRESS_REG_1__SCAN_IN,
         P1_ADDRESS_REG_0__SCAN_IN, P1_STATE_REG_2__SCAN_IN,
         P1_STATE_REG_1__SCAN_IN, P1_STATE_REG_0__SCAN_IN,
         P1_DATAWIDTH_REG_0__SCAN_IN, P1_DATAWIDTH_REG_1__SCAN_IN,
         P1_DATAWIDTH_REG_2__SCAN_IN, P1_DATAWIDTH_REG_3__SCAN_IN,
         P1_DATAWIDTH_REG_4__SCAN_IN, P1_DATAWIDTH_REG_5__SCAN_IN,
         P1_DATAWIDTH_REG_6__SCAN_IN, P1_DATAWIDTH_REG_7__SCAN_IN,
         P1_DATAWIDTH_REG_8__SCAN_IN, P1_DATAWIDTH_REG_9__SCAN_IN,
         P1_DATAWIDTH_REG_10__SCAN_IN, P1_DATAWIDTH_REG_11__SCAN_IN,
         P1_DATAWIDTH_REG_12__SCAN_IN, P1_DATAWIDTH_REG_13__SCAN_IN,
         P1_DATAWIDTH_REG_14__SCAN_IN, P1_DATAWIDTH_REG_15__SCAN_IN,
         P1_DATAWIDTH_REG_16__SCAN_IN, P1_DATAWIDTH_REG_17__SCAN_IN,
         P1_DATAWIDTH_REG_18__SCAN_IN, P1_DATAWIDTH_REG_19__SCAN_IN,
         P1_DATAWIDTH_REG_20__SCAN_IN, P1_DATAWIDTH_REG_21__SCAN_IN,
         P1_DATAWIDTH_REG_22__SCAN_IN, P1_DATAWIDTH_REG_23__SCAN_IN,
         P1_DATAWIDTH_REG_24__SCAN_IN, P1_DATAWIDTH_REG_25__SCAN_IN,
         P1_DATAWIDTH_REG_26__SCAN_IN, P1_DATAWIDTH_REG_27__SCAN_IN,
         P1_DATAWIDTH_REG_28__SCAN_IN, P1_DATAWIDTH_REG_29__SCAN_IN,
         P1_DATAWIDTH_REG_30__SCAN_IN, P1_DATAWIDTH_REG_31__SCAN_IN,
         P1_STATE2_REG_3__SCAN_IN, P1_STATE2_REG_2__SCAN_IN,
         P1_STATE2_REG_1__SCAN_IN, P1_STATE2_REG_0__SCAN_IN,
         P1_INSTQUEUE_REG_15__7__SCAN_IN, P1_INSTQUEUE_REG_15__6__SCAN_IN,
         P1_INSTQUEUE_REG_15__5__SCAN_IN, P1_INSTQUEUE_REG_15__4__SCAN_IN,
         P1_INSTQUEUE_REG_15__3__SCAN_IN, P1_INSTQUEUE_REG_15__2__SCAN_IN,
         P1_INSTQUEUE_REG_15__1__SCAN_IN, P1_INSTQUEUE_REG_15__0__SCAN_IN,
         P1_INSTQUEUE_REG_14__7__SCAN_IN, P1_INSTQUEUE_REG_14__6__SCAN_IN,
         P1_INSTQUEUE_REG_14__5__SCAN_IN, P1_INSTQUEUE_REG_14__4__SCAN_IN,
         P1_INSTQUEUE_REG_14__3__SCAN_IN, P1_INSTQUEUE_REG_14__2__SCAN_IN,
         P1_INSTQUEUE_REG_14__1__SCAN_IN, P1_INSTQUEUE_REG_14__0__SCAN_IN,
         P1_INSTQUEUE_REG_13__7__SCAN_IN, P1_INSTQUEUE_REG_13__6__SCAN_IN,
         P1_INSTQUEUE_REG_13__5__SCAN_IN, P1_INSTQUEUE_REG_13__4__SCAN_IN,
         P1_INSTQUEUE_REG_13__3__SCAN_IN, P1_INSTQUEUE_REG_13__2__SCAN_IN,
         P1_INSTQUEUE_REG_13__1__SCAN_IN, P1_INSTQUEUE_REG_13__0__SCAN_IN,
         P1_INSTQUEUE_REG_12__7__SCAN_IN, P1_INSTQUEUE_REG_12__6__SCAN_IN,
         P1_INSTQUEUE_REG_12__5__SCAN_IN, P1_INSTQUEUE_REG_12__4__SCAN_IN,
         P1_INSTQUEUE_REG_12__3__SCAN_IN, P1_INSTQUEUE_REG_12__2__SCAN_IN,
         P1_INSTQUEUE_REG_12__1__SCAN_IN, P1_INSTQUEUE_REG_12__0__SCAN_IN,
         P1_INSTQUEUE_REG_11__7__SCAN_IN, P1_INSTQUEUE_REG_11__6__SCAN_IN,
         P1_INSTQUEUE_REG_11__5__SCAN_IN, P1_INSTQUEUE_REG_11__4__SCAN_IN,
         P1_INSTQUEUE_REG_11__3__SCAN_IN, P1_INSTQUEUE_REG_11__2__SCAN_IN,
         P1_INSTQUEUE_REG_11__1__SCAN_IN, P1_INSTQUEUE_REG_11__0__SCAN_IN,
         P1_INSTQUEUE_REG_10__7__SCAN_IN, P1_INSTQUEUE_REG_10__6__SCAN_IN,
         P1_INSTQUEUE_REG_10__5__SCAN_IN, P1_INSTQUEUE_REG_10__4__SCAN_IN,
         P1_INSTQUEUE_REG_10__3__SCAN_IN, P1_INSTQUEUE_REG_10__2__SCAN_IN,
         P1_INSTQUEUE_REG_10__1__SCAN_IN, P1_INSTQUEUE_REG_10__0__SCAN_IN,
         P1_INSTQUEUE_REG_9__7__SCAN_IN, P1_INSTQUEUE_REG_9__6__SCAN_IN,
         P1_INSTQUEUE_REG_9__5__SCAN_IN, P1_INSTQUEUE_REG_9__4__SCAN_IN,
         P1_INSTQUEUE_REG_9__3__SCAN_IN, P1_INSTQUEUE_REG_9__2__SCAN_IN,
         P1_INSTQUEUE_REG_9__1__SCAN_IN, P1_INSTQUEUE_REG_9__0__SCAN_IN,
         P1_INSTQUEUE_REG_8__7__SCAN_IN, P1_INSTQUEUE_REG_8__6__SCAN_IN,
         P1_INSTQUEUE_REG_8__5__SCAN_IN, P1_INSTQUEUE_REG_8__4__SCAN_IN,
         P1_INSTQUEUE_REG_8__3__SCAN_IN, P1_INSTQUEUE_REG_8__2__SCAN_IN,
         P1_INSTQUEUE_REG_8__1__SCAN_IN, P1_INSTQUEUE_REG_8__0__SCAN_IN,
         P1_INSTQUEUE_REG_7__7__SCAN_IN, P1_INSTQUEUE_REG_7__6__SCAN_IN,
         P1_INSTQUEUE_REG_7__5__SCAN_IN, P1_INSTQUEUE_REG_7__4__SCAN_IN,
         P1_INSTQUEUE_REG_7__3__SCAN_IN, P1_INSTQUEUE_REG_7__2__SCAN_IN,
         P1_INSTQUEUE_REG_7__1__SCAN_IN, P1_INSTQUEUE_REG_7__0__SCAN_IN,
         P1_INSTQUEUE_REG_6__7__SCAN_IN, P1_INSTQUEUE_REG_6__6__SCAN_IN,
         P1_INSTQUEUE_REG_6__5__SCAN_IN, P1_INSTQUEUE_REG_6__4__SCAN_IN,
         P1_INSTQUEUE_REG_6__3__SCAN_IN, P1_INSTQUEUE_REG_6__2__SCAN_IN,
         P1_INSTQUEUE_REG_6__1__SCAN_IN, P1_INSTQUEUE_REG_6__0__SCAN_IN,
         P1_INSTQUEUE_REG_5__7__SCAN_IN, P1_INSTQUEUE_REG_5__6__SCAN_IN,
         P1_INSTQUEUE_REG_5__5__SCAN_IN, P1_INSTQUEUE_REG_5__4__SCAN_IN,
         P1_INSTQUEUE_REG_5__3__SCAN_IN, P1_INSTQUEUE_REG_5__2__SCAN_IN,
         P1_INSTQUEUE_REG_5__1__SCAN_IN, P1_INSTQUEUE_REG_5__0__SCAN_IN,
         P1_INSTQUEUE_REG_4__7__SCAN_IN, P1_INSTQUEUE_REG_4__6__SCAN_IN,
         P1_INSTQUEUE_REG_4__5__SCAN_IN, P1_INSTQUEUE_REG_4__4__SCAN_IN,
         P1_INSTQUEUE_REG_4__3__SCAN_IN, P1_INSTQUEUE_REG_4__2__SCAN_IN,
         P1_INSTQUEUE_REG_4__1__SCAN_IN, keyinput0, keyinput1, keyinput2,
         keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, keyinput8,
         keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, keyinput14,
         keyinput15, keyinput16, keyinput17, keyinput18, keyinput19,
         keyinput20, keyinput21, keyinput22, keyinput23, keyinput24,
         keyinput25, keyinput26, keyinput27, keyinput28, keyinput29,
         keyinput30, keyinput31, keyinput32, keyinput33, keyinput34,
         keyinput35, keyinput36, keyinput37, keyinput38, keyinput39,
         keyinput40, keyinput41, keyinput42, keyinput43, keyinput44,
         keyinput45, keyinput46, keyinput47, keyinput48, keyinput49,
         keyinput50, keyinput51, keyinput52, keyinput53, keyinput54,
         keyinput55, keyinput56, keyinput57, keyinput58, keyinput59,
         keyinput60, keyinput61, keyinput62, keyinput63, keyinput64,
         keyinput65, keyinput66, keyinput67, keyinput68, keyinput69,
         keyinput70, keyinput71, keyinput72, keyinput73, keyinput74,
         keyinput75, keyinput76, keyinput77, keyinput78, keyinput79,
         keyinput80, keyinput81, keyinput82, keyinput83, keyinput84,
         keyinput85, keyinput86, keyinput87, keyinput88, keyinput89,
         keyinput90, keyinput91, keyinput92, keyinput93, keyinput94,
         keyinput95, keyinput96, keyinput97, keyinput98, keyinput99,
         keyinput100, keyinput101, keyinput102, keyinput103, keyinput104,
         keyinput105, keyinput106, keyinput107, keyinput108, keyinput109,
         keyinput110, keyinput111, keyinput112, keyinput113, keyinput114,
         keyinput115, keyinput116, keyinput117, keyinput118, keyinput119,
         keyinput120, keyinput121, keyinput122, keyinput123, keyinput124,
         keyinput125, keyinput126, keyinput127, keyinput128, keyinput129,
         keyinput130, keyinput131, keyinput132, keyinput133, keyinput134,
         keyinput135, keyinput136, keyinput137, keyinput138, keyinput139,
         keyinput140, keyinput141, keyinput142, keyinput143, keyinput144,
         keyinput145, keyinput146, keyinput147, keyinput148, keyinput149,
         keyinput150, keyinput151, keyinput152, keyinput153, keyinput154,
         keyinput155, keyinput156, keyinput157, keyinput158, keyinput159,
         keyinput160, keyinput161, keyinput162, keyinput163, keyinput164,
         keyinput165, keyinput166, keyinput167, keyinput168, keyinput169,
         keyinput170, keyinput171, keyinput172, keyinput173, keyinput174,
         keyinput175, keyinput176, keyinput177, keyinput178, keyinput179,
         keyinput180, keyinput181, keyinput182, keyinput183, keyinput184,
         keyinput185, keyinput186, keyinput187, keyinput188, keyinput189,
         keyinput190, keyinput191, keyinput192, keyinput193, keyinput194,
         keyinput195, keyinput196, keyinput197, keyinput198, keyinput199,
         keyinput200, keyinput201, keyinput202, keyinput203, keyinput204,
         keyinput205, keyinput206, keyinput207, keyinput208, keyinput209,
         keyinput210, keyinput211, keyinput212, keyinput213, keyinput214,
         keyinput215, keyinput216, keyinput217, keyinput218, keyinput219,
         keyinput220, keyinput221, keyinput222, keyinput223, keyinput224,
         keyinput225, keyinput226, keyinput227, keyinput228, keyinput229,
         keyinput230, keyinput231, keyinput232, keyinput233, keyinput234,
         keyinput235, keyinput236, keyinput237, keyinput238, keyinput239,
         keyinput240, keyinput241, keyinput242, keyinput243, keyinput244,
         keyinput245, keyinput246, keyinput247, keyinput248, keyinput249,
         keyinput250, keyinput251, keyinput252, keyinput253, keyinput254,
         keyinput255;
  output U355, U356, U357, U358, U359, U360, U361, U362, U363, U364, U366,
         U367, U368, U369, U370, U371, U372, U373, U374, U375, U347, U348,
         U349, U350, U351, U352, U353, U354, U365, U376, U247, U246, U245,
         U244, U243, U242, U241, U240, U239, U238, U237, U236, U235, U234,
         U233, U232, U231, U230, U229, U228, U227, U226, U225, U224, U223,
         U222, U221, U220, U219, U218, U217, U216, U251, U252, U253, U254,
         U255, U256, U257, U258, U259, U260, U261, U262, U263, U264, U265,
         U266, U267, U268, U269, U270, U271, U272, U273, U274, U275, U276,
         U277, U278, U279, U280, U281, U282, U212, U215, U213, U214, P3_U3274,
         P3_U3275, P3_U3276, P3_U3277, P3_U3061, P3_U3060, P3_U3059, P3_U3058,
         P3_U3057, P3_U3056, P3_U3055, P3_U3054, P3_U3053, P3_U3052, P3_U3051,
         P3_U3050, P3_U3049, P3_U3048, P3_U3047, P3_U3046, P3_U3045, P3_U3044,
         P3_U3043, P3_U3042, P3_U3041, P3_U3040, P3_U3039, P3_U3038, P3_U3037,
         P3_U3036, P3_U3035, P3_U3034, P3_U3033, P3_U3032, P3_U3031, P3_U3030,
         P3_U3029, P3_U3280, P3_U3281, P3_U3028, P3_U3027, P3_U3026, P3_U3025,
         P3_U3024, P3_U3023, P3_U3022, P3_U3021, P3_U3020, P3_U3019, P3_U3018,
         P3_U3017, P3_U3016, P3_U3015, P3_U3014, P3_U3013, P3_U3012, P3_U3011,
         P3_U3010, P3_U3009, P3_U3008, P3_U3007, P3_U3006, P3_U3005, P3_U3004,
         P3_U3003, P3_U3002, P3_U3001, P3_U3000, P3_U2999, P3_U3282, P3_U2998,
         P3_U2997, P3_U2996, P3_U2995, P3_U2994, P3_U2993, P3_U2992, P3_U2991,
         P3_U2990, P3_U2989, P3_U2988, P3_U2987, P3_U2986, P3_U2985, P3_U2984,
         P3_U2983, P3_U2982, P3_U2981, P3_U2980, P3_U2979, P3_U2978, P3_U2977,
         P3_U2976, P3_U2975, P3_U2974, P3_U2973, P3_U2972, P3_U2971, P3_U2970,
         P3_U2969, P3_U2968, P3_U2967, P3_U2966, P3_U2965, P3_U2964, P3_U2963,
         P3_U2962, P3_U2961, P3_U2960, P3_U2959, P3_U2958, P3_U2957, P3_U2956,
         P3_U2955, P3_U2954, P3_U2953, P3_U2952, P3_U2951, P3_U2950, P3_U2949,
         P3_U2948, P3_U2947, P3_U2946, P3_U2945, P3_U2944, P3_U2943, P3_U2942,
         P3_U2941, P3_U2940, P3_U2939, P3_U2938, P3_U2937, P3_U2936, P3_U2935,
         P3_U2934, P3_U2933, P3_U2932, P3_U2931, P3_U2930, P3_U2929, P3_U2928,
         P3_U2927, P3_U2926, P3_U2925, P3_U2924, P3_U2923, P3_U2922, P3_U2921,
         P3_U2920, P3_U2919, P3_U2918, P3_U2917, P3_U2916, P3_U2915, P3_U2914,
         P3_U2913, P3_U2912, P3_U2911, P3_U2910, P3_U2909, P3_U2908, P3_U2907,
         P3_U2906, P3_U2905, P3_U2904, P3_U2903, P3_U2902, P3_U2901, P3_U2900,
         P3_U2899, P3_U2898, P3_U2897, P3_U2896, P3_U2895, P3_U2894, P3_U2893,
         P3_U2892, P3_U2891, P3_U2890, P3_U2889, P3_U2888, P3_U2887, P3_U2886,
         P3_U2885, P3_U2884, P3_U2883, P3_U2882, P3_U2881, P3_U2880, P3_U2879,
         P3_U2878, P3_U2877, P3_U2876, P3_U2875, P3_U2874, P3_U2873, P3_U2872,
         P3_U2871, P3_U2870, P3_U2869, P3_U2868, P3_U3284, P3_U3285, P3_U3288,
         P3_U3289, P3_U3290, P3_U2867, P3_U2866, P3_U2865, P3_U2864, P3_U2863,
         P3_U2862, P3_U2861, P3_U2860, P3_U2859, P3_U2858, P3_U2857, P3_U2856,
         P3_U2855, P3_U2854, P3_U2853, P3_U2852, P3_U2851, P3_U2850, P3_U2849,
         P3_U2848, P3_U2847, P3_U2846, P3_U2845, P3_U2844, P3_U2843, P3_U2842,
         P3_U2841, P3_U2840, P3_U2839, P3_U2838, P3_U2837, P3_U2836, P3_U2835,
         P3_U2834, P3_U2833, P3_U2832, P3_U2831, P3_U2830, P3_U2829, P3_U2828,
         P3_U2827, P3_U2826, P3_U2825, P3_U2824, P3_U2823, P3_U2822, P3_U2821,
         P3_U2820, P3_U2819, P3_U2818, P3_U2817, P3_U2816, P3_U2815, P3_U2814,
         P3_U2813, P3_U2812, P3_U2811, P3_U2810, P3_U2809, P3_U2808, P3_U2807,
         P3_U2806, P3_U2805, P3_U2804, P3_U2803, P3_U2802, P3_U2801, P3_U2800,
         P3_U2799, P3_U2798, P3_U2797, P3_U2796, P3_U2795, P3_U2794, P3_U2793,
         P3_U2792, P3_U2791, P3_U2790, P3_U2789, P3_U2788, P3_U2787, P3_U2786,
         P3_U2785, P3_U2784, P3_U2783, P3_U2782, P3_U2781, P3_U2780, P3_U2779,
         P3_U2778, P3_U2777, P3_U2776, P3_U2775, P3_U2774, P3_U2773, P3_U2772,
         P3_U2771, P3_U2770, P3_U2769, P3_U2768, P3_U2767, P3_U2766, P3_U2765,
         P3_U2764, P3_U2763, P3_U2762, P3_U2761, P3_U2760, P3_U2759, P3_U2758,
         P3_U2757, P3_U2756, P3_U2755, P3_U2754, P3_U2753, P3_U2752, P3_U2751,
         P3_U2750, P3_U2749, P3_U2748, P3_U2747, P3_U2746, P3_U2745, P3_U2744,
         P3_U2743, P3_U2742, P3_U2741, P3_U2740, P3_U2739, P3_U2738, P3_U2737,
         P3_U2736, P3_U2735, P3_U2734, P3_U2733, P3_U2732, P3_U2731, P3_U2730,
         P3_U2729, P3_U2728, P3_U2727, P3_U2726, P3_U2725, P3_U2724, P3_U2723,
         P3_U2722, P3_U2721, P3_U2720, P3_U2719, P3_U2718, P3_U2717, P3_U2716,
         P3_U2715, P3_U2714, P3_U2713, P3_U2712, P3_U2711, P3_U2710, P3_U2709,
         P3_U2708, P3_U2707, P3_U2706, P3_U2705, P3_U2704, P3_U2703, P3_U2702,
         P3_U2701, P3_U2700, P3_U2699, P3_U2698, P3_U2697, P3_U2696, P3_U2695,
         P3_U2694, P3_U2693, P3_U2692, P3_U2691, P3_U2690, P3_U2689, P3_U2688,
         P3_U2687, P3_U2686, P3_U2685, P3_U2684, P3_U2683, P3_U2682, P3_U2681,
         P3_U2680, P3_U2679, P3_U2678, P3_U2677, P3_U2676, P3_U2675, P3_U2674,
         P3_U2673, P3_U2672, P3_U2671, P3_U2670, P3_U2669, P3_U2668, P3_U2667,
         P3_U2666, P3_U2665, P3_U2664, P3_U2663, P3_U2662, P3_U2661, P3_U2660,
         P3_U2659, P3_U2658, P3_U2657, P3_U2656, P3_U2655, P3_U2654, P3_U2653,
         P3_U2652, P3_U2651, P3_U2650, P3_U2649, P3_U2648, P3_U2647, P3_U2646,
         P3_U2645, P3_U2644, P3_U2643, P3_U2642, P3_U2641, P3_U2640, P3_U2639,
         P3_U3292, P3_U2638, P3_U3293, P3_U3294, P3_U2637, P3_U3295, P3_U2636,
         P3_U3296, P3_U2635, P3_U3297, P3_U2634, P3_U2633, P3_U3298, P3_U3299,
         P2_U3585, P2_U3586, P2_U3587, P2_U3588, P2_U3241, P2_U3240, P2_U3239,
         P2_U3238, P2_U3237, P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232,
         P2_U3231, P2_U3230, P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225,
         P2_U3224, P2_U3223, P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218,
         P2_U3217, P2_U3216, P2_U3215, P2_U3214, P2_U3213, P2_U3212, P2_U3211,
         P2_U3210, P2_U3209, P2_U3591, P2_U3592, P2_U3208, P2_U3207, P2_U3206,
         P2_U3205, P2_U3204, P2_U3203, P2_U3202, P2_U3201, P2_U3200, P2_U3199,
         P2_U3198, P2_U3197, P2_U3196, P2_U3195, P2_U3194, P2_U3193, P2_U3192,
         P2_U3191, P2_U3190, P2_U3189, P2_U3188, P2_U3187, P2_U3186, P2_U3185,
         P2_U3184, P2_U3183, P2_U3182, P2_U3181, P2_U3180, P2_U3179, P2_U3593,
         P2_U3178, P2_U3177, P2_U3176, P2_U3175, P2_U3174, P2_U3173, P2_U3172,
         P2_U3171, P2_U3170, P2_U3169, P2_U3168, P2_U3167, P2_U3166, P2_U3165,
         P2_U3164, P2_U3163, P2_U3162, P2_U3161, P2_U3160, P2_U3159, P2_U3158,
         P2_U3157, P2_U3156, P2_U3155, P2_U3154, P2_U3153, P2_U3152, P2_U3151,
         P2_U3150, P2_U3149, P2_U3148, P2_U3147, P2_U3146, P2_U3145, P2_U3144,
         P2_U3143, P2_U3142, P2_U3141, P2_U3140, P2_U3139, P2_U3138, P2_U3137,
         P2_U3136, P2_U3135, P2_U3134, P2_U3133, P2_U3132, P2_U3131, P2_U3130,
         P2_U3129, P2_U3128, P2_U3127, P2_U3126, P2_U3125, P2_U3124, P2_U3123,
         P2_U3122, P2_U3121, P2_U3120, P2_U3119, P2_U3118, P2_U3117, P2_U3116,
         P2_U3115, P2_U3114, P2_U3113, P2_U3112, P2_U3111, P2_U3110, P2_U3109,
         P2_U3108, P2_U3107, P2_U3106, P2_U3105, P2_U3104, P2_U3103, P2_U3102,
         P2_U3101, P2_U3100, P2_U3099, P2_U3098, P2_U3097, P2_U3096, P2_U3095,
         P2_U3094, P2_U3093, P2_U3092, P2_U3091, P2_U3090, P2_U3089, P2_U3088,
         P2_U3087, P2_U3086, P2_U3085, P2_U3084, P2_U3083, P2_U3082, P2_U3081,
         P2_U3080, P2_U3079, P2_U3078, P2_U3077, P2_U3076, P2_U3075, P2_U3074,
         P2_U3073, P2_U3072, P2_U3071, P2_U3070, P2_U3069, P2_U3068, P2_U3067,
         P2_U3066, P2_U3065, P2_U3064, P2_U3063, P2_U3062, P2_U3061, P2_U3060,
         P2_U3059, P2_U3058, P2_U3057, P2_U3056, P2_U3055, P2_U3054, P2_U3053,
         P2_U3052, P2_U3051, P2_U3050, P2_U3049, P2_U3048, P2_U3595, P2_U3596,
         P2_U3599, P2_U3600, P2_U3601, P2_U3047, P2_U3602, P2_U3603, P2_U3604,
         P2_U3605, P2_U3046, P2_U3045, P2_U3044, P2_U3043, P2_U3042, P2_U3041,
         P2_U3040, P2_U3039, P2_U3038, P2_U3037, P2_U3036, P2_U3035, P2_U3034,
         P2_U3033, P2_U3032, P2_U3031, P2_U3030, P2_U3029, P2_U3028, P2_U3027,
         P2_U3026, P2_U3025, P2_U3024, P2_U3023, P2_U3022, P2_U3021, P2_U3020,
         P2_U3019, P2_U3018, P2_U3017, P2_U3016, P2_U3015, P2_U3014, P2_U3013,
         P2_U3012, P2_U3011, P2_U3010, P2_U3009, P2_U3008, P2_U3007, P2_U3006,
         P2_U3005, P2_U3004, P2_U3003, P2_U3002, P2_U3001, P2_U3000, P2_U2999,
         P2_U2998, P2_U2997, P2_U2996, P2_U2995, P2_U2994, P2_U2993, P2_U2992,
         P2_U2991, P2_U2990, P2_U2989, P2_U2988, P2_U2987, P2_U2986, P2_U2985,
         P2_U2984, P2_U2983, P2_U2982, P2_U2981, P2_U2980, P2_U2979, P2_U2978,
         P2_U2977, P2_U2976, P2_U2975, P2_U2974, P2_U2973, P2_U2972, P2_U2971,
         P2_U2970, P2_U2969, P2_U2968, P2_U2967, P2_U2966, P2_U2965, P2_U2964,
         P2_U2963, P2_U2962, P2_U2961, P2_U2960, P2_U2959, P2_U2958, P2_U2957,
         P2_U2956, P2_U2955, P2_U2954, P2_U2953, P2_U2952, P2_U2951, P2_U2950,
         P2_U2949, P2_U2948, P2_U2947, P2_U2946, P2_U2945, P2_U2944, P2_U2943,
         P2_U2942, P2_U2941, P2_U2940, P2_U2939, P2_U2938, P2_U2937, P2_U2936,
         P2_U2935, P2_U2934, P2_U2933, P2_U2932, P2_U2931, P2_U2930, P2_U2929,
         P2_U2928, P2_U2927, P2_U2926, P2_U2925, P2_U2924, P2_U2923, P2_U2922,
         P2_U2921, P2_U2920, P2_U2919, P2_U2918, P2_U2917, P2_U2916, P2_U2915,
         P2_U2914, P2_U2913, P2_U2912, P2_U2911, P2_U2910, P2_U2909, P2_U2908,
         P2_U2907, P2_U2906, P2_U2905, P2_U2904, P2_U2903, P2_U2902, P2_U2901,
         P2_U2900, P2_U2899, P2_U2898, P2_U2897, P2_U2896, P2_U2895, P2_U2894,
         P2_U2893, P2_U2892, P2_U2891, P2_U2890, P2_U2889, P2_U2888, P2_U2887,
         P2_U2886, P2_U2885, P2_U2884, P2_U2883, P2_U2882, P2_U2881, P2_U2880,
         P2_U2879, P2_U2878, P2_U2877, P2_U2876, P2_U2875, P2_U2874, P2_U2873,
         P2_U2872, P2_U2871, P2_U2870, P2_U2869, P2_U2868, P2_U2867, P2_U2866,
         P2_U2865, P2_U2864, P2_U2863, P2_U2862, P2_U2861, P2_U2860, P2_U2859,
         P2_U2858, P2_U2857, P2_U2856, P2_U2855, P2_U2854, P2_U2853, P2_U2852,
         P2_U2851, P2_U2850, P2_U2849, P2_U2848, P2_U2847, P2_U2846, P2_U2845,
         P2_U2844, P2_U2843, P2_U2842, P2_U2841, P2_U2840, P2_U2839, P2_U2838,
         P2_U2837, P2_U2836, P2_U2835, P2_U2834, P2_U2833, P2_U2832, P2_U2831,
         P2_U2830, P2_U2829, P2_U2828, P2_U2827, P2_U2826, P2_U2825, P2_U2824,
         P2_U2823, P2_U2822, P2_U2821, P2_U2820, P2_U3608, P2_U2819, P2_U3609,
         P2_U2818, P2_U3610, P2_U2817, P2_U3611, P2_U2816, P2_U2815, P2_U3612,
         P2_U2814, P1_U3458, P1_U3459, P1_U3460, P1_U3461, P1_U3226, P1_U3225,
         P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218,
         P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211,
         P1_U3210, P1_U3209, P1_U3208, P1_U3207, P1_U3206, P1_U3205, P1_U3204,
         P1_U3203, P1_U3202, P1_U3201, P1_U3200, P1_U3199, P1_U3198, P1_U3197,
         P1_U3196, P1_U3195, P1_U3194, P1_U3464, P1_U3465, P1_U3193, P1_U3192,
         P1_U3191, P1_U3190, P1_U3189, P1_U3188, P1_U3187, P1_U3186, P1_U3185,
         P1_U3184, P1_U3183, P1_U3182, P1_U3181, P1_U3180, P1_U3179, P1_U3178,
         P1_U3177, P1_U3176, P1_U3175, P1_U3174, P1_U3173, P1_U3172, P1_U3171,
         P1_U3170, P1_U3169, P1_U3168, P1_U3167, P1_U3166, P1_U3165, P1_U3164,
         P1_U3466, P1_U3163, P1_U3162, P1_U3161, P1_U3160, P1_U3159, P1_U3158,
         P1_U3157, P1_U3156, P1_U3155, P1_U3154, P1_U3153, P1_U3152, P1_U3151,
         P1_U3150, P1_U3149, P1_U3148, P1_U3147, P1_U3146, P1_U3145, P1_U3144,
         P1_U3143, P1_U3142, P1_U3141, P1_U3140, P1_U3139, P1_U3138, P1_U3137,
         P1_U3136, P1_U3135, P1_U3134, P1_U3133, P1_U3132, P1_U3131, P1_U3130,
         P1_U3129, P1_U3128, P1_U3127, P1_U3126, P1_U3125, P1_U3124, P1_U3123,
         P1_U3122, P1_U3121, P1_U3120, P1_U3119, P1_U3118, P1_U3117, P1_U3116,
         P1_U3115, P1_U3114, P1_U3113, P1_U3112, P1_U3111, P1_U3110, P1_U3109,
         P1_U3108, P1_U3107, P1_U3106, P1_U3105, P1_U3104, P1_U3103, P1_U3102,
         P1_U3101, P1_U3100, P1_U3099, P1_U3098, P1_U3097, P1_U3096, P1_U3095,
         P1_U3094, P1_U3093, P1_U3092, P1_U3091, P1_U3090, P1_U3089, P1_U3088,
         P1_U3087, P1_U3086, P1_U3085, P1_U3084, P1_U3083, P1_U3082, P1_U3081,
         P1_U3080, P1_U3079, P1_U3078, P1_U3077, P1_U3076, P1_U3075, P1_U3074,
         P1_U3073, P1_U3072, P1_U3071, P1_U3070, P1_U3069, P1_U3068, P1_U3067,
         P1_U3066, P1_U3065, P1_U3064, P1_U3063, P1_U3062, P1_U3061, P1_U3060,
         P1_U3059, P1_U3058, P1_U3057, P1_U3056, P1_U3055, P1_U3054, P1_U3053,
         P1_U3052, P1_U3051, P1_U3050, P1_U3049, P1_U3048, P1_U3047, P1_U3046,
         P1_U3045, P1_U3044, P1_U3043, P1_U3042, P1_U3041, P1_U3040, P1_U3039,
         P1_U3038, P1_U3037, P1_U3036, P1_U3035, P1_U3034, P1_U3033, P1_U3468,
         P1_U3469, P1_U3472, P1_U3473, P1_U3474, P1_U3032, P1_U3475, P1_U3476,
         P1_U3477, P1_U3478, P1_U3031, P1_U3030, P1_U3029, P1_U3028, P1_U3027,
         P1_U3026, P1_U3025, P1_U3024, P1_U3023, P1_U3022, P1_U3021, P1_U3020,
         P1_U3019, P1_U3018, P1_U3017, P1_U3016, P1_U3015, P1_U3014, P1_U3013,
         P1_U3012, P1_U3011, P1_U3010, P1_U3009, P1_U3008, P1_U3007, P1_U3006,
         P1_U3005, P1_U3004, P1_U3003, P1_U3002, P1_U3001, P1_U3000, P1_U2999,
         P1_U2998, P1_U2997, P1_U2996, P1_U2995, P1_U2994, P1_U2993, P1_U2992,
         P1_U2991, P1_U2990, P1_U2989, P1_U2988, P1_U2987, P1_U2986, P1_U2985,
         P1_U2984, P1_U2983, P1_U2982, P1_U2981, P1_U2980, P1_U2979, P1_U2978,
         P1_U2977, P1_U2976, P1_U2975, P1_U2974, P1_U2973, P1_U2972, P1_U2971,
         P1_U2970, P1_U2969, P1_U2968, P1_U2967, P1_U2966, P1_U2965, P1_U2964,
         P1_U2963, P1_U2962, P1_U2961, P1_U2960, P1_U2959, P1_U2958, P1_U2957,
         P1_U2956, P1_U2955, P1_U2954, P1_U2953, P1_U2952, P1_U2951, P1_U2950,
         P1_U2949, P1_U2948, P1_U2947, P1_U2946, P1_U2945, P1_U2944, P1_U2943,
         P1_U2942, P1_U2941, P1_U2940, P1_U2939, P1_U2938, P1_U2937, P1_U2936,
         P1_U2935, P1_U2934, P1_U2933, P1_U2932, P1_U2931, P1_U2930, P1_U2929,
         P1_U2928, P1_U2927, P1_U2926, P1_U2925, P1_U2924, P1_U2923, P1_U2922,
         P1_U2921, P1_U2920, P1_U2919, P1_U2918, P1_U2917, P1_U2916, P1_U2915,
         P1_U2914, P1_U2913, P1_U2912, P1_U2911, P1_U2910, P1_U2909, P1_U2908,
         P1_U2907, P1_U2906, P1_U2905, P1_U2904, P1_U2903, P1_U2902, P1_U2901,
         P1_U2900, P1_U2899, P1_U2898, P1_U2897, P1_U2896, P1_U2895, P1_U2894,
         P1_U2893, P1_U2892, P1_U2891, P1_U2890, P1_U2889, P1_U2888, P1_U2887,
         P1_U2886, P1_U2885, P1_U2884, P1_U2883, P1_U2882, P1_U2881, P1_U2880,
         P1_U2879, P1_U2878, P1_U2877, P1_U2876, P1_U2875, P1_U2874, P1_U2873,
         P1_U2872, P1_U2871, P1_U2870, P1_U2869, P1_U2868, P1_U2867, P1_U2866,
         P1_U2865, P1_U2864, P1_U2863, P1_U2862, P1_U2861, P1_U2860, P1_U2859,
         P1_U2858, P1_U2857, P1_U2856, P1_U2855, P1_U2854, P1_U2853, P1_U2852,
         P1_U2851, P1_U2850, P1_U2849, P1_U2848, P1_U2847, P1_U2846, P1_U2845,
         P1_U2844, P1_U2843, P1_U2842, P1_U2841, P1_U2840, P1_U2839, P1_U2838,
         P1_U2837, P1_U2836, P1_U2835, P1_U2834, P1_U2833, P1_U2832, P1_U2831,
         P1_U2830, P1_U2829, P1_U2828, P1_U2827, P1_U2826, P1_U2825, P1_U2824,
         P1_U2823, P1_U2822, P1_U2821, P1_U2820, P1_U2819, P1_U2818, P1_U2817,
         P1_U2816, P1_U2815, P1_U2814, P1_U2813, P1_U2812, P1_U2811, P1_U2810,
         P1_U2809, P1_U2808, P1_U3481, P1_U2807, P1_U3482, P1_U3483, P1_U2806,
         P1_U3484, P1_U2805, P1_U3485, P1_U2804, P1_U3486, P1_U2803, P1_U2802,
         P1_U3487, P1_U2801;
  wire   n9805, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9815, n9816,
         n9817, n9818, n9819, n9820, n9822, n9823, n9824, n9825, n9826, n9827,
         n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,
         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,
         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,
         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,
         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,
         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,
         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,
         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,
         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,
         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,
         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,
         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,
         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,
         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,
         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,
         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,
         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,
         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,
         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,
         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,
         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,
         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,
         n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
         n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,
         n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,
         n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,
         n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
         n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,
         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,
         n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
         n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,
         n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,
         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
         n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,
         n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
         n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
         n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,
         n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,
         n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176,
         n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,
         n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
         n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,
         n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208,
         n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
         n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,
         n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248,
         n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256,
         n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
         n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272,
         n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280,
         n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
         n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296,
         n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304,
         n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312,
         n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320,
         n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328,
         n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
         n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344,
         n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352,
         n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
         n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368,
         n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376,
         n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384,
         n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392,
         n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400,
         n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,
         n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416,
         n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424,
         n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
         n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440,
         n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
         n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456,
         n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464,
         n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472,
         n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
         n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488,
         n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
         n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,
         n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512,
         n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520,
         n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528,
         n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
         n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
         n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
         n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560,
         n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
         n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
         n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584,
         n19585, n19586, n19587, n19588, n19589, n19590, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19690,
         n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698,
         n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
         n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
         n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722,
         n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730,
         n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
         n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746,
         n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754,
         n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762,
         n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770,
         n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
         n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
         n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794,
         n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802,
         n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
         n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818,
         n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
         n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834,
         n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
         n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
         n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
         n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906,
         n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914,
         n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
         n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
         n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938,
         n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
         n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954,
         n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962,
         n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970,
         n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978,
         n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986,
         n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
         n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
         n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
         n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018,
         n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
         n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034,
         n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
         n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
         n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
         n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
         n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
         n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
         n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
         n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
         n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
         n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
         n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
         n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162,
         n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
         n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178,
         n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
         n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
         n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202,
         n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
         n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
         n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226,
         n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250,
         n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
         n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
         n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274,
         n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282,
         n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
         n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298,
         n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306,
         n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314,
         n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322,
         n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
         n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338,
         n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
         n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
         n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
         n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370,
         n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378,
         n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
         n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
         n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
         n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
         n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
         n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
         n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
         n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442,
         n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450,
         n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
         n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
         n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
         n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482,
         n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490,
         n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
         n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
         n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514,
         n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
         n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
         n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
         n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
         n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554,
         n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562,
         n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
         n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
         n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
         n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610,
         n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
         n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626,
         n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634,
         n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
         n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
         n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
         n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
         n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
         n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
         n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
         n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
         n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
         n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754,
         n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
         n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770,
         n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778,
         n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
         n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
         n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
         n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
         n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
         n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
         n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842,
         n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
         n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
         n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
         n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874,
         n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
         n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
         n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
         n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
         n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946,
         n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
         n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
         n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970,
         n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
         n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986,
         n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994,
         n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
         n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
         n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018,
         n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026,
         n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034,
         n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
         n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050,
         n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058,
         n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066,
         n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074,
         n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082,
         n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090,
         n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098,
         n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106,
         n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114,
         n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122,
         n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130,
         n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138,
         n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146,
         n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154,
         n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162,
         n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170,
         n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178,
         n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186,
         n21187, n21188, n21189, n21190, n21191, n21192;

  INV_X1 U11249 ( .A(n19941), .ZN(n19953) );
  AND2_X1 U11250 ( .A1(n9988), .A2(n9987), .ZN(n15095) );
  OR2_X1 U11251 ( .A1(n10828), .A2(n10827), .ZN(n15131) );
  AOI21_X1 U11252 ( .B1(n13503), .B2(n13501), .A(n12886), .ZN(n13508) );
  INV_X1 U11253 ( .A(n12695), .ZN(n12845) );
  CLKBUF_X2 U11254 ( .A(n10468), .Z(n12622) );
  INV_X1 U11255 ( .A(n12868), .ZN(n14914) );
  AND2_X1 U11256 ( .A1(n10527), .A2(n10521), .ZN(n19647) );
  OAI22_X1 U11257 ( .A1(n13654), .A2(P1_STATE2_REG_0__SCAN_IN), .B1(n11262), 
        .B2(n11278), .ZN(n11255) );
  OAI211_X1 U11258 ( .C1(n11233), .C2(n10036), .A(n10035), .B(n10031), .ZN(
        n13654) );
  CLKBUF_X1 U11259 ( .A(n11858), .Z(n17034) );
  AND2_X1 U11260 ( .A1(n10540), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12952) );
  AND2_X1 U11261 ( .A1(n9827), .A2(n16232), .ZN(n10690) );
  CLKBUF_X2 U11263 ( .A(n11677), .Z(n9815) );
  CLKBUF_X2 U11264 ( .A(n11806), .Z(n9813) );
  CLKBUF_X2 U11265 ( .A(n11677), .Z(n9816) );
  CLKBUF_X3 U11266 ( .A(n11805), .Z(n9818) );
  CLKBUF_X1 U11267 ( .A(n11110), .Z(n12458) );
  CLKBUF_X2 U11269 ( .A(n11147), .Z(n12275) );
  CLKBUF_X2 U11270 ( .A(n11098), .Z(n12466) );
  CLKBUF_X2 U11271 ( .A(n12465), .Z(n9831) );
  NAND2_X1 U11273 ( .A1(n10423), .A2(n12658), .ZN(n10472) );
  INV_X1 U11274 ( .A(n20122), .ZN(n13281) );
  CLKBUF_X2 U11275 ( .A(n10447), .Z(n16281) );
  AND4_X1 U11276 ( .A1(n11102), .A2(n11101), .A3(n11100), .A4(n11099), .ZN(
        n10313) );
  NAND2_X2 U11277 ( .A1(n10385), .A2(n10386), .ZN(n10443) );
  AND2_X1 U11278 ( .A1(n11004), .A2(n13673), .ZN(n11194) );
  AND2_X2 U11279 ( .A1(n11006), .A2(n11005), .ZN(n11245) );
  AND2_X2 U11280 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13672) );
  AND3_X2 U11281 ( .A1(n9959), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n9825) );
  CLKBUF_X1 U11282 ( .A(n18599), .Z(n9805) );
  NOR2_X1 U11283 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n18696), .ZN(n18599) );
  INV_X1 U11285 ( .A(n21192), .ZN(n9807) );
  AND2_X1 U11286 ( .A1(n10999), .A2(n13667), .ZN(n11098) );
  CLKBUF_X2 U11287 ( .A(n11194), .Z(n11167) );
  NAND2_X1 U11288 ( .A1(n11188), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n11228) );
  AND3_X1 U11289 ( .A1(n10594), .A2(n10593), .A3(n10592), .ZN(n10307) );
  AND2_X1 U11290 ( .A1(n12659), .A2(n10426), .ZN(n10423) );
  AND2_X1 U11291 ( .A1(n10353), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10572) );
  AND3_X1 U11292 ( .A1(n10438), .A2(n10437), .A3(n19838), .ZN(n12643) );
  AOI22_X1 U11293 ( .A1(n21101), .A2(keyinput44), .B1(keyinput120), .B2(n21100), .ZN(n21099) );
  INV_X1 U11294 ( .A(n11108), .ZN(n11491) );
  NAND2_X1 U11295 ( .A1(n10801), .A2(n10146), .ZN(n10809) );
  INV_X1 U11296 ( .A(n12710), .ZN(n12841) );
  OR3_X1 U11297 ( .A1(n16062), .A2(n15176), .A3(n15120), .ZN(n10829) );
  NAND4_X1 U11298 ( .A1(n10636), .A2(n10635), .A3(n10634), .A4(n10633), .ZN(
        n15187) );
  CLKBUF_X2 U11299 ( .A(n11806), .Z(n9812) );
  INV_X1 U11300 ( .A(n15611), .ZN(n17049) );
  INV_X1 U11301 ( .A(n18568), .ZN(n18549) );
  OAI221_X1 U11302 ( .B1(n21101), .B2(keyinput44), .C1(n21100), .C2(
        keyinput120), .A(n21099), .ZN(n21106) );
  NOR2_X1 U11303 ( .A1(n11501), .A2(n20122), .ZN(n13265) );
  INV_X1 U11304 ( .A(n11588), .ZN(n13516) );
  NAND2_X1 U11305 ( .A1(n14058), .A2(n14123), .ZN(n14122) );
  NOR2_X2 U11306 ( .A1(n10809), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10815) );
  BUF_X1 U11307 ( .A(n12571), .Z(n9839) );
  OR2_X1 U11308 ( .A1(n9977), .A2(n9976), .ZN(n9975) );
  NOR2_X1 U11309 ( .A1(n15110), .A2(n21005), .ZN(n15112) );
  AND2_X1 U11310 ( .A1(n12875), .A2(n12885), .ZN(n13503) );
  NAND2_X1 U11311 ( .A1(n10398), .A2(n10397), .ZN(n10427) );
  AND2_X1 U11312 ( .A1(n16567), .A2(n16797), .ZN(n16558) );
  INV_X1 U11313 ( .A(n11825), .ZN(n11658) );
  INV_X1 U11314 ( .A(n11500), .ZN(n12493) );
  AND2_X1 U11316 ( .A1(n14101), .A2(n9930), .ZN(n14998) );
  NAND2_X1 U11317 ( .A1(n10254), .A2(n10255), .ZN(n14100) );
  AND3_X1 U11318 ( .A1(n9970), .A2(n9969), .A3(n9968), .ZN(n9857) );
  INV_X1 U11319 ( .A(n17153), .ZN(n18134) );
  INV_X1 U11320 ( .A(n17598), .ZN(n17575) );
  INV_X1 U11321 ( .A(n17652), .ZN(n17579) );
  INV_X1 U11322 ( .A(n14069), .ZN(n14070) );
  INV_X1 U11323 ( .A(n19908), .ZN(n15796) );
  NOR2_X2 U11324 ( .A1(n17197), .A2(n17365), .ZN(n17191) );
  INV_X2 U11325 ( .A(n15667), .ZN(n11979) );
  NAND2_X1 U11326 ( .A1(n12498), .A2(n20122), .ZN(n14432) );
  AND2_X2 U11327 ( .A1(n10546), .A2(n10315), .ZN(n9808) );
  NAND2_X1 U11328 ( .A1(n14588), .A2(n15859), .ZN(n14575) );
  NAND2_X2 U11329 ( .A1(n16797), .A2(n10185), .ZN(n10184) );
  INV_X1 U11330 ( .A(n11812), .ZN(n9809) );
  INV_X1 U11331 ( .A(n11812), .ZN(n9810) );
  NOR2_X2 U11332 ( .A1(n11648), .A2(n11647), .ZN(n11857) );
  AND2_X4 U11333 ( .A1(n15542), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n10539) );
  NAND2_X2 U11334 ( .A1(n15140), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15119) );
  NOR2_X2 U11335 ( .A1(n14211), .A2(n9873), .ZN(n15140) );
  NOR2_X2 U11336 ( .A1(n14990), .A2(n14989), .ZN(n14988) );
  INV_X2 U11337 ( .A(n11658), .ZN(n9811) );
  NOR2_X1 U11338 ( .A1(n18563), .A2(n11639), .ZN(n11825) );
  AOI21_X2 U11339 ( .B1(n15374), .B2(n15217), .A(n15211), .ZN(n15376) );
  INV_X2 U11340 ( .A(n15195), .ZN(n15211) );
  NOR2_X1 U11342 ( .A1(n11649), .A2(n16793), .ZN(n11806) );
  OR2_X1 U11343 ( .A1(n14964), .A2(n14963), .ZN(n13083) );
  NAND2_X1 U11344 ( .A1(n10011), .A2(n10013), .ZN(n14685) );
  NOR2_X1 U11345 ( .A1(n14663), .A2(n15875), .ZN(n11404) );
  AND2_X1 U11346 ( .A1(n10038), .A2(n10012), .ZN(n10011) );
  NOR2_X1 U11347 ( .A1(n13637), .A2(n19156), .ZN(n13576) );
  NAND2_X1 U11348 ( .A1(n12889), .A2(n12888), .ZN(n13637) );
  INV_X4 U11349 ( .A(n14636), .ZN(n14688) );
  NOR2_X1 U11350 ( .A1(n18696), .A2(n16796), .ZN(n16754) );
  BUF_X1 U11351 ( .A(n11996), .Z(n9828) );
  CLKBUF_X2 U11352 ( .A(n10913), .Z(n9847) );
  INV_X1 U11353 ( .A(n18100), .ZN(n16313) );
  NAND2_X1 U11354 ( .A1(n15746), .A2(n17250), .ZN(n11953) );
  OR2_X1 U11355 ( .A1(n11686), .A2(n10078), .ZN(n17153) );
  NOR2_X1 U11356 ( .A1(n11707), .A2(n11706), .ZN(n18123) );
  NOR2_X1 U11357 ( .A1(n11802), .A2(n11801), .ZN(n17240) );
  INV_X2 U11359 ( .A(n10427), .ZN(n9817) );
  AND4_X1 U11360 ( .A1(n11003), .A2(n11002), .A3(n11001), .A4(n11000), .ZN(
        n11012) );
  CLKBUF_X2 U11361 ( .A(n11245), .Z(n12459) );
  CLKBUF_X2 U11362 ( .A(n11240), .Z(n11146) );
  BUF_X2 U11363 ( .A(n11299), .Z(n12440) );
  CLKBUF_X2 U11364 ( .A(n11356), .Z(n12299) );
  CLKBUF_X2 U11365 ( .A(n11193), .Z(n11154) );
  CLKBUF_X1 U11367 ( .A(n15560), .Z(n9841) );
  CLKBUF_X2 U11369 ( .A(n15560), .Z(n9822) );
  CLKBUF_X2 U11370 ( .A(n11691), .Z(n17048) );
  BUF_X1 U11371 ( .A(n11805), .Z(n9838) );
  CLKBUF_X2 U11372 ( .A(n11283), .Z(n11152) );
  BUF_X2 U11373 ( .A(n11153), .Z(n12460) );
  CLKBUF_X2 U11374 ( .A(n11246), .Z(n11155) );
  INV_X2 U11376 ( .A(n18074), .ZN(n9820) );
  INV_X2 U11378 ( .A(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11640) );
  INV_X4 U11379 ( .A(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18720) );
  INV_X2 U11380 ( .A(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n18727) );
  INV_X2 U11381 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n15554) );
  OAI21_X1 U11382 ( .B1(n12553), .B2(n12552), .A(n10309), .ZN(n12559) );
  XNOR2_X1 U11383 ( .A(n15192), .B(n15191), .ZN(n15351) );
  NAND2_X1 U11384 ( .A1(n9975), .A2(n9973), .ZN(n9969) );
  NAND2_X1 U11385 ( .A1(n9971), .A2(n9891), .ZN(n9970) );
  NAND2_X1 U11386 ( .A1(n10065), .A2(n10063), .ZN(n15366) );
  AND2_X1 U11387 ( .A1(n10242), .A2(n10241), .ZN(n14940) );
  AOI21_X1 U11388 ( .B1(n14352), .B2(n14359), .A(n14351), .ZN(n14599) );
  OR2_X1 U11389 ( .A1(n15219), .A2(n15183), .ZN(n10065) );
  NAND2_X1 U11390 ( .A1(n14590), .A2(n14699), .ZN(n14296) );
  NOR2_X1 U11391 ( .A1(n14590), .A2(n11413), .ZN(n14297) );
  NAND2_X1 U11392 ( .A1(n10021), .A2(n14603), .ZN(n14590) );
  NAND2_X1 U11393 ( .A1(n10240), .A2(n13111), .ZN(n10244) );
  OAI21_X1 U11394 ( .B1(n15251), .B2(n10049), .A(n10047), .ZN(n15182) );
  NAND2_X1 U11395 ( .A1(n10022), .A2(n10296), .ZN(n10021) );
  NOR2_X1 U11396 ( .A1(n14617), .A2(n10298), .ZN(n14578) );
  NAND2_X1 U11397 ( .A1(n15175), .A2(n16133), .ZN(n15251) );
  NAND2_X1 U11398 ( .A1(n13083), .A2(n13082), .ZN(n13113) );
  AOI211_X1 U11399 ( .C1(n16013), .C2(n16219), .A(n12858), .B(n12857), .ZN(
        n12859) );
  NAND2_X1 U11400 ( .A1(n15860), .A2(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n14588) );
  NAND2_X1 U11401 ( .A1(n14968), .A2(n13059), .ZN(n13081) );
  OAI21_X1 U11402 ( .B1(n10026), .B2(n10023), .A(n10206), .ZN(n10095) );
  AND2_X1 U11403 ( .A1(n14960), .A2(n14953), .ZN(n14947) );
  NOR2_X1 U11404 ( .A1(n14973), .A2(n14959), .ZN(n14960) );
  NOR2_X1 U11405 ( .A1(n14651), .A2(n11550), .ZN(n10023) );
  OR2_X1 U11406 ( .A1(n14651), .A2(n11550), .ZN(n10024) );
  NAND3_X1 U11407 ( .A1(n14685), .A2(n11404), .A3(n10209), .ZN(n14651) );
  OAI21_X1 U11408 ( .B1(n10275), .B2(n10060), .A(n10058), .ZN(n15452) );
  OR2_X1 U11409 ( .A1(n14985), .A2(n14971), .ZN(n14973) );
  OR2_X1 U11410 ( .A1(n10884), .A2(n10883), .ZN(n10886) );
  XNOR2_X1 U11411 ( .A(n10884), .B(n15176), .ZN(n14078) );
  OR2_X1 U11412 ( .A1(n12537), .A2(n12536), .ZN(n12554) );
  OR2_X1 U11413 ( .A1(n17418), .A2(n11896), .ZN(n11897) );
  OR2_X1 U11414 ( .A1(n10826), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15132) );
  AND2_X1 U11415 ( .A1(n10831), .A2(n10830), .ZN(n12534) );
  AND2_X1 U11416 ( .A1(n11394), .A2(n10016), .ZN(n10015) );
  AND2_X1 U11417 ( .A1(n11396), .A2(n10039), .ZN(n10038) );
  NOR2_X1 U11418 ( .A1(n19789), .A2(n19318), .ZN(n19372) );
  INV_X1 U11419 ( .A(n10824), .ZN(n10831) );
  NOR2_X1 U11420 ( .A1(n14662), .A2(n15872), .ZN(n11407) );
  OR3_X1 U11421 ( .A1(n14679), .A2(n14673), .A3(n14677), .ZN(n14812) );
  NOR2_X1 U11422 ( .A1(n10816), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10820) );
  OR2_X1 U11423 ( .A1(n13952), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11394) );
  INV_X1 U11424 ( .A(n17489), .ZN(n17502) );
  OR2_X1 U11425 ( .A1(n15680), .A2(n15176), .ZN(n10804) );
  AND3_X1 U11426 ( .A1(n13506), .A2(n12866), .A3(n13334), .ZN(n12889) );
  AOI21_X1 U11427 ( .B1(n12034), .B2(n12130), .A(n12033), .ZN(n13825) );
  NAND2_X1 U11428 ( .A1(n11388), .A2(n11387), .ZN(n11414) );
  OR2_X1 U11429 ( .A1(n10795), .A2(n15387), .ZN(n15222) );
  OR2_X1 U11430 ( .A1(n12867), .A2(n13505), .ZN(n13506) );
  OR2_X1 U11431 ( .A1(n10796), .A2(n15357), .ZN(n15186) );
  NAND2_X1 U11432 ( .A1(n10802), .A2(n12555), .ZN(n10801) );
  OR2_X1 U11433 ( .A1(n10532), .A2(n10523), .ZN(n19442) );
  NAND2_X1 U11434 ( .A1(n11340), .A2(n9867), .ZN(n11388) );
  NAND2_X1 U11435 ( .A1(n12865), .A2(n12864), .ZN(n12867) );
  OR2_X1 U11436 ( .A1(n18808), .A2(n15176), .ZN(n10795) );
  AOI21_X1 U11437 ( .B1(n17888), .B2(n17649), .A(n17528), .ZN(n11888) );
  OR2_X1 U11438 ( .A1(n10532), .A2(n10524), .ZN(n10581) );
  NAND2_X1 U11439 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(n17746), .ZN(n17598) );
  NOR2_X1 U11440 ( .A1(n10520), .A2(n10524), .ZN(n19321) );
  AND2_X1 U11441 ( .A1(n15179), .A2(n10756), .ZN(n15238) );
  OR2_X1 U11442 ( .A1(n18820), .A2(n15176), .ZN(n10798) );
  XNOR2_X1 U11443 ( .A(n11267), .B(n20069), .ZN(n13733) );
  INV_X1 U11444 ( .A(n11342), .ZN(n11340) );
  OR2_X1 U11445 ( .A1(n10778), .A2(n10777), .ZN(n10786) );
  NAND2_X1 U11446 ( .A1(n11216), .A2(n11215), .ZN(n11267) );
  NAND2_X1 U11447 ( .A1(n17646), .A2(n10165), .ZN(n17587) );
  AND2_X1 U11448 ( .A1(n10755), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10790) );
  NAND2_X1 U11449 ( .A1(n10770), .A2(n10769), .ZN(n10778) );
  AOI21_X1 U11450 ( .B1(n13362), .B2(n13361), .A(n12884), .ZN(n13501) );
  BUF_X2 U11451 ( .A(n12868), .Z(n19105) );
  NAND2_X1 U11452 ( .A1(n12555), .A2(n10753), .ZN(n10770) );
  AND2_X1 U11453 ( .A1(n11886), .A2(n17988), .ZN(n17646) );
  XNOR2_X1 U11454 ( .A(n11213), .B(n20041), .ZN(n13626) );
  OR2_X1 U11455 ( .A1(n10759), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10753) );
  XNOR2_X1 U11456 ( .A(n15523), .B(n12882), .ZN(n13362) );
  NOR2_X2 U11457 ( .A1(n17337), .A2(n17253), .ZN(n17251) );
  AND2_X1 U11458 ( .A1(n10745), .A2(n10142), .ZN(n10773) );
  NAND2_X1 U11459 ( .A1(n10097), .A2(n10099), .ZN(n20041) );
  NAND2_X2 U11460 ( .A1(n14529), .A2(n13492), .ZN(n14566) );
  NAND2_X1 U11461 ( .A1(n17111), .A2(P3_EAX_REG_0__SCAN_IN), .ZN(n17253) );
  NOR2_X2 U11462 ( .A1(n19125), .A2(n19613), .ZN(n19126) );
  NAND2_X1 U11463 ( .A1(n12877), .A2(n12876), .ZN(n15523) );
  NOR2_X2 U11464 ( .A1(n19119), .A2(n19613), .ZN(n19120) );
  NOR2_X2 U11465 ( .A1(n19115), .A2(n19613), .ZN(n19116) );
  INV_X2 U11466 ( .A(n13416), .ZN(n20026) );
  NOR2_X2 U11467 ( .A1(n16313), .A2(n16345), .ZN(n18052) );
  NOR2_X1 U11468 ( .A1(n10484), .A2(n10496), .ZN(n10228) );
  OR2_X1 U11469 ( .A1(n11226), .A2(n11225), .ZN(n11227) );
  NAND2_X1 U11470 ( .A1(n9884), .A2(n12555), .ZN(n10745) );
  NAND2_X1 U11471 ( .A1(n9955), .A2(n11192), .ZN(n11208) );
  NAND2_X1 U11472 ( .A1(n9956), .A2(n9952), .ZN(n9951) );
  AND2_X1 U11473 ( .A1(n10907), .A2(n10489), .ZN(n10490) );
  OR2_X1 U11474 ( .A1(n10494), .A2(n10495), .ZN(n10504) );
  INV_X1 U11475 ( .A(n18554), .ZN(n18566) );
  NOR2_X1 U11476 ( .A1(n10033), .A2(n11239), .ZN(n10032) );
  NOR2_X1 U11477 ( .A1(n10140), .A2(n10139), .ZN(n10733) );
  NAND2_X1 U11478 ( .A1(n13249), .A2(n13248), .ZN(n18951) );
  NAND4_X1 U11479 ( .A1(n10466), .A2(n10465), .A3(n10482), .A4(n10464), .ZN(
        n10494) );
  NAND2_X1 U11480 ( .A1(n11276), .A2(n11275), .ZN(n20257) );
  OAI21_X1 U11481 ( .B1(n10482), .B2(n15554), .A(n10483), .ZN(n10496) );
  NOR2_X1 U11482 ( .A1(n10705), .A2(n10704), .ZN(n10718) );
  AND2_X1 U11483 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n11960), .ZN(
        n11961) );
  NOR2_X1 U11484 ( .A1(n10659), .A2(n10658), .ZN(n10688) );
  OR2_X1 U11485 ( .A1(n11926), .A2(n17312), .ZN(n10073) );
  NOR2_X1 U11486 ( .A1(n17233), .A2(n11855), .ZN(n11880) );
  AND2_X1 U11487 ( .A1(n10440), .A2(n10441), .ZN(n12657) );
  NAND3_X1 U11488 ( .A1(n12613), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n10426), 
        .ZN(n10267) );
  OAI21_X1 U11489 ( .B1(n10422), .B2(n12641), .A(n10421), .ZN(n12658) );
  OR2_X1 U11490 ( .A1(n17727), .A2(n17726), .ZN(n10159) );
  NAND2_X1 U11491 ( .A1(n18106), .A2(n11917), .ZN(n11912) );
  NOR2_X1 U11492 ( .A1(n17240), .A2(n11950), .ZN(n11874) );
  OR2_X1 U11493 ( .A1(n13454), .A2(n11488), .ZN(n11597) );
  AND2_X1 U11494 ( .A1(n14432), .A2(n11608), .ZN(n11096) );
  AND2_X1 U11495 ( .A1(n14427), .A2(n12493), .ZN(n13280) );
  NOR2_X1 U11496 ( .A1(n13221), .A2(n16144), .ZN(n13223) );
  INV_X1 U11497 ( .A(n10434), .ZN(n12592) );
  NAND2_X1 U11498 ( .A1(n17244), .A2(n17250), .ZN(n11950) );
  NAND2_X1 U11499 ( .A1(n13281), .A2(n11501), .ZN(n20793) );
  NAND2_X1 U11500 ( .A1(n11109), .A2(n11600), .ZN(n11487) );
  INV_X2 U11501 ( .A(n11501), .ZN(n12498) );
  INV_X1 U11502 ( .A(n15187), .ZN(n15176) );
  AND2_X1 U11503 ( .A1(n10238), .A2(n10428), .ZN(n10237) );
  OR2_X1 U11504 ( .A1(n11818), .A2(n11817), .ZN(n17244) );
  INV_X1 U11505 ( .A(n18123), .ZN(n17115) );
  INV_X2 U11506 ( .A(n10416), .ZN(n19114) );
  INV_X1 U11507 ( .A(n12645), .ZN(n13942) );
  NAND4_X1 U11508 ( .A1(n11830), .A2(n11834), .A3(n11833), .A4(n9880), .ZN(
        n17250) );
  OR2_X1 U11509 ( .A1(n10565), .A2(n10564), .ZN(n10855) );
  OR2_X1 U11510 ( .A1(n10578), .A2(n10577), .ZN(n10641) );
  NOR2_X1 U11511 ( .A1(n11108), .A2(n20129), .ZN(n13656) );
  INV_X2 U11512 ( .A(U212), .ZN(n16404) );
  NAND2_X1 U11513 ( .A1(n10413), .A2(n10412), .ZN(n12645) );
  OR2_X1 U11514 ( .A1(n10701), .A2(n10700), .ZN(n12702) );
  OR2_X1 U11515 ( .A1(n11161), .A2(n11160), .ZN(n11390) );
  AND4_X1 U11516 ( .A1(n10620), .A2(n10619), .A3(n10618), .A4(n10617), .ZN(
        n10636) );
  AND2_X1 U11517 ( .A1(n10005), .A2(n10004), .ZN(n10447) );
  NAND2_X1 U11518 ( .A1(n9853), .A2(n9885), .ZN(n11121) );
  OR2_X1 U11519 ( .A1(n10715), .A2(n10714), .ZN(n12706) );
  INV_X1 U11520 ( .A(n11127), .ZN(n11176) );
  AND4_X1 U11521 ( .A1(n11061), .A2(n11060), .A3(n11059), .A4(n11058), .ZN(
        n11077) );
  AND4_X1 U11522 ( .A1(n11065), .A2(n11064), .A3(n11063), .A4(n11062), .ZN(
        n11076) );
  AND4_X1 U11523 ( .A1(n10998), .A2(n10997), .A3(n10996), .A4(n10995), .ZN(
        n11013) );
  AND4_X1 U11524 ( .A1(n10994), .A2(n10993), .A3(n10992), .A4(n10991), .ZN(
        n11014) );
  AND4_X1 U11525 ( .A1(n11030), .A2(n11029), .A3(n11028), .A4(n11027), .ZN(
        n11031) );
  NAND2_X2 U11526 ( .A1(n19853), .A2(n19735), .ZN(n19775) );
  NAND2_X2 U11527 ( .A1(P2_STATE_REG_2__SCAN_IN), .A2(n19853), .ZN(n19772) );
  AND4_X1 U11528 ( .A1(n11073), .A2(n11072), .A3(n11071), .A4(n11070), .ZN(
        n11074) );
  AND4_X1 U11529 ( .A1(n11038), .A2(n11037), .A3(n11036), .A4(n11035), .ZN(
        n11057) );
  AND4_X1 U11530 ( .A1(n11046), .A2(n11045), .A3(n11044), .A4(n11043), .ZN(
        n11053) );
  AND4_X1 U11531 ( .A1(n11018), .A2(n11017), .A3(n11016), .A4(n11015), .ZN(
        n11034) );
  AND4_X1 U11532 ( .A1(n11022), .A2(n11021), .A3(n11020), .A4(n11019), .ZN(
        n11033) );
  AND4_X1 U11533 ( .A1(n11026), .A2(n11025), .A3(n11024), .A4(n11023), .ZN(
        n11032) );
  AND4_X1 U11534 ( .A1(n10405), .A2(n10404), .A3(n10403), .A4(n10402), .ZN(
        n10406) );
  AND4_X1 U11535 ( .A1(n11106), .A2(n11105), .A3(n11104), .A4(n11103), .ZN(
        n11107) );
  INV_X1 U11536 ( .A(n11821), .ZN(n17006) );
  INV_X2 U11537 ( .A(n11792), .ZN(n9830) );
  CLKBUF_X3 U11538 ( .A(n17063), .Z(n17019) );
  BUF_X2 U11539 ( .A(n11691), .Z(n17024) );
  AND3_X1 U11540 ( .A1(n10363), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A3(
        n10362), .ZN(n10366) );
  AND2_X2 U11541 ( .A1(n9837), .A2(n16232), .ZN(n10671) );
  INV_X2 U11542 ( .A(n15622), .ZN(n15609) );
  BUF_X2 U11543 ( .A(n11858), .Z(n9842) );
  AND2_X1 U11544 ( .A1(n10392), .A2(n16232), .ZN(n10396) );
  INV_X2 U11545 ( .A(n16438), .ZN(U215) );
  INV_X2 U11546 ( .A(n19854), .ZN(n19853) );
  INV_X2 U11547 ( .A(n16441), .ZN(n16443) );
  NAND2_X2 U11548 ( .A1(n18682), .A2(n18625), .ZN(n18685) );
  AND2_X2 U11549 ( .A1(n11004), .A2(n11006), .ZN(n11193) );
  OR2_X2 U11550 ( .A1(n11647), .A2(n11639), .ZN(n15622) );
  NOR2_X1 U11551 ( .A1(n18563), .A2(n11648), .ZN(n11677) );
  BUF_X4 U11552 ( .A(n10539), .Z(n9837) );
  NOR2_X2 U11553 ( .A1(n11646), .A2(n18563), .ZN(n17063) );
  NOR2_X1 U11554 ( .A1(n16793), .A2(n11639), .ZN(n11691) );
  NOR2_X2 U11555 ( .A1(n18563), .A2(n11649), .ZN(n11827) );
  AND2_X2 U11556 ( .A1(n13594), .A2(n15554), .ZN(n13172) );
  AND2_X2 U11557 ( .A1(n10546), .A2(n10315), .ZN(n10541) );
  AND2_X2 U11558 ( .A1(n13687), .A2(n13672), .ZN(n11246) );
  AND2_X2 U11559 ( .A1(n11235), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11005) );
  NAND3_X2 U11560 ( .A1(n18604), .A2(n18603), .A3(n18723), .ZN(n18074) );
  NAND2_X1 U11561 ( .A1(n11640), .A2(n18713), .ZN(n11648) );
  INV_X2 U11562 ( .A(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11235) );
  AND2_X1 U11563 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18542) );
  NAND2_X1 U11564 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n11639) );
  NAND2_X2 U11565 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n18563) );
  NOR2_X2 U11566 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15532) );
  INV_X1 U11567 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9959) );
  AND2_X2 U11568 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10546) );
  AND2_X2 U11569 ( .A1(n10003), .A2(n10002), .ZN(n10416) );
  AND2_X4 U11570 ( .A1(n10999), .A2(n13672), .ZN(n11047) );
  NOR2_X1 U11571 ( .A1(n18563), .A2(n11649), .ZN(n9823) );
  NAND2_X2 U11572 ( .A1(n10239), .A2(n10237), .ZN(n12635) );
  NOR2_X1 U11573 ( .A1(n10267), .A2(n12635), .ZN(n9824) );
  NOR2_X2 U11574 ( .A1(n10267), .A2(n12635), .ZN(n10468) );
  AND2_X2 U11575 ( .A1(n10546), .A2(n10315), .ZN(n9826) );
  NAND2_X1 U11576 ( .A1(n11596), .A2(n20122), .ZN(n13466) );
  AND2_X2 U11577 ( .A1(n13594), .A2(n15554), .ZN(n9827) );
  AND2_X2 U11578 ( .A1(n14284), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11006) );
  XNOR2_X1 U11579 ( .A(n11218), .B(n11217), .ZN(n11996) );
  OAI21_X2 U11580 ( .B1(n11987), .B2(n12168), .A(n11986), .ZN(n11988) );
  AND2_X1 U11581 ( .A1(n11120), .A2(n11121), .ZN(n14171) );
  INV_X1 U11582 ( .A(n11792), .ZN(n9829) );
  OR2_X1 U11583 ( .A1(n11645), .A2(n11648), .ZN(n11792) );
  AND2_X2 U11584 ( .A1(n11005), .A2(n10999), .ZN(n12465) );
  INV_X1 U11585 ( .A(n11826), .ZN(n9844) );
  NAND2_X2 U11586 ( .A1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n11640), .ZN(
        n11646) );
  OR2_X1 U11587 ( .A1(n11144), .A2(n11143), .ZN(n11145) );
  NAND2_X1 U11588 ( .A1(n11144), .A2(n11143), .ZN(n9957) );
  INV_X1 U11589 ( .A(n15622), .ZN(n9832) );
  OAI21_X1 U11590 ( .B1(n11234), .B2(n11235), .A(n11238), .ZN(n11239) );
  OAI21_X2 U11591 ( .B1(n11234), .B2(n13661), .A(n11185), .ZN(n11189) );
  AND2_X4 U11592 ( .A1(n15532), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n9833) );
  AND3_X4 U11593 ( .A1(n10315), .A2(n15554), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n9834) );
  AND2_X2 U11594 ( .A1(n14372), .A2(n14547), .ZN(n14486) );
  NOR2_X2 U11595 ( .A1(n14147), .A2(n10211), .ZN(n14372) );
  NAND2_X1 U11596 ( .A1(n10874), .A2(n13925), .ZN(n13917) );
  OAI21_X1 U11597 ( .B1(n11987), .B2(n11423), .A(n11266), .ZN(n13732) );
  AND2_X1 U11598 ( .A1(n11176), .A2(n11180), .ZN(n13267) );
  NOR2_X2 U11599 ( .A1(n14100), .A2(n14102), .ZN(n14101) );
  XNOR2_X1 U11600 ( .A(n10869), .B(n10868), .ZN(n10874) );
  NAND2_X2 U11601 ( .A1(n11470), .A2(n13281), .ZN(n13453) );
  AND3_X2 U11602 ( .A1(n11125), .A2(n11124), .A3(n9902), .ZN(n11470) );
  AND2_X1 U11603 ( .A1(n11004), .A2(n13673), .ZN(n9835) );
  AND2_X1 U11604 ( .A1(n11004), .A2(n13673), .ZN(n9836) );
  INV_X2 U11605 ( .A(n16797), .ZN(n16770) );
  XNOR2_X1 U11607 ( .A(n14322), .B(n12486), .ZN(n14504) );
  AND2_X2 U11608 ( .A1(n10227), .A2(n9875), .ZN(n15160) );
  NOR2_X2 U11609 ( .A1(n10415), .A2(n12588), .ZN(n15659) );
  NOR2_X1 U11610 ( .A1(n11646), .A2(n11645), .ZN(n11805) );
  NAND2_X2 U11611 ( .A1(n14321), .A2(n14301), .ZN(n14305) );
  NAND2_X1 U11612 ( .A1(n12668), .A2(n19114), .ZN(n12571) );
  INV_X2 U11614 ( .A(n9839), .ZN(n12613) );
  AND2_X1 U11615 ( .A1(n10546), .A2(n10547), .ZN(n12975) );
  NOR2_X1 U11616 ( .A1(n11646), .A2(n11647), .ZN(n15560) );
  NAND2_X2 U11617 ( .A1(n14139), .A2(n12171), .ZN(n14147) );
  NAND2_X2 U11618 ( .A1(n14122), .A2(n12106), .ZN(n14139) );
  AND2_X4 U11619 ( .A1(n10092), .A2(n10091), .ZN(n18929) );
  NOR2_X1 U11620 ( .A1(n11640), .A2(n10084), .ZN(n11858) );
  AND2_X1 U11621 ( .A1(n10999), .A2(n13667), .ZN(n9843) );
  AND2_X4 U11622 ( .A1(n11006), .A2(n13667), .ZN(n11110) );
  NAND2_X4 U11623 ( .A1(n10906), .A2(n10285), .ZN(n10521) );
  NAND2_X2 U11624 ( .A1(n9992), .A2(n10490), .ZN(n10906) );
  NAND2_X2 U11625 ( .A1(n13453), .A2(n13466), .ZN(n10201) );
  INV_X1 U11626 ( .A(n9844), .ZN(n9845) );
  INV_X1 U11627 ( .A(n9844), .ZN(n9846) );
  NOR2_X1 U11628 ( .A1(n11649), .A2(n11647), .ZN(n11826) );
  NOR2_X1 U11629 ( .A1(n11961), .A2(n17690), .ZN(n17678) );
  NOR2_X4 U11630 ( .A1(n15440), .A2(n16196), .ZN(n15247) );
  NAND2_X2 U11631 ( .A1(n16146), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15440) );
  OAI211_X2 U11632 ( .C1(n9956), .C2(n9954), .A(n9953), .B(n9951), .ZN(n11989)
         );
  NAND2_X2 U11633 ( .A1(n11218), .A2(n11217), .ZN(n9956) );
  NOR2_X2 U11634 ( .A1(n10507), .A2(n19105), .ZN(n19159) );
  INV_X1 U11635 ( .A(n9899), .ZN(n10913) );
  AOI211_X1 U11636 ( .C1(n20766), .C2(n20765), .A(n20764), .B(n20763), .ZN(
        n20769) );
  XNOR2_X2 U11637 ( .A(n10220), .B(n10030), .ZN(n20766) );
  OAI22_X2 U11638 ( .A1(n10499), .A2(n10228), .B1(n10497), .B2(n10229), .ZN(
        n10492) );
  INV_X2 U11639 ( .A(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n10315) );
  NOR2_X4 U11640 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15542) );
  AND2_X2 U11641 ( .A1(n10538), .A2(n16232), .ZN(n10676) );
  AND2_X4 U11642 ( .A1(n15542), .A2(n10315), .ZN(n10538) );
  NAND2_X1 U11643 ( .A1(n14588), .A2(n14688), .ZN(n10296) );
  NAND2_X1 U11644 ( .A1(n10040), .A2(n9958), .ZN(n10026) );
  AND2_X1 U11645 ( .A1(n10027), .A2(n11407), .ZN(n9958) );
  NOR2_X1 U11646 ( .A1(n10096), .A2(n10028), .ZN(n10027) );
  NOR2_X1 U11647 ( .A1(n14688), .A2(n11550), .ZN(n10028) );
  AOI21_X1 U11648 ( .B1(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n19796), .A(
        n10670), .ZN(n10835) );
  NOR2_X1 U11649 ( .A1(n16052), .A2(n15176), .ZN(n15097) );
  INV_X1 U11650 ( .A(n16292), .ZN(n13386) );
  INV_X1 U11651 ( .A(n10059), .ZN(n10058) );
  OAI21_X1 U11652 ( .B1(n10061), .B2(n10060), .A(n15453), .ZN(n10059) );
  INV_X1 U11653 ( .A(n11341), .ZN(n11339) );
  NAND2_X1 U11654 ( .A1(n11997), .A2(n11180), .ZN(n11126) );
  OR2_X1 U11655 ( .A1(n11127), .A2(n11192), .ZN(n11278) );
  OR2_X1 U11656 ( .A1(n11501), .A2(n11192), .ZN(n11277) );
  NAND2_X1 U11657 ( .A1(n12493), .A2(n11588), .ZN(n11586) );
  INV_X1 U11658 ( .A(n11586), .ZN(n11581) );
  NAND3_X1 U11659 ( .A1(n11127), .A2(n11501), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11438) );
  NAND2_X1 U11660 ( .A1(n10815), .A2(n14974), .ZN(n10816) );
  NOR2_X1 U11661 ( .A1(n16039), .A2(n15176), .ZN(n15098) );
  INV_X1 U11662 ( .A(n14870), .ZN(n10954) );
  OAI21_X1 U11663 ( .B1(n15188), .B2(n9882), .A(n15187), .ZN(n10281) );
  NAND2_X1 U11664 ( .A1(n10420), .A2(n12641), .ZN(n10421) );
  NAND2_X1 U11665 ( .A1(n12664), .A2(n16281), .ZN(n12819) );
  AND2_X1 U11666 ( .A1(n9983), .A2(n19798), .ZN(n12664) );
  AND2_X1 U11667 ( .A1(n10471), .A2(n10446), .ZN(n13181) );
  NAND2_X1 U11668 ( .A1(n20789), .A2(n12489), .ZN(n14430) );
  OR2_X1 U11669 ( .A1(n14688), .A2(n14710), .ZN(n11413) );
  NAND2_X1 U11670 ( .A1(n10095), .A2(n14688), .ZN(n15860) );
  NOR2_X1 U11671 ( .A1(n10207), .A2(n9936), .ZN(n10206) );
  INV_X1 U11672 ( .A(n10026), .ZN(n10025) );
  AND2_X1 U11673 ( .A1(n11493), .A2(n11492), .ZN(n11620) );
  INV_X1 U11674 ( .A(n13829), .ZN(n10186) );
  NAND2_X1 U11675 ( .A1(n15096), .A2(n15097), .ZN(n9977) );
  AND2_X1 U11676 ( .A1(n10885), .A2(n10886), .ZN(n16172) );
  NOR2_X1 U11677 ( .A1(n15481), .A2(n10277), .ZN(n10276) );
  INV_X1 U11678 ( .A(n10278), .ZN(n10277) );
  OR2_X1 U11679 ( .A1(n14080), .A2(n10725), .ZN(n10279) );
  NAND2_X1 U11680 ( .A1(n15520), .A2(n10070), .ZN(n13591) );
  INV_X1 U11681 ( .A(n12657), .ZN(n10070) );
  NAND2_X1 U11682 ( .A1(n12612), .A2(n13386), .ZN(n12663) );
  AND2_X1 U11683 ( .A1(n10983), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n12881) );
  NAND2_X1 U11684 ( .A1(n12584), .A2(n12583), .ZN(n16257) );
  NAND2_X1 U11685 ( .A1(n11682), .A2(n9887), .ZN(n10078) );
  AND2_X1 U11686 ( .A1(n19113), .A2(n19807), .ZN(n19104) );
  NOR2_X1 U11687 ( .A1(n10983), .A2(n15530), .ZN(n9960) );
  AOI22_X1 U11688 ( .A1(n10538), .A2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n9827), .B2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n10405) );
  INV_X1 U11689 ( .A(n11366), .ZN(n10210) );
  NAND2_X1 U11690 ( .A1(n20771), .A2(n11192), .ZN(n11291) );
  AND2_X1 U11691 ( .A1(n10648), .A2(n10649), .ZN(n10670) );
  NOR2_X1 U11692 ( .A1(n10368), .A2(n10302), .ZN(n10372) );
  AOI21_X1 U11693 ( .B1(n9826), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10367) );
  NAND2_X1 U11694 ( .A1(n10424), .A2(n10472), .ZN(n9961) );
  NOR2_X1 U11695 ( .A1(n10453), .A2(n10291), .ZN(n10424) );
  OR2_X1 U11696 ( .A1(n18872), .A2(n15176), .ZN(n10768) );
  AND2_X1 U11697 ( .A1(n10587), .A2(n10586), .ZN(n10588) );
  NAND2_X1 U11698 ( .A1(n10467), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10482) );
  AND2_X1 U11699 ( .A1(n12613), .A2(n10426), .ZN(n10471) );
  AOI22_X1 U11700 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9825), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n10322) );
  INV_X1 U11701 ( .A(n14360), .ZN(n10218) );
  AND2_X1 U11702 ( .A1(n14454), .A2(n14462), .ZN(n10219) );
  NAND2_X1 U11703 ( .A1(n10213), .A2(n10212), .ZN(n10211) );
  INV_X1 U11704 ( .A(n10214), .ZN(n10213) );
  INV_X1 U11705 ( .A(n14374), .ZN(n10212) );
  OR2_X1 U11706 ( .A1(n10215), .A2(n14388), .ZN(n10214) );
  INV_X1 U11707 ( .A(n12481), .ZN(n12447) );
  NAND2_X1 U11708 ( .A1(n12172), .A2(P1_STATE2_REG_0__SCAN_IN), .ZN(n12481) );
  NAND2_X1 U11709 ( .A1(n10098), .A2(n11212), .ZN(n11213) );
  NAND2_X1 U11710 ( .A1(n11208), .A2(n10101), .ZN(n10098) );
  INV_X1 U11711 ( .A(n11120), .ZN(n11997) );
  NOR2_X1 U11712 ( .A1(n20145), .A2(n20691), .ZN(n11999) );
  AND2_X1 U11713 ( .A1(n11397), .A2(n14636), .ZN(n10174) );
  AND2_X1 U11714 ( .A1(n14151), .A2(n14180), .ZN(n10134) );
  INV_X1 U11715 ( .A(n11385), .ZN(n10018) );
  NAND2_X1 U11716 ( .A1(n10017), .A2(n11385), .ZN(n10016) );
  INV_X1 U11717 ( .A(n11384), .ZN(n10017) );
  NAND2_X1 U11718 ( .A1(n11395), .A2(n11394), .ZN(n10039) );
  INV_X1 U11719 ( .A(n11576), .ZN(n11591) );
  AND2_X1 U11720 ( .A1(n11500), .A2(n11588), .ZN(n11576) );
  NAND2_X1 U11721 ( .A1(n9948), .A2(n12498), .ZN(n11610) );
  XNOR2_X1 U11722 ( .A(n11255), .B(n11254), .ZN(n11257) );
  NAND2_X1 U11723 ( .A1(n11127), .A2(n11121), .ZN(n11123) );
  INV_X1 U11724 ( .A(n15059), .ZN(n10199) );
  AND2_X1 U11725 ( .A1(n15330), .A2(n15066), .ZN(n10200) );
  NOR2_X1 U11726 ( .A1(n15163), .A2(n10086), .ZN(n10085) );
  INV_X1 U11727 ( .A(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n10086) );
  NOR2_X1 U11728 ( .A1(n16157), .A2(n10088), .ZN(n10087) );
  INV_X1 U11729 ( .A(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n10088) );
  AND2_X1 U11730 ( .A1(n15025), .A2(n14234), .ZN(n14261) );
  INV_X1 U11731 ( .A(n15000), .ZN(n10258) );
  NAND2_X1 U11732 ( .A1(n10280), .A2(n9894), .ZN(n9985) );
  NAND2_X1 U11733 ( .A1(n13789), .A2(n13802), .ZN(n10193) );
  NOR2_X1 U11734 ( .A1(n10062), .A2(n15467), .ZN(n10061) );
  INV_X1 U11735 ( .A(n10272), .ZN(n10062) );
  NAND2_X1 U11736 ( .A1(n10278), .A2(n10725), .ZN(n10274) );
  AND4_X1 U11737 ( .A1(n10628), .A2(n10627), .A3(n10626), .A4(n10625), .ZN(
        n10634) );
  AND4_X1 U11738 ( .A1(n10632), .A2(n10631), .A3(n10630), .A4(n10629), .ZN(
        n10633) );
  AND4_X1 U11739 ( .A1(n10624), .A2(n10623), .A3(n10622), .A4(n10621), .ZN(
        n10635) );
  AOI21_X1 U11740 ( .B1(n12708), .B2(n9906), .A(n10197), .ZN(n10196) );
  INV_X1 U11741 ( .A(n13499), .ZN(n10197) );
  CLKBUF_X1 U11742 ( .A(n12598), .Z(n12599) );
  AOI21_X1 U11743 ( .B1(n13717), .B2(n12680), .A(n12679), .ZN(n12687) );
  INV_X1 U11744 ( .A(n12580), .ZN(n12584) );
  NOR2_X1 U11745 ( .A1(n12868), .A2(n15507), .ZN(n10522) );
  NAND2_X1 U11746 ( .A1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n18727), .ZN(
        n11645) );
  NAND2_X2 U11747 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18720), .ZN(
        n11647) );
  NOR2_X1 U11748 ( .A1(n16793), .A2(n11648), .ZN(n11821) );
  NAND2_X1 U11749 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n10080) );
  NOR2_X1 U11750 ( .A1(n15726), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16298) );
  NOR2_X1 U11751 ( .A1(n17668), .A2(n11885), .ZN(n11886) );
  AND2_X1 U11752 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n11875), .ZN(
        n11876) );
  INV_X1 U11753 ( .A(n11873), .ZN(n10153) );
  AOI211_X1 U11754 ( .C1(n18112), .C2(n11737), .A(n11736), .B(n11735), .ZN(
        n11924) );
  OAI21_X1 U11755 ( .B1(n18112), .B2(n11738), .A(n11924), .ZN(n11914) );
  AND3_X1 U11756 ( .A1(n11923), .A2(n11902), .A3(n18106), .ZN(n11738) );
  NOR3_X1 U11757 ( .A1(n18123), .A2(n11912), .A3(n11911), .ZN(n14225) );
  NOR2_X1 U11758 ( .A1(n9852), .A2(n10122), .ZN(n10121) );
  INV_X1 U11759 ( .A(n14056), .ZN(n10122) );
  AND2_X1 U11760 ( .A1(n12493), .A2(n11514), .ZN(n13522) );
  AND2_X1 U11761 ( .A1(n20691), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12485) );
  AND2_X1 U11762 ( .A1(n12457), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12490) );
  NOR2_X2 U11763 ( .A1(n14321), .A2(n14323), .ZN(n14322) );
  NOR2_X2 U11764 ( .A1(n14337), .A2(n14339), .ZN(n14338) );
  INV_X1 U11765 ( .A(n12057), .ZN(n12061) );
  INV_X1 U11766 ( .A(n13825), .ZN(n12035) );
  NAND2_X1 U11767 ( .A1(n12020), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12025) );
  INV_X1 U11768 ( .A(n13522), .ZN(n12495) );
  OR2_X1 U11769 ( .A1(n12523), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9944) );
  INV_X1 U11770 ( .A(n9938), .ZN(n9937) );
  OAI21_X1 U11771 ( .B1(n11415), .B2(n9939), .A(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n9938) );
  NAND2_X1 U11772 ( .A1(n9947), .A2(n11415), .ZN(n12522) );
  NOR3_X1 U11773 ( .A1(n14468), .A2(n10131), .A3(n10128), .ZN(n14336) );
  OR2_X1 U11774 ( .A1(n10129), .A2(n14334), .ZN(n10128) );
  INV_X1 U11775 ( .A(n14589), .ZN(n10022) );
  NOR2_X1 U11776 ( .A1(n14498), .A2(n14497), .ZN(n14499) );
  AND2_X1 U11777 ( .A1(n11397), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n10209) );
  INV_X1 U11778 ( .A(n20062), .ZN(n14786) );
  NOR2_X1 U11779 ( .A1(n14841), .A2(n14185), .ZN(n14186) );
  AND2_X1 U11780 ( .A1(n11535), .A2(n11534), .ZN(n14838) );
  NAND2_X1 U11781 ( .A1(n10014), .A2(n11385), .ZN(n13954) );
  NAND2_X1 U11782 ( .A1(n15898), .A2(n11384), .ZN(n10014) );
  NOR2_X1 U11783 ( .A1(n11611), .A2(n11603), .ZN(n13658) );
  AND2_X1 U11784 ( .A1(n9950), .A2(n20122), .ZN(n10169) );
  NAND2_X1 U11785 ( .A1(n10112), .A2(n9910), .ZN(n10111) );
  NOR2_X1 U11786 ( .A1(n10115), .A2(n10116), .ZN(n10112) );
  NAND2_X1 U11787 ( .A1(n13522), .A2(n20087), .ZN(n10114) );
  AOI21_X1 U11788 ( .B1(n11423), .B2(n11183), .A(n10100), .ZN(n10099) );
  INV_X1 U11789 ( .A(n20413), .ZN(n20549) );
  INV_X1 U11790 ( .A(n20434), .ZN(n20579) );
  NOR2_X1 U11791 ( .A1(n20378), .A2(n10030), .ZN(n20580) );
  OR2_X1 U11792 ( .A1(n11469), .A2(n11468), .ZN(n13698) );
  AND2_X1 U11793 ( .A1(n11479), .A2(n11467), .ZN(n11468) );
  AOI21_X1 U11794 ( .B1(n11466), .B2(n11479), .A(n11465), .ZN(n11469) );
  NOR2_X1 U11795 ( .A1(n9877), .A2(n15024), .ZN(n15025) );
  OAI21_X1 U11796 ( .B1(n10820), .B2(n10751), .A(n10821), .ZN(n10824) );
  INV_X1 U11797 ( .A(n14997), .ZN(n10250) );
  NAND2_X1 U11798 ( .A1(n10942), .A2(n9917), .ZN(n14870) );
  INV_X1 U11799 ( .A(n14955), .ZN(n10243) );
  XNOR2_X1 U11800 ( .A(n13081), .B(n10308), .ZN(n14964) );
  NOR2_X1 U11801 ( .A1(n15485), .A2(n15484), .ZN(n13739) );
  INV_X1 U11802 ( .A(n10433), .ZN(n10239) );
  XNOR2_X1 U11803 ( .A(n10094), .B(n10093), .ZN(n14289) );
  INV_X1 U11804 ( .A(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n10093) );
  NAND2_X1 U11805 ( .A1(n13228), .A2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n10094) );
  NOR2_X2 U11806 ( .A1(n15686), .A2(n15152), .ZN(n15151) );
  NAND2_X1 U11807 ( .A1(n13211), .A2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14867) );
  NOR2_X1 U11808 ( .A1(n14078), .A2(n10882), .ZN(n10001) );
  NAND2_X1 U11809 ( .A1(n14078), .A2(n10882), .ZN(n9966) );
  INV_X1 U11810 ( .A(n14077), .ZN(n9999) );
  NAND2_X1 U11811 ( .A1(n14077), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n10000) );
  INV_X1 U11812 ( .A(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n14901) );
  NAND2_X1 U11813 ( .A1(n10235), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10230) );
  NOR2_X1 U11814 ( .A1(n15098), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10271) );
  OR2_X1 U11815 ( .A1(n15097), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10299) );
  NOR2_X1 U11816 ( .A1(n9889), .A2(n15093), .ZN(n10270) );
  NAND2_X1 U11817 ( .A1(n21005), .A2(n15263), .ZN(n10145) );
  NAND2_X1 U11818 ( .A1(n15105), .A2(n10010), .ZN(n15265) );
  OR2_X1 U11819 ( .A1(n15112), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10010) );
  AOI21_X1 U11820 ( .B1(n15325), .B2(n15326), .A(n15328), .ZN(n15157) );
  NAND2_X1 U11821 ( .A1(n15182), .A2(n15181), .ZN(n15219) );
  INV_X1 U11822 ( .A(n10050), .ZN(n10049) );
  AOI21_X1 U11823 ( .B1(n10050), .B2(n10052), .A(n10048), .ZN(n10047) );
  AOI21_X1 U11824 ( .B1(n15249), .B2(n10053), .A(n10051), .ZN(n10050) );
  INV_X1 U11825 ( .A(n15179), .ZN(n10051) );
  INV_X1 U11826 ( .A(n15251), .ZN(n10056) );
  AND2_X1 U11827 ( .A1(n10728), .A2(n14214), .ZN(n10278) );
  NAND2_X1 U11828 ( .A1(n10194), .A2(n10196), .ZN(n14048) );
  AOI21_X1 U11829 ( .B1(n9854), .B2(n9982), .A(n9920), .ZN(n9979) );
  NAND2_X1 U11830 ( .A1(n13865), .A2(n13924), .ZN(n9998) );
  XNOR2_X1 U11831 ( .A(n10702), .B(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n13922) );
  OR2_X1 U11832 ( .A1(n12694), .A2(n12693), .ZN(n13829) );
  INV_X1 U11833 ( .A(n19808), .ZN(n19786) );
  AOI21_X1 U11834 ( .B1(n15536), .B2(n12881), .A(n12880), .ZN(n13361) );
  NAND2_X1 U11835 ( .A1(n19788), .A2(n19158), .ZN(n19347) );
  NAND4_X1 U11836 ( .A1(n10396), .A2(n10395), .A3(n10394), .A4(n10393), .ZN(
        n10397) );
  NAND2_X1 U11837 ( .A1(n19407), .A2(n19158), .ZN(n19556) );
  INV_X1 U11838 ( .A(n19648), .ZN(n19613) );
  OAI22_X2 U11839 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n16286), .B1(n13938), 
        .B2(n19841), .ZN(n19648) );
  AOI21_X1 U11840 ( .B1(n9878), .B2(n18528), .A(n17313), .ZN(n11753) );
  NAND2_X1 U11841 ( .A1(n18542), .A2(n18727), .ZN(n10084) );
  OAI21_X1 U11842 ( .B1(n18558), .B2(n10083), .A(n14224), .ZN(n15744) );
  AND2_X1 U11843 ( .A1(n17312), .A2(n16313), .ZN(n10083) );
  NOR4_X2 U11844 ( .A1(n18094), .A2(n11912), .A3(n17115), .A4(n11730), .ZN(
        n17312) );
  NOR2_X1 U11845 ( .A1(n17438), .A2(n17410), .ZN(n11633) );
  AND2_X1 U11846 ( .A1(n9855), .A2(n9923), .ZN(n10180) );
  NAND2_X1 U11847 ( .A1(n17559), .A2(n17558), .ZN(n17581) );
  INV_X1 U11848 ( .A(n17694), .ZN(n10177) );
  AND2_X1 U11849 ( .A1(n11892), .A2(n10167), .ZN(n10166) );
  OAI21_X1 U11850 ( .B1(n17689), .B2(n10161), .A(n10160), .ZN(n17673) );
  NAND2_X1 U11851 ( .A1(n10164), .A2(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10161) );
  NAND2_X1 U11852 ( .A1(n11879), .A2(n10164), .ZN(n10160) );
  INV_X1 U11853 ( .A(n17674), .ZN(n10164) );
  OR2_X1 U11854 ( .A1(n17689), .A2(n18026), .ZN(n10163) );
  NAND2_X1 U11855 ( .A1(n11741), .A2(n9878), .ZN(n18555) );
  INV_X1 U11856 ( .A(n18595), .ZN(n18741) );
  AND2_X1 U11857 ( .A1(n14430), .A2(n12492), .ZN(n19908) );
  NAND2_X1 U11858 ( .A1(n12512), .A2(n12511), .ZN(n19934) );
  XNOR2_X1 U11859 ( .A(n10106), .B(n10105), .ZN(n14320) );
  INV_X1 U11860 ( .A(n12494), .ZN(n10105) );
  NAND2_X1 U11861 ( .A1(n10108), .A2(n10107), .ZN(n10106) );
  NAND2_X1 U11862 ( .A1(n11592), .A2(n12493), .ZN(n10107) );
  AND2_X2 U11863 ( .A1(n13182), .A2(n13386), .ZN(n14993) );
  NAND2_X1 U11864 ( .A1(n14993), .A2(n10443), .ZN(n15009) );
  INV_X1 U11865 ( .A(n13452), .ZN(n19081) );
  INV_X1 U11866 ( .A(n15109), .ZN(n9971) );
  NAND2_X1 U11867 ( .A1(n9977), .A2(n9974), .ZN(n9973) );
  NAND2_X1 U11868 ( .A1(n15099), .A2(n21005), .ZN(n9974) );
  NAND2_X1 U11869 ( .A1(n15109), .A2(n9972), .ZN(n9968) );
  AND2_X1 U11870 ( .A1(n9976), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n9972) );
  NAND2_X1 U11871 ( .A1(n13260), .A2(n10979), .ZN(n19113) );
  INV_X1 U11872 ( .A(n19101), .ZN(n19098) );
  NAND2_X1 U11873 ( .A1(n14274), .A2(n14273), .ZN(n14275) );
  NOR2_X1 U11874 ( .A1(n14272), .A2(n14271), .ZN(n14273) );
  NAND2_X1 U11875 ( .A1(n16017), .A2(n16209), .ZN(n14274) );
  XNOR2_X1 U11876 ( .A(n12620), .B(n12621), .ZN(n16018) );
  INV_X1 U11877 ( .A(n15100), .ZN(n16041) );
  INV_X1 U11878 ( .A(n16197), .ZN(n15444) );
  OR2_X1 U11879 ( .A1(n12663), .A2(n12631), .ZN(n16212) );
  NAND2_X1 U11880 ( .A1(n9967), .A2(n10616), .ZN(n9997) );
  INV_X1 U11881 ( .A(n16212), .ZN(n16219) );
  NAND2_X1 U11882 ( .A1(n18950), .A2(n12881), .ZN(n12877) );
  NAND2_X1 U11883 ( .A1(n18741), .A2(n18586), .ZN(n16450) );
  NAND2_X1 U11884 ( .A1(n10184), .A2(n10183), .ZN(n16569) );
  NAND2_X1 U11885 ( .A1(n16797), .A2(n17449), .ZN(n10183) );
  NOR2_X2 U11886 ( .A1(n18588), .A2(n11760), .ZN(n16782) );
  INV_X1 U11887 ( .A(n16811), .ZN(n16779) );
  NAND2_X1 U11888 ( .A1(n17118), .A2(n10077), .ZN(n10076) );
  OR2_X1 U11889 ( .A1(n17155), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n10077) );
  OR2_X1 U11890 ( .A1(n17120), .A2(n17252), .ZN(n17118) );
  NOR2_X1 U11891 ( .A1(n17332), .A2(n17124), .ZN(n17120) );
  NAND2_X1 U11892 ( .A1(P3_EAX_REG_28__SCAN_IN), .A2(n17132), .ZN(n17124) );
  AND2_X1 U11893 ( .A1(n17144), .A2(P3_EAX_REG_24__SCAN_IN), .ZN(n17140) );
  NOR2_X1 U11894 ( .A1(n17153), .A2(n17149), .ZN(n17144) );
  NAND2_X1 U11895 ( .A1(n17150), .A2(P3_EAX_REG_23__SCAN_IN), .ZN(n17149) );
  NAND2_X1 U11896 ( .A1(n17111), .A2(n17153), .ZN(n17247) );
  NOR2_X2 U11897 ( .A1(n16313), .A2(n16450), .ZN(n17742) );
  NAND2_X1 U11898 ( .A1(n10442), .A2(n13942), .ZN(n12597) );
  NAND2_X1 U11899 ( .A1(n13942), .A2(n10443), .ZN(n10434) );
  AND2_X1 U11900 ( .A1(n11420), .A2(n11419), .ZN(n11444) );
  AND2_X1 U11901 ( .A1(n11338), .A2(n11337), .ZN(n11341) );
  AND2_X1 U11902 ( .A1(n11207), .A2(n20122), .ZN(n10101) );
  INV_X1 U11903 ( .A(n14653), .ZN(n10096) );
  OR2_X1 U11904 ( .A1(n11362), .A2(n11361), .ZN(n11379) );
  OR2_X1 U11905 ( .A1(n11289), .A2(n11288), .ZN(n11313) );
  OR2_X1 U11906 ( .A1(n13486), .A2(n11127), .ZN(n11129) );
  NAND2_X1 U11907 ( .A1(n11596), .A2(n11482), .ZN(n11186) );
  NAND2_X1 U11908 ( .A1(n11129), .A2(n11135), .ZN(n10172) );
  AND2_X2 U11909 ( .A1(n10990), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11004) );
  INV_X1 U11910 ( .A(n11438), .ZN(n11461) );
  AOI21_X1 U11911 ( .B1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n20184), .A(
        n11421), .ZN(n11450) );
  AND2_X1 U11912 ( .A1(n11452), .A2(n11453), .ZN(n11421) );
  XNOR2_X1 U11913 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n10649) );
  NOR2_X1 U11914 ( .A1(n10762), .A2(n10143), .ZN(n10142) );
  AOI21_X1 U11915 ( .B1(n12628), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10455), 
        .ZN(n10456) );
  NAND2_X1 U11916 ( .A1(n9961), .A2(n9960), .ZN(n10431) );
  OAI21_X1 U11917 ( .B1(n12625), .B2(n10009), .A(n10006), .ZN(n10487) );
  NOR2_X1 U11918 ( .A1(n10008), .A2(n10007), .ZN(n10006) );
  INV_X1 U11919 ( .A(n10486), .ZN(n10007) );
  NOR2_X1 U11920 ( .A1(n10913), .A2(n12690), .ZN(n10008) );
  NOR2_X1 U11921 ( .A1(n10136), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10135) );
  INV_X1 U11922 ( .A(n12702), .ZN(n10868) );
  AOI21_X1 U11923 ( .B1(n19250), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A(
        n10597), .ZN(n10598) );
  AND2_X1 U11924 ( .A1(n19377), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(
        n10597) );
  AOI21_X1 U11925 ( .B1(n19647), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A(
        n16281), .ZN(n10528) );
  INV_X1 U11926 ( .A(n10641), .ZN(n12683) );
  AOI22_X1 U11927 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_2__4__SCAN_IN), .B1(
        n10353), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10404) );
  AND4_X1 U11928 ( .A1(n12645), .A2(n10419), .A3(n12644), .A4(n10443), .ZN(
        n10439) );
  AOI21_X1 U11929 ( .B1(n20944), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(
        n11742), .ZN(n11748) );
  NOR2_X1 U11930 ( .A1(n11930), .A2(n11927), .ZN(n11742) );
  NOR2_X1 U11931 ( .A1(n11945), .A2(n17244), .ZN(n11951) );
  NAND2_X1 U11932 ( .A1(n18094), .A2(n17153), .ZN(n11737) );
  INV_X1 U11933 ( .A(n11731), .ZN(n11733) );
  NAND2_X1 U11934 ( .A1(n14206), .A2(n10216), .ZN(n10215) );
  AND2_X1 U11935 ( .A1(n12169), .A2(n14141), .ZN(n14140) );
  INV_X1 U11936 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n12149) );
  NOR2_X1 U11937 ( .A1(n11252), .A2(n11251), .ZN(n11262) );
  NAND2_X1 U11938 ( .A1(n10130), .A2(n14349), .ZN(n10129) );
  INV_X1 U11939 ( .A(n14457), .ZN(n10130) );
  INV_X1 U11940 ( .A(n14361), .ZN(n10131) );
  INV_X1 U11941 ( .A(n14645), .ZN(n10207) );
  NOR2_X1 U11942 ( .A1(n14759), .A2(n14758), .ZN(n10119) );
  XNOR2_X1 U11943 ( .A(n11388), .B(n11377), .ZN(n12044) );
  NAND2_X1 U11944 ( .A1(n10127), .A2(n10126), .ZN(n10125) );
  INV_X1 U11945 ( .A(n13712), .ZN(n10127) );
  INV_X1 U11946 ( .A(n13779), .ZN(n10126) );
  INV_X1 U11947 ( .A(n10172), .ZN(n10170) );
  NAND2_X1 U11948 ( .A1(n11129), .A2(n10168), .ZN(n11473) );
  AND2_X1 U11949 ( .A1(n11135), .A2(n11176), .ZN(n10168) );
  OR2_X1 U11950 ( .A1(n11173), .A2(n11172), .ZN(n11259) );
  NAND2_X1 U11951 ( .A1(n11278), .A2(n11277), .ZN(n11466) );
  NAND2_X1 U11952 ( .A1(n10745), .A2(n10746), .ZN(n10764) );
  NAND2_X1 U11953 ( .A1(n10722), .A2(n10717), .ZN(n10139) );
  NAND2_X1 U11954 ( .A1(n10137), .A2(n10720), .ZN(n10136) );
  INV_X1 U11955 ( .A(n10139), .ZN(n10137) );
  INV_X1 U11956 ( .A(n10718), .ZN(n10140) );
  OR2_X1 U11957 ( .A1(n10487), .A2(n10488), .ZN(n10907) );
  INV_X1 U11958 ( .A(n14869), .ZN(n10953) );
  AOI21_X1 U11959 ( .B1(n13002), .B2(n10247), .A(n13031), .ZN(n10246) );
  INV_X1 U11960 ( .A(n14978), .ZN(n10247) );
  NOR2_X1 U11961 ( .A1(n10253), .A2(n10252), .ZN(n10251) );
  INV_X1 U11962 ( .A(n15005), .ZN(n10253) );
  AND2_X1 U11963 ( .A1(n12927), .A2(n10256), .ZN(n10255) );
  INV_X1 U11964 ( .A(n10257), .ZN(n10256) );
  AND2_X1 U11965 ( .A1(n14111), .A2(n13997), .ZN(n12927) );
  NAND4_X1 U11966 ( .A1(n10372), .A2(n10371), .A3(n10370), .A4(n10369), .ZN(
        n10373) );
  NAND2_X1 U11967 ( .A1(n10366), .A2(n9881), .ZN(n10374) );
  NAND2_X1 U11968 ( .A1(n9817), .A2(n12645), .ZN(n10433) );
  AND2_X1 U11969 ( .A1(n12669), .A2(n12681), .ZN(n12670) );
  INV_X1 U11970 ( .A(n13841), .ZN(n10928) );
  INV_X1 U11971 ( .A(n13842), .ZN(n10260) );
  NAND2_X1 U11972 ( .A1(n10265), .A2(n13640), .ZN(n10264) );
  INV_X1 U11973 ( .A(n13630), .ZN(n10265) );
  INV_X1 U11974 ( .A(n10496), .ZN(n10229) );
  AND2_X1 U11975 ( .A1(n14948), .A2(n10977), .ZN(n10266) );
  NOR2_X1 U11976 ( .A1(n14239), .A2(n15263), .ZN(n10235) );
  AND2_X1 U11977 ( .A1(n14873), .A2(n9870), .ZN(n15044) );
  AND2_X1 U11978 ( .A1(n12853), .A2(n9875), .ZN(n10226) );
  AND2_X1 U11979 ( .A1(n12825), .A2(n12822), .ZN(n10198) );
  INV_X1 U11980 ( .A(n15231), .ZN(n10048) );
  NAND2_X1 U11981 ( .A1(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15162) );
  INV_X1 U11982 ( .A(n14001), .ZN(n10941) );
  INV_X1 U11983 ( .A(n13965), .ZN(n10942) );
  OR2_X1 U11984 ( .A1(n10264), .A2(n13527), .ZN(n10263) );
  OR2_X1 U11985 ( .A1(n13922), .A2(n9982), .ZN(n9981) );
  INV_X1 U11986 ( .A(n10703), .ZN(n9982) );
  NAND2_X1 U11987 ( .A1(n10684), .A2(n10045), .ZN(n10044) );
  INV_X1 U11988 ( .A(n14902), .ZN(n10045) );
  NAND2_X1 U11989 ( .A1(n9995), .A2(n10862), .ZN(n10863) );
  INV_X1 U11990 ( .A(n14249), .ZN(n9996) );
  OR2_X1 U11991 ( .A1(n10521), .A2(n10525), .ZN(n10511) );
  NOR2_X1 U11992 ( .A1(n10520), .A2(n15536), .ZN(n10519) );
  OR2_X1 U11993 ( .A1(n10521), .A2(n10512), .ZN(n10507) );
  NAND3_X1 U11994 ( .A1(n15507), .A2(n10284), .A3(n10521), .ZN(n10533) );
  AND2_X1 U11995 ( .A1(n10510), .A2(n10521), .ZN(n19543) );
  AOI22_X1 U11996 ( .A1(n13601), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n10541), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10392) );
  NOR2_X1 U11997 ( .A1(n20860), .A2(n21012), .ZN(n17609) );
  NAND2_X1 U11998 ( .A1(n15727), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16299) );
  NAND2_X1 U11999 ( .A1(n11880), .A2(n17680), .ZN(n11899) );
  AND2_X1 U12000 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n11881), .ZN(
        n11882) );
  NOR2_X1 U12001 ( .A1(n11739), .A2(n18106), .ZN(n11926) );
  INV_X1 U12002 ( .A(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n20860) );
  NOR2_X1 U12003 ( .A1(n13713), .A2(n10125), .ZN(n13815) );
  NOR2_X1 U12004 ( .A1(n10111), .A2(n10110), .ZN(n13652) );
  AND2_X1 U12005 ( .A1(n11506), .A2(n11505), .ZN(n13651) );
  NAND2_X1 U12006 ( .A1(n13649), .A2(n12006), .ZN(n13711) );
  AND2_X1 U12007 ( .A1(n13514), .A2(n13513), .ZN(n19969) );
  NAND2_X1 U12008 ( .A1(n11596), .A2(n13621), .ZN(n13284) );
  AND2_X1 U12009 ( .A1(n12428), .A2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n12429) );
  OR2_X1 U12010 ( .A1(n12433), .A2(n12432), .ZN(n14339) );
  AND2_X1 U12011 ( .A1(n9915), .A2(n12409), .ZN(n10217) );
  NOR2_X1 U12012 ( .A1(n12383), .A2(n15748), .ZN(n12384) );
  NAND2_X1 U12013 ( .A1(n12384), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12427) );
  NAND2_X1 U12014 ( .A1(n14463), .A2(n10219), .ZN(n14456) );
  NAND2_X1 U12015 ( .A1(n12342), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12383) );
  AND2_X1 U12016 ( .A1(n14463), .A2(n14462), .ZN(n14464) );
  NOR2_X1 U12017 ( .A1(n12290), .A2(n15802), .ZN(n12291) );
  AND2_X1 U12018 ( .A1(n12274), .A2(n12273), .ZN(n14488) );
  NOR2_X1 U12019 ( .A1(n11409), .A2(n10041), .ZN(n14630) );
  OR2_X1 U12020 ( .A1(n14637), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10041) );
  AND2_X1 U12021 ( .A1(n12259), .A2(n12258), .ZN(n14547) );
  CLKBUF_X1 U12022 ( .A(n14486), .Z(n14487) );
  NOR2_X1 U12023 ( .A1(n21101), .A2(n12238), .ZN(n12257) );
  CLKBUF_X1 U12024 ( .A(n14372), .Z(n14373) );
  NOR2_X1 U12025 ( .A1(n12221), .A2(n15810), .ZN(n12222) );
  NAND2_X1 U12026 ( .A1(n12222), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12238) );
  NOR2_X1 U12027 ( .A1(n12188), .A2(n12187), .ZN(n12189) );
  NAND2_X1 U12028 ( .A1(n12189), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12221) );
  OR2_X1 U12029 ( .A1(n12121), .A2(n15830), .ZN(n12188) );
  NAND2_X1 U12030 ( .A1(n12164), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n12121) );
  INV_X1 U12031 ( .A(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n15830) );
  NOR2_X1 U12032 ( .A1(n12148), .A2(n12149), .ZN(n12164) );
  AND2_X1 U12033 ( .A1(n12091), .A2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n12092) );
  NAND2_X1 U12034 ( .A1(n12092), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n12148) );
  NAND2_X1 U12035 ( .A1(n12061), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n12062) );
  NOR2_X1 U12036 ( .A1(n21011), .A2(n12062), .ZN(n12091) );
  CLKBUF_X1 U12037 ( .A(n13971), .Z(n13972) );
  AND3_X1 U12038 ( .A1(n12060), .A2(n12059), .A3(n12058), .ZN(n13900) );
  NAND2_X1 U12039 ( .A1(n12038), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n12057) );
  INV_X1 U12040 ( .A(n12037), .ZN(n12038) );
  NAND2_X1 U12041 ( .A1(n12029), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12037) );
  OAI211_X1 U12042 ( .C1(n12028), .C2(n12168), .A(n12027), .B(n12026), .ZN(
        n13806) );
  CLKBUF_X1 U12043 ( .A(n13804), .Z(n13805) );
  AOI21_X1 U12044 ( .B1(n12024), .B2(n12130), .A(n12023), .ZN(n13776) );
  CLKBUF_X1 U12045 ( .A(n13709), .Z(n13775) );
  NAND2_X1 U12046 ( .A1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n12008) );
  NOR2_X1 U12047 ( .A1(n12008), .A2(n12007), .ZN(n12020) );
  INV_X1 U12048 ( .A(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12007) );
  AND2_X1 U12049 ( .A1(n13698), .A2(n13520), .ZN(n13621) );
  NAND2_X1 U12050 ( .A1(n11594), .A2(n11593), .ZN(n10108) );
  NOR3_X1 U12051 ( .A1(n14468), .A2(n10131), .A3(n14457), .ZN(n14363) );
  NOR2_X1 U12052 ( .A1(n10205), .A2(n10204), .ZN(n10203) );
  INV_X1 U12053 ( .A(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10204) );
  OAI21_X1 U12054 ( .B1(n10020), .B2(n10019), .A(n14636), .ZN(n14603) );
  INV_X1 U12055 ( .A(n14588), .ZN(n10020) );
  NAND2_X1 U12056 ( .A1(n15859), .A2(n9874), .ZN(n10019) );
  NOR2_X1 U12057 ( .A1(n14468), .A2(n14457), .ZN(n14458) );
  OR2_X1 U12058 ( .A1(n14474), .A2(n14466), .ZN(n14468) );
  NAND2_X1 U12059 ( .A1(n14484), .A2(n14472), .ZN(n14474) );
  NOR2_X1 U12060 ( .A1(n14491), .A2(n14482), .ZN(n14484) );
  NAND2_X1 U12061 ( .A1(n10119), .A2(n10118), .ZN(n14491) );
  INV_X1 U12062 ( .A(n14489), .ZN(n10118) );
  INV_X1 U12063 ( .A(n10119), .ZN(n14761) );
  OR2_X1 U12064 ( .A1(n14688), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14637) );
  AND2_X1 U12065 ( .A1(n14499), .A2(n14392), .ZN(n14390) );
  AND2_X1 U12066 ( .A1(n11554), .A2(n11553), .ZN(n14497) );
  OR2_X1 U12067 ( .A1(n14688), .A2(n15937), .ZN(n14653) );
  AND2_X1 U12068 ( .A1(n10134), .A2(n10133), .ZN(n10132) );
  INV_X1 U12069 ( .A(n14169), .ZN(n10133) );
  AND2_X1 U12070 ( .A1(n14186), .A2(n14180), .ZN(n14182) );
  NAND2_X1 U12071 ( .A1(n14186), .A2(n10134), .ZN(n14168) );
  AND2_X1 U12072 ( .A1(n11414), .A2(n11607), .ZN(n14677) );
  OR2_X1 U12073 ( .A1(n14128), .A2(n11539), .ZN(n14841) );
  NAND2_X1 U12074 ( .A1(n15898), .A2(n10015), .ZN(n10013) );
  NAND2_X1 U12075 ( .A1(n10015), .A2(n10018), .ZN(n10012) );
  AND3_X1 U12076 ( .A1(n11530), .A2(n11558), .A3(n11529), .ZN(n13975) );
  NOR2_X1 U12077 ( .A1(n13902), .A2(n9852), .ZN(n14057) );
  OR2_X1 U12078 ( .A1(n13902), .A2(n13901), .ZN(n13976) );
  AND3_X1 U12079 ( .A1(n11523), .A2(n11558), .A3(n11522), .ZN(n13886) );
  NAND2_X1 U12080 ( .A1(n11525), .A2(n11524), .ZN(n13902) );
  INV_X1 U12081 ( .A(n13886), .ZN(n11524) );
  INV_X1 U12082 ( .A(n15985), .ZN(n11525) );
  NOR2_X1 U12083 ( .A1(n13713), .A2(n10123), .ZN(n15983) );
  NAND2_X1 U12084 ( .A1(n10124), .A2(n13814), .ZN(n10123) );
  INV_X1 U12085 ( .A(n10125), .ZN(n10124) );
  AND2_X1 U12086 ( .A1(n11521), .A2(n11520), .ZN(n15982) );
  OR2_X1 U12087 ( .A1(n13713), .A2(n13712), .ZN(n13778) );
  INV_X1 U12088 ( .A(n14845), .ZN(n20066) );
  INV_X1 U12089 ( .A(n11620), .ZN(n11613) );
  OAI21_X1 U12090 ( .B1(n11234), .B2(n14284), .A(n11134), .ZN(n11144) );
  INV_X1 U12091 ( .A(n11225), .ZN(n9954) );
  INV_X1 U12092 ( .A(n11239), .ZN(n10036) );
  NAND2_X1 U12093 ( .A1(n11233), .A2(n10032), .ZN(n10031) );
  INV_X1 U12094 ( .A(n20147), .ZN(n20262) );
  INV_X1 U12095 ( .A(n11123), .ZN(n9949) );
  AND3_X1 U12096 ( .A1(n13477), .A2(n13476), .A3(n13519), .ZN(n15699) );
  OR2_X1 U12097 ( .A1(n13700), .A2(n20105), .ZN(n20379) );
  NAND2_X1 U12098 ( .A1(n20256), .A2(n10030), .ZN(n20351) );
  OR2_X1 U12099 ( .A1(n13700), .A2(n20765), .ZN(n20554) );
  AND2_X1 U12100 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n20147), .ZN(n20144) );
  OAI21_X1 U12101 ( .B1(n13727), .B2(n20795), .A(n15722), .ZN(n20147) );
  AOI21_X1 U12102 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n20551), .A(n20262), 
        .ZN(n20636) );
  AOI221_X1 U12103 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n10835), 
        .C1(n15664), .C2(n10835), .A(n10834), .ZN(n12582) );
  NOR2_X1 U12104 ( .A1(n10807), .A2(n10147), .ZN(n10146) );
  INV_X1 U12105 ( .A(n10800), .ZN(n10147) );
  NOR2_X1 U12106 ( .A1(n13222), .A2(n10089), .ZN(n13225) );
  NAND2_X1 U12107 ( .A1(n10742), .A2(n10741), .ZN(n10743) );
  NOR2_X1 U12108 ( .A1(n10140), .A2(n10136), .ZN(n10730) );
  AND2_X1 U12109 ( .A1(n10906), .A2(n10907), .ZN(n13588) );
  NAND2_X1 U12110 ( .A1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n13212) );
  NAND2_X1 U12111 ( .A1(n10954), .A2(n10953), .ZN(n15001) );
  NAND2_X1 U12112 ( .A1(n12891), .A2(n13793), .ZN(n10257) );
  OR2_X1 U12113 ( .A1(n12735), .A2(n12734), .ZN(n12890) );
  OR2_X1 U12114 ( .A1(n14261), .A2(n14235), .ZN(n16027) );
  XNOR2_X1 U12115 ( .A(n10248), .B(n13057), .ZN(n14970) );
  NAND2_X1 U12116 ( .A1(n14970), .A2(n14969), .ZN(n14968) );
  NAND2_X1 U12117 ( .A1(n14873), .A2(n9862), .ZN(n15061) );
  AND2_X1 U12118 ( .A1(n14873), .A2(n15330), .ZN(n15332) );
  INV_X1 U12119 ( .A(n14066), .ZN(n12823) );
  AND2_X1 U12120 ( .A1(n10428), .A2(n10443), .ZN(n13388) );
  NOR2_X1 U12121 ( .A1(n10190), .A2(n12701), .ZN(n10187) );
  INV_X1 U12122 ( .A(n13930), .ZN(n10190) );
  AND2_X1 U12123 ( .A1(n13345), .A2(n13344), .ZN(n13343) );
  INV_X1 U12124 ( .A(n12581), .ZN(n19835) );
  INV_X1 U12125 ( .A(n13208), .ZN(n14069) );
  INV_X1 U12126 ( .A(n10235), .ZN(n10233) );
  NAND2_X1 U12127 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n10232) );
  NOR2_X1 U12128 ( .A1(n15113), .A2(n15101), .ZN(n15102) );
  OR2_X1 U12129 ( .A1(n15126), .A2(n16049), .ZN(n15113) );
  NOR2_X1 U12130 ( .A1(n15146), .A2(n15138), .ZN(n15136) );
  NAND2_X1 U12131 ( .A1(n15136), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15126) );
  NAND2_X1 U12132 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n15151), .ZN(
        n15146) );
  NAND2_X1 U12133 ( .A1(n13211), .A2(n9866), .ZN(n15686) );
  AND2_X1 U12134 ( .A1(n13225), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13227) );
  AND2_X1 U12135 ( .A1(n13227), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13211) );
  NOR2_X1 U12136 ( .A1(n13893), .A2(n13913), .ZN(n13967) );
  NAND2_X1 U12137 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n13223), .ZN(
        n13222) );
  NAND2_X1 U12138 ( .A1(n13220), .A2(n9865), .ZN(n13221) );
  NOR2_X1 U12139 ( .A1(n14217), .A2(n13217), .ZN(n13220) );
  NAND2_X1 U12140 ( .A1(n13220), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n13219) );
  NOR2_X1 U12141 ( .A1(n13215), .A2(n14082), .ZN(n13218) );
  NAND2_X1 U12142 ( .A1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n13218), .ZN(
        n13217) );
  NAND2_X1 U12143 ( .A1(n13216), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13215) );
  OR2_X1 U12144 ( .A1(n13629), .A2(n10264), .ZN(n13641) );
  NOR2_X1 U12145 ( .A1(n13629), .A2(n13630), .ZN(n13639) );
  NOR2_X1 U12146 ( .A1(n13213), .A2(n16191), .ZN(n13216) );
  NOR2_X1 U12147 ( .A1(n14901), .A2(n13212), .ZN(n13214) );
  NAND2_X1 U12148 ( .A1(n13214), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n13213) );
  XNOR2_X1 U12149 ( .A(n14266), .B(n12847), .ZN(n16012) );
  AND2_X1 U12150 ( .A1(n14266), .A2(n14265), .ZN(n16017) );
  NAND2_X1 U12151 ( .A1(n10269), .A2(n10268), .ZN(n12553) );
  AND2_X1 U12152 ( .A1(n12532), .A2(n10144), .ZN(n10268) );
  AND2_X1 U12153 ( .A1(n14947), .A2(n14948), .ZN(n14950) );
  NAND2_X1 U12154 ( .A1(n15112), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15105) );
  INV_X1 U12155 ( .A(n14983), .ZN(n10259) );
  NOR2_X1 U12156 ( .A1(n10280), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9986) );
  OAI21_X1 U12157 ( .B1(n15167), .B2(n15168), .A(n10785), .ZN(n10794) );
  NAND2_X1 U12158 ( .A1(n12823), .A2(n10198), .ZN(n15382) );
  NAND2_X1 U12159 ( .A1(n10942), .A2(n10941), .ZN(n14114) );
  INV_X1 U12160 ( .A(n13851), .ZN(n10191) );
  OR2_X1 U12161 ( .A1(n13738), .A2(n10193), .ZN(n14019) );
  NOR2_X1 U12162 ( .A1(n9892), .A2(n10273), .ZN(n10272) );
  NOR2_X1 U12163 ( .A1(n15481), .A2(n10274), .ZN(n10273) );
  INV_X1 U12164 ( .A(n15479), .ZN(n10740) );
  NOR2_X1 U12165 ( .A1(n13629), .A2(n10261), .ZN(n13705) );
  NAND2_X1 U12166 ( .A1(n10262), .A2(n13572), .ZN(n10261) );
  INV_X1 U12167 ( .A(n10263), .ZN(n10262) );
  AND2_X1 U12168 ( .A1(n13705), .A2(n13704), .ZN(n13742) );
  NAND2_X1 U12169 ( .A1(n16171), .A2(n10886), .ZN(n14212) );
  NAND3_X1 U12170 ( .A1(n10066), .A2(n10876), .A3(n10236), .ZN(n10069) );
  OR2_X1 U12171 ( .A1(n10878), .A2(n12706), .ZN(n10876) );
  NAND2_X1 U12172 ( .A1(n10069), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13981) );
  OR2_X1 U12173 ( .A1(n12663), .A2(n12650), .ZN(n15400) );
  OR2_X1 U12174 ( .A1(n12663), .A2(n16252), .ZN(n13875) );
  NAND2_X1 U12175 ( .A1(n12862), .A2(n19798), .ZN(n12878) );
  INV_X1 U12176 ( .A(n10520), .ZN(n10286) );
  NOR2_X2 U12177 ( .A1(n10507), .A2(n14914), .ZN(n19284) );
  OR2_X1 U12178 ( .A1(n19804), .A2(n19786), .ZN(n19408) );
  NOR2_X2 U12179 ( .A1(n14069), .A2(n13941), .ZN(n19152) );
  NOR2_X2 U12180 ( .A1(n14070), .A2(n13941), .ZN(n19151) );
  OR2_X1 U12181 ( .A1(n19607), .A2(n19789), .ZN(n19615) );
  INV_X1 U12182 ( .A(n19151), .ZN(n19146) );
  INV_X1 U12183 ( .A(n19139), .ZN(n19148) );
  AOI21_X1 U12184 ( .B1(n11752), .B2(n11932), .A(n11931), .ZN(n11935) );
  INV_X1 U12185 ( .A(n17312), .ZN(n10071) );
  NAND2_X1 U12186 ( .A1(n18552), .A2(n11908), .ZN(n18528) );
  NOR2_X1 U12187 ( .A1(n16498), .A2(n16770), .ZN(n16491) );
  NOR2_X1 U12188 ( .A1(n16492), .A2(n16491), .ZN(n16490) );
  NOR2_X1 U12189 ( .A1(n17416), .A2(n16515), .ZN(n16514) );
  OR2_X1 U12190 ( .A1(n16569), .A2(n17487), .ZN(n16567) );
  NAND3_X1 U12191 ( .A1(n11717), .A2(n11716), .A3(n11715), .ZN(n17112) );
  AOI211_X1 U12192 ( .C1(n9819), .C2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A(
        n11714), .B(n11713), .ZN(n11715) );
  AOI21_X1 U12193 ( .B1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B2(n9812), .A(n11808), .ZN(n11809) );
  NOR2_X1 U12194 ( .A1(n11832), .A2(n10151), .ZN(n10150) );
  AND2_X1 U12195 ( .A1(n11857), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11823) );
  AOI22_X1 U12196 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n11821), .B2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11822) );
  OR3_X1 U12197 ( .A1(n11664), .A2(n11663), .A3(n10079), .ZN(n18746) );
  AOI21_X1 U12198 ( .B1(n10072), .B2(n18589), .A(n18744), .ZN(n17259) );
  INV_X1 U12199 ( .A(n17309), .ZN(n17260) );
  NOR2_X1 U12200 ( .A1(n16307), .A2(n16479), .ZN(n11635) );
  NAND2_X1 U12201 ( .A1(n11638), .A2(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n16307) );
  NAND2_X1 U12202 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10182) );
  NOR2_X1 U12203 ( .A1(n17389), .A2(n9876), .ZN(n11638) );
  NOR3_X1 U12204 ( .A1(n17438), .A2(n17412), .A3(n17410), .ZN(n17366) );
  NAND2_X1 U12205 ( .A1(n17453), .A2(n10295), .ZN(n17442) );
  NOR2_X1 U12206 ( .A1(n17442), .A2(n17745), .ZN(n17409) );
  AND2_X1 U12207 ( .A1(n17532), .A2(n10179), .ZN(n17453) );
  AND2_X1 U12208 ( .A1(n10180), .A2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10179) );
  AND3_X1 U12209 ( .A1(n17609), .A2(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n17559) );
  AND3_X1 U12210 ( .A1(n10177), .A2(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A3(
        n10176), .ZN(n17558) );
  NOR2_X1 U12211 ( .A1(n17693), .A2(n17665), .ZN(n10176) );
  NOR2_X1 U12212 ( .A1(n17694), .A2(n17693), .ZN(n17684) );
  NAND2_X1 U12213 ( .A1(n15667), .A2(n15666), .ZN(n15726) );
  OR2_X1 U12214 ( .A1(n15668), .A2(n11899), .ZN(n11906) );
  NAND2_X1 U12215 ( .A1(n17378), .A2(n17379), .ZN(n17377) );
  NOR2_X1 U12216 ( .A1(n11898), .A2(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15667) );
  NOR2_X1 U12217 ( .A1(n11781), .A2(n11780), .ZN(n16315) );
  NOR2_X1 U12218 ( .A1(n17930), .A2(n17934), .ZN(n17557) );
  NAND2_X1 U12219 ( .A1(n17941), .A2(n17606), .ZN(n17930) );
  AND2_X1 U12220 ( .A1(n17630), .A2(n17608), .ZN(n10165) );
  INV_X1 U12221 ( .A(n18561), .ZN(n18540) );
  NAND2_X1 U12222 ( .A1(n10154), .A2(n10152), .ZN(n17702) );
  AOI211_X1 U12223 ( .C1(n11934), .C2(n11933), .A(n11932), .B(n11931), .ZN(
        n18535) );
  NAND2_X1 U12224 ( .A1(n17967), .A2(n18554), .ZN(n16345) );
  XNOR2_X1 U12225 ( .A(n17250), .B(n18708), .ZN(n17740) );
  NOR2_X1 U12226 ( .A1(n11739), .A2(n11914), .ZN(n11908) );
  NOR2_X1 U12227 ( .A1(n11941), .A2(n11922), .ZN(n18532) );
  INV_X1 U12228 ( .A(n18555), .ZN(n18552) );
  NAND2_X1 U12229 ( .A1(n18758), .A2(n14225), .ZN(n18561) );
  INV_X1 U12230 ( .A(n18528), .ZN(n18558) );
  INV_X1 U12231 ( .A(n18542), .ZN(n18557) );
  INV_X1 U12232 ( .A(n18746), .ZN(n18094) );
  NOR2_X2 U12233 ( .A1(n11655), .A2(n11654), .ZN(n18100) );
  NOR2_X1 U12234 ( .A1(n11697), .A2(n11696), .ZN(n18112) );
  NOR2_X1 U12235 ( .A1(n11727), .A2(n11726), .ZN(n18117) );
  INV_X1 U12236 ( .A(n17112), .ZN(n18128) );
  INV_X1 U12237 ( .A(n16306), .ZN(n18444) );
  INV_X1 U12238 ( .A(n13284), .ZN(n13282) );
  AND2_X1 U12239 ( .A1(n14430), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n19932) );
  NOR2_X1 U12240 ( .A1(n12507), .A2(n12509), .ZN(n15781) );
  INV_X1 U12241 ( .A(n19934), .ZN(n19955) );
  INV_X1 U12242 ( .A(n15881), .ZN(n14184) );
  NOR2_X1 U12243 ( .A1(n14558), .A2(n13492), .ZN(n14163) );
  AND2_X1 U12244 ( .A1(n13485), .A2(n13520), .ZN(n14529) );
  INV_X1 U12245 ( .A(n14163), .ZN(n14155) );
  INV_X1 U12246 ( .A(n20035), .ZN(n13569) );
  XNOR2_X1 U12247 ( .A(n12491), .B(n12513), .ZN(n14257) );
  INV_X1 U12248 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n15810) );
  INV_X1 U12249 ( .A(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n15916) );
  NAND2_X1 U12250 ( .A1(n19863), .A2(n13623), .ZN(n15915) );
  AND2_X1 U12251 ( .A1(n15915), .A2(n20037), .ZN(n15911) );
  INV_X1 U12252 ( .A(n15915), .ZN(n20038) );
  AND2_X1 U12253 ( .A1(n13621), .A2(n15709), .ZN(n20043) );
  XNOR2_X1 U12254 ( .A(n12497), .B(n12496), .ZN(n14447) );
  OR2_X1 U12255 ( .A1(n12523), .A2(n9941), .ZN(n9940) );
  NAND2_X1 U12256 ( .A1(n9945), .A2(n9944), .ZN(n9943) );
  NAND2_X1 U12257 ( .A1(n14578), .A2(n10301), .ZN(n14579) );
  NAND2_X1 U12258 ( .A1(n14617), .A2(n10173), .ZN(n14611) );
  OAI21_X1 U12259 ( .B1(n11409), .B2(n14645), .A(n14644), .ZN(n14797) );
  NAND2_X1 U12260 ( .A1(n10037), .A2(n11394), .ZN(n14005) );
  OR2_X1 U12261 ( .A1(n13954), .A2(n11395), .ZN(n10037) );
  INV_X1 U12262 ( .A(n20095), .ZN(n20077) );
  NOR2_X1 U12263 ( .A1(n11620), .A2(n11604), .ZN(n20062) );
  AND2_X1 U12264 ( .A1(n20099), .A2(n10100), .ZN(n20084) );
  XNOR2_X1 U12265 ( .A(n10113), .B(n13523), .ZN(n13542) );
  NAND2_X1 U12266 ( .A1(n10109), .A2(n10114), .ZN(n10113) );
  INV_X1 U12267 ( .A(n10111), .ZN(n10109) );
  OAI21_X1 U12268 ( .B1(n9828), .B2(n11423), .A(n11183), .ZN(n20039) );
  INV_X1 U12269 ( .A(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20440) );
  CLKBUF_X1 U12271 ( .A(n13654), .Z(n13655) );
  INV_X1 U12272 ( .A(n20581), .ZN(n20767) );
  OAI22_X1 U12273 ( .A1(n20116), .A2(n20115), .B1(n20383), .B2(n20259), .ZN(
        n20149) );
  OR2_X1 U12274 ( .A1(n20221), .A2(n20434), .ZN(n20250) );
  INV_X1 U12275 ( .A(n20278), .ZN(n20281) );
  INV_X1 U12276 ( .A(n20304), .ZN(n20307) );
  OAI22_X1 U12277 ( .A1(n20318), .A2(n20317), .B1(n20316), .B2(n20584), .ZN(
        n20344) );
  NOR2_X1 U12278 ( .A1(n20551), .A2(n20350), .ZN(n20372) );
  OR2_X1 U12279 ( .A1(n20351), .A2(n20434), .ZN(n20377) );
  INV_X1 U12280 ( .A(n20371), .ZN(n20405) );
  OAI211_X1 U12281 ( .C1(n20620), .C2(n20590), .A(n20589), .B(n20588), .ZN(
        n20624) );
  INV_X1 U12282 ( .A(n20441), .ZN(n20632) );
  INV_X1 U12283 ( .A(n20523), .ZN(n20633) );
  INV_X1 U12284 ( .A(n20526), .ZN(n20644) );
  INV_X1 U12285 ( .A(n20454), .ZN(n20649) );
  INV_X1 U12286 ( .A(n20529), .ZN(n20650) );
  INV_X1 U12287 ( .A(n20458), .ZN(n20655) );
  INV_X1 U12288 ( .A(n20532), .ZN(n20656) );
  INV_X1 U12289 ( .A(n20535), .ZN(n20662) );
  INV_X1 U12290 ( .A(n20333), .ZN(n20667) );
  INV_X1 U12291 ( .A(n20538), .ZN(n20668) );
  INV_X1 U12292 ( .A(n20337), .ZN(n20673) );
  INV_X1 U12293 ( .A(n20541), .ZN(n20674) );
  INV_X1 U12294 ( .A(n20472), .ZN(n20679) );
  INV_X1 U12295 ( .A(n20547), .ZN(n20680) );
  NAND3_X1 U12296 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n11192), .A3(n13698), 
        .ZN(n15722) );
  INV_X1 U12297 ( .A(P1_STATE2_REG_1__SCAN_IN), .ZN(n16000) );
  NAND2_X1 U12298 ( .A1(n16000), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20689) );
  INV_X1 U12299 ( .A(n10820), .ZN(n10822) );
  NAND2_X1 U12300 ( .A1(n18929), .A2(n9886), .ZN(n15687) );
  NAND2_X1 U12301 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n12616), .ZN(n10091) );
  NAND2_X1 U12302 ( .A1(n14289), .A2(n10983), .ZN(n10092) );
  NOR2_X1 U12303 ( .A1(n14905), .A2(n9927), .ZN(n14906) );
  OR3_X1 U12304 ( .A1(n19847), .A2(n16276), .A3(n13231), .ZN(n18954) );
  INV_X1 U12305 ( .A(n18831), .ZN(n18958) );
  OR2_X1 U12306 ( .A1(n13845), .A2(n13844), .ZN(n13909) );
  NAND2_X1 U12307 ( .A1(n10254), .A2(n12891), .ZN(n13747) );
  OR2_X1 U12308 ( .A1(n12720), .A2(n12719), .ZN(n13575) );
  INV_X1 U12309 ( .A(n15009), .ZN(n14965) );
  INV_X2 U12310 ( .A(n14993), .ZN(n15006) );
  NAND2_X1 U12311 ( .A1(n10244), .A2(n14944), .ZN(n14956) );
  INV_X1 U12312 ( .A(n13083), .ZN(n14962) );
  NOR2_X1 U12313 ( .A1(n14979), .A2(n14978), .ZN(n14977) );
  NOR2_X1 U12314 ( .A1(n14988), .A2(n13002), .ZN(n14979) );
  NAND2_X1 U12315 ( .A1(n10195), .A2(n9906), .ZN(n13500) );
  OR2_X1 U12316 ( .A1(n13395), .A2(n12708), .ZN(n10195) );
  AND2_X1 U12317 ( .A1(n13387), .A2(n13386), .ZN(n15083) );
  OR2_X1 U12318 ( .A1(n13608), .A2(n13385), .ZN(n13387) );
  AND2_X1 U12319 ( .A1(n18969), .A2(n19009), .ZN(n18995) );
  AND2_X1 U12320 ( .A1(n15084), .A2(n14071), .ZN(n19013) );
  NOR2_X1 U12321 ( .A1(n15523), .A2(n13336), .ZN(n19158) );
  AND2_X1 U12322 ( .A1(n15083), .A2(n10238), .ZN(n19005) );
  INV_X1 U12323 ( .A(n15083), .ZN(n19004) );
  AND2_X1 U12324 ( .A1(n19016), .A2(n19721), .ZN(n19057) );
  OR2_X1 U12325 ( .A1(n19081), .A2(n13288), .ZN(n13429) );
  NAND2_X1 U12326 ( .A1(n10234), .A2(n10231), .ZN(n12617) );
  NOR2_X1 U12327 ( .A1(n10233), .A2(n10232), .ZN(n10231) );
  INV_X1 U12328 ( .A(n15247), .ZN(n15402) );
  INV_X1 U12329 ( .A(P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16144) );
  INV_X1 U12330 ( .A(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n14217) );
  AND2_X1 U12331 ( .A1(n10222), .A2(n10221), .ZN(n16173) );
  NAND2_X1 U12332 ( .A1(n10000), .A2(n14078), .ZN(n10222) );
  NAND2_X1 U12333 ( .A1(n9999), .A2(n10882), .ZN(n10221) );
  INV_X1 U12334 ( .A(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n14082) );
  INV_X1 U12335 ( .A(n19104), .ZN(n16174) );
  XNOR2_X1 U12336 ( .A(n12627), .B(n12626), .ZN(n16013) );
  NAND2_X1 U12337 ( .A1(n15018), .A2(n16209), .ZN(n14243) );
  XNOR2_X1 U12338 ( .A(n12533), .B(n10310), .ZN(n14248) );
  OR2_X1 U12339 ( .A1(n14947), .A2(n14954), .ZN(n16048) );
  AND2_X1 U12340 ( .A1(n10064), .A2(n15184), .ZN(n10063) );
  INV_X1 U12341 ( .A(n15202), .ZN(n10064) );
  NAND2_X1 U12342 ( .A1(n10065), .A2(n15184), .ZN(n15203) );
  NAND2_X1 U12343 ( .A1(n10046), .A2(n10050), .ZN(n15230) );
  NAND2_X1 U12344 ( .A1(n15251), .A2(n10053), .ZN(n10046) );
  AND2_X1 U12345 ( .A1(n15247), .A2(n12618), .ZN(n15404) );
  NAND2_X1 U12346 ( .A1(n10055), .A2(n15248), .ZN(n15239) );
  NAND2_X1 U12347 ( .A1(n10056), .A2(n10057), .ZN(n10055) );
  NAND2_X1 U12348 ( .A1(n15167), .A2(n15466), .ZN(n15454) );
  INV_X1 U12349 ( .A(n15160), .ZN(n15469) );
  NAND2_X1 U12350 ( .A1(n10279), .A2(n10278), .ZN(n15480) );
  OR2_X1 U12351 ( .A1(n15514), .A2(n15511), .ZN(n15397) );
  NAND2_X1 U12352 ( .A1(n13921), .A2(n13922), .ZN(n9980) );
  AND2_X1 U12353 ( .A1(n9998), .A2(n13866), .ZN(n13918) );
  NAND2_X1 U12354 ( .A1(n16219), .A2(n10521), .ZN(n16220) );
  NOR2_X1 U12355 ( .A1(n13396), .A2(n12688), .ZN(n13830) );
  OR2_X1 U12356 ( .A1(n12663), .A2(n12662), .ZN(n16222) );
  NAND2_X1 U12357 ( .A1(n13875), .A2(n15400), .ZN(n15514) );
  INV_X1 U12358 ( .A(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19823) );
  INV_X1 U12359 ( .A(n19158), .ZN(n19818) );
  INV_X1 U12360 ( .A(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n19814) );
  INV_X1 U12361 ( .A(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n19796) );
  XNOR2_X1 U12362 ( .A(n13363), .B(n13362), .ZN(n19808) );
  NAND2_X1 U12363 ( .A1(n10521), .A2(n15541), .ZN(n13607) );
  INV_X1 U12364 ( .A(n19788), .ZN(n19407) );
  INV_X1 U12365 ( .A(n19179), .ZN(n19182) );
  NOR2_X1 U12366 ( .A1(n19408), .A2(n19347), .ZN(n19207) );
  NOR2_X1 U12367 ( .A1(n19347), .A2(n19468), .ZN(n19268) );
  INV_X1 U12368 ( .A(n19303), .ZN(n19315) );
  INV_X1 U12369 ( .A(n19325), .ZN(n19343) );
  AND2_X1 U12370 ( .A1(n19470), .A2(n19319), .ZN(n19382) );
  INV_X1 U12371 ( .A(n19430), .ZN(n19431) );
  OAI21_X1 U12372 ( .B1(n19445), .B2(n19462), .A(n19648), .ZN(n19464) );
  NOR2_X1 U12373 ( .A1(n19556), .A2(n19468), .ZN(n19531) );
  NOR2_X1 U12374 ( .A1(n19607), .A2(n19555), .ZN(n19587) );
  INV_X1 U12375 ( .A(n19685), .ZN(n19590) );
  INV_X1 U12376 ( .A(n19587), .ZN(n19605) );
  INV_X1 U12377 ( .A(n19699), .ZN(n19606) );
  OAI21_X1 U12378 ( .B1(n19620), .B2(n19619), .A(n19618), .ZN(n19642) );
  INV_X1 U12379 ( .A(n19565), .ZN(n19663) );
  AND2_X1 U12380 ( .A1(n13334), .A2(n19148), .ZN(n19661) );
  INV_X1 U12381 ( .A(n19571), .ZN(n19668) );
  AND2_X1 U12382 ( .A1(n19124), .A2(n19148), .ZN(n19666) );
  INV_X1 U12383 ( .A(n19578), .ZN(n19677) );
  INV_X1 U12384 ( .A(n19615), .ZN(n19700) );
  INV_X1 U12385 ( .A(n19436), .ZN(n19701) );
  AND2_X1 U12386 ( .A1(n16285), .A2(n16288), .ZN(n16294) );
  INV_X1 U12387 ( .A(P2_STATE2_REG_2__SCAN_IN), .ZN(n19842) );
  INV_X1 U12388 ( .A(P2_STATE2_REG_3__SCAN_IN), .ZN(n19798) );
  INV_X1 U12389 ( .A(n10073), .ZN(n16449) );
  NAND2_X1 U12390 ( .A1(n18741), .A2(n11935), .ZN(n17313) );
  NOR2_X1 U12391 ( .A1(n16499), .A2(n17384), .ZN(n16498) );
  AND2_X1 U12392 ( .A1(n16782), .A2(n11756), .ZN(n16518) );
  INV_X1 U12393 ( .A(n16782), .ZN(n16802) );
  INV_X1 U12394 ( .A(n16593), .ZN(n10185) );
  INV_X1 U12395 ( .A(n16810), .ZN(n16796) );
  NAND4_X1 U12396 ( .A1(n18741), .A2(n16313), .A3(n18746), .A4(n15742), .ZN(
        n17107) );
  AND2_X1 U12397 ( .A1(P3_EAX_REG_27__SCAN_IN), .A2(n17133), .ZN(n17132) );
  NOR2_X1 U12398 ( .A1(n17139), .A2(n17266), .ZN(n17133) );
  NAND2_X1 U12399 ( .A1(n17140), .A2(P3_EAX_REG_25__SCAN_IN), .ZN(n17139) );
  NOR2_X1 U12400 ( .A1(n17187), .A2(n10081), .ZN(n17150) );
  INV_X1 U12401 ( .A(n17160), .ZN(n10082) );
  NOR2_X1 U12402 ( .A1(n17280), .A2(n17175), .ZN(n17170) );
  NAND2_X1 U12403 ( .A1(n17191), .A2(P3_EAX_REG_16__SCAN_IN), .ZN(n17187) );
  NAND3_X1 U12404 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17221), .A3(n17196), 
        .ZN(n17197) );
  NAND2_X1 U12405 ( .A1(n17251), .A2(n17228), .ZN(n17222) );
  NOR2_X1 U12406 ( .A1(n17296), .A2(n17222), .ZN(n17221) );
  INV_X1 U12407 ( .A(n17247), .ZN(n17252) );
  INV_X1 U12408 ( .A(n17243), .ZN(n17255) );
  CLKBUF_X1 U12409 ( .A(n17361), .Z(n17349) );
  INV_X1 U12410 ( .A(n11633), .ZN(n11632) );
  NAND2_X1 U12411 ( .A1(n17532), .A2(n10180), .ZN(n17484) );
  NAND2_X1 U12412 ( .A1(n17532), .A2(n10297), .ZN(n17517) );
  INV_X1 U12413 ( .A(n17582), .ZN(n17531) );
  NOR2_X1 U12414 ( .A1(n17581), .A2(n11630), .ZN(n17532) );
  NAND2_X1 U12415 ( .A1(n11629), .A2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n11630) );
  INV_X1 U12416 ( .A(n17583), .ZN(n11629) );
  NOR2_X1 U12417 ( .A1(n17550), .A2(n17564), .ZN(n17896) );
  NAND2_X1 U12418 ( .A1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n17583) );
  INV_X1 U12419 ( .A(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n21012) );
  INV_X1 U12420 ( .A(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n17665) );
  NAND2_X1 U12421 ( .A1(n10177), .A2(n10175), .ZN(n17664) );
  NOR2_X1 U12422 ( .A1(n10178), .A2(n17693), .ZN(n10175) );
  INV_X1 U12423 ( .A(n17750), .ZN(n17708) );
  INV_X1 U12424 ( .A(P3_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n17693) );
  INV_X1 U12425 ( .A(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n17745) );
  OAI21_X1 U12426 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18740), .A(n16450), 
        .ZN(n17750) );
  INV_X1 U12427 ( .A(n17742), .ZN(n17755) );
  NAND2_X1 U12428 ( .A1(n17434), .A2(n11892), .ZN(n17427) );
  INV_X1 U12429 ( .A(n11879), .ZN(n10162) );
  INV_X1 U12430 ( .A(n10163), .ZN(n17688) );
  INV_X1 U12431 ( .A(n10157), .ZN(n17717) );
  AND2_X1 U12432 ( .A1(n10157), .A2(n10156), .ZN(n17715) );
  NAND2_X1 U12433 ( .A1(n10159), .A2(n10158), .ZN(n10157) );
  NOR2_X1 U12434 ( .A1(n9820), .A2(n18073), .ZN(n18055) );
  INV_X1 U12435 ( .A(n10159), .ZN(n17725) );
  NOR2_X2 U12436 ( .A1(n11908), .A2(n18555), .ZN(n18568) );
  INV_X1 U12437 ( .A(n18061), .ZN(n18073) );
  INV_X1 U12438 ( .A(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18576) );
  AOI211_X1 U12439 ( .C1(n18741), .C2(n18565), .A(n18093), .B(n14227), .ZN(
        n18728) );
  INV_X1 U12440 ( .A(P3_STATE2_REG_2__SCAN_IN), .ZN(n18603) );
  INV_X1 U12441 ( .A(P3_STATE2_REG_0__SCAN_IN), .ZN(n18604) );
  INV_X1 U12443 ( .A(n14320), .ZN(n14448) );
  NAND2_X1 U12444 ( .A1(n10104), .A2(n10102), .ZN(P1_U2842) );
  NAND2_X1 U12445 ( .A1(n14320), .A2(n15856), .ZN(n10104) );
  AOI21_X1 U12446 ( .B1(n14572), .B2(n19964), .A(n10103), .ZN(n10102) );
  NOR2_X1 U12447 ( .A1(n19968), .A2(n14449), .ZN(n10103) );
  AOI21_X1 U12448 ( .B1(n14993), .B2(n10521), .A(n13510), .ZN(n13511) );
  AOI21_X1 U12449 ( .B1(n16018), .B2(n19104), .A(n12547), .ZN(n12549) );
  AND2_X1 U12450 ( .A1(n19104), .A2(n10521), .ZN(n10249) );
  INV_X1 U12451 ( .A(n14277), .ZN(n14278) );
  AOI21_X1 U12452 ( .B1(n16018), .B2(n16219), .A(n14275), .ZN(n14276) );
  NAND2_X1 U12453 ( .A1(n9857), .A2(n16227), .ZN(n9993) );
  AOI211_X1 U12454 ( .C1(n16472), .C2(n16788), .A(n16471), .B(n16470), .ZN(
        n16475) );
  OAI211_X1 U12455 ( .C1(P3_EAX_REG_31__SCAN_IN), .C2(n17113), .A(n10075), .B(
        n10074), .ZN(P3_U2704) );
  NAND2_X1 U12456 ( .A1(n17185), .A2(BUF2_REG_31__SCAN_IN), .ZN(n10074) );
  NAND2_X1 U12457 ( .A1(n10076), .A2(P3_EAX_REG_31__SCAN_IN), .ZN(n10075) );
  INV_X1 U12458 ( .A(n17140), .ZN(n17143) );
  AND2_X1 U12459 ( .A1(n16317), .A2(n16318), .ZN(n10148) );
  AND2_X1 U12460 ( .A1(n16355), .A2(n16356), .ZN(n10149) );
  INV_X2 U12461 ( .A(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n16232) );
  AND2_X1 U12463 ( .A1(n10225), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n9848) );
  AND2_X1 U12464 ( .A1(n10954), .A2(n9861), .ZN(n9849) );
  NOR2_X1 U12465 ( .A1(n12688), .A2(n10186), .ZN(n10189) );
  AND2_X1 U12466 ( .A1(n12668), .A2(n19798), .ZN(n12684) );
  INV_X2 U12467 ( .A(n9983), .ZN(n19134) );
  INV_X1 U12468 ( .A(n11819), .ZN(n15599) );
  CLKBUF_X3 U12469 ( .A(n12668), .Z(n13334) );
  NAND2_X1 U12470 ( .A1(n11409), .A2(n14645), .ZN(n14644) );
  AND2_X1 U12471 ( .A1(n13172), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n12725) );
  AND2_X1 U12472 ( .A1(n14463), .A2(n9915), .ZN(n14350) );
  NAND2_X1 U12473 ( .A1(n10227), .A2(n10226), .ZN(n9850) );
  NOR2_X1 U12474 ( .A1(n13738), .A2(n9912), .ZN(n9851) );
  OR2_X1 U12475 ( .A1(n13975), .A2(n13901), .ZN(n9852) );
  AND4_X1 U12476 ( .A1(n11118), .A2(n11117), .A3(n11116), .A4(n11115), .ZN(
        n9853) );
  AND2_X1 U12477 ( .A1(n9981), .A2(n13983), .ZN(n9854) );
  OAI21_X1 U12478 ( .B1(n14077), .B2(n10001), .A(n9896), .ZN(n16171) );
  INV_X1 U12479 ( .A(n10227), .ZN(n14211) );
  AND2_X1 U12480 ( .A1(n10297), .A2(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n9855) );
  AND2_X1 U12481 ( .A1(n12644), .A2(n12588), .ZN(n9856) );
  INV_X1 U12482 ( .A(n12635), .ZN(n10446) );
  AND2_X1 U12483 ( .A1(n10196), .A2(n12724), .ZN(n9858) );
  AND2_X1 U12484 ( .A1(n10687), .A2(n10044), .ZN(n9859) );
  AND2_X1 U12485 ( .A1(n14101), .A2(n14118), .ZN(n9860) );
  INV_X1 U12486 ( .A(P2_STATE2_REG_0__SCAN_IN), .ZN(n10983) );
  INV_X1 U12487 ( .A(n13396), .ZN(n10188) );
  INV_X1 U12488 ( .A(n15249), .ZN(n10057) );
  AND2_X1 U12489 ( .A1(n10953), .A2(n10258), .ZN(n9861) );
  AND2_X1 U12490 ( .A1(n10200), .A2(n10199), .ZN(n9862) );
  AND2_X1 U12491 ( .A1(n10198), .A2(n15082), .ZN(n9863) );
  AND2_X1 U12492 ( .A1(n10941), .A2(n9964), .ZN(n9864) );
  NOR2_X1 U12493 ( .A1(n13738), .A2(n9919), .ZN(n13849) );
  AND2_X1 U12494 ( .A1(n10087), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n9865) );
  AND2_X1 U12495 ( .A1(n10085), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n9866) );
  AND2_X1 U12496 ( .A1(n10210), .A2(n11339), .ZN(n9867) );
  AND2_X1 U12497 ( .A1(n9861), .A2(n14992), .ZN(n9868) );
  AND2_X1 U12498 ( .A1(n9864), .A2(n14098), .ZN(n9869) );
  AND2_X1 U12499 ( .A1(n9862), .A2(n9934), .ZN(n9870) );
  AND2_X1 U12500 ( .A1(n9863), .A2(n13243), .ZN(n9871) );
  INV_X1 U12501 ( .A(n9837), .ZN(n13044) );
  INV_X1 U12502 ( .A(n10540), .ZN(n13009) );
  AND3_X1 U12503 ( .A1(n10188), .A2(n10189), .A3(n13835), .ZN(n9872) );
  NAND2_X1 U12504 ( .A1(n10226), .A2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n9873) );
  NOR2_X1 U12505 ( .A1(n11412), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n9874) );
  AND2_X1 U12506 ( .A1(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n9875) );
  INV_X1 U12507 ( .A(n18929), .ZN(n18917) );
  AND2_X1 U12508 ( .A1(n10353), .A2(n16232), .ZN(n12953) );
  OR3_X1 U12509 ( .A1(n17438), .A2(n17412), .A3(n10182), .ZN(n9876) );
  OR2_X1 U12510 ( .A1(n15033), .A2(n15034), .ZN(n9877) );
  AND2_X1 U12511 ( .A1(n10072), .A2(n10071), .ZN(n9878) );
  NAND2_X1 U12512 ( .A1(n10875), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10878) );
  OAI21_X1 U12514 ( .B1(n10825), .B2(n10271), .A(n10270), .ZN(n12533) );
  NAND2_X1 U12515 ( .A1(n14685), .A2(n11397), .ZN(n14661) );
  OR2_X1 U12516 ( .A1(n14147), .A2(n10215), .ZN(n14205) );
  AND2_X1 U12517 ( .A1(n10519), .A2(n14914), .ZN(n9879) );
  AND3_X1 U12518 ( .A1(n10150), .A2(n11831), .A3(n11829), .ZN(n9880) );
  INV_X1 U12519 ( .A(n11812), .ZN(n17068) );
  INV_X1 U12520 ( .A(n11857), .ZN(n11812) );
  AND2_X1 U12521 ( .A1(n10365), .A2(n10364), .ZN(n9881) );
  NAND4_X1 U12522 ( .A1(n10793), .A2(n10792), .A3(n15177), .A4(n10791), .ZN(
        n9882) );
  XOR2_X1 U12523 ( .A(n12615), .B(n12548), .Z(n9883) );
  NAND2_X1 U12524 ( .A1(n10029), .A2(n11258), .ZN(n11987) );
  OR2_X1 U12525 ( .A1(P2_EBX_REG_11__SCAN_IN), .A2(n10743), .ZN(n9884) );
  AND4_X1 U12526 ( .A1(n11114), .A2(n11113), .A3(n11112), .A4(n11111), .ZN(
        n9885) );
  NAND2_X1 U12527 ( .A1(n17519), .A2(n17604), .ZN(n17434) );
  NAND2_X1 U12528 ( .A1(n14463), .A2(n10217), .ZN(n14337) );
  OR2_X1 U12529 ( .A1(n15684), .A2(n15685), .ZN(n9886) );
  NAND2_X1 U12530 ( .A1(n10495), .A2(n10494), .ZN(n10493) );
  AND3_X1 U12531 ( .A1(n11683), .A2(n11684), .A3(n11685), .ZN(n9887) );
  NAND3_X1 U12532 ( .A1(n10452), .A2(n10450), .A3(n10451), .ZN(n10467) );
  OR3_X1 U12533 ( .A1(n14468), .A2(n10131), .A3(n10129), .ZN(n9888) );
  AND2_X1 U12534 ( .A1(n15098), .A2(n10145), .ZN(n9889) );
  AND3_X1 U12535 ( .A1(n10244), .A2(n14944), .A3(n10243), .ZN(n9890) );
  NAND2_X1 U12536 ( .A1(n13113), .A2(n13112), .ZN(n14944) );
  AND2_X1 U12537 ( .A1(n9977), .A2(n15099), .ZN(n9891) );
  INV_X1 U12538 ( .A(n11871), .ZN(n10158) );
  INV_X1 U12539 ( .A(n10468), .ZN(n10485) );
  NAND2_X1 U12540 ( .A1(n9983), .A2(n10427), .ZN(n10442) );
  INV_X1 U12541 ( .A(n10442), .ZN(n10420) );
  NAND2_X1 U12542 ( .A1(n10374), .A2(n10373), .ZN(n10428) );
  AOI21_X1 U12543 ( .B1(n14321), .B2(n14323), .A(n14322), .ZN(n14572) );
  OR2_X1 U12544 ( .A1(n10311), .A2(n10740), .ZN(n9892) );
  AND4_X1 U12545 ( .A1(n15222), .A2(n15186), .A3(n15206), .A4(n15181), .ZN(
        n9893) );
  OR2_X1 U12546 ( .A1(n9882), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9894) );
  AND2_X1 U12547 ( .A1(n12522), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n9895) );
  NAND2_X1 U12548 ( .A1(n10245), .A2(n10246), .ZN(n10248) );
  AND2_X1 U12549 ( .A1(n16172), .A2(n9966), .ZN(n9896) );
  OR2_X1 U12550 ( .A1(n14147), .A2(n10214), .ZN(n9897) );
  NAND2_X1 U12551 ( .A1(n14338), .A2(n14300), .ZN(n14321) );
  INV_X1 U12552 ( .A(n15536), .ZN(n15507) );
  NAND2_X1 U12553 ( .A1(n10502), .A2(n10503), .ZN(n15536) );
  INV_X1 U12554 ( .A(n15093), .ZN(n9987) );
  NOR2_X1 U12555 ( .A1(n9991), .A2(n9990), .ZN(n9898) );
  NOR2_X2 U12556 ( .A1(n12660), .A2(n13584), .ZN(n9899) );
  NOR2_X1 U12557 ( .A1(n15123), .A2(n9989), .ZN(n9900) );
  AND2_X1 U12558 ( .A1(n10040), .A2(n11407), .ZN(n9901) );
  AND2_X1 U12559 ( .A1(n13267), .A2(n12498), .ZN(n9902) );
  AND2_X1 U12560 ( .A1(n10684), .A2(n15176), .ZN(n9903) );
  AND2_X1 U12561 ( .A1(n20104), .A2(n11326), .ZN(n9904) );
  AND2_X1 U12562 ( .A1(n10493), .A2(n10504), .ZN(n18950) );
  INV_X1 U12563 ( .A(n18950), .ZN(n10284) );
  INV_X1 U12564 ( .A(n12644), .ZN(n19124) );
  AND2_X1 U12565 ( .A1(n10360), .A2(n10359), .ZN(n12644) );
  OR2_X1 U12566 ( .A1(n13267), .A2(n11491), .ZN(n9905) );
  INV_X1 U12567 ( .A(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n10178) );
  AND2_X2 U12568 ( .A1(n11005), .A2(n13673), .ZN(n11356) );
  INV_X1 U12569 ( .A(n12685), .ZN(n12695) );
  OR2_X1 U12570 ( .A1(n15176), .A2(n12819), .ZN(n9906) );
  NOR2_X1 U12571 ( .A1(n11886), .A2(n17988), .ZN(n17647) );
  NAND2_X1 U12572 ( .A1(n11291), .A2(n11290), .ZN(n20104) );
  INV_X1 U12573 ( .A(n20104), .ZN(n10030) );
  NAND2_X1 U12574 ( .A1(n10043), .A2(n14902), .ZN(n13868) );
  AND2_X1 U12575 ( .A1(n11501), .A2(n20122), .ZN(n11588) );
  NOR2_X1 U12576 ( .A1(n13883), .A2(n13900), .ZN(n9907) );
  INV_X1 U12577 ( .A(n10443), .ZN(n10238) );
  NAND2_X1 U12578 ( .A1(n13849), .A2(n15413), .ZN(n14066) );
  AND2_X1 U12579 ( .A1(n13211), .A2(n10085), .ZN(n9908) );
  AND2_X1 U12580 ( .A1(n13220), .A2(n10087), .ZN(n9909) );
  NAND2_X1 U12581 ( .A1(n11500), .A2(n13516), .ZN(n9910) );
  NOR2_X1 U12582 ( .A1(n15157), .A2(n15156), .ZN(n15155) );
  AND2_X1 U12583 ( .A1(n12823), .A2(n9871), .ZN(n13242) );
  NOR2_X1 U12584 ( .A1(n13743), .A2(n13795), .ZN(n13796) );
  NAND2_X1 U12585 ( .A1(n10260), .A2(n10928), .ZN(n13840) );
  NAND2_X1 U12586 ( .A1(n14101), .A2(n10251), .ZN(n14996) );
  AND2_X1 U12587 ( .A1(n10942), .A2(n9864), .ZN(n9911) );
  INV_X1 U12588 ( .A(n10441), .ZN(n12586) );
  NOR2_X1 U12589 ( .A1(n13574), .A2(n10257), .ZN(n13791) );
  OR2_X1 U12590 ( .A1(n10193), .A2(n14020), .ZN(n9912) );
  OAI21_X1 U12591 ( .B1(n10794), .B2(n9986), .A(n9984), .ZN(n15325) );
  NAND2_X1 U12592 ( .A1(n9980), .A2(n10703), .ZN(n13982) );
  NAND2_X1 U12593 ( .A1(n10275), .A2(n10272), .ZN(n15465) );
  AND2_X1 U12594 ( .A1(n10279), .A2(n10728), .ZN(n14213) );
  INV_X1 U12595 ( .A(n10746), .ZN(n10143) );
  AND3_X1 U12596 ( .A1(n14250), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A3(
        n10685), .ZN(n9913) );
  OR3_X1 U12597 ( .A1(n13222), .A2(n10090), .A3(n15253), .ZN(n9914) );
  NAND2_X1 U12598 ( .A1(n12823), .A2(n12822), .ZN(n14065) );
  AND2_X1 U12599 ( .A1(n10218), .A2(n10219), .ZN(n9915) );
  AND2_X1 U12600 ( .A1(n12823), .A2(n9863), .ZN(n9916) );
  AND2_X1 U12601 ( .A1(n9869), .A2(n13236), .ZN(n9917) );
  INV_X1 U12602 ( .A(n15248), .ZN(n10054) );
  INV_X1 U12603 ( .A(n10053), .ZN(n10052) );
  NOR2_X1 U12604 ( .A1(n10054), .A2(n15178), .ZN(n10053) );
  AND2_X1 U12605 ( .A1(n10942), .A2(n9869), .ZN(n13235) );
  OR2_X1 U12606 ( .A1(n12762), .A2(n12761), .ZN(n13793) );
  INV_X1 U12607 ( .A(n9964), .ZN(n14113) );
  OR2_X1 U12608 ( .A1(n10945), .A2(n9965), .ZN(n9964) );
  AND2_X1 U12609 ( .A1(n10171), .A2(n11608), .ZN(n9918) );
  NAND2_X1 U12610 ( .A1(n14873), .A2(n10200), .ZN(n15058) );
  INV_X1 U12611 ( .A(n10141), .ZN(n10742) );
  NAND2_X1 U12612 ( .A1(n10718), .A2(n10135), .ZN(n10141) );
  OR2_X1 U12613 ( .A1(n9912), .A2(n10191), .ZN(n9919) );
  AND2_X1 U12614 ( .A1(n18920), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n9920) );
  AND2_X1 U12615 ( .A1(n13242), .A2(n14872), .ZN(n14873) );
  NAND2_X1 U12616 ( .A1(n10954), .A2(n9868), .ZN(n14982) );
  AND2_X1 U12617 ( .A1(n10142), .A2(n10748), .ZN(n9921) );
  AND2_X1 U12618 ( .A1(n10579), .A2(n10612), .ZN(n9922) );
  NAND2_X1 U12619 ( .A1(n10073), .A2(n11910), .ZN(n10072) );
  AND2_X1 U12620 ( .A1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n9923) );
  AND2_X1 U12621 ( .A1(n9858), .A2(n14888), .ZN(n9924) );
  AND2_X1 U12622 ( .A1(n10928), .A2(n10932), .ZN(n9925) );
  INV_X1 U12623 ( .A(P1_EBX_REG_1__SCAN_IN), .ZN(n10117) );
  NOR2_X1 U12624 ( .A1(n20771), .A2(n20109), .ZN(n9926) );
  INV_X1 U12625 ( .A(n19962), .ZN(n15856) );
  INV_X1 U12626 ( .A(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n9963) );
  NAND2_X1 U12627 ( .A1(n13395), .A2(n9906), .ZN(n10194) );
  NAND2_X1 U12628 ( .A1(n10188), .A2(n10189), .ZN(n13831) );
  AND2_X1 U12629 ( .A1(n10194), .A2(n9858), .ZN(n14047) );
  NOR2_X1 U12630 ( .A1(n10533), .A2(n14914), .ZN(n19513) );
  NOR2_X1 U12631 ( .A1(n13629), .A2(n10263), .ZN(n13528) );
  NAND2_X1 U12632 ( .A1(n13742), .A2(n13741), .ZN(n13743) );
  NAND2_X1 U12633 ( .A1(n12586), .A2(n19114), .ZN(n12660) );
  XNOR2_X1 U12634 ( .A(n13343), .B(n12674), .ZN(n13717) );
  AND2_X1 U12635 ( .A1(n10521), .A2(n18949), .ZN(n9927) );
  INV_X1 U12636 ( .A(n15466), .ZN(n10060) );
  NOR2_X1 U12637 ( .A1(n10533), .A2(n19105), .ZN(n19377) );
  INV_X1 U12638 ( .A(n10184), .ZN(n16615) );
  NAND2_X1 U12639 ( .A1(n10733), .A2(n9983), .ZN(n12555) );
  NAND2_X1 U12640 ( .A1(n10286), .A2(n10522), .ZN(n19190) );
  INV_X1 U12642 ( .A(n11126), .ZN(n9950) );
  AND2_X1 U12643 ( .A1(n10163), .A2(n10162), .ZN(n9928) );
  INV_X1 U12644 ( .A(n10192), .ZN(n13801) );
  OR2_X1 U12645 ( .A1(n13738), .A2(n12780), .ZN(n10192) );
  OR2_X1 U12646 ( .A1(n10208), .A2(n13900), .ZN(n9929) );
  OR2_X1 U12647 ( .A1(n10682), .A2(n10681), .ZN(n12696) );
  AND2_X1 U12648 ( .A1(n10251), .A2(n10250), .ZN(n9930) );
  NOR2_X1 U12649 ( .A1(n14253), .A2(n10249), .ZN(n9931) );
  AND2_X1 U12650 ( .A1(n9868), .A2(n10259), .ZN(n9932) );
  AND2_X1 U12651 ( .A1(n10266), .A2(n12621), .ZN(n9933) );
  INV_X1 U12652 ( .A(n19108), .ZN(n19087) );
  INV_X1 U12653 ( .A(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n10100) );
  NOR2_X2 U12654 ( .A1(n16315), .A2(n11899), .ZN(n17649) );
  INV_X1 U12655 ( .A(n17649), .ZN(n17604) );
  NAND2_X1 U12656 ( .A1(n12835), .A2(n12834), .ZN(n9934) );
  AND2_X1 U12657 ( .A1(n10243), .A2(n14945), .ZN(n9935) );
  NAND2_X1 U12658 ( .A1(n17532), .A2(n9855), .ZN(n10181) );
  NAND2_X1 U12659 ( .A1(n14763), .A2(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(
        n9936) );
  INV_X1 U12660 ( .A(n14118), .ZN(n10252) );
  INV_X1 U12661 ( .A(n14601), .ZN(n10205) );
  INV_X1 U12662 ( .A(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n10009) );
  INV_X1 U12663 ( .A(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n10167) );
  INV_X1 U12664 ( .A(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n9939) );
  INV_X1 U12665 ( .A(P3_STATE2_REG_3__SCAN_IN), .ZN(n18696) );
  NOR3_X2 U12666 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n9805), .A3(
        n18233), .ZN(n18162) );
  NOR3_X2 U12667 ( .A1(n9805), .A2(n20944), .A3(n18233), .ZN(n18205) );
  NOR3_X2 U12668 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n9805), .A3(
        n18277), .ZN(n18249) );
  NOR3_X2 U12669 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n9805), .A3(
        n18371), .ZN(n18340) );
  OAI22_X2 U12670 ( .A1(n20121), .A2(n20120), .B1(n21054), .B2(n20119), .ZN(
        n20596) );
  AOI22_X2 U12671 ( .A1(DATAI_17_), .A2(n20143), .B1(BUF1_REG_17__SCAN_IN), 
        .B2(n20142), .ZN(n20599) );
  NOR3_X2 U12672 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n9805), .A3(
        n18323), .ZN(n18294) );
  NOR2_X4 U12673 ( .A1(n11119), .A2(n20798), .ZN(n20747) );
  NAND2_X1 U12674 ( .A1(n12543), .A2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10909) );
  INV_X2 U12675 ( .A(n12625), .ZN(n12543) );
  AOI22_X2 U12676 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n20142), .B1(DATAI_16_), 
        .B2(n20143), .ZN(n20595) );
  INV_X1 U12677 ( .A(n20120), .ZN(n20142) );
  INV_X1 U12678 ( .A(n20119), .ZN(n20143) );
  NOR2_X2 U12679 ( .A1(n19129), .A2(n19139), .ZN(n19671) );
  OAI21_X1 U12680 ( .B1(n9947), .B2(n9939), .A(n9937), .ZN(n9946) );
  NAND3_X1 U12681 ( .A1(n9943), .A2(n9942), .A3(n9940), .ZN(n14260) );
  NAND2_X1 U12682 ( .A1(n12524), .A2(n9939), .ZN(n9941) );
  NAND2_X1 U12683 ( .A1(n9895), .A2(n12524), .ZN(n9942) );
  INV_X1 U12684 ( .A(n9946), .ZN(n9945) );
  INV_X1 U12685 ( .A(n14296), .ZN(n9947) );
  NAND3_X1 U12686 ( .A1(n9905), .A2(n11125), .A3(n11124), .ZN(n9948) );
  NAND4_X4 U12687 ( .A1(n11014), .A2(n11012), .A3(n11013), .A4(n11011), .ZN(
        n11127) );
  NAND2_X2 U12688 ( .A1(n9950), .A2(n9949), .ZN(n14280) );
  INV_X1 U12689 ( .A(n20380), .ZN(n9955) );
  NAND2_X1 U12690 ( .A1(n9956), .A2(n11386), .ZN(n11226) );
  OAI21_X2 U12691 ( .B1(n11989), .B2(n11990), .A(n11227), .ZN(n11256) );
  NAND2_X2 U12692 ( .A1(n11208), .A2(n11207), .ZN(n11990) );
  NOR2_X1 U12693 ( .A1(n11225), .A2(n11219), .ZN(n9952) );
  NAND2_X1 U12694 ( .A1(n11225), .A2(n11219), .ZN(n9953) );
  INV_X1 U12695 ( .A(n9957), .ZN(n11191) );
  NAND2_X2 U12696 ( .A1(n11145), .A2(n9957), .ZN(n14282) );
  NAND2_X1 U12697 ( .A1(n11190), .A2(n9957), .ZN(n20153) );
  INV_X2 U12698 ( .A(n11414), .ZN(n14636) );
  OAI211_X2 U12699 ( .C1(n15859), .C2(n10205), .A(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .B(n10202), .ZN(n14589) );
  NAND3_X1 U12700 ( .A1(n14685), .A2(n10174), .A3(n11404), .ZN(n10040) );
  AND3_X4 U12701 ( .A1(n9959), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A3(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n10353) );
  NOR2_X1 U12702 ( .A1(n10983), .A2(n9959), .ZN(n10224) );
  AND2_X2 U12703 ( .A1(n9961), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n10477) );
  NOR2_X2 U12704 ( .A1(n10481), .A2(n9962), .ZN(n10497) );
  NOR2_X2 U12705 ( .A1(n12625), .A2(n9963), .ZN(n9962) );
  NOR2_X1 U12706 ( .A1(n12625), .A2(n15387), .ZN(n9965) );
  NAND2_X1 U12707 ( .A1(n10492), .A2(n10491), .ZN(n10285) );
  OR2_X2 U12708 ( .A1(n10872), .A2(n10871), .ZN(n10884) );
  NAND3_X1 U12709 ( .A1(n10616), .A2(n9967), .A3(n9996), .ZN(n9995) );
  NAND3_X1 U12710 ( .A1(n10616), .A2(n9967), .A3(n9903), .ZN(n10042) );
  NAND3_X1 U12711 ( .A1(n10616), .A2(n9967), .A3(n15176), .ZN(n10043) );
  INV_X2 U12712 ( .A(n10867), .ZN(n9967) );
  AND3_X2 U12713 ( .A1(n10580), .A2(n10613), .A3(n9922), .ZN(n10867) );
  AND2_X2 U12714 ( .A1(n14212), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10227) );
  NAND4_X1 U12715 ( .A1(n9970), .A2(n9969), .A3(n9968), .A4(n19087), .ZN(n9994) );
  INV_X1 U12716 ( .A(n15099), .ZN(n9976) );
  NAND2_X1 U12717 ( .A1(n13921), .A2(n9854), .ZN(n9978) );
  NAND2_X1 U12718 ( .A1(n9978), .A2(n9979), .ZN(n14080) );
  XNOR2_X1 U12719 ( .A(n10867), .B(n12697), .ZN(n10864) );
  INV_X1 U12720 ( .A(n12588), .ZN(n10432) );
  NAND2_X2 U12721 ( .A1(n9983), .A2(n9817), .ZN(n12588) );
  INV_X2 U12722 ( .A(n10428), .ZN(n9983) );
  AND2_X1 U12723 ( .A1(n9985), .A2(n9893), .ZN(n9984) );
  OR3_X1 U12724 ( .A1(n9991), .A2(n9990), .A3(n9989), .ZN(n15122) );
  INV_X1 U12725 ( .A(n9988), .ZN(n15094) );
  NAND3_X1 U12726 ( .A1(n10283), .A2(n10282), .A3(n9900), .ZN(n9988) );
  INV_X1 U12727 ( .A(n15132), .ZN(n9989) );
  INV_X1 U12728 ( .A(n10282), .ZN(n9990) );
  INV_X1 U12729 ( .A(n10283), .ZN(n9991) );
  INV_X1 U12730 ( .A(n10492), .ZN(n9992) );
  NAND2_X1 U12731 ( .A1(n15268), .A2(n9993), .ZN(P2_U3018) );
  NAND2_X1 U12732 ( .A1(n15108), .A2(n9994), .ZN(P2_U2986) );
  XNOR2_X1 U12733 ( .A(n9997), .B(n14249), .ZN(n16224) );
  NAND3_X2 U12734 ( .A1(n9998), .A2(n13917), .A3(n13866), .ZN(n10877) );
  NAND2_X2 U12735 ( .A1(n10866), .A2(n10865), .ZN(n13866) );
  INV_X1 U12736 ( .A(n10877), .ZN(n10067) );
  INV_X2 U12737 ( .A(n10447), .ZN(n12668) );
  NAND2_X1 U12738 ( .A1(n10447), .A2(n10416), .ZN(n12562) );
  NAND2_X1 U12739 ( .A1(n10325), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10002) );
  NAND2_X1 U12740 ( .A1(n10320), .A2(n16232), .ZN(n10003) );
  NAND2_X1 U12741 ( .A1(n10335), .A2(n16232), .ZN(n10004) );
  NAND2_X1 U12742 ( .A1(n10330), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10005) );
  NAND2_X2 U12743 ( .A1(n10890), .A2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15110) );
  NAND2_X2 U12744 ( .A1(n10025), .A2(n10024), .ZN(n11409) );
  OR2_X2 U12745 ( .A1(n11256), .A2(n11257), .ZN(n10029) );
  INV_X2 U12746 ( .A(n10029), .ZN(n10220) );
  INV_X1 U12747 ( .A(n11232), .ZN(n10033) );
  NAND2_X1 U12748 ( .A1(n10034), .A2(n11239), .ZN(n11270) );
  NAND2_X1 U12749 ( .A1(n11233), .A2(n11232), .ZN(n10034) );
  NAND2_X1 U12750 ( .A1(n10033), .A2(n11239), .ZN(n10035) );
  OAI21_X2 U12751 ( .B1(n11409), .B2(n11411), .A(n14636), .ZN(n15859) );
  NAND2_X1 U12752 ( .A1(n10042), .A2(n9859), .ZN(n13921) );
  NAND2_X1 U12753 ( .A1(n10275), .A2(n10061), .ZN(n15167) );
  NAND2_X2 U12754 ( .A1(n10500), .A2(n10493), .ZN(n10503) );
  NAND2_X1 U12755 ( .A1(n10067), .A2(n10068), .ZN(n10066) );
  INV_X1 U12756 ( .A(n10879), .ZN(n10068) );
  OAI21_X1 U12757 ( .B1(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n10069), .A(
        n13981), .ZN(n16179) );
  NAND3_X1 U12758 ( .A1(n11665), .A2(n11666), .A3(n10080), .ZN(n10079) );
  NAND2_X2 U12759 ( .A1(n10503), .A2(n10476), .ZN(n10499) );
  AND2_X2 U12760 ( .A1(n10476), .A2(n10461), .ZN(n10500) );
  NAND3_X1 U12761 ( .A1(n10082), .A2(P3_EAX_REG_22__SCAN_IN), .A3(
        P3_EAX_REG_17__SCAN_IN), .ZN(n10081) );
  NAND2_X1 U12762 ( .A1(n10863), .A2(n10864), .ZN(n13865) );
  AOI21_X2 U12763 ( .B1(n15744), .B2(n15743), .A(n18595), .ZN(n17111) );
  AND2_X2 U12764 ( .A1(n15160), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16146) );
  INV_X2 U12765 ( .A(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n18713) );
  NAND3_X1 U12766 ( .A1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .A3(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10089) );
  NOR2_X1 U12767 ( .A1(n13222), .A2(n15253), .ZN(n13224) );
  INV_X1 U12768 ( .A(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n10090) );
  NAND2_X1 U12769 ( .A1(n11996), .A2(n11183), .ZN(n10097) );
  NAND2_X1 U12770 ( .A1(n13626), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n11216) );
  OAI21_X1 U12771 ( .B1(n13523), .B2(n13516), .A(n10114), .ZN(n10110) );
  NOR2_X1 U12772 ( .A1(n11586), .A2(P1_EBX_REG_1__SCAN_IN), .ZN(n10115) );
  NOR2_X1 U12773 ( .A1(n12493), .A2(n10117), .ZN(n10116) );
  INV_X1 U12774 ( .A(n13902), .ZN(n10120) );
  NAND2_X1 U12775 ( .A1(n10120), .A2(n10121), .ZN(n14128) );
  NAND2_X1 U12776 ( .A1(n14186), .A2(n10132), .ZN(n14498) );
  NOR2_X1 U12777 ( .A1(n10140), .A2(n10138), .ZN(n10724) );
  INV_X1 U12778 ( .A(n10717), .ZN(n10138) );
  NAND2_X1 U12779 ( .A1(n10745), .A2(n9921), .ZN(n10759) );
  NAND2_X1 U12780 ( .A1(n9987), .A2(n10271), .ZN(n10144) );
  NAND2_X1 U12781 ( .A1(n10801), .A2(n10800), .ZN(n10808) );
  NOR2_X2 U12782 ( .A1(n17400), .A2(n11897), .ZN(n11898) );
  OAI21_X1 U12783 ( .B1(n16357), .B2(n17555), .A(n10148), .ZN(P3_U2799) );
  OAI21_X1 U12784 ( .B1(n16357), .B2(n17909), .A(n10149), .ZN(P3_U2831) );
  INV_X1 U12785 ( .A(n11828), .ZN(n10151) );
  INV_X1 U12786 ( .A(n17716), .ZN(n10156) );
  NAND2_X1 U12787 ( .A1(n17716), .A2(n10153), .ZN(n10152) );
  NAND2_X1 U12788 ( .A1(n10159), .A2(n10155), .ZN(n10154) );
  NOR2_X1 U12789 ( .A1(n11873), .A2(n11871), .ZN(n10155) );
  XNOR2_X1 U12790 ( .A(n11878), .B(n11877), .ZN(n17689) );
  NOR2_X2 U12791 ( .A1(n17587), .A2(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n17542) );
  NAND2_X1 U12792 ( .A1(n17434), .A2(n10166), .ZN(n17419) );
  INV_X1 U12793 ( .A(n17419), .ZN(n17426) );
  NAND2_X1 U12794 ( .A1(n10170), .A2(n10169), .ZN(n11603) );
  AND2_X1 U12795 ( .A1(n10170), .A2(n11475), .ZN(n13271) );
  NAND2_X1 U12796 ( .A1(n10172), .A2(n20122), .ZN(n10171) );
  INV_X1 U12797 ( .A(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n10173) );
  INV_X1 U12798 ( .A(n10181), .ZN(n17495) );
  NAND3_X1 U12799 ( .A1(n10188), .A2(n10189), .A3(n10187), .ZN(n13929) );
  NAND2_X1 U12800 ( .A1(n10194), .A2(n9924), .ZN(n15485) );
  INV_X1 U12801 ( .A(n10201), .ZN(n11497) );
  OR2_X1 U12802 ( .A1(n10201), .A2(n11187), .ZN(n11188) );
  OAI21_X2 U12803 ( .B1(n11132), .B2(n10201), .A(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11234) );
  NOR2_X2 U12804 ( .A1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n13667) );
  NAND2_X1 U12805 ( .A1(n15860), .A2(n10203), .ZN(n10202) );
  MUX2_X1 U12806 ( .A(n14636), .B(n14637), .S(n14644), .Z(n14638) );
  NOR2_X2 U12807 ( .A1(n13883), .A2(n9929), .ZN(n13971) );
  AND2_X2 U12808 ( .A1(n13971), .A2(n14060), .ZN(n14058) );
  INV_X1 U12809 ( .A(n13973), .ZN(n10208) );
  NAND2_X1 U12810 ( .A1(n11340), .A2(n11339), .ZN(n11365) );
  NOR2_X1 U12811 ( .A1(n14147), .A2(n14166), .ZN(n14165) );
  INV_X1 U12812 ( .A(n14166), .ZN(n10216) );
  NAND2_X1 U12813 ( .A1(n9904), .A2(n10220), .ZN(n11342) );
  NAND2_X1 U12814 ( .A1(n10220), .A2(n20104), .ZN(n11325) );
  AND2_X2 U12815 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13594) );
  NAND2_X1 U12816 ( .A1(n10467), .A2(n10224), .ZN(n10223) );
  NAND2_X1 U12817 ( .A1(n10456), .A2(n10223), .ZN(n10460) );
  CLKBUF_X1 U12818 ( .A(n10227), .Z(n10225) );
  NOR2_X1 U12819 ( .A1(n15110), .A2(n10230), .ZN(n12615) );
  INV_X1 U12820 ( .A(n15110), .ZN(n10234) );
  NAND2_X1 U12821 ( .A1(n10521), .A2(n10284), .ZN(n10532) );
  NAND3_X1 U12822 ( .A1(n10877), .A2(n10879), .A3(n10878), .ZN(n10236) );
  INV_X1 U12823 ( .A(n10460), .ZN(n10457) );
  NAND3_X1 U12824 ( .A1(n10244), .A2(n9935), .A3(n14944), .ZN(n10241) );
  INV_X1 U12825 ( .A(n13113), .ZN(n10240) );
  NAND2_X1 U12826 ( .A1(n13135), .A2(n14945), .ZN(n10242) );
  NAND2_X1 U12827 ( .A1(n14988), .A2(n10247), .ZN(n10245) );
  NAND2_X1 U12828 ( .A1(n10521), .A2(n12881), .ZN(n12865) );
  INV_X1 U12829 ( .A(n13574), .ZN(n10254) );
  NAND2_X1 U12830 ( .A1(n10954), .A2(n9932), .ZN(n14985) );
  NAND2_X1 U12831 ( .A1(n10260), .A2(n9925), .ZN(n13893) );
  NAND2_X1 U12832 ( .A1(n14947), .A2(n10266), .ZN(n12620) );
  NAND2_X1 U12833 ( .A1(n14947), .A2(n9933), .ZN(n12627) );
  NAND2_X1 U12834 ( .A1(n10825), .A2(n10270), .ZN(n10269) );
  NAND2_X1 U12835 ( .A1(n14080), .A2(n10276), .ZN(n10275) );
  NAND2_X1 U12836 ( .A1(n10580), .A2(n10579), .ZN(n10615) );
  NAND2_X1 U12837 ( .A1(n10613), .A2(n10612), .ZN(n10614) );
  INV_X1 U12838 ( .A(n10281), .ZN(n10280) );
  NAND2_X1 U12839 ( .A1(n15143), .A2(n15301), .ZN(n10282) );
  OAI21_X1 U12840 ( .B1(n15143), .B2(n15301), .A(n15144), .ZN(n10283) );
  NAND3_X1 U12841 ( .A1(n10906), .A2(n10285), .A3(n10284), .ZN(n10520) );
  NAND2_X1 U12842 ( .A1(n14504), .A2(n10287), .ZN(n14506) );
  NAND2_X1 U12843 ( .A1(n15173), .A2(n16132), .ZN(n15175) );
  AND2_X2 U12844 ( .A1(n13667), .A2(n13673), .ZN(n11153) );
  CLKBUF_X1 U12845 ( .A(n14058), .Z(n14124) );
  NAND2_X1 U12846 ( .A1(n9899), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n10430) );
  INV_X2 U12847 ( .A(n13668), .ZN(n12468) );
  NAND2_X1 U12848 ( .A1(n15210), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n15195) );
  NOR2_X1 U12849 ( .A1(n11127), .A2(n11180), .ZN(n13480) );
  CLKBUF_X1 U12850 ( .A(n13883), .Z(n13899) );
  XNOR2_X1 U12851 ( .A(n11296), .B(n13756), .ZN(n13753) );
  NAND2_X1 U12852 ( .A1(n11365), .A2(n11366), .ZN(n12034) );
  AND3_X4 U12853 ( .A1(n10315), .A2(n15554), .A3(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n10401) );
  NAND2_X1 U12854 ( .A1(n10519), .A2(n19105), .ZN(n19252) );
  XNOR2_X1 U12855 ( .A(n12617), .B(n12616), .ZN(n14292) );
  NAND2_X1 U12856 ( .A1(n19129), .A2(n12644), .ZN(n12595) );
  AND2_X1 U12857 ( .A1(n10596), .A2(n10595), .ZN(n10599) );
  AND2_X1 U12858 ( .A1(n14529), .A2(n14503), .ZN(n10287) );
  AND2_X1 U12859 ( .A1(n10806), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10288) );
  OR2_X1 U12860 ( .A1(n9883), .A2(n19092), .ZN(n10289) );
  AND2_X1 U12861 ( .A1(n13184), .A2(n13183), .ZN(n10290) );
  AND2_X1 U12862 ( .A1(n12586), .A2(n10843), .ZN(n10291) );
  AND2_X1 U12863 ( .A1(n17996), .A2(n17604), .ZN(n10292) );
  AND2_X1 U12864 ( .A1(n10442), .A2(n16281), .ZN(n10293) );
  INV_X1 U12865 ( .A(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15664) );
  OR2_X1 U12866 ( .A1(n11771), .A2(n11770), .ZN(P3_U2640) );
  AND2_X1 U12867 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10295) );
  INV_X1 U12868 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12616) );
  INV_X1 U12869 ( .A(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12548) );
  INV_X1 U12870 ( .A(n18682), .ZN(n18755) );
  AND2_X1 U12871 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10297) );
  AND2_X1 U12872 ( .A1(n11414), .A2(n14601), .ZN(n10298) );
  INV_X1 U12873 ( .A(n12684), .ZN(n12710) );
  INV_X1 U12874 ( .A(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n21011) );
  INV_X1 U12875 ( .A(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12524) );
  OR2_X1 U12876 ( .A1(n11627), .A2(n14568), .ZN(n10300) );
  AND2_X1 U12877 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n10301) );
  INV_X1 U12878 ( .A(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n17561) );
  NOR2_X1 U12879 ( .A1(n20066), .A2(n20084), .ZN(n20070) );
  AND2_X1 U12880 ( .A1(n13601), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n10302) );
  INV_X1 U12881 ( .A(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n13690) );
  AND2_X1 U12882 ( .A1(n12668), .A2(n12644), .ZN(n10303) );
  AND2_X1 U12883 ( .A1(n10389), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10304) );
  OR3_X1 U12884 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n17457), .ZN(n10305) );
  INV_X1 U12885 ( .A(n16315), .ZN(n11904) );
  AND2_X1 U12886 ( .A1(n12323), .A2(n12322), .ZN(n10306) );
  INV_X1 U12887 ( .A(n12452), .ZN(n12484) );
  INV_X1 U12888 ( .A(n14350), .ZN(n14359) );
  NOR2_X1 U12889 ( .A1(n17533), .A2(n17708), .ZN(n17452) );
  INV_X1 U12890 ( .A(n12672), .ZN(n12709) );
  INV_X1 U12891 ( .A(n10514), .ZN(n19412) );
  INV_X1 U12892 ( .A(n19252), .ZN(n19250) );
  INV_X1 U12893 ( .A(P2_STATE2_REG_1__SCAN_IN), .ZN(n15527) );
  AND2_X1 U12894 ( .A1(n13080), .A2(n13109), .ZN(n10308) );
  AND2_X1 U12895 ( .A1(n12551), .A2(n12550), .ZN(n10309) );
  AND2_X1 U12896 ( .A1(n12550), .A2(n12532), .ZN(n10310) );
  AND2_X1 U12897 ( .A1(n18898), .A2(n10737), .ZN(n10311) );
  NOR2_X1 U12898 ( .A1(n15155), .A2(n10288), .ZN(n15143) );
  AND4_X1 U12899 ( .A1(n11091), .A2(n11090), .A3(n11089), .A4(n11088), .ZN(
        n10312) );
  AND2_X2 U12900 ( .A1(n13667), .A2(n13687), .ZN(n11283) );
  AND4_X1 U12901 ( .A1(n11095), .A2(n11094), .A3(n11093), .A4(n11092), .ZN(
        n10314) );
  NAND2_X1 U12902 ( .A1(n19647), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(
        n10587) );
  AND2_X1 U12903 ( .A1(n11433), .A2(n11432), .ZN(n11442) );
  AND2_X1 U12904 ( .A1(n13388), .A2(n9817), .ZN(n10399) );
  AOI22_X1 U12905 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19224), .B1(
        n19284), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10592) );
  NAND2_X1 U12906 ( .A1(n10434), .A2(n10433), .ZN(n10436) );
  AOI22_X1 U12907 ( .A1(n9824), .A2(P2_EBX_REG_1__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n10429) );
  INV_X1 U12908 ( .A(n11424), .ZN(n11434) );
  INV_X1 U12909 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10990) );
  NOR2_X1 U12910 ( .A1(n11162), .A2(n11278), .ZN(n11219) );
  OR2_X1 U12911 ( .A1(n11336), .A2(n11335), .ZN(n11368) );
  AND2_X1 U12912 ( .A1(n13480), .A2(n11997), .ZN(n11109) );
  OR2_X1 U12913 ( .A1(n11205), .A2(n11204), .ZN(n11260) );
  OR2_X1 U12914 ( .A1(n10611), .A2(n10610), .ZN(n10655) );
  NOR2_X1 U12915 ( .A1(n9913), .A2(n10686), .ZN(n10687) );
  AND2_X1 U12916 ( .A1(n10407), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10411) );
  AND4_X1 U12917 ( .A1(n11051), .A2(n11050), .A3(n11049), .A4(n11048), .ZN(
        n11052) );
  AND2_X1 U12918 ( .A1(n11364), .A2(n11363), .ZN(n11366) );
  OR2_X1 U12919 ( .A1(n11309), .A2(n11308), .ZN(n11317) );
  INV_X1 U12920 ( .A(n11174), .ZN(n11175) );
  AND4_X1 U12921 ( .A1(n11010), .A2(n11009), .A3(n11008), .A4(n11007), .ZN(
        n11011) );
  NAND2_X1 U12922 ( .A1(n10439), .A2(n10418), .ZN(n10441) );
  AND2_X1 U12923 ( .A1(n19134), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10762) );
  INV_X1 U12924 ( .A(n13057), .ZN(n13058) );
  NOR2_X1 U12925 ( .A1(n14270), .A2(n14269), .ZN(n14272) );
  INV_X1 U12926 ( .A(n13895), .ZN(n10932) );
  NAND2_X1 U12927 ( .A1(n10689), .A2(n10688), .ZN(n10705) );
  OR2_X1 U12928 ( .A1(n11747), .A2(n11748), .ZN(n11743) );
  AND2_X1 U12929 ( .A1(n17649), .A2(n17757), .ZN(n11896) );
  AND2_X1 U12930 ( .A1(n11460), .A2(n11459), .ZN(n11480) );
  AND2_X1 U12931 ( .A1(n14312), .A2(n12452), .ZN(n12453) );
  INV_X1 U12932 ( .A(n14352), .ZN(n12409) );
  AND2_X1 U12933 ( .A1(n12170), .A2(n14140), .ZN(n12171) );
  INV_X1 U12934 ( .A(n11999), .ZN(n12424) );
  AND2_X1 U12935 ( .A1(n11414), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11415) );
  AND2_X1 U12936 ( .A1(n11510), .A2(n11509), .ZN(n13712) );
  AOI221_X1 U12937 ( .B1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n11450), 
        .C1(n13690), .C2(n11450), .A(n11422), .ZN(n11479) );
  NAND2_X1 U12938 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n19823), .ZN(
        n10836) );
  NAND2_X1 U12939 ( .A1(n10788), .A2(n15007), .ZN(n10802) );
  INV_X1 U12940 ( .A(n10657), .ZN(n10658) );
  NAND2_X1 U12941 ( .A1(n10248), .A2(n13058), .ZN(n13059) );
  AND2_X1 U12942 ( .A1(n12634), .A2(n12633), .ZN(n13592) );
  INV_X1 U12943 ( .A(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n16248) );
  INV_X1 U12944 ( .A(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n20918) );
  NOR2_X1 U12945 ( .A1(n18134), .A2(n18112), .ZN(n11917) );
  INV_X1 U12946 ( .A(n12340), .ZN(n12341) );
  AND2_X1 U12947 ( .A1(n11543), .A2(n11542), .ZN(n14185) );
  AND2_X1 U12948 ( .A1(n15754), .A2(n12452), .ZN(n12364) );
  NAND2_X1 U12949 ( .A1(n12490), .A2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12491) );
  INV_X1 U12950 ( .A(n12168), .ZN(n12130) );
  INV_X1 U12951 ( .A(n20793), .ZN(n11391) );
  INV_X1 U12952 ( .A(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13661) );
  INV_X1 U12953 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20514) );
  NOR2_X1 U12954 ( .A1(n13746), .A2(n13745), .ZN(n12891) );
  INV_X1 U12955 ( .A(n13111), .ZN(n13112) );
  AND2_X1 U12956 ( .A1(n14998), .A2(n13027), .ZN(n13002) );
  INV_X1 U12957 ( .A(n13793), .ZN(n12892) );
  INV_X1 U12958 ( .A(n14873), .ZN(n14874) );
  NAND2_X1 U12959 ( .A1(n13967), .A2(n13966), .ZN(n13965) );
  NOR2_X1 U12960 ( .A1(n19838), .A2(n13334), .ZN(n10843) );
  INV_X1 U12961 ( .A(n13718), .ZN(n12680) );
  OAI22_X1 U12962 ( .A1(n18720), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B1(
        n20944), .B2(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n11930) );
  NOR2_X1 U12963 ( .A1(n11895), .A2(n17604), .ZN(n17418) );
  NAND2_X1 U12964 ( .A1(n17434), .A2(n17471), .ZN(n17472) );
  OAI21_X1 U12965 ( .B1(n11917), .B2(n11916), .A(n11915), .ZN(n18543) );
  INV_X1 U12966 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n11869) );
  NAND2_X1 U12967 ( .A1(n18128), .A2(n18117), .ZN(n11730) );
  AND2_X1 U12968 ( .A1(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n12341), .ZN(
        n12342) );
  NOR2_X1 U12969 ( .A1(n14257), .A2(n16000), .ZN(n12492) );
  AND2_X1 U12970 ( .A1(n14257), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14198) );
  AND2_X1 U12971 ( .A1(n11545), .A2(n11544), .ZN(n14180) );
  OR2_X1 U12972 ( .A1(n14338), .A2(n14300), .ZN(n14301) );
  AND2_X1 U12973 ( .A1(n13482), .A2(n13481), .ZN(n13483) );
  NAND2_X1 U12974 ( .A1(n12429), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12456) );
  OR2_X1 U12975 ( .A1(n12389), .A2(n12388), .ZN(n14360) );
  INV_X1 U12976 ( .A(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n12187) );
  AND2_X1 U12977 ( .A1(n12130), .A2(n12105), .ZN(n14131) );
  INV_X1 U12978 ( .A(n12521), .ZN(n12523) );
  AND2_X1 U12979 ( .A1(n20099), .A2(n11616), .ZN(n14790) );
  INV_X1 U12980 ( .A(n20089), .ZN(n15975) );
  NAND2_X2 U12981 ( .A1(n20153), .A2(n11233), .ZN(n20380) );
  INV_X1 U12982 ( .A(n9828), .ZN(n20105) );
  NOR2_X1 U12983 ( .A1(n20262), .A2(n20513), .ZN(n20447) );
  NOR2_X1 U12984 ( .A1(n20262), .A2(n20438), .ZN(n20589) );
  AND2_X1 U12985 ( .A1(n13700), .A2(n20105), .ZN(n20486) );
  NAND3_X1 U12986 ( .A1(n10427), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n13334), 
        .ZN(n13584) );
  AND2_X1 U12987 ( .A1(n12926), .A2(n13811), .ZN(n13997) );
  AOI21_X1 U12988 ( .B1(n16013), .B2(n19104), .A(n14290), .ZN(n14291) );
  NOR2_X1 U12989 ( .A1(n14241), .A2(n14240), .ZN(n14242) );
  AND2_X1 U12990 ( .A1(n15181), .A2(n15180), .ZN(n15231) );
  INV_X1 U12991 ( .A(n19253), .ZN(n19318) );
  OR2_X1 U12992 ( .A1(n19804), .A2(n19808), .ZN(n19468) );
  NAND3_X1 U12993 ( .A1(n19612), .A2(P2_STATEBS16_REG_SCAN_IN), .A3(n19648), 
        .ZN(n13941) );
  INV_X1 U12994 ( .A(n19612), .ZN(n19790) );
  INV_X1 U12995 ( .A(n19152), .ZN(n19144) );
  AND3_X1 U12996 ( .A1(n13616), .A2(n13615), .A3(n13614), .ZN(n16268) );
  NOR2_X1 U12997 ( .A1(n18100), .A2(n18746), .ZN(n11910) );
  NOR2_X1 U12998 ( .A1(n11766), .A2(n11765), .ZN(n11767) );
  NOR2_X1 U12999 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16605), .ZN(n16596) );
  NOR2_X1 U13000 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16631), .ZN(n16619) );
  NOR2_X1 U13001 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n16721), .ZN(n16706) );
  NOR2_X1 U13002 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(n16747), .ZN(n16730) );
  NAND2_X1 U13003 ( .A1(n11753), .A2(n18746), .ZN(n11760) );
  INV_X1 U13004 ( .A(n17452), .ZN(n17483) );
  NAND2_X1 U13005 ( .A1(n17840), .A2(n17376), .ZN(n11976) );
  AND2_X1 U13006 ( .A1(n15673), .A2(n18062), .ZN(n11943) );
  NAND2_X1 U13007 ( .A1(n11891), .A2(n10305), .ZN(n11892) );
  NOR2_X1 U13008 ( .A1(n18549), .A2(n18566), .ZN(n17858) );
  AOI21_X2 U13009 ( .B1(n18544), .B2(n18552), .A(n18543), .ZN(n18554) );
  NOR2_X1 U13010 ( .A1(n18549), .A2(n18540), .ZN(n17967) );
  INV_X1 U13011 ( .A(n17996), .ZN(n17653) );
  NOR2_X1 U13012 ( .A1(n17692), .A2(n17691), .ZN(n17690) );
  INV_X1 U13013 ( .A(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20944) );
  INV_X1 U13014 ( .A(n11900), .ZN(n18106) );
  AOI22_X1 U13015 ( .A1(n18052), .A2(n18535), .B1(n18532), .B2(n16296), .ZN(
        n16297) );
  OR2_X1 U13016 ( .A1(n13263), .A2(n19857), .ZN(n13261) );
  OAI21_X1 U13017 ( .B1(n14447), .B2(n19937), .A(n12517), .ZN(n12518) );
  NAND2_X1 U13018 ( .A1(n12257), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n12290) );
  NOR2_X1 U13019 ( .A1(n14196), .A2(n19890), .ZN(n15849) );
  NOR2_X1 U13020 ( .A1(n19891), .A2(n19911), .ZN(n19898) );
  AND2_X1 U13021 ( .A1(n14430), .A2(n14198), .ZN(n19941) );
  AND2_X1 U13022 ( .A1(n11532), .A2(n11531), .ZN(n14056) );
  INV_X1 U13023 ( .A(n14529), .ZN(n14558) );
  INV_X1 U13024 ( .A(n20016), .ZN(n13555) );
  NAND2_X1 U13025 ( .A1(n12291), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12340) );
  AND2_X1 U13026 ( .A1(n14149), .A2(n14143), .ZN(n15881) );
  NOR2_X1 U13027 ( .A1(n12025), .A2(n15916), .ZN(n12029) );
  AND2_X1 U13028 ( .A1(n20581), .A2(n13620), .ZN(n20101) );
  AND2_X1 U13029 ( .A1(n14750), .A2(n10205), .ZN(n15922) );
  AND2_X1 U13030 ( .A1(n15930), .A2(n11615), .ZN(n14750) );
  INV_X1 U13031 ( .A(n14790), .ZN(n20076) );
  NOR2_X1 U13032 ( .A1(n20064), .A2(n14819), .ZN(n20057) );
  NOR2_X1 U13033 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n14858) );
  INV_X1 U13034 ( .A(n20169), .ZN(n20176) );
  OAI22_X1 U13035 ( .A1(n20187), .A2(n20186), .B1(n20383), .B2(n20316), .ZN(
        n20211) );
  NAND2_X1 U13036 ( .A1(n20103), .A2(n20378), .ZN(n20221) );
  OAI221_X1 U13037 ( .B1(n20279), .B2(n20388), .C1(n20279), .C2(n20263), .A(
        n20589), .ZN(n20282) );
  OR2_X1 U13038 ( .A1(n13700), .A2(n9828), .ZN(n20413) );
  INV_X1 U13039 ( .A(n20486), .ZN(n20348) );
  OAI211_X1 U13040 ( .C1(n20403), .C2(n20388), .A(n20447), .B(n20387), .ZN(
        n20406) );
  INV_X1 U13041 ( .A(n20379), .ZN(n20508) );
  AND2_X1 U13042 ( .A1(n20487), .A2(n20549), .ZN(n20475) );
  AND2_X1 U13043 ( .A1(n20766), .A2(n20378), .ZN(n20487) );
  AND2_X1 U13044 ( .A1(n20487), .A2(n20486), .ZN(n20543) );
  AND2_X1 U13045 ( .A1(n20580), .A2(n20508), .ZN(n20575) );
  INV_X1 U13046 ( .A(n20591), .ZN(n20623) );
  INV_X1 U13047 ( .A(n20450), .ZN(n20643) );
  INV_X1 U13048 ( .A(n20462), .ZN(n20661) );
  AND2_X1 U13049 ( .A1(n20580), .A2(n20486), .ZN(n20683) );
  INV_X1 U13050 ( .A(n18947), .ZN(n18933) );
  INV_X1 U13051 ( .A(n18954), .ZN(n18885) );
  INV_X1 U13052 ( .A(n18937), .ZN(n18949) );
  INV_X1 U13053 ( .A(n15254), .ZN(n18847) );
  OR2_X1 U13054 ( .A1(n12775), .A2(n12774), .ZN(n13811) );
  INV_X1 U13055 ( .A(n12890), .ZN(n13746) );
  OR2_X1 U13056 ( .A1(n13507), .A2(n13508), .ZN(n13583) );
  INV_X1 U13057 ( .A(n19013), .ZN(n18989) );
  INV_X1 U13058 ( .A(n13429), .ZN(n19082) );
  AND2_X1 U13059 ( .A1(n13798), .A2(n13797), .ZN(n18889) );
  AND2_X1 U13060 ( .A1(n19113), .A2(n13369), .ZN(n19101) );
  INV_X1 U13061 ( .A(n19113), .ZN(n19086) );
  AND2_X1 U13062 ( .A1(n15488), .A2(n12852), .ZN(n16197) );
  INV_X1 U13063 ( .A(n16222), .ZN(n16209) );
  INV_X1 U13064 ( .A(n16217), .ZN(n16227) );
  XNOR2_X1 U13065 ( .A(n13503), .B(n13502), .ZN(n19804) );
  NAND2_X1 U13066 ( .A1(n16257), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n16286) );
  OAI21_X1 U13067 ( .B1(n13947), .B2(n13946), .A(n13945), .ZN(n19153) );
  AND2_X1 U13068 ( .A1(n19788), .A2(n19818), .ZN(n19253) );
  AND2_X1 U13069 ( .A1(n19253), .A2(n19784), .ZN(n19238) );
  OAI21_X1 U13070 ( .B1(n19257), .B2(n19273), .A(n19256), .ZN(n19275) );
  NOR2_X1 U13071 ( .A1(n19318), .A2(n19555), .ZN(n19303) );
  NOR2_X1 U13072 ( .A1(n19347), .A2(n19789), .ZN(n19395) );
  NAND2_X1 U13073 ( .A1(n19407), .A2(n19818), .ZN(n19607) );
  INV_X1 U13074 ( .A(n19467), .ZN(n19457) );
  NOR2_X1 U13075 ( .A1(n19607), .A2(n19468), .ZN(n19499) );
  OR3_X1 U13076 ( .A1(n19520), .A2(n19519), .A3(n19613), .ZN(n19538) );
  NAND2_X1 U13077 ( .A1(n19804), .A2(n19808), .ZN(n19555) );
  INV_X1 U13078 ( .A(n19608), .ZN(n19641) );
  INV_X1 U13079 ( .A(n19484), .ZN(n19658) );
  INV_X1 U13080 ( .A(n19363), .ZN(n19674) );
  NAND2_X1 U13081 ( .A1(n19804), .A2(n19786), .ZN(n19789) );
  INV_X1 U13082 ( .A(n11753), .ZN(n18759) );
  NOR2_X1 U13083 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16541), .ZN(n16526) );
  NOR2_X1 U13084 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16561), .ZN(n16548) );
  NOR2_X1 U13085 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16579), .ZN(n16570) );
  NOR2_X1 U13086 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n16653), .ZN(n16636) );
  NOR2_X1 U13087 ( .A1(P3_EBX_REG_12__SCAN_IN), .A2(n16678), .ZN(n16658) );
  NOR2_X1 U13088 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n16699), .ZN(n16683) );
  NOR2_X1 U13089 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(n16775), .ZN(n16751) );
  NAND4_X1 U13090 ( .A1(n18074), .A2(n18759), .A3(n18602), .A4(n18593), .ZN(
        n16810) );
  INV_X1 U13091 ( .A(n16960), .ZN(n16937) );
  INV_X1 U13092 ( .A(P3_EBX_REG_3__SCAN_IN), .ZN(n17091) );
  NOR3_X1 U13093 ( .A1(n17153), .A2(n17316), .A3(n17187), .ZN(n17179) );
  INV_X1 U13094 ( .A(n17161), .ZN(n17185) );
  INV_X1 U13095 ( .A(n17257), .ZN(n17245) );
  INV_X1 U13096 ( .A(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n21050) );
  NOR2_X2 U13097 ( .A1(n18394), .A2(n18444), .ZN(n18476) );
  NOR2_X2 U13098 ( .A1(n17754), .A2(n16315), .ZN(n17655) );
  INV_X1 U13099 ( .A(n17754), .ZN(n17738) );
  NAND2_X1 U13100 ( .A1(n11977), .A2(n11976), .ZN(n11978) );
  INV_X1 U13101 ( .A(n17858), .ZN(n18045) );
  NAND2_X1 U13102 ( .A1(n17557), .A2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n17556) );
  INV_X1 U13103 ( .A(n17909), .ZN(n17994) );
  INV_X1 U13104 ( .A(n18079), .ZN(n18037) );
  INV_X1 U13105 ( .A(n17867), .ZN(n18035) );
  INV_X1 U13106 ( .A(n18077), .ZN(n18066) );
  NAND2_X1 U13107 ( .A1(n18604), .A2(n18092), .ZN(n18394) );
  NOR2_X1 U13108 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18696), .ZN(
        n18721) );
  CLKBUF_X1 U13109 ( .A(n18196), .Z(n18206) );
  INV_X1 U13110 ( .A(n16297), .ZN(n18586) );
  INV_X1 U13111 ( .A(P3_STATE_REG_1__SCAN_IN), .ZN(n20880) );
  INV_X1 U13112 ( .A(n14173), .ZN(n20102) );
  AND2_X1 U13113 ( .A1(n13284), .A2(n13261), .ZN(n20789) );
  INV_X1 U13114 ( .A(n12518), .ZN(n12519) );
  INV_X1 U13115 ( .A(n19932), .ZN(n19954) );
  INV_X1 U13116 ( .A(n19951), .ZN(n19937) );
  AND2_X1 U13117 ( .A1(n15796), .A2(n14428), .ZN(n19960) );
  NAND2_X1 U13118 ( .A1(n19968), .A2(n14503), .ZN(n19962) );
  AND2_X2 U13119 ( .A1(n13521), .A2(n13520), .ZN(n19968) );
  OAI21_X1 U13120 ( .B1(n10306), .B2(n14470), .A(n14471), .ZN(n15772) );
  INV_X1 U13121 ( .A(n14649), .ZN(n14567) );
  INV_X1 U13122 ( .A(n19969), .ZN(n19995) );
  NOR2_X1 U13123 ( .A1(n13284), .A2(n13283), .ZN(n13416) );
  INV_X1 U13124 ( .A(n15911), .ZN(n15909) );
  INV_X1 U13125 ( .A(n20043), .ZN(n19863) );
  OR2_X1 U13126 ( .A1(n13622), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20046) );
  NAND2_X1 U13127 ( .A1(n11613), .A2(n11498), .ZN(n20095) );
  INV_X1 U13128 ( .A(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n20551) );
  OR2_X1 U13129 ( .A1(n20221), .A2(n20379), .ZN(n20169) );
  OR2_X1 U13130 ( .A1(n20221), .A2(n20413), .ZN(n20209) );
  INV_X1 U13131 ( .A(n20220), .ZN(n20255) );
  OR2_X1 U13132 ( .A1(n20221), .A2(n20348), .ZN(n20278) );
  OR2_X1 U13133 ( .A1(n20351), .A2(n20379), .ZN(n20304) );
  OR2_X1 U13134 ( .A1(n20351), .A2(n20413), .ZN(n20342) );
  OR2_X1 U13135 ( .A1(n20351), .A2(n20348), .ZN(n20371) );
  NAND2_X1 U13136 ( .A1(n20487), .A2(n20508), .ZN(n20433) );
  AOI22_X1 U13137 ( .A1(n20445), .A2(n20443), .B1(n20439), .B2(n20438), .ZN(
        n20479) );
  NAND2_X1 U13138 ( .A1(n20487), .A2(n20579), .ZN(n20507) );
  AOI22_X1 U13139 ( .A1(n20518), .A2(n20515), .B1(n20520), .B2(n20513), .ZN(
        n20548) );
  NAND2_X1 U13140 ( .A1(n20580), .A2(n20549), .ZN(n20591) );
  NAND2_X1 U13141 ( .A1(n20580), .A2(n20579), .ZN(n20687) );
  INV_X1 U13142 ( .A(n20756), .ZN(n20693) );
  OR2_X1 U13143 ( .A1(n16255), .A2(n13241), .ZN(n13289) );
  AND2_X1 U13144 ( .A1(n13381), .A2(n13386), .ZN(n19847) );
  NAND2_X1 U13145 ( .A1(n19081), .A2(n16280), .ZN(n18945) );
  NAND2_X1 U13146 ( .A1(n13583), .A2(n13509), .ZN(n19788) );
  NAND2_X1 U13147 ( .A1(n15083), .A2(n10420), .ZN(n19009) );
  OR2_X1 U13148 ( .A1(n19057), .A2(n19850), .ZN(n19059) );
  INV_X1 U13149 ( .A(n19057), .ZN(n19078) );
  OR2_X1 U13150 ( .A1(n13289), .A2(n13334), .ZN(n13452) );
  INV_X1 U13151 ( .A(P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16157) );
  INV_X1 U13152 ( .A(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n16191) );
  OR2_X1 U13153 ( .A1(n12663), .A2(n19825), .ZN(n16217) );
  OR2_X1 U13154 ( .A1(n12663), .A2(n19826), .ZN(n16223) );
  INV_X1 U13155 ( .A(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20934) );
  AOI211_X2 U13156 ( .C1(n13940), .C2(n13946), .A(n13939), .B(n19613), .ZN(
        n19157) );
  INV_X1 U13157 ( .A(n19207), .ZN(n19217) );
  INV_X1 U13158 ( .A(n19238), .ZN(n19248) );
  INV_X1 U13159 ( .A(n19268), .ZN(n19278) );
  AND2_X1 U13160 ( .A1(n19283), .A2(n19282), .ZN(n19307) );
  INV_X1 U13161 ( .A(n19372), .ZN(n19370) );
  INV_X1 U13162 ( .A(n19395), .ZN(n19405) );
  OR2_X1 U13163 ( .A1(n19607), .A2(n19408), .ZN(n19430) );
  OR2_X1 U13164 ( .A1(n19556), .A2(n19408), .ZN(n19467) );
  INV_X1 U13165 ( .A(n19499), .ZN(n19511) );
  INV_X1 U13166 ( .A(n19531), .ZN(n19541) );
  OR2_X1 U13167 ( .A1(n19556), .A2(n19555), .ZN(n19608) );
  AOI211_X2 U13168 ( .C1(n19616), .C2(n19619), .A(n19614), .B(n19613), .ZN(
        n19646) );
  AND3_X1 U13169 ( .A1(n16274), .A2(n16273), .A3(n16272), .ZN(n16293) );
  INV_X1 U13170 ( .A(n19783), .ZN(n19716) );
  INV_X1 U13171 ( .A(P3_STATEBS16_REG_SCAN_IN), .ZN(n18745) );
  INV_X1 U13172 ( .A(n16812), .ZN(n16801) );
  INV_X1 U13173 ( .A(n16754), .ZN(n16798) );
  NOR2_X1 U13174 ( .A1(n16542), .A2(n16877), .ZN(n16883) );
  AND2_X1 U13175 ( .A1(P3_EBX_REG_18__SCAN_IN), .A2(n16937), .ZN(n16949) );
  NOR2_X1 U13176 ( .A1(n11791), .A2(n11790), .ZN(n17233) );
  NAND2_X1 U13177 ( .A1(n18567), .A2(n17111), .ZN(n17257) );
  NAND2_X1 U13178 ( .A1(n17311), .A2(n17259), .ZN(n17309) );
  INV_X1 U13179 ( .A(n17362), .ZN(n17352) );
  INV_X1 U13180 ( .A(n17350), .ZN(n17364) );
  NAND2_X1 U13181 ( .A1(n16315), .A2(n17738), .ZN(n17652) );
  INV_X1 U13182 ( .A(n17655), .ZN(n17555) );
  INV_X1 U13183 ( .A(n17741), .ZN(n17736) );
  NOR2_X1 U13184 ( .A1(n17708), .A2(n17721), .ZN(n17746) );
  NAND2_X1 U13185 ( .A1(n11904), .A2(n18066), .ZN(n17909) );
  INV_X1 U13186 ( .A(n18055), .ZN(n18062) );
  OAI21_X2 U13187 ( .B1(n14223), .B2(n11942), .A(n18741), .ZN(n18061) );
  INV_X1 U13188 ( .A(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18088) );
  INV_X1 U13189 ( .A(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n18580) );
  INV_X1 U13190 ( .A(n18139), .ZN(n18480) );
  INV_X1 U13191 ( .A(n18155), .ZN(n18510) );
  OAI21_X1 U13192 ( .B1(n14248), .B2(n19108), .A(n10989), .ZN(P2_U2985) );
  AOI22_X1 U13193 ( .A1(n10538), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n10319) );
  AND2_X4 U13194 ( .A1(n15532), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n10540) );
  AOI22_X1 U13195 ( .A1(n10539), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10540), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10318) );
  AOI22_X1 U13196 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10353), .B2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n10317) );
  AND2_X4 U13197 ( .A1(n13594), .A2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13601) );
  AOI22_X1 U13198 ( .A1(n13601), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n9808), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10316) );
  NAND4_X1 U13199 ( .A1(n10319), .A2(n10318), .A3(n10317), .A4(n10316), .ZN(
        n10320) );
  AOI22_X1 U13200 ( .A1(n10538), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9827), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n10324) );
  AOI22_X1 U13201 ( .A1(n10539), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9833), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10323) );
  AOI22_X1 U13202 ( .A1(n13601), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9826), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10321) );
  NAND4_X1 U13203 ( .A1(n10324), .A2(n10323), .A3(n10322), .A4(n10321), .ZN(
        n10325) );
  AOI22_X1 U13204 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n9825), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10329) );
  AOI22_X1 U13205 ( .A1(n10539), .A2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9827), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n10328) );
  AOI22_X1 U13206 ( .A1(n13601), .A2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n9826), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10327) );
  AOI22_X1 U13207 ( .A1(n10538), .A2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n10540), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10326) );
  NAND4_X1 U13208 ( .A1(n10329), .A2(n10328), .A3(n10327), .A4(n10326), .ZN(
        n10330) );
  AOI22_X1 U13209 ( .A1(n10538), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10334) );
  AOI22_X1 U13210 ( .A1(n13601), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9808), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10333) );
  AOI22_X1 U13211 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n10353), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n10332) );
  AOI22_X1 U13212 ( .A1(n10539), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n9833), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10331) );
  NAND4_X1 U13213 ( .A1(n10334), .A2(n10333), .A3(n10332), .A4(n10331), .ZN(
        n10335) );
  INV_X1 U13214 ( .A(n12562), .ZN(n10361) );
  AOI22_X1 U13215 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n10353), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10339) );
  AOI22_X1 U13216 ( .A1(n10539), .A2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n10540), .B2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n10338) );
  AOI22_X1 U13217 ( .A1(n10538), .A2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n9827), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n10337) );
  AOI22_X1 U13218 ( .A1(n13601), .A2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9826), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10336) );
  NAND4_X1 U13219 ( .A1(n10339), .A2(n10338), .A3(n10337), .A4(n10336), .ZN(
        n10340) );
  NAND2_X1 U13220 ( .A1(n10340), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10347) );
  AOI22_X1 U13221 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(n9825), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n10344) );
  AOI22_X1 U13222 ( .A1(n10538), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n10343) );
  AOI22_X1 U13223 ( .A1(n10539), .A2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9833), .B2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n10342) );
  AOI22_X1 U13224 ( .A1(n13601), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9808), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10341) );
  NAND4_X1 U13225 ( .A1(n10344), .A2(n10343), .A3(n10342), .A4(n10341), .ZN(
        n10345) );
  NAND2_X1 U13226 ( .A1(n10345), .A2(n16232), .ZN(n10346) );
  NAND2_X1 U13227 ( .A1(n10347), .A2(n10346), .ZN(n10419) );
  INV_X1 U13228 ( .A(n10419), .ZN(n19129) );
  AOI22_X1 U13229 ( .A1(n10538), .A2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n10351) );
  AOI22_X1 U13230 ( .A1(n13601), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n9808), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10350) );
  AOI22_X1 U13231 ( .A1(n10539), .A2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n9833), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10349) );
  AOI22_X1 U13232 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(n9825), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n10348) );
  NAND4_X1 U13233 ( .A1(n10351), .A2(n10350), .A3(n10349), .A4(n10348), .ZN(
        n10352) );
  NAND2_X1 U13234 ( .A1(n10352), .A2(n16232), .ZN(n10360) );
  AOI22_X1 U13235 ( .A1(n10538), .A2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9827), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n10357) );
  AOI22_X1 U13236 ( .A1(n10539), .A2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n10540), .B2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n10356) );
  AOI22_X1 U13237 ( .A1(n13601), .A2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9826), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10355) );
  AOI22_X1 U13238 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n10353), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10354) );
  NAND4_X1 U13239 ( .A1(n10357), .A2(n10356), .A3(n10355), .A4(n10354), .ZN(
        n10358) );
  NAND2_X1 U13240 ( .A1(n10358), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10359) );
  INV_X1 U13241 ( .A(n12595), .ZN(n10426) );
  NAND2_X1 U13242 ( .A1(n10361), .A2(n10426), .ZN(n13384) );
  INV_X1 U13243 ( .A(n13384), .ZN(n10400) );
  AOI22_X1 U13244 ( .A1(n10538), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n10363) );
  AOI22_X1 U13245 ( .A1(n13601), .A2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9826), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10362) );
  AOI22_X1 U13246 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n9825), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10365) );
  AOI22_X1 U13247 ( .A1(n10539), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n9833), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10364) );
  INV_X1 U13248 ( .A(n10367), .ZN(n10368) );
  AOI22_X1 U13249 ( .A1(n10538), .A2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n10371) );
  AOI22_X1 U13250 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9825), .B2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n10370) );
  AOI22_X1 U13251 ( .A1(n10539), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9833), .B2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n10369) );
  AOI22_X1 U13252 ( .A1(n10538), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9827), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n10378) );
  AOI22_X1 U13253 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9825), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n10377) );
  AOI22_X1 U13254 ( .A1(n10539), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n10540), .B2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n10376) );
  AOI22_X1 U13255 ( .A1(n13601), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n10541), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n10375) );
  NAND4_X1 U13256 ( .A1(n10378), .A2(n10377), .A3(n10376), .A4(n10375), .ZN(
        n10379) );
  NAND2_X1 U13257 ( .A1(n10379), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10386) );
  AOI22_X1 U13258 ( .A1(n10538), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n10383) );
  AOI22_X1 U13259 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10539), .B1(
        n9833), .B2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n10382) );
  AOI22_X1 U13260 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n9834), .B1(
        n10353), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n10381) );
  AOI22_X1 U13261 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n13601), .B1(
        n10541), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n10380) );
  NAND4_X1 U13262 ( .A1(n10383), .A2(n10382), .A3(n10381), .A4(n10380), .ZN(
        n10384) );
  NAND2_X1 U13263 ( .A1(n10384), .A2(n16232), .ZN(n10385) );
  AOI22_X1 U13264 ( .A1(n10538), .A2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n10388) );
  AOI22_X1 U13265 ( .A1(n10539), .A2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n9833), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10387) );
  AND2_X1 U13266 ( .A1(n10388), .A2(n10387), .ZN(n10391) );
  AOI22_X1 U13267 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10353), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10390) );
  AOI22_X1 U13268 ( .A1(n13601), .A2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n10541), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10389) );
  NAND3_X1 U13269 ( .A1(n10391), .A2(n10390), .A3(n10304), .ZN(n10398) );
  AOI22_X1 U13270 ( .A1(n10538), .A2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n9827), .B2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n10395) );
  AOI22_X1 U13271 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n10353), .B2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n10394) );
  AOI22_X1 U13272 ( .A1(n10539), .A2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n10540), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10393) );
  NAND2_X1 U13273 ( .A1(n10400), .A2(n10399), .ZN(n10417) );
  INV_X1 U13274 ( .A(n12644), .ZN(n10414) );
  AOI22_X1 U13275 ( .A1(n13601), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9808), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n10403) );
  AOI22_X1 U13276 ( .A1(n10539), .A2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n9833), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10402) );
  NAND2_X1 U13277 ( .A1(n10406), .A2(n16232), .ZN(n10413) );
  AOI22_X1 U13278 ( .A1(n13601), .A2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n9808), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10407) );
  AOI22_X1 U13279 ( .A1(n9837), .A2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n10540), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n10410) );
  AOI22_X1 U13280 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10353), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n10409) );
  AOI22_X1 U13281 ( .A1(n10538), .A2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10408) );
  NAND4_X1 U13282 ( .A1(n10411), .A2(n10410), .A3(n10409), .A4(n10408), .ZN(
        n10412) );
  NAND4_X1 U13283 ( .A1(n19129), .A2(n10414), .A3(n12645), .A4(n10443), .ZN(
        n10415) );
  NAND2_X1 U13284 ( .A1(n15659), .A2(n19838), .ZN(n12598) );
  NAND2_X1 U13285 ( .A1(n10417), .A2(n12598), .ZN(n10453) );
  NAND2_X1 U13286 ( .A1(n10428), .A2(n10427), .ZN(n12589) );
  INV_X1 U13287 ( .A(n12589), .ZN(n10418) );
  NAND2_X1 U13289 ( .A1(n10418), .A2(n19838), .ZN(n10422) );
  INV_X1 U13290 ( .A(P2_REIP_REG_1__SCAN_IN), .ZN(n10425) );
  NAND3_X1 U13291 ( .A1(n10431), .A2(n10430), .A3(n10429), .ZN(n10459) );
  INV_X1 U13292 ( .A(n10459), .ZN(n10458) );
  NAND2_X1 U13293 ( .A1(n10442), .A2(n12641), .ZN(n10435) );
  NAND3_X1 U13294 ( .A1(n9856), .A2(n10436), .A3(n10435), .ZN(n10438) );
  INV_X1 U13295 ( .A(n15659), .ZN(n10437) );
  INV_X1 U13296 ( .A(n12643), .ZN(n10452) );
  NAND2_X1 U13297 ( .A1(n10439), .A2(n10432), .ZN(n10842) );
  NAND2_X1 U13298 ( .A1(n10842), .A2(n10303), .ZN(n10440) );
  NAND2_X1 U13299 ( .A1(n12657), .A2(n19114), .ZN(n10451) );
  NAND3_X1 U13300 ( .A1(n12589), .A2(n12645), .A3(n12588), .ZN(n12596) );
  NAND3_X1 U13301 ( .A1(n12596), .A2(n12597), .A3(n10443), .ZN(n12639) );
  NAND2_X1 U13302 ( .A1(n12639), .A2(n12641), .ZN(n10445) );
  NAND2_X1 U13303 ( .A1(n19129), .A2(n12635), .ZN(n10444) );
  NAND3_X1 U13304 ( .A1(n10445), .A2(n10444), .A3(n19114), .ZN(n10449) );
  NAND2_X1 U13305 ( .A1(n12635), .A2(n10293), .ZN(n10448) );
  NAND2_X1 U13306 ( .A1(n10449), .A2(n10448), .ZN(n10450) );
  INV_X1 U13307 ( .A(n10453), .ZN(n10454) );
  NAND2_X1 U13308 ( .A1(n10454), .A2(n12660), .ZN(n12628) );
  NAND2_X1 U13309 ( .A1(n10983), .A2(n15527), .ZN(n19846) );
  NOR2_X1 U13310 ( .A1(n19846), .A2(n19814), .ZN(n10455) );
  NAND2_X1 U13311 ( .A1(n10458), .A2(n10457), .ZN(n10476) );
  NAND2_X1 U13312 ( .A1(n10460), .A2(n10459), .ZN(n10461) );
  NAND2_X1 U13313 ( .A1(n10477), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n10466) );
  NAND2_X1 U13314 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n10462) );
  NAND2_X1 U13315 ( .A1(n19846), .A2(n10462), .ZN(n10463) );
  AOI21_X1 U13316 ( .B1(n10468), .B2(P2_EBX_REG_0__SCAN_IN), .A(n10463), .ZN(
        n10465) );
  NAND2_X1 U13317 ( .A1(n9899), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n10464) );
  NAND2_X1 U13318 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_STATE2_REG_0__SCAN_IN), .ZN(n10469) );
  NAND2_X1 U13319 ( .A1(n10485), .A2(n10469), .ZN(n10470) );
  OAI21_X1 U13320 ( .B1(n10467), .B2(n10471), .A(n10470), .ZN(n10475) );
  INV_X1 U13321 ( .A(n10472), .ZN(n12629) );
  NOR2_X1 U13322 ( .A1(n19846), .A2(n19823), .ZN(n10473) );
  AOI21_X1 U13323 ( .B1(n12629), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n10473), 
        .ZN(n10474) );
  NAND2_X1 U13324 ( .A1(n10475), .A2(n10474), .ZN(n10495) );
  INV_X2 U13325 ( .A(n10477), .ZN(n12625) );
  INV_X1 U13326 ( .A(P2_REIP_REG_2__SCAN_IN), .ZN(n10480) );
  NAND2_X1 U13327 ( .A1(n10468), .A2(P2_EBX_REG_2__SCAN_IN), .ZN(n10479) );
  NAND2_X1 U13328 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n10478) );
  OAI211_X1 U13329 ( .C1(n10913), .C2(n10480), .A(n10479), .B(n10478), .ZN(
        n10481) );
  AOI21_X1 U13330 ( .B1(n10983), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n10483) );
  INV_X1 U13331 ( .A(n10497), .ZN(n10484) );
  OAI22_X1 U13332 ( .A1(n10482), .A2(n16232), .B1(n19846), .B2(n19796), .ZN(
        n10488) );
  INV_X1 U13333 ( .A(P2_REIP_REG_3__SCAN_IN), .ZN(n12690) );
  AOI22_X1 U13334 ( .A1(n10468), .A2(P2_EBX_REG_3__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10486) );
  NAND2_X1 U13335 ( .A1(n10488), .A2(n10487), .ZN(n10489) );
  INV_X1 U13336 ( .A(n10490), .ZN(n10491) );
  XNOR2_X1 U13337 ( .A(n10497), .B(n10496), .ZN(n10498) );
  XNOR2_X2 U13338 ( .A(n10499), .B(n10498), .ZN(n12868) );
  INV_X1 U13339 ( .A(n10500), .ZN(n10506) );
  INV_X1 U13340 ( .A(n10493), .ZN(n10501) );
  NAND2_X1 U13341 ( .A1(n10506), .A2(n10501), .ZN(n10502) );
  NAND2_X1 U13342 ( .A1(n12868), .A2(n15536), .ZN(n10524) );
  INV_X1 U13343 ( .A(n10503), .ZN(n10505) );
  NAND2_X1 U13344 ( .A1(n10505), .A2(n10504), .ZN(n10525) );
  NOR2_X2 U13345 ( .A1(n10511), .A2(n19105), .ZN(n19224) );
  AOI22_X1 U13346 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19321), .B1(
        n19224), .B2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n10518) );
  NAND2_X1 U13347 ( .A1(n10506), .A2(n18950), .ZN(n10512) );
  AOI22_X1 U13348 ( .A1(P2_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n19284), .B1(
        n19159), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n10517) );
  NOR2_X1 U13349 ( .A1(n12868), .A2(n10525), .ZN(n10508) );
  AND2_X1 U13350 ( .A1(n10521), .A2(n10508), .ZN(n19472) );
  INV_X1 U13351 ( .A(n10512), .ZN(n10509) );
  AND2_X1 U13352 ( .A1(n12868), .A2(n10509), .ZN(n10510) );
  AOI22_X1 U13353 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19472), .B1(
        n19543), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10516) );
  NOR2_X2 U13354 ( .A1(n10511), .A2(n14914), .ZN(n19348) );
  NOR2_X1 U13355 ( .A1(n12868), .A2(n10512), .ZN(n10513) );
  NAND2_X1 U13356 ( .A1(n10513), .A2(n10521), .ZN(n10514) );
  AOI22_X1 U13357 ( .A1(n19348), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_9__1__SCAN_IN), .B2(n19412), .ZN(n10515) );
  AND4_X1 U13358 ( .A1(n10518), .A2(n10517), .A3(n10516), .A4(n10515), .ZN(
        n10537) );
  AOI22_X1 U13359 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19250), .B1(
        n9879), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n10536) );
  INV_X1 U13360 ( .A(P2_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n13005) );
  INV_X1 U13361 ( .A(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n13015) );
  INV_X1 U13362 ( .A(n10522), .ZN(n10523) );
  OAI22_X1 U13363 ( .A1(n19190), .A2(n13005), .B1(n13015), .B2(n19442), .ZN(
        n10531) );
  INV_X1 U13364 ( .A(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10529) );
  INV_X1 U13365 ( .A(n10525), .ZN(n10526) );
  AND2_X1 U13366 ( .A1(n12868), .A2(n10526), .ZN(n10527) );
  OAI21_X1 U13367 ( .B1(n10581), .B2(n10529), .A(n10528), .ZN(n10530) );
  NOR2_X1 U13368 ( .A1(n10531), .A2(n10530), .ZN(n10535) );
  AOI22_X1 U13369 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19513), .B1(
        n19377), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10534) );
  NAND4_X1 U13370 ( .A1(n10537), .A2(n10536), .A3(n10535), .A4(n10534), .ZN(
        n10580) );
  AND2_X1 U13371 ( .A1(n10538), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10554) );
  AOI22_X1 U13372 ( .A1(n10554), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n10566), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n10545) );
  AND2_X2 U13373 ( .A1(n10401), .A2(n16232), .ZN(n10559) );
  AOI22_X1 U13374 ( .A1(n10559), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n10544) );
  AOI22_X1 U13375 ( .A1(n12952), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n10543) );
  AND2_X2 U13376 ( .A1(n9833), .A2(n16232), .ZN(n12954) );
  AND2_X1 U13377 ( .A1(n10541), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10567) );
  AOI22_X1 U13378 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10567), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n10542) );
  NAND4_X1 U13379 ( .A1(n10545), .A2(n10544), .A3(n10543), .A4(n10542), .ZN(
        n10553) );
  AOI22_X1 U13380 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n10551) );
  AND2_X2 U13381 ( .A1(n10401), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10695) );
  AND2_X1 U13382 ( .A1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n10547) );
  AOI22_X1 U13383 ( .A1(n10695), .A2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12975), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n10550) );
  AND2_X2 U13384 ( .A1(n13601), .A2(n16232), .ZN(n13593) );
  AND2_X1 U13385 ( .A1(n10541), .A2(n16232), .ZN(n10601) );
  AOI22_X1 U13386 ( .A1(n13593), .A2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n10549) );
  AOI22_X1 U13387 ( .A1(n10671), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n10548) );
  NAND4_X1 U13388 ( .A1(n10551), .A2(n10550), .A3(n10549), .A4(n10548), .ZN(
        n10552) );
  NOR2_X1 U13389 ( .A1(n10553), .A2(n10552), .ZN(n12671) );
  OR2_X1 U13390 ( .A1(n12671), .A2(n13334), .ZN(n10854) );
  INV_X1 U13391 ( .A(n10854), .ZN(n13340) );
  AOI22_X1 U13392 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10671), .B1(
        n10554), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n10558) );
  AOI22_X1 U13393 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n10557) );
  AOI22_X1 U13394 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n10601), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n10556) );
  AOI22_X1 U13395 ( .A1(P2_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n10567), .B1(
        n13593), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n10555) );
  NAND4_X1 U13396 ( .A1(n10558), .A2(n10557), .A3(n10556), .A4(n10555), .ZN(
        n10565) );
  AOI22_X1 U13397 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n10566), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n10563) );
  AOI22_X1 U13398 ( .A1(n10695), .A2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n12975), .ZN(n10562) );
  AOI22_X1 U13399 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10559), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n10561) );
  AOI22_X1 U13400 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n10560) );
  NAND4_X1 U13401 ( .A1(n10563), .A2(n10562), .A3(n10561), .A4(n10560), .ZN(
        n10564) );
  NAND2_X1 U13402 ( .A1(n13340), .A2(n10855), .ZN(n10858) );
  AOI22_X1 U13403 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n10566), .B1(
        n10554), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n10571) );
  AOI22_X1 U13404 ( .A1(n10671), .A2(P2_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n10567), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n10570) );
  AOI22_X1 U13405 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n10601), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n10569) );
  AOI22_X1 U13406 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n12725), .B1(
        n13593), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n10568) );
  NAND4_X1 U13407 ( .A1(n10571), .A2(n10570), .A3(n10569), .A4(n10568), .ZN(
        n10578) );
  AOI22_X1 U13408 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n10676), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n10576) );
  AOI22_X1 U13409 ( .A1(n10559), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__2__SCAN_IN), .B2(n12975), .ZN(n10575) );
  AOI22_X1 U13410 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n10695), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n10574) );
  AOI22_X1 U13411 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n10573) );
  NAND4_X1 U13412 ( .A1(n10576), .A2(n10575), .A3(n10574), .A4(n10573), .ZN(
        n10577) );
  NAND2_X1 U13413 ( .A1(n10858), .A2(n12683), .ZN(n10579) );
  INV_X1 U13414 ( .A(n10581), .ZN(n19617) );
  AOI22_X1 U13415 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19321), .B1(
        n19617), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10582) );
  INV_X1 U13416 ( .A(n10582), .ZN(n10591) );
  INV_X1 U13417 ( .A(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10584) );
  INV_X1 U13418 ( .A(n19472), .ZN(n10583) );
  INV_X1 U13419 ( .A(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n13072) );
  OAI22_X1 U13420 ( .A1(n10514), .A2(n10584), .B1(n10583), .B2(n13072), .ZN(
        n10585) );
  INV_X1 U13421 ( .A(n10585), .ZN(n10589) );
  NAND2_X1 U13422 ( .A1(n19543), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(
        n10586) );
  NAND2_X1 U13423 ( .A1(n10589), .A2(n10588), .ZN(n10590) );
  NOR2_X1 U13424 ( .A1(n10591), .A2(n10590), .ZN(n10600) );
  INV_X1 U13425 ( .A(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n19133) );
  NAND2_X1 U13426 ( .A1(n9879), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n10594) );
  AOI22_X1 U13427 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19348), .B1(
        n19159), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n10593) );
  INV_X1 U13428 ( .A(n19190), .ZN(n19186) );
  INV_X1 U13429 ( .A(n19442), .ZN(n19438) );
  AOI22_X1 U13430 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19186), .B1(
        n19438), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n10596) );
  NAND2_X1 U13431 ( .A1(n19513), .A2(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(
        n10595) );
  NAND4_X1 U13432 ( .A1(n10600), .A2(n10307), .A3(n10599), .A4(n10598), .ZN(
        n10613) );
  AOI22_X1 U13433 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n10676), .B1(
        n10554), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n10605) );
  AOI22_X1 U13434 ( .A1(n10671), .A2(P2_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n10604) );
  AOI22_X1 U13435 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n10690), .B1(
        n10567), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n10603) );
  AOI22_X1 U13436 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n12725), .B1(
        n13593), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n10602) );
  NAND4_X1 U13437 ( .A1(n10605), .A2(n10604), .A3(n10603), .A4(n10602), .ZN(
        n10611) );
  AOI22_X1 U13438 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n10566), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n10609) );
  AOI22_X1 U13439 ( .A1(n10559), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__3__SCAN_IN), .B2(n12975), .ZN(n10608) );
  AOI22_X1 U13440 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n10695), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n10607) );
  AOI22_X1 U13441 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n10606) );
  NAND4_X1 U13442 ( .A1(n10609), .A2(n10608), .A3(n10607), .A4(n10606), .ZN(
        n10610) );
  INV_X1 U13443 ( .A(n10655), .ZN(n12692) );
  NAND2_X1 U13444 ( .A1(n12692), .A2(n16281), .ZN(n10612) );
  NAND2_X1 U13445 ( .A1(n10615), .A2(n10614), .ZN(n10616) );
  NAND2_X1 U13446 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(
        n10620) );
  NAND2_X1 U13447 ( .A1(n10554), .A2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(
        n10619) );
  NAND2_X1 U13448 ( .A1(n10671), .A2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(
        n10618) );
  NAND2_X1 U13449 ( .A1(n10601), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(
        n10617) );
  NAND2_X1 U13450 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(
        n10624) );
  NAND2_X1 U13451 ( .A1(n10566), .A2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(
        n10623) );
  NAND2_X1 U13452 ( .A1(n12952), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(
        n10622) );
  NAND2_X1 U13453 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(
        n10621) );
  NAND2_X1 U13454 ( .A1(n10559), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(
        n10628) );
  NAND2_X1 U13455 ( .A1(n10695), .A2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(
        n10627) );
  NAND2_X1 U13456 ( .A1(n10572), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(
        n10626) );
  INV_X1 U13457 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n19156) );
  NAND2_X1 U13458 ( .A1(n12975), .A2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(
        n10625) );
  NAND2_X1 U13459 ( .A1(n10567), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(
        n10632) );
  NAND2_X1 U13460 ( .A1(n10690), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(
        n10631) );
  NAND2_X1 U13461 ( .A1(n13593), .A2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(
        n10630) );
  NAND2_X1 U13462 ( .A1(n12725), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(
        n10629) );
  XNOR2_X1 U13463 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n10846) );
  INV_X1 U13464 ( .A(n10836), .ZN(n10637) );
  NAND2_X1 U13465 ( .A1(n10846), .A2(n10637), .ZN(n10639) );
  NAND2_X1 U13466 ( .A1(n19814), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10638) );
  NAND2_X1 U13467 ( .A1(n10639), .A2(n10638), .ZN(n10645) );
  MUX2_X1 U13468 ( .A(n16248), .B(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .S(
        P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .Z(n10644) );
  XNOR2_X1 U13469 ( .A(n10645), .B(n10644), .ZN(n12569) );
  INV_X1 U13470 ( .A(n12569), .ZN(n10640) );
  MUX2_X1 U13471 ( .A(n10641), .B(n10640), .S(n9839), .Z(n10848) );
  INV_X1 U13472 ( .A(P2_EBX_REG_2__SCAN_IN), .ZN(n21020) );
  MUX2_X1 U13473 ( .A(n10848), .B(n21020), .S(n19134), .Z(n10668) );
  INV_X1 U13474 ( .A(P2_EBX_REG_0__SCAN_IN), .ZN(n13337) );
  AND2_X1 U13475 ( .A1(n19134), .A2(n13337), .ZN(n10662) );
  INV_X1 U13476 ( .A(P2_EBX_REG_1__SCAN_IN), .ZN(n14929) );
  NAND2_X1 U13477 ( .A1(n10662), .A2(n14929), .ZN(n10643) );
  NAND2_X1 U13478 ( .A1(n9983), .A2(n10855), .ZN(n10642) );
  NAND2_X1 U13479 ( .A1(n10643), .A2(n10642), .ZN(n10664) );
  NAND2_X1 U13480 ( .A1(n10668), .A2(n10664), .ZN(n10659) );
  NAND2_X1 U13481 ( .A1(n10645), .A2(n10644), .ZN(n10647) );
  NAND2_X1 U13482 ( .A1(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(n16248), .ZN(
        n10646) );
  NAND2_X1 U13483 ( .A1(n10647), .A2(n10646), .ZN(n10648) );
  INV_X1 U13484 ( .A(n10670), .ZN(n10653) );
  INV_X1 U13485 ( .A(n10648), .ZN(n10651) );
  INV_X1 U13486 ( .A(n10649), .ZN(n10650) );
  NAND2_X1 U13487 ( .A1(n10651), .A2(n10650), .ZN(n10652) );
  NAND2_X1 U13488 ( .A1(n10653), .A2(n10652), .ZN(n12572) );
  INV_X1 U13489 ( .A(n12572), .ZN(n10654) );
  MUX2_X1 U13490 ( .A(n10655), .B(n10654), .S(n9839), .Z(n10844) );
  INV_X1 U13491 ( .A(P2_EBX_REG_3__SCAN_IN), .ZN(n10656) );
  MUX2_X1 U13492 ( .A(n10844), .B(n10656), .S(n19134), .Z(n10657) );
  INV_X1 U13493 ( .A(n10688), .ZN(n10661) );
  NAND2_X1 U13494 ( .A1(n10659), .A2(n10658), .ZN(n10660) );
  NAND2_X1 U13495 ( .A1(n10661), .A2(n10660), .ZN(n14902) );
  OAI21_X1 U13496 ( .B1(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n19823), .A(
        n10836), .ZN(n12564) );
  MUX2_X1 U13497 ( .A(n12564), .B(n12671), .S(n12613), .Z(n10663) );
  AOI21_X1 U13498 ( .B1(n10663), .B2(n9983), .A(n10662), .ZN(n18943) );
  NAND2_X1 U13499 ( .A1(n18943), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13373) );
  INV_X1 U13500 ( .A(n10664), .ZN(n10667) );
  NAND3_X1 U13501 ( .A1(n19134), .A2(P2_EBX_REG_1__SCAN_IN), .A3(
        P2_EBX_REG_0__SCAN_IN), .ZN(n10665) );
  NAND2_X1 U13502 ( .A1(n10667), .A2(n10665), .ZN(n14930) );
  NOR2_X1 U13503 ( .A1(n13373), .A2(n14930), .ZN(n10666) );
  NAND2_X1 U13504 ( .A1(n13373), .A2(n14930), .ZN(n13372) );
  OAI21_X1 U13505 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n10666), .A(
        n13372), .ZN(n13403) );
  XNOR2_X1 U13506 ( .A(n10668), .B(n10667), .ZN(n14911) );
  XNOR2_X1 U13507 ( .A(n14911), .B(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n13402) );
  OR2_X1 U13508 ( .A1(n13403), .A2(n13402), .ZN(n13405) );
  NAND2_X1 U13509 ( .A1(n14911), .A2(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n10669) );
  NAND2_X1 U13510 ( .A1(n13405), .A2(n10669), .ZN(n14250) );
  NAND3_X1 U13511 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n10835), .A3(
        n15664), .ZN(n12560) );
  AOI22_X1 U13512 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10671), .B1(
        n10554), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n10675) );
  AOI22_X1 U13513 ( .A1(n10566), .A2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n10674) );
  AOI22_X1 U13514 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n12725), .B1(
        n13593), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n10673) );
  AOI22_X1 U13515 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n10601), .B1(
        n10567), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n10672) );
  NAND4_X1 U13516 ( .A1(n10675), .A2(n10674), .A3(n10673), .A4(n10672), .ZN(
        n10682) );
  AOI22_X1 U13517 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10676), .B1(
        n12954), .B2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n10680) );
  AOI22_X1 U13518 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__4__SCAN_IN), .B2(n12975), .ZN(n10679) );
  AOI22_X1 U13519 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10559), .B1(
        n10695), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n10678) );
  AOI22_X1 U13520 ( .A1(n12952), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n10677) );
  NAND4_X1 U13521 ( .A1(n10680), .A2(n10679), .A3(n10678), .A4(n10677), .ZN(
        n10681) );
  MUX2_X1 U13522 ( .A(n12560), .B(n12696), .S(n12613), .Z(n10845) );
  INV_X1 U13523 ( .A(P2_EBX_REG_4__SCAN_IN), .ZN(n14033) );
  MUX2_X1 U13524 ( .A(n10845), .B(n14033), .S(n19134), .Z(n10689) );
  XNOR2_X1 U13525 ( .A(n10689), .B(n10688), .ZN(n14038) );
  INV_X1 U13526 ( .A(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n13924) );
  NAND2_X1 U13527 ( .A1(n14038), .A2(n13924), .ZN(n10685) );
  OAI21_X1 U13528 ( .B1(n14250), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n10685), .ZN(n10683) );
  INV_X1 U13529 ( .A(n10683), .ZN(n10684) );
  NOR2_X1 U13530 ( .A1(n14038), .A2(n13924), .ZN(n10686) );
  AOI22_X1 U13531 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n10554), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n10694) );
  AOI22_X1 U13532 ( .A1(n10671), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n10693) );
  AOI22_X1 U13533 ( .A1(n10690), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10567), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n10692) );
  AOI22_X1 U13534 ( .A1(n13593), .A2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n10691) );
  NAND4_X1 U13535 ( .A1(n10694), .A2(n10693), .A3(n10692), .A4(n10691), .ZN(
        n10701) );
  AOI22_X1 U13536 ( .A1(n10566), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n10699) );
  INV_X1 U13537 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n19138) );
  AOI22_X1 U13538 ( .A1(n10559), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n12975), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n10698) );
  AOI22_X1 U13539 ( .A1(n10695), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n10697) );
  AOI22_X1 U13540 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n10696) );
  NAND4_X1 U13541 ( .A1(n10699), .A2(n10698), .A3(n10697), .A4(n10696), .ZN(
        n10700) );
  MUX2_X1 U13542 ( .A(n10868), .B(P2_EBX_REG_5__SCAN_IN), .S(n19134), .Z(
        n10704) );
  XNOR2_X1 U13543 ( .A(n10705), .B(n10704), .ZN(n10702) );
  INV_X1 U13544 ( .A(n10702), .ZN(n18932) );
  NAND2_X1 U13545 ( .A1(n18932), .A2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n10703) );
  AOI22_X1 U13546 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10671), .B1(
        n10554), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n10709) );
  AOI22_X1 U13547 ( .A1(n10566), .A2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n10708) );
  AOI22_X1 U13548 ( .A1(P2_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n10567), .B1(
        n13593), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n10707) );
  AOI22_X1 U13549 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n10601), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n10706) );
  NAND4_X1 U13550 ( .A1(n10709), .A2(n10708), .A3(n10707), .A4(n10706), .ZN(
        n10715) );
  AOI22_X1 U13551 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10676), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n10713) );
  AOI22_X1 U13552 ( .A1(n10559), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_0__6__SCAN_IN), .B2(n12975), .ZN(n10712) );
  AOI22_X1 U13553 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10695), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n10711) );
  AOI22_X1 U13554 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n10710) );
  NAND4_X1 U13555 ( .A1(n10713), .A2(n10712), .A3(n10711), .A4(n10710), .ZN(
        n10714) );
  INV_X1 U13556 ( .A(P2_EBX_REG_6__SCAN_IN), .ZN(n13645) );
  MUX2_X1 U13557 ( .A(n12706), .B(n13645), .S(n19134), .Z(n10717) );
  XNOR2_X1 U13558 ( .A(n10718), .B(n10717), .ZN(n10716) );
  XNOR2_X1 U13559 ( .A(n10716), .B(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n13983) );
  INV_X1 U13560 ( .A(n10716), .ZN(n18920) );
  INV_X1 U13561 ( .A(P2_EBX_REG_7__SCAN_IN), .ZN(n10719) );
  MUX2_X1 U13562 ( .A(n15187), .B(n10719), .S(n19134), .Z(n10722) );
  NAND2_X1 U13563 ( .A1(n19134), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10720) );
  NOR2_X1 U13564 ( .A1(n10733), .A2(n10720), .ZN(n10721) );
  NOR2_X1 U13565 ( .A1(n10730), .A2(n10721), .ZN(n14042) );
  NAND2_X1 U13566 ( .A1(n14042), .A2(n15187), .ZN(n10726) );
  INV_X1 U13567 ( .A(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n16207) );
  OR2_X1 U13568 ( .A1(n10726), .A2(n16207), .ZN(n16168) );
  INV_X1 U13569 ( .A(n10722), .ZN(n10723) );
  XNOR2_X1 U13570 ( .A(n10724), .B(n10723), .ZN(n18908) );
  NAND2_X1 U13571 ( .A1(n18908), .A2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n16164) );
  NAND2_X1 U13572 ( .A1(n16168), .A2(n16164), .ZN(n10725) );
  NAND2_X1 U13573 ( .A1(n10726), .A2(n16207), .ZN(n16167) );
  INV_X1 U13574 ( .A(n18908), .ZN(n10727) );
  INV_X1 U13575 ( .A(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n10882) );
  NAND2_X1 U13576 ( .A1(n10727), .A2(n10882), .ZN(n16166) );
  AND2_X1 U13577 ( .A1(n16167), .A2(n16166), .ZN(n10728) );
  INV_X1 U13578 ( .A(P2_EBX_REG_9__SCAN_IN), .ZN(n10729) );
  NAND2_X1 U13579 ( .A1(n19134), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n10731) );
  MUX2_X1 U13580 ( .A(n10731), .B(n19134), .S(n10730), .Z(n10732) );
  NAND2_X1 U13581 ( .A1(n10141), .A2(n10732), .ZN(n10738) );
  INV_X1 U13582 ( .A(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15497) );
  OAI21_X1 U13583 ( .B1(n10738), .B2(n15176), .A(n15497), .ZN(n14214) );
  INV_X1 U13584 ( .A(P2_EBX_REG_10__SCAN_IN), .ZN(n10741) );
  NOR2_X1 U13585 ( .A1(n10742), .A2(n10741), .ZN(n10734) );
  NAND2_X1 U13586 ( .A1(n19134), .A2(n10734), .ZN(n10735) );
  NAND2_X1 U13587 ( .A1(n12555), .A2(n10735), .ZN(n10736) );
  AOI21_X1 U13588 ( .B1(n10742), .B2(n10741), .A(n10736), .ZN(n18898) );
  AOI21_X1 U13589 ( .B1(n18898), .B2(n15187), .A(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15481) );
  AND2_X1 U13590 ( .A1(n15187), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10737) );
  INV_X1 U13591 ( .A(n10738), .ZN(n14893) );
  AND2_X1 U13592 ( .A1(n15187), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10739) );
  NAND2_X1 U13593 ( .A1(n14893), .A2(n10739), .ZN(n15479) );
  AND3_X1 U13594 ( .A1(n19134), .A2(P2_EBX_REG_11__SCAN_IN), .A3(n10743), .ZN(
        n10744) );
  OR2_X1 U13595 ( .A1(n10745), .A2(n10744), .ZN(n18883) );
  NOR2_X1 U13596 ( .A1(n18883), .A2(n15176), .ZN(n10766) );
  AND2_X1 U13597 ( .A1(n10766), .A2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n15467) );
  NAND2_X1 U13598 ( .A1(n19134), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10746) );
  NAND2_X1 U13599 ( .A1(n10143), .A2(n9884), .ZN(n10747) );
  NAND2_X1 U13600 ( .A1(n10764), .A2(n10747), .ZN(n18872) );
  INV_X1 U13601 ( .A(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15461) );
  XNOR2_X1 U13602 ( .A(n10768), .B(n15461), .ZN(n15168) );
  NAND2_X1 U13603 ( .A1(n19134), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10749) );
  OAI21_X1 U13604 ( .B1(P2_EBX_REG_15__SCAN_IN), .B2(P2_EBX_REG_14__SCAN_IN), 
        .A(n19134), .ZN(n10748) );
  NAND2_X1 U13605 ( .A1(n19134), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10769) );
  MUX2_X1 U13606 ( .A(n19134), .B(n10749), .S(n10778), .Z(n10750) );
  OR2_X1 U13607 ( .A1(n10778), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10781) );
  NAND2_X1 U13608 ( .A1(n10750), .A2(n10781), .ZN(n18808) );
  INV_X1 U13609 ( .A(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n15387) );
  NAND2_X1 U13610 ( .A1(n10795), .A2(n15387), .ZN(n15220) );
  AND2_X1 U13611 ( .A1(n19134), .A2(P2_EBX_REG_16__SCAN_IN), .ZN(n10752) );
  INV_X1 U13612 ( .A(n12555), .ZN(n10751) );
  AOI21_X1 U13613 ( .B1(n10759), .B2(n10752), .A(n10751), .ZN(n10754) );
  AND2_X1 U13614 ( .A1(n10754), .A2(n10753), .ZN(n10755) );
  NAND2_X1 U13615 ( .A1(n10790), .A2(n15187), .ZN(n15179) );
  INV_X1 U13616 ( .A(n10755), .ZN(n18832) );
  INV_X1 U13617 ( .A(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15405) );
  OAI21_X1 U13618 ( .B1(n18832), .B2(n15176), .A(n15405), .ZN(n10756) );
  INV_X1 U13619 ( .A(P2_EBX_REG_14__SCAN_IN), .ZN(n13898) );
  NAND2_X1 U13620 ( .A1(n10773), .A2(n13898), .ZN(n10758) );
  AND2_X1 U13621 ( .A1(n19134), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10757) );
  NAND2_X1 U13622 ( .A1(n10758), .A2(n10757), .ZN(n10760) );
  NAND2_X1 U13623 ( .A1(n10760), .A2(n10759), .ZN(n18841) );
  OR2_X1 U13624 ( .A1(n18841), .A2(n15176), .ZN(n10761) );
  INV_X1 U13625 ( .A(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15428) );
  NAND2_X1 U13626 ( .A1(n10761), .A2(n15428), .ZN(n15248) );
  INV_X1 U13627 ( .A(n10762), .ZN(n10763) );
  XNOR2_X1 U13628 ( .A(n10764), .B(n10763), .ZN(n18855) );
  NAND2_X1 U13629 ( .A1(n18855), .A2(n15187), .ZN(n10765) );
  INV_X1 U13630 ( .A(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n15443) );
  NAND2_X1 U13631 ( .A1(n10765), .A2(n15443), .ZN(n15172) );
  INV_X1 U13632 ( .A(n10766), .ZN(n10767) );
  INV_X1 U13633 ( .A(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n15470) );
  NAND2_X1 U13634 ( .A1(n10767), .A2(n15470), .ZN(n15466) );
  NAND2_X1 U13635 ( .A1(n10768), .A2(n15461), .ZN(n15169) );
  AND4_X1 U13636 ( .A1(n15248), .A2(n15172), .A3(n15466), .A4(n15169), .ZN(
        n10774) );
  OR2_X1 U13637 ( .A1(n10770), .A2(n10769), .ZN(n10771) );
  NAND2_X1 U13638 ( .A1(n10778), .A2(n10771), .ZN(n18820) );
  INV_X1 U13639 ( .A(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n15411) );
  NAND2_X1 U13640 ( .A1(n10798), .A2(n15411), .ZN(n15180) );
  AND2_X1 U13641 ( .A1(n19134), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10772) );
  XNOR2_X1 U13642 ( .A(n10773), .B(n10772), .ZN(n14017) );
  NAND2_X1 U13643 ( .A1(n14017), .A2(n15187), .ZN(n15174) );
  INV_X1 U13644 ( .A(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n16196) );
  NAND2_X1 U13645 ( .A1(n15174), .A2(n16196), .ZN(n16132) );
  AND4_X1 U13646 ( .A1(n15238), .A2(n10774), .A3(n15180), .A4(n16132), .ZN(
        n10784) );
  INV_X1 U13647 ( .A(P2_EBX_REG_19__SCAN_IN), .ZN(n10775) );
  INV_X1 U13648 ( .A(P2_EBX_REG_18__SCAN_IN), .ZN(n14116) );
  NAND2_X1 U13649 ( .A1(n10775), .A2(n14116), .ZN(n10776) );
  AND2_X1 U13650 ( .A1(n19134), .A2(n10776), .ZN(n10777) );
  NAND2_X1 U13651 ( .A1(n19134), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10779) );
  XNOR2_X1 U13652 ( .A(n10786), .B(n10779), .ZN(n13240) );
  NAND2_X1 U13653 ( .A1(n13240), .A2(n15187), .ZN(n10796) );
  INV_X1 U13654 ( .A(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n15357) );
  NAND2_X1 U13655 ( .A1(n10796), .A2(n15357), .ZN(n15185) );
  AND2_X1 U13656 ( .A1(n19134), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n10780) );
  NAND2_X1 U13657 ( .A1(n10781), .A2(n10780), .ZN(n10782) );
  NAND2_X1 U13658 ( .A1(n10782), .A2(n10786), .ZN(n18794) );
  OR2_X1 U13659 ( .A1(n18794), .A2(n15176), .ZN(n10783) );
  INV_X1 U13660 ( .A(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15374) );
  NAND2_X1 U13661 ( .A1(n10783), .A2(n15374), .ZN(n15207) );
  AND4_X1 U13662 ( .A1(n15220), .A2(n10784), .A3(n15185), .A4(n15207), .ZN(
        n10785) );
  INV_X1 U13663 ( .A(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n15189) );
  NOR2_X2 U13664 ( .A1(n10786), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n10788) );
  INV_X1 U13665 ( .A(P2_EBX_REG_21__SCAN_IN), .ZN(n15007) );
  NAND2_X1 U13666 ( .A1(n19134), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10787) );
  NOR2_X1 U13667 ( .A1(n10788), .A2(n10787), .ZN(n10789) );
  NOR2_X1 U13668 ( .A1(n10801), .A2(n10789), .ZN(n15188) );
  INV_X1 U13669 ( .A(n10790), .ZN(n10793) );
  NAND2_X1 U13670 ( .A1(n14017), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n10792) );
  OR2_X1 U13671 ( .A1(n18841), .A2(n15428), .ZN(n15177) );
  NAND2_X1 U13672 ( .A1(n18855), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n10791) );
  NAND2_X1 U13673 ( .A1(n15187), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10797) );
  OR2_X1 U13674 ( .A1(n18794), .A2(n10797), .ZN(n15206) );
  INV_X1 U13675 ( .A(n10798), .ZN(n10799) );
  NAND2_X1 U13676 ( .A1(n10799), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(
        n15181) );
  NAND2_X1 U13677 ( .A1(n19134), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10800) );
  NAND3_X1 U13678 ( .A1(n10802), .A2(n19134), .A3(P2_EBX_REG_22__SCAN_IN), 
        .ZN(n10803) );
  NAND2_X1 U13679 ( .A1(n10808), .A2(n10803), .ZN(n15680) );
  INV_X1 U13680 ( .A(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15338) );
  NAND2_X1 U13681 ( .A1(n10804), .A2(n15338), .ZN(n15326) );
  NOR2_X1 U13682 ( .A1(n10804), .A2(n15338), .ZN(n15328) );
  AND2_X1 U13683 ( .A1(n19134), .A2(P2_EBX_REG_23__SCAN_IN), .ZN(n10807) );
  XOR2_X1 U13684 ( .A(n10807), .B(n10808), .Z(n16094) );
  NAND2_X1 U13685 ( .A1(n16094), .A2(n15187), .ZN(n10805) );
  XOR2_X1 U13686 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B(n10805), .Z(
        n15156) );
  INV_X1 U13687 ( .A(n10805), .ZN(n10806) );
  NAND3_X1 U13688 ( .A1(n10809), .A2(P2_EBX_REG_24__SCAN_IN), .A3(n19134), 
        .ZN(n10810) );
  NAND2_X1 U13689 ( .A1(n10810), .A2(n12555), .ZN(n10811) );
  NOR2_X1 U13690 ( .A1(n10815), .A2(n10811), .ZN(n16083) );
  NAND2_X1 U13691 ( .A1(n16083), .A2(n15187), .ZN(n15144) );
  INV_X1 U13692 ( .A(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n15301) );
  INV_X1 U13693 ( .A(P2_EBX_REG_25__SCAN_IN), .ZN(n14974) );
  NOR2_X1 U13694 ( .A1(n10815), .A2(n14974), .ZN(n10812) );
  NAND2_X1 U13695 ( .A1(n19134), .A2(n10812), .ZN(n10813) );
  NAND2_X1 U13696 ( .A1(n12555), .A2(n10813), .ZN(n10814) );
  AOI21_X1 U13697 ( .B1(n10815), .B2(n14974), .A(n10814), .ZN(n16073) );
  AND2_X1 U13698 ( .A1(n16073), .A2(n15187), .ZN(n10826) );
  AND2_X1 U13699 ( .A1(P2_EBX_REG_26__SCAN_IN), .A2(n10816), .ZN(n10817) );
  AOI21_X1 U13700 ( .B1(n19134), .B2(n10817), .A(n10820), .ZN(n10818) );
  NAND2_X1 U13701 ( .A1(n12555), .A2(n10818), .ZN(n16062) );
  INV_X1 U13702 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n15120) );
  OAI21_X1 U13703 ( .B1(n16062), .B2(n15176), .A(n15120), .ZN(n10819) );
  NAND2_X1 U13704 ( .A1(n10819), .A2(n10829), .ZN(n15123) );
  NAND2_X1 U13705 ( .A1(n19134), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n10821) );
  NAND3_X1 U13706 ( .A1(n19134), .A2(P2_EBX_REG_27__SCAN_IN), .A3(n10822), 
        .ZN(n10823) );
  NAND2_X1 U13707 ( .A1(n10824), .A2(n10823), .ZN(n16052) );
  NAND2_X1 U13708 ( .A1(n15094), .A2(n10299), .ZN(n10825) );
  NAND2_X1 U13709 ( .A1(n19134), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n10830) );
  XNOR2_X1 U13710 ( .A(n10831), .B(n10830), .ZN(n16039) );
  INV_X1 U13711 ( .A(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n15263) );
  INV_X1 U13712 ( .A(n10826), .ZN(n10828) );
  INV_X1 U13713 ( .A(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n10827) );
  NAND2_X1 U13714 ( .A1(n15131), .A2(n10829), .ZN(n15093) );
  NAND2_X1 U13715 ( .A1(n19134), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n12535) );
  XNOR2_X1 U13716 ( .A(n12534), .B(n12535), .ZN(n10832) );
  INV_X1 U13717 ( .A(n10832), .ZN(n16026) );
  NAND3_X1 U13718 ( .A1(n16026), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A3(
        n15187), .ZN(n12550) );
  INV_X1 U13719 ( .A(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14239) );
  OAI21_X1 U13720 ( .B1(n10832), .B2(n15176), .A(n14239), .ZN(n12532) );
  INV_X1 U13721 ( .A(n12560), .ZN(n10833) );
  NOR3_X1 U13722 ( .A1(n12572), .A2(n12569), .A3(n10833), .ZN(n10837) );
  INV_X1 U13723 ( .A(n10837), .ZN(n10839) );
  NOR2_X1 U13724 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20934), .ZN(
        n10834) );
  XNOR2_X1 U13725 ( .A(n10846), .B(n10836), .ZN(n12565) );
  AND2_X1 U13726 ( .A1(n12565), .A2(n10837), .ZN(n10838) );
  OR2_X1 U13727 ( .A1(n12582), .A2(n10838), .ZN(n16255) );
  INV_X1 U13728 ( .A(n16255), .ZN(n12603) );
  OAI21_X1 U13729 ( .B1(n12564), .B2(n10839), .A(n12603), .ZN(n10841) );
  INV_X1 U13730 ( .A(n10572), .ZN(n10840) );
  AOI21_X1 U13731 ( .B1(n10546), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n15660) );
  AOI21_X1 U13732 ( .B1(n10840), .B2(n15660), .A(P2_FLUSH_REG_SCAN_IN), .ZN(
        n19816) );
  MUX2_X1 U13733 ( .A(n10841), .B(n19816), .S(P2_STATE2_REG_1__SCAN_IN), .Z(
        n19830) );
  INV_X1 U13734 ( .A(n10842), .ZN(n12614) );
  NAND2_X1 U13735 ( .A1(n12614), .A2(n13334), .ZN(n10851) );
  NAND2_X1 U13736 ( .A1(n12614), .A2(n10843), .ZN(n19826) );
  NAND2_X1 U13737 ( .A1(n10845), .A2(n10844), .ZN(n12576) );
  INV_X1 U13738 ( .A(n10846), .ZN(n12563) );
  NOR2_X1 U13739 ( .A1(n12563), .A2(n12564), .ZN(n10847) );
  NOR2_X1 U13740 ( .A1(n10848), .A2(n10847), .ZN(n10849) );
  NOR2_X1 U13741 ( .A1(n12576), .A2(n10849), .ZN(n10850) );
  OR2_X1 U13742 ( .A1(n10850), .A2(n12582), .ZN(n19827) );
  OAI22_X1 U13743 ( .A1(n19830), .A2(n10851), .B1(n19826), .B2(n19827), .ZN(
        n12608) );
  NAND2_X1 U13744 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15527), .ZN(n19707) );
  INV_X1 U13745 ( .A(n19707), .ZN(n10852) );
  NAND2_X1 U13746 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n10852), .ZN(n16292) );
  AND2_X1 U13747 ( .A1(n19114), .A2(n13386), .ZN(n10853) );
  NAND2_X1 U13748 ( .A1(n12608), .A2(n10853), .ZN(n13260) );
  INV_X1 U13749 ( .A(n13260), .ZN(n10891) );
  NAND2_X1 U13750 ( .A1(n10891), .A2(n13334), .ZN(n19108) );
  AND2_X1 U13751 ( .A1(n10854), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n13339) );
  INV_X1 U13752 ( .A(n10855), .ZN(n12677) );
  XOR2_X1 U13753 ( .A(n12671), .B(n12677), .Z(n10856) );
  NAND2_X1 U13754 ( .A1(n13339), .A2(n10856), .ZN(n10857) );
  XOR2_X1 U13755 ( .A(n10856), .B(n13339), .Z(n13376) );
  NAND2_X1 U13756 ( .A1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n13376), .ZN(
        n13375) );
  NAND2_X1 U13757 ( .A1(n10857), .A2(n13375), .ZN(n10859) );
  XNOR2_X1 U13758 ( .A(n9963), .B(n10859), .ZN(n13401) );
  XNOR2_X1 U13759 ( .A(n12683), .B(n10858), .ZN(n13400) );
  NAND2_X1 U13760 ( .A1(n13401), .A2(n13400), .ZN(n13399) );
  NAND2_X1 U13761 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n10859), .ZN(
        n10860) );
  NAND2_X1 U13762 ( .A1(n13399), .A2(n10860), .ZN(n10861) );
  XNOR2_X1 U13763 ( .A(n10861), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14249) );
  NAND2_X1 U13764 ( .A1(n10861), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n10862) );
  INV_X1 U13765 ( .A(n10863), .ZN(n10866) );
  INV_X1 U13766 ( .A(n10864), .ZN(n10865) );
  NAND2_X1 U13767 ( .A1(n10867), .A2(n12696), .ZN(n10869) );
  INV_X1 U13768 ( .A(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n13925) );
  INV_X1 U13769 ( .A(n10869), .ZN(n10870) );
  NAND2_X1 U13770 ( .A1(n10870), .A2(n12702), .ZN(n10872) );
  INV_X1 U13771 ( .A(n12706), .ZN(n10871) );
  NAND2_X1 U13772 ( .A1(n10872), .A2(n10871), .ZN(n10873) );
  INV_X1 U13774 ( .A(n10874), .ZN(n10875) );
  NAND2_X1 U13775 ( .A1(n10877), .A2(n10878), .ZN(n10880) );
  NAND2_X1 U13776 ( .A1(n10880), .A2(n10879), .ZN(n10881) );
  NAND2_X2 U13777 ( .A1(n13981), .A2(n10881), .ZN(n14077) );
  OAI21_X1 U13778 ( .B1(n10884), .B2(n15176), .A(n16207), .ZN(n10885) );
  NAND2_X1 U13779 ( .A1(n15187), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10883) );
  INV_X1 U13780 ( .A(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15487) );
  NOR2_X1 U13781 ( .A1(n15405), .A2(n15428), .ZN(n15161) );
  NAND3_X1 U13782 ( .A1(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n15403) );
  INV_X1 U13783 ( .A(n15403), .ZN(n10887) );
  NAND3_X1 U13784 ( .A1(n15161), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n10887), .ZN(n15379) );
  NOR2_X1 U13785 ( .A1(n15387), .A2(n15379), .ZN(n15358) );
  NAND3_X1 U13786 ( .A1(n15358), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n15347) );
  INV_X1 U13787 ( .A(n15347), .ZN(n10888) );
  AND2_X1 U13788 ( .A1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n10888), .ZN(
        n15312) );
  AND2_X1 U13789 ( .A1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n10889) );
  AND2_X1 U13790 ( .A1(n15312), .A2(n10889), .ZN(n12853) );
  INV_X1 U13791 ( .A(n15119), .ZN(n10890) );
  INV_X1 U13792 ( .A(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n21005) );
  AOI21_X1 U13793 ( .B1(n14239), .B2(n15105), .A(n12615), .ZN(n14246) );
  NAND2_X1 U13794 ( .A1(n10891), .A2(n16281), .ZN(n19092) );
  INV_X1 U13795 ( .A(n19092), .ZN(n19102) );
  NAND2_X1 U13796 ( .A1(n12543), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n10896) );
  INV_X1 U13797 ( .A(P2_REIP_REG_12__SCAN_IN), .ZN(n12779) );
  NAND2_X1 U13798 ( .A1(n12622), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n10893) );
  NAND2_X1 U13799 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n10892) );
  OAI211_X1 U13800 ( .C1(n9847), .C2(n12779), .A(n10893), .B(n10892), .ZN(
        n10894) );
  INV_X1 U13801 ( .A(n10894), .ZN(n10895) );
  NAND2_X1 U13802 ( .A1(n10896), .A2(n10895), .ZN(n13809) );
  NAND2_X1 U13803 ( .A1(n12543), .A2(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n10901) );
  INV_X1 U13804 ( .A(P2_REIP_REG_8__SCAN_IN), .ZN(n14050) );
  NAND2_X1 U13805 ( .A1(n12622), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n10898) );
  NAND2_X1 U13806 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n10897) );
  OAI211_X1 U13807 ( .C1(n9847), .C2(n14050), .A(n10898), .B(n10897), .ZN(
        n10899) );
  INV_X1 U13808 ( .A(n10899), .ZN(n10900) );
  NAND2_X1 U13809 ( .A1(n10901), .A2(n10900), .ZN(n13572) );
  INV_X1 U13810 ( .A(P2_REIP_REG_5__SCAN_IN), .ZN(n10904) );
  NAND2_X1 U13811 ( .A1(n12622), .A2(P2_EBX_REG_5__SCAN_IN), .ZN(n10903) );
  NAND2_X1 U13812 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n10902) );
  OAI211_X1 U13813 ( .C1(n9847), .C2(n10904), .A(n10903), .B(n10902), .ZN(
        n10905) );
  AOI21_X1 U13814 ( .B1(n12543), .B2(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .A(
        n10905), .ZN(n13630) );
  INV_X1 U13815 ( .A(P2_REIP_REG_4__SCAN_IN), .ZN(n12700) );
  AOI22_X1 U13816 ( .A1(n12622), .A2(P2_EBX_REG_4__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n10908) );
  OAI211_X1 U13817 ( .C1(n12700), .C2(n9847), .A(n10909), .B(n10908), .ZN(
        n13587) );
  NAND2_X1 U13818 ( .A1(n13588), .A2(n13587), .ZN(n13629) );
  INV_X1 U13819 ( .A(P2_REIP_REG_6__SCAN_IN), .ZN(n10912) );
  NAND2_X1 U13820 ( .A1(n12543), .A2(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10911) );
  AOI22_X1 U13821 ( .A1(n12622), .A2(P2_EBX_REG_6__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n10910) );
  OAI211_X1 U13822 ( .C1(n9847), .C2(n10912), .A(n10911), .B(n10910), .ZN(
        n13640) );
  INV_X1 U13823 ( .A(P2_REIP_REG_7__SCAN_IN), .ZN(n10916) );
  NAND2_X1 U13824 ( .A1(n12622), .A2(P2_EBX_REG_7__SCAN_IN), .ZN(n10915) );
  NAND2_X1 U13825 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n10914) );
  OAI211_X1 U13826 ( .C1(n9847), .C2(n10916), .A(n10915), .B(n10914), .ZN(
        n10917) );
  AOI21_X1 U13827 ( .B1(n12543), .B2(P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(
        n10917), .ZN(n13527) );
  INV_X1 U13828 ( .A(P2_REIP_REG_9__SCAN_IN), .ZN(n14218) );
  NAND2_X1 U13829 ( .A1(n12543), .A2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10919) );
  AOI22_X1 U13830 ( .A1(n12622), .A2(P2_EBX_REG_9__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n10918) );
  OAI211_X1 U13831 ( .C1(n9847), .C2(n14218), .A(n10919), .B(n10918), .ZN(
        n13704) );
  INV_X1 U13832 ( .A(P2_REIP_REG_10__SCAN_IN), .ZN(n12751) );
  NAND2_X1 U13833 ( .A1(n12543), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n10921) );
  AOI22_X1 U13834 ( .A1(n12622), .A2(P2_EBX_REG_10__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), 
        .ZN(n10920) );
  OAI211_X1 U13835 ( .C1(n9847), .C2(n12751), .A(n10921), .B(n10920), .ZN(
        n13741) );
  INV_X1 U13836 ( .A(P2_REIP_REG_11__SCAN_IN), .ZN(n12765) );
  NAND2_X1 U13837 ( .A1(n12622), .A2(P2_EBX_REG_11__SCAN_IN), .ZN(n10923) );
  NAND2_X1 U13838 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n10922) );
  OAI211_X1 U13839 ( .C1(n9847), .C2(n12765), .A(n10923), .B(n10922), .ZN(
        n10924) );
  AOI21_X1 U13840 ( .B1(n12543), .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        n10924), .ZN(n13795) );
  NAND2_X1 U13841 ( .A1(n13809), .A2(n13796), .ZN(n13842) );
  INV_X1 U13842 ( .A(P2_REIP_REG_13__SCAN_IN), .ZN(n12793) );
  NAND2_X1 U13843 ( .A1(n12622), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n10926) );
  NAND2_X1 U13844 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n10925) );
  OAI211_X1 U13845 ( .C1(n9847), .C2(n12793), .A(n10926), .B(n10925), .ZN(
        n10927) );
  AOI21_X1 U13846 ( .B1(n12543), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n10927), .ZN(n13841) );
  INV_X1 U13847 ( .A(P2_REIP_REG_14__SCAN_IN), .ZN(n14023) );
  NAND2_X1 U13848 ( .A1(n12622), .A2(P2_EBX_REG_14__SCAN_IN), .ZN(n10930) );
  NAND2_X1 U13849 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n10929) );
  OAI211_X1 U13850 ( .C1(n9847), .C2(n14023), .A(n10930), .B(n10929), .ZN(
        n10931) );
  AOI21_X1 U13851 ( .B1(n12543), .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n10931), .ZN(n13895) );
  INV_X1 U13852 ( .A(P2_REIP_REG_15__SCAN_IN), .ZN(n19747) );
  NAND2_X1 U13853 ( .A1(n12622), .A2(P2_EBX_REG_15__SCAN_IN), .ZN(n10934) );
  NAND2_X1 U13854 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n10933) );
  OAI211_X1 U13855 ( .C1(n9847), .C2(n19747), .A(n10934), .B(n10933), .ZN(
        n10935) );
  AOI21_X1 U13856 ( .B1(n12543), .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .A(
        n10935), .ZN(n13913) );
  INV_X1 U13857 ( .A(P2_REIP_REG_16__SCAN_IN), .ZN(n15415) );
  NAND2_X1 U13858 ( .A1(n12543), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n10937) );
  AOI22_X1 U13859 ( .A1(n12622), .A2(P2_EBX_REG_16__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n10936) );
  OAI211_X1 U13860 ( .C1(n9847), .C2(n15415), .A(n10937), .B(n10936), .ZN(
        n13966) );
  INV_X1 U13861 ( .A(P2_REIP_REG_17__SCAN_IN), .ZN(n19750) );
  NAND2_X1 U13862 ( .A1(n12622), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n10939) );
  NAND2_X1 U13863 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n10938) );
  OAI211_X1 U13864 ( .C1(n9847), .C2(n19750), .A(n10939), .B(n10938), .ZN(
        n10940) );
  AOI21_X1 U13865 ( .B1(n12543), .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A(
        n10940), .ZN(n14001) );
  INV_X1 U13866 ( .A(P2_REIP_REG_18__SCAN_IN), .ZN(n19752) );
  NAND2_X1 U13867 ( .A1(n12622), .A2(P2_EBX_REG_18__SCAN_IN), .ZN(n10944) );
  NAND2_X1 U13868 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n10943) );
  OAI211_X1 U13869 ( .C1(n9847), .C2(n19752), .A(n10944), .B(n10943), .ZN(
        n10945) );
  INV_X1 U13870 ( .A(P2_REIP_REG_19__SCAN_IN), .ZN(n19754) );
  NAND2_X1 U13871 ( .A1(n12543), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n10947) );
  AOI22_X1 U13872 ( .A1(n12622), .A2(P2_EBX_REG_19__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), 
        .ZN(n10946) );
  OAI211_X1 U13873 ( .C1(n9847), .C2(n19754), .A(n10947), .B(n10946), .ZN(
        n14098) );
  INV_X1 U13874 ( .A(P2_REIP_REG_20__SCAN_IN), .ZN(n19756) );
  NAND2_X1 U13875 ( .A1(n12543), .A2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n10949) );
  AOI22_X1 U13876 ( .A1(n12622), .A2(P2_EBX_REG_20__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), 
        .ZN(n10948) );
  OAI211_X1 U13877 ( .C1(n9847), .C2(n19756), .A(n10949), .B(n10948), .ZN(
        n13236) );
  INV_X1 U13878 ( .A(P2_REIP_REG_21__SCAN_IN), .ZN(n19758) );
  NAND2_X1 U13879 ( .A1(n12622), .A2(P2_EBX_REG_21__SCAN_IN), .ZN(n10951) );
  NAND2_X1 U13880 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n10950) );
  OAI211_X1 U13881 ( .C1(n9847), .C2(n19758), .A(n10951), .B(n10950), .ZN(
        n10952) );
  AOI21_X1 U13882 ( .B1(n12543), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n10952), .ZN(n14869) );
  INV_X1 U13883 ( .A(P2_REIP_REG_22__SCAN_IN), .ZN(n12830) );
  NAND2_X1 U13884 ( .A1(n12622), .A2(P2_EBX_REG_22__SCAN_IN), .ZN(n10956) );
  NAND2_X1 U13885 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n10955) );
  OAI211_X1 U13886 ( .C1(n9847), .C2(n12830), .A(n10956), .B(n10955), .ZN(
        n10957) );
  AOI21_X1 U13887 ( .B1(n12543), .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .A(
        n10957), .ZN(n15000) );
  INV_X1 U13888 ( .A(P2_REIP_REG_23__SCAN_IN), .ZN(n10960) );
  NAND2_X1 U13889 ( .A1(n12543), .A2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n10959) );
  AOI22_X1 U13890 ( .A1(n12622), .A2(P2_EBX_REG_23__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_23__SCAN_IN), 
        .ZN(n10958) );
  OAI211_X1 U13891 ( .C1(n9847), .C2(n10960), .A(n10959), .B(n10958), .ZN(
        n14992) );
  INV_X1 U13892 ( .A(P2_REIP_REG_24__SCAN_IN), .ZN(n10963) );
  NAND2_X1 U13893 ( .A1(n12622), .A2(P2_EBX_REG_24__SCAN_IN), .ZN(n10962) );
  NAND2_X1 U13894 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n10961) );
  OAI211_X1 U13895 ( .C1(n9847), .C2(n10963), .A(n10962), .B(n10961), .ZN(
        n10964) );
  AOI21_X1 U13896 ( .B1(n12543), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n10964), .ZN(n14983) );
  INV_X1 U13897 ( .A(P2_REIP_REG_25__SCAN_IN), .ZN(n19763) );
  NAND2_X1 U13898 ( .A1(n12622), .A2(P2_EBX_REG_25__SCAN_IN), .ZN(n10966) );
  NAND2_X1 U13899 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n10965) );
  OAI211_X1 U13900 ( .C1(n9847), .C2(n19763), .A(n10966), .B(n10965), .ZN(
        n10967) );
  AOI21_X1 U13901 ( .B1(n12543), .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n10967), .ZN(n14971) );
  INV_X1 U13902 ( .A(P2_REIP_REG_26__SCAN_IN), .ZN(n21017) );
  NAND2_X1 U13903 ( .A1(n12622), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n10969) );
  NAND2_X1 U13904 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(
        P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n10968) );
  OAI211_X1 U13905 ( .C1(n9847), .C2(n21017), .A(n10969), .B(n10968), .ZN(
        n10970) );
  AOI21_X1 U13906 ( .B1(n12543), .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        n10970), .ZN(n14959) );
  INV_X1 U13907 ( .A(P2_REIP_REG_27__SCAN_IN), .ZN(n19767) );
  NAND2_X1 U13908 ( .A1(n12543), .A2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n10972) );
  AOI22_X1 U13909 ( .A1(n12622), .A2(P2_EBX_REG_27__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_27__SCAN_IN), 
        .ZN(n10971) );
  OAI211_X1 U13910 ( .C1(n9847), .C2(n19767), .A(n10972), .B(n10971), .ZN(
        n14953) );
  INV_X1 U13911 ( .A(P2_REIP_REG_28__SCAN_IN), .ZN(n19768) );
  NAND2_X1 U13912 ( .A1(n12543), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n10974) );
  AOI22_X1 U13913 ( .A1(n12622), .A2(P2_EBX_REG_28__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), 
        .ZN(n10973) );
  OAI211_X1 U13914 ( .C1(n9847), .C2(n19768), .A(n10974), .B(n10973), .ZN(
        n14948) );
  INV_X1 U13915 ( .A(P2_REIP_REG_29__SCAN_IN), .ZN(n19770) );
  NAND2_X1 U13916 ( .A1(n12543), .A2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n10976) );
  AOI22_X1 U13917 ( .A1(n12622), .A2(P2_EBX_REG_29__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), 
        .ZN(n10975) );
  OAI211_X1 U13918 ( .C1(n9847), .C2(n19770), .A(n10976), .B(n10975), .ZN(
        n10977) );
  OR2_X1 U13919 ( .A1(n14950), .A2(n10977), .ZN(n10978) );
  NAND2_X1 U13920 ( .A1(n12620), .A2(n10978), .ZN(n16028) );
  NOR2_X2 U13921 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19612) );
  NOR2_X1 U13922 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n15552) );
  OR2_X1 U13923 ( .A1(n19612), .A2(n15552), .ZN(n19806) );
  NAND2_X1 U13924 ( .A1(n19806), .A2(n10983), .ZN(n10979) );
  INV_X1 U13925 ( .A(P2_STATEBS16_REG_SCAN_IN), .ZN(n19836) );
  NOR2_X1 U13926 ( .A1(n15527), .A2(n19836), .ZN(n19807) );
  NAND2_X1 U13927 ( .A1(n15552), .A2(n19842), .ZN(n18766) );
  INV_X1 U13928 ( .A(n18766), .ZN(n10980) );
  AND2_X2 U13929 ( .A1(n10980), .A2(n10983), .ZN(n19085) );
  INV_X2 U13930 ( .A(n19085), .ZN(n18934) );
  NOR2_X1 U13931 ( .A1(n18934), .A2(n19770), .ZN(n14237) );
  AOI21_X1 U13932 ( .B1(n19086), .B2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A(
        n14237), .ZN(n10987) );
  INV_X1 U13933 ( .A(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n10982) );
  INV_X1 U13934 ( .A(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n15152) );
  INV_X1 U13935 ( .A(P2_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15163) );
  INV_X1 U13936 ( .A(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n15253) );
  INV_X1 U13937 ( .A(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n18819) );
  INV_X1 U13938 ( .A(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15138) );
  INV_X1 U13939 ( .A(P2_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n16049) );
  INV_X1 U13940 ( .A(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n15101) );
  INV_X1 U13941 ( .A(n15102), .ZN(n10981) );
  AND2_X2 U13942 ( .A1(n15102), .A2(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n13228) );
  AOI21_X1 U13943 ( .B1(n10982), .B2(n10981), .A(n13228), .ZN(n16002) );
  INV_X1 U13944 ( .A(n12881), .ZN(n10985) );
  NAND2_X1 U13945 ( .A1(n19836), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n10984) );
  NAND2_X1 U13946 ( .A1(n10985), .A2(n10984), .ZN(n13369) );
  NAND2_X1 U13947 ( .A1(n16002), .A2(n19101), .ZN(n10986) );
  OAI211_X1 U13948 ( .C1(n16028), .C2(n16174), .A(n10987), .B(n10986), .ZN(
        n10988) );
  AOI21_X1 U13949 ( .B1(n14246), .B2(n19102), .A(n10988), .ZN(n10989) );
  NOR2_X4 U13950 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13687) );
  NAND2_X1 U13952 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(
        n10994) );
  INV_X2 U13953 ( .A(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n14284) );
  NAND2_X1 U13954 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(
        n10993) );
  NOR2_X2 U13955 ( .A1(n14284), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n10999) );
  AND2_X2 U13956 ( .A1(n11004), .A2(n10999), .ZN(n11147) );
  NAND2_X1 U13957 ( .A1(n11147), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(
        n10992) );
  AND2_X2 U13958 ( .A1(n11005), .A2(n13687), .ZN(n11199) );
  NAND2_X1 U13959 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(
        n10991) );
  AND2_X4 U13960 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n13673) );
  NAND2_X1 U13961 ( .A1(n11356), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(
        n10998) );
  NAND2_X1 U13962 ( .A1(n11047), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(
        n10997) );
  NAND2_X1 U13963 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(
        n10996) );
  NAND2_X1 U13964 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(
        n10995) );
  AND2_X2 U13965 ( .A1(n11006), .A2(n13672), .ZN(n11240) );
  NAND2_X1 U13966 ( .A1(n11240), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(
        n11003) );
  NAND2_X1 U13967 ( .A1(n12465), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(
        n11002) );
  NAND2_X1 U13968 ( .A1(n11098), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(
        n11001) );
  NAND2_X2 U13969 ( .A1(n13673), .A2(n13672), .ZN(n13668) );
  INV_X2 U13970 ( .A(n13668), .ZN(n12294) );
  NAND2_X1 U13971 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(
        n11000) );
  NAND2_X1 U13972 ( .A1(n11193), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(
        n11010) );
  NAND2_X1 U13973 ( .A1(n11245), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(
        n11009) );
  NAND2_X1 U13974 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(
        n11008) );
  NAND2_X1 U13975 ( .A1(n11246), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(
        n11007) );
  NAND2_X1 U13976 ( .A1(n11240), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(
        n11018) );
  NAND2_X1 U13977 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(
        n11017) );
  NAND2_X1 U13978 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(
        n11016) );
  NAND2_X1 U13979 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(
        n11015) );
  NAND2_X1 U13980 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(
        n11022) );
  NAND2_X1 U13981 ( .A1(n12465), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(
        n11021) );
  NAND2_X1 U13982 ( .A1(n11147), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(
        n11020) );
  NAND2_X1 U13983 ( .A1(n9843), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(
        n11019) );
  NAND2_X1 U13984 ( .A1(n11047), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(
        n11026) );
  NAND2_X1 U13985 ( .A1(n11245), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(
        n11025) );
  NAND2_X1 U13986 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(
        n11024) );
  NAND2_X1 U13987 ( .A1(n11246), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(
        n11023) );
  NAND2_X1 U13988 ( .A1(n11193), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(
        n11030) );
  NAND2_X1 U13989 ( .A1(n11356), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(
        n11029) );
  NAND2_X1 U13990 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n11028) );
  NAND2_X1 U13991 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(
        n11027) );
  NAND4_X4 U13992 ( .A1(n11034), .A2(n11033), .A3(n11032), .A4(n11031), .ZN(
        n20122) );
  NAND2_X1 U13993 ( .A1(n11193), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n11038) );
  NAND2_X1 U13994 ( .A1(n11356), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(
        n11037) );
  NAND2_X1 U13995 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n11036) );
  NAND2_X1 U13996 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(
        n11035) );
  NAND2_X1 U13997 ( .A1(n11240), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n11042) );
  NAND2_X1 U13998 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(
        n11041) );
  NAND2_X1 U13999 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(
        n11040) );
  NAND2_X1 U14000 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(
        n11039) );
  NAND4_X1 U14001 ( .A1(n11042), .A2(n11041), .A3(n11040), .A4(n11039), .ZN(
        n11055) );
  NAND2_X1 U14002 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(
        n11046) );
  NAND2_X1 U14003 ( .A1(n12465), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n11045) );
  NAND2_X1 U14004 ( .A1(n11147), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(
        n11044) );
  NAND2_X1 U14005 ( .A1(n11098), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n11043) );
  NAND2_X1 U14006 ( .A1(n11047), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(
        n11051) );
  NAND2_X1 U14007 ( .A1(n11245), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(
        n11050) );
  NAND2_X1 U14008 ( .A1(n9835), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(
        n11049) );
  NAND2_X1 U14009 ( .A1(n11246), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(
        n11048) );
  NAND2_X1 U14010 ( .A1(n11053), .A2(n11052), .ZN(n11054) );
  NOR2_X1 U14011 ( .A1(n11055), .A2(n11054), .ZN(n11056) );
  NAND2_X4 U14012 ( .A1(n11057), .A2(n11056), .ZN(n11501) );
  NAND2_X1 U14013 ( .A1(n11356), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(
        n11061) );
  NAND2_X1 U14014 ( .A1(n11047), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(
        n11060) );
  NAND2_X1 U14015 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(
        n11059) );
  NAND2_X1 U14016 ( .A1(n11153), .A2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(
        n11058) );
  NAND2_X1 U14017 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(
        n11065) );
  NAND2_X1 U14018 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(
        n11064) );
  NAND2_X1 U14019 ( .A1(n12465), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(
        n11063) );
  NAND2_X1 U14020 ( .A1(n11098), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(
        n11062) );
  NAND2_X1 U14021 ( .A1(n11240), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(
        n11069) );
  NAND2_X1 U14022 ( .A1(n11147), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(
        n11068) );
  NAND2_X1 U14023 ( .A1(n11199), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(
        n11067) );
  NAND2_X1 U14024 ( .A1(n12294), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(
        n11066) );
  AND4_X2 U14025 ( .A1(n11069), .A2(n11068), .A3(n11067), .A4(n11066), .ZN(
        n11075) );
  NAND2_X1 U14026 ( .A1(n11193), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(
        n11073) );
  NAND2_X1 U14027 ( .A1(n11245), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(
        n11072) );
  NAND2_X1 U14028 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11071) );
  NAND2_X1 U14029 ( .A1(n11246), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(
        n11070) );
  NAND4_X4 U14030 ( .A1(n11077), .A2(n11076), .A3(n11075), .A4(n11074), .ZN(
        n11180) );
  AOI22_X1 U14031 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .B1(
        n11240), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11081) );
  AOI22_X1 U14032 ( .A1(n12465), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11199), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11080) );
  AOI22_X1 U14033 ( .A1(n11147), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n9843), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11079) );
  AOI22_X1 U14034 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n12468), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11078) );
  NAND4_X1 U14035 ( .A1(n11081), .A2(n11080), .A3(n11079), .A4(n11078), .ZN(
        n11087) );
  AOI22_X1 U14036 ( .A1(n11047), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n11194), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n11085) );
  AOI22_X1 U14037 ( .A1(n11356), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11283), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11084) );
  AOI22_X1 U14038 ( .A1(n11193), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11153), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11083) );
  AOI22_X1 U14039 ( .A1(n11245), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n11246), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n11082) );
  NAND4_X1 U14040 ( .A1(n11085), .A2(n11084), .A3(n11083), .A4(n11082), .ZN(
        n11086) );
  OR2_X2 U14041 ( .A1(n11087), .A2(n11086), .ZN(n20129) );
  AND2_X2 U14042 ( .A1(n20129), .A2(n20122), .ZN(n11500) );
  NAND2_X1 U14043 ( .A1(n13267), .A2(n11500), .ZN(n11097) );
  AOI22_X1 U14044 ( .A1(n12465), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11110), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11091) );
  AOI22_X1 U14045 ( .A1(n11147), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11356), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11090) );
  AOI22_X1 U14046 ( .A1(n11193), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11047), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11089) );
  AOI22_X1 U14047 ( .A1(n11245), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n11246), .B2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11088) );
  AOI22_X1 U14048 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n11199), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11095) );
  AOI22_X1 U14049 ( .A1(n11098), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11283), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11094) );
  AOI22_X1 U14050 ( .A1(n11194), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11153), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11093) );
  AOI22_X1 U14051 ( .A1(n11240), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11092) );
  NAND2_X2 U14052 ( .A1(n10312), .A2(n10314), .ZN(n11108) );
  NAND2_X1 U14053 ( .A1(n11108), .A2(n11501), .ZN(n11608) );
  OAI211_X1 U14054 ( .C1(n11176), .C2(n20793), .A(n11097), .B(n11096), .ZN(
        n11139) );
  NOR2_X1 U14055 ( .A1(n11139), .A2(n13656), .ZN(n11131) );
  AOI22_X1 U14056 ( .A1(n11147), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11098), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11102) );
  AOI22_X1 U14057 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n11240), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11101) );
  AOI22_X1 U14058 ( .A1(n12465), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11199), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11100) );
  AOI22_X1 U14059 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11099) );
  AOI22_X1 U14060 ( .A1(n11047), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n9836), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n11106) );
  AOI22_X1 U14061 ( .A1(n11193), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11153), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11105) );
  AOI22_X1 U14062 ( .A1(n11356), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11283), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11104) );
  AOI22_X1 U14063 ( .A1(n11245), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11246), .B2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11103) );
  NAND2_X2 U14064 ( .A1(n10313), .A2(n11107), .ZN(n11120) );
  NOR2_X2 U14065 ( .A1(n11487), .A2(n12498), .ZN(n13269) );
  AOI22_X1 U14066 ( .A1(n11283), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11153), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11114) );
  AOI22_X1 U14067 ( .A1(n12465), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n11110), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11113) );
  AOI22_X1 U14068 ( .A1(n11193), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n11194), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n11112) );
  AOI22_X1 U14069 ( .A1(n11147), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n9843), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11111) );
  AOI22_X1 U14070 ( .A1(n11299), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n11199), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11118) );
  AOI22_X1 U14071 ( .A1(n11356), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11047), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11117) );
  AOI22_X1 U14072 ( .A1(n11240), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11116) );
  AOI22_X1 U14073 ( .A1(n11245), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11246), .B2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n11115) );
  AND2_X2 U14074 ( .A1(n13269), .A2(n20145), .ZN(n11596) );
  INV_X1 U14075 ( .A(P1_STATE_REG_2__SCAN_IN), .ZN(n11119) );
  XNOR2_X1 U14076 ( .A(n11119), .B(P1_STATE_REG_1__SCAN_IN), .ZN(n11482) );
  NAND2_X1 U14077 ( .A1(n14280), .A2(n20129), .ZN(n11125) );
  NAND2_X1 U14078 ( .A1(n11491), .A2(n11180), .ZN(n11210) );
  NAND2_X1 U14079 ( .A1(n11210), .A2(n14171), .ZN(n11122) );
  OAI21_X1 U14080 ( .B1(n11120), .B2(n11123), .A(n11122), .ZN(n11124) );
  INV_X1 U14081 ( .A(n11180), .ZN(n11428) );
  NAND2_X1 U14082 ( .A1(n11428), .A2(n11120), .ZN(n11128) );
  AND2_X1 U14083 ( .A1(n11128), .A2(n20145), .ZN(n11135) );
  NAND2_X1 U14084 ( .A1(n11473), .A2(n14280), .ZN(n11130) );
  NAND4_X1 U14085 ( .A1(n11131), .A2(n11186), .A3(n11610), .A4(n11130), .ZN(
        n11132) );
  INV_X1 U14086 ( .A(n20689), .ZN(n11133) );
  NAND2_X1 U14087 ( .A1(n14858), .A2(n11192), .ZN(n13622) );
  MUX2_X1 U14088 ( .A(n11133), .B(n13622), .S(n20551), .Z(n11134) );
  INV_X1 U14089 ( .A(n11135), .ZN(n11137) );
  INV_X1 U14090 ( .A(n13265), .ZN(n14427) );
  NAND2_X1 U14091 ( .A1(n13486), .A2(n20129), .ZN(n11136) );
  AOI22_X1 U14092 ( .A1(n11137), .A2(n11391), .B1(n13280), .B2(n11136), .ZN(
        n11142) );
  INV_X1 U14093 ( .A(n13656), .ZN(n13669) );
  OR2_X1 U14094 ( .A1(n13669), .A2(n11120), .ZN(n11601) );
  NAND3_X1 U14095 ( .A1(n11601), .A2(n14858), .A3(P1_STATE2_REG_0__SCAN_IN), 
        .ZN(n11138) );
  NOR2_X1 U14096 ( .A1(n11139), .A2(n11138), .ZN(n11141) );
  NAND3_X1 U14097 ( .A1(n11473), .A2(n20122), .A3(n14280), .ZN(n11140) );
  NAND4_X1 U14098 ( .A1(n11142), .A2(n11610), .A3(n11141), .A4(n11140), .ZN(
        n11143) );
  AOI22_X1 U14099 ( .A1(n12458), .A2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n11146), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11151) );
  AOI22_X1 U14100 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11150) );
  AOI22_X1 U14101 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n11149) );
  AOI22_X1 U14102 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n12468), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11148) );
  NAND4_X1 U14103 ( .A1(n11151), .A2(n11150), .A3(n11149), .A4(n11148), .ZN(
        n11161) );
  AOI22_X1 U14104 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11167), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n11159) );
  AOI22_X1 U14105 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n11158) );
  AOI22_X1 U14106 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11157) );
  AOI22_X1 U14107 ( .A1(n11245), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11156) );
  NAND4_X1 U14108 ( .A1(n11159), .A2(n11158), .A3(n11157), .A4(n11156), .ZN(
        n11160) );
  INV_X1 U14109 ( .A(n11390), .ZN(n11162) );
  NOR2_X1 U14110 ( .A1(n11278), .A2(n11390), .ZN(n11220) );
  AOI22_X1 U14111 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11166) );
  AOI22_X1 U14112 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11047), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11165) );
  AOI22_X1 U14113 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12468), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11164) );
  AOI22_X1 U14114 ( .A1(n12466), .A2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11163) );
  NAND4_X1 U14115 ( .A1(n11166), .A2(n11165), .A3(n11164), .A4(n11163), .ZN(
        n11173) );
  AOI22_X1 U14116 ( .A1(n12458), .A2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n11146), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11171) );
  AOI22_X1 U14117 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11167), .B2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n11170) );
  AOI22_X1 U14118 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11169) );
  AOI22_X1 U14119 ( .A1(n11245), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11168) );
  NAND4_X1 U14120 ( .A1(n11171), .A2(n11170), .A3(n11169), .A4(n11168), .ZN(
        n11172) );
  MUX2_X1 U14121 ( .A(n11219), .B(n11220), .S(n11259), .Z(n11174) );
  OAI21_X2 U14122 ( .B1(n14282), .B2(P1_STATE2_REG_0__SCAN_IN), .A(n11175), 
        .ZN(n11218) );
  INV_X1 U14123 ( .A(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n11179) );
  AOI21_X1 U14124 ( .B1(n11176), .B2(n11390), .A(n11192), .ZN(n11178) );
  NAND2_X1 U14125 ( .A1(n12498), .A2(n11259), .ZN(n11177) );
  OAI211_X1 U14126 ( .C1(n11438), .C2(n11179), .A(n11178), .B(n11177), .ZN(
        n11217) );
  NAND2_X1 U14127 ( .A1(n11180), .A2(n20122), .ZN(n11423) );
  INV_X1 U14128 ( .A(n11423), .ZN(n11181) );
  NAND2_X1 U14129 ( .A1(n12498), .A2(n20129), .ZN(n11263) );
  OAI21_X1 U14130 ( .B1(n20793), .B2(n11259), .A(n11263), .ZN(n11182) );
  INV_X1 U14131 ( .A(n11182), .ZN(n11183) );
  NAND2_X1 U14132 ( .A1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n11236) );
  OAI21_X1 U14133 ( .B1(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(
        P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A(n11236), .ZN(n20437) );
  NAND2_X1 U14134 ( .A1(n20689), .A2(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n11229) );
  OAI21_X1 U14135 ( .B1(n13622), .B2(n20437), .A(n11229), .ZN(n11184) );
  INV_X1 U14136 ( .A(n11184), .ZN(n11185) );
  NAND3_X1 U14137 ( .A1(n13656), .A2(n13265), .A3(n11428), .ZN(n13454) );
  INV_X1 U14138 ( .A(n14171), .ZN(n11488) );
  NAND2_X1 U14139 ( .A1(n11186), .A2(n11597), .ZN(n11187) );
  XNOR2_X2 U14140 ( .A(n11189), .B(n11228), .ZN(n20218) );
  INV_X1 U14141 ( .A(n20218), .ZN(n11190) );
  NAND2_X2 U14142 ( .A1(n20218), .A2(n11191), .ZN(n11233) );
  INV_X1 U14143 ( .A(P1_STATE2_REG_0__SCAN_IN), .ZN(n11192) );
  INV_X1 U14144 ( .A(n11278), .ZN(n11206) );
  AOI22_X1 U14145 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n12458), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11198) );
  AOI22_X1 U14146 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n11167), .B2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n11197) );
  AOI22_X1 U14147 ( .A1(n11245), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n11047), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n11196) );
  AOI22_X1 U14148 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n11195) );
  NAND4_X1 U14149 ( .A1(n11198), .A2(n11197), .A3(n11196), .A4(n11195), .ZN(
        n11205) );
  AOI22_X1 U14150 ( .A1(n12467), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n11203) );
  AOI22_X1 U14151 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12299), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n11202) );
  AOI22_X1 U14152 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n12468), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11201) );
  AOI22_X1 U14153 ( .A1(n12460), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11200) );
  NAND4_X1 U14154 ( .A1(n11203), .A2(n11202), .A3(n11201), .A4(n11200), .ZN(
        n11204) );
  NAND2_X1 U14155 ( .A1(n11206), .A2(n11260), .ZN(n11207) );
  INV_X1 U14156 ( .A(n11259), .ZN(n11209) );
  XNOR2_X1 U14157 ( .A(n11209), .B(n11260), .ZN(n11211) );
  AOI21_X1 U14158 ( .B1(n11211), .B2(n11391), .A(n11210), .ZN(n11212) );
  INV_X1 U14159 ( .A(n11213), .ZN(n11214) );
  OR2_X1 U14160 ( .A1(n20041), .A2(n11214), .ZN(n11215) );
  INV_X1 U14161 ( .A(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20069) );
  INV_X1 U14162 ( .A(n11219), .ZN(n11386) );
  INV_X1 U14163 ( .A(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11224) );
  INV_X1 U14164 ( .A(n11220), .ZN(n11223) );
  INV_X1 U14165 ( .A(n11277), .ZN(n11221) );
  NAND2_X1 U14166 ( .A1(n11221), .A2(n11260), .ZN(n11222) );
  OAI211_X1 U14167 ( .C1(n11224), .C2(n11438), .A(n11223), .B(n11222), .ZN(
        n11225) );
  INV_X1 U14168 ( .A(n11228), .ZN(n11231) );
  NAND2_X1 U14169 ( .A1(n11229), .A2(n13661), .ZN(n11230) );
  NAND2_X1 U14170 ( .A1(n11231), .A2(n11230), .ZN(n11232) );
  AND2_X1 U14171 ( .A1(n11236), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11237) );
  NOR2_X1 U14172 ( .A1(n11236), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n20480) );
  OR2_X1 U14173 ( .A1(n11237), .A2(n20480), .ZN(n20114) );
  INV_X1 U14174 ( .A(n13622), .ZN(n11274) );
  AOI22_X1 U14175 ( .A1(n20114), .A2(n11274), .B1(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n20689), .ZN(n11238) );
  AOI22_X1 U14176 ( .A1(n12458), .A2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n11146), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11244) );
  AOI22_X1 U14177 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n11243) );
  AOI22_X1 U14178 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11242) );
  AOI22_X1 U14179 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n12468), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11241) );
  NAND4_X1 U14180 ( .A1(n11244), .A2(n11243), .A3(n11242), .A4(n11241), .ZN(
        n11252) );
  AOI22_X1 U14181 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11167), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n11250) );
  AOI22_X1 U14182 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n11249) );
  AOI22_X1 U14183 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11248) );
  AOI22_X1 U14184 ( .A1(n11245), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11247) );
  NAND4_X1 U14185 ( .A1(n11250), .A2(n11249), .A3(n11248), .A4(n11247), .ZN(
        n11251) );
  INV_X1 U14186 ( .A(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n11253) );
  OAI22_X1 U14187 ( .A1(n11438), .A2(n11253), .B1(n11262), .B2(n11277), .ZN(
        n11254) );
  NAND2_X1 U14188 ( .A1(n11257), .A2(n11256), .ZN(n11258) );
  NAND2_X1 U14189 ( .A1(n11260), .A2(n11259), .ZN(n11261) );
  NAND2_X1 U14190 ( .A1(n11261), .A2(n11262), .ZN(n11314) );
  OAI21_X1 U14191 ( .B1(n11262), .B2(n11261), .A(n11314), .ZN(n11265) );
  INV_X1 U14192 ( .A(n11263), .ZN(n11264) );
  AOI21_X1 U14193 ( .B1(n11265), .B2(n11391), .A(n11264), .ZN(n11266) );
  NAND2_X1 U14194 ( .A1(n13733), .A2(n13732), .ZN(n11269) );
  NAND2_X1 U14195 ( .A1(n11267), .A2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n11268) );
  NAND2_X1 U14196 ( .A1(n11269), .A2(n11268), .ZN(n11296) );
  INV_X1 U14197 ( .A(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n13756) );
  INV_X1 U14198 ( .A(n11234), .ZN(n11271) );
  NAND2_X1 U14199 ( .A1(n11271), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n11276) );
  NAND3_X1 U14200 ( .A1(n20184), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20350) );
  INV_X1 U14201 ( .A(n20372), .ZN(n11273) );
  NOR3_X1 U14202 ( .A1(n20184), .A2(n20514), .A3(n20440), .ZN(n20638) );
  INV_X1 U14203 ( .A(n20638), .ZN(n20630) );
  NOR2_X1 U14204 ( .A1(n20551), .A2(n20630), .ZN(n11272) );
  AOI21_X1 U14205 ( .B1(n20184), .B2(n11273), .A(n11272), .ZN(n20381) );
  AOI22_X1 U14206 ( .A1(n20381), .A2(n11274), .B1(
        P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20689), .ZN(n11275) );
  XNOR2_X2 U14207 ( .A(n11270), .B(n20257), .ZN(n20771) );
  AOI22_X1 U14208 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n12458), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11282) );
  AOI22_X1 U14209 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n9831), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11281) );
  AOI22_X1 U14210 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11167), .B2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11280) );
  AOI22_X1 U14211 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11279) );
  NAND4_X1 U14212 ( .A1(n11282), .A2(n11281), .A3(n11280), .A4(n11279), .ZN(
        n11289) );
  AOI22_X1 U14213 ( .A1(n12467), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11287) );
  AOI22_X1 U14214 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11286) );
  AOI22_X1 U14215 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11285) );
  AOI22_X1 U14216 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n12468), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11284) );
  NAND4_X1 U14217 ( .A1(n11287), .A2(n11286), .A3(n11285), .A4(n11284), .ZN(
        n11288) );
  AOI22_X1 U14218 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n11461), .B1(
        n11466), .B2(n11313), .ZN(n11290) );
  NAND2_X1 U14219 ( .A1(n20766), .A2(n11181), .ZN(n11295) );
  INV_X1 U14220 ( .A(n11313), .ZN(n11292) );
  XNOR2_X1 U14221 ( .A(n11314), .B(n11292), .ZN(n11293) );
  NAND2_X1 U14222 ( .A1(n11293), .A2(n11391), .ZN(n11294) );
  NAND2_X1 U14223 ( .A1(n11295), .A2(n11294), .ZN(n13752) );
  NAND2_X1 U14224 ( .A1(n13753), .A2(n13752), .ZN(n11298) );
  NAND2_X1 U14225 ( .A1(n11296), .A2(P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n11297) );
  NAND2_X1 U14226 ( .A1(n11298), .A2(n11297), .ZN(n13820) );
  AOI22_X1 U14227 ( .A1(n12458), .A2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n11146), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11303) );
  AOI22_X1 U14228 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n11302) );
  AOI22_X1 U14229 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11301) );
  AOI22_X1 U14230 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12468), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11300) );
  NAND4_X1 U14231 ( .A1(n11303), .A2(n11302), .A3(n11301), .A4(n11300), .ZN(
        n11309) );
  AOI22_X1 U14232 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n11167), .B1(
        n11047), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11307) );
  AOI22_X1 U14233 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11306) );
  AOI22_X1 U14234 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11305) );
  AOI22_X1 U14235 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11304) );
  NAND4_X1 U14236 ( .A1(n11307), .A2(n11306), .A3(n11305), .A4(n11304), .ZN(
        n11308) );
  NAND2_X1 U14237 ( .A1(n11466), .A2(n11317), .ZN(n11312) );
  INV_X1 U14238 ( .A(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11310) );
  OR2_X1 U14239 ( .A1(n11438), .A2(n11310), .ZN(n11311) );
  NAND2_X1 U14240 ( .A1(n11312), .A2(n11311), .ZN(n11326) );
  XNOR2_X1 U14241 ( .A(n11325), .B(n11326), .ZN(n12024) );
  NAND2_X1 U14242 ( .A1(n12024), .A2(n11181), .ZN(n11320) );
  NAND2_X1 U14243 ( .A1(n11314), .A2(n11313), .ZN(n11316) );
  INV_X1 U14244 ( .A(n11316), .ZN(n11318) );
  INV_X1 U14245 ( .A(n11317), .ZN(n11315) );
  OR2_X1 U14246 ( .A1(n11316), .A2(n11315), .ZN(n11367) );
  OAI211_X1 U14247 ( .C1(n11318), .C2(n11317), .A(n11391), .B(n11367), .ZN(
        n11319) );
  NAND2_X1 U14248 ( .A1(n11320), .A2(n11319), .ZN(n11322) );
  INV_X1 U14249 ( .A(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n11321) );
  XNOR2_X1 U14250 ( .A(n11322), .B(n11321), .ZN(n13819) );
  NAND2_X1 U14251 ( .A1(n13820), .A2(n13819), .ZN(n11324) );
  NAND2_X1 U14252 ( .A1(n11322), .A2(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n11323) );
  NAND2_X1 U14253 ( .A1(n11324), .A2(n11323), .ZN(n13854) );
  NAND2_X1 U14254 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(
        n11338) );
  AOI22_X1 U14255 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12458), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11330) );
  AOI22_X1 U14256 ( .A1(n12467), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12299), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11329) );
  AOI22_X1 U14257 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n11047), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11328) );
  AOI22_X1 U14258 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11327) );
  NAND4_X1 U14259 ( .A1(n11330), .A2(n11329), .A3(n11328), .A4(n11327), .ZN(
        n11336) );
  AOI22_X1 U14260 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n11334) );
  AOI22_X1 U14261 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11333) );
  AOI22_X1 U14262 ( .A1(n11167), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11332) );
  AOI22_X1 U14263 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n12468), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11331) );
  NAND4_X1 U14264 ( .A1(n11334), .A2(n11333), .A3(n11332), .A4(n11331), .ZN(
        n11335) );
  NAND2_X1 U14265 ( .A1(n11466), .A2(n11368), .ZN(n11337) );
  NAND2_X1 U14266 ( .A1(n11342), .A2(n11341), .ZN(n11343) );
  NAND2_X1 U14267 ( .A1(n11365), .A2(n11343), .ZN(n12028) );
  INV_X1 U14268 ( .A(n12028), .ZN(n11344) );
  NAND2_X1 U14269 ( .A1(n11344), .A2(n11181), .ZN(n11347) );
  XNOR2_X1 U14270 ( .A(n11367), .B(n11368), .ZN(n11345) );
  NAND2_X1 U14271 ( .A1(n11345), .A2(n11391), .ZN(n11346) );
  NAND2_X1 U14272 ( .A1(n11347), .A2(n11346), .ZN(n11349) );
  INV_X1 U14273 ( .A(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n11348) );
  XNOR2_X1 U14274 ( .A(n11349), .B(n11348), .ZN(n13853) );
  NAND2_X1 U14275 ( .A1(n13854), .A2(n13853), .ZN(n11351) );
  NAND2_X1 U14276 ( .A1(n11349), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11350) );
  NAND2_X1 U14277 ( .A1(n11351), .A2(n11350), .ZN(n15906) );
  NAND2_X1 U14278 ( .A1(n11461), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(
        n11364) );
  AOI22_X1 U14279 ( .A1(n12458), .A2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n11146), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11355) );
  AOI22_X1 U14280 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n11354) );
  AOI22_X1 U14281 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n11353) );
  AOI22_X1 U14282 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12468), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n11352) );
  NAND4_X1 U14283 ( .A1(n11355), .A2(n11354), .A3(n11353), .A4(n11352), .ZN(
        n11362) );
  AOI22_X1 U14284 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11167), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n11360) );
  AOI22_X1 U14285 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11359) );
  AOI22_X1 U14286 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11358) );
  AOI22_X1 U14287 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11357) );
  NAND4_X1 U14288 ( .A1(n11360), .A2(n11359), .A3(n11358), .A4(n11357), .ZN(
        n11361) );
  NAND2_X1 U14289 ( .A1(n11466), .A2(n11379), .ZN(n11363) );
  NAND3_X1 U14290 ( .A1(n11388), .A2(n11181), .A3(n12034), .ZN(n11372) );
  INV_X1 U14291 ( .A(n11367), .ZN(n11369) );
  NAND2_X1 U14292 ( .A1(n11369), .A2(n11368), .ZN(n11378) );
  XNOR2_X1 U14293 ( .A(n11378), .B(n11379), .ZN(n11370) );
  NAND2_X1 U14294 ( .A1(n11370), .A2(n11391), .ZN(n11371) );
  NAND2_X1 U14295 ( .A1(n11372), .A2(n11371), .ZN(n11373) );
  OR2_X1 U14296 ( .A1(n11373), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15904) );
  NAND2_X1 U14297 ( .A1(n15906), .A2(n15904), .ZN(n11374) );
  NAND2_X1 U14298 ( .A1(n11373), .A2(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n15903) );
  NAND2_X1 U14299 ( .A1(n11374), .A2(n15903), .ZN(n15898) );
  INV_X1 U14300 ( .A(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11376) );
  NAND2_X1 U14301 ( .A1(n11466), .A2(n11390), .ZN(n11375) );
  OAI21_X1 U14302 ( .B1(n11376), .B2(n11438), .A(n11375), .ZN(n11377) );
  NAND2_X1 U14303 ( .A1(n12044), .A2(n11181), .ZN(n11383) );
  INV_X1 U14304 ( .A(n11378), .ZN(n11380) );
  NAND2_X1 U14305 ( .A1(n11380), .A2(n11379), .ZN(n11389) );
  XNOR2_X1 U14306 ( .A(n11389), .B(n11390), .ZN(n11381) );
  NAND2_X1 U14307 ( .A1(n11381), .A2(n11391), .ZN(n11382) );
  NAND2_X1 U14308 ( .A1(n11383), .A2(n11382), .ZN(n15899) );
  OR2_X1 U14309 ( .A1(n15899), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11384) );
  NAND2_X1 U14310 ( .A1(n15899), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11385) );
  NOR2_X1 U14311 ( .A1(n11386), .A2(n11423), .ZN(n11387) );
  INV_X1 U14312 ( .A(n11389), .ZN(n11392) );
  NAND3_X1 U14313 ( .A1(n11392), .A2(n11391), .A3(n11390), .ZN(n11393) );
  NAND2_X1 U14314 ( .A1(n11414), .A2(n11393), .ZN(n13952) );
  AND2_X1 U14315 ( .A1(n13952), .A2(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n11395) );
  INV_X1 U14316 ( .A(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n15954) );
  OR2_X1 U14317 ( .A1(n14688), .A2(n15954), .ZN(n11396) );
  NAND2_X1 U14318 ( .A1(n11414), .A2(n15954), .ZN(n11397) );
  INV_X1 U14319 ( .A(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14827) );
  OR2_X1 U14320 ( .A1(n11414), .A2(n14827), .ZN(n14811) );
  NAND2_X1 U14321 ( .A1(n11414), .A2(n14827), .ZN(n11398) );
  NAND2_X1 U14322 ( .A1(n14811), .A2(n11398), .ZN(n14679) );
  NAND2_X1 U14323 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11399) );
  AND2_X1 U14324 ( .A1(n11414), .A2(n11399), .ZN(n14673) );
  INV_X1 U14325 ( .A(P1_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n11607) );
  INV_X1 U14326 ( .A(n14812), .ZN(n11402) );
  INV_X1 U14327 ( .A(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n11400) );
  NAND2_X1 U14328 ( .A1(n11414), .A2(n11400), .ZN(n11401) );
  NAND2_X1 U14329 ( .A1(n11402), .A2(n11401), .ZN(n14663) );
  INV_X1 U14330 ( .A(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15937) );
  NAND2_X1 U14331 ( .A1(n14688), .A2(n15937), .ZN(n11403) );
  NAND2_X1 U14332 ( .A1(n14653), .A2(n11403), .ZN(n15875) );
  INV_X1 U14333 ( .A(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n14806) );
  NOR2_X1 U14334 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n11405) );
  OR2_X1 U14335 ( .A1(n14688), .A2(n11405), .ZN(n14674) );
  OR2_X1 U14336 ( .A1(n14688), .A2(n11607), .ZN(n14675) );
  NAND2_X1 U14337 ( .A1(n14674), .A2(n14675), .ZN(n14662) );
  NOR2_X1 U14338 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n14665) );
  AND2_X1 U14339 ( .A1(n14665), .A2(n14806), .ZN(n11406) );
  NOR2_X1 U14340 ( .A1(n11414), .A2(n11406), .ZN(n15872) );
  NAND2_X1 U14341 ( .A1(n11414), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11408) );
  NAND2_X1 U14342 ( .A1(n14637), .A2(n11408), .ZN(n14645) );
  AND2_X1 U14343 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14763) );
  NOR2_X1 U14344 ( .A1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n14764) );
  INV_X1 U14345 ( .A(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n11565) );
  INV_X1 U14346 ( .A(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n11410) );
  NAND3_X1 U14347 ( .A1(n14764), .A2(n11565), .A3(n11410), .ZN(n11411) );
  INV_X1 U14348 ( .A(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n14727) );
  INV_X1 U14349 ( .A(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14739) );
  NAND2_X1 U14350 ( .A1(n14727), .A2(n14739), .ZN(n11412) );
  AND2_X1 U14351 ( .A1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n14728) );
  NAND2_X1 U14352 ( .A1(n14728), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14601) );
  INV_X1 U14353 ( .A(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14581) );
  INV_X1 U14354 ( .A(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n14718) );
  NAND2_X1 U14355 ( .A1(n14581), .A2(n14718), .ZN(n14710) );
  INV_X1 U14356 ( .A(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n14698) );
  NAND2_X1 U14357 ( .A1(n14297), .A2(n14698), .ZN(n12521) );
  AND2_X1 U14358 ( .A1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n14699) );
  NAND2_X1 U14359 ( .A1(n12521), .A2(n12522), .ZN(n11416) );
  XNOR2_X1 U14360 ( .A(n11416), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14574) );
  MUX2_X1 U14361 ( .A(n20440), .B(P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .Z(n11435) );
  NAND2_X1 U14362 ( .A1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n20551), .ZN(
        n11424) );
  NAND2_X1 U14363 ( .A1(n11435), .A2(n11434), .ZN(n11418) );
  NAND2_X1 U14364 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n20440), .ZN(
        n11417) );
  NAND2_X1 U14365 ( .A1(n11418), .A2(n11417), .ZN(n11445) );
  NAND2_X1 U14366 ( .A1(n20514), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n11420) );
  NAND2_X1 U14367 ( .A1(n11235), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n11419) );
  NAND2_X1 U14368 ( .A1(n11445), .A2(n11444), .ZN(n11443) );
  NAND2_X1 U14369 ( .A1(n11443), .A2(n11420), .ZN(n11452) );
  MUX2_X1 U14370 ( .A(n20184), .B(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n11453) );
  INV_X1 U14371 ( .A(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n20100) );
  NOR2_X1 U14372 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n20100), .ZN(
        n11422) );
  NOR2_X1 U14373 ( .A1(n11438), .A2(n11423), .ZN(n11467) );
  INV_X1 U14374 ( .A(n11467), .ZN(n11427) );
  OAI21_X1 U14375 ( .B1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20551), .A(
        n11424), .ZN(n11425) );
  INV_X1 U14376 ( .A(n11425), .ZN(n11431) );
  NAND2_X1 U14377 ( .A1(n11466), .A2(n11431), .ZN(n11426) );
  NAND2_X1 U14378 ( .A1(n11427), .A2(n11426), .ZN(n11433) );
  AOI21_X1 U14379 ( .B1(n11428), .B2(n11501), .A(n20122), .ZN(n11455) );
  INV_X1 U14380 ( .A(n11455), .ZN(n11430) );
  NAND2_X1 U14381 ( .A1(n13267), .A2(n11501), .ZN(n11429) );
  NAND3_X1 U14382 ( .A1(n11431), .A2(n11430), .A3(n11429), .ZN(n11432) );
  XNOR2_X1 U14383 ( .A(n11435), .B(n11434), .ZN(n11477) );
  INV_X1 U14384 ( .A(n11477), .ZN(n11440) );
  NAND2_X1 U14385 ( .A1(n11466), .A2(n20122), .ZN(n11437) );
  NOR2_X1 U14386 ( .A1(n11180), .A2(n11192), .ZN(n11439) );
  INV_X1 U14387 ( .A(n11439), .ZN(n11436) );
  OAI211_X1 U14388 ( .C1(n11438), .C2(n11440), .A(n11437), .B(n11436), .ZN(
        n11441) );
  NOR3_X1 U14389 ( .A1(n11466), .A2(n11439), .A3(n13281), .ZN(n11451) );
  OAI22_X1 U14390 ( .A1(n11442), .A2(n11441), .B1(n11451), .B2(n11440), .ZN(
        n11449) );
  NAND2_X1 U14391 ( .A1(n11442), .A2(n11441), .ZN(n11448) );
  OAI21_X1 U14392 ( .B1(n11445), .B2(n11444), .A(n11443), .ZN(n11478) );
  INV_X1 U14393 ( .A(n11466), .ZN(n11446) );
  NOR2_X1 U14394 ( .A1(n11446), .A2(n11478), .ZN(n11456) );
  AOI211_X1 U14395 ( .C1(n11461), .C2(n11478), .A(n11455), .B(n11456), .ZN(
        n11447) );
  AOI21_X1 U14396 ( .B1(n11449), .B2(n11448), .A(n11447), .ZN(n11463) );
  NAND3_X1 U14397 ( .A1(P1_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n11450), .A3(
        n13690), .ZN(n11460) );
  INV_X1 U14398 ( .A(n11451), .ZN(n11458) );
  XOR2_X1 U14399 ( .A(n11453), .B(n11452), .Z(n11459) );
  INV_X1 U14400 ( .A(n11459), .ZN(n11454) );
  AOI22_X1 U14401 ( .A1(n11456), .A2(n11455), .B1(n11181), .B2(n11454), .ZN(
        n11457) );
  OAI21_X1 U14402 ( .B1(n11460), .B2(n11458), .A(n11457), .ZN(n11462) );
  OAI22_X1 U14403 ( .A1(n11463), .A2(n11462), .B1(n11461), .B2(n11480), .ZN(
        n11464) );
  OAI21_X1 U14404 ( .B1(P1_STATE2_REG_0__SCAN_IN), .B2(n13690), .A(n11464), 
        .ZN(n11465) );
  INV_X1 U14405 ( .A(n14280), .ZN(n12172) );
  NAND2_X1 U14406 ( .A1(n12172), .A2(n20122), .ZN(n11485) );
  INV_X1 U14407 ( .A(n11470), .ZN(n13272) );
  NAND2_X1 U14408 ( .A1(n13486), .A2(n11501), .ZN(n11471) );
  NAND2_X1 U14409 ( .A1(n11471), .A2(n20793), .ZN(n11472) );
  NAND2_X1 U14410 ( .A1(n11473), .A2(n11472), .ZN(n11609) );
  INV_X1 U14411 ( .A(n11600), .ZN(n11474) );
  AOI21_X1 U14412 ( .B1(n14280), .B2(n12498), .A(n11474), .ZN(n11475) );
  NAND2_X1 U14413 ( .A1(n11609), .A2(n13271), .ZN(n11476) );
  NAND2_X1 U14414 ( .A1(n13272), .A2(n11476), .ZN(n13473) );
  NOR2_X1 U14415 ( .A1(n11478), .A2(n11477), .ZN(n11481) );
  AOI21_X1 U14416 ( .B1(n11481), .B2(n11480), .A(n11479), .ZN(n13472) );
  NAND2_X1 U14417 ( .A1(READY1), .A2(READY11_REG_SCAN_IN), .ZN(n15993) );
  INV_X1 U14418 ( .A(P1_STATE_REG_0__SCAN_IN), .ZN(n20699) );
  NAND2_X1 U14419 ( .A1(n11482), .A2(n20699), .ZN(n15736) );
  NAND2_X1 U14420 ( .A1(n20122), .A2(n15736), .ZN(n11483) );
  NAND4_X1 U14421 ( .A1(n13472), .A2(n11108), .A3(n15993), .A4(n11483), .ZN(
        n11484) );
  OAI211_X1 U14422 ( .C1(n13698), .C2(n11485), .A(n13473), .B(n11484), .ZN(
        n11486) );
  NOR2_X1 U14423 ( .A1(n20689), .A2(n11192), .ZN(n13520) );
  NAND2_X1 U14424 ( .A1(n11486), .A2(n13520), .ZN(n11493) );
  INV_X1 U14425 ( .A(n15736), .ZN(n13513) );
  OR2_X1 U14426 ( .A1(n20122), .A2(n13513), .ZN(n12502) );
  NAND2_X1 U14427 ( .A1(n12502), .A2(n15993), .ZN(n11489) );
  OAI211_X1 U14428 ( .C1(n11487), .C2(n11489), .A(n11501), .B(n11488), .ZN(
        n11490) );
  NAND3_X1 U14429 ( .A1(n13621), .A2(n11491), .A3(n11490), .ZN(n11492) );
  AND2_X1 U14430 ( .A1(n13271), .A2(n13267), .ZN(n15709) );
  INV_X1 U14431 ( .A(n15709), .ZN(n11496) );
  NAND2_X1 U14432 ( .A1(n13271), .A2(n13265), .ZN(n13657) );
  INV_X1 U14433 ( .A(n11597), .ZN(n11494) );
  NAND2_X1 U14434 ( .A1(n11494), .A2(n11127), .ZN(n11495) );
  NAND4_X1 U14435 ( .A1(n11497), .A2(n11496), .A3(n13657), .A4(n11495), .ZN(
        n11498) );
  INV_X1 U14436 ( .A(n20129), .ZN(n11499) );
  NAND2_X1 U14437 ( .A1(n11499), .A2(n11501), .ZN(n11514) );
  INV_X1 U14438 ( .A(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n20087) );
  INV_X1 U14439 ( .A(P1_EBX_REG_0__SCAN_IN), .ZN(n11502) );
  OR2_X1 U14440 ( .A1(n11514), .A2(n11502), .ZN(n11504) );
  NAND2_X1 U14441 ( .A1(n11500), .A2(n11502), .ZN(n11503) );
  NAND2_X1 U14442 ( .A1(n11504), .A2(n11503), .ZN(n13523) );
  MUX2_X1 U14443 ( .A(n11586), .B(n12493), .S(P1_EBX_REG_2__SCAN_IN), .Z(
        n11506) );
  NAND2_X1 U14444 ( .A1(n20069), .A2(n13522), .ZN(n11505) );
  NAND2_X1 U14445 ( .A1(n13652), .A2(n13651), .ZN(n13713) );
  INV_X1 U14446 ( .A(P1_EBX_REG_3__SCAN_IN), .ZN(n19935) );
  NAND2_X1 U14447 ( .A1(n11576), .A2(n19935), .ZN(n11510) );
  NAND2_X1 U14448 ( .A1(n11514), .A2(n13756), .ZN(n11508) );
  NAND2_X1 U14449 ( .A1(n11588), .A2(n19935), .ZN(n11507) );
  NAND3_X1 U14450 ( .A1(n11508), .A2(n12493), .A3(n11507), .ZN(n11509) );
  INV_X1 U14451 ( .A(P1_EBX_REG_4__SCAN_IN), .ZN(n19924) );
  NAND2_X1 U14452 ( .A1(n11581), .A2(n19924), .ZN(n11513) );
  NAND2_X1 U14453 ( .A1(n11588), .A2(n19924), .ZN(n11511) );
  OAI211_X1 U14454 ( .C1(n11500), .C2(n11321), .A(n11511), .B(n11514), .ZN(
        n11512) );
  NAND2_X1 U14455 ( .A1(n11513), .A2(n11512), .ZN(n13779) );
  MUX2_X1 U14456 ( .A(n11591), .B(n11514), .S(P1_EBX_REG_5__SCAN_IN), .Z(
        n11518) );
  INV_X1 U14457 ( .A(n11514), .ZN(n11515) );
  NAND2_X1 U14458 ( .A1(n11515), .A2(n13516), .ZN(n11558) );
  NAND2_X1 U14459 ( .A1(n13516), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n11516) );
  AND2_X1 U14460 ( .A1(n11558), .A2(n11516), .ZN(n11517) );
  NAND2_X1 U14461 ( .A1(n11518), .A2(n11517), .ZN(n13814) );
  INV_X1 U14462 ( .A(P1_EBX_REG_6__SCAN_IN), .ZN(n19967) );
  NAND2_X1 U14463 ( .A1(n11581), .A2(n19967), .ZN(n11521) );
  INV_X1 U14464 ( .A(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n15974) );
  NAND2_X1 U14465 ( .A1(n11588), .A2(n19967), .ZN(n11519) );
  OAI211_X1 U14466 ( .C1(n11500), .C2(n15974), .A(n11519), .B(n11514), .ZN(
        n11520) );
  NAND2_X1 U14467 ( .A1(n15983), .A2(n15982), .ZN(n15985) );
  MUX2_X1 U14468 ( .A(n11591), .B(n11514), .S(P1_EBX_REG_7__SCAN_IN), .Z(
        n11523) );
  NAND2_X1 U14469 ( .A1(n13516), .A2(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n11522) );
  INV_X1 U14470 ( .A(P1_EBX_REG_8__SCAN_IN), .ZN(n14421) );
  NAND2_X1 U14471 ( .A1(n11581), .A2(n14421), .ZN(n11528) );
  INV_X1 U14472 ( .A(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n15973) );
  NAND2_X1 U14473 ( .A1(n11588), .A2(n14421), .ZN(n11526) );
  OAI211_X1 U14474 ( .C1(n11500), .C2(n15973), .A(n11526), .B(n11514), .ZN(
        n11527) );
  NAND2_X1 U14475 ( .A1(n11528), .A2(n11527), .ZN(n13901) );
  MUX2_X1 U14476 ( .A(n11591), .B(n11514), .S(P1_EBX_REG_9__SCAN_IN), .Z(
        n11530) );
  NAND2_X1 U14477 ( .A1(n13516), .A2(P1_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n11529) );
  MUX2_X1 U14478 ( .A(n11586), .B(n12493), .S(P1_EBX_REG_10__SCAN_IN), .Z(
        n11532) );
  INV_X1 U14479 ( .A(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15960) );
  NAND2_X1 U14480 ( .A1(n13522), .A2(n15960), .ZN(n11531) );
  INV_X1 U14481 ( .A(P1_EBX_REG_12__SCAN_IN), .ZN(n15858) );
  NAND2_X1 U14482 ( .A1(n11581), .A2(n15858), .ZN(n11535) );
  NAND2_X1 U14483 ( .A1(n11588), .A2(n15858), .ZN(n11533) );
  OAI211_X1 U14484 ( .C1(n11500), .C2(n11607), .A(n11533), .B(n11514), .ZN(
        n11534) );
  MUX2_X1 U14485 ( .A(n11591), .B(n11514), .S(P1_EBX_REG_11__SCAN_IN), .Z(
        n11538) );
  NAND2_X1 U14486 ( .A1(n13516), .A2(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(
        n11536) );
  AND2_X1 U14487 ( .A1(n11558), .A2(n11536), .ZN(n11537) );
  NAND2_X1 U14488 ( .A1(n11538), .A2(n11537), .ZN(n14839) );
  NAND2_X1 U14489 ( .A1(n14838), .A2(n14839), .ZN(n11539) );
  INV_X1 U14490 ( .A(P1_EBX_REG_13__SCAN_IN), .ZN(n14188) );
  NAND2_X1 U14491 ( .A1(n11576), .A2(n14188), .ZN(n11543) );
  NAND2_X1 U14492 ( .A1(n11514), .A2(n14827), .ZN(n11541) );
  NAND2_X1 U14493 ( .A1(n11588), .A2(n14188), .ZN(n11540) );
  NAND3_X1 U14494 ( .A1(n11541), .A2(n12493), .A3(n11540), .ZN(n11542) );
  MUX2_X1 U14495 ( .A(n11586), .B(n12493), .S(P1_EBX_REG_14__SCAN_IN), .Z(
        n11545) );
  NAND2_X1 U14496 ( .A1(n13522), .A2(n11400), .ZN(n11544) );
  MUX2_X1 U14497 ( .A(n11591), .B(n11514), .S(P1_EBX_REG_15__SCAN_IN), .Z(
        n11548) );
  NAND2_X1 U14498 ( .A1(n13516), .A2(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n11546) );
  AND2_X1 U14499 ( .A1(n11558), .A2(n11546), .ZN(n11547) );
  NAND2_X1 U14500 ( .A1(n11548), .A2(n11547), .ZN(n14151) );
  MUX2_X1 U14501 ( .A(n11586), .B(n12493), .S(P1_EBX_REG_16__SCAN_IN), .Z(
        n11549) );
  OAI21_X1 U14502 ( .B1(P1_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n12495), .A(
        n11549), .ZN(n14169) );
  INV_X1 U14503 ( .A(P1_EBX_REG_17__SCAN_IN), .ZN(n15811) );
  NAND2_X1 U14504 ( .A1(n11576), .A2(n15811), .ZN(n11554) );
  INV_X1 U14505 ( .A(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n11550) );
  NAND2_X1 U14506 ( .A1(n11514), .A2(n11550), .ZN(n11552) );
  NAND2_X1 U14507 ( .A1(n11588), .A2(n15811), .ZN(n11551) );
  NAND3_X1 U14508 ( .A1(n11552), .A2(n12493), .A3(n11551), .ZN(n11553) );
  MUX2_X1 U14509 ( .A(n11581), .B(n11500), .S(P1_EBX_REG_18__SCAN_IN), .Z(
        n11556) );
  NOR2_X1 U14510 ( .A1(n12495), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n11555) );
  NOR2_X1 U14511 ( .A1(n11556), .A2(n11555), .ZN(n14392) );
  MUX2_X1 U14512 ( .A(n11591), .B(n11514), .S(P1_EBX_REG_19__SCAN_IN), .Z(
        n11560) );
  NAND2_X1 U14513 ( .A1(n13516), .A2(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n11557) );
  AND2_X1 U14514 ( .A1(n11558), .A2(n11557), .ZN(n11559) );
  NAND2_X1 U14515 ( .A1(n11560), .A2(n11559), .ZN(n14381) );
  NAND2_X1 U14516 ( .A1(n14390), .A2(n14381), .ZN(n14759) );
  INV_X1 U14517 ( .A(P1_EBX_REG_20__SCAN_IN), .ZN(n15854) );
  NAND2_X1 U14518 ( .A1(n11581), .A2(n15854), .ZN(n11564) );
  INV_X1 U14519 ( .A(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n11562) );
  NAND2_X1 U14520 ( .A1(n11588), .A2(n15854), .ZN(n11561) );
  OAI211_X1 U14521 ( .C1(n11500), .C2(n11562), .A(n11561), .B(n11514), .ZN(
        n11563) );
  NAND2_X1 U14522 ( .A1(n11564), .A2(n11563), .ZN(n14758) );
  INV_X1 U14523 ( .A(P1_EBX_REG_21__SCAN_IN), .ZN(n11566) );
  NAND2_X1 U14524 ( .A1(n11576), .A2(n11566), .ZN(n11570) );
  NAND2_X1 U14525 ( .A1(n11514), .A2(n11565), .ZN(n11568) );
  NAND2_X1 U14526 ( .A1(n11588), .A2(n11566), .ZN(n11567) );
  NAND3_X1 U14527 ( .A1(n11568), .A2(n12493), .A3(n11567), .ZN(n11569) );
  AND2_X1 U14528 ( .A1(n11570), .A2(n11569), .ZN(n14489) );
  MUX2_X1 U14529 ( .A(n11586), .B(n12493), .S(P1_EBX_REG_22__SCAN_IN), .Z(
        n11571) );
  OAI21_X1 U14530 ( .B1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n12495), .A(
        n11571), .ZN(n14482) );
  NAND2_X1 U14531 ( .A1(n11514), .A2(n10173), .ZN(n11573) );
  INV_X1 U14532 ( .A(P1_EBX_REG_23__SCAN_IN), .ZN(n14475) );
  NAND2_X1 U14533 ( .A1(n11588), .A2(n14475), .ZN(n11572) );
  NAND3_X1 U14534 ( .A1(n11573), .A2(n12493), .A3(n11572), .ZN(n11574) );
  OAI21_X1 U14535 ( .B1(n11591), .B2(P1_EBX_REG_23__SCAN_IN), .A(n11574), .ZN(
        n14472) );
  MUX2_X1 U14536 ( .A(n11586), .B(n12493), .S(P1_EBX_REG_24__SCAN_IN), .Z(
        n11575) );
  OAI21_X1 U14537 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n12495), .A(
        n11575), .ZN(n14466) );
  INV_X1 U14538 ( .A(P1_EBX_REG_25__SCAN_IN), .ZN(n15749) );
  NAND2_X1 U14539 ( .A1(n11576), .A2(n15749), .ZN(n11580) );
  NAND2_X1 U14540 ( .A1(n11514), .A2(n14727), .ZN(n11578) );
  NAND2_X1 U14541 ( .A1(n11588), .A2(n15749), .ZN(n11577) );
  NAND3_X1 U14542 ( .A1(n11578), .A2(n12493), .A3(n11577), .ZN(n11579) );
  AND2_X1 U14543 ( .A1(n11580), .A2(n11579), .ZN(n14457) );
  MUX2_X1 U14544 ( .A(n11581), .B(n11500), .S(P1_EBX_REG_26__SCAN_IN), .Z(
        n11583) );
  NOR2_X1 U14545 ( .A1(n12495), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n11582) );
  NOR2_X1 U14546 ( .A1(n11583), .A2(n11582), .ZN(n14361) );
  NAND2_X1 U14547 ( .A1(n11514), .A2(n14718), .ZN(n11584) );
  OAI211_X1 U14548 ( .C1(P1_EBX_REG_27__SCAN_IN), .C2(n13516), .A(n11584), .B(
        n12493), .ZN(n11585) );
  OAI21_X1 U14549 ( .B1(n11591), .B2(P1_EBX_REG_27__SCAN_IN), .A(n11585), .ZN(
        n14349) );
  MUX2_X1 U14550 ( .A(n11586), .B(n12493), .S(P1_EBX_REG_28__SCAN_IN), .Z(
        n11587) );
  OAI21_X1 U14551 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n12495), .A(
        n11587), .ZN(n14334) );
  OR2_X1 U14552 ( .A1(n12495), .A2(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n11590) );
  INV_X1 U14553 ( .A(P1_EBX_REG_29__SCAN_IN), .ZN(n14319) );
  NAND2_X1 U14554 ( .A1(n11588), .A2(n14319), .ZN(n11589) );
  NAND2_X1 U14555 ( .A1(n11590), .A2(n11589), .ZN(n11593) );
  OAI22_X1 U14556 ( .A1(n11593), .A2(n11500), .B1(P1_EBX_REG_29__SCAN_IN), 
        .B2(n11591), .ZN(n14311) );
  NAND2_X1 U14557 ( .A1(n14336), .A2(n14311), .ZN(n14310) );
  NAND2_X1 U14558 ( .A1(n14310), .A2(n11500), .ZN(n11594) );
  INV_X1 U14559 ( .A(n14336), .ZN(n11592) );
  AND2_X1 U14560 ( .A1(n13516), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n11595) );
  AOI21_X1 U14561 ( .B1(n12495), .B2(P1_EBX_REG_30__SCAN_IN), .A(n11595), .ZN(
        n12494) );
  NOR2_X1 U14562 ( .A1(n11597), .A2(n11127), .ZN(n11598) );
  AOI21_X1 U14563 ( .B1(n11596), .B2(n13281), .A(n11598), .ZN(n11599) );
  NOR2_X2 U14564 ( .A1(n11620), .A2(n11599), .ZN(n20089) );
  NAND2_X1 U14565 ( .A1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n15936) );
  NOR3_X1 U14566 ( .A1(n11400), .A2(n11550), .A3(n15936), .ZN(n14789) );
  AND2_X1 U14567 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n14789), .ZN(
        n11619) );
  OR2_X1 U14568 ( .A1(n13522), .A2(n11600), .ZN(n13457) );
  OR2_X1 U14569 ( .A1(n13267), .A2(n14432), .ZN(n13456) );
  AND2_X1 U14570 ( .A1(n13456), .A2(n11601), .ZN(n11602) );
  NAND2_X1 U14571 ( .A1(n13457), .A2(n11602), .ZN(n11611) );
  INV_X1 U14572 ( .A(n13658), .ZN(n11604) );
  AOI21_X1 U14573 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n20064) );
  NAND2_X1 U14574 ( .A1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n20056) );
  NOR2_X1 U14575 ( .A1(n11348), .A2(n20056), .ZN(n14006) );
  INV_X1 U14576 ( .A(n14006), .ZN(n11605) );
  NOR2_X1 U14577 ( .A1(n20064), .A2(n11605), .ZN(n14008) );
  INV_X1 U14578 ( .A(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15980) );
  NOR3_X1 U14579 ( .A1(n15973), .A2(n15980), .A3(n15974), .ZN(n14009) );
  NOR2_X1 U14580 ( .A1(n15960), .A2(n15954), .ZN(n15953) );
  AND2_X1 U14581 ( .A1(n14009), .A2(n15953), .ZN(n11606) );
  NAND3_X1 U14582 ( .A1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n14008), .A3(
        n11606), .ZN(n14846) );
  NOR2_X1 U14583 ( .A1(n11607), .A2(n14846), .ZN(n11617) );
  INV_X1 U14584 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n14848) );
  NAND4_X1 U14585 ( .A1(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n14006), .A4(n11606), .ZN(
        n14844) );
  NOR3_X1 U14586 ( .A1(n11607), .A2(n14848), .A3(n14844), .ZN(n11618) );
  AND2_X1 U14587 ( .A1(n11470), .A2(n20122), .ZN(n15697) );
  NAND2_X1 U14588 ( .A1(n11613), .A2(n15697), .ZN(n20099) );
  NAND3_X1 U14589 ( .A1(n11610), .A2(n9918), .A3(n11609), .ZN(n13459) );
  OR2_X1 U14590 ( .A1(n13459), .A2(n11611), .ZN(n11612) );
  NAND2_X1 U14591 ( .A1(n11613), .A2(n11612), .ZN(n11621) );
  NAND2_X1 U14592 ( .A1(n20099), .A2(n11621), .ZN(n14845) );
  AOI22_X1 U14593 ( .A1(n20062), .A2(n11617), .B1(n11618), .B2(n20070), .ZN(
        n14828) );
  NOR2_X1 U14594 ( .A1(n14828), .A2(n14827), .ZN(n14784) );
  NAND2_X1 U14595 ( .A1(n11619), .A2(n14784), .ZN(n14779) );
  INV_X1 U14596 ( .A(n14763), .ZN(n11614) );
  NOR2_X1 U14597 ( .A1(n14779), .A2(n11614), .ZN(n15930) );
  AND2_X1 U14598 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n11615) );
  NAND2_X1 U14599 ( .A1(n15922), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n14697) );
  INV_X1 U14600 ( .A(n14699), .ZN(n14709) );
  OR3_X1 U14601 ( .A1(n14697), .A2(n14709), .A3(n14698), .ZN(n12528) );
  NAND2_X1 U14602 ( .A1(n11621), .A2(n14786), .ZN(n20075) );
  INV_X1 U14603 ( .A(n20075), .ZN(n11616) );
  NAND2_X1 U14604 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n15929) );
  AND2_X1 U14605 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n11617), .ZN(
        n14820) );
  AOI21_X1 U14606 ( .B1(n14820), .B2(n11619), .A(n14786), .ZN(n11623) );
  AND2_X1 U14607 ( .A1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n11618), .ZN(
        n14785) );
  AOI21_X1 U14608 ( .B1(n11619), .B2(n14785), .A(n20066), .ZN(n11622) );
  NAND2_X1 U14609 ( .A1(n11620), .A2(n20046), .ZN(n20098) );
  OAI21_X1 U14610 ( .B1(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(n11621), .A(
        n20098), .ZN(n14788) );
  NOR3_X1 U14611 ( .A1(n11623), .A2(n11622), .A3(n14788), .ZN(n14777) );
  INV_X1 U14612 ( .A(n14788), .ZN(n20065) );
  AOI22_X1 U14613 ( .A1(n14763), .A2(n14777), .B1(n14790), .B2(n20065), .ZN(
        n15926) );
  AOI21_X1 U14614 ( .B1(n20076), .B2(n15929), .A(n15926), .ZN(n14746) );
  OAI21_X1 U14615 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n14786), .A(
        n14746), .ZN(n14736) );
  OAI22_X1 U14616 ( .A1(n20066), .A2(n14728), .B1(
        P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14786), .ZN(n11624) );
  NOR2_X1 U14617 ( .A1(n14736), .A2(n11624), .ZN(n14726) );
  NAND2_X1 U14618 ( .A1(n14726), .A2(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15920) );
  INV_X1 U14619 ( .A(n15920), .ZN(n11625) );
  NAND2_X1 U14620 ( .A1(n11625), .A2(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14708) );
  NAND2_X1 U14621 ( .A1(n14726), .A2(n14790), .ZN(n14707) );
  OAI21_X1 U14622 ( .B1(n14708), .B2(n14709), .A(n14707), .ZN(n14696) );
  OAI211_X1 U14623 ( .C1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .C2(n14790), .A(
        n14696), .B(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12525) );
  INV_X1 U14624 ( .A(n12525), .ZN(n11626) );
  AOI21_X1 U14625 ( .B1(n9939), .B2(n12528), .A(n11626), .ZN(n11627) );
  INV_X1 U14626 ( .A(P1_REIP_REG_30__SCAN_IN), .ZN(n14324) );
  NOR2_X1 U14627 ( .A1(n20046), .A2(n14324), .ZN(n14568) );
  AOI21_X1 U14628 ( .B1(n14320), .B2(n20089), .A(n10300), .ZN(n11628) );
  OAI21_X1 U14629 ( .B1(n14574), .B2(n20095), .A(n11628), .ZN(P1_U3001) );
  INV_X1 U14630 ( .A(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16469) );
  INV_X1 U14631 ( .A(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n17389) );
  NAND3_X1 U14632 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17694) );
  INV_X1 U14633 ( .A(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n16607) );
  INV_X1 U14634 ( .A(n17409), .ZN(n17438) );
  INV_X1 U14635 ( .A(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n17410) );
  NAND2_X1 U14636 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17412) );
  INV_X1 U14637 ( .A(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n16479) );
  XNOR2_X1 U14638 ( .A(n16469), .B(n11635), .ZN(n16468) );
  AOI21_X1 U14639 ( .B1(n16479), .B2(n16307), .A(n11635), .ZN(n16478) );
  OAI21_X1 U14640 ( .B1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .B2(n11638), .A(
        n16307), .ZN(n17371) );
  INV_X1 U14641 ( .A(n17371), .ZN(n16492) );
  INV_X1 U14642 ( .A(P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17414) );
  NAND2_X1 U14643 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n11633), .ZN(
        n11631) );
  AOI21_X1 U14644 ( .B1(n17414), .B2(n11631), .A(n17366), .ZN(n17416) );
  INV_X1 U14645 ( .A(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n17424) );
  AOI22_X1 U14646 ( .A1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n11633), .B1(
        n11632), .B2(n17424), .ZN(n17431) );
  AOI21_X1 U14647 ( .B1(n17410), .B2(n17438), .A(n11633), .ZN(n17439) );
  INV_X1 U14648 ( .A(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n17465) );
  NAND2_X1 U14649 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(n17495), .ZN(
        n16601) );
  INV_X1 U14650 ( .A(n16601), .ZN(n17493) );
  NAND3_X1 U14651 ( .A1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A3(n17493), .ZN(n17449) );
  NOR2_X1 U14652 ( .A1(n21050), .A2(n17449), .ZN(n11637) );
  NAND2_X1 U14653 ( .A1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .A2(n11637), .ZN(
        n11634) );
  AOI21_X1 U14654 ( .B1(n17465), .B2(n11634), .A(n17409), .ZN(n17455) );
  XOR2_X1 U14655 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n11637), .Z(
        n17470) );
  INV_X1 U14656 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n16310) );
  NAND2_X1 U14657 ( .A1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n11635), .ZN(
        n11636) );
  XOR2_X2 U14658 ( .A(n16310), .B(n11636), .Z(n16797) );
  OR2_X1 U14659 ( .A1(n17745), .A2(n17664), .ZN(n16731) );
  NOR2_X1 U14660 ( .A1(n17665), .A2(n16731), .ZN(n16718) );
  NAND2_X1 U14661 ( .A1(n17559), .A2(n16718), .ZN(n17571) );
  OR2_X1 U14662 ( .A1(n17583), .A2(n17571), .ZN(n16646) );
  NOR2_X1 U14663 ( .A1(n17561), .A2(n16646), .ZN(n17534) );
  NAND2_X1 U14664 ( .A1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n17534), .ZN(
        n16627) );
  NOR2_X1 U14665 ( .A1(n16627), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16593) );
  AOI21_X1 U14666 ( .B1(n21050), .B2(n17449), .A(n11637), .ZN(n17487) );
  NOR2_X1 U14667 ( .A1(n17470), .A2(n16558), .ZN(n16557) );
  NOR2_X1 U14668 ( .A1(n16557), .A2(n16770), .ZN(n16550) );
  NOR2_X1 U14669 ( .A1(n17455), .A2(n16550), .ZN(n16549) );
  NOR2_X1 U14670 ( .A1(n16549), .A2(n16770), .ZN(n16535) );
  NOR2_X1 U14671 ( .A1(n17439), .A2(n16535), .ZN(n16534) );
  NOR2_X1 U14672 ( .A1(n16534), .A2(n16770), .ZN(n16528) );
  NOR2_X1 U14673 ( .A1(n17431), .A2(n16528), .ZN(n16527) );
  NOR2_X1 U14674 ( .A1(n16527), .A2(n16770), .ZN(n16515) );
  OAI21_X1 U14675 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17366), .A(
        n9876), .ZN(n17399) );
  AOI21_X1 U14676 ( .B1(n16514), .B2(n17399), .A(n16770), .ZN(n16499) );
  AOI21_X1 U14677 ( .B1(n17389), .B2(n9876), .A(n11638), .ZN(n17384) );
  NOR2_X1 U14678 ( .A1(n16490), .A2(n16770), .ZN(n16477) );
  NOR2_X1 U14679 ( .A1(n16478), .A2(n16477), .ZN(n16476) );
  NOR2_X1 U14680 ( .A1(n16476), .A2(n16770), .ZN(n16467) );
  NAND4_X1 U14681 ( .A1(n18603), .A2(n18604), .A3(n18745), .A4(
        P3_STATE2_REG_1__SCAN_IN), .ZN(n18602) );
  INV_X1 U14682 ( .A(n18602), .ZN(n16788) );
  NAND2_X1 U14683 ( .A1(n16797), .A2(n16788), .ZN(n16799) );
  NOR3_X1 U14684 ( .A1(n16468), .A2(n16467), .A3(n16799), .ZN(n11771) );
  INV_X1 U14685 ( .A(P3_REIP_REG_27__SCAN_IN), .ZN(n18675) );
  NAND2_X2 U14686 ( .A1(n18720), .A2(n18727), .ZN(n16793) );
  OR2_X2 U14687 ( .A1(n11646), .A2(n16793), .ZN(n15611) );
  INV_X2 U14688 ( .A(n15611), .ZN(n17035) );
  AOI22_X1 U14689 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n9845), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n11644) );
  AOI22_X1 U14690 ( .A1(n17024), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11825), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n11643) );
  AOI22_X1 U14691 ( .A1(n15609), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(n17034), .ZN(n11642) );
  INV_X4 U14692 ( .A(n15599), .ZN(n15640) );
  AOI22_X1 U14693 ( .A1(n9815), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11641) );
  NAND4_X1 U14694 ( .A1(n11644), .A2(n11643), .A3(n11642), .A4(n11641), .ZN(
        n11655) );
  AOI22_X1 U14696 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n17069), .B2(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n11653) );
  AOI22_X1 U14697 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n9818), .B2(P3_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n11652) );
  AOI22_X1 U14698 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(n9841), .B2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n11651) );
  AOI22_X1 U14699 ( .A1(n9809), .A2(P3_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11827), .B2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n11650) );
  NAND4_X1 U14700 ( .A1(n11653), .A2(n11652), .A3(n11651), .A4(n11650), .ZN(
        n11654) );
  INV_X1 U14701 ( .A(P3_STATE_REG_0__SCAN_IN), .ZN(n18623) );
  NOR2_X2 U14702 ( .A1(n20880), .A2(P3_STATE_REG_0__SCAN_IN), .ZN(n18682) );
  NAND2_X2 U14703 ( .A1(n18682), .A2(P3_STATE_REG_2__SCAN_IN), .ZN(n18680) );
  NOR2_X1 U14704 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(P3_STATE_REG_2__SCAN_IN), 
        .ZN(n18609) );
  INV_X1 U14705 ( .A(n18609), .ZN(n11656) );
  NAND3_X1 U14706 ( .A1(n18623), .A2(n18680), .A3(n11656), .ZN(n18744) );
  NAND2_X1 U14707 ( .A1(READY2), .A2(READY22_REG_SCAN_IN), .ZN(n18747) );
  INV_X1 U14708 ( .A(n18747), .ZN(n18615) );
  AOI211_X1 U14709 ( .C1(n18100), .C2(n18744), .A(n18615), .B(
        P3_STATEBS16_REG_SCAN_IN), .ZN(n11761) );
  INV_X1 U14710 ( .A(n11761), .ZN(n18588) );
  AOI22_X1 U14711 ( .A1(n9815), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11666) );
  AOI22_X1 U14712 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(n9841), .B2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n11665) );
  INV_X1 U14713 ( .A(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n18098) );
  AOI22_X1 U14714 ( .A1(n9838), .A2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n17024), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n11657) );
  OAI21_X1 U14715 ( .B1(n17006), .B2(n18098), .A(n11657), .ZN(n11664) );
  AOI22_X1 U14716 ( .A1(n11825), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11662) );
  AOI22_X1 U14717 ( .A1(n9810), .A2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n11827), .B2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n11661) );
  AOI22_X1 U14718 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(n9845), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n11660) );
  AOI22_X1 U14719 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9842), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11659) );
  NAND4_X1 U14720 ( .A1(n11662), .A2(n11661), .A3(n11660), .A4(n11659), .ZN(
        n11663) );
  AOI22_X1 U14721 ( .A1(n9811), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11676) );
  AOI22_X1 U14722 ( .A1(n9809), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17024), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11675) );
  INV_X1 U14723 ( .A(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n18110) );
  AOI22_X1 U14724 ( .A1(n9845), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(n9842), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11667) );
  OAI21_X1 U14725 ( .B1(n17006), .B2(n18110), .A(n11667), .ZN(n11673) );
  AOI22_X1 U14726 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n9830), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n11671) );
  AOI22_X1 U14727 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(n9822), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11670) );
  AOI22_X1 U14728 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9816), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n11669) );
  AOI22_X1 U14729 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n11668) );
  NAND4_X1 U14730 ( .A1(n11671), .A2(n11670), .A3(n11669), .A4(n11668), .ZN(
        n11672) );
  AOI211_X1 U14731 ( .C1(n9819), .C2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A(
        n11673), .B(n11672), .ZN(n11674) );
  NAND3_X1 U14732 ( .A1(n11676), .A2(n11675), .A3(n11674), .ZN(n11900) );
  AOI22_X1 U14733 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n9841), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11681) );
  AOI22_X1 U14734 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(n9815), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11680) );
  AOI22_X1 U14735 ( .A1(n9838), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(n9842), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11679) );
  AOI22_X1 U14736 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11678) );
  NAND4_X1 U14737 ( .A1(n11681), .A2(n11680), .A3(n11679), .A4(n11678), .ZN(
        n11686) );
  AOI22_X1 U14738 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n11826), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n11685) );
  AOI22_X1 U14739 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n11684) );
  AOI22_X1 U14740 ( .A1(n17024), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11825), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11683) );
  AOI22_X1 U14741 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n17069), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11682) );
  AOI22_X1 U14742 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n9815), .B2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n11690) );
  AOI22_X1 U14743 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11689) );
  AOI22_X1 U14744 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .B1(n9813), .B2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n11688) );
  AOI22_X1 U14745 ( .A1(n9811), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9842), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11687) );
  NAND4_X1 U14746 ( .A1(n11690), .A2(n11689), .A3(n11688), .A4(n11687), .ZN(
        n11697) );
  AOI22_X1 U14747 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n11695) );
  AOI22_X1 U14748 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .B1(
        n9809), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n11694) );
  AOI22_X1 U14749 ( .A1(n17048), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n9846), .B2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n11693) );
  AOI22_X1 U14750 ( .A1(n9841), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11692) );
  NAND4_X1 U14751 ( .A1(n11695), .A2(n11694), .A3(n11693), .A4(n11692), .ZN(
        n11696) );
  AOI22_X1 U14752 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(n9819), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11701) );
  AOI22_X1 U14753 ( .A1(n9838), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11825), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11700) );
  AOI22_X1 U14754 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n17024), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11699) );
  AOI22_X1 U14755 ( .A1(n9841), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11698) );
  NAND4_X1 U14756 ( .A1(n11701), .A2(n11700), .A3(n11699), .A4(n11698), .ZN(
        n11707) );
  AOI22_X1 U14757 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9809), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n11705) );
  AOI22_X1 U14758 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n11704) );
  AOI22_X1 U14759 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n9845), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n11703) );
  AOI22_X1 U14760 ( .A1(n9815), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n11702) );
  NAND4_X1 U14761 ( .A1(n11705), .A2(n11704), .A3(n11703), .A4(n11702), .ZN(
        n11706) );
  AOI22_X1 U14762 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17024), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11717) );
  AOI22_X1 U14763 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11716) );
  AOI22_X1 U14764 ( .A1(n9845), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n9815), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11708) );
  OAI21_X1 U14765 ( .B1(n11792), .B2(n20918), .A(n11708), .ZN(n11714) );
  AOI22_X1 U14766 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11825), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11712) );
  AOI22_X1 U14767 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n11711) );
  AOI22_X1 U14768 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11857), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n11710) );
  AOI22_X1 U14769 ( .A1(n15640), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9842), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11709) );
  NAND4_X1 U14770 ( .A1(n11712), .A2(n11711), .A3(n11710), .A4(n11709), .ZN(
        n11713) );
  AOI22_X1 U14771 ( .A1(n9809), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n17024), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n11721) );
  AOI22_X1 U14772 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n11720) );
  AOI22_X1 U14773 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(n9811), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11719) );
  AOI22_X1 U14774 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n9842), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n11718) );
  NAND4_X1 U14775 ( .A1(n11721), .A2(n11720), .A3(n11719), .A4(n11718), .ZN(
        n11727) );
  AOI22_X1 U14776 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11725) );
  AOI22_X1 U14777 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n17069), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11724) );
  AOI22_X1 U14778 ( .A1(n15640), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n11723) );
  AOI22_X1 U14779 ( .A1(n9845), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n9816), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11722) );
  NAND4_X1 U14780 ( .A1(n11725), .A2(n11724), .A3(n11723), .A4(n11722), .ZN(
        n11726) );
  INV_X1 U14781 ( .A(n11737), .ZN(n11740) );
  NAND2_X1 U14782 ( .A1(n17115), .A2(n17112), .ZN(n11731) );
  NAND4_X1 U14783 ( .A1(n18112), .A2(n18117), .A3(n11740), .A4(n11733), .ZN(
        n11739) );
  NOR2_X1 U14784 ( .A1(n18123), .A2(n17112), .ZN(n18567) );
  NOR2_X1 U14785 ( .A1(n18134), .A2(n18567), .ZN(n15745) );
  INV_X1 U14786 ( .A(n15745), .ZN(n11728) );
  NOR2_X1 U14787 ( .A1(n16313), .A2(n18094), .ZN(n11909) );
  NAND2_X1 U14788 ( .A1(n11728), .A2(n11909), .ZN(n11923) );
  NAND2_X1 U14789 ( .A1(n18123), .A2(n11730), .ZN(n11902) );
  AOI21_X1 U14790 ( .B1(n18106), .B2(n18094), .A(n18567), .ZN(n11729) );
  AOI21_X1 U14791 ( .B1(n11731), .B2(n11730), .A(n11729), .ZN(n11736) );
  NOR2_X1 U14792 ( .A1(n18134), .A2(n11733), .ZN(n11734) );
  NOR2_X1 U14793 ( .A1(n11910), .A2(n11900), .ZN(n11732) );
  OAI22_X1 U14794 ( .A1(n18117), .A2(n11734), .B1(n11733), .B2(n11732), .ZN(
        n11735) );
  NAND2_X1 U14795 ( .A1(n18106), .A2(n18112), .ZN(n11913) );
  NOR3_X1 U14796 ( .A1(n18128), .A2(n17115), .A3(n11913), .ZN(n15633) );
  NAND3_X1 U14797 ( .A1(n11740), .A2(n15633), .A3(n18100), .ZN(n11741) );
  NOR2_X1 U14798 ( .A1(n18604), .A2(P3_STATE2_REG_1__SCAN_IN), .ZN(n17751) );
  NAND2_X1 U14799 ( .A1(P3_STATE2_REG_2__SCAN_IN), .A2(n17751), .ZN(n18595) );
  NAND2_X1 U14800 ( .A1(n18088), .A2(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n11927) );
  XOR2_X1 U14801 ( .A(n11930), .B(n11927), .Z(n11752) );
  OAI22_X1 U14802 ( .A1(n18713), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B1(
        n18576), .B2(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n11747) );
  OAI21_X1 U14803 ( .B1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n18713), .A(
        n11743), .ZN(n11744) );
  OAI22_X1 U14804 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18580), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n11744), .ZN(n11750) );
  NOR2_X1 U14805 ( .A1(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n18580), .ZN(
        n11745) );
  NAND2_X1 U14806 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n11744), .ZN(
        n11749) );
  AOI22_X1 U14807 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n11750), .B1(
        n11745), .B2(n11749), .ZN(n11934) );
  NAND2_X1 U14808 ( .A1(n11748), .A2(n11747), .ZN(n11746) );
  OAI211_X1 U14809 ( .C1(n11748), .C2(n11747), .A(n11934), .B(n11746), .ZN(
        n11928) );
  INV_X1 U14810 ( .A(n11928), .ZN(n11932) );
  INV_X1 U14811 ( .A(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n18539) );
  AND2_X1 U14812 ( .A1(n11749), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n11751) );
  OAI22_X1 U14813 ( .A1(P3_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n18539), .B1(
        n11751), .B2(n11750), .ZN(n11931) );
  NAND2_X1 U14814 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .ZN(n11755) );
  INV_X1 U14815 ( .A(P3_REIP_REG_26__SCAN_IN), .ZN(n18672) );
  INV_X1 U14816 ( .A(P3_REIP_REG_25__SCAN_IN), .ZN(n18670) );
  NOR2_X1 U14817 ( .A1(n18672), .A2(n18670), .ZN(n11754) );
  INV_X1 U14818 ( .A(P3_REIP_REG_24__SCAN_IN), .ZN(n18669) );
  INV_X1 U14819 ( .A(P3_REIP_REG_23__SCAN_IN), .ZN(n20919) );
  INV_X1 U14820 ( .A(P3_REIP_REG_21__SCAN_IN), .ZN(n18663) );
  INV_X1 U14821 ( .A(P3_REIP_REG_19__SCAN_IN), .ZN(n18659) );
  INV_X1 U14822 ( .A(P3_REIP_REG_17__SCAN_IN), .ZN(n18655) );
  INV_X1 U14823 ( .A(P3_REIP_REG_15__SCAN_IN), .ZN(n18651) );
  INV_X1 U14824 ( .A(P3_REIP_REG_12__SCAN_IN), .ZN(n18645) );
  INV_X1 U14825 ( .A(P3_REIP_REG_5__SCAN_IN), .ZN(n18634) );
  INV_X1 U14826 ( .A(P3_REIP_REG_3__SCAN_IN), .ZN(n18629) );
  NAND2_X1 U14827 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_2__SCAN_IN), 
        .ZN(n16781) );
  NOR2_X1 U14828 ( .A1(n18629), .A2(n16781), .ZN(n16766) );
  NAND2_X1 U14829 ( .A1(P3_REIP_REG_4__SCAN_IN), .A2(n16766), .ZN(n16670) );
  NOR2_X1 U14830 ( .A1(n18634), .A2(n16670), .ZN(n16687) );
  INV_X1 U14831 ( .A(P3_REIP_REG_10__SCAN_IN), .ZN(n18641) );
  INV_X1 U14832 ( .A(P3_REIP_REG_9__SCAN_IN), .ZN(n18640) );
  NAND3_X1 U14833 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(P3_REIP_REG_6__SCAN_IN), 
        .A3(P3_REIP_REG_7__SCAN_IN), .ZN(n16688) );
  NOR3_X1 U14834 ( .A1(n18641), .A2(n18640), .A3(n16688), .ZN(n16671) );
  NAND3_X1 U14835 ( .A1(P3_REIP_REG_11__SCAN_IN), .A2(n16687), .A3(n16671), 
        .ZN(n16665) );
  NOR2_X1 U14836 ( .A1(n18645), .A2(n16665), .ZN(n16638) );
  NAND3_X1 U14837 ( .A1(P3_REIP_REG_14__SCAN_IN), .A2(P3_REIP_REG_13__SCAN_IN), 
        .A3(n16638), .ZN(n16622) );
  NOR2_X1 U14838 ( .A1(n18651), .A2(n16622), .ZN(n16614) );
  NAND2_X1 U14839 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n16614), .ZN(n16604) );
  NOR2_X1 U14840 ( .A1(n18655), .A2(n16604), .ZN(n16578) );
  NAND2_X1 U14841 ( .A1(P3_REIP_REG_18__SCAN_IN), .A2(n16578), .ZN(n16583) );
  NOR2_X1 U14842 ( .A1(n18659), .A2(n16583), .ZN(n16574) );
  NAND2_X1 U14843 ( .A1(P3_REIP_REG_20__SCAN_IN), .A2(n16574), .ZN(n16565) );
  NOR2_X1 U14844 ( .A1(n18663), .A2(n16565), .ZN(n16547) );
  NAND2_X1 U14845 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16547), .ZN(n16538) );
  NOR2_X1 U14846 ( .A1(n20919), .A2(n16538), .ZN(n16525) );
  INV_X1 U14847 ( .A(n16525), .ZN(n16536) );
  NOR2_X1 U14848 ( .A1(n18669), .A2(n16536), .ZN(n11756) );
  NOR2_X1 U14849 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(P3_STATE2_REG_3__SCAN_IN), .ZN(n18723) );
  NAND2_X1 U14850 ( .A1(n17751), .A2(n9805), .ZN(n18593) );
  OAI221_X1 U14851 ( .B1(n16802), .B2(n11754), .C1(n16802), .C2(n11756), .A(
        n16810), .ZN(n16488) );
  AOI221_X1 U14852 ( .B1(n18675), .B2(n16782), .C1(n11755), .C2(n16782), .A(
        n16488), .ZN(n16480) );
  NAND3_X1 U14853 ( .A1(P3_REIP_REG_26__SCAN_IN), .A2(n16518), .A3(
        P3_REIP_REG_25__SCAN_IN), .ZN(n16500) );
  NOR2_X1 U14854 ( .A1(n18675), .A2(n16500), .ZN(n16487) );
  NAND3_X1 U14855 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(P3_REIP_REG_29__SCAN_IN), 
        .A3(n16487), .ZN(n11762) );
  NOR2_X1 U14856 ( .A1(P3_REIP_REG_30__SCAN_IN), .A2(n11762), .ZN(n16471) );
  INV_X1 U14857 ( .A(n16471), .ZN(n11757) );
  INV_X1 U14858 ( .A(P3_REIP_REG_31__SCAN_IN), .ZN(n18684) );
  AOI21_X1 U14859 ( .B1(n16480), .B2(n11757), .A(n18684), .ZN(n11758) );
  INV_X1 U14860 ( .A(n11758), .ZN(n11769) );
  NAND2_X1 U14861 ( .A1(P3_EBX_REG_31__SCAN_IN), .A2(n16313), .ZN(n11759) );
  AOI211_X4 U14862 ( .C1(n18747), .C2(n18745), .A(n11760), .B(n11759), .ZN(
        n16811) );
  NOR3_X1 U14863 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(P3_EBX_REG_1__SCAN_IN), 
        .A3(P3_EBX_REG_2__SCAN_IN), .ZN(n16780) );
  NAND2_X1 U14864 ( .A1(n16780), .A2(n17091), .ZN(n16775) );
  INV_X1 U14865 ( .A(P3_EBX_REG_5__SCAN_IN), .ZN(n16748) );
  NAND2_X1 U14866 ( .A1(n16751), .A2(n16748), .ZN(n16747) );
  INV_X1 U14867 ( .A(P3_EBX_REG_7__SCAN_IN), .ZN(n17080) );
  NAND2_X1 U14868 ( .A1(n16730), .A2(n17080), .ZN(n16721) );
  INV_X1 U14869 ( .A(P3_EBX_REG_9__SCAN_IN), .ZN(n16701) );
  NAND2_X1 U14870 ( .A1(n16706), .A2(n16701), .ZN(n16699) );
  INV_X1 U14871 ( .A(P3_EBX_REG_11__SCAN_IN), .ZN(n16679) );
  NAND2_X1 U14872 ( .A1(n16683), .A2(n16679), .ZN(n16678) );
  INV_X1 U14873 ( .A(P3_EBX_REG_13__SCAN_IN), .ZN(n16654) );
  NAND2_X1 U14874 ( .A1(n16658), .A2(n16654), .ZN(n16653) );
  INV_X1 U14875 ( .A(P3_EBX_REG_15__SCAN_IN), .ZN(n16632) );
  NAND2_X1 U14876 ( .A1(n16636), .A2(n16632), .ZN(n16631) );
  INV_X1 U14877 ( .A(P3_EBX_REG_17__SCAN_IN), .ZN(n16612) );
  NAND2_X1 U14878 ( .A1(n16619), .A2(n16612), .ZN(n16605) );
  INV_X1 U14879 ( .A(P3_EBX_REG_19__SCAN_IN), .ZN(n16580) );
  NAND2_X1 U14880 ( .A1(n16596), .A2(n16580), .ZN(n16579) );
  INV_X1 U14881 ( .A(P3_EBX_REG_21__SCAN_IN), .ZN(n16562) );
  NAND2_X1 U14882 ( .A1(n16570), .A2(n16562), .ZN(n16561) );
  INV_X1 U14883 ( .A(P3_EBX_REG_23__SCAN_IN), .ZN(n16542) );
  NAND2_X1 U14884 ( .A1(n16548), .A2(n16542), .ZN(n16541) );
  INV_X1 U14885 ( .A(P3_EBX_REG_25__SCAN_IN), .ZN(n16520) );
  NAND2_X1 U14886 ( .A1(n16526), .A2(n16520), .ZN(n16519) );
  NOR2_X1 U14887 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16519), .ZN(n16507) );
  INV_X1 U14888 ( .A(P3_EBX_REG_27__SCAN_IN), .ZN(n16818) );
  NAND2_X1 U14889 ( .A1(n16507), .A2(n16818), .ZN(n16503) );
  NOR2_X1 U14890 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16503), .ZN(n16489) );
  INV_X1 U14891 ( .A(P3_EBX_REG_29__SCAN_IN), .ZN(n16856) );
  NAND2_X1 U14892 ( .A1(n16489), .A2(n16856), .ZN(n16466) );
  NOR2_X1 U14893 ( .A1(n16779), .A2(n16466), .ZN(n16473) );
  INV_X1 U14894 ( .A(P3_EBX_REG_30__SCAN_IN), .ZN(n16846) );
  NAND2_X1 U14895 ( .A1(n16473), .A2(n16846), .ZN(n11768) );
  AOI211_X4 U14896 ( .C1(P3_EBX_REG_31__SCAN_IN), .C2(n16313), .A(n11761), .B(
        n11760), .ZN(n16812) );
  INV_X1 U14897 ( .A(P3_REIP_REG_30__SCAN_IN), .ZN(n18681) );
  NOR3_X1 U14898 ( .A1(P3_REIP_REG_31__SCAN_IN), .A2(n18681), .A3(n11762), 
        .ZN(n11763) );
  AOI21_X1 U14899 ( .B1(n16812), .B2(P3_EBX_REG_31__SCAN_IN), .A(n11763), .ZN(
        n11764) );
  INV_X1 U14900 ( .A(n11764), .ZN(n11766) );
  NOR2_X1 U14901 ( .A1(n16798), .A2(n16310), .ZN(n11765) );
  NAND3_X1 U14902 ( .A1(n11769), .A2(n11768), .A3(n11767), .ZN(n11770) );
  AOI22_X1 U14903 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n11775) );
  AOI22_X1 U14904 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n11774) );
  AOI22_X1 U14905 ( .A1(n9841), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n11773) );
  AOI22_X1 U14906 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9846), .B2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n11772) );
  NAND4_X1 U14907 ( .A1(n11775), .A2(n11774), .A3(n11773), .A4(n11772), .ZN(
        n11781) );
  AOI22_X1 U14908 ( .A1(n17024), .A2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n11779) );
  AOI22_X1 U14909 ( .A1(n9810), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(n9816), .B2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n11778) );
  AOI22_X1 U14910 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n11777) );
  INV_X2 U14911 ( .A(n17006), .ZN(n16983) );
  AOI22_X1 U14912 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n11776) );
  NAND4_X1 U14913 ( .A1(n11779), .A2(n11778), .A3(n11777), .A4(n11776), .ZN(
        n11780) );
  AOI22_X1 U14914 ( .A1(n17048), .A2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n11785) );
  AOI22_X1 U14915 ( .A1(n9846), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n11784) );
  AOI22_X1 U14916 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(n9811), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n11783) );
  AOI22_X1 U14917 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n11782) );
  NAND4_X1 U14918 ( .A1(n11785), .A2(n11784), .A3(n11783), .A4(n11782), .ZN(
        n11791) );
  AOI22_X1 U14919 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n11789) );
  AOI22_X1 U14920 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n9819), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n11788) );
  AOI22_X1 U14921 ( .A1(n9810), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(n9830), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n11787) );
  AOI22_X1 U14922 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n9815), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n11786) );
  NAND4_X1 U14923 ( .A1(n11789), .A2(n11788), .A3(n11787), .A4(n11786), .ZN(
        n11790) );
  AOI22_X1 U14924 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n17024), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n11796) );
  AOI22_X1 U14925 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n9815), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n11795) );
  AOI22_X1 U14926 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n9810), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n11794) );
  AOI22_X1 U14927 ( .A1(n9845), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9842), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n11793) );
  NAND4_X1 U14928 ( .A1(n11796), .A2(n11795), .A3(n11794), .A4(n11793), .ZN(
        n11802) );
  AOI22_X1 U14929 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n11800) );
  AOI22_X1 U14930 ( .A1(n11827), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n11799) );
  AOI22_X1 U14931 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n11825), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n11798) );
  AOI22_X1 U14932 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(n9822), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n11797) );
  NAND4_X1 U14933 ( .A1(n11800), .A2(n11799), .A3(n11798), .A4(n11797), .ZN(
        n11801) );
  AOI22_X1 U14934 ( .A1(n11821), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11827), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n11803) );
  OAI21_X1 U14935 ( .B1(n11658), .B2(n18110), .A(n11803), .ZN(n11804) );
  INV_X1 U14936 ( .A(n11804), .ZN(n11811) );
  AOI22_X1 U14937 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11826), .B2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n11810) );
  AOI22_X1 U14938 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n11677), .B2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n11807) );
  INV_X1 U14939 ( .A(n11807), .ZN(n11808) );
  NAND3_X1 U14940 ( .A1(n11811), .A2(n11810), .A3(n11809), .ZN(n11818) );
  AOI22_X1 U14941 ( .A1(n17048), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n11816) );
  AOI22_X1 U14942 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n11815) );
  AOI22_X1 U14943 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n11819), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n11814) );
  AOI22_X1 U14944 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n9842), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n11813) );
  NAND4_X1 U14945 ( .A1(n11816), .A2(n11815), .A3(n11814), .A4(n11813), .ZN(
        n11817) );
  AOI22_X1 U14946 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n9818), .B1(
        P3_INSTQUEUE_REG_4__1__SCAN_IN), .B2(n9816), .ZN(n11834) );
  AOI22_X1 U14947 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n17049), .ZN(n11833) );
  INV_X1 U14948 ( .A(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n15598) );
  AOI22_X1 U14949 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n11819), .B1(
        n11691), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n11820) );
  OAI21_X1 U14950 ( .B1(n15622), .B2(n15598), .A(n11820), .ZN(n11832) );
  INV_X1 U14951 ( .A(n11822), .ZN(n11824) );
  NOR2_X1 U14952 ( .A1(n11824), .A2(n11823), .ZN(n11831) );
  AOI22_X1 U14953 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n11825), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n9842), .ZN(n11830) );
  AOI22_X1 U14954 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9822), .B1(n9829), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n11829) );
  AOI22_X1 U14955 ( .A1(n9823), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11826), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n11828) );
  AOI22_X1 U14956 ( .A1(n17024), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17049), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n11844) );
  AOI22_X1 U14957 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n17069), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n11843) );
  INV_X1 U14958 ( .A(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n20907) );
  AOI22_X1 U14959 ( .A1(n9845), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n11835) );
  OAI21_X1 U14960 ( .B1(n11812), .B2(n20907), .A(n11835), .ZN(n11841) );
  AOI22_X1 U14961 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(n9815), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n11839) );
  AOI22_X1 U14962 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11825), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n11838) );
  AOI22_X1 U14963 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n11837) );
  AOI22_X1 U14964 ( .A1(n15609), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9842), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n11836) );
  NAND4_X1 U14965 ( .A1(n11839), .A2(n11838), .A3(n11837), .A4(n11836), .ZN(
        n11840) );
  AOI211_X1 U14966 ( .C1(n9838), .C2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A(
        n11841), .B(n11840), .ZN(n11842) );
  NAND3_X1 U14967 ( .A1(n11844), .A2(n11843), .A3(n11842), .ZN(n11948) );
  NAND2_X1 U14968 ( .A1(n11874), .A2(n11948), .ZN(n11855) );
  AOI22_X1 U14969 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n11854) );
  AOI22_X1 U14970 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9815), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n11853) );
  AOI22_X1 U14971 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n11845) );
  OAI21_X1 U14972 ( .B1(n11812), .B2(n20918), .A(n11845), .ZN(n11851) );
  AOI22_X1 U14973 ( .A1(n9841), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n9846), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n11849) );
  AOI22_X1 U14974 ( .A1(n17024), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n11848) );
  AOI22_X1 U14975 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n9819), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n11847) );
  AOI22_X1 U14976 ( .A1(n9811), .A2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n11846) );
  NAND4_X1 U14977 ( .A1(n11849), .A2(n11848), .A3(n11847), .A4(n11846), .ZN(
        n11850) );
  AOI211_X1 U14978 ( .C1(n17019), .C2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A(
        n11851), .B(n11850), .ZN(n11852) );
  NAND3_X1 U14979 ( .A1(n11854), .A2(n11853), .A3(n11852), .ZN(n17680) );
  INV_X1 U14980 ( .A(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n17781) );
  INV_X1 U14981 ( .A(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n18026) );
  XNOR2_X1 U14982 ( .A(n17233), .B(n11855), .ZN(n11877) );
  INV_X1 U14983 ( .A(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18708) );
  NOR2_X1 U14984 ( .A1(n17250), .A2(n18708), .ZN(n11868) );
  AOI22_X1 U14985 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n17069), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n11867) );
  AOI22_X1 U14986 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(n9816), .B2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n11866) );
  AOI22_X1 U14987 ( .A1(n9823), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11691), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n11856) );
  OAI21_X1 U14988 ( .B1(n11658), .B2(n18098), .A(n11856), .ZN(n11864) );
  AOI22_X1 U14989 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n9832), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n11862) );
  AOI22_X1 U14990 ( .A1(n11857), .A2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n15560), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n11861) );
  AOI22_X1 U14991 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n11826), .B2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n11860) );
  AOI22_X1 U14992 ( .A1(n11819), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9842), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n11859) );
  NAND4_X1 U14993 ( .A1(n11862), .A2(n11861), .A3(n11860), .A4(n11859), .ZN(
        n11863) );
  AOI211_X1 U14994 ( .C1(n9818), .C2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A(
        n11864), .B(n11863), .ZN(n11865) );
  NAND3_X1 U14995 ( .A1(n11867), .A2(n11866), .A3(n11865), .ZN(n15746) );
  NAND2_X1 U14996 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15746), .ZN(
        n17747) );
  NOR2_X1 U14997 ( .A1(n17740), .A2(n17747), .ZN(n17737) );
  NOR2_X1 U14998 ( .A1(n11868), .A2(n17737), .ZN(n17727) );
  XNOR2_X1 U14999 ( .A(n17244), .B(n17250), .ZN(n11870) );
  XNOR2_X1 U15000 ( .A(n11870), .B(n11869), .ZN(n17726) );
  NOR2_X1 U15001 ( .A1(n11869), .A2(n11870), .ZN(n11871) );
  INV_X1 U15002 ( .A(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18041) );
  XOR2_X1 U15003 ( .A(n17240), .B(n11950), .Z(n11872) );
  XOR2_X1 U15004 ( .A(n18041), .B(n11872), .Z(n17716) );
  AND2_X1 U15005 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n11872), .ZN(
        n11873) );
  INV_X1 U15006 ( .A(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18021) );
  XOR2_X1 U15007 ( .A(n11948), .B(n11874), .Z(n11875) );
  XOR2_X1 U15008 ( .A(n18021), .B(n11875), .Z(n17701) );
  NOR2_X1 U15009 ( .A1(n17702), .A2(n17701), .ZN(n17700) );
  NOR2_X1 U15010 ( .A1(n17700), .A2(n11876), .ZN(n11878) );
  NOR2_X1 U15011 ( .A1(n11878), .A2(n11877), .ZN(n11879) );
  INV_X1 U15012 ( .A(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n18019) );
  XOR2_X1 U15013 ( .A(n17680), .B(n11880), .Z(n11881) );
  XOR2_X1 U15014 ( .A(n18019), .B(n11881), .Z(n17674) );
  NOR2_X2 U15015 ( .A1(n17673), .A2(n11882), .ZN(n17603) );
  AOI21_X1 U15016 ( .B1(n11899), .B2(n16315), .A(n17649), .ZN(n11883) );
  INV_X1 U15017 ( .A(n11883), .ZN(n11884) );
  NOR2_X1 U15018 ( .A1(n17603), .A2(n11884), .ZN(n11885) );
  INV_X1 U15019 ( .A(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n18009) );
  XNOR2_X1 U15020 ( .A(n11884), .B(n17603), .ZN(n17669) );
  NOR2_X1 U15021 ( .A1(n18009), .A2(n17669), .ZN(n17668) );
  INV_X1 U15022 ( .A(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n17988) );
  INV_X1 U15023 ( .A(n17647), .ZN(n17576) );
  INV_X1 U15024 ( .A(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17910) );
  NAND2_X1 U15025 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17959) );
  INV_X1 U15026 ( .A(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n17608) );
  NOR2_X1 U15027 ( .A1(n17959), .A2(n17608), .ZN(n17926) );
  NAND2_X1 U15028 ( .A1(n17926), .A2(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n17911) );
  INV_X1 U15029 ( .A(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n17934) );
  NOR2_X1 U15030 ( .A1(n17911), .A2(n17934), .ZN(n17916) );
  INV_X1 U15031 ( .A(n17916), .ZN(n17914) );
  NOR2_X1 U15032 ( .A1(n17910), .A2(n17914), .ZN(n17894) );
  NAND2_X1 U15033 ( .A1(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n17894), .ZN(
        n17870) );
  NOR2_X1 U15034 ( .A1(n17576), .A2(n17870), .ZN(n11893) );
  INV_X1 U15035 ( .A(n11893), .ZN(n17529) );
  INV_X1 U15036 ( .A(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n17888) );
  NOR2_X1 U15037 ( .A1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17630) );
  NOR3_X1 U15038 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n11887) );
  AOI21_X1 U15039 ( .B1(n17542), .B2(n11887), .A(n17649), .ZN(n17528) );
  INV_X1 U15040 ( .A(n11888), .ZN(n11889) );
  AOI21_X1 U15041 ( .B1(n17529), .B2(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n11889), .ZN(n17520) );
  INV_X1 U15042 ( .A(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17866) );
  NAND2_X1 U15043 ( .A1(n17520), .A2(n17866), .ZN(n17519) );
  NOR2_X1 U15044 ( .A1(n17888), .A2(n17866), .ZN(n17865) );
  NAND2_X1 U15045 ( .A1(n17865), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n17480) );
  INV_X1 U15046 ( .A(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n17478) );
  NAND2_X1 U15047 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17475) );
  NOR2_X1 U15048 ( .A1(n17478), .A2(n17475), .ZN(n17815) );
  NAND2_X1 U15049 ( .A1(n17815), .A2(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n11918) );
  NOR2_X1 U15050 ( .A1(n17480), .A2(n11918), .ZN(n17792) );
  INV_X1 U15051 ( .A(n17792), .ZN(n17808) );
  INV_X1 U15052 ( .A(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n17798) );
  NOR2_X1 U15053 ( .A1(n17808), .A2(n17798), .ZN(n17769) );
  NAND2_X1 U15054 ( .A1(n11893), .A2(n17769), .ZN(n11891) );
  NOR2_X1 U15055 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17649), .ZN(
        n17511) );
  INV_X1 U15056 ( .A(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n17855) );
  NAND2_X1 U15057 ( .A1(n17511), .A2(n17855), .ZN(n11890) );
  NOR2_X1 U15058 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n11890), .ZN(
        n17473) );
  NAND2_X1 U15059 ( .A1(n17473), .A2(n17478), .ZN(n17457) );
  INV_X1 U15060 ( .A(n11918), .ZN(n17433) );
  NAND2_X1 U15061 ( .A1(n17865), .A2(n11893), .ZN(n17471) );
  NAND3_X1 U15062 ( .A1(n17433), .A2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n17472), .ZN(n17435) );
  NOR3_X1 U15063 ( .A1(n17426), .A2(n17435), .A3(n17798), .ZN(n11895) );
  NAND2_X1 U15064 ( .A1(n17604), .A2(n17419), .ZN(n11894) );
  OAI221_X1 U15065 ( .B1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n17604), 
        .C1(n17781), .C2(n11895), .A(n11894), .ZN(n17401) );
  NOR2_X1 U15066 ( .A1(n17401), .A2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n17400) );
  NAND2_X1 U15067 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17757) );
  NAND2_X1 U15068 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n11898), .ZN(
        n15668) );
  AND2_X2 U15069 ( .A1(n11979), .A2(n15668), .ZN(n17387) );
  NAND2_X1 U15070 ( .A1(n17387), .A2(n17649), .ZN(n17386) );
  NAND2_X1 U15071 ( .A1(n17386), .A2(n11979), .ZN(n17378) );
  INV_X1 U15072 ( .A(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n17375) );
  AOI22_X1 U15073 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17649), .B1(
        n17604), .B2(n17375), .ZN(n17379) );
  NOR2_X1 U15074 ( .A1(n18100), .A2(n11900), .ZN(n11901) );
  NAND2_X1 U15075 ( .A1(n11901), .A2(n17112), .ZN(n11941) );
  NOR2_X1 U15076 ( .A1(n11910), .A2(n11912), .ZN(n11903) );
  OAI211_X1 U15077 ( .C1(n18128), .C2(n18117), .A(n11903), .B(n11902), .ZN(
        n11922) );
  AND2_X1 U15078 ( .A1(n18532), .A2(n11904), .ZN(n11905) );
  AND2_X1 U15079 ( .A1(n11906), .A2(n11905), .ZN(n11907) );
  NAND2_X1 U15080 ( .A1(n17377), .A2(n11907), .ZN(n11944) );
  NOR2_X1 U15081 ( .A1(n11910), .A2(n11909), .ZN(n18758) );
  NOR2_X1 U15082 ( .A1(n17112), .A2(n18117), .ZN(n18545) );
  INV_X1 U15083 ( .A(n18545), .ZN(n11911) );
  INV_X1 U15084 ( .A(n17967), .ZN(n17933) );
  INV_X1 U15085 ( .A(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n17768) );
  INV_X1 U15086 ( .A(n11913), .ZN(n18544) );
  NAND2_X1 U15087 ( .A1(n16313), .A2(n9878), .ZN(n11916) );
  INV_X1 U15088 ( .A(n11914), .ZN(n11915) );
  NAND4_X1 U15089 ( .A1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n11919) );
  NOR3_X1 U15090 ( .A1(n11918), .A2(n11919), .A3(n17768), .ZN(n17376) );
  NOR2_X1 U15091 ( .A1(n17808), .A2(n11919), .ZN(n15675) );
  INV_X1 U15092 ( .A(n15675), .ZN(n17756) );
  INV_X1 U15093 ( .A(n17870), .ZN(n11975) );
  NAND4_X1 U15094 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A4(
        P3_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n18000) );
  NOR2_X1 U15095 ( .A1(n18009), .A2(n18000), .ZN(n17992) );
  NAND2_X1 U15096 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17992), .ZN(
        n17868) );
  NAND2_X1 U15097 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n17985) );
  NOR2_X1 U15098 ( .A1(n17868), .A2(n17985), .ZN(n17882) );
  NAND2_X1 U15099 ( .A1(n11975), .A2(n17882), .ZN(n17818) );
  AOI21_X1 U15100 ( .B1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n17984) );
  OR2_X1 U15101 ( .A1(n17868), .A2(n17984), .ZN(n17881) );
  NOR2_X1 U15102 ( .A1(n17870), .A2(n17881), .ZN(n17820) );
  INV_X1 U15103 ( .A(n17820), .ZN(n17861) );
  OAI21_X1 U15104 ( .B1(n17756), .B2(n17861), .A(n18540), .ZN(n17758) );
  INV_X1 U15105 ( .A(n17758), .ZN(n11920) );
  AOI221_X1 U15106 ( .B1(n17756), .B2(n18549), .C1(n17818), .C2(n18549), .A(
        n11920), .ZN(n11921) );
  NAND3_X1 U15107 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18049) );
  NOR2_X1 U15108 ( .A1(n18049), .A2(n17868), .ZN(n17974) );
  NAND2_X1 U15109 ( .A1(n11975), .A2(n17974), .ZN(n17885) );
  OAI21_X1 U15110 ( .B1(n17480), .B2(n17885), .A(n18566), .ZN(n17841) );
  OAI211_X1 U15111 ( .C1(n18554), .C2(n17376), .A(n11921), .B(n17841), .ZN(
        n15730) );
  AOI21_X1 U15112 ( .B1(n17933), .B2(n17768), .A(n15730), .ZN(n15673) );
  INV_X1 U15113 ( .A(n11922), .ZN(n11925) );
  OAI211_X1 U15114 ( .C1(n11926), .C2(n11925), .A(n11924), .B(n11923), .ZN(
        n14223) );
  OAI21_X1 U15115 ( .B1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n18088), .A(
        n11927), .ZN(n11929) );
  OAI21_X1 U15116 ( .B1(n11928), .B2(n11929), .A(n11935), .ZN(n18531) );
  NOR2_X1 U15117 ( .A1(n11930), .A2(n11929), .ZN(n11933) );
  NAND2_X1 U15118 ( .A1(n18106), .A2(n17115), .ZN(n11939) );
  INV_X1 U15119 ( .A(n11935), .ZN(n18530) );
  XNOR2_X1 U15120 ( .A(n18100), .B(n18106), .ZN(n11936) );
  AOI21_X1 U15121 ( .B1(n11936), .B2(n18744), .A(n18615), .ZN(n16448) );
  INV_X1 U15122 ( .A(n16448), .ZN(n11937) );
  OAI21_X1 U15123 ( .B1(n18530), .B2(n11937), .A(n11939), .ZN(n11938) );
  OAI21_X1 U15124 ( .B1(n18535), .B2(n11939), .A(n11938), .ZN(n11940) );
  OAI21_X1 U15125 ( .B1(n11941), .B2(n18531), .A(n11940), .ZN(n11942) );
  NAND2_X1 U15126 ( .A1(n11944), .A2(n11943), .ZN(n11973) );
  INV_X1 U15127 ( .A(n17911), .ZN(n17941) );
  INV_X1 U15128 ( .A(n11953), .ZN(n11945) );
  NOR2_X1 U15129 ( .A1(n11951), .A2(n17240), .ZN(n11949) );
  NAND2_X1 U15130 ( .A1(n11949), .A2(n11948), .ZN(n11947) );
  NOR2_X1 U15131 ( .A1(n17233), .A2(n11947), .ZN(n17679) );
  NAND2_X1 U15132 ( .A1(n17679), .A2(n17680), .ZN(n11946) );
  NOR2_X1 U15133 ( .A1(n16315), .A2(n11946), .ZN(n11967) );
  XNOR2_X1 U15134 ( .A(n11904), .B(n11946), .ZN(n11964) );
  XOR2_X1 U15135 ( .A(n11947), .B(n17233), .Z(n11960) );
  INV_X1 U15136 ( .A(n11948), .ZN(n17236) );
  XOR2_X1 U15137 ( .A(n11949), .B(n17236), .Z(n11958) );
  NOR2_X1 U15138 ( .A1(n11958), .A2(n18021), .ZN(n11959) );
  XNOR2_X1 U15139 ( .A(n17240), .B(n11951), .ZN(n11956) );
  NOR2_X1 U15140 ( .A1(n11956), .A2(n18041), .ZN(n11957) );
  INV_X1 U15141 ( .A(n11950), .ZN(n11952) );
  AOI21_X1 U15142 ( .B1(n11952), .B2(n15746), .A(n11951), .ZN(n11954) );
  NOR2_X1 U15143 ( .A1(n11954), .A2(n11869), .ZN(n11955) );
  NOR2_X1 U15144 ( .A1(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A2(n15746), .ZN(
        n17749) );
  NAND2_X1 U15145 ( .A1(n17749), .A2(n17740), .ZN(n17739) );
  OAI211_X1 U15146 ( .C1(P3_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(n17250), .A(
        n11953), .B(n17739), .ZN(n17730) );
  XOR2_X1 U15147 ( .A(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n11954), .Z(
        n17729) );
  NOR2_X1 U15148 ( .A1(n17730), .A2(n17729), .ZN(n17728) );
  NOR2_X1 U15149 ( .A1(n11955), .A2(n17728), .ZN(n17714) );
  XOR2_X1 U15150 ( .A(n11956), .B(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .Z(
        n17713) );
  NOR2_X1 U15151 ( .A1(n17714), .A2(n17713), .ZN(n17712) );
  NOR2_X1 U15152 ( .A1(n11957), .A2(n17712), .ZN(n17707) );
  XOR2_X1 U15153 ( .A(n11958), .B(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .Z(
        n17706) );
  NOR2_X1 U15154 ( .A1(n17707), .A2(n17706), .ZN(n17705) );
  NOR2_X1 U15155 ( .A1(n11959), .A2(n17705), .ZN(n17692) );
  XOR2_X1 U15156 ( .A(n18026), .B(n11960), .Z(n17691) );
  INV_X1 U15157 ( .A(n17679), .ZN(n17677) );
  INV_X1 U15158 ( .A(n17680), .ZN(n17681) );
  XNOR2_X1 U15159 ( .A(n17677), .B(n17681), .ZN(n11962) );
  AOI222_X1 U15160 ( .A1(n17678), .A2(n18019), .B1(n17678), .B2(n11962), .C1(
        n18019), .C2(n11962), .ZN(n11965) );
  NOR2_X1 U15161 ( .A1(n11964), .A2(n11965), .ZN(n17659) );
  NOR2_X1 U15162 ( .A1(n17659), .A2(n18009), .ZN(n11963) );
  NAND2_X1 U15163 ( .A1(n11967), .A2(n11963), .ZN(n11968) );
  INV_X1 U15164 ( .A(n11963), .ZN(n17660) );
  AND2_X1 U15165 ( .A1(n11965), .A2(n11964), .ZN(n17661) );
  AOI21_X1 U15166 ( .B1(n11967), .B2(n17660), .A(n17661), .ZN(n11966) );
  OAI21_X1 U15167 ( .B1(n11967), .B2(n17660), .A(n11966), .ZN(n17651) );
  NAND2_X1 U15168 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n17651), .ZN(
        n17650) );
  NAND2_X2 U15169 ( .A1(n11968), .A2(n17650), .ZN(n17606) );
  INV_X1 U15170 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17550) );
  NOR2_X2 U15171 ( .A1(n17556), .A2(n17550), .ZN(n17902) );
  NAND2_X1 U15172 ( .A1(n17902), .A2(n15675), .ZN(n17762) );
  NOR2_X1 U15173 ( .A1(n17375), .A2(n17768), .ZN(n15677) );
  INV_X1 U15174 ( .A(n15677), .ZN(n11969) );
  NOR2_X1 U15175 ( .A1(n17762), .A2(n11969), .ZN(n16341) );
  INV_X1 U15176 ( .A(n18052), .ZN(n18534) );
  NAND2_X1 U15177 ( .A1(n17647), .A2(n17894), .ZN(n17564) );
  NAND2_X1 U15178 ( .A1(n15675), .A2(n17896), .ZN(n17374) );
  INV_X1 U15179 ( .A(n17374), .ZN(n17760) );
  NAND2_X1 U15180 ( .A1(n15677), .A2(n17760), .ZN(n16330) );
  INV_X1 U15181 ( .A(n16330), .ZN(n11970) );
  NAND2_X1 U15182 ( .A1(n16315), .A2(n18532), .ZN(n17897) );
  OAI22_X1 U15183 ( .A1(n16341), .A2(n18534), .B1(n11970), .B2(n17897), .ZN(
        n11972) );
  NOR2_X1 U15184 ( .A1(n9820), .A2(n17375), .ZN(n11971) );
  OAI21_X1 U15185 ( .B1(n11973), .B2(n11972), .A(n11971), .ZN(n11982) );
  NAND2_X1 U15186 ( .A1(n18532), .A2(n18073), .ZN(n18077) );
  AND2_X1 U15187 ( .A1(n18066), .A2(n17649), .ZN(n11974) );
  NAND2_X1 U15188 ( .A1(n17377), .A2(n11974), .ZN(n11977) );
  INV_X1 U15189 ( .A(n17606), .ZN(n17954) );
  OAI22_X1 U15190 ( .A1(n17954), .A2(n18534), .B1(n17897), .B2(n17576), .ZN(
        n17869) );
  INV_X1 U15191 ( .A(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n18724) );
  NAND2_X1 U15192 ( .A1(n18568), .A2(n18724), .ZN(n18067) );
  NAND2_X1 U15193 ( .A1(n18067), .A2(n18045), .ZN(n18044) );
  OAI22_X1 U15194 ( .A1(n18561), .A2(n17861), .B1(n17818), .B2(n18044), .ZN(
        n17779) );
  AOI21_X1 U15195 ( .B1(n11975), .B2(n17869), .A(n17779), .ZN(n17809) );
  NOR3_X1 U15196 ( .A1(n17809), .A2(n18061), .A3(n17480), .ZN(n17840) );
  NAND2_X1 U15197 ( .A1(n11978), .A2(n17375), .ZN(n11981) );
  NAND2_X1 U15198 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n9820), .ZN(n17370) );
  OR3_X1 U15199 ( .A1(n11979), .A2(n17909), .A3(n17379), .ZN(n11980) );
  NAND4_X1 U15200 ( .A1(n11982), .A2(n11981), .A3(n17370), .A4(n11980), .ZN(
        P3_U2834) );
  NAND2_X1 U15201 ( .A1(n11997), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12168) );
  NAND2_X1 U15202 ( .A1(n14171), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n12018) );
  NOR2_X2 U15203 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n12452) );
  XNOR2_X1 U15204 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .B(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n14431) );
  INV_X2 U15205 ( .A(P1_STATE2_REG_2__SCAN_IN), .ZN(n20691) );
  AOI21_X1 U15206 ( .B1(n12452), .B2(n14431), .A(n12485), .ZN(n11984) );
  INV_X1 U15207 ( .A(n12424), .ZN(n12451) );
  NAND2_X1 U15208 ( .A1(n12451), .A2(P1_EAX_REG_2__SCAN_IN), .ZN(n11983) );
  OAI211_X1 U15209 ( .C1(n12018), .C2(n11235), .A(n11984), .B(n11983), .ZN(
        n11985) );
  INV_X1 U15210 ( .A(n11985), .ZN(n11986) );
  NAND2_X1 U15211 ( .A1(n12485), .A2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(
        n12006) );
  NAND2_X1 U15212 ( .A1(n11988), .A2(n12006), .ZN(n13647) );
  INV_X1 U15213 ( .A(n13647), .ZN(n12005) );
  XNOR2_X2 U15214 ( .A(n11989), .B(n11990), .ZN(n13700) );
  NAND2_X1 U15215 ( .A1(n13700), .A2(n12130), .ZN(n11995) );
  AOI22_X1 U15216 ( .A1(n12451), .A2(P1_EAX_REG_1__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n20691), .ZN(n11993) );
  INV_X1 U15217 ( .A(n12018), .ZN(n11991) );
  NAND2_X1 U15218 ( .A1(n11991), .A2(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n11992) );
  AND2_X1 U15219 ( .A1(n11993), .A2(n11992), .ZN(n11994) );
  NAND2_X1 U15220 ( .A1(n11995), .A2(n11994), .ZN(n13540) );
  NAND2_X1 U15221 ( .A1(n9828), .A2(n11997), .ZN(n11998) );
  NAND2_X1 U15222 ( .A1(n11998), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n13487) );
  INV_X1 U15223 ( .A(n14282), .ZN(n20217) );
  NAND2_X1 U15224 ( .A1(n20691), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n12001) );
  NAND2_X1 U15225 ( .A1(n11999), .A2(P1_EAX_REG_0__SCAN_IN), .ZN(n12000) );
  OAI211_X1 U15226 ( .C1(n12018), .C2(n14284), .A(n12001), .B(n12000), .ZN(
        n12002) );
  AOI21_X1 U15227 ( .B1(n20217), .B2(n12130), .A(n12002), .ZN(n13488) );
  OR2_X1 U15228 ( .A1(n13487), .A2(n13488), .ZN(n13489) );
  NAND2_X1 U15229 ( .A1(n13488), .A2(n12452), .ZN(n12003) );
  NAND2_X1 U15230 ( .A1(n13489), .A2(n12003), .ZN(n13539) );
  NAND2_X1 U15231 ( .A1(n13540), .A2(n13539), .ZN(n13646) );
  INV_X1 U15232 ( .A(n13646), .ZN(n12004) );
  NAND2_X1 U15233 ( .A1(n12005), .A2(n12004), .ZN(n13649) );
  NAND2_X1 U15234 ( .A1(n20766), .A2(n12130), .ZN(n12015) );
  INV_X1 U15235 ( .A(n12008), .ZN(n12010) );
  INV_X1 U15236 ( .A(n12020), .ZN(n12009) );
  OAI21_X1 U15237 ( .B1(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n12010), .A(
        n12009), .ZN(n19940) );
  AOI22_X1 U15238 ( .A1(n12452), .A2(n19940), .B1(n12485), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n12012) );
  NAND2_X1 U15239 ( .A1(n12451), .A2(P1_EAX_REG_3__SCAN_IN), .ZN(n12011) );
  OAI211_X1 U15240 ( .C1(n12018), .C2(n10990), .A(n12012), .B(n12011), .ZN(
        n12013) );
  INV_X1 U15241 ( .A(n12013), .ZN(n12014) );
  NAND2_X1 U15242 ( .A1(n12015), .A2(n12014), .ZN(n13710) );
  NAND2_X1 U15243 ( .A1(n13711), .A2(n13710), .ZN(n13709) );
  NAND2_X1 U15244 ( .A1(n20691), .A2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(
        n12017) );
  NAND2_X1 U15245 ( .A1(n12451), .A2(P1_EAX_REG_4__SCAN_IN), .ZN(n12016) );
  OAI211_X1 U15246 ( .C1(n12018), .C2(n13690), .A(n12017), .B(n12016), .ZN(
        n12019) );
  NAND2_X1 U15247 ( .A1(n12019), .A2(n12484), .ZN(n12022) );
  OAI21_X1 U15248 ( .B1(n12020), .B2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n12025), .ZN(n19925) );
  NAND2_X1 U15249 ( .A1(n19925), .A2(n12452), .ZN(n12021) );
  NAND2_X1 U15250 ( .A1(n12022), .A2(n12021), .ZN(n12023) );
  NOR2_X2 U15251 ( .A1(n13709), .A2(n13776), .ZN(n13774) );
  AOI22_X1 U15252 ( .A1(n11999), .A2(P1_EAX_REG_5__SCAN_IN), .B1(n12485), .B2(
        P1_PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n12027) );
  AOI21_X1 U15253 ( .B1(n12025), .B2(n15916), .A(n12029), .ZN(n15912) );
  INV_X1 U15254 ( .A(n15912), .ZN(n19921) );
  NAND2_X1 U15255 ( .A1(n19921), .A2(n12452), .ZN(n12026) );
  NAND2_X1 U15256 ( .A1(n13774), .A2(n13806), .ZN(n13804) );
  INV_X1 U15257 ( .A(n13804), .ZN(n12036) );
  INV_X1 U15258 ( .A(P1_EAX_REG_6__SCAN_IN), .ZN(n12032) );
  OAI21_X1 U15259 ( .B1(n12029), .B2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n12037), .ZN(n19906) );
  NAND2_X1 U15260 ( .A1(n19906), .A2(n12452), .ZN(n12031) );
  NAND2_X1 U15261 ( .A1(n12485), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(
        n12030) );
  OAI211_X1 U15262 ( .C1(n12424), .C2(n12032), .A(n12031), .B(n12030), .ZN(
        n12033) );
  NAND2_X1 U15263 ( .A1(n12036), .A2(n12035), .ZN(n13824) );
  INV_X1 U15264 ( .A(n13824), .ZN(n12046) );
  INV_X1 U15265 ( .A(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n12042) );
  INV_X1 U15266 ( .A(n12485), .ZN(n12203) );
  NAND2_X1 U15267 ( .A1(n11999), .A2(P1_EAX_REG_7__SCAN_IN), .ZN(n12041) );
  NAND2_X1 U15268 ( .A1(n12037), .A2(n12042), .ZN(n12039) );
  NAND2_X1 U15269 ( .A1(n12039), .A2(n12057), .ZN(n19901) );
  NAND2_X1 U15270 ( .A1(n19901), .A2(n12452), .ZN(n12040) );
  OAI211_X1 U15271 ( .C1(n12042), .C2(n12203), .A(n12041), .B(n12040), .ZN(
        n12043) );
  AOI21_X1 U15272 ( .B1(n12044), .B2(n12130), .A(n12043), .ZN(n13884) );
  INV_X1 U15273 ( .A(n13884), .ZN(n12045) );
  NAND2_X1 U15274 ( .A1(n12046), .A2(n12045), .ZN(n13883) );
  AOI22_X1 U15275 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11146), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12050) );
  AOI22_X1 U15276 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12049) );
  AOI22_X1 U15277 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12048) );
  AOI22_X1 U15278 ( .A1(n11167), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12047) );
  NAND4_X1 U15279 ( .A1(n12050), .A2(n12049), .A3(n12048), .A4(n12047), .ZN(
        n12056) );
  AOI22_X1 U15280 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12054) );
  AOI22_X1 U15281 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n11047), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12053) );
  AOI22_X1 U15282 ( .A1(n12458), .A2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n12468), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12052) );
  AOI22_X1 U15283 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12051) );
  NAND4_X1 U15284 ( .A1(n12054), .A2(n12053), .A3(n12052), .A4(n12051), .ZN(
        n12055) );
  OAI21_X1 U15285 ( .B1(n12056), .B2(n12055), .A(n12130), .ZN(n12060) );
  XNOR2_X1 U15286 ( .A(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .B(n12061), .ZN(
        n14417) );
  AOI22_X1 U15287 ( .A1(n12452), .A2(n14417), .B1(n12485), .B2(
        P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n12059) );
  NAND2_X1 U15288 ( .A1(n11999), .A2(P1_EAX_REG_8__SCAN_IN), .ZN(n12058) );
  AOI21_X1 U15289 ( .B1(n21011), .B2(n12062), .A(n12091), .ZN(n19886) );
  OR2_X1 U15290 ( .A1(n19886), .A2(n12484), .ZN(n12077) );
  AOI22_X1 U15291 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12066) );
  AOI22_X1 U15292 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12299), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12065) );
  AOI22_X1 U15293 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11167), .B2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12064) );
  AOI22_X1 U15294 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n12468), .B2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12063) );
  NAND4_X1 U15295 ( .A1(n12066), .A2(n12065), .A3(n12064), .A4(n12063), .ZN(
        n12072) );
  AOI22_X1 U15296 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11146), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12070) );
  AOI22_X1 U15297 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12069) );
  AOI22_X1 U15298 ( .A1(n11152), .A2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12068) );
  AOI22_X1 U15299 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12067) );
  NAND4_X1 U15300 ( .A1(n12070), .A2(n12069), .A3(n12068), .A4(n12067), .ZN(
        n12071) );
  OAI21_X1 U15301 ( .B1(n12072), .B2(n12071), .A(n12130), .ZN(n12075) );
  NAND2_X1 U15302 ( .A1(n11999), .A2(P1_EAX_REG_9__SCAN_IN), .ZN(n12074) );
  NAND2_X1 U15303 ( .A1(n12485), .A2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n12073) );
  AND3_X1 U15304 ( .A1(n12075), .A2(n12074), .A3(n12073), .ZN(n12076) );
  NAND2_X1 U15305 ( .A1(n12077), .A2(n12076), .ZN(n13973) );
  AOI22_X1 U15306 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n12458), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12081) );
  AOI22_X1 U15307 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11047), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12080) );
  AOI22_X1 U15308 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12079) );
  AOI22_X1 U15309 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12078) );
  NAND4_X1 U15310 ( .A1(n12081), .A2(n12080), .A3(n12079), .A4(n12078), .ZN(
        n12087) );
  AOI22_X1 U15311 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n11154), .B2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12085) );
  AOI22_X1 U15312 ( .A1(n12467), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12084) );
  AOI22_X1 U15313 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12083) );
  AOI22_X1 U15314 ( .A1(n11167), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12082) );
  NAND4_X1 U15315 ( .A1(n12085), .A2(n12084), .A3(n12083), .A4(n12082), .ZN(
        n12086) );
  NOR2_X1 U15316 ( .A1(n12087), .A2(n12086), .ZN(n12090) );
  XNOR2_X1 U15317 ( .A(n12091), .B(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14691) );
  NAND2_X1 U15318 ( .A1(n14691), .A2(n12452), .ZN(n12089) );
  AOI22_X1 U15319 ( .A1(n11999), .A2(P1_EAX_REG_10__SCAN_IN), .B1(n12485), 
        .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n12088) );
  OAI211_X1 U15320 ( .C1(n12090), .C2(n12168), .A(n12089), .B(n12088), .ZN(
        n14060) );
  NAND2_X1 U15321 ( .A1(n12451), .A2(P1_EAX_REG_11__SCAN_IN), .ZN(n12094) );
  OAI21_X1 U15322 ( .B1(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n12092), .A(
        n12148), .ZN(n15897) );
  AOI22_X1 U15323 ( .A1(n12452), .A2(n15897), .B1(n12485), .B2(
        P1_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n12093) );
  NAND2_X1 U15324 ( .A1(n12094), .A2(n12093), .ZN(n14123) );
  AOI22_X1 U15325 ( .A1(n12458), .A2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n11146), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12098) );
  AOI22_X1 U15326 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12097) );
  AOI22_X1 U15327 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12299), .B2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12096) );
  AOI22_X1 U15328 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n11167), .B2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12095) );
  NAND4_X1 U15329 ( .A1(n12098), .A2(n12097), .A3(n12096), .A4(n12095), .ZN(
        n12104) );
  AOI22_X1 U15330 ( .A1(n12466), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12102) );
  AOI22_X1 U15331 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12101) );
  AOI22_X1 U15332 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12100) );
  AOI22_X1 U15333 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12099) );
  NAND4_X1 U15334 ( .A1(n12102), .A2(n12101), .A3(n12100), .A4(n12099), .ZN(
        n12103) );
  OR2_X1 U15335 ( .A1(n12104), .A2(n12103), .ZN(n12105) );
  NAND2_X1 U15336 ( .A1(n14058), .A2(n14131), .ZN(n12106) );
  XNOR2_X1 U15337 ( .A(n12188), .B(n12187), .ZN(n14669) );
  AOI22_X1 U15338 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12440), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12110) );
  AOI22_X1 U15339 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11167), .B2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12109) );
  AOI22_X1 U15340 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12108) );
  AOI22_X1 U15341 ( .A1(n11152), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12107) );
  NAND4_X1 U15342 ( .A1(n12110), .A2(n12109), .A3(n12108), .A4(n12107), .ZN(
        n12116) );
  AOI22_X1 U15343 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n11146), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12114) );
  AOI22_X1 U15344 ( .A1(n12467), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12113) );
  AOI22_X1 U15345 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12299), .B2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12112) );
  AOI22_X1 U15346 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12111) );
  NAND4_X1 U15347 ( .A1(n12114), .A2(n12113), .A3(n12112), .A4(n12111), .ZN(
        n12115) );
  OAI21_X1 U15348 ( .B1(n12116), .B2(n12115), .A(n12130), .ZN(n12119) );
  NAND2_X1 U15349 ( .A1(n11999), .A2(P1_EAX_REG_15__SCAN_IN), .ZN(n12118) );
  NAND2_X1 U15350 ( .A1(n12485), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n12117) );
  NAND3_X1 U15351 ( .A1(n12119), .A2(n12118), .A3(n12117), .ZN(n12120) );
  AOI21_X1 U15352 ( .B1(n14669), .B2(n12452), .A(n12120), .ZN(n14150) );
  INV_X1 U15353 ( .A(n14150), .ZN(n12170) );
  XOR2_X1 U15354 ( .A(n15830), .B(n12121), .Z(n15880) );
  INV_X1 U15355 ( .A(n15880), .ZN(n12137) );
  AOI22_X1 U15356 ( .A1(n12458), .A2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n11146), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12125) );
  AOI22_X1 U15357 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n12440), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12124) );
  AOI22_X1 U15358 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12123) );
  AOI22_X1 U15359 ( .A1(n12460), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12122) );
  NAND4_X1 U15360 ( .A1(n12125), .A2(n12124), .A3(n12123), .A4(n12122), .ZN(
        n12132) );
  AOI22_X1 U15361 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n11167), .B2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12129) );
  AOI22_X1 U15362 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11047), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12128) );
  AOI22_X1 U15363 ( .A1(n12467), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n12468), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12127) );
  AOI22_X1 U15364 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12126) );
  NAND4_X1 U15365 ( .A1(n12129), .A2(n12128), .A3(n12127), .A4(n12126), .ZN(
        n12131) );
  OAI21_X1 U15366 ( .B1(n12132), .B2(n12131), .A(n12130), .ZN(n12135) );
  NAND2_X1 U15367 ( .A1(n11999), .A2(P1_EAX_REG_14__SCAN_IN), .ZN(n12134) );
  NAND2_X1 U15368 ( .A1(n12485), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(
        n12133) );
  NAND3_X1 U15369 ( .A1(n12135), .A2(n12134), .A3(n12133), .ZN(n12136) );
  AOI21_X1 U15370 ( .B1(n12137), .B2(n12452), .A(n12136), .ZN(n14142) );
  INV_X1 U15371 ( .A(n14142), .ZN(n12169) );
  AOI22_X1 U15372 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n9831), .B1(
        n12440), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12141) );
  AOI22_X1 U15373 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12140) );
  AOI22_X1 U15374 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11167), .B2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12139) );
  AOI22_X1 U15375 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12138) );
  NAND4_X1 U15376 ( .A1(n12141), .A2(n12140), .A3(n12139), .A4(n12138), .ZN(
        n12147) );
  AOI22_X1 U15377 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12458), .B1(
        n11146), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12145) );
  AOI22_X1 U15378 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n12144) );
  AOI22_X1 U15379 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12143) );
  AOI22_X1 U15380 ( .A1(n12467), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n12468), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12142) );
  NAND4_X1 U15381 ( .A1(n12145), .A2(n12144), .A3(n12143), .A4(n12142), .ZN(
        n12146) );
  NOR2_X1 U15382 ( .A1(n12147), .A2(n12146), .ZN(n12153) );
  XNOR2_X1 U15383 ( .A(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B(n12148), .ZN(
        n15886) );
  OAI22_X1 U15384 ( .A1(n15886), .A2(n12484), .B1(n12203), .B2(n12149), .ZN(
        n12150) );
  INV_X1 U15385 ( .A(n12150), .ZN(n12152) );
  NAND2_X1 U15386 ( .A1(n11999), .A2(P1_EAX_REG_12__SCAN_IN), .ZN(n12151) );
  OAI211_X1 U15387 ( .C1(n12168), .C2(n12153), .A(n12152), .B(n12151), .ZN(
        n14134) );
  AOI22_X1 U15388 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12157) );
  AOI22_X1 U15389 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12156) );
  AOI22_X1 U15390 ( .A1(n11167), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12155) );
  AOI22_X1 U15391 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12154) );
  NAND4_X1 U15392 ( .A1(n12157), .A2(n12156), .A3(n12155), .A4(n12154), .ZN(
        n12163) );
  AOI22_X1 U15393 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12161) );
  AOI22_X1 U15394 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12440), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12160) );
  AOI22_X1 U15395 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n12468), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12159) );
  AOI22_X1 U15396 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12158) );
  NAND4_X1 U15397 ( .A1(n12161), .A2(n12160), .A3(n12159), .A4(n12158), .ZN(
        n12162) );
  NOR2_X1 U15398 ( .A1(n12163), .A2(n12162), .ZN(n12167) );
  XNOR2_X1 U15399 ( .A(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B(n12164), .ZN(
        n14681) );
  AOI22_X1 U15400 ( .A1(n12452), .A2(n14681), .B1(n12485), .B2(
        P1_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n12166) );
  NAND2_X1 U15401 ( .A1(n11999), .A2(P1_EAX_REG_13__SCAN_IN), .ZN(n12165) );
  OAI211_X1 U15402 ( .C1(n12168), .C2(n12167), .A(n12166), .B(n12165), .ZN(
        n14156) );
  AND2_X1 U15403 ( .A1(n14134), .A2(n14156), .ZN(n14141) );
  AOI22_X1 U15404 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12458), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12176) );
  AOI22_X1 U15405 ( .A1(n12467), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12175) );
  AOI22_X1 U15406 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12299), .B2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12174) );
  AOI22_X1 U15407 ( .A1(n11167), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12173) );
  NAND4_X1 U15408 ( .A1(n12176), .A2(n12175), .A3(n12174), .A4(n12173), .ZN(
        n12182) );
  AOI22_X1 U15409 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12306), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12180) );
  AOI22_X1 U15410 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12179) );
  AOI22_X1 U15411 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12178) );
  AOI22_X1 U15412 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12177) );
  NAND4_X1 U15413 ( .A1(n12180), .A2(n12179), .A3(n12178), .A4(n12177), .ZN(
        n12181) );
  NOR2_X1 U15414 ( .A1(n12182), .A2(n12181), .ZN(n12186) );
  NAND2_X1 U15415 ( .A1(n20691), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n12183) );
  NAND2_X1 U15416 ( .A1(n12484), .A2(n12183), .ZN(n12184) );
  AOI21_X1 U15417 ( .B1(n12451), .B2(P1_EAX_REG_16__SCAN_IN), .A(n12184), .ZN(
        n12185) );
  OAI21_X1 U15418 ( .B1(n12481), .B2(n12186), .A(n12185), .ZN(n12191) );
  OAI21_X1 U15419 ( .B1(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n12189), .A(
        n12221), .ZN(n15879) );
  OR2_X1 U15420 ( .A1(n12484), .A2(n15879), .ZN(n12190) );
  NAND2_X1 U15421 ( .A1(n12191), .A2(n12190), .ZN(n14166) );
  AOI22_X1 U15422 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12458), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12195) );
  AOI22_X1 U15423 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12194) );
  AOI22_X1 U15424 ( .A1(n12467), .A2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12193) );
  AOI22_X1 U15425 ( .A1(n11152), .A2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n12192) );
  NAND4_X1 U15426 ( .A1(n12195), .A2(n12194), .A3(n12193), .A4(n12192), .ZN(
        n12201) );
  AOI22_X1 U15427 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n9831), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12199) );
  AOI22_X1 U15428 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11167), .B2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12198) );
  AOI22_X1 U15429 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12197) );
  AOI22_X1 U15430 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12196) );
  NAND4_X1 U15431 ( .A1(n12199), .A2(n12198), .A3(n12197), .A4(n12196), .ZN(
        n12200) );
  OR2_X1 U15432 ( .A1(n12201), .A2(n12200), .ZN(n12202) );
  NAND2_X1 U15433 ( .A1(n12447), .A2(n12202), .ZN(n12206) );
  XNOR2_X1 U15434 ( .A(P1_PHYADDRPOINTER_REG_17__SCAN_IN), .B(n12221), .ZN(
        n15813) );
  OAI22_X1 U15435 ( .A1(n15813), .A2(n12484), .B1(n12203), .B2(n15810), .ZN(
        n12204) );
  AOI21_X1 U15436 ( .B1(n12451), .B2(P1_EAX_REG_17__SCAN_IN), .A(n12204), .ZN(
        n12205) );
  NAND2_X1 U15437 ( .A1(n12206), .A2(n12205), .ZN(n14206) );
  AOI22_X1 U15438 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12210) );
  AOI22_X1 U15439 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12209) );
  AOI22_X1 U15440 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12208) );
  AOI22_X1 U15441 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12207) );
  NAND4_X1 U15442 ( .A1(n12210), .A2(n12209), .A3(n12208), .A4(n12207), .ZN(
        n12216) );
  AOI22_X1 U15443 ( .A1(n12458), .A2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n11146), .B2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12214) );
  AOI22_X1 U15444 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12306), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12213) );
  AOI22_X1 U15445 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n12212) );
  AOI22_X1 U15446 ( .A1(n11167), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12211) );
  NAND4_X1 U15447 ( .A1(n12214), .A2(n12213), .A3(n12212), .A4(n12211), .ZN(
        n12215) );
  NOR2_X1 U15448 ( .A1(n12216), .A2(n12215), .ZN(n12220) );
  NAND2_X1 U15449 ( .A1(n20691), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n12217) );
  NAND2_X1 U15450 ( .A1(n12484), .A2(n12217), .ZN(n12218) );
  AOI21_X1 U15451 ( .B1(n12451), .B2(P1_EAX_REG_18__SCAN_IN), .A(n12218), .ZN(
        n12219) );
  OAI21_X1 U15452 ( .B1(n12481), .B2(n12220), .A(n12219), .ZN(n12224) );
  OAI21_X1 U15453 ( .B1(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n12222), .A(
        n12238), .ZN(n14647) );
  OR2_X1 U15454 ( .A1(n12484), .A2(n14647), .ZN(n12223) );
  NAND2_X1 U15455 ( .A1(n12224), .A2(n12223), .ZN(n14388) );
  AOI22_X1 U15456 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12458), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12228) );
  AOI22_X1 U15457 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n11167), .B2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12227) );
  AOI22_X1 U15458 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12306), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12226) );
  AOI22_X1 U15459 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n12225) );
  NAND4_X1 U15460 ( .A1(n12228), .A2(n12227), .A3(n12226), .A4(n12225), .ZN(
        n12234) );
  AOI22_X1 U15461 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12232) );
  AOI22_X1 U15462 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12231) );
  AOI22_X1 U15463 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n12468), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12230) );
  AOI22_X1 U15464 ( .A1(n11152), .A2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12229) );
  NAND4_X1 U15465 ( .A1(n12232), .A2(n12231), .A3(n12230), .A4(n12229), .ZN(
        n12233) );
  NOR2_X1 U15466 ( .A1(n12234), .A2(n12233), .ZN(n12237) );
  INV_X1 U15467 ( .A(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n21101) );
  OAI21_X1 U15468 ( .B1(P1_STATE2_REG_2__SCAN_IN), .B2(n21101), .A(n12484), 
        .ZN(n12235) );
  AOI21_X1 U15469 ( .B1(n12451), .B2(P1_EAX_REG_19__SCAN_IN), .A(n12235), .ZN(
        n12236) );
  OAI21_X1 U15470 ( .B1(n12481), .B2(n12237), .A(n12236), .ZN(n12242) );
  INV_X1 U15471 ( .A(n12238), .ZN(n12240) );
  INV_X1 U15472 ( .A(n12257), .ZN(n12239) );
  OAI21_X1 U15473 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n12240), .A(
        n12239), .ZN(n14640) );
  OR2_X1 U15474 ( .A1(n12484), .A2(n14640), .ZN(n12241) );
  NAND2_X1 U15475 ( .A1(n12242), .A2(n12241), .ZN(n14374) );
  AOI22_X1 U15476 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .B1(
        n11146), .B2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n12246) );
  AOI22_X1 U15477 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .B1(
        n11167), .B2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12245) );
  AOI22_X1 U15478 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n12466), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12244) );
  AOI22_X1 U15479 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12243) );
  NAND4_X1 U15480 ( .A1(n12246), .A2(n12245), .A3(n12244), .A4(n12243), .ZN(
        n12252) );
  AOI22_X1 U15481 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12250) );
  AOI22_X1 U15482 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12299), .B2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12249) );
  AOI22_X1 U15483 ( .A1(n12458), .A2(P1_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n12468), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12248) );
  AOI22_X1 U15484 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12247) );
  NAND4_X1 U15485 ( .A1(n12250), .A2(n12249), .A3(n12248), .A4(n12247), .ZN(
        n12251) );
  NOR2_X1 U15486 ( .A1(n12252), .A2(n12251), .ZN(n12256) );
  INV_X1 U15487 ( .A(P1_STATEBS16_REG_SCAN_IN), .ZN(n20765) );
  OAI21_X1 U15488 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n20765), .A(
        n20691), .ZN(n12253) );
  INV_X1 U15489 ( .A(n12253), .ZN(n12254) );
  AOI21_X1 U15490 ( .B1(n12451), .B2(P1_EAX_REG_20__SCAN_IN), .A(n12254), .ZN(
        n12255) );
  OAI21_X1 U15491 ( .B1(n12481), .B2(n12256), .A(n12255), .ZN(n12259) );
  OAI21_X1 U15492 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n12257), .A(
        n12290), .ZN(n15866) );
  OR2_X1 U15493 ( .A1(n12484), .A2(n15866), .ZN(n12258) );
  AOI22_X1 U15494 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n11146), .B2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12263) );
  AOI22_X1 U15495 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n11167), .B2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12262) );
  AOI22_X1 U15496 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n12261) );
  AOI22_X1 U15497 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12260) );
  NAND4_X1 U15498 ( .A1(n12263), .A2(n12262), .A3(n12261), .A4(n12260), .ZN(
        n12269) );
  AOI22_X1 U15499 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12267) );
  AOI22_X1 U15500 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12299), .B2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12266) );
  AOI22_X1 U15501 ( .A1(n12458), .A2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12468), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12265) );
  AOI22_X1 U15502 ( .A1(n12466), .A2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12264) );
  NAND4_X1 U15503 ( .A1(n12267), .A2(n12266), .A3(n12265), .A4(n12264), .ZN(
        n12268) );
  NOR2_X1 U15504 ( .A1(n12269), .A2(n12268), .ZN(n12272) );
  INV_X1 U15505 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n15802) );
  AOI21_X1 U15506 ( .B1(P1_STATEBS16_REG_SCAN_IN), .B2(n15802), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12270) );
  AOI21_X1 U15507 ( .B1(n12451), .B2(P1_EAX_REG_21__SCAN_IN), .A(n12270), .ZN(
        n12271) );
  OAI21_X1 U15508 ( .B1(n12481), .B2(n12272), .A(n12271), .ZN(n12274) );
  XNOR2_X1 U15509 ( .A(P1_PHYADDRPOINTER_REG_21__SCAN_IN), .B(n12290), .ZN(
        n15799) );
  NAND2_X1 U15510 ( .A1(n15799), .A2(n12452), .ZN(n12273) );
  NAND2_X1 U15511 ( .A1(n14486), .A2(n14488), .ZN(n14478) );
  AOI22_X1 U15512 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12279) );
  AOI22_X1 U15513 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12278) );
  AOI22_X1 U15514 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .B1(
        n11167), .B2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12277) );
  AOI22_X1 U15515 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12276) );
  NAND4_X1 U15516 ( .A1(n12279), .A2(n12278), .A3(n12277), .A4(n12276), .ZN(
        n12285) );
  AOI22_X1 U15517 ( .A1(n12458), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n11146), .B2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n12283) );
  AOI22_X1 U15518 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12282) );
  AOI22_X1 U15519 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12281) );
  AOI22_X1 U15520 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12280) );
  NAND4_X1 U15521 ( .A1(n12283), .A2(n12282), .A3(n12281), .A4(n12280), .ZN(
        n12284) );
  NOR2_X1 U15522 ( .A1(n12285), .A2(n12284), .ZN(n12289) );
  NAND2_X1 U15523 ( .A1(n20691), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n12286) );
  NAND2_X1 U15524 ( .A1(n12484), .A2(n12286), .ZN(n12287) );
  AOI21_X1 U15525 ( .B1(n12451), .B2(P1_EAX_REG_22__SCAN_IN), .A(n12287), .ZN(
        n12288) );
  OAI21_X1 U15526 ( .B1(n12481), .B2(n12289), .A(n12288), .ZN(n12293) );
  OAI21_X1 U15527 ( .B1(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n12291), .A(
        n12340), .ZN(n15865) );
  OR2_X1 U15528 ( .A1(n12484), .A2(n15865), .ZN(n12292) );
  NAND2_X1 U15529 ( .A1(n12293), .A2(n12292), .ZN(n14479) );
  NOR2_X2 U15530 ( .A1(n14478), .A2(n14479), .ZN(n14470) );
  AOI22_X1 U15531 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n11146), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12298) );
  AOI22_X1 U15532 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12297) );
  AOI22_X1 U15533 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n12296) );
  AOI22_X1 U15534 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n12295) );
  NAND4_X1 U15535 ( .A1(n12298), .A2(n12297), .A3(n12296), .A4(n12295), .ZN(
        n12305) );
  AOI22_X1 U15536 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n11167), .B2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12303) );
  AOI22_X1 U15537 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12302) );
  AOI22_X1 U15538 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12301) );
  AOI22_X1 U15539 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12300) );
  NAND4_X1 U15540 ( .A1(n12303), .A2(n12302), .A3(n12301), .A4(n12300), .ZN(
        n12304) );
  NOR2_X1 U15541 ( .A1(n12305), .A2(n12304), .ZN(n12324) );
  AOI22_X1 U15542 ( .A1(n12458), .A2(P1_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n11146), .B2(P1_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12310) );
  AOI22_X1 U15543 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n12309) );
  AOI22_X1 U15544 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12306), .B2(P1_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12308) );
  AOI22_X1 U15545 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12307) );
  NAND4_X1 U15546 ( .A1(n12310), .A2(n12309), .A3(n12308), .A4(n12307), .ZN(
        n12316) );
  AOI22_X1 U15547 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n12314) );
  AOI22_X1 U15548 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12313) );
  AOI22_X1 U15549 ( .A1(n11167), .A2(P1_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12312) );
  AOI22_X1 U15550 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n12311) );
  NAND4_X1 U15551 ( .A1(n12314), .A2(n12313), .A3(n12312), .A4(n12311), .ZN(
        n12315) );
  NOR2_X1 U15552 ( .A1(n12316), .A2(n12315), .ZN(n12325) );
  XOR2_X1 U15553 ( .A(n12324), .B(n12325), .Z(n12317) );
  NAND2_X1 U15554 ( .A1(n12317), .A2(n12447), .ZN(n12321) );
  NAND2_X1 U15555 ( .A1(n20691), .A2(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n12318) );
  NAND2_X1 U15556 ( .A1(n12484), .A2(n12318), .ZN(n12319) );
  AOI21_X1 U15557 ( .B1(n12451), .B2(P1_EAX_REG_23__SCAN_IN), .A(n12319), .ZN(
        n12320) );
  NAND2_X1 U15558 ( .A1(n12321), .A2(n12320), .ZN(n12323) );
  XNOR2_X1 U15559 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B(n12340), .ZN(
        n15774) );
  NAND2_X1 U15560 ( .A1(n15774), .A2(n12452), .ZN(n12322) );
  AND2_X2 U15561 ( .A1(n14470), .A2(n10306), .ZN(n14463) );
  NOR2_X1 U15562 ( .A1(n12325), .A2(n12324), .ZN(n12350) );
  AOI22_X1 U15563 ( .A1(n12458), .A2(P1_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n11146), .B2(P1_INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n12329) );
  AOI22_X1 U15564 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n12328) );
  AOI22_X1 U15565 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12327) );
  AOI22_X1 U15566 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        n12468), .B2(P1_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n12326) );
  NAND4_X1 U15567 ( .A1(n12329), .A2(n12328), .A3(n12327), .A4(n12326), .ZN(
        n12335) );
  AOI22_X1 U15568 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_1__1__SCAN_IN), .B1(
        n11167), .B2(P1_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12333) );
  AOI22_X1 U15569 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_15__1__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n12332) );
  AOI22_X1 U15570 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12331) );
  AOI22_X1 U15571 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12330) );
  NAND4_X1 U15572 ( .A1(n12333), .A2(n12332), .A3(n12331), .A4(n12330), .ZN(
        n12334) );
  OR2_X1 U15573 ( .A1(n12335), .A2(n12334), .ZN(n12349) );
  INV_X1 U15574 ( .A(n12349), .ZN(n12336) );
  XNOR2_X1 U15575 ( .A(n12350), .B(n12336), .ZN(n12337) );
  NAND2_X1 U15576 ( .A1(n12337), .A2(n12447), .ZN(n12348) );
  NAND2_X1 U15577 ( .A1(n20691), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n12338) );
  NAND2_X1 U15578 ( .A1(n12484), .A2(n12338), .ZN(n12339) );
  AOI21_X1 U15579 ( .B1(n12451), .B2(P1_EAX_REG_24__SCAN_IN), .A(n12339), .ZN(
        n12347) );
  INV_X1 U15580 ( .A(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n12344) );
  INV_X1 U15581 ( .A(n12342), .ZN(n12343) );
  NAND2_X1 U15582 ( .A1(n12344), .A2(n12343), .ZN(n12345) );
  NAND2_X1 U15583 ( .A1(n12383), .A2(n12345), .ZN(n15769) );
  NOR2_X1 U15584 ( .A1(n15769), .A2(n12484), .ZN(n12346) );
  AOI21_X1 U15585 ( .B1(n12348), .B2(n12347), .A(n12346), .ZN(n14462) );
  NAND2_X1 U15586 ( .A1(n12350), .A2(n12349), .ZN(n12367) );
  AOI22_X1 U15587 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12354) );
  AOI22_X1 U15588 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n12459), .B2(P1_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12353) );
  AOI22_X1 U15589 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n12299), .B2(P1_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12352) );
  AOI22_X1 U15590 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n12294), .B2(P1_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n12351) );
  NAND4_X1 U15591 ( .A1(n12354), .A2(n12353), .A3(n12352), .A4(n12351), .ZN(
        n12360) );
  AOI22_X1 U15592 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n12458), .B2(P1_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12358) );
  AOI22_X1 U15593 ( .A1(n12467), .A2(P1_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n12357) );
  AOI22_X1 U15594 ( .A1(n11167), .A2(P1_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12356) );
  AOI22_X1 U15595 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12355) );
  NAND4_X1 U15596 ( .A1(n12358), .A2(n12357), .A3(n12356), .A4(n12355), .ZN(
        n12359) );
  NOR2_X1 U15597 ( .A1(n12360), .A2(n12359), .ZN(n12368) );
  XOR2_X1 U15598 ( .A(n12367), .B(n12368), .Z(n12361) );
  NAND2_X1 U15599 ( .A1(n12361), .A2(n12447), .ZN(n12366) );
  NAND2_X1 U15600 ( .A1(n20691), .A2(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n12362) );
  NAND2_X1 U15601 ( .A1(n12484), .A2(n12362), .ZN(n12363) );
  AOI21_X1 U15602 ( .B1(n12451), .B2(P1_EAX_REG_25__SCAN_IN), .A(n12363), .ZN(
        n12365) );
  XNOR2_X1 U15603 ( .A(n12383), .B(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15754) );
  AOI21_X1 U15604 ( .B1(n12366), .B2(n12365), .A(n12364), .ZN(n14454) );
  NOR2_X1 U15605 ( .A1(n12368), .A2(n12367), .ZN(n12391) );
  AOI22_X1 U15606 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n11146), .B2(P1_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n12372) );
  AOI22_X1 U15607 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n12371) );
  AOI22_X1 U15608 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12370) );
  AOI22_X1 U15609 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n12468), .B2(P1_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n12369) );
  NAND4_X1 U15610 ( .A1(n12372), .A2(n12371), .A3(n12370), .A4(n12369), .ZN(
        n12378) );
  AOI22_X1 U15611 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_1__3__SCAN_IN), .B1(
        n11167), .B2(P1_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12376) );
  AOI22_X1 U15612 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n12375) );
  AOI22_X1 U15613 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12374) );
  AOI22_X1 U15614 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12373) );
  NAND4_X1 U15615 ( .A1(n12376), .A2(n12375), .A3(n12374), .A4(n12373), .ZN(
        n12377) );
  OR2_X1 U15616 ( .A1(n12378), .A2(n12377), .ZN(n12390) );
  INV_X1 U15617 ( .A(n12390), .ZN(n12379) );
  XNOR2_X1 U15618 ( .A(n12391), .B(n12379), .ZN(n12382) );
  INV_X1 U15619 ( .A(P1_EAX_REG_26__SCAN_IN), .ZN(n14521) );
  NAND2_X1 U15620 ( .A1(n20691), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n12380) );
  OAI211_X1 U15621 ( .C1(n12424), .C2(n14521), .A(n12484), .B(n12380), .ZN(
        n12381) );
  AOI21_X1 U15622 ( .B1(n12382), .B2(n12447), .A(n12381), .ZN(n12389) );
  INV_X1 U15623 ( .A(P1_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n15748) );
  INV_X1 U15624 ( .A(n12384), .ZN(n12386) );
  INV_X1 U15625 ( .A(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n12385) );
  NAND2_X1 U15626 ( .A1(n12386), .A2(n12385), .ZN(n12387) );
  NAND2_X1 U15627 ( .A1(n12427), .A2(n12387), .ZN(n14607) );
  NOR2_X1 U15628 ( .A1(n14607), .A2(n12484), .ZN(n12388) );
  NAND2_X1 U15629 ( .A1(n12391), .A2(n12390), .ZN(n12410) );
  AOI22_X1 U15630 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n9831), .B1(
        n12299), .B2(P1_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12395) );
  AOI22_X1 U15631 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n11167), .B2(P1_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12394) );
  AOI22_X1 U15632 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n12468), .B2(P1_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n12393) );
  AOI22_X1 U15633 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12392) );
  NAND4_X1 U15634 ( .A1(n12395), .A2(n12394), .A3(n12393), .A4(n12392), .ZN(
        n12401) );
  AOI22_X1 U15635 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n11146), .B2(P1_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n12399) );
  AOI22_X1 U15636 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n12466), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12398) );
  AOI22_X1 U15637 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n12397) );
  AOI22_X1 U15638 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n12396) );
  NAND4_X1 U15639 ( .A1(n12399), .A2(n12398), .A3(n12397), .A4(n12396), .ZN(
        n12400) );
  NOR2_X1 U15640 ( .A1(n12401), .A2(n12400), .ZN(n12411) );
  XOR2_X1 U15641 ( .A(n12410), .B(n12411), .Z(n12402) );
  NAND2_X1 U15642 ( .A1(n12402), .A2(n12447), .ZN(n12406) );
  INV_X1 U15643 ( .A(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n12403) );
  AOI21_X1 U15644 ( .B1(n12403), .B2(P1_STATEBS16_REG_SCAN_IN), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n12404) );
  AOI21_X1 U15645 ( .B1(n12451), .B2(P1_EAX_REG_27__SCAN_IN), .A(n12404), .ZN(
        n12405) );
  NAND2_X1 U15646 ( .A1(n12406), .A2(n12405), .ZN(n12408) );
  XNOR2_X1 U15647 ( .A(n12427), .B(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14594) );
  NAND2_X1 U15648 ( .A1(n14594), .A2(n12452), .ZN(n12407) );
  NAND2_X1 U15649 ( .A1(n12408), .A2(n12407), .ZN(n14352) );
  NOR2_X1 U15650 ( .A1(n12411), .A2(n12410), .ZN(n12435) );
  AOI22_X1 U15651 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n11146), .B2(P1_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12415) );
  AOI22_X1 U15652 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n12467), .B2(P1_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n12414) );
  AOI22_X1 U15653 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n12413) );
  AOI22_X1 U15654 ( .A1(n12440), .A2(P1_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n12468), .B2(P1_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n12412) );
  NAND4_X1 U15655 ( .A1(n12415), .A2(n12414), .A3(n12413), .A4(n12412), .ZN(
        n12421) );
  AOI22_X1 U15656 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_1__5__SCAN_IN), .B1(
        n11167), .B2(P1_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12419) );
  AOI22_X1 U15657 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n12418) );
  AOI22_X1 U15658 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12417) );
  AOI22_X1 U15659 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12416) );
  NAND4_X1 U15660 ( .A1(n12419), .A2(n12418), .A3(n12417), .A4(n12416), .ZN(
        n12420) );
  OR2_X1 U15661 ( .A1(n12421), .A2(n12420), .ZN(n12434) );
  INV_X1 U15662 ( .A(n12434), .ZN(n12422) );
  XNOR2_X1 U15663 ( .A(n12435), .B(n12422), .ZN(n12426) );
  INV_X1 U15664 ( .A(P1_EAX_REG_28__SCAN_IN), .ZN(n14512) );
  NAND2_X1 U15665 ( .A1(n20691), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n12423) );
  OAI211_X1 U15666 ( .C1(n12424), .C2(n14512), .A(n12484), .B(n12423), .ZN(
        n12425) );
  AOI21_X1 U15667 ( .B1(n12426), .B2(n12447), .A(n12425), .ZN(n12433) );
  INV_X1 U15668 ( .A(n12427), .ZN(n12428) );
  INV_X1 U15669 ( .A(n12429), .ZN(n12430) );
  INV_X1 U15670 ( .A(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n14340) );
  NAND2_X1 U15671 ( .A1(n12430), .A2(n14340), .ZN(n12431) );
  NAND2_X1 U15672 ( .A1(n12456), .A2(n12431), .ZN(n14584) );
  NOR2_X1 U15673 ( .A1(n14584), .A2(n12484), .ZN(n12432) );
  NAND2_X1 U15674 ( .A1(n12435), .A2(n12434), .ZN(n12475) );
  AOI22_X1 U15675 ( .A1(n11110), .A2(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n11146), .B2(P1_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n12439) );
  AOI22_X1 U15676 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n12299), .B2(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12438) );
  AOI22_X1 U15677 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n11167), .B2(P1_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12437) );
  AOI22_X1 U15678 ( .A1(n12466), .A2(P1_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n12468), .B2(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n12436) );
  NAND4_X1 U15679 ( .A1(n12439), .A2(n12438), .A3(n12437), .A4(n12436), .ZN(
        n12446) );
  AOI22_X1 U15680 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n12440), .B2(P1_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12444) );
  AOI22_X1 U15681 ( .A1(n12467), .A2(P1_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n11152), .B2(P1_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n12443) );
  AOI22_X1 U15682 ( .A1(n12306), .A2(P1_INSTQUEUE_REG_1__6__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n12442) );
  AOI22_X1 U15683 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12441) );
  NAND4_X1 U15684 ( .A1(n12444), .A2(n12443), .A3(n12442), .A4(n12441), .ZN(
        n12445) );
  NOR2_X1 U15685 ( .A1(n12446), .A2(n12445), .ZN(n12476) );
  XOR2_X1 U15686 ( .A(n12475), .B(n12476), .Z(n12448) );
  NAND2_X1 U15687 ( .A1(n12448), .A2(n12447), .ZN(n12455) );
  NAND2_X1 U15688 ( .A1(n20691), .A2(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n12449) );
  NAND2_X1 U15689 ( .A1(n12484), .A2(n12449), .ZN(n12450) );
  AOI21_X1 U15690 ( .B1(n12451), .B2(P1_EAX_REG_29__SCAN_IN), .A(n12450), .ZN(
        n12454) );
  XNOR2_X1 U15691 ( .A(n12456), .B(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14312) );
  AOI21_X1 U15692 ( .B1(n12455), .B2(n12454), .A(n12453), .ZN(n14300) );
  INV_X1 U15693 ( .A(n12456), .ZN(n12457) );
  XNOR2_X1 U15694 ( .A(n12490), .B(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n14570) );
  AOI22_X1 U15695 ( .A1(n12275), .A2(P1_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n12458), .B2(P1_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12464) );
  AOI22_X1 U15696 ( .A1(n11154), .A2(P1_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n11167), .B2(P1_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12463) );
  AOI22_X1 U15697 ( .A1(n12459), .A2(P1_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n11047), .B2(P1_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n12462) );
  AOI22_X1 U15698 ( .A1(n11152), .A2(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n12460), .B2(P1_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12461) );
  NAND4_X1 U15699 ( .A1(n12464), .A2(n12463), .A3(n12462), .A4(n12461), .ZN(
        n12474) );
  AOI22_X1 U15700 ( .A1(n9831), .A2(P1_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n12440), .B2(P1_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12472) );
  AOI22_X1 U15701 ( .A1(n12467), .A2(P1_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n12466), .B2(P1_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12471) );
  AOI22_X1 U15702 ( .A1(n11146), .A2(P1_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n12468), .B2(P1_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n12470) );
  AOI22_X1 U15703 ( .A1(n12299), .A2(P1_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n11155), .B2(P1_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12469) );
  NAND4_X1 U15704 ( .A1(n12472), .A2(n12471), .A3(n12470), .A4(n12469), .ZN(
        n12473) );
  NOR2_X1 U15705 ( .A1(n12474), .A2(n12473), .ZN(n12478) );
  NOR2_X1 U15706 ( .A1(n12476), .A2(n12475), .ZN(n12477) );
  XOR2_X1 U15707 ( .A(n12478), .B(n12477), .Z(n12482) );
  AOI21_X1 U15708 ( .B1(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n20691), .A(
        n12452), .ZN(n12480) );
  NAND2_X1 U15709 ( .A1(n12451), .A2(P1_EAX_REG_30__SCAN_IN), .ZN(n12479) );
  OAI211_X1 U15710 ( .C1(n12482), .C2(n12481), .A(n12480), .B(n12479), .ZN(
        n12483) );
  OAI21_X1 U15711 ( .B1(n12484), .B2(n14570), .A(n12483), .ZN(n14323) );
  AOI22_X1 U15712 ( .A1(n12451), .A2(P1_EAX_REG_31__SCAN_IN), .B1(n12485), 
        .B2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12486) );
  NAND2_X1 U15713 ( .A1(n13472), .A2(n11470), .ZN(n13263) );
  INV_X1 U15714 ( .A(n13520), .ZN(n19857) );
  INV_X1 U15715 ( .A(P1_STATE2_REG_3__SCAN_IN), .ZN(n20388) );
  NAND2_X1 U15716 ( .A1(n20691), .A2(n16000), .ZN(n15723) );
  OR2_X1 U15717 ( .A1(n20388), .A2(n15723), .ZN(n15718) );
  NOR2_X1 U15718 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n16000), .ZN(n15725) );
  NAND2_X1 U15719 ( .A1(n12452), .A2(n15725), .ZN(n12487) );
  OAI211_X1 U15720 ( .C1(n15718), .C2(n11192), .A(n20046), .B(n12487), .ZN(
        n12488) );
  INV_X1 U15721 ( .A(n12488), .ZN(n12489) );
  INV_X1 U15722 ( .A(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n12513) );
  NAND2_X1 U15723 ( .A1(n14504), .A2(n19908), .ZN(n12520) );
  MUX2_X1 U15724 ( .A(n12494), .B(n12493), .S(n14310), .Z(n12497) );
  AOI22_X1 U15725 ( .A1(n12495), .A2(P1_EBX_REG_31__SCAN_IN), .B1(
        P1_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n13516), .ZN(n12496) );
  OR2_X1 U15726 ( .A1(n20789), .A2(n12498), .ZN(n12507) );
  AND2_X1 U15727 ( .A1(n20122), .A2(P1_EBX_REG_31__SCAN_IN), .ZN(n12508) );
  NAND2_X1 U15728 ( .A1(n15993), .A2(n20765), .ZN(n12500) );
  NAND2_X1 U15729 ( .A1(n12508), .A2(n12500), .ZN(n12499) );
  NOR2_X2 U15730 ( .A1(n12507), .A2(n12499), .ZN(n19951) );
  AND2_X1 U15731 ( .A1(P1_REIP_REG_29__SCAN_IN), .A2(P1_REIP_REG_30__SCAN_IN), 
        .ZN(n12506) );
  INV_X1 U15732 ( .A(n12500), .ZN(n12501) );
  NAND2_X1 U15733 ( .A1(n12502), .A2(n12501), .ZN(n12509) );
  INV_X1 U15734 ( .A(n15781), .ZN(n19892) );
  INV_X1 U15735 ( .A(P1_REIP_REG_24__SCAN_IN), .ZN(n20739) );
  INV_X1 U15736 ( .A(P1_REIP_REG_19__SCAN_IN), .ZN(n14379) );
  INV_X1 U15737 ( .A(P1_REIP_REG_18__SCAN_IN), .ZN(n20729) );
  NAND4_X1 U15738 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_4__SCAN_IN), 
        .A3(P1_REIP_REG_3__SCAN_IN), .A4(P1_REIP_REG_2__SCAN_IN), .ZN(n14192)
         );
  NAND4_X1 U15739 ( .A1(P1_REIP_REG_14__SCAN_IN), .A2(P1_REIP_REG_13__SCAN_IN), 
        .A3(P1_REIP_REG_12__SCAN_IN), .A4(P1_REIP_REG_11__SCAN_IN), .ZN(n14400) );
  NAND4_X1 U15740 ( .A1(P1_REIP_REG_6__SCAN_IN), .A2(P1_REIP_REG_5__SCAN_IN), 
        .A3(P1_REIP_REG_8__SCAN_IN), .A4(P1_REIP_REG_7__SCAN_IN), .ZN(n14191)
         );
  NAND2_X1 U15741 ( .A1(P1_REIP_REG_16__SCAN_IN), .A2(P1_REIP_REG_15__SCAN_IN), 
        .ZN(n15814) );
  NOR4_X1 U15742 ( .A1(n14192), .A2(n14400), .A3(n14191), .A4(n15814), .ZN(
        n12503) );
  NAND4_X1 U15743 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(P1_REIP_REG_10__SCAN_IN), 
        .A3(P1_REIP_REG_9__SCAN_IN), .A4(n12503), .ZN(n14375) );
  NOR3_X1 U15744 ( .A1(n14379), .A2(n20729), .A3(n14375), .ZN(n15779) );
  INV_X1 U15745 ( .A(P1_REIP_REG_22__SCAN_IN), .ZN(n20736) );
  NAND2_X1 U15746 ( .A1(P1_REIP_REG_21__SCAN_IN), .A2(P1_REIP_REG_20__SCAN_IN), 
        .ZN(n15782) );
  NOR2_X1 U15747 ( .A1(n20736), .A2(n15782), .ZN(n15770) );
  NAND3_X1 U15748 ( .A1(P1_REIP_REG_23__SCAN_IN), .A2(n15779), .A3(n15770), 
        .ZN(n15761) );
  NOR2_X1 U15749 ( .A1(n20739), .A2(n15761), .ZN(n12514) );
  AND3_X1 U15750 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(P1_REIP_REG_26__SCAN_IN), 
        .A3(n12514), .ZN(n12504) );
  NAND2_X1 U15751 ( .A1(n14430), .A2(n12504), .ZN(n14353) );
  NAND2_X1 U15752 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(P1_REIP_REG_27__SCAN_IN), 
        .ZN(n12505) );
  INV_X1 U15753 ( .A(n14430), .ZN(n15780) );
  OR2_X1 U15754 ( .A1(n15781), .A2(n15780), .ZN(n19952) );
  OAI21_X1 U15755 ( .B1(n14353), .B2(n12505), .A(n19952), .ZN(n14342) );
  OAI21_X1 U15756 ( .B1(n12506), .B2(n19892), .A(n14342), .ZN(n14330) );
  INV_X1 U15757 ( .A(n12507), .ZN(n12512) );
  INV_X1 U15758 ( .A(n12508), .ZN(n12510) );
  AND2_X1 U15759 ( .A1(n12510), .A2(n12509), .ZN(n12511) );
  INV_X1 U15760 ( .A(P1_EBX_REG_31__SCAN_IN), .ZN(n14446) );
  OAI22_X1 U15761 ( .A1(n19934), .A2(n14446), .B1(n12513), .B2(n19954), .ZN(
        n12516) );
  AND2_X1 U15762 ( .A1(n15781), .A2(n12514), .ZN(n15753) );
  NAND2_X1 U15763 ( .A1(P1_REIP_REG_25__SCAN_IN), .A2(n15753), .ZN(n14364) );
  INV_X1 U15764 ( .A(P1_REIP_REG_26__SCAN_IN), .ZN(n15925) );
  INV_X1 U15765 ( .A(P1_REIP_REG_27__SCAN_IN), .ZN(n14595) );
  NOR3_X1 U15766 ( .A1(n14364), .A2(n15925), .A3(n14595), .ZN(n14341) );
  NAND2_X1 U15767 ( .A1(n14341), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14326) );
  INV_X1 U15768 ( .A(P1_REIP_REG_29__SCAN_IN), .ZN(n14325) );
  NOR4_X1 U15769 ( .A1(n14326), .A2(P1_REIP_REG_31__SCAN_IN), .A3(n14325), 
        .A4(n14324), .ZN(n12515) );
  AOI211_X1 U15770 ( .C1(P1_REIP_REG_31__SCAN_IN), .C2(n14330), .A(n12516), 
        .B(n12515), .ZN(n12517) );
  NAND2_X1 U15771 ( .A1(n12520), .A2(n12519), .ZN(P1_U2809) );
  INV_X1 U15772 ( .A(n14447), .ZN(n12530) );
  NAND2_X1 U15773 ( .A1(n12524), .A2(P1_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12527) );
  NAND3_X1 U15774 ( .A1(n12525), .A2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .A3(
        n14707), .ZN(n12526) );
  INV_X2 U15775 ( .A(n20046), .ZN(n15986) );
  NAND2_X1 U15776 ( .A1(n15986), .A2(P1_REIP_REG_31__SCAN_IN), .ZN(n14256) );
  OAI211_X1 U15777 ( .C1(n12528), .C2(n12527), .A(n12526), .B(n14256), .ZN(
        n12529) );
  AOI21_X1 U15778 ( .B1(n12530), .B2(n20089), .A(n12529), .ZN(n12531) );
  OAI21_X1 U15779 ( .B1(n14260), .B2(n20095), .A(n12531), .ZN(P1_U3000) );
  NAND2_X1 U15780 ( .A1(n12553), .A2(n12550), .ZN(n12542) );
  INV_X1 U15781 ( .A(n12534), .ZN(n12537) );
  INV_X1 U15782 ( .A(n12535), .ZN(n12536) );
  NAND2_X1 U15783 ( .A1(n19134), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n12538) );
  XNOR2_X1 U15784 ( .A(n12554), .B(n12538), .ZN(n16016) );
  AOI21_X1 U15785 ( .B1(n16016), .B2(n15187), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12552) );
  AND2_X1 U15786 ( .A1(n15187), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12539) );
  NAND2_X1 U15787 ( .A1(n16016), .A2(n12539), .ZN(n12551) );
  INV_X1 U15788 ( .A(n12551), .ZN(n12540) );
  NOR2_X1 U15789 ( .A1(n12552), .A2(n12540), .ZN(n12541) );
  XNOR2_X1 U15790 ( .A(n12542), .B(n12541), .ZN(n14279) );
  INV_X1 U15791 ( .A(P2_REIP_REG_30__SCAN_IN), .ZN(n12844) );
  NAND2_X1 U15792 ( .A1(n12543), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n12545) );
  AOI22_X1 U15793 ( .A1(n12622), .A2(P2_EBX_REG_30__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), 
        .ZN(n12544) );
  OAI211_X1 U15794 ( .C1(n9847), .C2(n12844), .A(n12545), .B(n12544), .ZN(
        n12621) );
  XNOR2_X1 U15795 ( .A(n13228), .B(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16021) );
  NOR2_X1 U15796 ( .A1(n18934), .A2(n12844), .ZN(n14271) );
  AOI21_X1 U15797 ( .B1(n19086), .B2(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14271), .ZN(n12546) );
  OAI21_X1 U15798 ( .B1(n16021), .B2(n19098), .A(n12546), .ZN(n12547) );
  OAI211_X1 U15799 ( .C1(n14279), .C2(n19108), .A(n12549), .B(n10289), .ZN(
        P2_U2984) );
  OAI21_X1 U15800 ( .B1(n12554), .B2(P2_EBX_REG_30__SCAN_IN), .A(n19134), .ZN(
        n12556) );
  NAND2_X1 U15801 ( .A1(n12556), .A2(n12555), .ZN(n16010) );
  NOR2_X1 U15802 ( .A1(n16010), .A2(n15176), .ZN(n12557) );
  XOR2_X1 U15803 ( .A(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B(n12557), .Z(
        n12558) );
  XNOR2_X1 U15804 ( .A(n12559), .B(n12558), .ZN(n14295) );
  NOR2_X1 U15805 ( .A1(n12560), .A2(n9839), .ZN(n12561) );
  OR2_X1 U15806 ( .A1(n12582), .A2(n12561), .ZN(n12578) );
  OAI21_X1 U15807 ( .B1(n12563), .B2(n12564), .A(n12613), .ZN(n12568) );
  INV_X1 U15808 ( .A(n12564), .ZN(n12566) );
  OAI211_X1 U15809 ( .C1(n13334), .C2(n12566), .A(n19838), .B(n12565), .ZN(
        n12567) );
  OAI211_X1 U15810 ( .C1(n12562), .C2(n12569), .A(n12568), .B(n12567), .ZN(
        n12574) );
  NAND2_X1 U15811 ( .A1(n19114), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12581) );
  NAND2_X1 U15812 ( .A1(n12581), .A2(n13334), .ZN(n12570) );
  MUX2_X1 U15813 ( .A(n9839), .B(n12570), .S(n12569), .Z(n12573) );
  AOI21_X1 U15814 ( .B1(n12574), .B2(n12573), .A(n12572), .ZN(n12575) );
  AOI21_X1 U15815 ( .B1(n12576), .B2(n9839), .A(n12575), .ZN(n12577) );
  NOR2_X1 U15816 ( .A1(n12578), .A2(n12577), .ZN(n12579) );
  MUX2_X1 U15817 ( .A(n15664), .B(n12579), .S(P2_STATE2_REG_0__SCAN_IN), .Z(
        n12580) );
  NAND2_X1 U15818 ( .A1(n12582), .A2(n19835), .ZN(n12583) );
  NAND2_X1 U15819 ( .A1(n16257), .A2(n13334), .ZN(n19015) );
  NAND2_X1 U15820 ( .A1(READY21_REG_SCAN_IN), .A2(READY12_REG_SCAN_IN), .ZN(
        n19849) );
  INV_X1 U15821 ( .A(n19849), .ZN(n19843) );
  INV_X1 U15822 ( .A(P2_STATE_REG_1__SCAN_IN), .ZN(n18764) );
  INV_X1 U15823 ( .A(P2_STATE_REG_2__SCAN_IN), .ZN(n19735) );
  NOR2_X1 U15824 ( .A1(n18764), .A2(n19735), .ZN(n19727) );
  NOR2_X1 U15825 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(P2_STATE_REG_2__SCAN_IN), 
        .ZN(n19728) );
  NOR3_X1 U15826 ( .A1(P2_STATE_REG_0__SCAN_IN), .A2(n19727), .A3(n19728), 
        .ZN(n19721) );
  INV_X1 U15827 ( .A(n19721), .ZN(n19837) );
  NOR2_X1 U15828 ( .A1(n19843), .A2(n19837), .ZN(n13611) );
  NAND2_X1 U15829 ( .A1(n19124), .A2(n13611), .ZN(n12611) );
  AOI21_X1 U15830 ( .B1(n12584), .B2(n19838), .A(n12645), .ZN(n12585) );
  NAND2_X1 U15831 ( .A1(n19015), .A2(n12585), .ZN(n12610) );
  MUX2_X1 U15832 ( .A(n12586), .B(n19124), .S(n16281), .Z(n12587) );
  NAND2_X1 U15833 ( .A1(n12587), .A2(n19849), .ZN(n12606) );
  NAND2_X1 U15834 ( .A1(n12589), .A2(n12588), .ZN(n12590) );
  NAND2_X1 U15835 ( .A1(n12590), .A2(n10443), .ZN(n12591) );
  NAND2_X1 U15836 ( .A1(n12591), .A2(n10843), .ZN(n12640) );
  NAND2_X1 U15837 ( .A1(n12592), .A2(n16281), .ZN(n12632) );
  AOI21_X1 U15838 ( .B1(n19114), .B2(n10443), .A(n19124), .ZN(n12593) );
  NAND2_X1 U15839 ( .A1(n12632), .A2(n12593), .ZN(n12594) );
  AND4_X1 U15840 ( .A1(n12596), .A2(n12640), .A3(n12595), .A4(n12594), .ZN(
        n12602) );
  INV_X1 U15841 ( .A(n12597), .ZN(n12600) );
  OAI21_X1 U15842 ( .B1(n12600), .B2(n19124), .A(n12599), .ZN(n12601) );
  AND2_X1 U15843 ( .A1(n12602), .A2(n12601), .ZN(n12634) );
  AND2_X1 U15844 ( .A1(n12603), .A2(n13611), .ZN(n12604) );
  NAND2_X1 U15845 ( .A1(n12586), .A2(n12604), .ZN(n12605) );
  AND2_X1 U15846 ( .A1(n12634), .A2(n12605), .ZN(n13609) );
  OAI21_X1 U15847 ( .B1(n16255), .B2(n12606), .A(n13609), .ZN(n12607) );
  NOR2_X1 U15848 ( .A1(n12608), .A2(n12607), .ZN(n12609) );
  OAI211_X1 U15849 ( .C1(n19015), .C2(n12611), .A(n12610), .B(n12609), .ZN(
        n12612) );
  NAND2_X1 U15850 ( .A1(n12614), .A2(n12613), .ZN(n19825) );
  INV_X1 U15851 ( .A(n14292), .ZN(n12619) );
  INV_X1 U15852 ( .A(n16223), .ZN(n12618) );
  NAND2_X1 U15853 ( .A1(n12619), .A2(n12618), .ZN(n12860) );
  AOI22_X1 U15854 ( .A1(n12622), .A2(P2_EBX_REG_31__SCAN_IN), .B1(
        P2_STATE2_REG_1__SCAN_IN), .B2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), 
        .ZN(n12624) );
  NAND2_X1 U15855 ( .A1(n9899), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n12623) );
  OAI211_X1 U15856 ( .C1(n12625), .C2(n12616), .A(n12624), .B(n12623), .ZN(
        n12626) );
  NAND2_X1 U15857 ( .A1(n12628), .A2(n16281), .ZN(n12630) );
  AND2_X1 U15858 ( .A1(n12630), .A2(n10472), .ZN(n12631) );
  INV_X1 U15859 ( .A(n12632), .ZN(n12633) );
  INV_X1 U15860 ( .A(n13592), .ZN(n16252) );
  MUX2_X1 U15861 ( .A(n12562), .B(n10293), .S(n12635), .Z(n12637) );
  NAND2_X1 U15862 ( .A1(n12637), .A2(n12636), .ZN(n12638) );
  NAND2_X1 U15863 ( .A1(n12638), .A2(n10426), .ZN(n12649) );
  NAND2_X1 U15864 ( .A1(n12639), .A2(n13334), .ZN(n15518) );
  NAND2_X1 U15865 ( .A1(n15518), .A2(n12640), .ZN(n12642) );
  NAND2_X1 U15866 ( .A1(n12642), .A2(n12641), .ZN(n12648) );
  OAI22_X1 U15867 ( .A1(n12636), .A2(n12645), .B1(n12644), .B2(n19838), .ZN(
        n12646) );
  NOR2_X1 U15868 ( .A1(n12643), .A2(n12646), .ZN(n12647) );
  NAND3_X1 U15869 ( .A1(n12649), .A2(n12648), .A3(n12647), .ZN(n15541) );
  NOR2_X1 U15870 ( .A1(n15541), .A2(n13181), .ZN(n12650) );
  NAND3_X1 U15871 ( .A1(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12848) );
  AND2_X1 U15872 ( .A1(n12663), .A2(n18934), .ZN(n15511) );
  INV_X1 U15873 ( .A(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n20914) );
  INV_X1 U15874 ( .A(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15530) );
  NOR2_X1 U15875 ( .A1(n20914), .A2(n15530), .ZN(n13408) );
  NOR2_X1 U15876 ( .A1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n13408), .ZN(
        n12849) );
  NOR2_X1 U15877 ( .A1(n13925), .A2(n13924), .ZN(n13991) );
  NAND3_X1 U15878 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n13991), .ZN(n14087) );
  NAND2_X1 U15879 ( .A1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n16202) );
  OR3_X1 U15880 ( .A1(n12849), .A2(n14087), .A3(n16202), .ZN(n12653) );
  AOI21_X1 U15881 ( .B1(P2_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n13408), .A(
        n15400), .ZN(n12651) );
  NOR2_X1 U15882 ( .A1(n15511), .A2(n12651), .ZN(n13873) );
  NAND2_X1 U15883 ( .A1(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A2(n13873), .ZN(
        n12652) );
  AOI21_X1 U15884 ( .B1(n15514), .B2(n12653), .A(n12652), .ZN(n15495) );
  AND2_X1 U15885 ( .A1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12852) );
  NAND2_X1 U15886 ( .A1(n15495), .A2(n12852), .ZN(n15396) );
  INV_X1 U15887 ( .A(n15396), .ZN(n12654) );
  AND2_X1 U15888 ( .A1(n12853), .A2(n12654), .ZN(n15280) );
  NAND2_X1 U15889 ( .A1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12655) );
  NOR2_X1 U15890 ( .A1(n15301), .A2(n12655), .ZN(n12855) );
  NAND2_X1 U15891 ( .A1(n15280), .A2(n12855), .ZN(n12656) );
  AND2_X1 U15892 ( .A1(n15397), .A2(n12656), .ZN(n15273) );
  AOI211_X1 U15893 ( .C1(n15514), .C2(n12848), .A(n12548), .B(n15273), .ZN(
        n14269) );
  INV_X1 U15894 ( .A(n15397), .ZN(n15471) );
  NOR3_X1 U15895 ( .A1(n14269), .A2(n15471), .A3(n12616), .ZN(n12858) );
  AND2_X1 U15896 ( .A1(n12659), .A2(n12658), .ZN(n15520) );
  AND2_X1 U15897 ( .A1(n12660), .A2(n12599), .ZN(n16253) );
  OR2_X1 U15898 ( .A1(n16253), .A2(n16281), .ZN(n12661) );
  AND2_X1 U15899 ( .A1(n13591), .A2(n12661), .ZN(n12662) );
  INV_X1 U15900 ( .A(n12819), .ZN(n12736) );
  NOR2_X1 U15901 ( .A1(n13334), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12665) );
  NAND2_X1 U15902 ( .A1(n13388), .A2(n12665), .ZN(n12685) );
  INV_X1 U15903 ( .A(P2_REIP_REG_0__SCAN_IN), .ZN(n18955) );
  AOI21_X1 U15904 ( .B1(n13334), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12667) );
  NAND2_X1 U15905 ( .A1(n10238), .A2(P2_EAX_REG_0__SCAN_IN), .ZN(n12666) );
  OAI211_X1 U15906 ( .C1(n12685), .C2(n18955), .A(n12667), .B(n12666), .ZN(
        n13345) );
  MUX2_X1 U15907 ( .A(n10443), .B(n19823), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12669) );
  NAND2_X1 U15908 ( .A1(n10420), .A2(n12684), .ZN(n12681) );
  OAI21_X1 U15909 ( .B1(n12819), .B2(n12671), .A(n12670), .ZN(n13344) );
  NOR2_X1 U15910 ( .A1(n10443), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n12672) );
  AOI22_X1 U15911 ( .A1(n12672), .A2(P2_EAX_REG_1__SCAN_IN), .B1(n12684), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n12673) );
  OAI21_X1 U15912 ( .B1(n12685), .B2(n10425), .A(n12673), .ZN(n12678) );
  INV_X1 U15913 ( .A(n12678), .ZN(n12674) );
  NAND2_X1 U15914 ( .A1(n10442), .A2(n10443), .ZN(n12675) );
  MUX2_X1 U15915 ( .A(n12675), .B(n19814), .S(P2_STATE2_REG_3__SCAN_IN), .Z(
        n12676) );
  OAI21_X1 U15916 ( .B1(n12677), .B2(n12819), .A(n12676), .ZN(n13718) );
  NOR2_X1 U15917 ( .A1(n13343), .A2(n12678), .ZN(n12679) );
  NAND2_X1 U15918 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n12682) );
  OAI211_X1 U15919 ( .C1(n12819), .C2(n12683), .A(n12682), .B(n12681), .ZN(
        n12686) );
  XNOR2_X1 U15920 ( .A(n12687), .B(n12686), .ZN(n13398) );
  INV_X1 U15921 ( .A(P2_EAX_REG_2__SCAN_IN), .ZN(n20879) );
  OAI222_X1 U15922 ( .A1(n12710), .A2(n9963), .B1(n12709), .B2(n20879), .C1(
        n12845), .C2(n10480), .ZN(n13397) );
  NOR2_X1 U15923 ( .A1(n13398), .A2(n13397), .ZN(n13396) );
  NOR2_X1 U15924 ( .A1(n12687), .A2(n12686), .ZN(n12688) );
  AOI22_X1 U15925 ( .A1(n12841), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .B1(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(P2_STATE2_REG_3__SCAN_IN), 
        .ZN(n12689) );
  OAI21_X1 U15926 ( .B1(n12845), .B2(n12690), .A(n12689), .ZN(n12694) );
  INV_X2 U15927 ( .A(n12709), .ZN(n12846) );
  NAND2_X1 U15928 ( .A1(n12846), .A2(P2_EAX_REG_3__SCAN_IN), .ZN(n12691) );
  OAI21_X1 U15929 ( .B1(n12819), .B2(n12692), .A(n12691), .ZN(n12693) );
  AOI22_X1 U15930 ( .A1(n12846), .A2(P2_EAX_REG_4__SCAN_IN), .B1(n12841), .B2(
        P2_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n12699) );
  INV_X1 U15931 ( .A(n12696), .ZN(n12697) );
  OR2_X1 U15932 ( .A1(n12819), .A2(n12697), .ZN(n12698) );
  OAI211_X1 U15933 ( .C1(n12845), .C2(n12700), .A(n12699), .B(n12698), .ZN(
        n13835) );
  INV_X1 U15934 ( .A(n13835), .ZN(n12701) );
  AOI22_X1 U15935 ( .A1(n12695), .A2(P2_REIP_REG_5__SCAN_IN), .B1(n12736), 
        .B2(n12702), .ZN(n12704) );
  AOI22_X1 U15936 ( .A1(n12846), .A2(P2_EAX_REG_5__SCAN_IN), .B1(n12841), .B2(
        P2_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n12703) );
  NAND2_X1 U15937 ( .A1(n12704), .A2(n12703), .ZN(n13930) );
  INV_X1 U15938 ( .A(n13929), .ZN(n12705) );
  AOI21_X1 U15939 ( .B1(n12736), .B2(n12706), .A(n12705), .ZN(n13395) );
  AOI22_X1 U15940 ( .A1(n12846), .A2(P2_EAX_REG_6__SCAN_IN), .B1(n12841), .B2(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n12707) );
  OAI21_X1 U15941 ( .B1(n12845), .B2(n10912), .A(n12707), .ZN(n13394) );
  INV_X1 U15942 ( .A(n13394), .ZN(n12708) );
  INV_X1 U15943 ( .A(P2_EAX_REG_7__SCAN_IN), .ZN(n19065) );
  OAI222_X1 U15944 ( .A1(n12710), .A2(n10882), .B1(n12709), .B2(n19065), .C1(
        n12845), .C2(n10916), .ZN(n13499) );
  AOI22_X1 U15945 ( .A1(n12846), .A2(P2_EAX_REG_8__SCAN_IN), .B1(n12841), .B2(
        P2_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n12723) );
  AOI22_X1 U15946 ( .A1(n10554), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n10566), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12714) );
  AOI22_X1 U15947 ( .A1(n10671), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10567), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12713) );
  AOI22_X1 U15948 ( .A1(n10690), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12712) );
  AOI22_X1 U15949 ( .A1(n13593), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12711) );
  NAND4_X1 U15950 ( .A1(n12714), .A2(n12713), .A3(n12712), .A4(n12711), .ZN(
        n12720) );
  AOI22_X1 U15951 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .B1(
        n12954), .B2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n12718) );
  AOI22_X1 U15952 ( .A1(n10695), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12975), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12717) );
  AOI22_X1 U15953 ( .A1(n10559), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12716) );
  AOI22_X1 U15954 ( .A1(n12952), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12715) );
  NAND4_X1 U15955 ( .A1(n12718), .A2(n12717), .A3(n12716), .A4(n12715), .ZN(
        n12719) );
  INV_X1 U15956 ( .A(n13575), .ZN(n12721) );
  OR2_X1 U15957 ( .A1(n12819), .A2(n12721), .ZN(n12722) );
  OAI211_X1 U15958 ( .C1(n12845), .C2(n14050), .A(n12723), .B(n12722), .ZN(
        n12724) );
  INV_X1 U15959 ( .A(n12724), .ZN(n14049) );
  AOI22_X1 U15960 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n10676), .B1(
        n10554), .B2(P2_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n12729) );
  AOI22_X1 U15961 ( .A1(n10671), .A2(P2_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12728) );
  AOI22_X1 U15962 ( .A1(P2_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n10567), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n12727) );
  AOI22_X1 U15963 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n13593), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n12726) );
  NAND4_X1 U15964 ( .A1(n12729), .A2(n12728), .A3(n12727), .A4(n12726), .ZN(
        n12735) );
  AOI22_X1 U15965 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n10566), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12733) );
  AOI22_X1 U15966 ( .A1(n10559), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n12975), .ZN(n12732) );
  AOI22_X1 U15967 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10695), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12731) );
  AOI22_X1 U15968 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n12730) );
  NAND4_X1 U15969 ( .A1(n12733), .A2(n12732), .A3(n12731), .A4(n12730), .ZN(
        n12734) );
  AOI22_X1 U15970 ( .A1(P2_REIP_REG_9__SCAN_IN), .A2(n12695), .B1(n12736), 
        .B2(n12890), .ZN(n12738) );
  AOI22_X1 U15971 ( .A1(n12846), .A2(P2_EAX_REG_9__SCAN_IN), .B1(n12841), .B2(
        P2_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n12737) );
  NAND2_X1 U15972 ( .A1(n12738), .A2(n12737), .ZN(n14888) );
  AOI22_X1 U15973 ( .A1(n12846), .A2(P2_EAX_REG_10__SCAN_IN), .B1(n12841), 
        .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n12750) );
  AOI22_X1 U15974 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n10676), .B1(
        n10554), .B2(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n12742) );
  AOI22_X1 U15975 ( .A1(n10671), .A2(P2_INSTQUEUE_REG_3__2__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12741) );
  AOI22_X1 U15976 ( .A1(P2_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n10567), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n12740) );
  AOI22_X1 U15977 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n12725), .B1(
        n13593), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12739) );
  NAND4_X1 U15978 ( .A1(n12742), .A2(n12741), .A3(n12740), .A4(n12739), .ZN(
        n12748) );
  AOI22_X1 U15979 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n10566), .B1(
        n12954), .B2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n12746) );
  AOI22_X1 U15980 ( .A1(n10559), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__2__SCAN_IN), .B2(n12975), .ZN(n12745) );
  AOI22_X1 U15981 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n10695), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n12744) );
  AOI22_X1 U15982 ( .A1(n12952), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12743) );
  NAND4_X1 U15983 ( .A1(n12746), .A2(n12745), .A3(n12744), .A4(n12743), .ZN(
        n12747) );
  NOR2_X1 U15984 ( .A1(n12748), .A2(n12747), .ZN(n13745) );
  OR2_X1 U15985 ( .A1(n12819), .A2(n13745), .ZN(n12749) );
  OAI211_X1 U15986 ( .C1(n12845), .C2(n12751), .A(n12750), .B(n12749), .ZN(
        n12752) );
  INV_X1 U15987 ( .A(n12752), .ZN(n15484) );
  AOI22_X1 U15988 ( .A1(n12846), .A2(P2_EAX_REG_11__SCAN_IN), .B1(n12841), 
        .B2(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n12764) );
  AOI22_X1 U15989 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n10676), .B1(
        n10554), .B2(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n12756) );
  AOI22_X1 U15990 ( .A1(n10671), .A2(P2_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12755) );
  AOI22_X1 U15991 ( .A1(P2_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n10567), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n12754) );
  AOI22_X1 U15992 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n13593), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n12753) );
  NAND4_X1 U15993 ( .A1(n12756), .A2(n12755), .A3(n12754), .A4(n12753), .ZN(
        n12762) );
  AOI22_X1 U15994 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n10566), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12760) );
  AOI22_X1 U15995 ( .A1(n10559), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__3__SCAN_IN), .B2(n12975), .ZN(n12759) );
  AOI22_X1 U15996 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n10695), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12758) );
  AOI22_X1 U15997 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n12757) );
  NAND4_X1 U15998 ( .A1(n12760), .A2(n12759), .A3(n12758), .A4(n12757), .ZN(
        n12761) );
  OR2_X1 U15999 ( .A1(n12819), .A2(n12892), .ZN(n12763) );
  OAI211_X1 U16000 ( .C1(n12845), .C2(n12765), .A(n12764), .B(n12763), .ZN(
        n13740) );
  NAND2_X1 U16001 ( .A1(n13739), .A2(n13740), .ZN(n13738) );
  AOI22_X1 U16002 ( .A1(n12846), .A2(P2_EAX_REG_12__SCAN_IN), .B1(n12841), 
        .B2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n12778) );
  AOI22_X1 U16003 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n10676), .B1(
        n10554), .B2(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n12769) );
  AOI22_X1 U16004 ( .A1(n10671), .A2(P2_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n10567), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12768) );
  AOI22_X1 U16005 ( .A1(P2_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n10690), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12767) );
  AOI22_X1 U16006 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n13593), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n12766) );
  NAND4_X1 U16007 ( .A1(n12769), .A2(n12768), .A3(n12767), .A4(n12766), .ZN(
        n12775) );
  AOI22_X1 U16008 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n10566), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12773) );
  AOI22_X1 U16009 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__4__SCAN_IN), .B2(n12975), .ZN(n12772) );
  AOI22_X1 U16010 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n10559), .B1(
        n10695), .B2(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n12771) );
  AOI22_X1 U16011 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12770) );
  NAND4_X1 U16012 ( .A1(n12773), .A2(n12772), .A3(n12771), .A4(n12770), .ZN(
        n12774) );
  INV_X1 U16013 ( .A(n13811), .ZN(n12776) );
  OR2_X1 U16014 ( .A1(n12819), .A2(n12776), .ZN(n12777) );
  OAI211_X1 U16015 ( .C1(n12845), .C2(n12779), .A(n12778), .B(n12777), .ZN(
        n13789) );
  INV_X1 U16016 ( .A(n13789), .ZN(n12780) );
  AOI22_X1 U16017 ( .A1(n12846), .A2(P2_EAX_REG_13__SCAN_IN), .B1(n12841), 
        .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n12792) );
  AOI22_X1 U16018 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n10554), .B2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n12784) );
  AOI22_X1 U16019 ( .A1(n10671), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12783) );
  AOI22_X1 U16020 ( .A1(n10690), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n10567), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12782) );
  AOI22_X1 U16021 ( .A1(n13593), .A2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n12781) );
  NAND4_X1 U16022 ( .A1(n12784), .A2(n12783), .A3(n12782), .A4(n12781), .ZN(
        n12790) );
  AOI22_X1 U16023 ( .A1(n10566), .A2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12788) );
  AOI22_X1 U16024 ( .A1(n10559), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n12975), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12787) );
  AOI22_X1 U16025 ( .A1(n10695), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12786) );
  AOI22_X1 U16026 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n12785) );
  NAND4_X1 U16027 ( .A1(n12788), .A2(n12787), .A3(n12786), .A4(n12785), .ZN(
        n12789) );
  OR2_X1 U16028 ( .A1(n12790), .A2(n12789), .ZN(n13846) );
  INV_X1 U16029 ( .A(n13846), .ZN(n13844) );
  OR2_X1 U16030 ( .A1(n12819), .A2(n13844), .ZN(n12791) );
  OAI211_X1 U16031 ( .C1(n12845), .C2(n12793), .A(n12792), .B(n12791), .ZN(
        n13802) );
  AOI22_X1 U16032 ( .A1(n12846), .A2(P2_EAX_REG_14__SCAN_IN), .B1(n12841), 
        .B2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n12805) );
  AOI22_X1 U16033 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n10676), .B1(
        n10554), .B2(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n12797) );
  AOI22_X1 U16034 ( .A1(n10671), .A2(P2_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n10567), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12796) );
  AOI22_X1 U16035 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n10690), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12795) );
  AOI22_X1 U16036 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n13593), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n12794) );
  NAND4_X1 U16037 ( .A1(n12797), .A2(n12796), .A3(n12795), .A4(n12794), .ZN(
        n12803) );
  AOI22_X1 U16038 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n10566), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12801) );
  AOI22_X1 U16039 ( .A1(n12953), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__6__SCAN_IN), .B2(n12975), .ZN(n12800) );
  AOI22_X1 U16040 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n10559), .B1(
        n10695), .B2(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n12799) );
  AOI22_X1 U16041 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12798) );
  NAND4_X1 U16042 ( .A1(n12801), .A2(n12800), .A3(n12799), .A4(n12798), .ZN(
        n12802) );
  OR2_X1 U16043 ( .A1(n12803), .A2(n12802), .ZN(n13891) );
  INV_X1 U16044 ( .A(n13891), .ZN(n13890) );
  OR2_X1 U16045 ( .A1(n12819), .A2(n13890), .ZN(n12804) );
  OAI211_X1 U16046 ( .C1(n12845), .C2(n14023), .A(n12805), .B(n12804), .ZN(
        n12806) );
  INV_X1 U16047 ( .A(n12806), .ZN(n14020) );
  AOI22_X1 U16048 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n10676), .B1(
        n10554), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n12810) );
  AOI22_X1 U16049 ( .A1(n10671), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12809) );
  AOI22_X1 U16050 ( .A1(P2_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n10567), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n12808) );
  AOI22_X1 U16051 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n13593), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n12807) );
  NAND4_X1 U16052 ( .A1(n12810), .A2(n12809), .A3(n12808), .A4(n12807), .ZN(
        n12816) );
  AOI22_X1 U16053 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n10566), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12814) );
  AOI22_X1 U16054 ( .A1(n10559), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_1__7__SCAN_IN), .B2(n12975), .ZN(n12813) );
  AOI22_X1 U16055 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n10695), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12812) );
  AOI22_X1 U16056 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n12811) );
  NAND4_X1 U16057 ( .A1(n12814), .A2(n12813), .A3(n12812), .A4(n12811), .ZN(
        n12815) );
  OR2_X1 U16058 ( .A1(n12816), .A2(n12815), .ZN(n13911) );
  INV_X1 U16059 ( .A(n13911), .ZN(n12923) );
  NAND2_X1 U16060 ( .A1(n12695), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n12818) );
  AOI22_X1 U16061 ( .A1(n12846), .A2(P2_EAX_REG_15__SCAN_IN), .B1(n12841), 
        .B2(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n12817) );
  OAI211_X1 U16062 ( .C1(n12923), .C2(n12819), .A(n12818), .B(n12817), .ZN(
        n13851) );
  AOI22_X1 U16063 ( .A1(n12846), .A2(P2_EAX_REG_16__SCAN_IN), .B1(n12684), 
        .B2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n12820) );
  OAI21_X1 U16064 ( .B1(n12845), .B2(n15415), .A(n12820), .ZN(n15413) );
  AOI22_X1 U16065 ( .A1(n12846), .A2(P2_EAX_REG_17__SCAN_IN), .B1(n12841), 
        .B2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n12821) );
  OAI21_X1 U16066 ( .B1(n12845), .B2(n19750), .A(n12821), .ZN(n12822) );
  INV_X1 U16067 ( .A(n12822), .ZN(n14067) );
  AOI22_X1 U16068 ( .A1(n12846), .A2(P2_EAX_REG_18__SCAN_IN), .B1(n12841), 
        .B2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n12824) );
  OAI21_X1 U16069 ( .B1(n12845), .B2(n19752), .A(n12824), .ZN(n12825) );
  INV_X1 U16070 ( .A(n12825), .ZN(n15380) );
  AOI22_X1 U16071 ( .A1(n12846), .A2(P2_EAX_REG_19__SCAN_IN), .B1(n12841), 
        .B2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n12826) );
  OAI21_X1 U16072 ( .B1(n12845), .B2(n19754), .A(n12826), .ZN(n15082) );
  AOI22_X1 U16073 ( .A1(n12846), .A2(P2_EAX_REG_20__SCAN_IN), .B1(n12841), 
        .B2(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n12827) );
  OAI21_X1 U16074 ( .B1(n12845), .B2(n19756), .A(n12827), .ZN(n13243) );
  AOI22_X1 U16075 ( .A1(n12846), .A2(P2_EAX_REG_21__SCAN_IN), .B1(n12841), 
        .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n12828) );
  OAI21_X1 U16076 ( .B1(n12845), .B2(n19758), .A(n12828), .ZN(n14872) );
  AOI22_X1 U16077 ( .A1(n12846), .A2(P2_EAX_REG_22__SCAN_IN), .B1(n12841), 
        .B2(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n12829) );
  OAI21_X1 U16078 ( .B1(n12845), .B2(n12830), .A(n12829), .ZN(n15330) );
  AOI22_X1 U16079 ( .A1(n12846), .A2(P2_EAX_REG_23__SCAN_IN), .B1(n12684), 
        .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n12831) );
  OAI21_X1 U16080 ( .B1(n12845), .B2(n10960), .A(n12831), .ZN(n15066) );
  NAND2_X1 U16081 ( .A1(n12695), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n12833) );
  AOI22_X1 U16082 ( .A1(n12846), .A2(P2_EAX_REG_24__SCAN_IN), .B1(n12841), 
        .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n12832) );
  AND2_X1 U16083 ( .A1(n12833), .A2(n12832), .ZN(n15059) );
  NAND2_X1 U16084 ( .A1(n12695), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n12835) );
  AOI22_X1 U16085 ( .A1(n12846), .A2(P2_EAX_REG_25__SCAN_IN), .B1(n12684), 
        .B2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n12834) );
  AOI22_X1 U16086 ( .A1(n12846), .A2(P2_EAX_REG_26__SCAN_IN), .B1(n12841), 
        .B2(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n12836) );
  OAI21_X1 U16087 ( .B1(n12845), .B2(n21017), .A(n12836), .ZN(n15043) );
  NAND2_X1 U16088 ( .A1(n15044), .A2(n15043), .ZN(n15033) );
  NAND2_X1 U16089 ( .A1(n12695), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n12838) );
  AOI22_X1 U16090 ( .A1(n12846), .A2(P2_EAX_REG_27__SCAN_IN), .B1(n12841), 
        .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n12837) );
  AND2_X1 U16091 ( .A1(n12838), .A2(n12837), .ZN(n15034) );
  NAND2_X1 U16092 ( .A1(n12695), .A2(P2_REIP_REG_28__SCAN_IN), .ZN(n12840) );
  AOI22_X1 U16093 ( .A1(n12846), .A2(P2_EAX_REG_28__SCAN_IN), .B1(n12841), 
        .B2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n12839) );
  AND2_X1 U16094 ( .A1(n12840), .A2(n12839), .ZN(n15024) );
  AOI22_X1 U16095 ( .A1(n12846), .A2(P2_EAX_REG_29__SCAN_IN), .B1(n12841), 
        .B2(P2_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n12842) );
  OAI21_X1 U16096 ( .B1(n12845), .B2(n19770), .A(n12842), .ZN(n14234) );
  AOI22_X1 U16097 ( .A1(n12846), .A2(P2_EAX_REG_30__SCAN_IN), .B1(n12841), 
        .B2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n12843) );
  OAI21_X1 U16098 ( .B1(n12845), .B2(n12844), .A(n12843), .ZN(n14262) );
  NAND2_X1 U16099 ( .A1(n14261), .A2(n14262), .ZN(n14266) );
  AOI222_X1 U16100 ( .A1(n12695), .A2(P2_REIP_REG_31__SCAN_IN), .B1(n12846), 
        .B2(P2_EAX_REG_31__SCAN_IN), .C1(n12841), .C2(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n12847) );
  NAND2_X1 U16101 ( .A1(n19085), .A2(P2_REIP_REG_31__SCAN_IN), .ZN(n14288) );
  INV_X1 U16102 ( .A(n12848), .ZN(n14268) );
  INV_X1 U16103 ( .A(n13875), .ZN(n15395) );
  INV_X1 U16104 ( .A(n13408), .ZN(n15513) );
  NOR2_X1 U16105 ( .A1(n9963), .A2(n15513), .ZN(n12850) );
  INV_X1 U16106 ( .A(n12849), .ZN(n13874) );
  OAI211_X1 U16107 ( .C1(n15395), .C2(n12850), .A(n13874), .B(n15514), .ZN(
        n16230) );
  NOR2_X1 U16108 ( .A1(n16230), .A2(n14087), .ZN(n16203) );
  INV_X1 U16109 ( .A(n16202), .ZN(n12851) );
  NAND2_X1 U16110 ( .A1(n16203), .A2(n12851), .ZN(n15496) );
  NOR2_X1 U16111 ( .A1(n15497), .A2(n15496), .ZN(n15488) );
  INV_X1 U16112 ( .A(n12853), .ZN(n12854) );
  NOR2_X1 U16113 ( .A1(n15444), .A2(n12854), .ZN(n15302) );
  NAND2_X1 U16114 ( .A1(n15302), .A2(n12855), .ZN(n15258) );
  INV_X1 U16115 ( .A(n15258), .ZN(n14267) );
  NAND4_X1 U16116 ( .A1(n14268), .A2(P2_INSTADDRPOINTER_REG_30__SCAN_IN), .A3(
        n12616), .A4(n14267), .ZN(n12856) );
  OAI211_X1 U16117 ( .C1(n16222), .C2(n16012), .A(n14288), .B(n12856), .ZN(
        n12857) );
  AND2_X1 U16118 ( .A1(n12860), .A2(n12859), .ZN(n12861) );
  OAI21_X1 U16119 ( .B1(n14295), .B2(n16217), .A(n12861), .ZN(P2_U3015) );
  NAND2_X1 U16120 ( .A1(n9817), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n12862) );
  AND2_X1 U16121 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n19470) );
  NOR2_X1 U16122 ( .A1(n16248), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19319) );
  INV_X1 U16123 ( .A(n19382), .ZN(n19379) );
  NOR2_X1 U16124 ( .A1(n16248), .A2(n19814), .ZN(n19610) );
  NAND2_X1 U16125 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19610), .ZN(
        n13937) );
  NAND2_X1 U16126 ( .A1(n13937), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n12863) );
  AOI21_X1 U16127 ( .B1(n19379), .B2(n12863), .A(n19790), .ZN(n19512) );
  AOI21_X1 U16128 ( .B1(n12878), .B2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A(
        n19512), .ZN(n12864) );
  NOR2_X1 U16129 ( .A1(n13584), .A2(n19133), .ZN(n13505) );
  AND3_X1 U16130 ( .A1(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A2(
        P2_INSTQUEUE_REG_0__5__SCAN_IN), .A3(P2_INSTQUEUE_REG_0__4__SCAN_IN), 
        .ZN(n12866) );
  NAND2_X1 U16131 ( .A1(n12867), .A2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(
        n12887) );
  NAND2_X1 U16132 ( .A1(n12868), .A2(n12881), .ZN(n12871) );
  OAI21_X1 U16133 ( .B1(n19470), .B2(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A(
        n13937), .ZN(n19249) );
  NOR2_X1 U16134 ( .A1(n19249), .A2(n19790), .ZN(n12869) );
  AOI21_X1 U16135 ( .B1(n12878), .B2(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(
        n12869), .ZN(n12870) );
  NAND2_X1 U16136 ( .A1(n12871), .A2(n12870), .ZN(n12874) );
  INV_X1 U16137 ( .A(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12872) );
  NOR2_X1 U16138 ( .A1(n13584), .A2(n12872), .ZN(n12873) );
  OR2_X1 U16139 ( .A1(n12874), .A2(n12873), .ZN(n12875) );
  NAND2_X1 U16140 ( .A1(n12874), .A2(n12873), .ZN(n12885) );
  AOI22_X1 U16141 ( .A1(n12878), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B1(
        n19612), .B2(n19823), .ZN(n12876) );
  INV_X1 U16142 ( .A(n13584), .ZN(n13109) );
  NAND2_X1 U16143 ( .A1(n13109), .A2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(
        n12882) );
  NAND2_X1 U16144 ( .A1(n12878), .A2(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(
        n12879) );
  NAND2_X1 U16145 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19814), .ZN(
        n19406) );
  NAND2_X1 U16146 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n19823), .ZN(
        n19437) );
  NAND2_X1 U16147 ( .A1(n19406), .A2(n19437), .ZN(n19320) );
  NAND2_X1 U16148 ( .A1(n19612), .A2(n19320), .ZN(n19440) );
  NAND2_X1 U16149 ( .A1(n12879), .A2(n19440), .ZN(n12880) );
  INV_X1 U16150 ( .A(n12882), .ZN(n12883) );
  NOR2_X1 U16151 ( .A1(n15523), .A2(n12883), .ZN(n12884) );
  INV_X1 U16152 ( .A(n12885), .ZN(n12886) );
  NAND2_X1 U16153 ( .A1(n12887), .A2(n13508), .ZN(n12888) );
  NAND2_X1 U16154 ( .A1(n13576), .A2(n13575), .ZN(n13574) );
  AOI22_X1 U16155 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n10676), .B1(
        n10554), .B2(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n12896) );
  AOI22_X1 U16156 ( .A1(n10671), .A2(P2_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n12895) );
  AOI22_X1 U16157 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n10690), .B1(
        n10567), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n12894) );
  AOI22_X1 U16158 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n13593), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n12893) );
  NAND4_X1 U16159 ( .A1(n12896), .A2(n12895), .A3(n12894), .A4(n12893), .ZN(
        n12902) );
  AOI22_X1 U16160 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n10566), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n12900) );
  AOI22_X1 U16161 ( .A1(n10559), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__2__SCAN_IN), .B2(n12975), .ZN(n12899) );
  AOI22_X1 U16162 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n10695), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n12898) );
  AOI22_X1 U16163 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n12897) );
  NAND4_X1 U16164 ( .A1(n12900), .A2(n12899), .A3(n12898), .A4(n12897), .ZN(
        n12901) );
  OR2_X1 U16165 ( .A1(n12902), .A2(n12901), .ZN(n14111) );
  AOI22_X1 U16166 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n10676), .B1(
        n10554), .B2(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n12906) );
  AOI22_X1 U16167 ( .A1(n10671), .A2(P2_INSTQUEUE_REG_4__1__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n12905) );
  AOI22_X1 U16168 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n10690), .B1(
        n10567), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n12904) );
  AOI22_X1 U16169 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n13593), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n12903) );
  NAND4_X1 U16170 ( .A1(n12906), .A2(n12905), .A3(n12904), .A4(n12903), .ZN(
        n12912) );
  AOI22_X1 U16171 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n10566), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n12910) );
  AOI22_X1 U16172 ( .A1(n10559), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n12975), .ZN(n12909) );
  AOI22_X1 U16173 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n10695), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n12908) );
  AOI22_X1 U16174 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_7__1__SCAN_IN), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n12907) );
  NAND4_X1 U16175 ( .A1(n12910), .A2(n12909), .A3(n12908), .A4(n12907), .ZN(
        n12911) );
  OR2_X1 U16176 ( .A1(n12912), .A2(n12911), .ZN(n13998) );
  AOI22_X1 U16177 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10554), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12916) );
  AOI22_X1 U16178 ( .A1(n10671), .A2(P2_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n12915) );
  AOI22_X1 U16179 ( .A1(n10690), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .B1(
        n10567), .B2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n12914) );
  AOI22_X1 U16180 ( .A1(n13593), .A2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n12913) );
  NAND4_X1 U16181 ( .A1(n12916), .A2(n12915), .A3(n12914), .A4(n12913), .ZN(
        n12922) );
  AOI22_X1 U16182 ( .A1(n10566), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n12920) );
  AOI22_X1 U16183 ( .A1(n10559), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n12975), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12919) );
  AOI22_X1 U16184 ( .A1(n10695), .A2(P2_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n12918) );
  AOI22_X1 U16185 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12917) );
  NAND4_X1 U16186 ( .A1(n12920), .A2(n12919), .A3(n12918), .A4(n12917), .ZN(
        n12921) );
  OR2_X1 U16187 ( .A1(n12922), .A2(n12921), .ZN(n13962) );
  INV_X1 U16188 ( .A(n13962), .ZN(n12924) );
  OR2_X1 U16189 ( .A1(n12923), .A2(n13890), .ZN(n13908) );
  OR2_X1 U16190 ( .A1(n12924), .A2(n13908), .ZN(n12925) );
  NOR2_X1 U16191 ( .A1(n12925), .A2(n13844), .ZN(n13960) );
  AND2_X1 U16192 ( .A1(n13998), .A2(n13960), .ZN(n12926) );
  AOI22_X1 U16193 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n10676), .B1(
        n10554), .B2(P2_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n12931) );
  AOI22_X1 U16194 ( .A1(n10671), .A2(P2_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n12930) );
  AOI22_X1 U16195 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n10690), .B1(
        n10567), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n12929) );
  AOI22_X1 U16196 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n13593), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n12928) );
  NAND4_X1 U16197 ( .A1(n12931), .A2(n12930), .A3(n12929), .A4(n12928), .ZN(
        n12937) );
  AOI22_X1 U16198 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n10566), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n12935) );
  AOI22_X1 U16199 ( .A1(n10559), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__3__SCAN_IN), .B2(n12975), .ZN(n12934) );
  AOI22_X1 U16200 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n10695), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n12933) );
  AOI22_X1 U16201 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n12932) );
  NAND4_X1 U16202 ( .A1(n12935), .A2(n12934), .A3(n12933), .A4(n12932), .ZN(
        n12936) );
  NOR2_X1 U16203 ( .A1(n12937), .A2(n12936), .ZN(n14102) );
  AOI22_X1 U16204 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n10676), .B1(
        n10554), .B2(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n12941) );
  AOI22_X1 U16205 ( .A1(n10671), .A2(P2_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n12940) );
  AOI22_X1 U16206 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n10567), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n12939) );
  AOI22_X1 U16207 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n13593), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n12938) );
  NAND4_X1 U16208 ( .A1(n12941), .A2(n12940), .A3(n12939), .A4(n12938), .ZN(
        n12947) );
  AOI22_X1 U16209 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n10566), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n12945) );
  AOI22_X1 U16210 ( .A1(n10559), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__4__SCAN_IN), .B2(n12975), .ZN(n12944) );
  AOI22_X1 U16211 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n10695), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n12943) );
  AOI22_X1 U16212 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_7__4__SCAN_IN), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n12942) );
  NAND4_X1 U16213 ( .A1(n12945), .A2(n12944), .A3(n12943), .A4(n12942), .ZN(
        n12946) );
  OR2_X1 U16214 ( .A1(n12947), .A2(n12946), .ZN(n14118) );
  AOI22_X1 U16215 ( .A1(n10676), .A2(P2_INSTQUEUE_REG_3__5__SCAN_IN), .B1(
        n10554), .B2(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n12951) );
  AOI22_X1 U16216 ( .A1(n10671), .A2(P2_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n12950) );
  AOI22_X1 U16217 ( .A1(n10690), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(
        n10567), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n12949) );
  AOI22_X1 U16218 ( .A1(n13593), .A2(P2_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n12948) );
  NAND4_X1 U16219 ( .A1(n12951), .A2(n12950), .A3(n12949), .A4(n12948), .ZN(
        n12960) );
  AOI22_X1 U16220 ( .A1(n10566), .A2(P2_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n12958) );
  AOI22_X1 U16221 ( .A1(n10559), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(
        n12975), .B2(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n12957) );
  AOI22_X1 U16222 ( .A1(n10695), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n12956) );
  AOI22_X1 U16223 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n12955) );
  NAND4_X1 U16224 ( .A1(n12958), .A2(n12957), .A3(n12956), .A4(n12955), .ZN(
        n12959) );
  OR2_X1 U16225 ( .A1(n12960), .A2(n12959), .ZN(n15005) );
  AOI22_X1 U16226 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n10676), .B1(
        n10554), .B2(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n12964) );
  AOI22_X1 U16227 ( .A1(n10671), .A2(P2_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n12963) );
  AOI22_X1 U16228 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n10567), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n12962) );
  AOI22_X1 U16229 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n13593), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n12961) );
  NAND4_X1 U16230 ( .A1(n12964), .A2(n12963), .A3(n12962), .A4(n12961), .ZN(
        n12970) );
  AOI22_X1 U16231 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n10566), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n12968) );
  AOI22_X1 U16232 ( .A1(n10559), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__6__SCAN_IN), .B2(n12975), .ZN(n12967) );
  AOI22_X1 U16233 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n10695), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n12966) );
  AOI22_X1 U16234 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n12965) );
  NAND4_X1 U16235 ( .A1(n12968), .A2(n12967), .A3(n12966), .A4(n12965), .ZN(
        n12969) );
  NOR2_X1 U16236 ( .A1(n12970), .A2(n12969), .ZN(n14997) );
  AOI22_X1 U16237 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n10671), .B1(
        n10554), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n12974) );
  AOI22_X1 U16238 ( .A1(n10566), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10690), .B2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n12973) );
  AOI22_X1 U16239 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n13593), .B1(
        n10601), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n12972) );
  AOI22_X1 U16240 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n10567), .B1(
        n12725), .B2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n12971) );
  NAND4_X1 U16241 ( .A1(n12974), .A2(n12973), .A3(n12972), .A4(n12971), .ZN(
        n12981) );
  AOI22_X1 U16242 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n10676), .B1(
        n12952), .B2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n12979) );
  AOI22_X1 U16243 ( .A1(n10559), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        P2_INSTQUEUE_REG_2__7__SCAN_IN), .B2(n12975), .ZN(n12978) );
  AOI22_X1 U16244 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n10695), .B1(
        n10572), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n12977) );
  AOI22_X1 U16245 ( .A1(n12954), .A2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .B1(
        n12953), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n12976) );
  NAND4_X1 U16246 ( .A1(n12979), .A2(n12978), .A3(n12977), .A4(n12976), .ZN(
        n12980) );
  OR2_X1 U16247 ( .A1(n12981), .A2(n12980), .ZN(n13025) );
  INV_X1 U16248 ( .A(n10538), .ZN(n13148) );
  INV_X1 U16249 ( .A(P2_INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n12982) );
  OR2_X1 U16250 ( .A1(n13148), .A2(n12982), .ZN(n12986) );
  INV_X1 U16251 ( .A(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n20891) );
  OR2_X1 U16252 ( .A1(n13009), .A2(n20891), .ZN(n12985) );
  NAND2_X1 U16253 ( .A1(n10353), .A2(P2_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(
        n12984) );
  NAND2_X1 U16254 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(
        n12983) );
  AND4_X1 U16255 ( .A1(n12986), .A2(n12985), .A3(n12984), .A4(n12983), .ZN(
        n12989) );
  AOI22_X1 U16256 ( .A1(n9837), .A2(P2_INSTQUEUE_REG_5__0__SCAN_IN), .B1(n9827), .B2(P2_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n12988) );
  AOI22_X1 U16257 ( .A1(n13601), .A2(P2_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n10541), .B2(P2_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n12987) );
  XNOR2_X1 U16258 ( .A(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n13166) );
  NAND4_X1 U16259 ( .A1(n12989), .A2(n12988), .A3(n12987), .A4(n13166), .ZN(
        n13000) );
  INV_X1 U16260 ( .A(P2_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n12990) );
  OR2_X1 U16261 ( .A1(n13044), .A2(n12990), .ZN(n12995) );
  INV_X1 U16262 ( .A(P2_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n12991) );
  OR2_X1 U16263 ( .A1(n13009), .A2(n12991), .ZN(n12994) );
  NAND2_X1 U16264 ( .A1(n9825), .A2(P2_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(
        n12993) );
  NAND2_X1 U16265 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(
        n12992) );
  AND4_X1 U16266 ( .A1(n12995), .A2(n12994), .A3(n12993), .A4(n12992), .ZN(
        n12998) );
  AOI22_X1 U16267 ( .A1(n10538), .A2(P2_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n13601), .B2(P2_INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n12997) );
  AOI22_X1 U16268 ( .A1(n9827), .A2(P2_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n10541), .B2(P2_INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n12996) );
  INV_X1 U16269 ( .A(n13166), .ZN(n13170) );
  NAND4_X1 U16270 ( .A1(n12998), .A2(n12997), .A3(n12996), .A4(n13170), .ZN(
        n12999) );
  NAND2_X1 U16271 ( .A1(n13000), .A2(n12999), .ZN(n13029) );
  NOR2_X1 U16272 ( .A1(n16281), .A2(n13029), .ZN(n13001) );
  XOR2_X1 U16273 ( .A(n13025), .B(n13001), .Z(n13027) );
  XNOR2_X1 U16274 ( .A(n14998), .B(n13027), .ZN(n14990) );
  INV_X1 U16275 ( .A(n13029), .ZN(n13024) );
  NAND2_X1 U16276 ( .A1(n16281), .A2(n13024), .ZN(n14989) );
  INV_X1 U16277 ( .A(P2_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n13004) );
  INV_X1 U16278 ( .A(n13172), .ZN(n13152) );
  INV_X1 U16279 ( .A(P2_INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n13003) );
  OAI22_X1 U16280 ( .A1(n13148), .A2(n13004), .B1(n13152), .B2(n13003), .ZN(
        n13008) );
  INV_X1 U16281 ( .A(n13601), .ZN(n15540) );
  INV_X1 U16282 ( .A(P2_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n13006) );
  INV_X1 U16283 ( .A(n10541), .ZN(n13150) );
  OAI22_X1 U16284 ( .A1(n15540), .A2(n13006), .B1(n13150), .B2(n13005), .ZN(
        n13007) );
  NOR2_X1 U16285 ( .A1(n13008), .A2(n13007), .ZN(n13012) );
  AOI22_X1 U16286 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B1(n9825), .B2(P2_INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n13011) );
  AOI22_X1 U16287 ( .A1(n9837), .A2(P2_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n10540), .B2(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n13010) );
  NAND4_X1 U16288 ( .A1(n13012), .A2(n13011), .A3(n13010), .A4(n13166), .ZN(
        n13023) );
  INV_X1 U16289 ( .A(P2_INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n13014) );
  INV_X1 U16290 ( .A(P2_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n13013) );
  OAI22_X1 U16291 ( .A1(n13148), .A2(n13014), .B1(n13152), .B2(n13013), .ZN(
        n13018) );
  INV_X1 U16292 ( .A(P2_INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n13016) );
  OAI22_X1 U16293 ( .A1(n15540), .A2(n13016), .B1(n13150), .B2(n13015), .ZN(
        n13017) );
  NOR2_X1 U16294 ( .A1(n13018), .A2(n13017), .ZN(n13021) );
  AOI22_X1 U16295 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_14__1__SCAN_IN), .B1(
        n9825), .B2(P2_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n13020) );
  AOI22_X1 U16296 ( .A1(n9837), .A2(P2_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        n9833), .B2(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n13019) );
  NAND4_X1 U16297 ( .A1(n13021), .A2(n13170), .A3(n13020), .A4(n13019), .ZN(
        n13022) );
  NAND2_X1 U16298 ( .A1(n13023), .A2(n13022), .ZN(n13032) );
  NAND2_X1 U16299 ( .A1(n13025), .A2(n13024), .ZN(n13033) );
  XOR2_X1 U16300 ( .A(n13032), .B(n13033), .Z(n13026) );
  NAND2_X1 U16301 ( .A1(n13026), .A2(n13109), .ZN(n14978) );
  INV_X1 U16302 ( .A(n13027), .ZN(n13030) );
  INV_X1 U16303 ( .A(n13032), .ZN(n13028) );
  NAND2_X1 U16304 ( .A1(n16281), .A2(n13028), .ZN(n14981) );
  NOR3_X1 U16305 ( .A1(n13030), .A2(n13029), .A3(n14981), .ZN(n13031) );
  NOR2_X1 U16306 ( .A1(n13033), .A2(n13032), .ZN(n13054) );
  INV_X1 U16307 ( .A(P2_INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n21084) );
  INV_X1 U16308 ( .A(P2_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n13034) );
  OAI22_X1 U16309 ( .A1(n13148), .A2(n21084), .B1(n13152), .B2(n13034), .ZN(
        n13038) );
  INV_X1 U16310 ( .A(P2_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n13036) );
  INV_X1 U16311 ( .A(P2_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n13035) );
  OAI22_X1 U16312 ( .A1(n15540), .A2(n13036), .B1(n13150), .B2(n13035), .ZN(
        n13037) );
  NOR2_X1 U16313 ( .A1(n13038), .A2(n13037), .ZN(n13041) );
  AOI22_X1 U16314 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n10353), .B2(P2_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n13040) );
  INV_X1 U16315 ( .A(P2_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n19296) );
  AOI22_X1 U16316 ( .A1(n9837), .A2(P2_INSTQUEUE_REG_5__2__SCAN_IN), .B1(n9833), .B2(P2_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n13039) );
  NAND4_X1 U16317 ( .A1(n13041), .A2(n13040), .A3(n13039), .A4(n13166), .ZN(
        n13053) );
  INV_X1 U16318 ( .A(P2_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n13043) );
  INV_X1 U16319 ( .A(P2_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n13042) );
  OAI22_X1 U16320 ( .A1(n13044), .A2(n13043), .B1(n13152), .B2(n13042), .ZN(
        n13048) );
  INV_X1 U16321 ( .A(P2_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n13046) );
  INV_X1 U16322 ( .A(P2_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n13045) );
  OAI22_X1 U16323 ( .A1(n15540), .A2(n13046), .B1(n13150), .B2(n13045), .ZN(
        n13047) );
  NOR2_X1 U16324 ( .A1(n13048), .A2(n13047), .ZN(n13051) );
  AOI22_X1 U16325 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_14__2__SCAN_IN), .B1(
        n9825), .B2(P2_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n13050) );
  AOI22_X1 U16326 ( .A1(n10538), .A2(P2_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n10540), .B2(P2_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n13049) );
  NAND4_X1 U16327 ( .A1(n13051), .A2(n13170), .A3(n13050), .A4(n13049), .ZN(
        n13052) );
  AND2_X1 U16328 ( .A1(n13053), .A2(n13052), .ZN(n13055) );
  NAND2_X1 U16329 ( .A1(n13054), .A2(n13055), .ZN(n13106) );
  OAI211_X1 U16330 ( .C1(n13054), .C2(n13055), .A(n13109), .B(n13106), .ZN(
        n13057) );
  INV_X1 U16331 ( .A(n13055), .ZN(n13056) );
  NOR2_X1 U16332 ( .A1(n13334), .A2(n13056), .ZN(n14969) );
  INV_X1 U16333 ( .A(P2_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n13061) );
  INV_X1 U16334 ( .A(P2_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n13060) );
  OAI22_X1 U16335 ( .A1(n13148), .A2(n13061), .B1(n13152), .B2(n13060), .ZN(
        n13065) );
  INV_X1 U16336 ( .A(P2_INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n13063) );
  INV_X1 U16337 ( .A(P2_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n13062) );
  OAI22_X1 U16338 ( .A1(n15540), .A2(n13063), .B1(n13150), .B2(n13062), .ZN(
        n13064) );
  NOR2_X1 U16339 ( .A1(n13065), .A2(n13064), .ZN(n13068) );
  AOI22_X1 U16340 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_6__3__SCAN_IN), .B1(
        n10353), .B2(P2_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n13067) );
  AOI22_X1 U16341 ( .A1(n9837), .A2(P2_INSTQUEUE_REG_5__3__SCAN_IN), .B1(n9833), .B2(P2_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n13066) );
  NAND4_X1 U16342 ( .A1(n13068), .A2(n13067), .A3(n13066), .A4(n13166), .ZN(
        n13079) );
  INV_X1 U16343 ( .A(P2_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n13070) );
  INV_X1 U16344 ( .A(P2_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n13069) );
  OAI22_X1 U16345 ( .A1(n13148), .A2(n13070), .B1(n13152), .B2(n13069), .ZN(
        n13074) );
  INV_X1 U16346 ( .A(P2_INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n13071) );
  OAI22_X1 U16347 ( .A1(n15540), .A2(n13072), .B1(n13150), .B2(n13071), .ZN(
        n13073) );
  NOR2_X1 U16348 ( .A1(n13074), .A2(n13073), .ZN(n13077) );
  AOI22_X1 U16349 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n9825), .B2(P2_INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n13076) );
  AOI22_X1 U16350 ( .A1(n9837), .A2(P2_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n10540), .B2(P2_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n13075) );
  NAND4_X1 U16351 ( .A1(n13077), .A2(n13170), .A3(n13076), .A4(n13075), .ZN(
        n13078) );
  AND2_X1 U16352 ( .A1(n13079), .A2(n13078), .ZN(n13104) );
  XNOR2_X1 U16353 ( .A(n13106), .B(n13104), .ZN(n13080) );
  NAND2_X1 U16354 ( .A1(n16281), .A2(n13104), .ZN(n14963) );
  NAND2_X1 U16355 ( .A1(n13081), .A2(n10308), .ZN(n13082) );
  INV_X1 U16356 ( .A(P2_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n13085) );
  INV_X1 U16357 ( .A(P2_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n13084) );
  OAI22_X1 U16358 ( .A1(n13148), .A2(n13085), .B1(n13152), .B2(n13084), .ZN(
        n13089) );
  INV_X1 U16359 ( .A(P2_INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n13087) );
  INV_X1 U16360 ( .A(P2_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n13086) );
  OAI22_X1 U16361 ( .A1(n15540), .A2(n13087), .B1(n13150), .B2(n13086), .ZN(
        n13088) );
  NOR2_X1 U16362 ( .A1(n13089), .A2(n13088), .ZN(n13092) );
  AOI22_X1 U16363 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n10353), .B2(P2_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n13091) );
  AOI22_X1 U16364 ( .A1(n9837), .A2(P2_INSTQUEUE_REG_5__4__SCAN_IN), .B1(
        n10540), .B2(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13090) );
  NAND4_X1 U16365 ( .A1(n13092), .A2(n13091), .A3(n13090), .A4(n13166), .ZN(
        n13103) );
  INV_X1 U16366 ( .A(P2_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n13094) );
  INV_X1 U16367 ( .A(P2_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n13093) );
  OAI22_X1 U16368 ( .A1(n13148), .A2(n13094), .B1(n13152), .B2(n13093), .ZN(
        n13098) );
  INV_X1 U16369 ( .A(P2_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n13096) );
  INV_X1 U16370 ( .A(P2_INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n13095) );
  OAI22_X1 U16371 ( .A1(n15540), .A2(n13096), .B1(n13150), .B2(n13095), .ZN(
        n13097) );
  NOR2_X1 U16372 ( .A1(n13098), .A2(n13097), .ZN(n13101) );
  AOI22_X1 U16373 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9825), .B2(P2_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n13100) );
  AOI22_X1 U16374 ( .A1(n9837), .A2(P2_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n9833), .B2(P2_INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n13099) );
  NAND4_X1 U16375 ( .A1(n13101), .A2(n13170), .A3(n13100), .A4(n13099), .ZN(
        n13102) );
  NAND2_X1 U16376 ( .A1(n13103), .A2(n13102), .ZN(n13107) );
  INV_X1 U16377 ( .A(n13107), .ZN(n13114) );
  INV_X1 U16378 ( .A(n13104), .ZN(n13105) );
  OR2_X1 U16379 ( .A1(n13106), .A2(n13105), .ZN(n13108) );
  INV_X1 U16380 ( .A(n13108), .ZN(n13110) );
  OR2_X1 U16381 ( .A1(n13108), .A2(n13107), .ZN(n14943) );
  OAI211_X1 U16382 ( .C1(n13114), .C2(n13110), .A(n14943), .B(n13109), .ZN(
        n13111) );
  NAND2_X1 U16383 ( .A1(n16281), .A2(n13114), .ZN(n14955) );
  INV_X1 U16384 ( .A(n14944), .ZN(n13135) );
  INV_X1 U16385 ( .A(P2_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n13116) );
  INV_X1 U16386 ( .A(P2_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n13115) );
  OAI22_X1 U16387 ( .A1(n13148), .A2(n13116), .B1(n13152), .B2(n13115), .ZN(
        n13120) );
  INV_X1 U16388 ( .A(P2_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n13118) );
  INV_X1 U16389 ( .A(P2_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n13117) );
  OAI22_X1 U16390 ( .A1(n15540), .A2(n13118), .B1(n13150), .B2(n13117), .ZN(
        n13119) );
  NOR2_X1 U16391 ( .A1(n13120), .A2(n13119), .ZN(n13123) );
  AOI22_X1 U16392 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_6__5__SCAN_IN), .B1(n9825), .B2(P2_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n13122) );
  AOI22_X1 U16393 ( .A1(n9837), .A2(P2_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n9833), .B2(P2_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n13121) );
  NAND4_X1 U16394 ( .A1(n13123), .A2(n13122), .A3(n13121), .A4(n13166), .ZN(
        n13134) );
  INV_X1 U16395 ( .A(P2_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n13125) );
  INV_X1 U16396 ( .A(P2_INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n13124) );
  OAI22_X1 U16397 ( .A1(n13148), .A2(n13125), .B1(n13152), .B2(n13124), .ZN(
        n13129) );
  INV_X1 U16398 ( .A(P2_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n13127) );
  INV_X1 U16399 ( .A(P2_INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n13126) );
  OAI22_X1 U16400 ( .A1(n15540), .A2(n13127), .B1(n13150), .B2(n13126), .ZN(
        n13128) );
  NOR2_X1 U16401 ( .A1(n13129), .A2(n13128), .ZN(n13132) );
  AOI22_X1 U16402 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9825), .B2(P2_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n13131) );
  AOI22_X1 U16403 ( .A1(n9837), .A2(P2_INSTQUEUE_REG_13__5__SCAN_IN), .B1(
        n10540), .B2(P2_INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n13130) );
  NAND4_X1 U16404 ( .A1(n13132), .A2(n13170), .A3(n13131), .A4(n13130), .ZN(
        n13133) );
  AND2_X1 U16405 ( .A1(n13134), .A2(n13133), .ZN(n14945) );
  NAND2_X1 U16406 ( .A1(n13334), .A2(n14945), .ZN(n13136) );
  NOR2_X1 U16407 ( .A1(n14943), .A2(n13136), .ZN(n13161) );
  INV_X1 U16408 ( .A(P2_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n13138) );
  INV_X1 U16409 ( .A(P2_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n13137) );
  OAI22_X1 U16410 ( .A1(n13148), .A2(n13138), .B1(n13152), .B2(n13137), .ZN(
        n13142) );
  INV_X1 U16411 ( .A(P2_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n13140) );
  INV_X1 U16412 ( .A(P2_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n13139) );
  OAI22_X1 U16413 ( .A1(n15540), .A2(n13140), .B1(n13150), .B2(n13139), .ZN(
        n13141) );
  NOR2_X1 U16414 ( .A1(n13142), .A2(n13141), .ZN(n13145) );
  AOI22_X1 U16415 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_6__6__SCAN_IN), .B1(n9825), .B2(P2_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n13144) );
  AOI22_X1 U16416 ( .A1(n9837), .A2(P2_INSTQUEUE_REG_5__6__SCAN_IN), .B1(n9833), .B2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n13143) );
  NAND4_X1 U16417 ( .A1(n13145), .A2(n13144), .A3(n13143), .A4(n13166), .ZN(
        n13159) );
  INV_X1 U16418 ( .A(P2_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n13147) );
  INV_X1 U16419 ( .A(P2_INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n13146) );
  OAI22_X1 U16420 ( .A1(n13148), .A2(n13147), .B1(n15540), .B2(n13146), .ZN(
        n13154) );
  INV_X1 U16421 ( .A(P2_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n13151) );
  INV_X1 U16422 ( .A(P2_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n13149) );
  OAI22_X1 U16423 ( .A1(n13152), .A2(n13151), .B1(n13150), .B2(n13149), .ZN(
        n13153) );
  NOR2_X1 U16424 ( .A1(n13154), .A2(n13153), .ZN(n13157) );
  AOI22_X1 U16425 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n10353), .B2(P2_INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n13156) );
  AOI22_X1 U16426 ( .A1(n9837), .A2(P2_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n10540), .B2(P2_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n13155) );
  NAND4_X1 U16427 ( .A1(n13157), .A2(n13170), .A3(n13156), .A4(n13155), .ZN(
        n13158) );
  AND2_X1 U16428 ( .A1(n13159), .A2(n13158), .ZN(n13160) );
  NAND2_X1 U16429 ( .A1(n13161), .A2(n13160), .ZN(n13162) );
  OAI21_X1 U16430 ( .B1(n13161), .B2(n13160), .A(n13162), .ZN(n14939) );
  NOR2_X1 U16431 ( .A1(n14940), .A2(n14939), .ZN(n14938) );
  INV_X1 U16432 ( .A(n13162), .ZN(n13163) );
  NOR2_X1 U16433 ( .A1(n14938), .A2(n13163), .ZN(n13180) );
  AOI22_X1 U16434 ( .A1(n10538), .A2(P2_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n13172), .B2(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n13165) );
  AOI22_X1 U16435 ( .A1(n13601), .A2(P2_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n10541), .B2(P2_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n13164) );
  NAND2_X1 U16436 ( .A1(n13165), .A2(n13164), .ZN(n13178) );
  AOI22_X1 U16437 ( .A1(n9837), .A2(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B1(
        n10540), .B2(P2_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n13168) );
  AOI22_X1 U16438 ( .A1(n10401), .A2(P2_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n10353), .B2(P2_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n13167) );
  NAND3_X1 U16439 ( .A1(n13168), .A2(n13167), .A3(n13166), .ZN(n13177) );
  AOI22_X1 U16440 ( .A1(n9837), .A2(P2_INSTQUEUE_REG_13__7__SCAN_IN), .B1(
        n9833), .B2(P2_INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n13171) );
  AOI22_X1 U16441 ( .A1(n9834), .A2(P2_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n9825), .B2(P2_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n13169) );
  NAND3_X1 U16442 ( .A1(n13171), .A2(n13170), .A3(n13169), .ZN(n13176) );
  AOI22_X1 U16443 ( .A1(n10538), .A2(P2_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n10541), .B2(P2_INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n13174) );
  AOI22_X1 U16444 ( .A1(n9827), .A2(P2_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n13601), .B2(P2_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n13173) );
  NAND2_X1 U16445 ( .A1(n13174), .A2(n13173), .ZN(n13175) );
  OAI22_X1 U16446 ( .A1(n13178), .A2(n13177), .B1(n13176), .B2(n13175), .ZN(
        n13179) );
  XNOR2_X1 U16447 ( .A(n13180), .B(n13179), .ZN(n15015) );
  OR2_X1 U16448 ( .A1(n16257), .A2(n13591), .ZN(n13610) );
  INV_X1 U16449 ( .A(n13181), .ZN(n13597) );
  NAND2_X1 U16450 ( .A1(n13610), .A2(n13597), .ZN(n13182) );
  NAND2_X1 U16451 ( .A1(n16018), .A2(n14993), .ZN(n13184) );
  NAND2_X1 U16452 ( .A1(n15006), .A2(P2_EBX_REG_30__SCAN_IN), .ZN(n13183) );
  OAI21_X1 U16453 ( .B1(n15015), .B2(n15009), .A(n10290), .ZN(P2_U2857) );
  NOR2_X1 U16454 ( .A1(P2_BE_N_REG_0__SCAN_IN), .A2(P2_BE_N_REG_1__SCAN_IN), 
        .ZN(n13186) );
  NOR4_X1 U16455 ( .A1(P2_BE_N_REG_2__SCAN_IN), .A2(P2_BE_N_REG_3__SCAN_IN), 
        .A3(P2_D_C_N_REG_SCAN_IN), .A4(P2_ADS_N_REG_SCAN_IN), .ZN(n13185) );
  NAND4_X1 U16456 ( .A1(P2_M_IO_N_REG_SCAN_IN), .A2(P2_W_R_N_REG_SCAN_IN), 
        .A3(n13186), .A4(n13185), .ZN(n13209) );
  NOR2_X1 U16457 ( .A1(P2_ADDRESS_REG_29__SCAN_IN), .A2(n13209), .ZN(n16422)
         );
  NOR4_X1 U16458 ( .A1(P1_ADDRESS_REG_14__SCAN_IN), .A2(
        P1_ADDRESS_REG_13__SCAN_IN), .A3(P1_ADDRESS_REG_12__SCAN_IN), .A4(
        P1_ADDRESS_REG_11__SCAN_IN), .ZN(n13190) );
  NOR4_X1 U16459 ( .A1(P1_ADDRESS_REG_19__SCAN_IN), .A2(
        P1_ADDRESS_REG_18__SCAN_IN), .A3(P1_ADDRESS_REG_17__SCAN_IN), .A4(
        P1_ADDRESS_REG_15__SCAN_IN), .ZN(n13189) );
  NOR4_X1 U16460 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(
        P1_ADDRESS_REG_5__SCAN_IN), .A3(P1_ADDRESS_REG_4__SCAN_IN), .A4(
        P1_ADDRESS_REG_3__SCAN_IN), .ZN(n13188) );
  NOR4_X1 U16461 ( .A1(P1_ADDRESS_REG_10__SCAN_IN), .A2(
        P1_ADDRESS_REG_9__SCAN_IN), .A3(P1_ADDRESS_REG_8__SCAN_IN), .A4(
        P1_ADDRESS_REG_7__SCAN_IN), .ZN(n13187) );
  AND4_X1 U16462 ( .A1(n13190), .A2(n13189), .A3(n13188), .A4(n13187), .ZN(
        n13195) );
  NOR4_X1 U16463 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(
        P1_ADDRESS_REG_0__SCAN_IN), .A3(P1_ADDRESS_REG_16__SCAN_IN), .A4(
        P1_ADDRESS_REG_28__SCAN_IN), .ZN(n13193) );
  NOR4_X1 U16464 ( .A1(P1_ADDRESS_REG_23__SCAN_IN), .A2(
        P1_ADDRESS_REG_22__SCAN_IN), .A3(P1_ADDRESS_REG_21__SCAN_IN), .A4(
        P1_ADDRESS_REG_20__SCAN_IN), .ZN(n13192) );
  NOR4_X1 U16465 ( .A1(P1_ADDRESS_REG_27__SCAN_IN), .A2(
        P1_ADDRESS_REG_26__SCAN_IN), .A3(P1_ADDRESS_REG_25__SCAN_IN), .A4(
        P1_ADDRESS_REG_24__SCAN_IN), .ZN(n13191) );
  INV_X1 U16466 ( .A(P1_ADDRESS_REG_2__SCAN_IN), .ZN(n20711) );
  AND4_X1 U16467 ( .A1(n13193), .A2(n13192), .A3(n13191), .A4(n20711), .ZN(
        n13194) );
  NAND2_X1 U16468 ( .A1(n13195), .A2(n13194), .ZN(n13196) );
  AND2_X2 U16469 ( .A1(n13196), .A2(P1_ADDRESS_REG_29__SCAN_IN), .ZN(n14173)
         );
  INV_X1 U16470 ( .A(P1_W_R_N_REG_SCAN_IN), .ZN(n20785) );
  NOR3_X1 U16471 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(P1_BE_N_REG_0__SCAN_IN), 
        .A3(n20785), .ZN(n13198) );
  NOR4_X1 U16472 ( .A1(P1_BE_N_REG_1__SCAN_IN), .A2(P1_BE_N_REG_3__SCAN_IN), 
        .A3(P1_D_C_N_REG_SCAN_IN), .A4(P1_ADS_N_REG_SCAN_IN), .ZN(n13197) );
  NAND4_X1 U16473 ( .A1(n14173), .A2(P1_M_IO_N_REG_SCAN_IN), .A3(n13198), .A4(
        n13197), .ZN(U214) );
  NOR4_X1 U16474 ( .A1(P2_ADDRESS_REG_17__SCAN_IN), .A2(
        P2_ADDRESS_REG_16__SCAN_IN), .A3(P2_ADDRESS_REG_15__SCAN_IN), .A4(
        P2_ADDRESS_REG_14__SCAN_IN), .ZN(n13202) );
  NOR4_X1 U16475 ( .A1(P2_ADDRESS_REG_21__SCAN_IN), .A2(
        P2_ADDRESS_REG_20__SCAN_IN), .A3(P2_ADDRESS_REG_19__SCAN_IN), .A4(
        P2_ADDRESS_REG_18__SCAN_IN), .ZN(n13201) );
  NOR4_X1 U16476 ( .A1(P2_ADDRESS_REG_8__SCAN_IN), .A2(
        P2_ADDRESS_REG_7__SCAN_IN), .A3(P2_ADDRESS_REG_6__SCAN_IN), .A4(
        P2_ADDRESS_REG_4__SCAN_IN), .ZN(n13200) );
  NOR4_X1 U16477 ( .A1(P2_ADDRESS_REG_13__SCAN_IN), .A2(
        P2_ADDRESS_REG_12__SCAN_IN), .A3(P2_ADDRESS_REG_11__SCAN_IN), .A4(
        P2_ADDRESS_REG_9__SCAN_IN), .ZN(n13199) );
  NAND4_X1 U16478 ( .A1(n13202), .A2(n13201), .A3(n13200), .A4(n13199), .ZN(
        n13207) );
  NOR4_X1 U16479 ( .A1(P2_ADDRESS_REG_1__SCAN_IN), .A2(
        P2_ADDRESS_REG_0__SCAN_IN), .A3(P2_ADDRESS_REG_5__SCAN_IN), .A4(
        P2_ADDRESS_REG_10__SCAN_IN), .ZN(n13205) );
  NOR4_X1 U16480 ( .A1(P2_ADDRESS_REG_25__SCAN_IN), .A2(
        P2_ADDRESS_REG_24__SCAN_IN), .A3(P2_ADDRESS_REG_23__SCAN_IN), .A4(
        P2_ADDRESS_REG_22__SCAN_IN), .ZN(n13204) );
  NOR4_X1 U16481 ( .A1(P2_ADDRESS_REG_3__SCAN_IN), .A2(
        P2_ADDRESS_REG_27__SCAN_IN), .A3(P2_ADDRESS_REG_28__SCAN_IN), .A4(
        P2_ADDRESS_REG_26__SCAN_IN), .ZN(n13203) );
  INV_X1 U16482 ( .A(P2_ADDRESS_REG_2__SCAN_IN), .ZN(n19738) );
  NAND4_X1 U16483 ( .A1(n13205), .A2(n13204), .A3(n13203), .A4(n19738), .ZN(
        n13206) );
  OAI21_X1 U16484 ( .B1(n13207), .B2(n13206), .A(P2_ADDRESS_REG_29__SCAN_IN), 
        .ZN(n13208) );
  NOR2_X1 U16485 ( .A1(n14070), .A2(n13209), .ZN(n16360) );
  NAND2_X1 U16486 ( .A1(n16360), .A2(U214), .ZN(U212) );
  OAI21_X1 U16487 ( .B1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n13211), .A(
        n14867), .ZN(n15199) );
  INV_X1 U16488 ( .A(n15199), .ZN(n13232) );
  NOR2_X1 U16489 ( .A1(n13227), .A2(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(
        n13210) );
  NOR2_X1 U16490 ( .A1(n13211), .A2(n13210), .ZN(n18792) );
  AOI21_X1 U16491 ( .B1(n18819), .B2(n9914), .A(n13225), .ZN(n18818) );
  AOI21_X1 U16492 ( .B1(n15253), .B2(n13222), .A(n13224), .ZN(n15252) );
  AOI21_X1 U16493 ( .B1(n16144), .B2(n13221), .A(n13223), .ZN(n18863) );
  AOI21_X1 U16494 ( .B1(n16157), .B2(n13219), .A(n9909), .ZN(n18888) );
  AOI21_X1 U16495 ( .B1(n14217), .B2(n13217), .A(n13220), .ZN(n14216) );
  AOI21_X1 U16496 ( .B1(n14082), .B2(n13215), .A(n13218), .ZN(n18906) );
  AOI21_X1 U16497 ( .B1(n16191), .B2(n13213), .A(n13216), .ZN(n18930) );
  AOI21_X1 U16498 ( .B1(n14901), .B2(n13212), .A(n13214), .ZN(n14900) );
  OAI22_X1 U16499 ( .A1(n10983), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(P2_STATE2_REG_0__SCAN_IN), .ZN(
        n14927) );
  INV_X1 U16500 ( .A(n14927), .ZN(n18942) );
  AOI22_X1 U16501 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n15530), .B1(
        P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n10983), .ZN(n14924) );
  NOR2_X1 U16502 ( .A1(n18942), .A2(n14924), .ZN(n14918) );
  OAI21_X1 U16503 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n13212), .ZN(n14920) );
  NAND2_X1 U16504 ( .A1(n14918), .A2(n14920), .ZN(n14898) );
  NOR2_X1 U16505 ( .A1(n14900), .A2(n14898), .ZN(n14028) );
  OAI21_X1 U16506 ( .B1(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n13214), .A(
        n13213), .ZN(n19097) );
  NAND2_X1 U16507 ( .A1(n14028), .A2(n19097), .ZN(n18928) );
  NOR2_X1 U16508 ( .A1(n18930), .A2(n18928), .ZN(n18916) );
  OAI21_X1 U16509 ( .B1(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n13216), .A(
        n13215), .ZN(n18919) );
  NAND2_X1 U16510 ( .A1(n18916), .A2(n18919), .ZN(n18905) );
  NOR2_X1 U16511 ( .A1(n18906), .A2(n18905), .ZN(n14043) );
  OAI21_X1 U16512 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n13218), .A(
        n13217), .ZN(n16178) );
  NAND2_X1 U16513 ( .A1(n14043), .A2(n16178), .ZN(n14885) );
  NOR2_X1 U16514 ( .A1(n14216), .A2(n14885), .ZN(n18895) );
  OAI21_X1 U16515 ( .B1(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n13220), .A(
        n13219), .ZN(n18897) );
  NAND2_X1 U16516 ( .A1(n18895), .A2(n18897), .ZN(n18886) );
  NOR2_X1 U16517 ( .A1(n18888), .A2(n18886), .ZN(n18868) );
  OAI21_X1 U16518 ( .B1(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n9909), .A(
        n13221), .ZN(n18869) );
  NAND2_X1 U16519 ( .A1(n18868), .A2(n18869), .ZN(n18854) );
  NOR2_X1 U16520 ( .A1(n18863), .A2(n18854), .ZN(n18853) );
  OAI21_X1 U16521 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n13223), .A(
        n13222), .ZN(n16138) );
  NAND2_X1 U16522 ( .A1(n18853), .A2(n16138), .ZN(n18844) );
  NOR2_X1 U16523 ( .A1(n15252), .A2(n18844), .ZN(n18828) );
  OAI21_X1 U16524 ( .B1(P2_PHYADDRPOINTER_REG_16__SCAN_IN), .B2(n13224), .A(
        n9914), .ZN(n18829) );
  NAND2_X1 U16525 ( .A1(n18828), .A2(n18829), .ZN(n18816) );
  NOR2_X1 U16526 ( .A1(n18818), .A2(n18816), .ZN(n18804) );
  NOR2_X1 U16527 ( .A1(n13225), .A2(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n13226) );
  OR2_X1 U16528 ( .A1(n13227), .A2(n13226), .ZN(n18805) );
  NAND2_X1 U16529 ( .A1(n18804), .A2(n18805), .ZN(n18790) );
  OR2_X1 U16530 ( .A1(n18792), .A2(n18790), .ZN(n13229) );
  NAND4_X1 U16531 ( .A1(n19842), .A2(n10983), .A3(n19836), .A4(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19714) );
  INV_X1 U16532 ( .A(n19714), .ZN(n18890) );
  NAND2_X1 U16533 ( .A1(n18890), .A2(n18929), .ZN(n18852) );
  NOR2_X1 U16534 ( .A1(n13229), .A2(n13232), .ZN(n14868) );
  OR2_X1 U16535 ( .A1(n18852), .A2(n14868), .ZN(n14880) );
  AOI21_X1 U16536 ( .B1(n13232), .B2(n13229), .A(n14880), .ZN(n13255) );
  NOR2_X1 U16537 ( .A1(n16255), .A2(n16253), .ZN(n13381) );
  NOR2_X1 U16538 ( .A1(n19798), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19708) );
  INV_X1 U16539 ( .A(n19708), .ZN(n13230) );
  NOR2_X1 U16540 ( .A1(n19707), .A2(n13230), .ZN(n16276) );
  NAND2_X1 U16541 ( .A1(n19714), .A2(n18934), .ZN(n13231) );
  NAND2_X1 U16542 ( .A1(n18954), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n18831) );
  NOR2_X1 U16543 ( .A1(n18929), .A2(n19714), .ZN(n18864) );
  AOI22_X1 U16544 ( .A1(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n18958), .B1(
        n13232), .B2(n18864), .ZN(n13233) );
  INV_X1 U16545 ( .A(n13233), .ZN(n13254) );
  NOR2_X1 U16546 ( .A1(P2_STATEBS16_REG_SCAN_IN), .A2(n19843), .ZN(n13245) );
  INV_X1 U16547 ( .A(n13245), .ZN(n13237) );
  NOR2_X1 U16548 ( .A1(n9839), .A2(n13237), .ZN(n13234) );
  NAND2_X1 U16549 ( .A1(n19847), .A2(n13234), .ZN(n18937) );
  OAI21_X1 U16550 ( .B1(n13235), .B2(n13236), .A(n14870), .ZN(n15362) );
  NAND2_X1 U16551 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n13237), .ZN(n13238) );
  NOR2_X1 U16552 ( .A1(n9839), .A2(n13238), .ZN(n13239) );
  NAND2_X1 U16553 ( .A1(n19847), .A2(n13239), .ZN(n18947) );
  NAND2_X1 U16554 ( .A1(n13240), .A2(n18933), .ZN(n13252) );
  OR2_X1 U16555 ( .A1(n12660), .A2(n16292), .ZN(n13241) );
  NAND2_X1 U16556 ( .A1(n13611), .A2(n19836), .ZN(n16007) );
  INV_X1 U16557 ( .A(n16007), .ZN(n16280) );
  INV_X1 U16558 ( .A(n18945), .ZN(n18877) );
  NOR2_X1 U16559 ( .A1(n9916), .A2(n13243), .ZN(n13244) );
  NOR2_X1 U16560 ( .A1(n13242), .A2(n13244), .ZN(n16113) );
  NAND2_X1 U16561 ( .A1(n19081), .A2(n16007), .ZN(n13249) );
  INV_X1 U16562 ( .A(n13289), .ZN(n13247) );
  NOR2_X1 U16563 ( .A1(P2_EBX_REG_31__SCAN_IN), .A2(n13245), .ZN(n13246) );
  NAND2_X1 U16564 ( .A1(n13247), .A2(n13246), .ZN(n13248) );
  INV_X1 U16565 ( .A(n18951), .ZN(n18840) );
  INV_X1 U16566 ( .A(P2_EBX_REG_20__SCAN_IN), .ZN(n20952) );
  OAI22_X1 U16567 ( .A1(n18840), .A2(n20952), .B1(n19756), .B2(n18954), .ZN(
        n13250) );
  AOI21_X1 U16568 ( .B1(n18877), .B2(n16113), .A(n13250), .ZN(n13251) );
  OAI211_X1 U16569 ( .C1(n18937), .C2(n15362), .A(n13252), .B(n13251), .ZN(
        n13253) );
  OR3_X1 U16570 ( .A1(n13255), .A2(n13254), .A3(n13253), .ZN(P2_U2835) );
  OR2_X1 U16571 ( .A1(n12599), .A2(n16292), .ZN(n19014) );
  NOR2_X1 U16572 ( .A1(n16255), .A2(n19014), .ZN(n18957) );
  INV_X1 U16573 ( .A(P2_MEMORYFETCH_REG_SCAN_IN), .ZN(n13256) );
  OAI211_X1 U16574 ( .C1(n18957), .C2(n13256), .A(n18766), .B(n13289), .ZN(
        P2_U2814) );
  NOR2_X1 U16575 ( .A1(n19847), .A2(P2_READREQUEST_REG_SCAN_IN), .ZN(n13258)
         );
  INV_X1 U16576 ( .A(n12636), .ZN(n13257) );
  AOI22_X1 U16577 ( .A1(n13258), .A2(n18766), .B1(n13257), .B2(n19847), .ZN(
        P2_U3612) );
  AND2_X1 U16578 ( .A1(n12636), .A2(n19849), .ZN(n13380) );
  NOR2_X1 U16579 ( .A1(n13380), .A2(n13611), .ZN(n13259) );
  AND2_X1 U16580 ( .A1(n13381), .A2(n13259), .ZN(n16265) );
  NOR2_X1 U16581 ( .A1(n16265), .A2(n16292), .ZN(n19833) );
  INV_X1 U16582 ( .A(P2_FLUSH_REG_SCAN_IN), .ZN(n15741) );
  OAI21_X1 U16583 ( .B1(n19833), .B2(n15741), .A(n13260), .ZN(P2_U2819) );
  NOR2_X2 U16584 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n20581) );
  NAND2_X1 U16585 ( .A1(n20581), .A2(n16000), .ZN(n19860) );
  INV_X1 U16586 ( .A(n19860), .ZN(n13278) );
  AOI211_X1 U16587 ( .C1(P1_MEMORYFETCH_REG_SCAN_IN), .C2(n13261), .A(n13278), 
        .B(n13282), .ZN(n13262) );
  INV_X1 U16588 ( .A(n13262), .ZN(P1_U2801) );
  INV_X1 U16589 ( .A(n11596), .ZN(n15692) );
  NAND2_X1 U16590 ( .A1(n13263), .A2(n15692), .ZN(n13264) );
  OAI21_X1 U16591 ( .B1(n13698), .B2(n13265), .A(n13264), .ZN(n19858) );
  NAND3_X1 U16592 ( .A1(n14427), .A2(n15736), .A3(n13516), .ZN(n13266) );
  AND2_X1 U16593 ( .A1(n13266), .A2(n15993), .ZN(n20792) );
  NOR2_X1 U16594 ( .A1(n19858), .A2(n20792), .ZN(n15711) );
  NOR2_X1 U16595 ( .A1(n15711), .A2(n19857), .ZN(n19865) );
  INV_X1 U16596 ( .A(P1_MORE_REG_SCAN_IN), .ZN(n13277) );
  INV_X1 U16597 ( .A(n13267), .ZN(n13268) );
  NAND2_X1 U16598 ( .A1(n13268), .A2(n14427), .ZN(n13270) );
  AOI21_X1 U16599 ( .B1(n13271), .B2(n13270), .A(n13269), .ZN(n13273) );
  OAI22_X1 U16600 ( .A1(n13698), .A2(n13273), .B1(n13472), .B2(n13272), .ZN(
        n13274) );
  AOI21_X1 U16601 ( .B1(n13658), .B2(n13698), .A(n13274), .ZN(n13275) );
  INV_X1 U16602 ( .A(n20145), .ZN(n14503) );
  NOR2_X1 U16603 ( .A1(n13275), .A2(n14503), .ZN(n15710) );
  NAND2_X1 U16604 ( .A1(n19865), .A2(n15710), .ZN(n13276) );
  OAI21_X1 U16605 ( .B1(n19865), .B2(n13277), .A(n13276), .ZN(P1_U3484) );
  OAI21_X1 U16606 ( .B1(n13278), .B2(P1_READREQUEST_REG_SCAN_IN), .A(n20789), 
        .ZN(n13279) );
  OAI21_X1 U16607 ( .B1(n13280), .B2(n20789), .A(n13279), .ZN(P1_U3487) );
  NAND2_X1 U16608 ( .A1(n13282), .A2(n13281), .ZN(n20035) );
  INV_X1 U16609 ( .A(P1_EAX_REG_15__SCAN_IN), .ZN(n19971) );
  INV_X1 U16610 ( .A(n15993), .ZN(n20791) );
  AND2_X1 U16611 ( .A1(n20793), .A2(n20791), .ZN(n13283) );
  NAND2_X1 U16612 ( .A1(n13416), .A2(n20122), .ZN(n20016) );
  INV_X1 U16613 ( .A(DATAI_15_), .ZN(n13286) );
  INV_X1 U16614 ( .A(BUF1_REG_15__SCAN_IN), .ZN(n13285) );
  MUX2_X1 U16615 ( .A(n13286), .B(n13285), .S(n14173), .Z(n14154) );
  INV_X1 U16616 ( .A(P1_LWORD_REG_15__SCAN_IN), .ZN(n13287) );
  OAI222_X1 U16617 ( .A1(n20035), .A2(n19971), .B1(n20016), .B2(n14154), .C1(
        n13416), .C2(n13287), .ZN(P1_U2967) );
  NOR2_X1 U16618 ( .A1(n13289), .A2(n19843), .ZN(n13288) );
  INV_X1 U16619 ( .A(P2_UWORD_REG_1__SCAN_IN), .ZN(n13291) );
  NOR3_X2 U16620 ( .A1(n13289), .A2(n16281), .A3(n19843), .ZN(n13448) );
  INV_X1 U16621 ( .A(n13448), .ZN(n13359) );
  AOI22_X1 U16622 ( .A1(n14069), .A2(BUF1_REG_1__SCAN_IN), .B1(
        BUF2_REG_1__SCAN_IN), .B2(n14070), .ZN(n19119) );
  NOR2_X1 U16623 ( .A1(n13359), .A2(n19119), .ZN(n13302) );
  AOI21_X1 U16624 ( .B1(n19081), .B2(P2_EAX_REG_17__SCAN_IN), .A(n13302), .ZN(
        n13290) );
  OAI21_X1 U16625 ( .B1(n13429), .B2(n13291), .A(n13290), .ZN(P2_U2953) );
  INV_X1 U16626 ( .A(P2_UWORD_REG_2__SCAN_IN), .ZN(n13293) );
  OAI22_X1 U16627 ( .A1(n14070), .A2(BUF1_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n14069), .ZN(n19125) );
  NOR2_X1 U16628 ( .A1(n13359), .A2(n19125), .ZN(n13305) );
  AOI21_X1 U16629 ( .B1(n19081), .B2(P2_EAX_REG_18__SCAN_IN), .A(n13305), .ZN(
        n13292) );
  OAI21_X1 U16630 ( .B1(n13429), .B2(n13293), .A(n13292), .ZN(P2_U2954) );
  INV_X1 U16631 ( .A(P2_UWORD_REG_3__SCAN_IN), .ZN(n13295) );
  AOI22_X1 U16632 ( .A1(n14069), .A2(BUF1_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n14070), .ZN(n19130) );
  NOR2_X1 U16633 ( .A1(n13359), .A2(n19130), .ZN(n13308) );
  AOI21_X1 U16634 ( .B1(n19081), .B2(P2_EAX_REG_19__SCAN_IN), .A(n13308), .ZN(
        n13294) );
  OAI21_X1 U16635 ( .B1(n13429), .B2(n13295), .A(n13294), .ZN(P2_U2955) );
  INV_X1 U16636 ( .A(P2_UWORD_REG_5__SCAN_IN), .ZN(n13297) );
  AOI22_X1 U16637 ( .A1(n14069), .A2(BUF1_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n14070), .ZN(n19135) );
  NOR2_X1 U16638 ( .A1(n13359), .A2(n19135), .ZN(n13314) );
  AOI21_X1 U16639 ( .B1(n19081), .B2(P2_EAX_REG_21__SCAN_IN), .A(n13314), .ZN(
        n13296) );
  OAI21_X1 U16640 ( .B1(n13429), .B2(n13297), .A(n13296), .ZN(P2_U2957) );
  INV_X1 U16641 ( .A(P2_UWORD_REG_4__SCAN_IN), .ZN(n13299) );
  OAI22_X1 U16642 ( .A1(n14070), .A2(BUF1_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n14069), .ZN(n13948) );
  NOR2_X1 U16643 ( .A1(n13359), .A2(n13948), .ZN(n13311) );
  AOI21_X1 U16644 ( .B1(n19081), .B2(P2_EAX_REG_20__SCAN_IN), .A(n13311), .ZN(
        n13298) );
  OAI21_X1 U16645 ( .B1(n13429), .B2(n13299), .A(n13298), .ZN(P2_U2956) );
  INV_X1 U16646 ( .A(P2_UWORD_REG_6__SCAN_IN), .ZN(n13301) );
  OAI22_X1 U16647 ( .A1(n14070), .A2(BUF1_REG_6__SCAN_IN), .B1(
        BUF2_REG_6__SCAN_IN), .B2(n14069), .ZN(n19140) );
  NOR2_X1 U16648 ( .A1(n13359), .A2(n19140), .ZN(n13317) );
  AOI21_X1 U16649 ( .B1(n19081), .B2(P2_EAX_REG_22__SCAN_IN), .A(n13317), .ZN(
        n13300) );
  OAI21_X1 U16650 ( .B1(n13429), .B2(n13301), .A(n13300), .ZN(P2_U2958) );
  INV_X1 U16651 ( .A(P2_LWORD_REG_1__SCAN_IN), .ZN(n13304) );
  AOI21_X1 U16652 ( .B1(P2_EAX_REG_1__SCAN_IN), .B2(n19081), .A(n13302), .ZN(
        n13303) );
  OAI21_X1 U16653 ( .B1(n13429), .B2(n13304), .A(n13303), .ZN(P2_U2968) );
  INV_X1 U16654 ( .A(P2_LWORD_REG_2__SCAN_IN), .ZN(n13307) );
  AOI21_X1 U16655 ( .B1(P2_EAX_REG_2__SCAN_IN), .B2(n19081), .A(n13305), .ZN(
        n13306) );
  OAI21_X1 U16656 ( .B1(n13429), .B2(n13307), .A(n13306), .ZN(P2_U2969) );
  INV_X1 U16657 ( .A(P2_LWORD_REG_3__SCAN_IN), .ZN(n13310) );
  AOI21_X1 U16658 ( .B1(P2_EAX_REG_3__SCAN_IN), .B2(n19081), .A(n13308), .ZN(
        n13309) );
  OAI21_X1 U16659 ( .B1(n13429), .B2(n13310), .A(n13309), .ZN(P2_U2970) );
  INV_X1 U16660 ( .A(P2_LWORD_REG_4__SCAN_IN), .ZN(n13313) );
  AOI21_X1 U16661 ( .B1(P2_EAX_REG_4__SCAN_IN), .B2(n19081), .A(n13311), .ZN(
        n13312) );
  OAI21_X1 U16662 ( .B1(n13429), .B2(n13313), .A(n13312), .ZN(P2_U2971) );
  INV_X1 U16663 ( .A(P2_LWORD_REG_5__SCAN_IN), .ZN(n13316) );
  AOI21_X1 U16664 ( .B1(P2_EAX_REG_5__SCAN_IN), .B2(n19081), .A(n13314), .ZN(
        n13315) );
  OAI21_X1 U16665 ( .B1(n13429), .B2(n13316), .A(n13315), .ZN(P2_U2972) );
  INV_X1 U16666 ( .A(P2_LWORD_REG_6__SCAN_IN), .ZN(n13319) );
  AOI21_X1 U16667 ( .B1(n19081), .B2(P2_EAX_REG_6__SCAN_IN), .A(n13317), .ZN(
        n13318) );
  OAI21_X1 U16668 ( .B1(n13429), .B2(n13319), .A(n13318), .ZN(P2_U2973) );
  INV_X1 U16669 ( .A(P2_LWORD_REG_7__SCAN_IN), .ZN(n13321) );
  AOI22_X1 U16670 ( .A1(n14069), .A2(BUF1_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n14070), .ZN(n19150) );
  NOR2_X1 U16671 ( .A1(n13359), .A2(n19150), .ZN(n13322) );
  AOI21_X1 U16672 ( .B1(n19081), .B2(P2_EAX_REG_7__SCAN_IN), .A(n13322), .ZN(
        n13320) );
  OAI21_X1 U16673 ( .B1(n13429), .B2(n13321), .A(n13320), .ZN(P2_U2974) );
  INV_X1 U16674 ( .A(P2_UWORD_REG_7__SCAN_IN), .ZN(n13324) );
  AOI21_X1 U16675 ( .B1(n19081), .B2(P2_EAX_REG_23__SCAN_IN), .A(n13322), .ZN(
        n13323) );
  OAI21_X1 U16676 ( .B1(n13429), .B2(n13324), .A(n13323), .ZN(P2_U2959) );
  INV_X1 U16677 ( .A(P2_LWORD_REG_11__SCAN_IN), .ZN(n13329) );
  INV_X1 U16678 ( .A(BUF1_REG_11__SCAN_IN), .ZN(n14125) );
  OR2_X1 U16679 ( .A1(n14070), .A2(n14125), .ZN(n13326) );
  NAND2_X1 U16680 ( .A1(n14070), .A2(BUF2_REG_11__SCAN_IN), .ZN(n13325) );
  AND2_X1 U16681 ( .A1(n13326), .A2(n13325), .ZN(n15039) );
  INV_X1 U16682 ( .A(n15039), .ZN(n13327) );
  NAND2_X1 U16683 ( .A1(n13448), .A2(n13327), .ZN(n13430) );
  NAND2_X1 U16684 ( .A1(n19081), .A2(P2_EAX_REG_11__SCAN_IN), .ZN(n13328) );
  OAI211_X1 U16685 ( .C1(n13429), .C2(n13329), .A(n13430), .B(n13328), .ZN(
        P2_U2978) );
  INV_X1 U16686 ( .A(P2_LWORD_REG_13__SCAN_IN), .ZN(n13331) );
  MUX2_X1 U16687 ( .A(BUF1_REG_13__SCAN_IN), .B(BUF2_REG_13__SCAN_IN), .S(
        n14070), .Z(n15019) );
  NAND2_X1 U16688 ( .A1(n13448), .A2(n15019), .ZN(n13434) );
  NAND2_X1 U16689 ( .A1(n19081), .A2(P2_EAX_REG_13__SCAN_IN), .ZN(n13330) );
  OAI211_X1 U16690 ( .C1(n13429), .C2(n13331), .A(n13434), .B(n13330), .ZN(
        P2_U2980) );
  INV_X1 U16691 ( .A(P2_LWORD_REG_12__SCAN_IN), .ZN(n13333) );
  MUX2_X1 U16692 ( .A(BUF1_REG_12__SCAN_IN), .B(BUF2_REG_12__SCAN_IN), .S(
        n14070), .Z(n15029) );
  NAND2_X1 U16693 ( .A1(n13448), .A2(n15029), .ZN(n13432) );
  NAND2_X1 U16694 ( .A1(n19081), .A2(P2_EAX_REG_12__SCAN_IN), .ZN(n13332) );
  OAI211_X1 U16695 ( .C1(n13429), .C2(n13333), .A(n13432), .B(n13332), .ZN(
        P2_U2979) );
  NAND2_X1 U16696 ( .A1(n13334), .A2(P2_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(
        n13335) );
  AND4_X1 U16697 ( .A1(n10427), .A2(n13335), .A3(P2_STATE2_REG_0__SCAN_IN), 
        .A4(n19798), .ZN(n13336) );
  MUX2_X1 U16698 ( .A(n13337), .B(n10284), .S(n14993), .Z(n13338) );
  OAI21_X1 U16699 ( .B1(n15009), .B2(n19818), .A(n13338), .ZN(P2_U2887) );
  INV_X1 U16700 ( .A(n15514), .ZN(n13354) );
  AND2_X1 U16701 ( .A1(n19085), .A2(P2_REIP_REG_0__SCAN_IN), .ZN(n13367) );
  INV_X1 U16702 ( .A(n13339), .ZN(n13342) );
  NAND2_X1 U16703 ( .A1(n13340), .A2(n20914), .ZN(n13341) );
  NAND2_X1 U16704 ( .A1(n13342), .A2(n13341), .ZN(n13365) );
  INV_X1 U16705 ( .A(n13343), .ZN(n13349) );
  INV_X1 U16706 ( .A(n13344), .ZN(n13347) );
  INV_X1 U16707 ( .A(n13345), .ZN(n13346) );
  NAND2_X1 U16708 ( .A1(n13347), .A2(n13346), .ZN(n13348) );
  NAND2_X1 U16709 ( .A1(n13349), .A2(n13348), .ZN(n18944) );
  OAI22_X1 U16710 ( .A1(n16223), .A2(n13365), .B1(n16222), .B2(n18944), .ZN(
        n13350) );
  AOI211_X1 U16711 ( .C1(n16219), .C2(n18950), .A(n13367), .B(n13350), .ZN(
        n13353) );
  OAI21_X1 U16712 ( .B1(n18943), .B2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13373), .ZN(n13351) );
  INV_X1 U16713 ( .A(n13351), .ZN(n13368) );
  AOI22_X1 U16714 ( .A1(n16227), .A2(n13368), .B1(n15511), .B2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n13352) );
  OAI211_X1 U16715 ( .C1(n13354), .C2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(
        n13353), .B(n13352), .ZN(P2_U3046) );
  INV_X1 U16716 ( .A(P2_LWORD_REG_15__SCAN_IN), .ZN(n13356) );
  AOI22_X1 U16717 ( .A1(n14069), .A2(BUF1_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n14070), .ZN(n13852) );
  INV_X1 U16718 ( .A(P2_EAX_REG_15__SCAN_IN), .ZN(n13355) );
  OAI222_X1 U16719 ( .A1(n13356), .A2(n13429), .B1(n13359), .B2(n13852), .C1(
        n13355), .C2(n13452), .ZN(P2_U2982) );
  INV_X1 U16720 ( .A(P2_UWORD_REG_0__SCAN_IN), .ZN(n13357) );
  INV_X1 U16721 ( .A(P2_EAX_REG_16__SCAN_IN), .ZN(n19047) );
  OAI22_X1 U16722 ( .A1(n14070), .A2(BUF1_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n14069), .ZN(n19115) );
  OAI222_X1 U16723 ( .A1(n13357), .A2(n13429), .B1(n13452), .B2(n19047), .C1(
        n19115), .C2(n13359), .ZN(P2_U2952) );
  INV_X1 U16724 ( .A(P2_LWORD_REG_0__SCAN_IN), .ZN(n13360) );
  INV_X1 U16725 ( .A(P2_EAX_REG_0__SCAN_IN), .ZN(n13358) );
  OAI222_X1 U16726 ( .A1(n13360), .A2(n13429), .B1(n13359), .B2(n19115), .C1(
        n13452), .C2(n13358), .ZN(P2_U2967) );
  INV_X1 U16727 ( .A(n13361), .ZN(n13363) );
  MUX2_X1 U16728 ( .A(n14929), .B(n15507), .S(n14993), .Z(n13364) );
  OAI21_X1 U16729 ( .B1(n19808), .B2(n15009), .A(n13364), .ZN(P2_U2886) );
  NOR2_X1 U16730 ( .A1(n19092), .A2(n13365), .ZN(n13366) );
  AOI211_X1 U16731 ( .C1(n19087), .C2(n13368), .A(n13367), .B(n13366), .ZN(
        n13371) );
  OAI21_X1 U16732 ( .B1(n19086), .B2(n13369), .A(
        P2_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n13370) );
  OAI211_X1 U16733 ( .C1(n16174), .C2(n10284), .A(n13371), .B(n13370), .ZN(
        P2_U3014) );
  OAI21_X1 U16734 ( .B1(n14930), .B2(n13373), .A(n13372), .ZN(n13374) );
  XOR2_X1 U16735 ( .A(n13374), .B(n15530), .Z(n15512) );
  AND2_X1 U16736 ( .A1(n19085), .A2(P2_REIP_REG_1__SCAN_IN), .ZN(n15509) );
  OAI21_X1 U16737 ( .B1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n13376), .A(
        n13375), .ZN(n15506) );
  NOR2_X1 U16738 ( .A1(n19092), .A2(n15506), .ZN(n13377) );
  AOI211_X1 U16739 ( .C1(n19087), .C2(n15512), .A(n15509), .B(n13377), .ZN(
        n13379) );
  MUX2_X1 U16740 ( .A(n19098), .B(n19113), .S(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .Z(n13378) );
  OAI211_X1 U16741 ( .C1(n15507), .C2(n16174), .A(n13379), .B(n13378), .ZN(
        P2_U3013) );
  NAND2_X1 U16742 ( .A1(n16257), .A2(n13592), .ZN(n13383) );
  NAND2_X1 U16743 ( .A1(n13381), .A2(n13380), .ZN(n13382) );
  NAND2_X1 U16744 ( .A1(n13383), .A2(n13382), .ZN(n13608) );
  NOR2_X1 U16745 ( .A1(n13384), .A2(n12635), .ZN(n13385) );
  NAND2_X1 U16746 ( .A1(n15083), .A2(n13388), .ZN(n15084) );
  AND2_X1 U16747 ( .A1(n9817), .A2(n10443), .ZN(n13389) );
  NAND2_X1 U16748 ( .A1(n15083), .A2(n13389), .ZN(n14071) );
  INV_X1 U16749 ( .A(n18944), .ZN(n13391) );
  NOR2_X1 U16750 ( .A1(n19818), .A2(n18944), .ZN(n19008) );
  INV_X1 U16751 ( .A(n19008), .ZN(n13390) );
  INV_X1 U16752 ( .A(n19009), .ZN(n16121) );
  OAI211_X1 U16753 ( .C1(n19158), .C2(n13391), .A(n13390), .B(n16121), .ZN(
        n13393) );
  AOI22_X1 U16754 ( .A1(n19005), .A2(n13391), .B1(n19004), .B2(
        P2_EAX_REG_0__SCAN_IN), .ZN(n13392) );
  OAI211_X1 U16755 ( .C1(n19013), .C2(n19115), .A(n13393), .B(n13392), .ZN(
        P2_U2919) );
  XNOR2_X1 U16756 ( .A(n13395), .B(n13394), .ZN(n13990) );
  INV_X1 U16757 ( .A(n13990), .ZN(n18923) );
  INV_X1 U16758 ( .A(n19005), .ZN(n18969) );
  INV_X1 U16759 ( .A(P2_EAX_REG_6__SCAN_IN), .ZN(n19067) );
  OAI222_X1 U16760 ( .A1(n18923), .A2(n18995), .B1(n15083), .B2(n19067), .C1(
        n19140), .C2(n19013), .ZN(P2_U2913) );
  AOI21_X1 U16761 ( .B1(n13398), .B2(n13397), .A(n13396), .ZN(n19799) );
  OAI21_X1 U16762 ( .B1(n13401), .B2(n13400), .A(n13399), .ZN(n19099) );
  NAND2_X1 U16763 ( .A1(n19085), .A2(P2_REIP_REG_2__SCAN_IN), .ZN(n19111) );
  OAI21_X1 U16764 ( .B1(n16223), .B2(n19099), .A(n19111), .ZN(n13407) );
  NAND2_X1 U16765 ( .A1(n13403), .A2(n13402), .ZN(n13404) );
  NAND2_X1 U16766 ( .A1(n13405), .A2(n13404), .ZN(n19109) );
  OAI22_X1 U16767 ( .A1(n16217), .A2(n19109), .B1(n13875), .B2(n13874), .ZN(
        n13406) );
  AOI211_X1 U16768 ( .C1(n19105), .C2(n16219), .A(n13407), .B(n13406), .ZN(
        n13415) );
  NOR2_X1 U16769 ( .A1(n15400), .A2(n15513), .ZN(n13412) );
  INV_X1 U16770 ( .A(n15511), .ZN(n13410) );
  OR2_X1 U16771 ( .A1(n15400), .A2(n13408), .ZN(n13409) );
  OAI211_X1 U16772 ( .C1(n15513), .C2(n13875), .A(n13410), .B(n13409), .ZN(
        n13411) );
  MUX2_X1 U16773 ( .A(n13412), .B(n13411), .S(
        P2_INSTADDRPOINTER_REG_2__SCAN_IN), .Z(n13413) );
  INV_X1 U16774 ( .A(n13413), .ZN(n13414) );
  OAI211_X1 U16775 ( .C1(n19799), .C2(n16222), .A(n13415), .B(n13414), .ZN(
        P2_U3044) );
  AOI22_X1 U16776 ( .A1(P1_EAX_REG_3__SCAN_IN), .A2(n13569), .B1(n20026), .B2(
        P1_LWORD_REG_3__SCAN_IN), .ZN(n13419) );
  INV_X1 U16777 ( .A(DATAI_3_), .ZN(n13418) );
  NAND2_X1 U16778 ( .A1(n14173), .A2(BUF1_REG_3__SCAN_IN), .ZN(n13417) );
  OAI21_X1 U16779 ( .B1(n14173), .B2(n13418), .A(n13417), .ZN(n20130) );
  NAND2_X1 U16780 ( .A1(n13555), .A2(n20130), .ZN(n13547) );
  NAND2_X1 U16781 ( .A1(n13419), .A2(n13547), .ZN(P1_U2955) );
  AOI22_X1 U16782 ( .A1(P1_EAX_REG_6__SCAN_IN), .A2(n13569), .B1(n20026), .B2(
        P1_LWORD_REG_6__SCAN_IN), .ZN(n13422) );
  INV_X1 U16783 ( .A(DATAI_6_), .ZN(n13421) );
  NAND2_X1 U16784 ( .A1(n14173), .A2(BUF1_REG_6__SCAN_IN), .ZN(n13420) );
  OAI21_X1 U16785 ( .B1(n14173), .B2(n13421), .A(n13420), .ZN(n20139) );
  NAND2_X1 U16786 ( .A1(n13555), .A2(n20139), .ZN(n13570) );
  NAND2_X1 U16787 ( .A1(n13422), .A2(n13570), .ZN(P1_U2958) );
  AOI22_X1 U16788 ( .A1(P1_EAX_REG_5__SCAN_IN), .A2(n13569), .B1(n20026), .B2(
        P1_LWORD_REG_5__SCAN_IN), .ZN(n13425) );
  INV_X1 U16789 ( .A(DATAI_5_), .ZN(n13424) );
  NAND2_X1 U16790 ( .A1(n14173), .A2(BUF1_REG_5__SCAN_IN), .ZN(n13423) );
  OAI21_X1 U16791 ( .B1(n14173), .B2(n13424), .A(n13423), .ZN(n20136) );
  NAND2_X1 U16792 ( .A1(n13555), .A2(n20136), .ZN(n13563) );
  NAND2_X1 U16793 ( .A1(n13425), .A2(n13563), .ZN(P1_U2957) );
  AOI22_X1 U16794 ( .A1(P1_EAX_REG_4__SCAN_IN), .A2(n13569), .B1(n20026), .B2(
        P1_LWORD_REG_4__SCAN_IN), .ZN(n13428) );
  INV_X1 U16795 ( .A(DATAI_4_), .ZN(n13427) );
  NAND2_X1 U16796 ( .A1(n14173), .A2(BUF1_REG_4__SCAN_IN), .ZN(n13426) );
  OAI21_X1 U16797 ( .B1(n14173), .B2(n13427), .A(n13426), .ZN(n20133) );
  NAND2_X1 U16798 ( .A1(n13555), .A2(n20133), .ZN(n13559) );
  NAND2_X1 U16799 ( .A1(n13428), .A2(n13559), .ZN(P1_U2956) );
  INV_X1 U16800 ( .A(P2_EAX_REG_27__SCAN_IN), .ZN(n19025) );
  NAND2_X1 U16801 ( .A1(n19082), .A2(P2_UWORD_REG_11__SCAN_IN), .ZN(n13431) );
  OAI211_X1 U16802 ( .C1(n13452), .C2(n19025), .A(n13431), .B(n13430), .ZN(
        P2_U2963) );
  INV_X1 U16803 ( .A(P2_EAX_REG_28__SCAN_IN), .ZN(n19023) );
  NAND2_X1 U16804 ( .A1(n19082), .A2(P2_UWORD_REG_12__SCAN_IN), .ZN(n13433) );
  OAI211_X1 U16805 ( .C1(n13452), .C2(n19023), .A(n13433), .B(n13432), .ZN(
        P2_U2964) );
  INV_X1 U16806 ( .A(P2_EAX_REG_29__SCAN_IN), .ZN(n19021) );
  NAND2_X1 U16807 ( .A1(n19082), .A2(P2_UWORD_REG_13__SCAN_IN), .ZN(n13435) );
  OAI211_X1 U16808 ( .C1(n13452), .C2(n19021), .A(n13435), .B(n13434), .ZN(
        P2_U2965) );
  INV_X1 U16809 ( .A(P2_EAX_REG_9__SCAN_IN), .ZN(n19061) );
  NAND2_X1 U16810 ( .A1(n19082), .A2(P2_LWORD_REG_9__SCAN_IN), .ZN(n13438) );
  INV_X1 U16811 ( .A(BUF1_REG_9__SCAN_IN), .ZN(n16388) );
  OR2_X1 U16812 ( .A1(n14070), .A2(n16388), .ZN(n13437) );
  NAND2_X1 U16813 ( .A1(n14070), .A2(BUF2_REG_9__SCAN_IN), .ZN(n13436) );
  AND2_X1 U16814 ( .A1(n13437), .A2(n13436), .ZN(n15054) );
  INV_X1 U16815 ( .A(n15054), .ZN(n18982) );
  NAND2_X1 U16816 ( .A1(n13448), .A2(n18982), .ZN(n13450) );
  OAI211_X1 U16817 ( .C1(n19061), .C2(n13452), .A(n13438), .B(n13450), .ZN(
        P2_U2976) );
  INV_X1 U16818 ( .A(P2_EAX_REG_24__SCAN_IN), .ZN(n19031) );
  NAND2_X1 U16819 ( .A1(n19082), .A2(P2_UWORD_REG_8__SCAN_IN), .ZN(n13439) );
  MUX2_X1 U16820 ( .A(BUF1_REG_8__SCAN_IN), .B(BUF2_REG_8__SCAN_IN), .S(n14070), .Z(n18985) );
  NAND2_X1 U16821 ( .A1(n13448), .A2(n18985), .ZN(n13440) );
  OAI211_X1 U16822 ( .C1(n19031), .C2(n13452), .A(n13439), .B(n13440), .ZN(
        P2_U2960) );
  INV_X1 U16823 ( .A(P2_EAX_REG_8__SCAN_IN), .ZN(n19063) );
  NAND2_X1 U16824 ( .A1(n19082), .A2(P2_LWORD_REG_8__SCAN_IN), .ZN(n13441) );
  OAI211_X1 U16825 ( .C1(n19063), .C2(n13452), .A(n13441), .B(n13440), .ZN(
        P2_U2975) );
  INV_X1 U16826 ( .A(P2_EAX_REG_30__SCAN_IN), .ZN(n19019) );
  NAND2_X1 U16827 ( .A1(n19082), .A2(P2_UWORD_REG_14__SCAN_IN), .ZN(n13445) );
  INV_X1 U16828 ( .A(BUF1_REG_14__SCAN_IN), .ZN(n13442) );
  OR2_X1 U16829 ( .A1(n14070), .A2(n13442), .ZN(n13444) );
  NAND2_X1 U16830 ( .A1(n14070), .A2(BUF2_REG_14__SCAN_IN), .ZN(n13443) );
  AND2_X1 U16831 ( .A1(n13444), .A2(n13443), .ZN(n15012) );
  INV_X1 U16832 ( .A(n15012), .ZN(n18976) );
  NAND2_X1 U16833 ( .A1(n13448), .A2(n18976), .ZN(n19083) );
  OAI211_X1 U16834 ( .C1(n19019), .C2(n13452), .A(n13445), .B(n19083), .ZN(
        P2_U2966) );
  INV_X1 U16835 ( .A(P2_EAX_REG_26__SCAN_IN), .ZN(n19027) );
  NAND2_X1 U16836 ( .A1(n19082), .A2(P2_UWORD_REG_10__SCAN_IN), .ZN(n13449) );
  INV_X1 U16837 ( .A(BUF1_REG_10__SCAN_IN), .ZN(n14062) );
  OR2_X1 U16838 ( .A1(n14070), .A2(n14062), .ZN(n13447) );
  NAND2_X1 U16839 ( .A1(n14070), .A2(BUF2_REG_10__SCAN_IN), .ZN(n13446) );
  AND2_X1 U16840 ( .A1(n13447), .A2(n13446), .ZN(n15048) );
  INV_X1 U16841 ( .A(n15048), .ZN(n18979) );
  NAND2_X1 U16842 ( .A1(n13448), .A2(n18979), .ZN(n19079) );
  OAI211_X1 U16843 ( .C1(n19027), .C2(n13452), .A(n13449), .B(n19079), .ZN(
        P2_U2962) );
  INV_X1 U16844 ( .A(P2_EAX_REG_25__SCAN_IN), .ZN(n19029) );
  NAND2_X1 U16845 ( .A1(n19082), .A2(P2_UWORD_REG_9__SCAN_IN), .ZN(n13451) );
  OAI211_X1 U16846 ( .C1(n13452), .C2(n19029), .A(n13451), .B(n13450), .ZN(
        P2_U2961) );
  NOR3_X1 U16847 ( .A1(n14280), .A2(n13687), .A3(n13673), .ZN(n13462) );
  AND2_X1 U16848 ( .A1(n11487), .A2(n13454), .ZN(n13455) );
  AND3_X1 U16849 ( .A1(n13457), .A2(n13456), .A3(n13455), .ZN(n13458) );
  NAND2_X1 U16850 ( .A1(n13453), .A2(n13458), .ZN(n13460) );
  NOR2_X1 U16851 ( .A1(n13460), .A2(n13459), .ZN(n14281) );
  NOR2_X1 U16852 ( .A1(n20380), .A2(n14281), .ZN(n13461) );
  AOI211_X1 U16853 ( .C1(n15697), .C2(n13661), .A(n13462), .B(n13461), .ZN(
        n15700) );
  INV_X1 U16854 ( .A(n15700), .ZN(n13465) );
  NAND2_X1 U16855 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n14862) );
  OAI22_X1 U16856 ( .A1(n12524), .A2(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B1(
        n20087), .B2(P1_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n14860) );
  NOR2_X1 U16857 ( .A1(n14862), .A2(n14860), .ZN(n13464) );
  NAND2_X1 U16858 ( .A1(P1_STATE2_REG_3__SCAN_IN), .A2(n13698), .ZN(n20758) );
  NOR3_X1 U16859 ( .A1(n13687), .A2(n13673), .A3(n20758), .ZN(n13463) );
  AOI211_X1 U16860 ( .C1(n13465), .C2(n14858), .A(n13464), .B(n13463), .ZN(
        n13479) );
  OAI21_X1 U16861 ( .B1(n13466), .B2(n20791), .A(n13657), .ZN(n13467) );
  NAND2_X1 U16862 ( .A1(n13698), .A2(n13467), .ZN(n13484) );
  NOR2_X1 U16863 ( .A1(n15736), .A2(n20791), .ZN(n13468) );
  NAND2_X1 U16864 ( .A1(n13698), .A2(n13468), .ZN(n15693) );
  NAND2_X1 U16865 ( .A1(n13484), .A2(n15693), .ZN(n13470) );
  INV_X1 U16866 ( .A(n15697), .ZN(n13680) );
  NAND3_X1 U16867 ( .A1(n13680), .A2(n11487), .A3(n13657), .ZN(n13469) );
  NAND2_X1 U16868 ( .A1(n13470), .A2(n13469), .ZN(n13477) );
  NOR2_X1 U16869 ( .A1(n13453), .A2(n20791), .ZN(n13471) );
  NAND2_X1 U16870 ( .A1(n13472), .A2(n13471), .ZN(n13482) );
  OAI211_X1 U16871 ( .C1(n14432), .C2(n11108), .A(n13482), .B(n13473), .ZN(
        n13474) );
  INV_X1 U16872 ( .A(n13474), .ZN(n13476) );
  INV_X1 U16873 ( .A(n13698), .ZN(n13475) );
  NAND2_X1 U16874 ( .A1(n13475), .A2(n13658), .ZN(n13519) );
  NAND2_X1 U16875 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .ZN(n15997) );
  INV_X1 U16876 ( .A(n15997), .ZN(n13727) );
  NAND2_X1 U16877 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(n13727), .ZN(n16001) );
  INV_X1 U16878 ( .A(P1_FLUSH_REG_SCAN_IN), .ZN(n19864) );
  OAI22_X1 U16879 ( .A1(n15699), .A2(n19857), .B1(n16001), .B2(n19864), .ZN(
        n13497) );
  AOI21_X1 U16880 ( .B1(P1_STATE2_REG_3__SCAN_IN), .B2(n11192), .A(n13497), 
        .ZN(n14865) );
  NAND2_X1 U16881 ( .A1(P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(n14865), .ZN(
        n13478) );
  OAI21_X1 U16882 ( .B1(n13479), .B2(n14865), .A(n13478), .ZN(P1_U3473) );
  NAND4_X1 U16883 ( .A1(n13656), .A2(n14503), .A3(n13480), .A4(n11120), .ZN(
        n13517) );
  OR2_X1 U16884 ( .A1(n13517), .A2(n14427), .ZN(n13481) );
  NAND2_X1 U16885 ( .A1(n13484), .A2(n13483), .ZN(n13485) );
  NAND2_X1 U16886 ( .A1(n13486), .A2(n20145), .ZN(n13492) );
  INV_X1 U16887 ( .A(n13487), .ZN(n13491) );
  INV_X1 U16888 ( .A(n13488), .ZN(n13490) );
  OAI21_X1 U16889 ( .B1(n13491), .B2(n13490), .A(n13489), .ZN(n20049) );
  INV_X1 U16890 ( .A(P1_EAX_REG_0__SCAN_IN), .ZN(n19996) );
  INV_X1 U16891 ( .A(DATAI_0_), .ZN(n13494) );
  NAND2_X1 U16892 ( .A1(n14173), .A2(BUF1_REG_0__SCAN_IN), .ZN(n13493) );
  OAI21_X1 U16893 ( .B1(n14173), .B2(n13494), .A(n13493), .ZN(n20112) );
  INV_X1 U16894 ( .A(n20112), .ZN(n13495) );
  OAI222_X1 U16895 ( .A1(n14566), .A2(n20049), .B1(n14529), .B2(n19996), .C1(
        n14155), .C2(n13495), .ZN(P1_U2904) );
  INV_X1 U16896 ( .A(n14865), .ZN(n20761) );
  INV_X1 U16897 ( .A(n13453), .ZN(n13689) );
  INV_X1 U16898 ( .A(n20257), .ZN(n20512) );
  OR2_X1 U16899 ( .A1(n11270), .A2(n20512), .ZN(n13496) );
  XNOR2_X1 U16900 ( .A(n13496), .B(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(
        n19922) );
  NAND4_X1 U16901 ( .A1(n13497), .A2(n14858), .A3(n13689), .A4(n19922), .ZN(
        n13498) );
  OAI21_X1 U16902 ( .B1(n13690), .B2(n20761), .A(n13498), .ZN(P1_U3468) );
  OAI21_X1 U16903 ( .B1(n13500), .B2(n13499), .A(n14048), .ZN(n18911) );
  OAI222_X1 U16904 ( .A1(n18911), .A2(n18995), .B1(n19150), .B2(n19013), .C1(
        n19065), .C2(n15083), .ZN(P2_U2912) );
  INV_X1 U16905 ( .A(n13501), .ZN(n13502) );
  INV_X1 U16906 ( .A(n19804), .ZN(n13834) );
  MUX2_X1 U16907 ( .A(n21020), .B(n14914), .S(n14993), .Z(n13504) );
  OAI21_X1 U16908 ( .B1(n13834), .B2(n15009), .A(n13504), .ZN(P2_U2885) );
  NAND2_X1 U16909 ( .A1(n12867), .A2(n13505), .ZN(n13581) );
  NAND2_X1 U16910 ( .A1(n13506), .A2(n13581), .ZN(n13507) );
  NAND2_X1 U16911 ( .A1(n13508), .A2(n13507), .ZN(n13509) );
  NOR2_X1 U16912 ( .A1(n14993), .A2(n10656), .ZN(n13510) );
  OAI21_X1 U16913 ( .B1(n19788), .B2(n15009), .A(n13511), .ZN(P2_U2884) );
  INV_X1 U16914 ( .A(P1_EAX_REG_30__SCAN_IN), .ZN(n20018) );
  NAND2_X1 U16915 ( .A1(n13621), .A2(n15697), .ZN(n13512) );
  NAND2_X1 U16916 ( .A1(n20035), .A2(n13512), .ZN(n13514) );
  NAND2_X1 U16917 ( .A1(n19969), .A2(n11501), .ZN(n13772) );
  NAND2_X1 U16918 ( .A1(n11192), .A2(n13727), .ZN(n20790) );
  INV_X2 U16919 ( .A(n20790), .ZN(n19993) );
  NOR2_X4 U16920 ( .A1(n19969), .A2(n19993), .ZN(n19978) );
  AOI22_X1 U16921 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n19978), .B1(n19993), 
        .B2(P1_UWORD_REG_14__SCAN_IN), .ZN(n13515) );
  OAI21_X1 U16922 ( .B1(n20018), .B2(n13772), .A(n13515), .ZN(P1_U2906) );
  OR2_X1 U16923 ( .A1(n13517), .A2(n13516), .ZN(n13518) );
  NAND2_X1 U16924 ( .A1(n13519), .A2(n13518), .ZN(n13521) );
  NAND2_X2 U16925 ( .A1(n19968), .A2(n20145), .ZN(n14496) );
  NAND2_X1 U16926 ( .A1(n13522), .A2(n10100), .ZN(n13525) );
  INV_X1 U16927 ( .A(n13523), .ZN(n13524) );
  AND2_X1 U16928 ( .A1(n13525), .A2(n13524), .ZN(n20088) );
  INV_X1 U16929 ( .A(n20088), .ZN(n13526) );
  OAI222_X1 U16930 ( .A1(n20049), .A2(n14496), .B1(n11502), .B2(n19968), .C1(
        n13526), .C2(n19962), .ZN(P1_U2872) );
  XOR2_X1 U16931 ( .A(P2_INSTQUEUE_REG_0__7__SCAN_IN), .B(n13637), .Z(n13532)
         );
  NAND2_X1 U16932 ( .A1(n13527), .A2(n13641), .ZN(n13530) );
  INV_X1 U16933 ( .A(n13528), .ZN(n13529) );
  NAND2_X1 U16934 ( .A1(n13530), .A2(n13529), .ZN(n18910) );
  MUX2_X1 U16935 ( .A(n10719), .B(n18910), .S(n14993), .Z(n13531) );
  OAI21_X1 U16936 ( .B1(n13532), .B2(n15009), .A(n13531), .ZN(P2_U2880) );
  INV_X1 U16937 ( .A(P1_EAX_REG_27__SCAN_IN), .ZN(n20007) );
  AOI22_X1 U16938 ( .A1(n19993), .A2(P1_UWORD_REG_11__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_27__SCAN_IN), .ZN(n13533) );
  OAI21_X1 U16939 ( .B1(n20007), .B2(n13772), .A(n13533), .ZN(P1_U2909) );
  INV_X1 U16940 ( .A(P1_EAX_REG_25__SCAN_IN), .ZN(n20002) );
  AOI22_X1 U16941 ( .A1(n19993), .A2(P1_UWORD_REG_9__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_25__SCAN_IN), .ZN(n13534) );
  OAI21_X1 U16942 ( .B1(n20002), .B2(n13772), .A(n13534), .ZN(P1_U2911) );
  INV_X1 U16943 ( .A(P1_EAX_REG_24__SCAN_IN), .ZN(n19999) );
  AOI22_X1 U16944 ( .A1(n19993), .A2(P1_UWORD_REG_8__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_24__SCAN_IN), .ZN(n13535) );
  OAI21_X1 U16945 ( .B1(n19999), .B2(n13772), .A(n13535), .ZN(P1_U2912) );
  AOI22_X1 U16946 ( .A1(n19993), .A2(P1_UWORD_REG_12__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_28__SCAN_IN), .ZN(n13536) );
  OAI21_X1 U16947 ( .B1(n14512), .B2(n13772), .A(n13536), .ZN(P1_U2908) );
  INV_X1 U16948 ( .A(P1_EAX_REG_23__SCAN_IN), .ZN(n13538) );
  AOI22_X1 U16949 ( .A1(n19993), .A2(P1_UWORD_REG_7__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_23__SCAN_IN), .ZN(n13537) );
  OAI21_X1 U16950 ( .B1(n13538), .B2(n13772), .A(n13537), .ZN(P1_U2913) );
  OR2_X1 U16951 ( .A1(n13540), .A2(n13539), .ZN(n13541) );
  NAND2_X1 U16952 ( .A1(n13646), .A2(n13541), .ZN(n14445) );
  XNOR2_X1 U16953 ( .A(n13542), .B(n11588), .ZN(n20080) );
  INV_X1 U16954 ( .A(n19968), .ZN(n14492) );
  AOI22_X1 U16955 ( .A1(n15856), .A2(n20080), .B1(P1_EBX_REG_1__SCAN_IN), .B2(
        n14492), .ZN(n13543) );
  OAI21_X1 U16956 ( .B1(n14445), .B2(n14496), .A(n13543), .ZN(P1_U2871) );
  AOI22_X1 U16957 ( .A1(P1_EAX_REG_18__SCAN_IN), .A2(n13569), .B1(n20026), 
        .B2(P1_UWORD_REG_2__SCAN_IN), .ZN(n13546) );
  INV_X1 U16958 ( .A(DATAI_2_), .ZN(n13545) );
  NAND2_X1 U16959 ( .A1(n14173), .A2(BUF1_REG_2__SCAN_IN), .ZN(n13544) );
  OAI21_X1 U16960 ( .B1(n14173), .B2(n13545), .A(n13544), .ZN(n20126) );
  NAND2_X1 U16961 ( .A1(n13555), .A2(n20126), .ZN(n13557) );
  NAND2_X1 U16962 ( .A1(n13546), .A2(n13557), .ZN(P1_U2939) );
  AOI22_X1 U16963 ( .A1(P1_EAX_REG_19__SCAN_IN), .A2(n13569), .B1(n20026), 
        .B2(P1_UWORD_REG_3__SCAN_IN), .ZN(n13548) );
  NAND2_X1 U16964 ( .A1(n13548), .A2(n13547), .ZN(P1_U2940) );
  AOI22_X1 U16965 ( .A1(P1_EAX_REG_1__SCAN_IN), .A2(n13569), .B1(n20026), .B2(
        P1_LWORD_REG_1__SCAN_IN), .ZN(n13551) );
  INV_X1 U16966 ( .A(DATAI_1_), .ZN(n13550) );
  NAND2_X1 U16967 ( .A1(n14173), .A2(BUF1_REG_1__SCAN_IN), .ZN(n13549) );
  OAI21_X1 U16968 ( .B1(n14173), .B2(n13550), .A(n13549), .ZN(n20123) );
  NAND2_X1 U16969 ( .A1(n13555), .A2(n20123), .ZN(n13567) );
  NAND2_X1 U16970 ( .A1(n13551), .A2(n13567), .ZN(P1_U2953) );
  AOI22_X1 U16971 ( .A1(P1_EAX_REG_0__SCAN_IN), .A2(n13569), .B1(n20026), .B2(
        P1_LWORD_REG_0__SCAN_IN), .ZN(n13552) );
  NAND2_X1 U16972 ( .A1(n13555), .A2(n20112), .ZN(n13565) );
  NAND2_X1 U16973 ( .A1(n13552), .A2(n13565), .ZN(P1_U2952) );
  AOI22_X1 U16974 ( .A1(P1_EAX_REG_7__SCAN_IN), .A2(n13569), .B1(n20026), .B2(
        P1_LWORD_REG_7__SCAN_IN), .ZN(n13556) );
  INV_X1 U16975 ( .A(DATAI_7_), .ZN(n13554) );
  NAND2_X1 U16976 ( .A1(n14173), .A2(BUF1_REG_7__SCAN_IN), .ZN(n13553) );
  OAI21_X1 U16977 ( .B1(n14173), .B2(n13554), .A(n13553), .ZN(n20148) );
  NAND2_X1 U16978 ( .A1(n13555), .A2(n20148), .ZN(n13561) );
  NAND2_X1 U16979 ( .A1(n13556), .A2(n13561), .ZN(P1_U2959) );
  AOI22_X1 U16980 ( .A1(P1_EAX_REG_2__SCAN_IN), .A2(n13569), .B1(n20026), .B2(
        P1_LWORD_REG_2__SCAN_IN), .ZN(n13558) );
  NAND2_X1 U16981 ( .A1(n13558), .A2(n13557), .ZN(P1_U2954) );
  AOI22_X1 U16982 ( .A1(P1_EAX_REG_20__SCAN_IN), .A2(n13569), .B1(n20026), 
        .B2(P1_UWORD_REG_4__SCAN_IN), .ZN(n13560) );
  NAND2_X1 U16983 ( .A1(n13560), .A2(n13559), .ZN(P1_U2941) );
  AOI22_X1 U16984 ( .A1(P1_EAX_REG_23__SCAN_IN), .A2(n13569), .B1(n20026), 
        .B2(P1_UWORD_REG_7__SCAN_IN), .ZN(n13562) );
  NAND2_X1 U16985 ( .A1(n13562), .A2(n13561), .ZN(P1_U2944) );
  AOI22_X1 U16986 ( .A1(P1_EAX_REG_21__SCAN_IN), .A2(n13569), .B1(n20026), 
        .B2(P1_UWORD_REG_5__SCAN_IN), .ZN(n13564) );
  NAND2_X1 U16987 ( .A1(n13564), .A2(n13563), .ZN(P1_U2942) );
  AOI22_X1 U16988 ( .A1(P1_EAX_REG_16__SCAN_IN), .A2(n13569), .B1(n20026), 
        .B2(P1_UWORD_REG_0__SCAN_IN), .ZN(n13566) );
  NAND2_X1 U16989 ( .A1(n13566), .A2(n13565), .ZN(P1_U2937) );
  AOI22_X1 U16990 ( .A1(P1_EAX_REG_17__SCAN_IN), .A2(n13569), .B1(n20026), 
        .B2(P1_UWORD_REG_1__SCAN_IN), .ZN(n13568) );
  NAND2_X1 U16991 ( .A1(n13568), .A2(n13567), .ZN(P1_U2938) );
  AOI22_X1 U16992 ( .A1(P1_EAX_REG_22__SCAN_IN), .A2(n13569), .B1(n20026), 
        .B2(P1_UWORD_REG_6__SCAN_IN), .ZN(n13571) );
  NAND2_X1 U16993 ( .A1(n13571), .A2(n13570), .ZN(P1_U2943) );
  NOR2_X1 U16994 ( .A1(n13572), .A2(n13528), .ZN(n13573) );
  OR2_X1 U16995 ( .A1(n13705), .A2(n13573), .ZN(n16211) );
  OAI211_X1 U16996 ( .C1(n13576), .C2(n13575), .A(n13574), .B(n14965), .ZN(
        n13578) );
  NAND2_X1 U16997 ( .A1(n15006), .A2(P2_EBX_REG_8__SCAN_IN), .ZN(n13577) );
  OAI211_X1 U16998 ( .C1(n16211), .C2(n15006), .A(n13578), .B(n13577), .ZN(
        P2_U2879) );
  INV_X1 U16999 ( .A(P1_EAX_REG_1__SCAN_IN), .ZN(n19992) );
  INV_X1 U17000 ( .A(n20123), .ZN(n13579) );
  OAI222_X1 U17001 ( .A1(n14566), .A2(n14445), .B1(n14529), .B2(n19992), .C1(
        n14155), .C2(n13579), .ZN(P1_U2903) );
  NAND2_X1 U17002 ( .A1(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n9817), .ZN(
        n13580) );
  AND2_X1 U17003 ( .A1(n13581), .A2(n13580), .ZN(n13582) );
  NAND2_X1 U17004 ( .A1(n13583), .A2(n13582), .ZN(n13586) );
  INV_X1 U17005 ( .A(P2_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n13951) );
  NOR2_X1 U17006 ( .A1(n13584), .A2(n13951), .ZN(n13585) );
  NAND2_X1 U17007 ( .A1(n13586), .A2(n13585), .ZN(n13636) );
  OAI21_X1 U17008 ( .B1(n13586), .B2(n13585), .A(n13636), .ZN(n18990) );
  OR2_X1 U17009 ( .A1(n13588), .A2(n13587), .ZN(n13589) );
  AND2_X1 U17010 ( .A1(n13589), .A2(n13629), .ZN(n19089) );
  INV_X1 U17011 ( .A(n19089), .ZN(n13878) );
  MUX2_X1 U17012 ( .A(n13878), .B(n14033), .S(n15006), .Z(n13590) );
  OAI21_X1 U17013 ( .B1(n18990), .B2(n15009), .A(n13590), .ZN(P2_U2883) );
  INV_X1 U17014 ( .A(n16286), .ZN(n15551) );
  INV_X1 U17015 ( .A(n13591), .ZN(n16256) );
  OR2_X1 U17016 ( .A1(n16256), .A2(n13592), .ZN(n15544) );
  NAND2_X1 U17017 ( .A1(n15544), .A2(n16232), .ZN(n13596) );
  INV_X1 U17018 ( .A(n13593), .ZN(n13595) );
  INV_X1 U17019 ( .A(n13594), .ZN(n15535) );
  NAND2_X1 U17020 ( .A1(n15535), .A2(n15554), .ZN(n15539) );
  INV_X1 U17021 ( .A(n15539), .ZN(n13598) );
  AOI21_X1 U17022 ( .B1(n13596), .B2(n13595), .A(n13598), .ZN(n13605) );
  AND2_X1 U17023 ( .A1(n10472), .A2(n13597), .ZN(n15548) );
  INV_X1 U17024 ( .A(n10546), .ZN(n13599) );
  AOI21_X1 U17025 ( .B1(n12628), .B2(n13599), .A(n13598), .ZN(n13600) );
  OAI21_X1 U17026 ( .B1(n15548), .B2(n13601), .A(n13600), .ZN(n13603) );
  AND2_X1 U17027 ( .A1(n12628), .A2(n10546), .ZN(n13602) );
  MUX2_X1 U17028 ( .A(n13603), .B(n13602), .S(n16232), .Z(n13604) );
  NOR2_X1 U17029 ( .A1(n13605), .A2(n13604), .ZN(n13606) );
  NAND2_X1 U17030 ( .A1(n13607), .A2(n13606), .ZN(n16245) );
  AOI22_X1 U17031 ( .A1(n19407), .A2(n15551), .B1(n15552), .B2(n16245), .ZN(
        n13619) );
  NAND2_X1 U17032 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(
        P2_STATE2_REG_1__SCAN_IN), .ZN(n19815) );
  INV_X1 U17033 ( .A(n19815), .ZN(n13938) );
  NAND2_X1 U17034 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n13938), .ZN(n16295) );
  INV_X1 U17035 ( .A(n16295), .ZN(n16277) );
  INV_X1 U17036 ( .A(n13608), .ZN(n13616) );
  AND2_X1 U17037 ( .A1(n13610), .A2(n13609), .ZN(n13615) );
  INV_X1 U17038 ( .A(n13611), .ZN(n13612) );
  OR2_X1 U17039 ( .A1(n12599), .A2(n13612), .ZN(n13613) );
  OR2_X1 U17040 ( .A1(n19015), .A2(n13613), .ZN(n13614) );
  OAI22_X1 U17041 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19798), .B1(n16268), 
        .B2(n16292), .ZN(n13617) );
  AOI21_X1 U17042 ( .B1(P2_FLUSH_REG_SCAN_IN), .B2(n16277), .A(n13617), .ZN(
        n15662) );
  NAND2_X1 U17043 ( .A1(n15662), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13618) );
  OAI21_X1 U17044 ( .B1(n13619), .B2(n15662), .A(n13618), .ZN(P2_U3596) );
  NAND2_X1 U17045 ( .A1(P1_STATEBS16_REG_SCAN_IN), .A2(n15725), .ZN(n15995) );
  INV_X1 U17046 ( .A(n15995), .ZN(n13620) );
  INV_X1 U17047 ( .A(n20101), .ZN(n20048) );
  NAND2_X1 U17048 ( .A1(n20767), .A2(n13622), .ZN(n20787) );
  NAND2_X1 U17049 ( .A1(n20787), .A2(n11192), .ZN(n13623) );
  INV_X1 U17050 ( .A(P1_REIP_REG_1__SCAN_IN), .ZN(n20776) );
  NOR2_X1 U17051 ( .A1(n20046), .A2(n20776), .ZN(n20079) );
  NAND2_X1 U17052 ( .A1(n11192), .A2(P1_STATE2_REG_2__SCAN_IN), .ZN(n15695) );
  NAND2_X1 U17053 ( .A1(n20765), .A2(P1_STATE2_REG_1__SCAN_IN), .ZN(n13624) );
  NAND2_X1 U17054 ( .A1(n15695), .A2(n13624), .ZN(n20037) );
  NOR2_X1 U17055 ( .A1(n15909), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(
        n13625) );
  AOI211_X1 U17056 ( .C1(n20038), .C2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .A(
        n20079), .B(n13625), .ZN(n13628) );
  XNOR2_X1 U17057 ( .A(n13626), .B(n20087), .ZN(n20078) );
  NAND2_X1 U17058 ( .A1(n20078), .A2(n20043), .ZN(n13627) );
  OAI211_X1 U17059 ( .C1(n20048), .C2(n14445), .A(n13628), .B(n13627), .ZN(
        P1_U2998) );
  XOR2_X1 U17060 ( .A(P2_INSTQUEUE_REG_0__5__SCAN_IN), .B(n13636), .Z(n13635)
         );
  INV_X1 U17061 ( .A(P2_EBX_REG_5__SCAN_IN), .ZN(n13633) );
  NAND2_X1 U17062 ( .A1(n13630), .A2(n13629), .ZN(n13632) );
  INV_X1 U17063 ( .A(n13639), .ZN(n13631) );
  AND2_X1 U17064 ( .A1(n13632), .A2(n13631), .ZN(n16188) );
  INV_X1 U17065 ( .A(n16188), .ZN(n18936) );
  MUX2_X1 U17066 ( .A(n13633), .B(n18936), .S(n14993), .Z(n13634) );
  OAI21_X1 U17067 ( .B1(n13635), .B2(n15009), .A(n13634), .ZN(P2_U2882) );
  NOR2_X1 U17068 ( .A1(n13636), .A2(n19138), .ZN(n13638) );
  OAI211_X1 U17069 ( .C1(n13638), .C2(P2_INSTQUEUE_REG_0__6__SCAN_IN), .A(
        n14965), .B(n13637), .ZN(n13644) );
  OR2_X1 U17070 ( .A1(n13640), .A2(n13639), .ZN(n13642) );
  AND2_X1 U17071 ( .A1(n13642), .A2(n13641), .ZN(n16180) );
  NAND2_X1 U17072 ( .A1(n14993), .A2(n16180), .ZN(n13643) );
  OAI211_X1 U17073 ( .C1(n14993), .C2(n13645), .A(n13644), .B(n13643), .ZN(
        P2_U2881) );
  NAND2_X1 U17074 ( .A1(n13647), .A2(n13646), .ZN(n13648) );
  NAND2_X1 U17075 ( .A1(n13649), .A2(n13648), .ZN(n14438) );
  INV_X1 U17076 ( .A(P1_EAX_REG_2__SCAN_IN), .ZN(n19990) );
  INV_X1 U17077 ( .A(n20126), .ZN(n13650) );
  OAI222_X1 U17078 ( .A1(n14566), .A2(n14438), .B1(n14529), .B2(n19990), .C1(
        n14155), .C2(n13650), .ZN(P1_U2902) );
  OAI21_X1 U17079 ( .B1(n13652), .B2(n13651), .A(n13713), .ZN(n14429) );
  INV_X1 U17080 ( .A(P1_EBX_REG_2__SCAN_IN), .ZN(n13653) );
  OAI222_X1 U17081 ( .A1(n14429), .A2(n19962), .B1(n13653), .B2(n19968), .C1(
        n14438), .C2(n14496), .ZN(P1_U2870) );
  NOR2_X1 U17082 ( .A1(P1_FLUSH_REG_SCAN_IN), .A2(n16000), .ZN(n13693) );
  OR2_X1 U17083 ( .A1(n13655), .A2(n14281), .ZN(n13666) );
  XNOR2_X1 U17084 ( .A(n13673), .B(n11235), .ZN(n13660) );
  NAND3_X1 U17085 ( .A1(n14281), .A2(n13656), .A3(n13660), .ZN(n13664) );
  INV_X1 U17086 ( .A(n13657), .ZN(n13659) );
  OR2_X1 U17087 ( .A1(n13659), .A2(n13658), .ZN(n13677) );
  INV_X1 U17088 ( .A(n13660), .ZN(n14864) );
  XNOR2_X1 U17089 ( .A(n13661), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(
        n13662) );
  AOI22_X1 U17090 ( .A1(n13677), .A2(n14864), .B1(n15697), .B2(n13662), .ZN(
        n13663) );
  AND2_X1 U17091 ( .A1(n13664), .A2(n13663), .ZN(n13665) );
  NAND2_X1 U17092 ( .A1(n13666), .A2(n13665), .ZN(n14859) );
  MUX2_X1 U17093 ( .A(n14859), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n15699), .Z(n15703) );
  AOI22_X1 U17094 ( .A1(n13693), .A2(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B1(
        n15703), .B2(n16000), .ZN(n13686) );
  INV_X1 U17095 ( .A(n14281), .ZN(n13683) );
  INV_X1 U17096 ( .A(n13667), .ZN(n13674) );
  OAI211_X1 U17097 ( .C1(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(n13673), .A(
        n13668), .B(n13674), .ZN(n20757) );
  NOR3_X1 U17098 ( .A1(n13683), .A2(n13669), .A3(n20757), .ZN(n13682) );
  NAND2_X1 U17099 ( .A1(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        P1_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n13671) );
  INV_X1 U17100 ( .A(n13671), .ZN(n13670) );
  MUX2_X1 U17101 ( .A(n13671), .B(n13670), .S(
        P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .Z(n13679) );
  INV_X1 U17102 ( .A(n13672), .ZN(n13676) );
  MUX2_X1 U17103 ( .A(n13674), .B(n10990), .S(n13673), .Z(n13675) );
  NAND3_X1 U17104 ( .A1(n13677), .A2(n13676), .A3(n13675), .ZN(n13678) );
  OAI21_X1 U17105 ( .B1(n13680), .B2(n13679), .A(n13678), .ZN(n13681) );
  AOI211_X1 U17106 ( .C1(n20771), .C2(n13683), .A(n13682), .B(n13681), .ZN(
        n20760) );
  NAND2_X1 U17107 ( .A1(n15699), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n13684) );
  OAI21_X1 U17108 ( .B1(n15699), .B2(n20760), .A(n13684), .ZN(n15708) );
  AOI22_X1 U17109 ( .A1(n13693), .A2(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B1(
        n16000), .B2(n15708), .ZN(n13685) );
  NOR2_X1 U17110 ( .A1(n13686), .A2(n13685), .ZN(n15717) );
  INV_X1 U17111 ( .A(n13687), .ZN(n13688) );
  NAND2_X1 U17112 ( .A1(n15717), .A2(n13688), .ZN(n13728) );
  AND2_X1 U17113 ( .A1(n19922), .A2(n13689), .ZN(n13692) );
  NAND2_X1 U17114 ( .A1(n15699), .A2(n13690), .ZN(n13691) );
  OAI211_X1 U17115 ( .C1(n15699), .C2(n13692), .A(n13691), .B(n16000), .ZN(
        n13695) );
  NAND2_X1 U17116 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n13693), .ZN(
        n13694) );
  AND2_X1 U17117 ( .A1(n13695), .A2(n13694), .ZN(n15714) );
  NAND3_X1 U17118 ( .A1(n13728), .A2(n15714), .A3(n19864), .ZN(n13697) );
  INV_X1 U17119 ( .A(n16001), .ZN(n13696) );
  NAND2_X1 U17120 ( .A1(n13697), .A2(n13696), .ZN(n13699) );
  NAND2_X1 U17121 ( .A1(n11192), .A2(n15723), .ZN(n20795) );
  NAND2_X1 U17122 ( .A1(n13699), .A2(n20262), .ZN(n20773) );
  NAND2_X1 U17123 ( .A1(P1_STATE2_REG_1__SCAN_IN), .A2(n20388), .ZN(n20772) );
  INV_X1 U17124 ( .A(n20772), .ZN(n14855) );
  NAND2_X1 U17125 ( .A1(n13700), .A2(P1_STATEBS16_REG_SCAN_IN), .ZN(n20634) );
  OAI211_X1 U17126 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n13700), .A(n20634), 
        .B(n20581), .ZN(n13701) );
  OAI21_X1 U17127 ( .B1(n14855), .B2(n20380), .A(n13701), .ZN(n13702) );
  NAND2_X1 U17128 ( .A1(n20773), .A2(n13702), .ZN(n13703) );
  OAI21_X1 U17129 ( .B1(n20773), .B2(n20440), .A(n13703), .ZN(P1_U3477) );
  XNOR2_X1 U17130 ( .A(n13574), .B(n13746), .ZN(n13708) );
  NOR2_X1 U17131 ( .A1(n13705), .A2(n13704), .ZN(n13706) );
  OR2_X1 U17132 ( .A1(n13742), .A2(n13706), .ZN(n15498) );
  MUX2_X1 U17133 ( .A(n10729), .B(n15498), .S(n14993), .Z(n13707) );
  OAI21_X1 U17134 ( .B1(n13708), .B2(n15009), .A(n13707), .ZN(P2_U2878) );
  OAI21_X1 U17135 ( .B1(n13711), .B2(n13710), .A(n13775), .ZN(n13781) );
  NAND2_X1 U17136 ( .A1(n13713), .A2(n13712), .ZN(n13714) );
  NAND2_X1 U17137 ( .A1(n13778), .A2(n13714), .ZN(n19936) );
  INV_X1 U17138 ( .A(n19936), .ZN(n13715) );
  AOI22_X1 U17139 ( .A1(n15856), .A2(n13715), .B1(P1_EBX_REG_3__SCAN_IN), .B2(
        n14492), .ZN(n13716) );
  OAI21_X1 U17140 ( .B1(n13781), .B2(n14496), .A(n13716), .ZN(P1_U2869) );
  XOR2_X1 U17141 ( .A(n19799), .B(n19804), .Z(n13722) );
  XNOR2_X1 U17142 ( .A(n13717), .B(n13718), .ZN(n19003) );
  NAND2_X1 U17143 ( .A1(n19808), .A2(n19003), .ZN(n13719) );
  OAI21_X1 U17144 ( .B1(n19808), .B2(n19003), .A(n13719), .ZN(n19007) );
  NOR2_X1 U17145 ( .A1(n19007), .A2(n19008), .ZN(n19006) );
  INV_X1 U17146 ( .A(n13719), .ZN(n13720) );
  NOR2_X1 U17147 ( .A1(n19006), .A2(n13720), .ZN(n13721) );
  NOR2_X1 U17148 ( .A1(n13722), .A2(n13721), .ZN(n13833) );
  AOI21_X1 U17149 ( .B1(n13722), .B2(n13721), .A(n13833), .ZN(n13726) );
  INV_X1 U17150 ( .A(n19125), .ZN(n16118) );
  AOI22_X1 U17151 ( .A1(n18989), .A2(n16118), .B1(P2_EAX_REG_2__SCAN_IN), .B2(
        n19004), .ZN(n13725) );
  INV_X1 U17152 ( .A(n19799), .ZN(n13723) );
  NAND2_X1 U17153 ( .A1(n13723), .A2(n19005), .ZN(n13724) );
  OAI211_X1 U17154 ( .C1(n13726), .C2(n19009), .A(n13725), .B(n13724), .ZN(
        P2_U2917) );
  NAND3_X1 U17155 ( .A1(n13728), .A2(n15714), .A3(n13727), .ZN(n15719) );
  INV_X1 U17156 ( .A(n15719), .ZN(n13730) );
  OAI22_X1 U17157 ( .A1(n9828), .A2(n20767), .B1(n14282), .B2(n14855), .ZN(
        n13729) );
  OAI21_X1 U17158 ( .B1(n13730), .B2(n13729), .A(n20773), .ZN(n13731) );
  OAI21_X1 U17159 ( .B1(n20773), .B2(n20551), .A(n13731), .ZN(P1_U3478) );
  XOR2_X1 U17160 ( .A(n13733), .B(n13732), .Z(n20068) );
  NAND2_X1 U17161 ( .A1(n20068), .A2(n20043), .ZN(n13737) );
  INV_X1 U17162 ( .A(P1_REIP_REG_2__SCAN_IN), .ZN(n13734) );
  NOR2_X1 U17163 ( .A1(n20046), .A2(n13734), .ZN(n20060) );
  NOR2_X1 U17164 ( .A1(n15909), .A2(n14431), .ZN(n13735) );
  AOI211_X1 U17165 ( .C1(n20038), .C2(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .A(
        n20060), .B(n13735), .ZN(n13736) );
  OAI211_X1 U17166 ( .C1(n20048), .C2(n14438), .A(n13737), .B(n13736), .ZN(
        P1_U2997) );
  OAI21_X1 U17167 ( .B1(n13740), .B2(n13739), .A(n13738), .ZN(n18894) );
  INV_X1 U17168 ( .A(P2_EAX_REG_11__SCAN_IN), .ZN(n19055) );
  OAI222_X1 U17169 ( .A1(n18894), .A2(n18995), .B1(n15039), .B2(n19013), .C1(
        n19055), .C2(n15083), .ZN(P2_U2908) );
  OR2_X1 U17170 ( .A1(n13742), .A2(n13741), .ZN(n13744) );
  NAND2_X1 U17171 ( .A1(n13744), .A2(n13743), .ZN(n18900) );
  OAI21_X1 U17172 ( .B1(n13574), .B2(n13746), .A(n13745), .ZN(n13748) );
  NAND3_X1 U17173 ( .A1(n13748), .A2(n14965), .A3(n13747), .ZN(n13750) );
  NAND2_X1 U17174 ( .A1(n15006), .A2(P2_EBX_REG_10__SCAN_IN), .ZN(n13749) );
  OAI211_X1 U17175 ( .C1(n18900), .C2(n15006), .A(n13750), .B(n13749), .ZN(
        P2_U2877) );
  INV_X1 U17176 ( .A(P1_EAX_REG_3__SCAN_IN), .ZN(n19988) );
  INV_X1 U17177 ( .A(n20130), .ZN(n13751) );
  OAI222_X1 U17178 ( .A1(n14566), .A2(n13781), .B1(n14529), .B2(n19988), .C1(
        n14155), .C2(n13751), .ZN(P1_U2901) );
  XNOR2_X1 U17179 ( .A(n13753), .B(n13752), .ZN(n13786) );
  NOR2_X1 U17180 ( .A1(n20069), .A2(n20087), .ZN(n14010) );
  AOI21_X1 U17181 ( .B1(n14010), .B2(n20070), .A(n20062), .ZN(n14819) );
  NAND2_X1 U17182 ( .A1(n15986), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n13783) );
  OAI21_X1 U17183 ( .B1(n15975), .B2(n19936), .A(n13783), .ZN(n13755) );
  NOR2_X1 U17184 ( .A1(n20066), .A2(n14010), .ZN(n13856) );
  AOI211_X1 U17185 ( .C1(n20062), .C2(n20064), .A(n14788), .B(n13856), .ZN(
        n20053) );
  NOR2_X1 U17186 ( .A1(n20053), .A2(n13756), .ZN(n13754) );
  AOI211_X1 U17187 ( .C1(n20057), .C2(n13756), .A(n13755), .B(n13754), .ZN(
        n13757) );
  OAI21_X1 U17188 ( .B1(n20095), .B2(n13786), .A(n13757), .ZN(P1_U3028) );
  INV_X1 U17189 ( .A(P1_EAX_REG_16__SCAN_IN), .ZN(n21034) );
  AOI22_X1 U17190 ( .A1(n19993), .A2(P1_UWORD_REG_0__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_16__SCAN_IN), .ZN(n13758) );
  OAI21_X1 U17191 ( .B1(n21034), .B2(n13772), .A(n13758), .ZN(P1_U2920) );
  INV_X1 U17192 ( .A(P1_EAX_REG_29__SCAN_IN), .ZN(n20013) );
  AOI22_X1 U17193 ( .A1(n19993), .A2(P1_UWORD_REG_13__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_29__SCAN_IN), .ZN(n13759) );
  OAI21_X1 U17194 ( .B1(n20013), .B2(n13772), .A(n13759), .ZN(P1_U2907) );
  INV_X1 U17195 ( .A(P1_EAX_REG_22__SCAN_IN), .ZN(n13761) );
  AOI22_X1 U17196 ( .A1(n19993), .A2(P1_UWORD_REG_6__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_22__SCAN_IN), .ZN(n13760) );
  OAI21_X1 U17197 ( .B1(n13761), .B2(n13772), .A(n13760), .ZN(P1_U2914) );
  INV_X1 U17198 ( .A(P1_EAX_REG_18__SCAN_IN), .ZN(n13763) );
  AOI22_X1 U17199 ( .A1(n19993), .A2(P1_UWORD_REG_2__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_18__SCAN_IN), .ZN(n13762) );
  OAI21_X1 U17200 ( .B1(n13763), .B2(n13772), .A(n13762), .ZN(P1_U2918) );
  INV_X1 U17201 ( .A(P1_EAX_REG_17__SCAN_IN), .ZN(n13765) );
  AOI22_X1 U17202 ( .A1(n19993), .A2(P1_UWORD_REG_1__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_17__SCAN_IN), .ZN(n13764) );
  OAI21_X1 U17203 ( .B1(n13765), .B2(n13772), .A(n13764), .ZN(P1_U2919) );
  AOI22_X1 U17204 ( .A1(n19993), .A2(P1_UWORD_REG_10__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_26__SCAN_IN), .ZN(n13766) );
  OAI21_X1 U17205 ( .B1(n14521), .B2(n13772), .A(n13766), .ZN(P1_U2910) );
  INV_X1 U17206 ( .A(P1_EAX_REG_21__SCAN_IN), .ZN(n13768) );
  AOI22_X1 U17207 ( .A1(n19993), .A2(P1_UWORD_REG_5__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_21__SCAN_IN), .ZN(n13767) );
  OAI21_X1 U17208 ( .B1(n13768), .B2(n13772), .A(n13767), .ZN(P1_U2915) );
  INV_X1 U17209 ( .A(P1_EAX_REG_20__SCAN_IN), .ZN(n13770) );
  AOI22_X1 U17210 ( .A1(n19993), .A2(P1_UWORD_REG_4__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_20__SCAN_IN), .ZN(n13769) );
  OAI21_X1 U17211 ( .B1(n13770), .B2(n13772), .A(n13769), .ZN(P1_U2916) );
  INV_X1 U17212 ( .A(P1_EAX_REG_19__SCAN_IN), .ZN(n13773) );
  AOI22_X1 U17213 ( .A1(n19993), .A2(P1_UWORD_REG_3__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_19__SCAN_IN), .ZN(n13771) );
  OAI21_X1 U17214 ( .B1(n13773), .B2(n13772), .A(n13771), .ZN(P1_U2917) );
  AOI21_X1 U17215 ( .B1(n13776), .B2(n13775), .A(n13774), .ZN(n13777) );
  INV_X1 U17216 ( .A(n13777), .ZN(n19926) );
  AOI21_X1 U17217 ( .B1(n13779), .B2(n13778), .A(n13815), .ZN(n20051) );
  AOI22_X1 U17218 ( .A1(n15856), .A2(n20051), .B1(P1_EBX_REG_4__SCAN_IN), .B2(
        n14492), .ZN(n13780) );
  OAI21_X1 U17219 ( .B1(n19926), .B2(n14496), .A(n13780), .ZN(P1_U2868) );
  INV_X1 U17220 ( .A(n13781), .ZN(n19944) );
  NAND2_X1 U17221 ( .A1(n20038), .A2(P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13782) );
  OAI211_X1 U17222 ( .C1(n15909), .C2(n19940), .A(n13783), .B(n13782), .ZN(
        n13784) );
  AOI21_X1 U17223 ( .B1(n19944), .B2(n20101), .A(n13784), .ZN(n13785) );
  OAI21_X1 U17224 ( .B1(n13786), .B2(n19863), .A(n13785), .ZN(P1_U2996) );
  INV_X1 U17225 ( .A(P1_EAX_REG_4__SCAN_IN), .ZN(n19986) );
  INV_X1 U17226 ( .A(n20133), .ZN(n13787) );
  OAI222_X1 U17227 ( .A1(n14566), .A2(n19926), .B1(n14529), .B2(n19986), .C1(
        n14155), .C2(n13787), .ZN(P1_U2900) );
  INV_X1 U17228 ( .A(n13738), .ZN(n13788) );
  OAI21_X1 U17229 ( .B1(n13789), .B2(n13788), .A(n10192), .ZN(n18875) );
  INV_X1 U17230 ( .A(n15029), .ZN(n13790) );
  INV_X1 U17231 ( .A(P2_EAX_REG_12__SCAN_IN), .ZN(n19053) );
  OAI222_X1 U17232 ( .A1(n18875), .A2(n18995), .B1(n13790), .B2(n19013), .C1(
        n19053), .C2(n15083), .ZN(P2_U2907) );
  INV_X1 U17233 ( .A(P2_EBX_REG_11__SCAN_IN), .ZN(n21018) );
  INV_X1 U17234 ( .A(n13747), .ZN(n13794) );
  INV_X1 U17235 ( .A(n13791), .ZN(n13792) );
  OAI211_X1 U17236 ( .C1(n13794), .C2(n13793), .A(n13792), .B(n14965), .ZN(
        n13800) );
  NAND2_X1 U17237 ( .A1(n13795), .A2(n13743), .ZN(n13798) );
  INV_X1 U17238 ( .A(n13796), .ZN(n13797) );
  NAND2_X1 U17239 ( .A1(n14993), .A2(n18889), .ZN(n13799) );
  OAI211_X1 U17240 ( .C1(n14993), .C2(n21018), .A(n13800), .B(n13799), .ZN(
        P2_U2876) );
  OAI21_X1 U17241 ( .B1(n13802), .B2(n13801), .A(n14019), .ZN(n18867) );
  INV_X1 U17242 ( .A(n15019), .ZN(n13803) );
  INV_X1 U17243 ( .A(P2_EAX_REG_13__SCAN_IN), .ZN(n19051) );
  OAI222_X1 U17244 ( .A1(n18867), .A2(n18995), .B1(n13803), .B2(n19013), .C1(
        n19051), .C2(n15083), .ZN(P2_U2906) );
  OR2_X1 U17245 ( .A1(n13774), .A2(n13806), .ZN(n13807) );
  AND2_X1 U17246 ( .A1(n13805), .A2(n13807), .ZN(n19918) );
  INV_X1 U17247 ( .A(n19918), .ZN(n13817) );
  AOI22_X1 U17248 ( .A1(n14163), .A2(n20136), .B1(P1_EAX_REG_5__SCAN_IN), .B2(
        n14558), .ZN(n13808) );
  OAI21_X1 U17249 ( .B1(n13817), .B2(n14566), .A(n13808), .ZN(P1_U2899) );
  OR2_X1 U17250 ( .A1(n13809), .A2(n13796), .ZN(n13810) );
  NAND2_X1 U17251 ( .A1(n13842), .A2(n13810), .ZN(n18874) );
  NAND2_X1 U17252 ( .A1(n13791), .A2(n13811), .ZN(n13845) );
  OAI211_X1 U17253 ( .C1(n13791), .C2(n13811), .A(n13845), .B(n14965), .ZN(
        n13813) );
  NAND2_X1 U17254 ( .A1(n15006), .A2(P2_EBX_REG_12__SCAN_IN), .ZN(n13812) );
  OAI211_X1 U17255 ( .C1(n18874), .C2(n15006), .A(n13813), .B(n13812), .ZN(
        P2_U2875) );
  NOR2_X1 U17256 ( .A1(n13815), .A2(n13814), .ZN(n13816) );
  OR2_X1 U17257 ( .A1(n15983), .A2(n13816), .ZN(n19916) );
  INV_X1 U17258 ( .A(P1_EBX_REG_5__SCAN_IN), .ZN(n13818) );
  OAI222_X1 U17259 ( .A1(n19916), .A2(n19962), .B1(n13818), .B2(n19968), .C1(
        n13817), .C2(n14496), .ZN(P1_U2867) );
  XOR2_X1 U17260 ( .A(n13820), .B(n13819), .Z(n20055) );
  NAND2_X1 U17261 ( .A1(n20055), .A2(n20043), .ZN(n13823) );
  INV_X1 U17262 ( .A(P1_REIP_REG_4__SCAN_IN), .ZN(n20710) );
  NOR2_X1 U17263 ( .A1(n20046), .A2(n20710), .ZN(n20050) );
  NOR2_X1 U17264 ( .A1(n15909), .A2(n19925), .ZN(n13821) );
  AOI211_X1 U17265 ( .C1(n20038), .C2(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n20050), .B(n13821), .ZN(n13822) );
  OAI211_X1 U17266 ( .C1(n20048), .C2(n19926), .A(n13823), .B(n13822), .ZN(
        P1_U2995) );
  NAND2_X1 U17267 ( .A1(n13805), .A2(n13825), .ZN(n13826) );
  AND2_X1 U17268 ( .A1(n13824), .A2(n13826), .ZN(n19965) );
  INV_X1 U17269 ( .A(n19965), .ZN(n13828) );
  INV_X1 U17270 ( .A(n20139), .ZN(n13827) );
  OAI222_X1 U17271 ( .A1(n14566), .A2(n13828), .B1(n14529), .B2(n12032), .C1(
        n14155), .C2(n13827), .ZN(P1_U2898) );
  OR2_X1 U17272 ( .A1(n13830), .A2(n13829), .ZN(n13832) );
  NAND2_X1 U17273 ( .A1(n13832), .A2(n13831), .ZN(n18996) );
  AOI21_X1 U17274 ( .B1(n19799), .B2(n13834), .A(n13833), .ZN(n18999) );
  XNOR2_X1 U17275 ( .A(n19788), .B(n18996), .ZN(n18998) );
  NOR2_X1 U17276 ( .A1(n18999), .A2(n18998), .ZN(n18997) );
  AOI21_X1 U17277 ( .B1(n18996), .B2(n19788), .A(n18997), .ZN(n13836) );
  XNOR2_X1 U17278 ( .A(n13831), .B(n13835), .ZN(n14036) );
  NOR2_X1 U17279 ( .A1(n13836), .A2(n14036), .ZN(n18991) );
  XNOR2_X1 U17280 ( .A(n18991), .B(n18990), .ZN(n13839) );
  AOI22_X1 U17281 ( .A1(n19005), .A2(n14036), .B1(n19004), .B2(
        P2_EAX_REG_4__SCAN_IN), .ZN(n13838) );
  INV_X1 U17282 ( .A(n13948), .ZN(n16112) );
  NAND2_X1 U17283 ( .A1(n18989), .A2(n16112), .ZN(n13837) );
  OAI211_X1 U17284 ( .C1(n13839), .C2(n19009), .A(n13838), .B(n13837), .ZN(
        P2_U2915) );
  NAND2_X1 U17285 ( .A1(n13842), .A2(n13841), .ZN(n13843) );
  AND2_X1 U17286 ( .A1(n13840), .A2(n13843), .ZN(n18862) );
  INV_X1 U17287 ( .A(n18862), .ZN(n15447) );
  INV_X1 U17288 ( .A(n13845), .ZN(n13961) );
  OAI211_X1 U17289 ( .C1(n13961), .C2(n13846), .A(n14965), .B(n13909), .ZN(
        n13848) );
  NAND2_X1 U17290 ( .A1(n15006), .A2(P2_EBX_REG_13__SCAN_IN), .ZN(n13847) );
  OAI211_X1 U17291 ( .C1(n15447), .C2(n15006), .A(n13848), .B(n13847), .ZN(
        P2_U2874) );
  INV_X1 U17292 ( .A(n13849), .ZN(n13850) );
  OAI21_X1 U17293 ( .B1(n13851), .B2(n9851), .A(n13850), .ZN(n18851) );
  OAI222_X1 U17294 ( .A1(n18851), .A2(n18995), .B1(n15083), .B2(n13355), .C1(
        n13852), .C2(n19013), .ZN(P2_U2904) );
  XOR2_X1 U17295 ( .A(n13854), .B(n13853), .Z(n15910) );
  OAI21_X1 U17296 ( .B1(n14008), .B2(n14786), .A(n20065), .ZN(n14011) );
  AND2_X1 U17297 ( .A1(n14845), .A2(n20056), .ZN(n13855) );
  OR2_X1 U17298 ( .A1(n13856), .A2(n13855), .ZN(n13857) );
  NOR2_X1 U17299 ( .A1(n14011), .A2(n13857), .ZN(n15963) );
  NOR2_X1 U17300 ( .A1(n20056), .A2(P1_INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(
        n15962) );
  NAND2_X1 U17301 ( .A1(n20057), .A2(n15962), .ZN(n13862) );
  INV_X1 U17302 ( .A(n19916), .ZN(n13860) );
  INV_X1 U17303 ( .A(P1_REIP_REG_5__SCAN_IN), .ZN(n13858) );
  OR2_X1 U17304 ( .A1(n20046), .A2(n13858), .ZN(n15913) );
  INV_X1 U17305 ( .A(n15913), .ZN(n13859) );
  AOI21_X1 U17306 ( .B1(n20089), .B2(n13860), .A(n13859), .ZN(n13861) );
  OAI211_X1 U17307 ( .C1(n11348), .C2(n15963), .A(n13862), .B(n13861), .ZN(
        n13863) );
  AOI21_X1 U17308 ( .B1(n15910), .B2(n20077), .A(n13863), .ZN(n13864) );
  INV_X1 U17309 ( .A(n13864), .ZN(P1_U3026) );
  NAND2_X1 U17310 ( .A1(n13866), .A2(n13865), .ZN(n13867) );
  XNOR2_X1 U17311 ( .A(n13867), .B(n13924), .ZN(n19093) );
  OAI21_X1 U17312 ( .B1(n13868), .B2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A(
        n14250), .ZN(n13870) );
  NAND2_X1 U17313 ( .A1(n13868), .A2(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n13869) );
  NAND2_X1 U17314 ( .A1(n13870), .A2(n13869), .ZN(n13872) );
  XNOR2_X1 U17315 ( .A(n14038), .B(n13924), .ZN(n13871) );
  XNOR2_X1 U17316 ( .A(n13872), .B(n13871), .ZN(n19088) );
  NOR2_X1 U17317 ( .A1(n10009), .A2(n16230), .ZN(n13986) );
  INV_X1 U17318 ( .A(n13986), .ZN(n13923) );
  OAI21_X1 U17319 ( .B1(n13875), .B2(n13874), .A(n13873), .ZN(n14088) );
  NOR2_X1 U17320 ( .A1(n10009), .A2(n14088), .ZN(n16231) );
  NOR2_X1 U17321 ( .A1(n15471), .A2(n16231), .ZN(n13928) );
  NOR2_X1 U17322 ( .A1(n12700), .A2(n18934), .ZN(n13876) );
  AOI21_X1 U17323 ( .B1(n16209), .B2(n14036), .A(n13876), .ZN(n13877) );
  OAI21_X1 U17324 ( .B1(n13878), .B2(n16212), .A(n13877), .ZN(n13879) );
  AOI21_X1 U17325 ( .B1(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n13928), .A(
        n13879), .ZN(n13880) );
  OAI21_X1 U17326 ( .B1(n13923), .B2(P2_INSTADDRPOINTER_REG_4__SCAN_IN), .A(
        n13880), .ZN(n13881) );
  AOI21_X1 U17327 ( .B1(n19088), .B2(n16227), .A(n13881), .ZN(n13882) );
  OAI21_X1 U17328 ( .B1(n16223), .B2(n19093), .A(n13882), .ZN(P2_U3042) );
  NAND2_X1 U17329 ( .A1(n13824), .A2(n13884), .ZN(n13885) );
  AND2_X1 U17330 ( .A1(n13899), .A2(n13885), .ZN(n19897) );
  INV_X1 U17331 ( .A(n19897), .ZN(n13889) );
  INV_X1 U17332 ( .A(P1_EBX_REG_7__SCAN_IN), .ZN(n21080) );
  NAND2_X1 U17333 ( .A1(n15985), .A2(n13886), .ZN(n13887) );
  NAND2_X1 U17334 ( .A1(n13902), .A2(n13887), .ZN(n19895) );
  OAI222_X1 U17335 ( .A1(n13889), .A2(n14496), .B1(n19968), .B2(n21080), .C1(
        n19895), .C2(n19962), .ZN(P1_U2865) );
  INV_X1 U17336 ( .A(P1_EAX_REG_7__SCAN_IN), .ZN(n19981) );
  INV_X1 U17337 ( .A(n20148), .ZN(n13888) );
  OAI222_X1 U17338 ( .A1(n14566), .A2(n13889), .B1(n14529), .B2(n19981), .C1(
        n14155), .C2(n13888), .ZN(P1_U2897) );
  INV_X1 U17339 ( .A(n13909), .ZN(n13892) );
  OR2_X1 U17340 ( .A1(n13909), .A2(n13890), .ZN(n13907) );
  OAI211_X1 U17341 ( .C1(n13892), .C2(n13891), .A(n14965), .B(n13907), .ZN(
        n13897) );
  INV_X1 U17342 ( .A(n13893), .ZN(n13894) );
  AOI21_X1 U17343 ( .B1(n13895), .B2(n13840), .A(n13894), .ZN(n16193) );
  NAND2_X1 U17344 ( .A1(n16193), .A2(n14993), .ZN(n13896) );
  OAI211_X1 U17345 ( .C1(n14993), .C2(n13898), .A(n13897), .B(n13896), .ZN(
        P2_U2873) );
  AOI21_X1 U17346 ( .B1(n13900), .B2(n13899), .A(n9907), .ZN(n13957) );
  INV_X1 U17347 ( .A(n13957), .ZN(n14426) );
  NAND2_X1 U17348 ( .A1(n13902), .A2(n13901), .ZN(n13903) );
  AND2_X1 U17349 ( .A1(n13976), .A2(n13903), .ZN(n15967) );
  AOI22_X1 U17350 ( .A1(n15856), .A2(n15967), .B1(P1_EBX_REG_8__SCAN_IN), .B2(
        n14492), .ZN(n13904) );
  OAI21_X1 U17351 ( .B1(n14426), .B2(n14496), .A(n13904), .ZN(P1_U2864) );
  INV_X1 U17352 ( .A(P1_EAX_REG_8__SCAN_IN), .ZN(n13906) );
  INV_X1 U17353 ( .A(DATAI_8_), .ZN(n13905) );
  INV_X1 U17354 ( .A(BUF1_REG_8__SCAN_IN), .ZN(n16390) );
  MUX2_X1 U17355 ( .A(n13905), .B(n16390), .S(n14173), .Z(n19997) );
  OAI222_X1 U17356 ( .A1(n14426), .A2(n14566), .B1(n13906), .B2(n14529), .C1(
        n14155), .C2(n19997), .ZN(P1_U2896) );
  INV_X1 U17357 ( .A(P2_EBX_REG_15__SCAN_IN), .ZN(n21015) );
  INV_X1 U17358 ( .A(n13907), .ZN(n13912) );
  NOR2_X1 U17359 ( .A1(n13909), .A2(n13908), .ZN(n13963) );
  INV_X1 U17360 ( .A(n13963), .ZN(n13910) );
  OAI211_X1 U17361 ( .C1(n13912), .C2(n13911), .A(n13910), .B(n14965), .ZN(
        n13916) );
  AND2_X1 U17362 ( .A1(n13893), .A2(n13913), .ZN(n13914) );
  OR2_X1 U17363 ( .A1(n13914), .A2(n13967), .ZN(n15254) );
  NAND2_X1 U17364 ( .A1(n18847), .A2(n14993), .ZN(n13915) );
  OAI211_X1 U17365 ( .C1(n14993), .C2(n21015), .A(n13916), .B(n13915), .ZN(
        P2_U2872) );
  INV_X1 U17366 ( .A(n10878), .ZN(n13920) );
  AND2_X1 U17367 ( .A1(n10878), .A2(n13917), .ZN(n13919) );
  OAI22_X1 U17368 ( .A1(n10877), .A2(n13920), .B1(n13919), .B2(n13918), .ZN(
        n16186) );
  XNOR2_X1 U17369 ( .A(n13921), .B(n13922), .ZN(n16185) );
  NOR2_X1 U17370 ( .A1(n10904), .A2(n18934), .ZN(n13927) );
  AOI211_X1 U17371 ( .C1(n13925), .C2(n13924), .A(n13991), .B(n13923), .ZN(
        n13926) );
  AOI211_X1 U17372 ( .C1(P2_INSTADDRPOINTER_REG_5__SCAN_IN), .C2(n13928), .A(
        n13927), .B(n13926), .ZN(n13933) );
  OAI21_X1 U17373 ( .B1(n9872), .B2(n13930), .A(n13929), .ZN(n18994) );
  OAI22_X1 U17374 ( .A1(n18994), .A2(n16222), .B1(n16212), .B2(n18936), .ZN(
        n13931) );
  INV_X1 U17375 ( .A(n13931), .ZN(n13932) );
  OAI211_X1 U17376 ( .C1(n16185), .C2(n16217), .A(n13933), .B(n13932), .ZN(
        n13934) );
  INV_X1 U17377 ( .A(n13934), .ZN(n13935) );
  OAI21_X1 U17378 ( .B1(n16186), .B2(n16223), .A(n13935), .ZN(P2_U3041) );
  NOR2_X2 U17379 ( .A1(n19556), .A2(n19789), .ZN(n19702) );
  INV_X1 U17380 ( .A(n19408), .ZN(n19160) );
  NAND2_X1 U17381 ( .A1(n19160), .A2(n19253), .ZN(n19179) );
  OAI21_X1 U17382 ( .B1(n19702), .B2(n19182), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n13936) );
  NAND2_X1 U17383 ( .A1(n13936), .A2(n19612), .ZN(n13947) );
  INV_X1 U17384 ( .A(n13947), .ZN(n13940) );
  NOR2_X1 U17385 ( .A1(n13937), .A2(n19796), .ZN(n19695) );
  NAND2_X1 U17386 ( .A1(n19796), .A2(n16248), .ZN(n19219) );
  OR2_X1 U17387 ( .A1(n19219), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19162) );
  NOR2_X1 U17388 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19162), .ZN(
        n19149) );
  NOR2_X1 U17389 ( .A1(n19695), .A2(n19149), .ZN(n13946) );
  AOI211_X1 U17390 ( .C1(n9879), .C2(n19798), .A(n19149), .B(n19612), .ZN(
        n13939) );
  OAI21_X1 U17391 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(
        P2_STATE2_REG_1__SCAN_IN), .A(n10983), .ZN(n19841) );
  INV_X1 U17392 ( .A(BUF2_REG_28__SCAN_IN), .ZN(n18118) );
  INV_X1 U17393 ( .A(BUF1_REG_28__SCAN_IN), .ZN(n16364) );
  OAI22_X2 U17394 ( .A1(n18118), .A2(n19144), .B1(n16364), .B2(n19146), .ZN(
        n19680) );
  AOI22_X2 U17395 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n19151), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n19152), .ZN(n19583) );
  INV_X1 U17396 ( .A(n19149), .ZN(n13943) );
  NAND2_X1 U17397 ( .A1(P2_STATE2_REG_3__SCAN_IN), .A2(n19648), .ZN(n19139) );
  NAND2_X1 U17398 ( .A1(n13942), .A2(n19148), .ZN(n19578) );
  OAI22_X1 U17399 ( .A1(n19583), .A2(n19179), .B1(n13943), .B2(n19578), .ZN(
        n13944) );
  AOI21_X1 U17400 ( .B1(n19702), .B2(n19680), .A(n13944), .ZN(n13950) );
  OAI21_X1 U17401 ( .B1(n9879), .B2(n19149), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n13945) );
  NOR2_X2 U17402 ( .A1(n13948), .A2(n19613), .ZN(n19678) );
  NAND2_X1 U17403 ( .A1(n19153), .A2(n19678), .ZN(n13949) );
  OAI211_X1 U17404 ( .C1(n19157), .C2(n13951), .A(n13950), .B(n13949), .ZN(
        P2_U3052) );
  XNOR2_X1 U17405 ( .A(n13952), .B(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13953) );
  XNOR2_X1 U17406 ( .A(n13954), .B(n13953), .ZN(n15970) );
  INV_X1 U17407 ( .A(n15970), .ZN(n13959) );
  NAND2_X1 U17408 ( .A1(n20038), .A2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(
        n13955) );
  NAND2_X1 U17409 ( .A1(n15986), .A2(P1_REIP_REG_8__SCAN_IN), .ZN(n15965) );
  OAI211_X1 U17410 ( .C1(n15909), .C2(n14417), .A(n13955), .B(n15965), .ZN(
        n13956) );
  AOI21_X1 U17411 ( .B1(n13957), .B2(n20101), .A(n13956), .ZN(n13958) );
  OAI21_X1 U17412 ( .B1(n13959), .B2(n19863), .A(n13958), .ZN(P1_U2991) );
  AND2_X1 U17413 ( .A1(n13961), .A2(n13960), .ZN(n13999) );
  NOR2_X1 U17414 ( .A1(n13963), .A2(n13962), .ZN(n13964) );
  OR2_X1 U17415 ( .A1(n13999), .A2(n13964), .ZN(n18970) );
  OR2_X1 U17416 ( .A1(n13967), .A2(n13966), .ZN(n13968) );
  NAND2_X1 U17417 ( .A1(n13965), .A2(n13968), .ZN(n18835) );
  NOR2_X1 U17418 ( .A1(n15006), .A2(n18835), .ZN(n13969) );
  AOI21_X1 U17419 ( .B1(P2_EBX_REG_16__SCAN_IN), .B2(n15006), .A(n13969), .ZN(
        n13970) );
  OAI21_X1 U17420 ( .B1(n18970), .B2(n15009), .A(n13970), .ZN(P2_U2871) );
  NOR2_X1 U17421 ( .A1(n9907), .A2(n13973), .ZN(n13974) );
  OR2_X1 U17422 ( .A1(n13972), .A2(n13974), .ZN(n19885) );
  INV_X1 U17423 ( .A(P1_EBX_REG_9__SCAN_IN), .ZN(n13978) );
  AND2_X1 U17424 ( .A1(n13976), .A2(n13975), .ZN(n13977) );
  OR2_X1 U17425 ( .A1(n13977), .A2(n14057), .ZN(n19883) );
  OAI222_X1 U17426 ( .A1(n19885), .A2(n14496), .B1(n13978), .B2(n19968), .C1(
        n19883), .C2(n19962), .ZN(P1_U2863) );
  INV_X1 U17427 ( .A(P1_EAX_REG_9__SCAN_IN), .ZN(n13980) );
  INV_X1 U17428 ( .A(DATAI_9_), .ZN(n13979) );
  MUX2_X1 U17429 ( .A(n13979), .B(n16388), .S(n14173), .Z(n20000) );
  OAI222_X1 U17430 ( .A1(n19885), .A2(n14566), .B1(n13980), .B2(n14529), .C1(
        n14155), .C2(n20000), .ZN(P1_U2895) );
  INV_X1 U17431 ( .A(n13983), .ZN(n13984) );
  XNOR2_X1 U17432 ( .A(n13982), .B(n13984), .ZN(n16181) );
  INV_X1 U17433 ( .A(n16180), .ZN(n18922) );
  INV_X1 U17434 ( .A(P2_INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n13985) );
  NAND3_X1 U17435 ( .A1(n13991), .A2(n13986), .A3(n13985), .ZN(n13988) );
  NAND2_X1 U17436 ( .A1(n19085), .A2(P2_REIP_REG_6__SCAN_IN), .ZN(n13987) );
  OAI211_X1 U17437 ( .C1(n18922), .C2(n16212), .A(n13988), .B(n13987), .ZN(
        n13989) );
  AOI21_X1 U17438 ( .B1(n16209), .B2(n13990), .A(n13989), .ZN(n13994) );
  NAND2_X1 U17439 ( .A1(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n13991), .ZN(
        n13992) );
  OAI211_X1 U17440 ( .C1(n14088), .C2(n13992), .A(
        P2_INSTADDRPOINTER_REG_6__SCAN_IN), .B(n15397), .ZN(n13993) );
  NAND2_X1 U17441 ( .A1(n13994), .A2(n13993), .ZN(n13995) );
  AOI21_X1 U17442 ( .B1(n16181), .B2(n16227), .A(n13995), .ZN(n13996) );
  OAI21_X1 U17443 ( .B1(n16179), .B2(n16223), .A(n13996), .ZN(P2_U3040) );
  NAND2_X1 U17444 ( .A1(n13791), .A2(n13997), .ZN(n14110) );
  OAI21_X1 U17445 ( .B1(n13999), .B2(n13998), .A(n14110), .ZN(n14076) );
  NAND2_X1 U17446 ( .A1(n15006), .A2(P2_EBX_REG_17__SCAN_IN), .ZN(n14003) );
  INV_X1 U17447 ( .A(n14114), .ZN(n14000) );
  AOI21_X1 U17448 ( .B1(n14001), .B2(n13965), .A(n14000), .ZN(n18824) );
  NAND2_X1 U17449 ( .A1(n18824), .A2(n14993), .ZN(n14002) );
  OAI211_X1 U17450 ( .C1(n14076), .C2(n15009), .A(n14003), .B(n14002), .ZN(
        P2_U2870) );
  XNOR2_X1 U17451 ( .A(n14688), .B(n15954), .ZN(n14004) );
  XNOR2_X1 U17452 ( .A(n14005), .B(n14004), .ZN(n14109) );
  INV_X1 U17453 ( .A(n14009), .ZN(n14007) );
  NAND2_X1 U17454 ( .A1(n14006), .A2(n20057), .ZN(n15992) );
  NOR2_X1 U17455 ( .A1(n14007), .A2(n15992), .ZN(n15955) );
  OAI211_X1 U17456 ( .C1(n20066), .C2(n14010), .A(n14009), .B(n14008), .ZN(
        n14012) );
  AOI21_X1 U17457 ( .B1(n20076), .B2(n14012), .A(n14011), .ZN(n15961) );
  NOR2_X1 U17458 ( .A1(n15961), .A2(n15954), .ZN(n14014) );
  NAND2_X1 U17459 ( .A1(n15986), .A2(P1_REIP_REG_9__SCAN_IN), .ZN(n14105) );
  OAI21_X1 U17460 ( .B1(n15975), .B2(n19883), .A(n14105), .ZN(n14013) );
  AOI211_X1 U17461 ( .C1(n15955), .C2(n15954), .A(n14014), .B(n14013), .ZN(
        n14015) );
  OAI21_X1 U17462 ( .B1(n14109), .B2(n20095), .A(n14015), .ZN(P1_U3022) );
  NOR2_X1 U17463 ( .A1(n18917), .A2(n18853), .ZN(n14016) );
  XNOR2_X1 U17464 ( .A(n14016), .B(n16138), .ZN(n14026) );
  INV_X1 U17465 ( .A(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n20975) );
  AOI22_X1 U17466 ( .A1(n14017), .A2(n18933), .B1(P2_EBX_REG_14__SCAN_IN), 
        .B2(n18951), .ZN(n14018) );
  OAI21_X1 U17467 ( .B1(n20975), .B2(n18831), .A(n14018), .ZN(n14025) );
  NAND2_X1 U17468 ( .A1(n16193), .A2(n18949), .ZN(n14022) );
  AOI21_X1 U17469 ( .B1(n14020), .B2(n14019), .A(n9851), .ZN(n18975) );
  AOI21_X1 U17470 ( .B1(n18877), .B2(n18975), .A(n19085), .ZN(n14021) );
  OAI211_X1 U17471 ( .C1(n18954), .C2(n14023), .A(n14022), .B(n14021), .ZN(
        n14024) );
  AOI211_X1 U17472 ( .C1(n14026), .C2(n18890), .A(n14025), .B(n14024), .ZN(
        n14027) );
  INV_X1 U17473 ( .A(n14027), .ZN(P2_U2841) );
  INV_X1 U17474 ( .A(n18957), .ZN(n14937) );
  INV_X1 U17475 ( .A(n19097), .ZN(n14031) );
  NOR2_X1 U17476 ( .A1(n18917), .A2(n14028), .ZN(n14030) );
  AOI21_X1 U17477 ( .B1(n14031), .B2(n14030), .A(n19714), .ZN(n14029) );
  OAI21_X1 U17478 ( .B1(n14031), .B2(n14030), .A(n14029), .ZN(n14041) );
  INV_X1 U17479 ( .A(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n14032) );
  OAI21_X1 U17480 ( .B1(n18831), .B2(n14032), .A(n18934), .ZN(n14035) );
  OAI22_X1 U17481 ( .A1(n18840), .A2(n14033), .B1(n12700), .B2(n18954), .ZN(
        n14034) );
  AOI211_X1 U17482 ( .C1(n18877), .C2(n14036), .A(n14035), .B(n14034), .ZN(
        n14037) );
  OAI21_X1 U17483 ( .B1(n14038), .B2(n18947), .A(n14037), .ZN(n14039) );
  AOI21_X1 U17484 ( .B1(n19089), .B2(n18949), .A(n14039), .ZN(n14040) );
  OAI211_X1 U17485 ( .C1(n14937), .C2(n18990), .A(n14041), .B(n14040), .ZN(
        P2_U2851) );
  INV_X1 U17486 ( .A(n14042), .ZN(n14055) );
  NOR2_X1 U17487 ( .A1(n18917), .A2(n14043), .ZN(n14044) );
  XNOR2_X1 U17488 ( .A(n14044), .B(n16178), .ZN(n14045) );
  NAND2_X1 U17489 ( .A1(n14045), .A2(n18890), .ZN(n14054) );
  AOI21_X1 U17490 ( .B1(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n18958), .A(
        n19085), .ZN(n14046) );
  OAI21_X1 U17491 ( .B1(n18937), .B2(n16211), .A(n14046), .ZN(n14052) );
  AOI21_X1 U17492 ( .B1(n14049), .B2(n14048), .A(n14047), .ZN(n16210) );
  INV_X1 U17493 ( .A(n16210), .ZN(n18987) );
  OAI22_X1 U17494 ( .A1(n14050), .A2(n18954), .B1(n18945), .B2(n18987), .ZN(
        n14051) );
  AOI211_X1 U17495 ( .C1(P2_EBX_REG_8__SCAN_IN), .C2(n18951), .A(n14052), .B(
        n14051), .ZN(n14053) );
  OAI211_X1 U17496 ( .C1(n18947), .C2(n14055), .A(n14054), .B(n14053), .ZN(
        P2_U2847) );
  OAI21_X1 U17497 ( .B1(n14057), .B2(n14056), .A(n14128), .ZN(n14411) );
  INV_X1 U17498 ( .A(P1_EBX_REG_10__SCAN_IN), .ZN(n14061) );
  INV_X1 U17499 ( .A(n14124), .ZN(n14059) );
  OAI21_X1 U17500 ( .B1(n13972), .B2(n14060), .A(n14059), .ZN(n14695) );
  OAI222_X1 U17501 ( .A1(n14411), .A2(n19962), .B1(n14061), .B2(n19968), .C1(
        n14695), .C2(n14496), .ZN(P1_U2862) );
  NAND2_X1 U17502 ( .A1(n14173), .A2(n14062), .ZN(n14063) );
  OAI21_X1 U17503 ( .B1(n14173), .B2(DATAI_10_), .A(n14063), .ZN(n20003) );
  INV_X1 U17504 ( .A(P1_EAX_REG_10__SCAN_IN), .ZN(n14064) );
  OAI222_X1 U17505 ( .A1(n14155), .A2(n20003), .B1(n14064), .B2(n14529), .C1(
        n14695), .C2(n14566), .ZN(P1_U2894) );
  NAND2_X1 U17506 ( .A1(n14066), .A2(n14067), .ZN(n14068) );
  NAND2_X1 U17507 ( .A1(n14065), .A2(n14068), .ZN(n15401) );
  INV_X1 U17508 ( .A(n15401), .ZN(n18823) );
  INV_X1 U17509 ( .A(P2_EAX_REG_17__SCAN_IN), .ZN(n19044) );
  OAI22_X1 U17510 ( .A1(n15084), .A2(n19119), .B1(n15083), .B2(n19044), .ZN(
        n14074) );
  NOR2_X2 U17511 ( .A1(n14071), .A2(n14069), .ZN(n18966) );
  INV_X1 U17512 ( .A(n18966), .ZN(n15088) );
  INV_X1 U17513 ( .A(BUF2_REG_17__SCAN_IN), .ZN(n14072) );
  NOR2_X2 U17514 ( .A1(n14071), .A2(n14070), .ZN(n18967) );
  INV_X1 U17515 ( .A(n18967), .ZN(n15086) );
  INV_X1 U17516 ( .A(BUF1_REG_17__SCAN_IN), .ZN(n14208) );
  OAI22_X1 U17517 ( .A1(n15088), .A2(n14072), .B1(n15086), .B2(n14208), .ZN(
        n14073) );
  AOI211_X1 U17518 ( .C1(n19005), .C2(n18823), .A(n14074), .B(n14073), .ZN(
        n14075) );
  OAI21_X1 U17519 ( .B1(n14076), .B2(n19009), .A(n14075), .ZN(P2_U2902) );
  XOR2_X1 U17520 ( .A(n10882), .B(n14078), .Z(n14079) );
  XNOR2_X1 U17521 ( .A(n14077), .B(n14079), .ZN(n14097) );
  NAND2_X1 U17522 ( .A1(n16164), .A2(n16166), .ZN(n14081) );
  XNOR2_X1 U17523 ( .A(n14080), .B(n14081), .ZN(n14095) );
  OAI22_X1 U17524 ( .A1(n19113), .A2(n14082), .B1(n10916), .B2(n18934), .ZN(
        n14085) );
  INV_X1 U17525 ( .A(n18906), .ZN(n14083) );
  OAI22_X1 U17526 ( .A1(n16174), .A2(n18910), .B1(n19098), .B2(n14083), .ZN(
        n14084) );
  AOI211_X1 U17527 ( .C1(n14095), .C2(n19087), .A(n14085), .B(n14084), .ZN(
        n14086) );
  OAI21_X1 U17528 ( .B1(n14097), .B2(n19092), .A(n14086), .ZN(P2_U3007) );
  OAI21_X1 U17529 ( .B1(n14088), .B2(n14087), .A(n15397), .ZN(n16206) );
  INV_X1 U17530 ( .A(n18910), .ZN(n14090) );
  NOR2_X1 U17531 ( .A1(n10916), .A2(n18934), .ZN(n14089) );
  AOI21_X1 U17532 ( .B1(n16219), .B2(n14090), .A(n14089), .ZN(n14091) );
  OAI21_X1 U17533 ( .B1(n18911), .B2(n16222), .A(n14091), .ZN(n14092) );
  AOI21_X1 U17534 ( .B1(n10882), .B2(n16203), .A(n14092), .ZN(n14093) );
  OAI21_X1 U17535 ( .B1(n10882), .B2(n16206), .A(n14093), .ZN(n14094) );
  AOI21_X1 U17536 ( .B1(n14095), .B2(n16227), .A(n14094), .ZN(n14096) );
  OAI21_X1 U17537 ( .B1(n14097), .B2(n16223), .A(n14096), .ZN(P2_U3039) );
  NOR2_X1 U17538 ( .A1(n9911), .A2(n14098), .ZN(n14099) );
  OR2_X1 U17539 ( .A1(n13235), .A2(n14099), .ZN(n18799) );
  AOI21_X1 U17540 ( .B1(n14102), .B2(n14100), .A(n14101), .ZN(n15081) );
  NAND2_X1 U17541 ( .A1(n15081), .A2(n14965), .ZN(n14104) );
  NAND2_X1 U17542 ( .A1(n15006), .A2(P2_EBX_REG_19__SCAN_IN), .ZN(n14103) );
  OAI211_X1 U17543 ( .C1(n18799), .C2(n15006), .A(n14104), .B(n14103), .ZN(
        P2_U2868) );
  OAI21_X1 U17544 ( .B1(n15915), .B2(n21011), .A(n14105), .ZN(n14107) );
  NOR2_X1 U17545 ( .A1(n19885), .A2(n20048), .ZN(n14106) );
  AOI211_X1 U17546 ( .C1(n15911), .C2(n19886), .A(n14107), .B(n14106), .ZN(
        n14108) );
  OAI21_X1 U17547 ( .B1(n19863), .B2(n14109), .A(n14108), .ZN(P1_U2990) );
  INV_X1 U17548 ( .A(n14110), .ZN(n14112) );
  OAI21_X1 U17549 ( .B1(n14112), .B2(n14111), .A(n14100), .ZN(n16119) );
  AND2_X1 U17550 ( .A1(n14114), .A2(n14113), .ZN(n14115) );
  OR2_X1 U17551 ( .A1(n14115), .A2(n9911), .ZN(n18811) );
  MUX2_X1 U17552 ( .A(n18811), .B(n14116), .S(n15006), .Z(n14117) );
  OAI21_X1 U17553 ( .B1(n16119), .B2(n15009), .A(n14117), .ZN(P2_U2869) );
  INV_X1 U17554 ( .A(n14101), .ZN(n14119) );
  AOI21_X1 U17555 ( .B1(n10252), .B2(n14119), .A(n9860), .ZN(n16114) );
  NAND2_X1 U17556 ( .A1(n16114), .A2(n14965), .ZN(n14121) );
  NAND2_X1 U17557 ( .A1(n15006), .A2(P2_EBX_REG_20__SCAN_IN), .ZN(n14120) );
  OAI211_X1 U17558 ( .C1(n15362), .C2(n15006), .A(n14121), .B(n14120), .ZN(
        P2_U2867) );
  OAI21_X1 U17559 ( .B1(n14124), .B2(n14123), .A(n14122), .ZN(n14133) );
  XNOR2_X1 U17560 ( .A(n14133), .B(n14131), .ZN(n15894) );
  INV_X1 U17561 ( .A(n15894), .ZN(n14130) );
  INV_X1 U17562 ( .A(P1_EAX_REG_11__SCAN_IN), .ZN(n14127) );
  INV_X1 U17563 ( .A(DATAI_11_), .ZN(n14126) );
  MUX2_X1 U17564 ( .A(n14126), .B(n14125), .S(n14173), .Z(n20005) );
  OAI222_X1 U17565 ( .A1(n14130), .A2(n14566), .B1(n14127), .B2(n14529), .C1(
        n14155), .C2(n20005), .ZN(P1_U2893) );
  INV_X1 U17566 ( .A(P1_EBX_REG_11__SCAN_IN), .ZN(n14129) );
  INV_X1 U17567 ( .A(n14128), .ZN(n14840) );
  XNOR2_X1 U17568 ( .A(n14840), .B(n14839), .ZN(n15844) );
  OAI222_X1 U17569 ( .A1(n14496), .A2(n14130), .B1(n14129), .B2(n19968), .C1(
        n19962), .C2(n15844), .ZN(P1_U2861) );
  INV_X1 U17570 ( .A(n14131), .ZN(n14132) );
  OAI21_X1 U17571 ( .B1(n14133), .B2(n14132), .A(n14122), .ZN(n14135) );
  NAND2_X1 U17572 ( .A1(n14135), .A2(n14134), .ZN(n14160) );
  OAI21_X1 U17573 ( .B1(n14135), .B2(n14134), .A(n14160), .ZN(n15838) );
  INV_X1 U17574 ( .A(P1_EAX_REG_12__SCAN_IN), .ZN(n14138) );
  INV_X1 U17575 ( .A(DATAI_12_), .ZN(n14137) );
  INV_X1 U17576 ( .A(BUF1_REG_12__SCAN_IN), .ZN(n14136) );
  MUX2_X1 U17577 ( .A(n14137), .B(n14136), .S(n14173), .Z(n20008) );
  OAI222_X1 U17578 ( .A1(n15838), .A2(n14566), .B1(n14138), .B2(n14529), .C1(
        n14155), .C2(n20008), .ZN(P1_U2892) );
  NAND2_X1 U17579 ( .A1(n14139), .A2(n14140), .ZN(n14149) );
  NAND2_X1 U17580 ( .A1(n14139), .A2(n14141), .ZN(n14157) );
  NAND2_X1 U17581 ( .A1(n14157), .A2(n14142), .ZN(n14143) );
  INV_X1 U17582 ( .A(DATAI_14_), .ZN(n14145) );
  NAND2_X1 U17583 ( .A1(n14173), .A2(BUF1_REG_14__SCAN_IN), .ZN(n14144) );
  OAI21_X1 U17584 ( .B1(n14173), .B2(n14145), .A(n14144), .ZN(n20014) );
  AOI22_X1 U17585 ( .A1(n14163), .A2(n20014), .B1(P1_EAX_REG_14__SCAN_IN), 
        .B2(n14558), .ZN(n14146) );
  OAI21_X1 U17586 ( .B1(n14184), .B2(n14566), .A(n14146), .ZN(P1_U2890) );
  INV_X1 U17587 ( .A(n14147), .ZN(n14148) );
  AOI21_X1 U17588 ( .B1(n14150), .B2(n14149), .A(n14148), .ZN(n14671) );
  INV_X1 U17589 ( .A(n14671), .ZN(n14409) );
  INV_X1 U17590 ( .A(P1_EBX_REG_15__SCAN_IN), .ZN(n14153) );
  OR2_X1 U17591 ( .A1(n14182), .A2(n14151), .ZN(n14152) );
  AND2_X1 U17592 ( .A1(n14168), .A2(n14152), .ZN(n14808) );
  INV_X1 U17593 ( .A(n14808), .ZN(n14404) );
  OAI222_X1 U17594 ( .A1(n14409), .A2(n14496), .B1(n19968), .B2(n14153), .C1(
        n14404), .C2(n19962), .ZN(P1_U2857) );
  OAI222_X1 U17595 ( .A1(n14409), .A2(n14566), .B1(n14529), .B2(n19971), .C1(
        n14155), .C2(n14154), .ZN(P1_U2889) );
  INV_X1 U17596 ( .A(n14156), .ZN(n14159) );
  INV_X1 U17597 ( .A(n14157), .ZN(n14158) );
  AOI21_X1 U17598 ( .B1(n14160), .B2(n14159), .A(n14158), .ZN(n14683) );
  INV_X1 U17599 ( .A(n14683), .ZN(n14204) );
  INV_X1 U17600 ( .A(DATAI_13_), .ZN(n14162) );
  NAND2_X1 U17601 ( .A1(n14173), .A2(BUF1_REG_13__SCAN_IN), .ZN(n14161) );
  OAI21_X1 U17602 ( .B1(n14173), .B2(n14162), .A(n14161), .ZN(n20010) );
  AOI22_X1 U17603 ( .A1(n14163), .A2(n20010), .B1(P1_EAX_REG_13__SCAN_IN), 
        .B2(n14558), .ZN(n14164) );
  OAI21_X1 U17604 ( .B1(n14204), .B2(n14566), .A(n14164), .ZN(P1_U2891) );
  AOI21_X1 U17605 ( .B1(n14166), .B2(n14147), .A(n14165), .ZN(n15876) );
  INV_X1 U17606 ( .A(n15876), .ZN(n14179) );
  INV_X1 U17607 ( .A(n14498), .ZN(n14167) );
  AOI21_X1 U17608 ( .B1(n14169), .B2(n14168), .A(n14167), .ZN(n15934) );
  AOI22_X1 U17609 ( .A1(n15934), .A2(n15856), .B1(P1_EBX_REG_16__SCAN_IN), 
        .B2(n14492), .ZN(n14170) );
  OAI21_X1 U17610 ( .B1(n14179), .B2(n14496), .A(n14170), .ZN(P1_U2856) );
  NAND2_X1 U17611 ( .A1(n14529), .A2(n14171), .ZN(n14172) );
  NOR2_X2 U17612 ( .A1(n14172), .A2(n14173), .ZN(n14564) );
  INV_X1 U17613 ( .A(n14172), .ZN(n14174) );
  NAND2_X1 U17614 ( .A1(n14174), .A2(n14173), .ZN(n14562) );
  INV_X1 U17615 ( .A(BUF1_REG_16__SCAN_IN), .ZN(n14176) );
  NOR3_X2 U17616 ( .A1(n14558), .A2(n14503), .A3(n11180), .ZN(n14559) );
  AOI22_X1 U17617 ( .A1(n14559), .A2(n20112), .B1(P1_EAX_REG_16__SCAN_IN), 
        .B2(n14558), .ZN(n14175) );
  OAI21_X1 U17618 ( .B1(n14562), .B2(n14176), .A(n14175), .ZN(n14177) );
  AOI21_X1 U17619 ( .B1(n14564), .B2(DATAI_16_), .A(n14177), .ZN(n14178) );
  OAI21_X1 U17620 ( .B1(n14179), .B2(n14566), .A(n14178), .ZN(P1_U2888) );
  INV_X1 U17621 ( .A(P1_EBX_REG_14__SCAN_IN), .ZN(n14183) );
  NOR2_X1 U17622 ( .A1(n14186), .A2(n14180), .ZN(n14181) );
  OR2_X1 U17623 ( .A1(n14182), .A2(n14181), .ZN(n15831) );
  OAI222_X1 U17624 ( .A1(n14184), .A2(n14496), .B1(n14183), .B2(n19968), .C1(
        n15831), .C2(n19962), .ZN(P1_U2858) );
  INV_X1 U17625 ( .A(n14496), .ZN(n19964) );
  AND2_X1 U17626 ( .A1(n14841), .A2(n14185), .ZN(n14187) );
  OR2_X1 U17627 ( .A1(n14187), .A2(n14186), .ZN(n14824) );
  OAI22_X1 U17628 ( .A1(n14824), .A2(n19962), .B1(n14188), .B2(n19968), .ZN(
        n14189) );
  AOI21_X1 U17629 ( .B1(n14683), .B2(n19964), .A(n14189), .ZN(n14190) );
  INV_X1 U17630 ( .A(n14190), .ZN(P1_U2859) );
  NAND2_X1 U17631 ( .A1(P1_REIP_REG_12__SCAN_IN), .A2(P1_REIP_REG_11__SCAN_IN), 
        .ZN(n15828) );
  NAND2_X1 U17632 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(P1_REIP_REG_9__SCAN_IN), 
        .ZN(n14196) );
  INV_X1 U17633 ( .A(n14191), .ZN(n14193) );
  AOI21_X1 U17634 ( .B1(n15781), .B2(n14192), .A(n15780), .ZN(n19931) );
  OAI21_X1 U17635 ( .B1(n14193), .B2(n19892), .A(n19931), .ZN(n19881) );
  AOI21_X1 U17636 ( .B1(n15781), .B2(n14196), .A(n19881), .ZN(n15846) );
  INV_X1 U17637 ( .A(n15846), .ZN(n14399) );
  AOI21_X1 U17638 ( .B1(n15828), .B2(n15781), .A(n14399), .ZN(n14194) );
  INV_X1 U17639 ( .A(n14194), .ZN(n15839) );
  INV_X1 U17640 ( .A(P1_REIP_REG_6__SCAN_IN), .ZN(n19891) );
  NAND3_X1 U17641 ( .A1(P1_REIP_REG_4__SCAN_IN), .A2(P1_REIP_REG_3__SCAN_IN), 
        .A3(P1_REIP_REG_2__SCAN_IN), .ZN(n14195) );
  NAND2_X1 U17642 ( .A1(n15781), .A2(P1_REIP_REG_1__SCAN_IN), .ZN(n19933) );
  NOR2_X1 U17643 ( .A1(n14195), .A2(n19933), .ZN(n19912) );
  NAND2_X1 U17644 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19912), .ZN(n19911) );
  NAND3_X1 U17645 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(P1_REIP_REG_7__SCAN_IN), 
        .A3(n19898), .ZN(n19890) );
  NOR2_X1 U17646 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n15828), .ZN(n14197) );
  AOI22_X1 U17647 ( .A1(P1_REIP_REG_13__SCAN_IN), .A2(n15839), .B1(n15849), 
        .B2(n14197), .ZN(n14203) );
  INV_X1 U17648 ( .A(n14681), .ZN(n14199) );
  AOI22_X1 U17649 ( .A1(n14199), .A2(n19941), .B1(n19955), .B2(
        P1_EBX_REG_13__SCAN_IN), .ZN(n14200) );
  OAI21_X1 U17650 ( .B1(n19937), .B2(n14824), .A(n14200), .ZN(n14201) );
  AOI211_X1 U17651 ( .C1(n19932), .C2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .A(
        n14201), .B(n15986), .ZN(n14202) );
  OAI211_X1 U17652 ( .C1(n14204), .C2(n15796), .A(n14203), .B(n14202), .ZN(
        P1_U2827) );
  OAI21_X1 U17653 ( .B1(n14165), .B2(n14206), .A(n14205), .ZN(n14660) );
  AOI22_X1 U17654 ( .A1(n14559), .A2(n20123), .B1(P1_EAX_REG_17__SCAN_IN), 
        .B2(n14558), .ZN(n14207) );
  OAI21_X1 U17655 ( .B1(n14562), .B2(n14208), .A(n14207), .ZN(n14209) );
  AOI21_X1 U17656 ( .B1(n14564), .B2(DATAI_17_), .A(n14209), .ZN(n14210) );
  OAI21_X1 U17657 ( .B1(n14660), .B2(n14566), .A(n14210), .ZN(P1_U2887) );
  OAI21_X1 U17658 ( .B1(n14212), .B2(P2_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n14211), .ZN(n15505) );
  NAND2_X1 U17659 ( .A1(n14214), .A2(n15479), .ZN(n14215) );
  XNOR2_X1 U17660 ( .A(n14213), .B(n14215), .ZN(n15502) );
  INV_X1 U17661 ( .A(n14216), .ZN(n14887) );
  OAI22_X1 U17662 ( .A1(n19113), .A2(n14217), .B1(n19098), .B2(n14887), .ZN(
        n14220) );
  OAI22_X1 U17663 ( .A1(n16174), .A2(n15498), .B1(n18934), .B2(n14218), .ZN(
        n14219) );
  AOI211_X1 U17664 ( .C1(n15502), .C2(n19087), .A(n14220), .B(n14219), .ZN(
        n14221) );
  OAI21_X1 U17665 ( .B1(n15505), .B2(n19092), .A(n14221), .ZN(P2_U3005) );
  INV_X1 U17666 ( .A(n18723), .ZN(n18757) );
  OAI21_X1 U17667 ( .B1(n18557), .B2(n11640), .A(n18539), .ZN(n14222) );
  NAND2_X1 U17668 ( .A1(n18558), .A2(n14222), .ZN(n18537) );
  NOR2_X1 U17669 ( .A1(n18757), .A2(n18537), .ZN(n14228) );
  NOR2_X1 U17670 ( .A1(n18615), .A2(n18530), .ZN(n14224) );
  NAND2_X1 U17671 ( .A1(n18100), .A2(n17312), .ZN(n18589) );
  AOI21_X1 U17672 ( .B1(n14224), .B2(n17259), .A(n14223), .ZN(n14226) );
  NAND2_X1 U17673 ( .A1(n14225), .A2(n18535), .ZN(n15634) );
  NAND3_X1 U17674 ( .A1(n14226), .A2(n15744), .A3(n15634), .ZN(n18565) );
  NOR2_X1 U17675 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(n18696), .ZN(n18093) );
  INV_X1 U17676 ( .A(P3_FLUSH_REG_SCAN_IN), .ZN(n18082) );
  NAND3_X1 U17677 ( .A1(P3_STATE2_REG_1__SCAN_IN), .A2(
        P3_STATE2_REG_0__SCAN_IN), .A3(P3_STATE2_REG_2__SCAN_IN), .ZN(n18694)
         );
  NOR2_X1 U17678 ( .A1(n18082), .A2(n18694), .ZN(n14227) );
  MUX2_X1 U17679 ( .A(n14228), .B(P3_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .S(
        n18728), .Z(P3_U3284) );
  OAI211_X1 U17680 ( .C1(n11640), .C2(n18557), .A(n15622), .B(n18539), .ZN(
        n18081) );
  NOR2_X1 U17681 ( .A1(P3_FLUSH_REG_SCAN_IN), .A2(n18081), .ZN(n14230) );
  INV_X1 U17682 ( .A(P3_STATE2_REG_1__SCAN_IN), .ZN(n18706) );
  AOI221_X1 U17683 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18706), .C1(n18603), 
        .C2(P3_STATE2_REG_1__SCAN_IN), .A(n18721), .ZN(n14229) );
  INV_X1 U17684 ( .A(n14229), .ZN(n18092) );
  OAI21_X1 U17685 ( .B1(n14230), .B2(n18694), .A(n18394), .ZN(n18087) );
  INV_X1 U17686 ( .A(n18087), .ZN(n14231) );
  OAI21_X1 U17687 ( .B1(n18706), .B2(n18603), .A(n18696), .ZN(n18740) );
  NOR2_X1 U17688 ( .A1(n18706), .A2(n18745), .ZN(n17721) );
  NOR2_X1 U17689 ( .A1(n18740), .A2(n17721), .ZN(n15656) );
  AOI21_X1 U17690 ( .B1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(
        P3_STATE2_REG_3__SCAN_IN), .A(n15656), .ZN(n15657) );
  NOR2_X1 U17691 ( .A1(n14231), .A2(n15657), .ZN(n14233) );
  NAND2_X1 U17692 ( .A1(n18696), .A2(n18603), .ZN(n16446) );
  NOR2_X1 U17693 ( .A1(n18745), .A2(n16446), .ZN(n16306) );
  NOR2_X1 U17694 ( .A1(n18696), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18140) );
  OR2_X1 U17695 ( .A1(n18140), .A2(n14231), .ZN(n15655) );
  OR2_X1 U17696 ( .A1(n16306), .A2(n15655), .ZN(n14232) );
  MUX2_X1 U17697 ( .A(n14233), .B(n14232), .S(
        P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .Z(P3_U2864) );
  NOR2_X1 U17698 ( .A1(n16028), .A2(n16212), .ZN(n14245) );
  NOR2_X1 U17699 ( .A1(n15025), .A2(n14234), .ZN(n14235) );
  INV_X1 U17700 ( .A(n16027), .ZN(n15018) );
  AOI21_X1 U17701 ( .B1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14239), .A(
        n15263), .ZN(n14236) );
  AOI211_X1 U17702 ( .C1(n14239), .C2(n15263), .A(n15258), .B(n14236), .ZN(
        n14238) );
  OR2_X1 U17703 ( .A1(n14238), .A2(n14237), .ZN(n14241) );
  NOR2_X1 U17704 ( .A1(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n15258), .ZN(
        n15269) );
  NOR2_X1 U17705 ( .A1(n15273), .A2(n15269), .ZN(n15264) );
  NOR2_X1 U17706 ( .A1(n15264), .A2(n14239), .ZN(n14240) );
  NAND2_X1 U17707 ( .A1(n14243), .A2(n14242), .ZN(n14244) );
  AOI211_X1 U17708 ( .C1(n14246), .C2(n12618), .A(n14245), .B(n14244), .ZN(
        n14247) );
  OAI21_X1 U17709 ( .B1(n14248), .B2(n16217), .A(n14247), .ZN(P2_U3017) );
  XNOR2_X1 U17710 ( .A(n14250), .B(P2_INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(
        n14251) );
  XNOR2_X1 U17711 ( .A(n13868), .B(n14251), .ZN(n16228) );
  NAND2_X1 U17712 ( .A1(n16228), .A2(n19087), .ZN(n14254) );
  NAND2_X1 U17713 ( .A1(n19101), .A2(n14900), .ZN(n14252) );
  NAND2_X1 U17714 ( .A1(n19085), .A2(P2_REIP_REG_3__SCAN_IN), .ZN(n16221) );
  OAI211_X1 U17715 ( .C1(n14901), .C2(n19113), .A(n14252), .B(n16221), .ZN(
        n14253) );
  OAI211_X1 U17716 ( .C1(n16224), .C2(n19092), .A(n14254), .B(n9931), .ZN(
        P2_U3011) );
  NAND2_X1 U17717 ( .A1(n20038), .A2(P1_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14255) );
  OAI211_X1 U17718 ( .C1(n15909), .C2(n14257), .A(n14256), .B(n14255), .ZN(
        n14258) );
  AOI21_X1 U17719 ( .B1(n14504), .B2(n20101), .A(n14258), .ZN(n14259) );
  OAI21_X1 U17720 ( .B1(n14260), .B2(n19863), .A(n14259), .ZN(P1_U2968) );
  INV_X1 U17721 ( .A(n14261), .ZN(n14264) );
  INV_X1 U17722 ( .A(n14262), .ZN(n14263) );
  NAND2_X1 U17723 ( .A1(n14264), .A2(n14263), .ZN(n14265) );
  AOI21_X1 U17724 ( .B1(n14268), .B2(n14267), .A(
        P2_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n14270) );
  OAI21_X1 U17725 ( .B1(n9883), .B2(n16223), .A(n14276), .ZN(n14277) );
  OAI21_X1 U17726 ( .B1(n14279), .B2(n16217), .A(n14278), .ZN(P2_U3016) );
  OAI22_X1 U17727 ( .A1(n14282), .A2(n14281), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n14280), .ZN(n15696) );
  OAI22_X1 U17728 ( .A1(n16000), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n20758), .ZN(n14283) );
  AOI21_X1 U17729 ( .B1(n15696), .B2(n14858), .A(n14283), .ZN(n14286) );
  AOI21_X1 U17730 ( .B1(n15697), .B2(n14858), .A(n14865), .ZN(n14285) );
  OAI22_X1 U17731 ( .A1(n14286), .A2(n14865), .B1(n14285), .B2(n14284), .ZN(
        P1_U3474) );
  NAND2_X1 U17732 ( .A1(n19086), .A2(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(
        n14287) );
  OAI211_X1 U17733 ( .C1(n14289), .C2(n19098), .A(n14288), .B(n14287), .ZN(
        n14290) );
  OAI21_X1 U17734 ( .B1(n14292), .B2(n19092), .A(n14291), .ZN(n14293) );
  INV_X1 U17735 ( .A(n14293), .ZN(n14294) );
  OAI21_X1 U17736 ( .B1(n14295), .B2(n19108), .A(n14294), .ZN(P2_U2983) );
  MUX2_X1 U17737 ( .A(n14688), .B(n14297), .S(n14296), .Z(n14298) );
  XNOR2_X1 U17738 ( .A(n14298), .B(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n14706) );
  INV_X1 U17739 ( .A(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n14299) );
  NAND2_X1 U17740 ( .A1(n15986), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14701) );
  OAI21_X1 U17741 ( .B1(n15915), .B2(n14299), .A(n14701), .ZN(n14303) );
  NOR2_X1 U17742 ( .A1(n14305), .A2(n20048), .ZN(n14302) );
  AOI211_X2 U17743 ( .C1(n14312), .C2(n15911), .A(n14303), .B(n14302), .ZN(
        n14304) );
  OAI21_X1 U17744 ( .B1(n14706), .B2(n19863), .A(n14304), .ZN(P1_U2970) );
  INV_X1 U17745 ( .A(BUF1_REG_29__SCAN_IN), .ZN(n14307) );
  AOI22_X1 U17746 ( .A1(n14559), .A2(n20010), .B1(P1_EAX_REG_29__SCAN_IN), 
        .B2(n14558), .ZN(n14306) );
  OAI21_X1 U17747 ( .B1(n14307), .B2(n14562), .A(n14306), .ZN(n14308) );
  AOI21_X1 U17748 ( .B1(n14564), .B2(DATAI_29_), .A(n14308), .ZN(n14309) );
  OAI21_X1 U17749 ( .B1(n14305), .B2(n14566), .A(n14309), .ZN(P1_U2875) );
  OAI21_X1 U17750 ( .B1(n14336), .B2(n14311), .A(n14310), .ZN(n14702) );
  INV_X1 U17751 ( .A(n14702), .ZN(n14317) );
  NOR2_X1 U17752 ( .A1(n14326), .A2(P1_REIP_REG_29__SCAN_IN), .ZN(n14316) );
  AOI22_X1 U17753 ( .A1(P1_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n19932), .B1(
        n19941), .B2(n14312), .ZN(n14314) );
  NAND2_X1 U17754 ( .A1(n19955), .A2(P1_EBX_REG_29__SCAN_IN), .ZN(n14313) );
  OAI211_X1 U17755 ( .C1(n14342), .C2(n14325), .A(n14314), .B(n14313), .ZN(
        n14315) );
  AOI211_X1 U17756 ( .C1(n14317), .C2(n19951), .A(n14316), .B(n14315), .ZN(
        n14318) );
  OAI21_X1 U17757 ( .B1(n14305), .B2(n15796), .A(n14318), .ZN(P1_U2811) );
  OAI222_X1 U17758 ( .A1(n14496), .A2(n14305), .B1(n14319), .B2(n19968), .C1(
        n14702), .C2(n19962), .ZN(P1_U2843) );
  NAND2_X1 U17759 ( .A1(n14572), .A2(n19908), .ZN(n14333) );
  OAI21_X1 U17760 ( .B1(n14326), .B2(n14325), .A(n14324), .ZN(n14331) );
  INV_X1 U17761 ( .A(P1_EBX_REG_30__SCAN_IN), .ZN(n14449) );
  NOR2_X1 U17762 ( .A1(n19934), .A2(n14449), .ZN(n14329) );
  INV_X1 U17763 ( .A(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n14327) );
  OAI22_X1 U17764 ( .A1(n14327), .A2(n19954), .B1(n19953), .B2(n14570), .ZN(
        n14328) );
  AOI211_X1 U17765 ( .C1(n14331), .C2(n14330), .A(n14329), .B(n14328), .ZN(
        n14332) );
  OAI211_X1 U17766 ( .C1(n14448), .C2(n19937), .A(n14333), .B(n14332), .ZN(
        P1_U2810) );
  AND2_X1 U17767 ( .A1(n9888), .A2(n14334), .ZN(n14335) );
  OR2_X1 U17768 ( .A1(n14336), .A2(n14335), .ZN(n14713) );
  AOI21_X1 U17769 ( .B1(n14339), .B2(n14337), .A(n14338), .ZN(n14586) );
  NAND2_X1 U17770 ( .A1(n14586), .A2(n19908), .ZN(n14348) );
  OAI22_X1 U17771 ( .A1(n14340), .A2(n19954), .B1(n19953), .B2(n14584), .ZN(
        n14346) );
  INV_X1 U17772 ( .A(n14341), .ZN(n14344) );
  INV_X1 U17773 ( .A(P1_REIP_REG_28__SCAN_IN), .ZN(n14343) );
  AOI21_X1 U17774 ( .B1(n14344), .B2(n14343), .A(n14342), .ZN(n14345) );
  AOI211_X1 U17775 ( .C1(n19955), .C2(P1_EBX_REG_28__SCAN_IN), .A(n14346), .B(
        n14345), .ZN(n14347) );
  OAI211_X1 U17776 ( .C1(n19937), .C2(n14713), .A(n14348), .B(n14347), .ZN(
        P1_U2812) );
  OAI21_X1 U17777 ( .B1(n14363), .B2(n14349), .A(n9888), .ZN(n14721) );
  INV_X1 U17778 ( .A(n14337), .ZN(n14351) );
  NAND2_X1 U17779 ( .A1(n14599), .A2(n19908), .ZN(n14358) );
  AND2_X1 U17780 ( .A1(n19952), .A2(n14353), .ZN(n14365) );
  INV_X1 U17781 ( .A(P1_EBX_REG_27__SCAN_IN), .ZN(n14451) );
  AOI22_X1 U17782 ( .A1(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n19932), .B1(
        n19941), .B2(n14594), .ZN(n14354) );
  OAI21_X1 U17783 ( .B1(n19934), .B2(n14451), .A(n14354), .ZN(n14356) );
  NOR3_X1 U17784 ( .A1(n14364), .A2(P1_REIP_REG_27__SCAN_IN), .A3(n15925), 
        .ZN(n14355) );
  AOI211_X1 U17785 ( .C1(P1_REIP_REG_27__SCAN_IN), .C2(n14365), .A(n14356), 
        .B(n14355), .ZN(n14357) );
  OAI211_X1 U17786 ( .C1(n19937), .C2(n14721), .A(n14358), .B(n14357), .ZN(
        P1_U2813) );
  AOI21_X1 U17787 ( .B1(n14360), .B2(n14456), .A(n14350), .ZN(n14609) );
  INV_X1 U17788 ( .A(n14609), .ZN(n14525) );
  NOR2_X1 U17789 ( .A1(n14458), .A2(n14361), .ZN(n14362) );
  OR2_X1 U17790 ( .A1(n14363), .A2(n14362), .ZN(n14452) );
  INV_X1 U17791 ( .A(n14452), .ZN(n15918) );
  INV_X1 U17792 ( .A(P1_EBX_REG_26__SCAN_IN), .ZN(n14453) );
  INV_X1 U17793 ( .A(n14364), .ZN(n14366) );
  OAI21_X1 U17794 ( .B1(n14366), .B2(P1_REIP_REG_26__SCAN_IN), .A(n14365), 
        .ZN(n14369) );
  INV_X1 U17795 ( .A(n14607), .ZN(n14367) );
  AOI22_X1 U17796 ( .A1(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n19932), .B1(
        n19941), .B2(n14367), .ZN(n14368) );
  OAI211_X1 U17797 ( .C1(n14453), .C2(n19934), .A(n14369), .B(n14368), .ZN(
        n14370) );
  AOI21_X1 U17798 ( .B1(n15918), .B2(n19951), .A(n14370), .ZN(n14371) );
  OAI21_X1 U17799 ( .B1(n14525), .B2(n15796), .A(n14371), .ZN(P1_U2814) );
  AOI21_X1 U17800 ( .B1(n14374), .B2(n9897), .A(n14373), .ZN(n14642) );
  INV_X1 U17801 ( .A(n14642), .ZN(n14557) );
  INV_X1 U17802 ( .A(n14375), .ZN(n14377) );
  INV_X1 U17803 ( .A(n19952), .ZN(n14376) );
  AOI21_X1 U17804 ( .B1(n14430), .B2(n14377), .A(n14376), .ZN(n15816) );
  INV_X1 U17805 ( .A(n14400), .ZN(n14378) );
  NAND2_X1 U17806 ( .A1(n14378), .A2(n15849), .ZN(n15827) );
  NOR3_X1 U17807 ( .A1(n14656), .A2(n15814), .A3(n15827), .ZN(n14397) );
  XOR2_X1 U17808 ( .A(n14379), .B(n20729), .Z(n14380) );
  AOI22_X1 U17809 ( .A1(P1_REIP_REG_19__SCAN_IN), .A2(n15816), .B1(n14397), 
        .B2(n14380), .ZN(n14387) );
  OR2_X1 U17810 ( .A1(n14390), .A2(n14381), .ZN(n14382) );
  NAND2_X1 U17811 ( .A1(n14759), .A2(n14382), .ZN(n14775) );
  INV_X1 U17812 ( .A(n14640), .ZN(n14383) );
  AOI22_X1 U17813 ( .A1(P1_EBX_REG_19__SCAN_IN), .A2(n19955), .B1(n14383), 
        .B2(n19941), .ZN(n14384) );
  OAI21_X1 U17814 ( .B1(n19937), .B2(n14775), .A(n14384), .ZN(n14385) );
  AOI211_X1 U17815 ( .C1(n19932), .C2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A(
        n14385), .B(n15986), .ZN(n14386) );
  OAI211_X1 U17816 ( .C1(n14557), .C2(n15796), .A(n14387), .B(n14386), .ZN(
        P1_U2821) );
  NAND2_X1 U17817 ( .A1(n14205), .A2(n14388), .ZN(n14389) );
  AND2_X1 U17818 ( .A1(n9897), .A2(n14389), .ZN(n14649) );
  INV_X1 U17819 ( .A(n14390), .ZN(n14391) );
  OAI21_X1 U17820 ( .B1(n14392), .B2(n14499), .A(n14391), .ZN(n14793) );
  AOI22_X1 U17821 ( .A1(n19955), .A2(P1_EBX_REG_18__SCAN_IN), .B1(
        P1_REIP_REG_18__SCAN_IN), .B2(n15816), .ZN(n14393) );
  OAI21_X1 U17822 ( .B1(n14647), .B2(n19953), .A(n14393), .ZN(n14394) );
  AOI211_X1 U17823 ( .C1(n19932), .C2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n14394), .B(n15986), .ZN(n14395) );
  OAI21_X1 U17824 ( .B1(n14793), .B2(n19937), .A(n14395), .ZN(n14396) );
  AOI21_X1 U17825 ( .B1(n14397), .B2(n20729), .A(n14396), .ZN(n14398) );
  OAI21_X1 U17826 ( .B1(n14567), .B2(n15796), .A(n14398), .ZN(P1_U2822) );
  NOR2_X1 U17827 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n15827), .ZN(n14407) );
  AOI21_X1 U17828 ( .B1(n14400), .B2(n19952), .A(n14399), .ZN(n15837) );
  INV_X1 U17829 ( .A(P1_REIP_REG_15__SCAN_IN), .ZN(n20726) );
  NOR2_X1 U17830 ( .A1(n15837), .A2(n20726), .ZN(n14406) );
  AOI21_X1 U17831 ( .B1(n19932), .B2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .A(
        n15986), .ZN(n14401) );
  OAI21_X1 U17832 ( .B1(n14669), .B2(n19953), .A(n14401), .ZN(n14402) );
  AOI21_X1 U17833 ( .B1(P1_EBX_REG_15__SCAN_IN), .B2(n19955), .A(n14402), .ZN(
        n14403) );
  OAI21_X1 U17834 ( .B1(n14404), .B2(n19937), .A(n14403), .ZN(n14405) );
  NOR3_X1 U17835 ( .A1(n14407), .A2(n14406), .A3(n14405), .ZN(n14408) );
  OAI21_X1 U17836 ( .B1(n14409), .B2(n15796), .A(n14408), .ZN(P1_U2825) );
  NOR2_X1 U17837 ( .A1(P1_REIP_REG_10__SCAN_IN), .A2(n19890), .ZN(n14415) );
  AOI21_X1 U17838 ( .B1(n19932), .B2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n15986), .ZN(n14410) );
  OAI21_X1 U17839 ( .B1(n14691), .B2(n19953), .A(n14410), .ZN(n14414) );
  INV_X1 U17840 ( .A(n14411), .ZN(n15952) );
  AOI22_X1 U17841 ( .A1(n19955), .A2(P1_EBX_REG_10__SCAN_IN), .B1(n19951), 
        .B2(n15952), .ZN(n14412) );
  OAI21_X1 U17842 ( .B1(n15846), .B2(n14690), .A(n14412), .ZN(n14413) );
  AOI211_X1 U17843 ( .C1(n14415), .C2(P1_REIP_REG_9__SCAN_IN), .A(n14414), .B(
        n14413), .ZN(n14416) );
  OAI21_X1 U17844 ( .B1(n14695), .B2(n15796), .A(n14416), .ZN(P1_U2830) );
  NOR2_X1 U17845 ( .A1(n19953), .A2(n14417), .ZN(n14418) );
  AOI211_X1 U17846 ( .C1(n19932), .C2(P1_PHYADDRPOINTER_REG_8__SCAN_IN), .A(
        n15986), .B(n14418), .ZN(n14420) );
  NAND2_X1 U17847 ( .A1(n19951), .A2(n15967), .ZN(n14419) );
  OAI211_X1 U17848 ( .C1(n14421), .C2(n19934), .A(n14420), .B(n14419), .ZN(
        n14422) );
  AOI21_X1 U17849 ( .B1(n19881), .B2(P1_REIP_REG_8__SCAN_IN), .A(n14422), .ZN(
        n14425) );
  INV_X1 U17850 ( .A(P1_REIP_REG_7__SCAN_IN), .ZN(n20717) );
  NOR2_X1 U17851 ( .A1(P1_REIP_REG_8__SCAN_IN), .A2(n20717), .ZN(n14423) );
  NAND2_X1 U17852 ( .A1(n19898), .A2(n14423), .ZN(n14424) );
  OAI211_X1 U17853 ( .C1(n14426), .C2(n15796), .A(n14425), .B(n14424), .ZN(
        P1_U2832) );
  OR2_X1 U17854 ( .A1(n20789), .A2(n14427), .ZN(n14428) );
  INV_X1 U17855 ( .A(n14429), .ZN(n20061) );
  OAI21_X1 U17856 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19892), .A(n14430), .ZN(
        n19945) );
  AOI22_X1 U17857 ( .A1(n19951), .A2(n20061), .B1(P1_REIP_REG_2__SCAN_IN), 
        .B2(n19945), .ZN(n14437) );
  INV_X1 U17858 ( .A(P1_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n21048) );
  OAI22_X1 U17859 ( .A1(n14431), .A2(n19953), .B1(n19954), .B2(n21048), .ZN(
        n14435) );
  NOR2_X1 U17860 ( .A1(n20789), .A2(n14432), .ZN(n19956) );
  INV_X1 U17861 ( .A(n19956), .ZN(n14433) );
  NOR2_X1 U17862 ( .A1(n14433), .A2(n13655), .ZN(n14434) );
  AOI211_X1 U17863 ( .C1(P1_EBX_REG_2__SCAN_IN), .C2(n19955), .A(n14435), .B(
        n14434), .ZN(n14436) );
  OAI211_X1 U17864 ( .C1(n19960), .C2(n14438), .A(n14437), .B(n14436), .ZN(
        n14439) );
  NOR2_X1 U17865 ( .A1(P1_REIP_REG_2__SCAN_IN), .A2(n19933), .ZN(n19946) );
  OR2_X1 U17866 ( .A1(n14439), .A2(n19946), .ZN(P1_U2838) );
  INV_X1 U17867 ( .A(n20380), .ZN(n20586) );
  NAND2_X1 U17868 ( .A1(n19956), .A2(n20586), .ZN(n14441) );
  AOI22_X1 U17869 ( .A1(n19932), .A2(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .B1(
        n15780), .B2(P1_REIP_REG_1__SCAN_IN), .ZN(n14440) );
  OAI211_X1 U17870 ( .C1(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n19953), .A(
        n14441), .B(n14440), .ZN(n14442) );
  AOI21_X1 U17871 ( .B1(n19951), .B2(n20080), .A(n14442), .ZN(n14444) );
  AOI22_X1 U17872 ( .A1(n19955), .A2(P1_EBX_REG_1__SCAN_IN), .B1(n15781), .B2(
        n20776), .ZN(n14443) );
  OAI211_X1 U17873 ( .C1(n19960), .C2(n14445), .A(n14444), .B(n14443), .ZN(
        P1_U2839) );
  OAI22_X1 U17874 ( .A1(n14447), .A2(n19962), .B1(n19968), .B2(n14446), .ZN(
        P1_U2841) );
  INV_X1 U17875 ( .A(n14572), .ZN(n14511) );
  INV_X1 U17876 ( .A(n14586), .ZN(n14516) );
  INV_X1 U17877 ( .A(P1_EBX_REG_28__SCAN_IN), .ZN(n14450) );
  OAI222_X1 U17878 ( .A1(n14496), .A2(n14516), .B1(n14450), .B2(n19968), .C1(
        n14713), .C2(n19962), .ZN(P1_U2844) );
  INV_X1 U17879 ( .A(n14599), .ZN(n14520) );
  OAI222_X1 U17880 ( .A1(n14496), .A2(n14520), .B1(n14451), .B2(n19968), .C1(
        n14721), .C2(n19962), .ZN(P1_U2845) );
  OAI222_X1 U17881 ( .A1(n14496), .A2(n14525), .B1(n14453), .B2(n19968), .C1(
        n14452), .C2(n19962), .ZN(P1_U2846) );
  OR2_X1 U17882 ( .A1(n14464), .A2(n14454), .ZN(n14455) );
  NAND2_X1 U17883 ( .A1(n14456), .A2(n14455), .ZN(n15756) );
  AND2_X1 U17884 ( .A1(n14468), .A2(n14457), .ZN(n14459) );
  OR2_X1 U17885 ( .A1(n14459), .A2(n14458), .ZN(n15760) );
  OAI22_X1 U17886 ( .A1(n15760), .A2(n19962), .B1(n15749), .B2(n19968), .ZN(
        n14460) );
  INV_X1 U17887 ( .A(n14460), .ZN(n14461) );
  OAI21_X1 U17888 ( .B1(n15756), .B2(n14496), .A(n14461), .ZN(P1_U2847) );
  INV_X1 U17889 ( .A(n14462), .ZN(n14465) );
  INV_X1 U17890 ( .A(n14463), .ZN(n14471) );
  AOI21_X1 U17891 ( .B1(n14465), .B2(n14471), .A(n14464), .ZN(n15766) );
  INV_X1 U17892 ( .A(n15766), .ZN(n14535) );
  INV_X1 U17893 ( .A(P1_EBX_REG_24__SCAN_IN), .ZN(n14469) );
  NAND2_X1 U17894 ( .A1(n14474), .A2(n14466), .ZN(n14467) );
  NAND2_X1 U17895 ( .A1(n14468), .A2(n14467), .ZN(n15764) );
  OAI222_X1 U17896 ( .A1(n14496), .A2(n14535), .B1(n14469), .B2(n19968), .C1(
        n15764), .C2(n19962), .ZN(P1_U2848) );
  INV_X1 U17897 ( .A(n14470), .ZN(n14481) );
  OR2_X1 U17898 ( .A1(n14484), .A2(n14472), .ZN(n14473) );
  NAND2_X1 U17899 ( .A1(n14474), .A2(n14473), .ZN(n15771) );
  OAI22_X1 U17900 ( .A1(n15771), .A2(n19962), .B1(n14475), .B2(n19968), .ZN(
        n14476) );
  INV_X1 U17901 ( .A(n14476), .ZN(n14477) );
  OAI21_X1 U17902 ( .B1(n15772), .B2(n14496), .A(n14477), .ZN(P1_U2849) );
  NAND2_X1 U17903 ( .A1(n14478), .A2(n14479), .ZN(n14480) );
  AND2_X1 U17904 ( .A1(n14481), .A2(n14480), .ZN(n15862) );
  INV_X1 U17905 ( .A(n15862), .ZN(n14543) );
  AND2_X1 U17906 ( .A1(n14491), .A2(n14482), .ZN(n14483) );
  NOR2_X1 U17907 ( .A1(n14484), .A2(n14483), .ZN(n15927) );
  AOI22_X1 U17908 ( .A1(n15927), .A2(n15856), .B1(P1_EBX_REG_22__SCAN_IN), 
        .B2(n14492), .ZN(n14485) );
  OAI21_X1 U17909 ( .B1(n14543), .B2(n14496), .A(n14485), .ZN(P1_U2850) );
  OAI21_X1 U17910 ( .B1(n14487), .B2(n14488), .A(n14478), .ZN(n15797) );
  NAND2_X1 U17911 ( .A1(n14761), .A2(n14489), .ZN(n14490) );
  NAND2_X1 U17912 ( .A1(n14491), .A2(n14490), .ZN(n15795) );
  INV_X1 U17913 ( .A(n15795), .ZN(n14493) );
  AOI22_X1 U17914 ( .A1(n14493), .A2(n15856), .B1(P1_EBX_REG_21__SCAN_IN), 
        .B2(n14492), .ZN(n14494) );
  OAI21_X1 U17915 ( .B1(n15797), .B2(n14496), .A(n14494), .ZN(P1_U2851) );
  INV_X1 U17916 ( .A(P1_EBX_REG_19__SCAN_IN), .ZN(n21014) );
  OAI222_X1 U17917 ( .A1(n14496), .A2(n14557), .B1(n19968), .B2(n21014), .C1(
        n14775), .C2(n19962), .ZN(P1_U2853) );
  INV_X1 U17918 ( .A(P1_EBX_REG_18__SCAN_IN), .ZN(n14495) );
  OAI222_X1 U17919 ( .A1(n14567), .A2(n14496), .B1(n14495), .B2(n19968), .C1(
        n14793), .C2(n19962), .ZN(P1_U2854) );
  INV_X1 U17920 ( .A(n14660), .ZN(n15817) );
  AND2_X1 U17921 ( .A1(n14498), .A2(n14497), .ZN(n14500) );
  OR2_X1 U17922 ( .A1(n14500), .A2(n14499), .ZN(n15820) );
  OAI22_X1 U17923 ( .A1(n15820), .A2(n19962), .B1(n15811), .B2(n19968), .ZN(
        n14501) );
  AOI21_X1 U17924 ( .B1(n15817), .B2(n19964), .A(n14501), .ZN(n14502) );
  INV_X1 U17925 ( .A(n14502), .ZN(P1_U2855) );
  INV_X1 U17926 ( .A(BUF1_REG_31__SCAN_IN), .ZN(n19147) );
  AOI22_X1 U17927 ( .A1(n14564), .A2(DATAI_31_), .B1(P1_EAX_REG_31__SCAN_IN), 
        .B2(n14558), .ZN(n14505) );
  OAI211_X1 U17928 ( .C1(n14562), .C2(n19147), .A(n14506), .B(n14505), .ZN(
        P1_U2873) );
  INV_X1 U17929 ( .A(BUF1_REG_30__SCAN_IN), .ZN(n14508) );
  AOI22_X1 U17930 ( .A1(n14559), .A2(n20014), .B1(P1_EAX_REG_30__SCAN_IN), 
        .B2(n14558), .ZN(n14507) );
  OAI21_X1 U17931 ( .B1(n14508), .B2(n14562), .A(n14507), .ZN(n14509) );
  AOI21_X1 U17932 ( .B1(n14564), .B2(DATAI_30_), .A(n14509), .ZN(n14510) );
  OAI21_X1 U17933 ( .B1(n14511), .B2(n14566), .A(n14510), .ZN(P1_U2874) );
  INV_X1 U17934 ( .A(n14562), .ZN(n14532) );
  INV_X1 U17935 ( .A(n14559), .ZN(n14530) );
  OAI22_X1 U17936 ( .A1(n14530), .A2(n20008), .B1(n14529), .B2(n14512), .ZN(
        n14513) );
  AOI21_X1 U17937 ( .B1(BUF1_REG_28__SCAN_IN), .B2(n14532), .A(n14513), .ZN(
        n14515) );
  NAND2_X1 U17938 ( .A1(n14564), .A2(DATAI_28_), .ZN(n14514) );
  OAI211_X1 U17939 ( .C1(n14516), .C2(n14566), .A(n14515), .B(n14514), .ZN(
        P1_U2876) );
  OAI22_X1 U17940 ( .A1(n14530), .A2(n20005), .B1(n14529), .B2(n20007), .ZN(
        n14517) );
  AOI21_X1 U17941 ( .B1(BUF1_REG_27__SCAN_IN), .B2(n14532), .A(n14517), .ZN(
        n14519) );
  NAND2_X1 U17942 ( .A1(n14564), .A2(DATAI_27_), .ZN(n14518) );
  OAI211_X1 U17943 ( .C1(n14520), .C2(n14566), .A(n14519), .B(n14518), .ZN(
        P1_U2877) );
  OAI22_X1 U17944 ( .A1(n14530), .A2(n20003), .B1(n14529), .B2(n14521), .ZN(
        n14522) );
  AOI21_X1 U17945 ( .B1(BUF1_REG_26__SCAN_IN), .B2(n14532), .A(n14522), .ZN(
        n14524) );
  NAND2_X1 U17946 ( .A1(n14564), .A2(DATAI_26_), .ZN(n14523) );
  OAI211_X1 U17947 ( .C1(n14525), .C2(n14566), .A(n14524), .B(n14523), .ZN(
        P1_U2878) );
  OAI22_X1 U17948 ( .A1(n14530), .A2(n20000), .B1(n14529), .B2(n20002), .ZN(
        n14526) );
  AOI21_X1 U17949 ( .B1(n14532), .B2(BUF1_REG_25__SCAN_IN), .A(n14526), .ZN(
        n14528) );
  NAND2_X1 U17950 ( .A1(n14564), .A2(DATAI_25_), .ZN(n14527) );
  OAI211_X1 U17951 ( .C1(n15756), .C2(n14566), .A(n14528), .B(n14527), .ZN(
        P1_U2879) );
  OAI22_X1 U17952 ( .A1(n14530), .A2(n19997), .B1(n14529), .B2(n19999), .ZN(
        n14531) );
  AOI21_X1 U17953 ( .B1(n14532), .B2(BUF1_REG_24__SCAN_IN), .A(n14531), .ZN(
        n14534) );
  NAND2_X1 U17954 ( .A1(n14564), .A2(DATAI_24_), .ZN(n14533) );
  OAI211_X1 U17955 ( .C1(n14535), .C2(n14566), .A(n14534), .B(n14533), .ZN(
        P1_U2880) );
  INV_X1 U17956 ( .A(BUF1_REG_23__SCAN_IN), .ZN(n15068) );
  AOI22_X1 U17957 ( .A1(n14559), .A2(n20148), .B1(P1_EAX_REG_23__SCAN_IN), 
        .B2(n14558), .ZN(n14536) );
  OAI21_X1 U17958 ( .B1(n14562), .B2(n15068), .A(n14536), .ZN(n14537) );
  AOI21_X1 U17959 ( .B1(n14564), .B2(DATAI_23_), .A(n14537), .ZN(n14538) );
  OAI21_X1 U17960 ( .B1(n15772), .B2(n14566), .A(n14538), .ZN(P1_U2881) );
  INV_X1 U17961 ( .A(BUF1_REG_22__SCAN_IN), .ZN(n14540) );
  AOI22_X1 U17962 ( .A1(n14559), .A2(n20139), .B1(P1_EAX_REG_22__SCAN_IN), 
        .B2(n14558), .ZN(n14539) );
  OAI21_X1 U17963 ( .B1(n14562), .B2(n14540), .A(n14539), .ZN(n14541) );
  AOI21_X1 U17964 ( .B1(n14564), .B2(DATAI_22_), .A(n14541), .ZN(n14542) );
  OAI21_X1 U17965 ( .B1(n14543), .B2(n14566), .A(n14542), .ZN(P1_U2882) );
  INV_X1 U17966 ( .A(BUF1_REG_21__SCAN_IN), .ZN(n15074) );
  AOI22_X1 U17967 ( .A1(n14559), .A2(n20136), .B1(P1_EAX_REG_21__SCAN_IN), 
        .B2(n14558), .ZN(n14544) );
  OAI21_X1 U17968 ( .B1(n14562), .B2(n15074), .A(n14544), .ZN(n14545) );
  AOI21_X1 U17969 ( .B1(n14564), .B2(DATAI_21_), .A(n14545), .ZN(n14546) );
  OAI21_X1 U17970 ( .B1(n15797), .B2(n14566), .A(n14546), .ZN(P1_U2883) );
  INV_X1 U17971 ( .A(n14547), .ZN(n14549) );
  INV_X1 U17972 ( .A(n14373), .ZN(n14548) );
  AOI21_X1 U17973 ( .B1(n14549), .B2(n14548), .A(n14487), .ZN(n15868) );
  INV_X1 U17974 ( .A(n15868), .ZN(n14553) );
  INV_X1 U17975 ( .A(BUF1_REG_20__SCAN_IN), .ZN(n16375) );
  AOI22_X1 U17976 ( .A1(n14559), .A2(n20133), .B1(P1_EAX_REG_20__SCAN_IN), 
        .B2(n14558), .ZN(n14550) );
  OAI21_X1 U17977 ( .B1(n16375), .B2(n14562), .A(n14550), .ZN(n14551) );
  AOI21_X1 U17978 ( .B1(n14564), .B2(DATAI_20_), .A(n14551), .ZN(n14552) );
  OAI21_X1 U17979 ( .B1(n14553), .B2(n14566), .A(n14552), .ZN(P1_U2884) );
  INV_X1 U17980 ( .A(BUF1_REG_19__SCAN_IN), .ZN(n15085) );
  AOI22_X1 U17981 ( .A1(n14559), .A2(n20130), .B1(P1_EAX_REG_19__SCAN_IN), 
        .B2(n14558), .ZN(n14554) );
  OAI21_X1 U17982 ( .B1(n14562), .B2(n15085), .A(n14554), .ZN(n14555) );
  AOI21_X1 U17983 ( .B1(n14564), .B2(DATAI_19_), .A(n14555), .ZN(n14556) );
  OAI21_X1 U17984 ( .B1(n14557), .B2(n14566), .A(n14556), .ZN(P1_U2885) );
  INV_X1 U17985 ( .A(BUF1_REG_18__SCAN_IN), .ZN(n14561) );
  AOI22_X1 U17986 ( .A1(n14559), .A2(n20126), .B1(P1_EAX_REG_18__SCAN_IN), 
        .B2(n14558), .ZN(n14560) );
  OAI21_X1 U17987 ( .B1(n14562), .B2(n14561), .A(n14560), .ZN(n14563) );
  AOI21_X1 U17988 ( .B1(n14564), .B2(DATAI_18_), .A(n14563), .ZN(n14565) );
  OAI21_X1 U17989 ( .B1(n14567), .B2(n14566), .A(n14565), .ZN(P1_U2886) );
  AOI21_X1 U17990 ( .B1(n20038), .B2(P1_PHYADDRPOINTER_REG_30__SCAN_IN), .A(
        n14568), .ZN(n14569) );
  OAI21_X1 U17991 ( .B1(n15909), .B2(n14570), .A(n14569), .ZN(n14571) );
  AOI21_X1 U17992 ( .B1(n14572), .B2(n20101), .A(n14571), .ZN(n14573) );
  OAI21_X1 U17993 ( .B1(n14574), .B2(n19863), .A(n14573), .ZN(P1_U2969) );
  INV_X1 U17994 ( .A(n14575), .ZN(n14617) );
  INV_X1 U17995 ( .A(n14578), .ZN(n14577) );
  INV_X1 U17996 ( .A(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n14604) );
  AND3_X1 U17997 ( .A1(n14604), .A2(n14727), .A3(n14718), .ZN(n14576) );
  NAND4_X1 U17998 ( .A1(n14577), .A2(n14576), .A3(n10173), .A4(n14739), .ZN(
        n14580) );
  MUX2_X1 U17999 ( .A(n14580), .B(n14579), .S(n11414), .Z(n14582) );
  XNOR2_X1 U18000 ( .A(n14582), .B(n14581), .ZN(n14716) );
  NAND2_X1 U18001 ( .A1(n15986), .A2(P1_REIP_REG_28__SCAN_IN), .ZN(n14712) );
  NAND2_X1 U18002 ( .A1(n20038), .A2(P1_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n14583) );
  OAI211_X1 U18003 ( .C1(n15909), .C2(n14584), .A(n14712), .B(n14583), .ZN(
        n14585) );
  AOI21_X1 U18004 ( .B1(n14586), .B2(n20101), .A(n14585), .ZN(n14587) );
  OAI21_X1 U18005 ( .B1(n19863), .B2(n14716), .A(n14587), .ZN(P1_U2971) );
  NOR2_X1 U18006 ( .A1(n14589), .A2(n14588), .ZN(n14592) );
  INV_X1 U18007 ( .A(n14590), .ZN(n14591) );
  MUX2_X1 U18008 ( .A(n14592), .B(n14591), .S(n14636), .Z(n14593) );
  XNOR2_X1 U18009 ( .A(n14593), .B(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n14725) );
  INV_X1 U18010 ( .A(n14594), .ZN(n14597) );
  NOR2_X1 U18011 ( .A1(n20046), .A2(n14595), .ZN(n14717) );
  AOI21_X1 U18012 ( .B1(n20038), .B2(P1_PHYADDRPOINTER_REG_27__SCAN_IN), .A(
        n14717), .ZN(n14596) );
  OAI21_X1 U18013 ( .B1(n15909), .B2(n14597), .A(n14596), .ZN(n14598) );
  AOI21_X1 U18014 ( .B1(n14599), .B2(n20101), .A(n14598), .ZN(n14600) );
  OAI21_X1 U18015 ( .B1(n19863), .B2(n14725), .A(n14600), .ZN(P1_U2972) );
  OAI21_X1 U18016 ( .B1(n14617), .B2(n14601), .A(n11414), .ZN(n14602) );
  NAND2_X1 U18017 ( .A1(n14603), .A2(n14602), .ZN(n14605) );
  XNOR2_X1 U18018 ( .A(n14605), .B(n14604), .ZN(n15917) );
  AOI22_X1 U18019 ( .A1(n20038), .A2(P1_PHYADDRPOINTER_REG_26__SCAN_IN), .B1(
        n15986), .B2(P1_REIP_REG_26__SCAN_IN), .ZN(n14606) );
  OAI21_X1 U18020 ( .B1(n15909), .B2(n14607), .A(n14606), .ZN(n14608) );
  AOI21_X1 U18021 ( .B1(n14609), .B2(n20101), .A(n14608), .ZN(n14610) );
  OAI21_X1 U18022 ( .B1(n19863), .B2(n15917), .A(n14610), .ZN(P1_U2973) );
  NAND2_X1 U18023 ( .A1(n10296), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14619) );
  MUX2_X1 U18024 ( .A(n14739), .B(n14611), .S(n14636), .Z(n14612) );
  AOI21_X1 U18025 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14619), .A(
        n14612), .ZN(n14613) );
  XNOR2_X1 U18026 ( .A(n14613), .B(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n14735) );
  NAND2_X1 U18027 ( .A1(n15986), .A2(P1_REIP_REG_25__SCAN_IN), .ZN(n14731) );
  OAI21_X1 U18028 ( .B1(n15915), .B2(n15748), .A(n14731), .ZN(n14615) );
  NOR2_X1 U18029 ( .A1(n15756), .A2(n20048), .ZN(n14614) );
  AOI211_X1 U18030 ( .C1(n15911), .C2(n15754), .A(n14615), .B(n14614), .ZN(
        n14616) );
  OAI21_X1 U18031 ( .B1(n19863), .B2(n14735), .A(n14616), .ZN(P1_U2974) );
  NAND2_X1 U18032 ( .A1(n14619), .A2(n14617), .ZN(n14618) );
  MUX2_X1 U18033 ( .A(n14619), .B(n14618), .S(n14636), .Z(n14620) );
  XNOR2_X1 U18034 ( .A(n14620), .B(n14739), .ZN(n14745) );
  OR2_X1 U18035 ( .A1(n20046), .A2(n20739), .ZN(n14741) );
  NAND2_X1 U18036 ( .A1(n20038), .A2(P1_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n14621) );
  OAI211_X1 U18037 ( .C1(n15909), .C2(n15769), .A(n14741), .B(n14621), .ZN(
        n14622) );
  AOI21_X1 U18038 ( .B1(n15766), .B2(n20101), .A(n14622), .ZN(n14623) );
  OAI21_X1 U18039 ( .B1(n19863), .B2(n14745), .A(n14623), .ZN(P1_U2975) );
  XNOR2_X1 U18040 ( .A(n14688), .B(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(
        n14624) );
  XNOR2_X1 U18041 ( .A(n14575), .B(n14624), .ZN(n14752) );
  INV_X1 U18042 ( .A(P1_PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n14626) );
  INV_X1 U18043 ( .A(P1_REIP_REG_23__SCAN_IN), .ZN(n14625) );
  OAI22_X1 U18044 ( .A1(n15915), .A2(n14626), .B1(n20046), .B2(n14625), .ZN(
        n14628) );
  NOR2_X1 U18045 ( .A1(n15772), .A2(n20048), .ZN(n14627) );
  AOI211_X1 U18046 ( .C1(n15911), .C2(n15774), .A(n14628), .B(n14627), .ZN(
        n14629) );
  OAI21_X1 U18047 ( .B1(n14752), .B2(n19863), .A(n14629), .ZN(P1_U2976) );
  INV_X1 U18048 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n14778) );
  NOR3_X1 U18049 ( .A1(n14644), .A2(n14636), .A3(n14778), .ZN(n14631) );
  NOR2_X1 U18050 ( .A1(n14631), .A2(n14630), .ZN(n14770) );
  NOR2_X1 U18051 ( .A1(n14770), .A2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(
        n14769) );
  AOI22_X1 U18052 ( .A1(n14769), .A2(n14636), .B1(
        P1_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n14631), .ZN(n14632) );
  XNOR2_X1 U18053 ( .A(n14632), .B(n11565), .ZN(n14757) );
  NAND2_X1 U18054 ( .A1(n15986), .A2(P1_REIP_REG_21__SCAN_IN), .ZN(n14754) );
  OAI21_X1 U18055 ( .B1(n15915), .B2(n15802), .A(n14754), .ZN(n14634) );
  NOR2_X1 U18056 ( .A1(n15797), .A2(n20048), .ZN(n14633) );
  AOI211_X1 U18057 ( .C1(n15911), .C2(n15799), .A(n14634), .B(n14633), .ZN(
        n14635) );
  OAI21_X1 U18058 ( .B1(n14757), .B2(n19863), .A(n14635), .ZN(P1_U2978) );
  XOR2_X1 U18059 ( .A(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B(n14638), .Z(
        n14783) );
  AOI22_X1 U18060 ( .A1(n20038), .A2(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B1(
        n15986), .B2(P1_REIP_REG_19__SCAN_IN), .ZN(n14639) );
  OAI21_X1 U18061 ( .B1(n15909), .B2(n14640), .A(n14639), .ZN(n14641) );
  AOI21_X1 U18062 ( .B1(n14642), .B2(n20101), .A(n14641), .ZN(n14643) );
  OAI21_X1 U18063 ( .B1(n14783), .B2(n19863), .A(n14643), .ZN(P1_U2980) );
  NAND2_X1 U18064 ( .A1(n15986), .A2(P1_REIP_REG_18__SCAN_IN), .ZN(n14792) );
  NAND2_X1 U18065 ( .A1(n20038), .A2(P1_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14646) );
  OAI211_X1 U18066 ( .C1(n15909), .C2(n14647), .A(n14792), .B(n14646), .ZN(
        n14648) );
  AOI21_X1 U18067 ( .B1(n14649), .B2(n20101), .A(n14648), .ZN(n14650) );
  OAI21_X1 U18068 ( .B1(n14797), .B2(n19863), .A(n14650), .ZN(P1_U2981) );
  NAND2_X1 U18069 ( .A1(n9901), .A2(n14651), .ZN(n14652) );
  XNOR2_X1 U18070 ( .A(n14652), .B(n14688), .ZN(n14654) );
  NAND2_X1 U18071 ( .A1(n14654), .A2(n14653), .ZN(n14655) );
  XOR2_X1 U18072 ( .A(n11550), .B(n14655), .Z(n14803) );
  NAND2_X1 U18073 ( .A1(n14803), .A2(n20043), .ZN(n14659) );
  INV_X1 U18074 ( .A(P1_REIP_REG_17__SCAN_IN), .ZN(n14656) );
  OR2_X1 U18075 ( .A1(n20046), .A2(n14656), .ZN(n14800) );
  OAI21_X1 U18076 ( .B1(n15915), .B2(n15810), .A(n14800), .ZN(n14657) );
  AOI21_X1 U18077 ( .B1(n15911), .B2(n15813), .A(n14657), .ZN(n14658) );
  OAI211_X1 U18078 ( .C1(n20048), .C2(n14660), .A(n14659), .B(n14658), .ZN(
        P1_U2982) );
  INV_X1 U18079 ( .A(n14661), .ZN(n15890) );
  NOR2_X1 U18080 ( .A1(n15890), .A2(n14662), .ZN(n14813) );
  NOR2_X1 U18081 ( .A1(n14813), .A2(n14663), .ZN(n15873) );
  INV_X1 U18082 ( .A(n15873), .ZN(n14664) );
  OAI21_X1 U18083 ( .B1(n14665), .B2(n14688), .A(n14664), .ZN(n14667) );
  XNOR2_X1 U18084 ( .A(n14688), .B(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n14666) );
  XNOR2_X1 U18085 ( .A(n14667), .B(n14666), .ZN(n14810) );
  AOI22_X1 U18086 ( .A1(n20038), .A2(P1_PHYADDRPOINTER_REG_15__SCAN_IN), .B1(
        n15986), .B2(P1_REIP_REG_15__SCAN_IN), .ZN(n14668) );
  OAI21_X1 U18087 ( .B1(n15909), .B2(n14669), .A(n14668), .ZN(n14670) );
  AOI21_X1 U18088 ( .B1(n14671), .B2(n20101), .A(n14670), .ZN(n14672) );
  OAI21_X1 U18089 ( .B1(n14810), .B2(n19863), .A(n14672), .ZN(P1_U2984) );
  NOR2_X1 U18090 ( .A1(n14661), .A2(n14673), .ZN(n14834) );
  INV_X1 U18091 ( .A(n14674), .ZN(n14833) );
  INV_X1 U18092 ( .A(n14677), .ZN(n14676) );
  NAND2_X1 U18093 ( .A1(n14676), .A2(n14675), .ZN(n14837) );
  NOR3_X1 U18094 ( .A1(n14834), .A2(n14833), .A3(n14837), .ZN(n14835) );
  NOR2_X1 U18095 ( .A1(n14835), .A2(n14677), .ZN(n14678) );
  XOR2_X1 U18096 ( .A(n14679), .B(n14678), .Z(n14832) );
  AOI22_X1 U18097 ( .A1(n20038), .A2(P1_PHYADDRPOINTER_REG_13__SCAN_IN), .B1(
        n15986), .B2(P1_REIP_REG_13__SCAN_IN), .ZN(n14680) );
  OAI21_X1 U18098 ( .B1(n15909), .B2(n14681), .A(n14680), .ZN(n14682) );
  AOI21_X1 U18099 ( .B1(n14683), .B2(n20101), .A(n14682), .ZN(n14684) );
  OAI21_X1 U18100 ( .B1(n14832), .B2(n19863), .A(n14684), .ZN(P1_U2986) );
  NAND2_X1 U18101 ( .A1(n14685), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14687) );
  XNOR2_X1 U18102 ( .A(n15890), .B(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n14686) );
  MUX2_X1 U18103 ( .A(n14687), .B(n14686), .S(n11414), .Z(n14689) );
  OR3_X1 U18104 ( .A1(n14685), .A2(P1_INSTADDRPOINTER_REG_10__SCAN_IN), .A3(
        n14688), .ZN(n15891) );
  NAND2_X1 U18105 ( .A1(n14689), .A2(n15891), .ZN(n15957) );
  NAND2_X1 U18106 ( .A1(n15957), .A2(n20043), .ZN(n14694) );
  INV_X1 U18107 ( .A(P1_REIP_REG_10__SCAN_IN), .ZN(n14690) );
  NOR2_X1 U18108 ( .A1(n20046), .A2(n14690), .ZN(n15951) );
  NOR2_X1 U18109 ( .A1(n15909), .A2(n14691), .ZN(n14692) );
  AOI211_X1 U18110 ( .C1(n20038), .C2(P1_PHYADDRPOINTER_REG_10__SCAN_IN), .A(
        n15951), .B(n14692), .ZN(n14693) );
  OAI211_X1 U18111 ( .C1(n20048), .C2(n14695), .A(n14694), .B(n14693), .ZN(
        P1_U2989) );
  INV_X1 U18112 ( .A(n14696), .ZN(n14704) );
  INV_X1 U18113 ( .A(n14697), .ZN(n14719) );
  NAND3_X1 U18114 ( .A1(n14719), .A2(n14699), .A3(n14698), .ZN(n14700) );
  OAI211_X1 U18115 ( .C1(n14702), .C2(n15975), .A(n14701), .B(n14700), .ZN(
        n14703) );
  AOI21_X1 U18116 ( .B1(P1_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n14704), .A(
        n14703), .ZN(n14705) );
  OAI21_X1 U18117 ( .B1(n14706), .B2(n20095), .A(n14705), .ZN(P1_U3002) );
  AND2_X1 U18118 ( .A1(n14708), .A2(n14707), .ZN(n14723) );
  NAND3_X1 U18119 ( .A1(n14719), .A2(n14710), .A3(n14709), .ZN(n14711) );
  OAI211_X1 U18120 ( .C1(n14713), .C2(n15975), .A(n14712), .B(n14711), .ZN(
        n14714) );
  AOI21_X1 U18121 ( .B1(P1_INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n14723), .A(
        n14714), .ZN(n14715) );
  OAI21_X1 U18122 ( .B1(n14716), .B2(n20095), .A(n14715), .ZN(P1_U3003) );
  AOI21_X1 U18123 ( .B1(n14719), .B2(n14718), .A(n14717), .ZN(n14720) );
  OAI21_X1 U18124 ( .B1(n14721), .B2(n15975), .A(n14720), .ZN(n14722) );
  AOI21_X1 U18125 ( .B1(P1_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n14723), .A(
        n14722), .ZN(n14724) );
  OAI21_X1 U18126 ( .B1(n14725), .B2(n20095), .A(n14724), .ZN(P1_U3004) );
  INV_X1 U18127 ( .A(n14726), .ZN(n14733) );
  AND2_X1 U18128 ( .A1(n14728), .A2(n14727), .ZN(n14729) );
  AND2_X1 U18129 ( .A1(n14750), .A2(n14729), .ZN(n15921) );
  INV_X1 U18130 ( .A(n15921), .ZN(n14730) );
  OAI211_X1 U18131 ( .C1(n15760), .C2(n15975), .A(n14731), .B(n14730), .ZN(
        n14732) );
  AOI21_X1 U18132 ( .B1(P1_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n14733), .A(
        n14732), .ZN(n14734) );
  OAI21_X1 U18133 ( .B1(n14735), .B2(n20095), .A(n14734), .ZN(P1_U3006) );
  INV_X1 U18134 ( .A(n20070), .ZN(n14738) );
  INV_X1 U18135 ( .A(n14736), .ZN(n14737) );
  OAI21_X1 U18136 ( .B1(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n14738), .A(
        n14737), .ZN(n14743) );
  NAND3_X1 U18137 ( .A1(n14750), .A2(P1_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n14739), .ZN(n14740) );
  OAI211_X1 U18138 ( .C1(n15764), .C2(n15975), .A(n14741), .B(n14740), .ZN(
        n14742) );
  AOI21_X1 U18139 ( .B1(P1_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n14743), .A(
        n14742), .ZN(n14744) );
  OAI21_X1 U18140 ( .B1(n14745), .B2(n20095), .A(n14744), .ZN(P1_U3007) );
  NOR2_X1 U18141 ( .A1(n14746), .A2(n10173), .ZN(n14749) );
  NAND2_X1 U18142 ( .A1(n15986), .A2(P1_REIP_REG_23__SCAN_IN), .ZN(n14747) );
  OAI21_X1 U18143 ( .B1(n15771), .B2(n15975), .A(n14747), .ZN(n14748) );
  AOI211_X1 U18144 ( .C1(n14750), .C2(n10173), .A(n14749), .B(n14748), .ZN(
        n14751) );
  OAI21_X1 U18145 ( .B1(n14752), .B2(n20095), .A(n14751), .ZN(P1_U3008) );
  NAND2_X1 U18146 ( .A1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n15926), .ZN(
        n14753) );
  OAI211_X1 U18147 ( .C1(n15795), .C2(n15975), .A(n14754), .B(n14753), .ZN(
        n14755) );
  AOI21_X1 U18148 ( .B1(n15930), .B2(n11565), .A(n14755), .ZN(n14756) );
  OAI21_X1 U18149 ( .B1(n14757), .B2(n20095), .A(n14756), .ZN(P1_U3010) );
  INV_X1 U18150 ( .A(n14777), .ZN(n14773) );
  NAND2_X1 U18151 ( .A1(n14759), .A2(n14758), .ZN(n14760) );
  NAND2_X1 U18152 ( .A1(n14761), .A2(n14760), .ZN(n15807) );
  INV_X1 U18153 ( .A(P1_REIP_REG_20__SCAN_IN), .ZN(n14762) );
  OR2_X1 U18154 ( .A1(n20046), .A2(n14762), .ZN(n14768) );
  INV_X1 U18155 ( .A(n14779), .ZN(n14766) );
  NOR2_X1 U18156 ( .A1(n14764), .A2(n14763), .ZN(n14765) );
  NAND2_X1 U18157 ( .A1(n14766), .A2(n14765), .ZN(n14767) );
  OAI211_X1 U18158 ( .C1(n15807), .C2(n15975), .A(n14768), .B(n14767), .ZN(
        n14772) );
  AOI21_X1 U18159 ( .B1(n14770), .B2(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n14769), .ZN(n15871) );
  NOR2_X1 U18160 ( .A1(n15871), .A2(n20095), .ZN(n14771) );
  AOI211_X1 U18161 ( .C1(P1_INSTADDRPOINTER_REG_20__SCAN_IN), .C2(n14773), .A(
        n14772), .B(n14771), .ZN(n14774) );
  INV_X1 U18162 ( .A(n14774), .ZN(P1_U3011) );
  INV_X1 U18163 ( .A(n14775), .ZN(n14781) );
  NAND2_X1 U18164 ( .A1(n15986), .A2(P1_REIP_REG_19__SCAN_IN), .ZN(n14776) );
  OAI221_X1 U18165 ( .B1(P1_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n14779), 
        .C1(n14778), .C2(n14777), .A(n14776), .ZN(n14780) );
  AOI21_X1 U18166 ( .B1(n14781), .B2(n20089), .A(n14780), .ZN(n14782) );
  OAI21_X1 U18167 ( .B1(n14783), .B2(n20095), .A(n14782), .ZN(P1_U3012) );
  NAND2_X1 U18168 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n14784), .ZN(
        n15939) );
  NOR2_X1 U18169 ( .A1(n15936), .A2(n15939), .ZN(n14799) );
  NOR2_X1 U18170 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n11550), .ZN(
        n14795) );
  OAI22_X1 U18171 ( .A1(n14820), .A2(n14786), .B1(n20066), .B2(n14785), .ZN(
        n14787) );
  NOR2_X1 U18172 ( .A1(n14788), .A2(n14787), .ZN(n14826) );
  OAI21_X1 U18173 ( .B1(n14790), .B2(n14789), .A(n14826), .ZN(n14798) );
  NAND2_X1 U18174 ( .A1(n14798), .A2(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(
        n14791) );
  OAI211_X1 U18175 ( .C1(n14793), .C2(n15975), .A(n14792), .B(n14791), .ZN(
        n14794) );
  AOI21_X1 U18176 ( .B1(n14799), .B2(n14795), .A(n14794), .ZN(n14796) );
  OAI21_X1 U18177 ( .B1(n14797), .B2(n20095), .A(n14796), .ZN(P1_U3013) );
  OAI21_X1 U18178 ( .B1(P1_INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n14799), .A(
        n14798), .ZN(n14801) );
  OAI211_X1 U18179 ( .C1(n15820), .C2(n15975), .A(n14801), .B(n14800), .ZN(
        n14802) );
  AOI21_X1 U18180 ( .B1(n14803), .B2(n20077), .A(n14802), .ZN(n14804) );
  INV_X1 U18181 ( .A(n14804), .ZN(P1_U3014) );
  INV_X1 U18182 ( .A(n14826), .ZN(n14818) );
  AOI21_X1 U18183 ( .B1(n11400), .B2(n20076), .A(n14818), .ZN(n15938) );
  NAND2_X1 U18184 ( .A1(n15986), .A2(P1_REIP_REG_15__SCAN_IN), .ZN(n14805) );
  OAI221_X1 U18185 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n15939), 
        .C1(n14806), .C2(n15938), .A(n14805), .ZN(n14807) );
  AOI21_X1 U18186 ( .B1(n14808), .B2(n20089), .A(n14807), .ZN(n14809) );
  OAI21_X1 U18187 ( .B1(n14810), .B2(n20095), .A(n14809), .ZN(P1_U3016) );
  OAI21_X1 U18188 ( .B1(n14813), .B2(n14812), .A(n14811), .ZN(n14815) );
  MUX2_X1 U18189 ( .A(n11400), .B(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .S(
        n11414), .Z(n14814) );
  XNOR2_X1 U18190 ( .A(n14815), .B(n14814), .ZN(n15884) );
  INV_X1 U18191 ( .A(P1_REIP_REG_14__SCAN_IN), .ZN(n14816) );
  OAI22_X1 U18192 ( .A1(n15831), .A2(n15975), .B1(n20046), .B2(n14816), .ZN(
        n14817) );
  AOI21_X1 U18193 ( .B1(n14818), .B2(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n14817), .ZN(n14823) );
  NOR2_X1 U18194 ( .A1(P1_INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n14819), .ZN(
        n14821) );
  NAND2_X1 U18195 ( .A1(n14821), .A2(n14820), .ZN(n14822) );
  OAI211_X1 U18196 ( .C1(n15884), .C2(n20095), .A(n14823), .B(n14822), .ZN(
        P1_U3017) );
  INV_X1 U18197 ( .A(n14824), .ZN(n14830) );
  NAND2_X1 U18198 ( .A1(n15986), .A2(P1_REIP_REG_13__SCAN_IN), .ZN(n14825) );
  OAI221_X1 U18199 ( .B1(P1_INSTADDRPOINTER_REG_13__SCAN_IN), .B2(n14828), 
        .C1(n14827), .C2(n14826), .A(n14825), .ZN(n14829) );
  AOI21_X1 U18200 ( .B1(n14830), .B2(n20089), .A(n14829), .ZN(n14831) );
  OAI21_X1 U18201 ( .B1(n14832), .B2(n20095), .A(n14831), .ZN(P1_U3018) );
  OR2_X1 U18202 ( .A1(n14834), .A2(n14833), .ZN(n14836) );
  AOI21_X1 U18203 ( .B1(n14837), .B2(n14836), .A(n14835), .ZN(n15889) );
  AOI21_X1 U18204 ( .B1(n14840), .B2(n14839), .A(n14838), .ZN(n14843) );
  INV_X1 U18205 ( .A(n14841), .ZN(n14842) );
  NOR2_X1 U18206 ( .A1(n14843), .A2(n14842), .ZN(n15855) );
  AOI22_X1 U18207 ( .A1(n15855), .A2(n20089), .B1(n15986), .B2(
        P1_REIP_REG_12__SCAN_IN), .ZN(n14854) );
  NAND2_X1 U18208 ( .A1(n15953), .A2(n15955), .ZN(n15950) );
  NOR2_X1 U18209 ( .A1(n14848), .A2(n15950), .ZN(n14851) );
  AOI22_X1 U18210 ( .A1(n20062), .A2(n14846), .B1(n14845), .B2(n14844), .ZN(
        n14847) );
  NAND2_X1 U18211 ( .A1(n20065), .A2(n14847), .ZN(n15946) );
  AOI21_X1 U18212 ( .B1(n20070), .B2(n14848), .A(n15946), .ZN(n14849) );
  INV_X1 U18213 ( .A(n14849), .ZN(n14850) );
  MUX2_X1 U18214 ( .A(n14851), .B(n14850), .S(
        P1_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(n14852) );
  INV_X1 U18215 ( .A(n14852), .ZN(n14853) );
  OAI211_X1 U18216 ( .C1(n15889), .C2(n20095), .A(n14854), .B(n14853), .ZN(
        P1_U3019) );
  XNOR2_X1 U18217 ( .A(n20378), .B(n20634), .ZN(n14856) );
  OAI22_X1 U18218 ( .A1(n14856), .A2(n20767), .B1(n13655), .B2(n14855), .ZN(
        n14857) );
  MUX2_X1 U18219 ( .A(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n14857), .S(
        n20773), .Z(P1_U3476) );
  INV_X1 U18220 ( .A(n14858), .ZN(n20759) );
  INV_X1 U18221 ( .A(n14859), .ZN(n14863) );
  INV_X1 U18222 ( .A(n14860), .ZN(n14861) );
  OAI222_X1 U18223 ( .A1(n14864), .A2(n20758), .B1(n20759), .B2(n14863), .C1(
        n14862), .C2(n14861), .ZN(n14866) );
  MUX2_X1 U18224 ( .A(n14866), .B(P1_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n14865), .Z(P1_U3472) );
  AOI21_X1 U18225 ( .B1(n15163), .B2(n14867), .A(n9908), .ZN(n15685) );
  INV_X1 U18226 ( .A(n14868), .ZN(n15684) );
  AOI21_X1 U18227 ( .B1(n18929), .B2(n15684), .A(n19714), .ZN(n14883) );
  INV_X1 U18228 ( .A(n15188), .ZN(n14879) );
  NAND2_X1 U18229 ( .A1(n14870), .A2(n14869), .ZN(n14871) );
  NAND2_X1 U18230 ( .A1(n15001), .A2(n14871), .ZN(n15164) );
  INV_X1 U18231 ( .A(n15164), .ZN(n15343) );
  OR2_X1 U18232 ( .A1(n13242), .A2(n14872), .ZN(n14875) );
  NAND2_X1 U18233 ( .A1(n14875), .A2(n14874), .ZN(n15346) );
  AOI22_X1 U18234 ( .A1(n18951), .A2(P2_EBX_REG_21__SCAN_IN), .B1(
        P2_REIP_REG_21__SCAN_IN), .B2(n18885), .ZN(n14876) );
  OAI21_X1 U18235 ( .B1(n18945), .B2(n15346), .A(n14876), .ZN(n14877) );
  AOI21_X1 U18236 ( .B1(n15343), .B2(n18949), .A(n14877), .ZN(n14878) );
  OAI21_X1 U18237 ( .B1(n14879), .B2(n18947), .A(n14878), .ZN(n14882) );
  OAI22_X1 U18238 ( .A1(n15685), .A2(n14880), .B1(n15163), .B2(n18831), .ZN(
        n14881) );
  AOI211_X1 U18239 ( .C1(n15685), .C2(n14883), .A(n14882), .B(n14881), .ZN(
        n14884) );
  INV_X1 U18240 ( .A(n14884), .ZN(P2_U2834) );
  NAND2_X1 U18241 ( .A1(n18929), .A2(n14885), .ZN(n14886) );
  XOR2_X1 U18242 ( .A(n14887), .B(n14886), .Z(n14896) );
  XNOR2_X1 U18243 ( .A(n14047), .B(n14888), .ZN(n18984) );
  OAI21_X1 U18244 ( .B1(n14218), .B2(n18954), .A(n18934), .ZN(n14889) );
  AOI21_X1 U18245 ( .B1(P2_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n18958), .A(
        n14889), .ZN(n14891) );
  NAND2_X1 U18246 ( .A1(n18951), .A2(P2_EBX_REG_9__SCAN_IN), .ZN(n14890) );
  OAI211_X1 U18247 ( .C1(n15498), .C2(n18937), .A(n14891), .B(n14890), .ZN(
        n14892) );
  AOI21_X1 U18248 ( .B1(n14893), .B2(n18933), .A(n14892), .ZN(n14894) );
  OAI21_X1 U18249 ( .B1(n18984), .B2(n18945), .A(n14894), .ZN(n14895) );
  AOI21_X1 U18250 ( .B1(n14896), .B2(n18890), .A(n14895), .ZN(n14897) );
  INV_X1 U18251 ( .A(n14897), .ZN(P2_U2846) );
  NAND2_X1 U18252 ( .A1(n18929), .A2(n14898), .ZN(n14899) );
  XNOR2_X1 U18253 ( .A(n14900), .B(n14899), .ZN(n14909) );
  NOR2_X1 U18254 ( .A1(n19788), .A2(n14937), .ZN(n14908) );
  OAI22_X1 U18255 ( .A1(n18840), .A2(n10656), .B1(n12690), .B2(n18954), .ZN(
        n14904) );
  OAI22_X1 U18256 ( .A1(n18947), .A2(n14902), .B1(n18831), .B2(n14901), .ZN(
        n14903) );
  OR2_X1 U18257 ( .A1(n14904), .A2(n14903), .ZN(n14905) );
  OAI21_X1 U18258 ( .B1(n18996), .B2(n18945), .A(n14906), .ZN(n14907) );
  AOI211_X1 U18259 ( .C1(n14909), .C2(n18890), .A(n14908), .B(n14907), .ZN(
        n14910) );
  INV_X1 U18260 ( .A(n14910), .ZN(P2_U2852) );
  INV_X1 U18261 ( .A(n14911), .ZN(n14913) );
  AOI22_X1 U18262 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(n18958), .B1(
        P2_REIP_REG_2__SCAN_IN), .B2(n18885), .ZN(n14912) );
  OAI21_X1 U18263 ( .B1(n18947), .B2(n14913), .A(n14912), .ZN(n14916) );
  NOR2_X1 U18264 ( .A1(n14914), .A2(n18937), .ZN(n14915) );
  AOI211_X1 U18265 ( .C1(P2_EBX_REG_2__SCAN_IN), .C2(n18951), .A(n14916), .B(
        n14915), .ZN(n14917) );
  OAI21_X1 U18266 ( .B1(n19799), .B2(n18945), .A(n14917), .ZN(n14922) );
  INV_X1 U18267 ( .A(n14920), .ZN(n19100) );
  NOR2_X1 U18268 ( .A1(n18917), .A2(n14918), .ZN(n14925) );
  INV_X1 U18269 ( .A(n14925), .ZN(n14919) );
  AOI221_X1 U18270 ( .B1(n19100), .B2(n14925), .C1(n14920), .C2(n14919), .A(
        n19714), .ZN(n14921) );
  AOI211_X1 U18271 ( .C1(n19804), .C2(n18957), .A(n14922), .B(n14921), .ZN(
        n14923) );
  INV_X1 U18272 ( .A(n14923), .ZN(P2_U2853) );
  INV_X1 U18273 ( .A(n14924), .ZN(n14926) );
  OAI21_X1 U18274 ( .B1(n14927), .B2(n14926), .A(n14925), .ZN(n15529) );
  OAI21_X1 U18275 ( .B1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n18929), .A(
        n15529), .ZN(n14928) );
  NAND2_X1 U18276 ( .A1(n14928), .A2(n18890), .ZN(n14936) );
  OAI22_X1 U18277 ( .A1(n18840), .A2(n14929), .B1(n19003), .B2(n18945), .ZN(
        n14932) );
  NOR2_X1 U18278 ( .A1(n18947), .A2(n14930), .ZN(n14931) );
  AOI211_X1 U18279 ( .C1(P2_PHYADDRPOINTER_REG_1__SCAN_IN), .C2(n18958), .A(
        n14932), .B(n14931), .ZN(n14933) );
  OAI21_X1 U18280 ( .B1(n10425), .B2(n18954), .A(n14933), .ZN(n14934) );
  AOI21_X1 U18281 ( .B1(n18949), .B2(n15536), .A(n14934), .ZN(n14935) );
  OAI211_X1 U18282 ( .C1(n14937), .C2(n19808), .A(n14936), .B(n14935), .ZN(
        P2_U2854) );
  MUX2_X1 U18283 ( .A(P2_EBX_REG_31__SCAN_IN), .B(n16013), .S(n14993), .Z(
        P2_U2856) );
  INV_X1 U18284 ( .A(n14938), .ZN(n15017) );
  NAND2_X1 U18285 ( .A1(n14940), .A2(n14939), .ZN(n15016) );
  NAND3_X1 U18286 ( .A1(n15017), .A2(n14965), .A3(n15016), .ZN(n14942) );
  NAND2_X1 U18287 ( .A1(n15006), .A2(P2_EBX_REG_29__SCAN_IN), .ZN(n14941) );
  OAI211_X1 U18288 ( .C1(n15006), .C2(n16028), .A(n14942), .B(n14941), .ZN(
        P2_U2858) );
  NAND2_X1 U18289 ( .A1(n14944), .A2(n14943), .ZN(n14946) );
  XNOR2_X1 U18290 ( .A(n14946), .B(n14945), .ZN(n15032) );
  NOR2_X1 U18291 ( .A1(n14947), .A2(n14948), .ZN(n14949) );
  OR2_X1 U18292 ( .A1(n14950), .A2(n14949), .ZN(n15100) );
  NOR2_X1 U18293 ( .A1(n15100), .A2(n15006), .ZN(n14951) );
  AOI21_X1 U18294 ( .B1(P2_EBX_REG_28__SCAN_IN), .B2(n15006), .A(n14951), .ZN(
        n14952) );
  OAI21_X1 U18295 ( .B1(n15032), .B2(n15009), .A(n14952), .ZN(P2_U2859) );
  NOR2_X1 U18296 ( .A1(n14960), .A2(n14953), .ZN(n14954) );
  AOI21_X1 U18297 ( .B1(n14956), .B2(n14955), .A(n9890), .ZN(n15041) );
  NAND2_X1 U18298 ( .A1(n15041), .A2(n14965), .ZN(n14958) );
  NAND2_X1 U18299 ( .A1(n15006), .A2(P2_EBX_REG_27__SCAN_IN), .ZN(n14957) );
  OAI211_X1 U18300 ( .C1(n15006), .C2(n16048), .A(n14958), .B(n14957), .ZN(
        P2_U2860) );
  AND2_X1 U18301 ( .A1(n14973), .A2(n14959), .ZN(n14961) );
  OR2_X1 U18302 ( .A1(n14961), .A2(n14960), .ZN(n15285) );
  AOI21_X1 U18303 ( .B1(n14964), .B2(n14963), .A(n14962), .ZN(n15050) );
  NAND2_X1 U18304 ( .A1(n15050), .A2(n14965), .ZN(n14967) );
  NAND2_X1 U18305 ( .A1(n15006), .A2(P2_EBX_REG_26__SCAN_IN), .ZN(n14966) );
  OAI211_X1 U18306 ( .C1(n15006), .C2(n15285), .A(n14967), .B(n14966), .ZN(
        P2_U2861) );
  OAI21_X1 U18307 ( .B1(n14970), .B2(n14969), .A(n14968), .ZN(n15057) );
  NAND2_X1 U18308 ( .A1(n14985), .A2(n14971), .ZN(n14972) );
  AND2_X1 U18309 ( .A1(n14973), .A2(n14972), .ZN(n16075) );
  NOR2_X1 U18310 ( .A1(n14993), .A2(n14974), .ZN(n14975) );
  AOI21_X1 U18311 ( .B1(n16075), .B2(n14993), .A(n14975), .ZN(n14976) );
  OAI21_X1 U18312 ( .B1(n15057), .B2(n15009), .A(n14976), .ZN(P2_U2862) );
  AOI21_X1 U18313 ( .B1(n14979), .B2(n14978), .A(n14977), .ZN(n14980) );
  XOR2_X1 U18314 ( .A(n14981), .B(n14980), .Z(n15065) );
  NAND2_X1 U18315 ( .A1(n14982), .A2(n14983), .ZN(n14984) );
  NAND2_X1 U18316 ( .A1(n14985), .A2(n14984), .ZN(n16085) );
  NOR2_X1 U18317 ( .A1(n16085), .A2(n15006), .ZN(n14986) );
  AOI21_X1 U18318 ( .B1(P2_EBX_REG_24__SCAN_IN), .B2(n15006), .A(n14986), .ZN(
        n14987) );
  OAI21_X1 U18319 ( .B1(n15065), .B2(n15009), .A(n14987), .ZN(P2_U2863) );
  AOI21_X1 U18320 ( .B1(n14990), .B2(n14989), .A(n14988), .ZN(n14991) );
  INV_X1 U18321 ( .A(n14991), .ZN(n15073) );
  INV_X1 U18322 ( .A(P2_EBX_REG_23__SCAN_IN), .ZN(n14994) );
  OAI21_X1 U18323 ( .B1(n9849), .B2(n14992), .A(n14982), .ZN(n16095) );
  MUX2_X1 U18324 ( .A(n14994), .B(n16095), .S(n14993), .Z(n14995) );
  OAI21_X1 U18325 ( .B1(n15073), .B2(n15009), .A(n14995), .ZN(P2_U2864) );
  AND2_X1 U18326 ( .A1(n14996), .A2(n14997), .ZN(n14999) );
  OR2_X1 U18327 ( .A1(n14999), .A2(n14998), .ZN(n16107) );
  AND2_X1 U18328 ( .A1(n15001), .A2(n15000), .ZN(n15002) );
  OR2_X1 U18329 ( .A1(n15002), .A2(n9849), .ZN(n15682) );
  INV_X1 U18330 ( .A(P2_EBX_REG_22__SCAN_IN), .ZN(n15003) );
  MUX2_X1 U18331 ( .A(n15682), .B(n15003), .S(n15006), .Z(n15004) );
  OAI21_X1 U18332 ( .B1(n16107), .B2(n15009), .A(n15004), .ZN(P2_U2865) );
  OAI21_X1 U18333 ( .B1(n9860), .B2(n15005), .A(n14996), .ZN(n15080) );
  MUX2_X1 U18334 ( .A(n15164), .B(n15007), .S(n15006), .Z(n15008) );
  OAI21_X1 U18335 ( .B1(n15080), .B2(n15009), .A(n15008), .ZN(P2_U2866) );
  AOI22_X1 U18336 ( .A1(n18966), .A2(BUF2_REG_30__SCAN_IN), .B1(n18967), .B2(
        BUF1_REG_30__SCAN_IN), .ZN(n15011) );
  AOI22_X1 U18337 ( .A1(n19005), .A2(n16017), .B1(P2_EAX_REG_30__SCAN_IN), 
        .B2(n19004), .ZN(n15010) );
  OAI211_X1 U18338 ( .C1(n15012), .C2(n15084), .A(n15011), .B(n15010), .ZN(
        n15013) );
  INV_X1 U18339 ( .A(n15013), .ZN(n15014) );
  OAI21_X1 U18340 ( .B1(n15015), .B2(n19009), .A(n15014), .ZN(P2_U2889) );
  NAND3_X1 U18341 ( .A1(n15017), .A2(n16121), .A3(n15016), .ZN(n15023) );
  AOI22_X1 U18342 ( .A1(n19005), .A2(n15018), .B1(n19004), .B2(
        P2_EAX_REG_29__SCAN_IN), .ZN(n15022) );
  AOI22_X1 U18343 ( .A1(n18966), .A2(BUF2_REG_29__SCAN_IN), .B1(n18967), .B2(
        BUF1_REG_29__SCAN_IN), .ZN(n15021) );
  INV_X1 U18344 ( .A(n15084), .ZN(n18965) );
  NAND2_X1 U18345 ( .A1(n18965), .A2(n15019), .ZN(n15020) );
  NAND4_X1 U18346 ( .A1(n15023), .A2(n15022), .A3(n15021), .A4(n15020), .ZN(
        P2_U2890) );
  AND2_X1 U18347 ( .A1(n9877), .A2(n15024), .ZN(n15026) );
  OR2_X1 U18348 ( .A1(n15026), .A2(n15025), .ZN(n16047) );
  INV_X1 U18349 ( .A(n16047), .ZN(n15261) );
  NAND2_X1 U18350 ( .A1(n19005), .A2(n15261), .ZN(n15027) );
  OAI21_X1 U18351 ( .B1(n15083), .B2(n19023), .A(n15027), .ZN(n15028) );
  AOI21_X1 U18352 ( .B1(n18965), .B2(n15029), .A(n15028), .ZN(n15031) );
  AOI22_X1 U18353 ( .A1(n18966), .A2(BUF2_REG_28__SCAN_IN), .B1(n18967), .B2(
        BUF1_REG_28__SCAN_IN), .ZN(n15030) );
  OAI211_X1 U18354 ( .C1(n15032), .C2(n19009), .A(n15031), .B(n15030), .ZN(
        P2_U2891) );
  AOI22_X1 U18355 ( .A1(n18966), .A2(BUF2_REG_27__SCAN_IN), .B1(n18967), .B2(
        BUF1_REG_27__SCAN_IN), .ZN(n15038) );
  NAND2_X1 U18356 ( .A1(n15033), .A2(n15034), .ZN(n15035) );
  NAND2_X1 U18357 ( .A1(n9877), .A2(n15035), .ZN(n16060) );
  INV_X1 U18358 ( .A(n16060), .ZN(n15036) );
  AOI22_X1 U18359 ( .A1(n19005), .A2(n15036), .B1(n19004), .B2(
        P2_EAX_REG_27__SCAN_IN), .ZN(n15037) );
  OAI211_X1 U18360 ( .C1(n15039), .C2(n15084), .A(n15038), .B(n15037), .ZN(
        n15040) );
  AOI21_X1 U18361 ( .B1(n15041), .B2(n16121), .A(n15040), .ZN(n15042) );
  INV_X1 U18362 ( .A(n15042), .ZN(P2_U2892) );
  AOI22_X1 U18363 ( .A1(n18966), .A2(BUF2_REG_26__SCAN_IN), .B1(n18967), .B2(
        BUF1_REG_26__SCAN_IN), .ZN(n15047) );
  OR2_X1 U18364 ( .A1(n15044), .A2(n15043), .ZN(n15045) );
  AND2_X1 U18365 ( .A1(n15033), .A2(n15045), .ZN(n16064) );
  AOI22_X1 U18366 ( .A1(n19005), .A2(n16064), .B1(n19004), .B2(
        P2_EAX_REG_26__SCAN_IN), .ZN(n15046) );
  OAI211_X1 U18367 ( .C1(n15048), .C2(n15084), .A(n15047), .B(n15046), .ZN(
        n15049) );
  AOI21_X1 U18368 ( .B1(n15050), .B2(n16121), .A(n15049), .ZN(n15051) );
  INV_X1 U18369 ( .A(n15051), .ZN(P2_U2893) );
  AOI22_X1 U18370 ( .A1(n18966), .A2(BUF2_REG_25__SCAN_IN), .B1(n18967), .B2(
        BUF1_REG_25__SCAN_IN), .ZN(n15053) );
  XNOR2_X1 U18371 ( .A(n15061), .B(n9934), .ZN(n16074) );
  AOI22_X1 U18372 ( .A1(n19005), .A2(n16074), .B1(n19004), .B2(
        P2_EAX_REG_25__SCAN_IN), .ZN(n15052) );
  OAI211_X1 U18373 ( .C1(n15054), .C2(n15084), .A(n15053), .B(n15052), .ZN(
        n15055) );
  INV_X1 U18374 ( .A(n15055), .ZN(n15056) );
  OAI21_X1 U18375 ( .B1(n15057), .B2(n19009), .A(n15056), .ZN(P2_U2894) );
  NAND2_X1 U18376 ( .A1(n15058), .A2(n15059), .ZN(n15060) );
  NAND2_X1 U18377 ( .A1(n15061), .A2(n15060), .ZN(n16084) );
  OAI22_X1 U18378 ( .A1(n18969), .A2(n16084), .B1(n15083), .B2(n19031), .ZN(
        n15062) );
  AOI21_X1 U18379 ( .B1(n18965), .B2(n18985), .A(n15062), .ZN(n15064) );
  AOI22_X1 U18380 ( .A1(n18966), .A2(BUF2_REG_24__SCAN_IN), .B1(n18967), .B2(
        BUF1_REG_24__SCAN_IN), .ZN(n15063) );
  OAI211_X1 U18381 ( .C1(n15065), .C2(n19009), .A(n15064), .B(n15063), .ZN(
        P2_U2895) );
  OR2_X1 U18382 ( .A1(n15332), .A2(n15066), .ZN(n15067) );
  AND2_X1 U18383 ( .A1(n15058), .A2(n15067), .ZN(n16096) );
  INV_X1 U18384 ( .A(P2_EAX_REG_23__SCAN_IN), .ZN(n21103) );
  OAI22_X1 U18385 ( .A1(n15084), .A2(n19150), .B1(n15083), .B2(n21103), .ZN(
        n15071) );
  INV_X1 U18386 ( .A(BUF2_REG_23__SCAN_IN), .ZN(n15069) );
  OAI22_X1 U18387 ( .A1(n15088), .A2(n15069), .B1(n15086), .B2(n15068), .ZN(
        n15070) );
  AOI211_X1 U18388 ( .C1(n19005), .C2(n16096), .A(n15071), .B(n15070), .ZN(
        n15072) );
  OAI21_X1 U18389 ( .B1(n15073), .B2(n19009), .A(n15072), .ZN(P2_U2896) );
  INV_X1 U18390 ( .A(n15346), .ZN(n15078) );
  INV_X1 U18391 ( .A(P2_EAX_REG_21__SCAN_IN), .ZN(n19036) );
  OAI22_X1 U18392 ( .A1(n15084), .A2(n19135), .B1(n15083), .B2(n19036), .ZN(
        n15077) );
  INV_X1 U18393 ( .A(BUF2_REG_21__SCAN_IN), .ZN(n15075) );
  OAI22_X1 U18394 ( .A1(n15088), .A2(n15075), .B1(n15086), .B2(n15074), .ZN(
        n15076) );
  AOI211_X1 U18395 ( .C1(n19005), .C2(n15078), .A(n15077), .B(n15076), .ZN(
        n15079) );
  OAI21_X1 U18396 ( .B1(n15080), .B2(n19009), .A(n15079), .ZN(P2_U2898) );
  INV_X1 U18397 ( .A(n15081), .ZN(n15092) );
  XNOR2_X1 U18398 ( .A(n15382), .B(n15082), .ZN(n18797) );
  INV_X1 U18399 ( .A(P2_EAX_REG_19__SCAN_IN), .ZN(n19040) );
  OAI22_X1 U18400 ( .A1(n15084), .A2(n19130), .B1(n15083), .B2(n19040), .ZN(
        n15090) );
  INV_X1 U18401 ( .A(BUF2_REG_19__SCAN_IN), .ZN(n15087) );
  OAI22_X1 U18402 ( .A1(n15088), .A2(n15087), .B1(n15086), .B2(n15085), .ZN(
        n15089) );
  AOI211_X1 U18403 ( .C1(n19005), .C2(n18797), .A(n15090), .B(n15089), .ZN(
        n15091) );
  OAI21_X1 U18404 ( .B1(n15092), .B2(n19009), .A(n15091), .ZN(P2_U2900) );
  XNOR2_X1 U18405 ( .A(n15095), .B(n15097), .ZN(n15109) );
  INV_X1 U18406 ( .A(n15095), .ZN(n15096) );
  XNOR2_X1 U18407 ( .A(n15098), .B(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15099) );
  AND2_X1 U18408 ( .A1(n15113), .A2(n15101), .ZN(n15103) );
  OR2_X1 U18409 ( .A1(n15103), .A2(n15102), .ZN(n16044) );
  NOR2_X1 U18410 ( .A1(n18934), .A2(n19768), .ZN(n15260) );
  AOI21_X1 U18411 ( .B1(n19086), .B2(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A(
        n15260), .ZN(n15104) );
  OAI21_X1 U18412 ( .B1(n16044), .B2(n19098), .A(n15104), .ZN(n15107) );
  NOR2_X1 U18413 ( .A1(n15265), .A2(n19092), .ZN(n15106) );
  AOI211_X2 U18414 ( .C1(n16041), .C2(n19104), .A(n15107), .B(n15106), .ZN(
        n15108) );
  XNOR2_X1 U18415 ( .A(n15109), .B(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(
        n15278) );
  AOI21_X1 U18417 ( .B1(n21005), .B2(n15111), .A(n15112), .ZN(n15276) );
  INV_X1 U18418 ( .A(n15113), .ZN(n15114) );
  AOI21_X1 U18419 ( .B1(n16049), .B2(n15126), .A(n15114), .ZN(n16003) );
  NAND2_X1 U18420 ( .A1(n19085), .A2(P2_REIP_REG_27__SCAN_IN), .ZN(n15270) );
  OAI21_X1 U18421 ( .B1(n19113), .B2(n16049), .A(n15270), .ZN(n15115) );
  AOI21_X1 U18422 ( .B1(n16003), .B2(n19101), .A(n15115), .ZN(n15116) );
  OAI21_X1 U18423 ( .B1(n16048), .B2(n16174), .A(n15116), .ZN(n15117) );
  AOI21_X1 U18424 ( .B1(n15276), .B2(n19102), .A(n15117), .ZN(n15118) );
  OAI21_X1 U18425 ( .B1(n15278), .B2(n19108), .A(n15118), .ZN(P2_U2987) );
  NAND2_X1 U18426 ( .A1(n15119), .A2(n15120), .ZN(n15121) );
  NAND2_X1 U18427 ( .A1(n15111), .A2(n15121), .ZN(n15290) );
  NAND2_X1 U18428 ( .A1(n15122), .A2(n15131), .ZN(n15124) );
  XNOR2_X1 U18429 ( .A(n15124), .B(n15123), .ZN(n15279) );
  NAND2_X1 U18430 ( .A1(n15279), .A2(n19087), .ZN(n15130) );
  INV_X1 U18431 ( .A(n15285), .ZN(n16065) );
  OR2_X1 U18432 ( .A1(n15136), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15125) );
  NAND2_X1 U18433 ( .A1(n15126), .A2(n15125), .ZN(n16068) );
  NAND2_X1 U18434 ( .A1(n19085), .A2(P2_REIP_REG_26__SCAN_IN), .ZN(n15282) );
  NAND2_X1 U18435 ( .A1(n19086), .A2(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(
        n15127) );
  OAI211_X1 U18436 ( .C1(n16068), .C2(n19098), .A(n15282), .B(n15127), .ZN(
        n15128) );
  AOI21_X1 U18437 ( .B1(n16065), .B2(n19104), .A(n15128), .ZN(n15129) );
  OAI211_X1 U18438 ( .C1(n19092), .C2(n15290), .A(n15130), .B(n15129), .ZN(
        P2_U2988) );
  INV_X1 U18439 ( .A(n15131), .ZN(n15134) );
  AND2_X1 U18440 ( .A1(n15132), .A2(n15131), .ZN(n15133) );
  OAI22_X1 U18441 ( .A1(n15122), .A2(n15134), .B1(n9898), .B2(n15133), .ZN(
        n15300) );
  AND2_X1 U18442 ( .A1(n15146), .A2(n15138), .ZN(n15135) );
  NOR2_X1 U18443 ( .A1(n15136), .A2(n15135), .ZN(n16004) );
  NAND2_X1 U18444 ( .A1(n16004), .A2(n19101), .ZN(n15137) );
  NAND2_X1 U18445 ( .A1(n19085), .A2(P2_REIP_REG_25__SCAN_IN), .ZN(n15291) );
  OAI211_X1 U18446 ( .C1(n19113), .C2(n15138), .A(n15137), .B(n15291), .ZN(
        n15139) );
  AOI21_X1 U18447 ( .B1(n16075), .B2(n19104), .A(n15139), .ZN(n15142) );
  OR2_X1 U18448 ( .A1(n15140), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15297) );
  NAND3_X1 U18449 ( .A1(n15297), .A2(n15119), .A3(n19102), .ZN(n15141) );
  OAI211_X1 U18450 ( .C1(n15300), .C2(n19108), .A(n15142), .B(n15141), .ZN(
        P2_U2989) );
  XNOR2_X1 U18451 ( .A(n15144), .B(n15301), .ZN(n15145) );
  XNOR2_X1 U18452 ( .A(n15143), .B(n15145), .ZN(n15311) );
  AOI21_X1 U18453 ( .B1(n15301), .B2(n9850), .A(n15140), .ZN(n15309) );
  NOR2_X1 U18454 ( .A1(n16085), .A2(n16174), .ZN(n15149) );
  OAI21_X1 U18455 ( .B1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n15151), .A(
        n15146), .ZN(n16089) );
  NAND2_X1 U18456 ( .A1(n19085), .A2(P2_REIP_REG_24__SCAN_IN), .ZN(n15303) );
  NAND2_X1 U18457 ( .A1(n19086), .A2(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(
        n15147) );
  OAI211_X1 U18458 ( .C1(n16089), .C2(n19098), .A(n15303), .B(n15147), .ZN(
        n15148) );
  AOI211_X1 U18459 ( .C1(n15309), .C2(n19102), .A(n15149), .B(n15148), .ZN(
        n15150) );
  OAI21_X1 U18460 ( .B1(n15311), .B2(n19108), .A(n15150), .ZN(P2_U2990) );
  NAND2_X1 U18461 ( .A1(n15160), .A2(n15312), .ZN(n15324) );
  NOR2_X1 U18462 ( .A1(n15324), .A2(n15338), .ZN(n15323) );
  OAI21_X1 U18463 ( .B1(n15323), .B2(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        n9850), .ZN(n15322) );
  AOI21_X1 U18464 ( .B1(n15152), .B2(n15686), .A(n15151), .ZN(n16005) );
  OAI22_X1 U18465 ( .A1(n19113), .A2(n15152), .B1(n10960), .B2(n18934), .ZN(
        n15154) );
  NOR2_X1 U18466 ( .A1(n16095), .A2(n16174), .ZN(n15153) );
  AOI211_X1 U18467 ( .C1(n16005), .C2(n19101), .A(n15154), .B(n15153), .ZN(
        n15159) );
  INV_X1 U18468 ( .A(n15155), .ZN(n15319) );
  NAND2_X1 U18469 ( .A1(n15157), .A2(n15156), .ZN(n15318) );
  NAND3_X1 U18470 ( .A1(n15319), .A2(n19087), .A3(n15318), .ZN(n15158) );
  OAI211_X1 U18471 ( .C1(n15322), .C2(n19092), .A(n15159), .B(n15158), .ZN(
        P2_U2991) );
  NAND2_X2 U18472 ( .A1(n15247), .A2(n15161), .ZN(n15394) );
  NOR2_X2 U18473 ( .A1(n15394), .A2(n15162), .ZN(n15210) );
  NOR2_X2 U18474 ( .A1(n15195), .A2(n15357), .ZN(n15196) );
  OAI21_X1 U18475 ( .B1(n15196), .B2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A(
        n15324), .ZN(n15354) );
  NAND2_X1 U18476 ( .A1(n19085), .A2(P2_REIP_REG_21__SCAN_IN), .ZN(n15344) );
  OAI21_X1 U18477 ( .B1(n19113), .B2(n15163), .A(n15344), .ZN(n15166) );
  NOR2_X1 U18478 ( .A1(n15164), .A2(n16174), .ZN(n15165) );
  AOI211_X1 U18479 ( .C1(n19101), .C2(n15685), .A(n15166), .B(n15165), .ZN(
        n15194) );
  INV_X1 U18480 ( .A(n15168), .ZN(n15453) );
  NAND2_X1 U18481 ( .A1(n15452), .A2(n15169), .ZN(n15436) );
  AND2_X1 U18482 ( .A1(n15187), .A2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(
        n15170) );
  NAND2_X1 U18483 ( .A1(n18855), .A2(n15170), .ZN(n15434) );
  AND2_X1 U18484 ( .A1(n15172), .A2(n15434), .ZN(n15171) );
  NAND2_X1 U18485 ( .A1(n15436), .A2(n15171), .ZN(n15437) );
  NAND2_X1 U18486 ( .A1(n15437), .A2(n15172), .ZN(n16134) );
  INV_X1 U18487 ( .A(n16134), .ZN(n15173) );
  OR2_X1 U18488 ( .A1(n15174), .A2(n16196), .ZN(n16133) );
  NOR2_X1 U18489 ( .A1(n15177), .A2(n15176), .ZN(n15249) );
  INV_X1 U18490 ( .A(n15238), .ZN(n15178) );
  NAND2_X1 U18491 ( .A1(n15222), .A2(n15206), .ZN(n15183) );
  AND2_X1 U18492 ( .A1(n15220), .A2(n15207), .ZN(n15184) );
  NAND2_X1 U18493 ( .A1(n15186), .A2(n15185), .ZN(n15202) );
  NAND2_X1 U18494 ( .A1(n15366), .A2(n15186), .ZN(n15192) );
  NAND2_X1 U18495 ( .A1(n15188), .A2(n15187), .ZN(n15190) );
  XNOR2_X1 U18496 ( .A(n15190), .B(n15189), .ZN(n15191) );
  NAND2_X1 U18497 ( .A1(n15351), .A2(n19087), .ZN(n15193) );
  OAI211_X1 U18498 ( .C1(n15354), .C2(n19092), .A(n15194), .B(n15193), .ZN(
        P2_U2993) );
  INV_X1 U18499 ( .A(n15196), .ZN(n15197) );
  OAI21_X1 U18500 ( .B1(P2_INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n15211), .A(
        n15197), .ZN(n15369) );
  INV_X1 U18501 ( .A(n15362), .ZN(n15201) );
  NOR2_X1 U18502 ( .A1(n18934), .A2(n19756), .ZN(n15359) );
  AOI21_X1 U18503 ( .B1(n19086), .B2(P2_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n15359), .ZN(n15198) );
  OAI21_X1 U18504 ( .B1(n19098), .B2(n15199), .A(n15198), .ZN(n15200) );
  AOI21_X1 U18505 ( .B1(n15201), .B2(n19104), .A(n15200), .ZN(n15205) );
  NAND2_X1 U18506 ( .A1(n15203), .A2(n15202), .ZN(n15365) );
  NAND3_X1 U18507 ( .A1(n15366), .A2(n19087), .A3(n15365), .ZN(n15204) );
  OAI211_X1 U18508 ( .C1(n15369), .C2(n19092), .A(n15205), .B(n15204), .ZN(
        P2_U2994) );
  NAND2_X1 U18509 ( .A1(n15207), .A2(n15206), .ZN(n15209) );
  NAND2_X1 U18510 ( .A1(n15219), .A2(n15220), .ZN(n15218) );
  NAND2_X1 U18511 ( .A1(n15218), .A2(n15222), .ZN(n15208) );
  XOR2_X1 U18512 ( .A(n15209), .B(n15208), .Z(n15378) );
  INV_X1 U18513 ( .A(n15210), .ZN(n15217) );
  INV_X1 U18514 ( .A(P2_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n18793) );
  NAND2_X1 U18515 ( .A1(n19085), .A2(P2_REIP_REG_19__SCAN_IN), .ZN(n15370) );
  OAI21_X1 U18516 ( .B1(n19113), .B2(n18793), .A(n15370), .ZN(n15212) );
  AOI21_X1 U18517 ( .B1(n18792), .B2(n19101), .A(n15212), .ZN(n15213) );
  OAI21_X1 U18518 ( .B1(n18799), .B2(n16174), .A(n15213), .ZN(n15214) );
  AOI21_X1 U18519 ( .B1(n15376), .B2(n19102), .A(n15214), .ZN(n15215) );
  OAI21_X1 U18520 ( .B1(n15378), .B2(n19108), .A(n15215), .ZN(P2_U2995) );
  OAI21_X1 U18521 ( .B1(n15394), .B2(n15411), .A(n15387), .ZN(n15216) );
  NAND2_X1 U18522 ( .A1(n15217), .A2(n15216), .ZN(n15393) );
  INV_X1 U18523 ( .A(n15218), .ZN(n15223) );
  AOI21_X1 U18524 ( .B1(n15220), .B2(n15222), .A(n15219), .ZN(n15221) );
  AOI21_X1 U18525 ( .B1(n15223), .B2(n15222), .A(n15221), .ZN(n15391) );
  INV_X1 U18526 ( .A(n18805), .ZN(n15226) );
  INV_X1 U18527 ( .A(P2_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n15224) );
  NAND2_X1 U18528 ( .A1(n19085), .A2(P2_REIP_REG_18__SCAN_IN), .ZN(n15383) );
  OAI21_X1 U18529 ( .B1(n19113), .B2(n15224), .A(n15383), .ZN(n15225) );
  AOI21_X1 U18530 ( .B1(n15226), .B2(n19101), .A(n15225), .ZN(n15227) );
  OAI21_X1 U18531 ( .B1(n18811), .B2(n16174), .A(n15227), .ZN(n15228) );
  AOI21_X1 U18532 ( .B1(n15391), .B2(n19087), .A(n15228), .ZN(n15229) );
  OAI21_X1 U18533 ( .B1(n15393), .B2(n19092), .A(n15229), .ZN(P2_U2996) );
  XNOR2_X1 U18534 ( .A(n15394), .B(n15411), .ZN(n15237) );
  XOR2_X1 U18535 ( .A(n15231), .B(n15230), .Z(n15408) );
  AOI22_X1 U18536 ( .A1(n19086), .A2(P2_PHYADDRPOINTER_REG_17__SCAN_IN), .B1(
        n19101), .B2(n18818), .ZN(n15234) );
  NOR2_X1 U18537 ( .A1(n19750), .A2(n18934), .ZN(n15232) );
  AOI21_X1 U18538 ( .B1(n18824), .B2(n19104), .A(n15232), .ZN(n15233) );
  NAND2_X1 U18539 ( .A1(n15234), .A2(n15233), .ZN(n15235) );
  AOI21_X1 U18540 ( .B1(n15408), .B2(n19087), .A(n15235), .ZN(n15236) );
  OAI21_X1 U18541 ( .B1(n15237), .B2(n19092), .A(n15236), .ZN(P2_U2997) );
  XNOR2_X1 U18542 ( .A(n15239), .B(n15238), .ZN(n15418) );
  INV_X1 U18543 ( .A(n15418), .ZN(n15246) );
  OAI21_X1 U18544 ( .B1(n15402), .B2(n15428), .A(n15405), .ZN(n15240) );
  NAND3_X1 U18545 ( .A1(n15240), .A2(n19102), .A3(n15394), .ZN(n15245) );
  INV_X1 U18546 ( .A(n18835), .ZN(n15243) );
  NOR2_X1 U18547 ( .A1(n15415), .A2(n18934), .ZN(n15242) );
  OAI22_X1 U18548 ( .A1(n19113), .A2(n10090), .B1(n19098), .B2(n18829), .ZN(
        n15241) );
  AOI211_X1 U18549 ( .C1(n15243), .C2(n19104), .A(n15242), .B(n15241), .ZN(
        n15244) );
  OAI211_X1 U18550 ( .C1(n15246), .C2(n19108), .A(n15245), .B(n15244), .ZN(
        P2_U2998) );
  XNOR2_X1 U18551 ( .A(n15247), .B(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n15433) );
  OR2_X1 U18552 ( .A1(n15249), .A2(n10054), .ZN(n15250) );
  XNOR2_X1 U18553 ( .A(n15251), .B(n15250), .ZN(n15431) );
  INV_X1 U18554 ( .A(n15252), .ZN(n18846) );
  OAI22_X1 U18555 ( .A1(n19113), .A2(n15253), .B1(n19098), .B2(n18846), .ZN(
        n15256) );
  NAND2_X1 U18556 ( .A1(n19085), .A2(P2_REIP_REG_15__SCAN_IN), .ZN(n15424) );
  OAI21_X1 U18557 ( .B1(n16174), .B2(n15254), .A(n15424), .ZN(n15255) );
  AOI211_X1 U18558 ( .C1(n15431), .C2(n19087), .A(n15256), .B(n15255), .ZN(
        n15257) );
  OAI21_X1 U18559 ( .B1(n15433), .B2(n19092), .A(n15257), .ZN(P2_U2999) );
  NOR3_X1 U18560 ( .A1(n21005), .A2(P2_INSTADDRPOINTER_REG_28__SCAN_IN), .A3(
        n15258), .ZN(n15259) );
  AOI211_X1 U18561 ( .C1(n16209), .C2(n15261), .A(n15260), .B(n15259), .ZN(
        n15262) );
  OAI21_X1 U18562 ( .B1(n15264), .B2(n15263), .A(n15262), .ZN(n15267) );
  NOR2_X1 U18563 ( .A1(n15265), .A2(n16223), .ZN(n15266) );
  AOI211_X2 U18564 ( .C1(n16041), .C2(n16219), .A(n15267), .B(n15266), .ZN(
        n15268) );
  INV_X1 U18565 ( .A(n15269), .ZN(n15271) );
  OAI211_X1 U18566 ( .C1(n16222), .C2(n16060), .A(n15271), .B(n15270), .ZN(
        n15272) );
  AOI21_X1 U18567 ( .B1(n15273), .B2(P2_INSTADDRPOINTER_REG_27__SCAN_IN), .A(
        n15272), .ZN(n15274) );
  OAI21_X1 U18568 ( .B1(n16048), .B2(n16212), .A(n15274), .ZN(n15275) );
  AOI21_X1 U18569 ( .B1(n15276), .B2(n12618), .A(n15275), .ZN(n15277) );
  OAI21_X1 U18570 ( .B1(n15278), .B2(n16217), .A(n15277), .ZN(P2_U3019) );
  NAND2_X1 U18571 ( .A1(n15279), .A2(n16227), .ZN(n15289) );
  NAND2_X1 U18572 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15280), .ZN(
        n15281) );
  AND2_X1 U18573 ( .A1(n15397), .A2(n15281), .ZN(n15305) );
  NAND2_X1 U18574 ( .A1(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n15302), .ZN(
        n15292) );
  XNOR2_X1 U18575 ( .A(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .B(
        P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n15284) );
  NAND2_X1 U18576 ( .A1(n16209), .A2(n16064), .ZN(n15283) );
  OAI211_X1 U18577 ( .C1(n15292), .C2(n15284), .A(n15283), .B(n15282), .ZN(
        n15287) );
  NOR2_X1 U18578 ( .A1(n15285), .A2(n16212), .ZN(n15286) );
  AOI211_X1 U18579 ( .C1(P2_INSTADDRPOINTER_REG_26__SCAN_IN), .C2(n15305), .A(
        n15287), .B(n15286), .ZN(n15288) );
  OAI211_X1 U18580 ( .C1(n15290), .C2(n16223), .A(n15289), .B(n15288), .ZN(
        P2_U3020) );
  NAND2_X1 U18581 ( .A1(n15305), .A2(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(
        n15295) );
  OAI21_X1 U18582 ( .B1(P2_INSTADDRPOINTER_REG_25__SCAN_IN), .B2(n15292), .A(
        n15291), .ZN(n15293) );
  AOI21_X1 U18583 ( .B1(n16209), .B2(n16074), .A(n15293), .ZN(n15294) );
  NAND2_X1 U18584 ( .A1(n15295), .A2(n15294), .ZN(n15296) );
  AOI21_X1 U18585 ( .B1(n16075), .B2(n16219), .A(n15296), .ZN(n15299) );
  NAND3_X1 U18586 ( .A1(n15297), .A2(n15119), .A3(n12618), .ZN(n15298) );
  OAI211_X1 U18587 ( .C1(n15300), .C2(n16217), .A(n15299), .B(n15298), .ZN(
        P2_U3021) );
  NAND2_X1 U18588 ( .A1(n15302), .A2(n15301), .ZN(n15307) );
  OAI21_X1 U18589 ( .B1(n16222), .B2(n16084), .A(n15303), .ZN(n15304) );
  AOI21_X1 U18590 ( .B1(n15305), .B2(P2_INSTADDRPOINTER_REG_24__SCAN_IN), .A(
        n15304), .ZN(n15306) );
  OAI211_X1 U18591 ( .C1(n16085), .C2(n16212), .A(n15307), .B(n15306), .ZN(
        n15308) );
  AOI21_X1 U18592 ( .B1(n15309), .B2(n12618), .A(n15308), .ZN(n15310) );
  OAI21_X1 U18593 ( .B1(n15311), .B2(n16217), .A(n15310), .ZN(P2_U3022) );
  NAND2_X1 U18594 ( .A1(n15396), .A2(n15397), .ZN(n15455) );
  OAI21_X1 U18595 ( .B1(n15312), .B2(n15471), .A(n15455), .ZN(n15350) );
  INV_X1 U18596 ( .A(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n15313) );
  NAND2_X1 U18597 ( .A1(n15312), .A2(n16197), .ZN(n15334) );
  AOI221_X1 U18598 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(
        P2_INSTADDRPOINTER_REG_22__SCAN_IN), .C1(n15313), .C2(n15338), .A(
        n15334), .ZN(n15315) );
  NOR2_X1 U18599 ( .A1(n18934), .A2(n10960), .ZN(n15314) );
  AOI211_X1 U18600 ( .C1(n16209), .C2(n16096), .A(n15315), .B(n15314), .ZN(
        n15316) );
  OAI21_X1 U18601 ( .B1(n16095), .B2(n16212), .A(n15316), .ZN(n15317) );
  AOI21_X1 U18602 ( .B1(P2_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n15350), .A(
        n15317), .ZN(n15321) );
  NAND3_X1 U18603 ( .A1(n15319), .A2(n16227), .A3(n15318), .ZN(n15320) );
  OAI211_X1 U18604 ( .C1(n15322), .C2(n16223), .A(n15321), .B(n15320), .ZN(
        P2_U3023) );
  AOI21_X1 U18605 ( .B1(n15338), .B2(n15324), .A(n15323), .ZN(n16126) );
  INV_X1 U18606 ( .A(n16126), .ZN(n15342) );
  INV_X1 U18607 ( .A(n15326), .ZN(n15327) );
  OR2_X1 U18608 ( .A1(n15328), .A2(n15327), .ZN(n15329) );
  XNOR2_X1 U18609 ( .A(n15325), .B(n15329), .ZN(n16128) );
  INV_X1 U18610 ( .A(n15350), .ZN(n15339) );
  INV_X1 U18611 ( .A(n15682), .ZN(n16127) );
  NOR2_X1 U18612 ( .A1(n15330), .A2(n14873), .ZN(n15331) );
  OR2_X1 U18613 ( .A1(n15332), .A2(n15331), .ZN(n16106) );
  NOR2_X1 U18614 ( .A1(n16222), .A2(n16106), .ZN(n15336) );
  NAND2_X1 U18615 ( .A1(P2_REIP_REG_22__SCAN_IN), .A2(n19085), .ZN(n15333) );
  OAI21_X1 U18616 ( .B1(P2_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n15334), .A(
        n15333), .ZN(n15335) );
  AOI211_X1 U18617 ( .C1(n16127), .C2(n16219), .A(n15336), .B(n15335), .ZN(
        n15337) );
  OAI21_X1 U18618 ( .B1(n15339), .B2(n15338), .A(n15337), .ZN(n15340) );
  AOI21_X1 U18619 ( .B1(n16128), .B2(n16227), .A(n15340), .ZN(n15341) );
  OAI21_X1 U18620 ( .B1(n15342), .B2(n16223), .A(n15341), .ZN(P2_U3024) );
  NAND2_X1 U18621 ( .A1(n15343), .A2(n16219), .ZN(n15345) );
  OAI211_X1 U18622 ( .C1(n16222), .C2(n15346), .A(n15345), .B(n15344), .ZN(
        n15349) );
  NOR3_X1 U18623 ( .A1(n15444), .A2(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .A3(
        n15347), .ZN(n15348) );
  AOI211_X1 U18624 ( .C1(P2_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(n15350), .A(
        n15349), .B(n15348), .ZN(n15353) );
  NAND2_X1 U18625 ( .A1(n15351), .A2(n16227), .ZN(n15352) );
  OAI211_X1 U18626 ( .C1(n15354), .C2(n16223), .A(n15353), .B(n15352), .ZN(
        P2_U3025) );
  NAND3_X1 U18627 ( .A1(n16197), .A2(n15358), .A3(n15374), .ZN(n15373) );
  INV_X1 U18628 ( .A(n15358), .ZN(n15355) );
  NAND2_X1 U18629 ( .A1(n15397), .A2(n15355), .ZN(n15356) );
  AND2_X1 U18630 ( .A1(n15455), .A2(n15356), .ZN(n15388) );
  AOI21_X1 U18631 ( .B1(n15373), .B2(n15388), .A(n15357), .ZN(n15364) );
  NAND4_X1 U18632 ( .A1(n16197), .A2(P2_INSTADDRPOINTER_REG_19__SCAN_IN), .A3(
        n15358), .A4(n15357), .ZN(n15361) );
  AOI21_X1 U18633 ( .B1(n16209), .B2(n16113), .A(n15359), .ZN(n15360) );
  OAI211_X1 U18634 ( .C1(n15362), .C2(n16212), .A(n15361), .B(n15360), .ZN(
        n15363) );
  NOR2_X1 U18635 ( .A1(n15364), .A2(n15363), .ZN(n15368) );
  NAND3_X1 U18636 ( .A1(n15366), .A2(n16227), .A3(n15365), .ZN(n15367) );
  OAI211_X1 U18637 ( .C1(n15369), .C2(n16223), .A(n15368), .B(n15367), .ZN(
        P2_U3026) );
  OAI21_X1 U18638 ( .B1(n18799), .B2(n16212), .A(n15370), .ZN(n15371) );
  AOI21_X1 U18639 ( .B1(n16209), .B2(n18797), .A(n15371), .ZN(n15372) );
  OAI211_X1 U18640 ( .C1(n15388), .C2(n15374), .A(n15373), .B(n15372), .ZN(
        n15375) );
  AOI21_X1 U18641 ( .B1(n15376), .B2(n12618), .A(n15375), .ZN(n15377) );
  OAI21_X1 U18642 ( .B1(n15378), .B2(n16217), .A(n15377), .ZN(P2_U3027) );
  NOR3_X1 U18643 ( .A1(n15444), .A2(P2_INSTADDRPOINTER_REG_18__SCAN_IN), .A3(
        n15379), .ZN(n15390) );
  INV_X1 U18644 ( .A(n18811), .ZN(n15385) );
  NAND2_X1 U18645 ( .A1(n14065), .A2(n15380), .ZN(n15381) );
  NAND2_X1 U18646 ( .A1(n15382), .A2(n15381), .ZN(n18810) );
  OAI21_X1 U18647 ( .B1(n16222), .B2(n18810), .A(n15383), .ZN(n15384) );
  AOI21_X1 U18648 ( .B1(n15385), .B2(n16219), .A(n15384), .ZN(n15386) );
  OAI21_X1 U18649 ( .B1(n15388), .B2(n15387), .A(n15386), .ZN(n15389) );
  AOI211_X1 U18650 ( .C1(n15391), .C2(n16227), .A(n15390), .B(n15389), .ZN(
        n15392) );
  OAI21_X1 U18651 ( .B1(n15393), .B2(n16223), .A(n15392), .ZN(P2_U3028) );
  OAI21_X1 U18652 ( .B1(n12618), .B2(n15395), .A(n15394), .ZN(n15399) );
  OR2_X1 U18653 ( .A1(n15396), .A2(n15403), .ZN(n15398) );
  NAND2_X1 U18654 ( .A1(n15398), .A2(n15397), .ZN(n15429) );
  OAI211_X1 U18655 ( .C1(P2_INSTADDRPOINTER_REG_15__SCAN_IN), .C2(n15400), .A(
        n15399), .B(n15429), .ZN(n15419) );
  AOI21_X1 U18656 ( .B1(n15405), .B2(n15514), .A(n15419), .ZN(n15412) );
  OAI22_X1 U18657 ( .A1(n16222), .A2(n15401), .B1(n19750), .B2(n18934), .ZN(
        n15407) );
  NOR2_X1 U18658 ( .A1(n15444), .A2(n15403), .ZN(n15423) );
  OAI21_X2 U18659 ( .B1(n15404), .B2(n15423), .A(
        P2_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15422) );
  NOR3_X1 U18660 ( .A1(n15422), .A2(P2_INSTADDRPOINTER_REG_17__SCAN_IN), .A3(
        n15405), .ZN(n15406) );
  AOI211_X1 U18661 ( .C1(n18824), .C2(n16219), .A(n15407), .B(n15406), .ZN(
        n15410) );
  NAND2_X1 U18662 ( .A1(n15408), .A2(n16227), .ZN(n15409) );
  OAI211_X1 U18663 ( .C1(n15412), .C2(n15411), .A(n15410), .B(n15409), .ZN(
        P2_U3029) );
  NOR2_X1 U18664 ( .A1(n16212), .A2(n18835), .ZN(n15417) );
  OR2_X1 U18665 ( .A1(n15413), .A2(n13849), .ZN(n15414) );
  NAND2_X1 U18666 ( .A1(n14066), .A2(n15414), .ZN(n18968) );
  OAI22_X1 U18667 ( .A1(n16222), .A2(n18968), .B1(n15415), .B2(n18934), .ZN(
        n15416) );
  AOI211_X1 U18668 ( .C1(n15418), .C2(n16227), .A(n15417), .B(n15416), .ZN(
        n15421) );
  NAND2_X1 U18669 ( .A1(n15419), .A2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(
        n15420) );
  OAI211_X1 U18670 ( .C1(n15422), .C2(P2_INSTADDRPOINTER_REG_16__SCAN_IN), .A(
        n15421), .B(n15420), .ZN(P2_U3030) );
  NAND2_X1 U18671 ( .A1(n15423), .A2(n15428), .ZN(n15427) );
  OAI21_X1 U18672 ( .B1(n16222), .B2(n18851), .A(n15424), .ZN(n15425) );
  AOI21_X1 U18673 ( .B1(n16219), .B2(n18847), .A(n15425), .ZN(n15426) );
  OAI211_X1 U18674 ( .C1(n15429), .C2(n15428), .A(n15427), .B(n15426), .ZN(
        n15430) );
  AOI21_X1 U18675 ( .B1(n15431), .B2(n16227), .A(n15430), .ZN(n15432) );
  OAI21_X1 U18676 ( .B1(n15433), .B2(n16223), .A(n15432), .ZN(P2_U3031) );
  INV_X1 U18677 ( .A(n15434), .ZN(n15435) );
  OR2_X1 U18678 ( .A1(n16134), .A2(n15435), .ZN(n15439) );
  NAND2_X1 U18679 ( .A1(n15437), .A2(n15436), .ZN(n15438) );
  NAND2_X1 U18680 ( .A1(n15439), .A2(n15438), .ZN(n16139) );
  OAI21_X1 U18681 ( .B1(n16146), .B2(P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A(
        n15440), .ZN(n16140) );
  OR2_X1 U18682 ( .A1(n16140), .A2(n16223), .ZN(n15451) );
  OR2_X1 U18683 ( .A1(n15461), .A2(n15443), .ZN(n15441) );
  NAND2_X1 U18684 ( .A1(n16197), .A2(n15441), .ZN(n15442) );
  NAND2_X1 U18685 ( .A1(n15442), .A2(n15455), .ZN(n16192) );
  OAI21_X1 U18686 ( .B1(n15461), .B2(n15444), .A(n15443), .ZN(n15449) );
  OR2_X1 U18687 ( .A1(n16222), .A2(n18867), .ZN(n15446) );
  NAND2_X1 U18688 ( .A1(n19085), .A2(P2_REIP_REG_13__SCAN_IN), .ZN(n15445) );
  OAI211_X1 U18689 ( .C1(n15447), .C2(n16212), .A(n15446), .B(n15445), .ZN(
        n15448) );
  AOI21_X1 U18690 ( .B1(n16192), .B2(n15449), .A(n15448), .ZN(n15450) );
  OAI211_X1 U18691 ( .C1(n16139), .C2(n16217), .A(n15451), .B(n15450), .ZN(
        P2_U3033) );
  OAI21_X1 U18692 ( .B1(n15454), .B2(n15453), .A(n15452), .ZN(n16149) );
  INV_X1 U18693 ( .A(n16149), .ZN(n15464) );
  NOR2_X1 U18694 ( .A1(n15160), .A2(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(
        n16145) );
  OR3_X1 U18695 ( .A1(n16146), .A2(n16145), .A3(n16223), .ZN(n15463) );
  NOR2_X1 U18696 ( .A1(n16212), .A2(n18874), .ZN(n15460) );
  NAND2_X1 U18697 ( .A1(P2_REIP_REG_12__SCAN_IN), .A2(n19085), .ZN(n15458) );
  INV_X1 U18698 ( .A(n15455), .ZN(n15456) );
  NAND2_X1 U18699 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n15456), .ZN(
        n15457) );
  OAI211_X1 U18700 ( .C1(n16222), .C2(n18875), .A(n15458), .B(n15457), .ZN(
        n15459) );
  AOI211_X1 U18701 ( .C1(n16197), .C2(n15461), .A(n15460), .B(n15459), .ZN(
        n15462) );
  OAI211_X1 U18702 ( .C1(n15464), .C2(n16217), .A(n15463), .B(n15462), .ZN(
        P2_U3034) );
  NOR2_X1 U18703 ( .A1(n10060), .A2(n15467), .ZN(n15468) );
  XNOR2_X1 U18704 ( .A(n15465), .B(n15468), .ZN(n16152) );
  OAI21_X1 U18705 ( .B1(P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n9848), .A(
        n15469), .ZN(n16153) );
  OR2_X1 U18706 ( .A1(n16153), .A2(n16223), .ZN(n15478) );
  XNOR2_X1 U18707 ( .A(n15470), .B(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n15476) );
  INV_X1 U18708 ( .A(n18889), .ZN(n15474) );
  OR2_X1 U18709 ( .A1(n16222), .A2(n18894), .ZN(n15473) );
  NOR2_X1 U18710 ( .A1(n15471), .A2(n15495), .ZN(n15489) );
  AOI22_X1 U18711 ( .A1(n19085), .A2(P2_REIP_REG_11__SCAN_IN), .B1(
        P2_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15489), .ZN(n15472) );
  OAI211_X1 U18712 ( .C1(n15474), .C2(n16212), .A(n15473), .B(n15472), .ZN(
        n15475) );
  AOI21_X1 U18713 ( .B1(n15488), .B2(n15476), .A(n15475), .ZN(n15477) );
  OAI211_X1 U18714 ( .C1(n16152), .C2(n16217), .A(n15478), .B(n15477), .ZN(
        P2_U3035) );
  NAND2_X1 U18715 ( .A1(n15480), .A2(n15479), .ZN(n15483) );
  NOR2_X1 U18716 ( .A1(n15481), .A2(n10311), .ZN(n15482) );
  XNOR2_X1 U18717 ( .A(n15483), .B(n15482), .ZN(n16159) );
  NOR2_X1 U18718 ( .A1(n10225), .A2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(
        n16158) );
  OR3_X1 U18719 ( .A1(n9848), .A2(n16158), .A3(n16223), .ZN(n15494) );
  XNOR2_X1 U18720 ( .A(n15485), .B(n15484), .ZN(n18981) );
  INV_X1 U18721 ( .A(n18981), .ZN(n15492) );
  NOR2_X1 U18722 ( .A1(n12751), .A2(n18934), .ZN(n15486) );
  AOI221_X1 U18723 ( .B1(n15489), .B2(P2_INSTADDRPOINTER_REG_10__SCAN_IN), 
        .C1(n15488), .C2(n15487), .A(n15486), .ZN(n15490) );
  OAI21_X1 U18724 ( .B1(n16212), .B2(n18900), .A(n15490), .ZN(n15491) );
  AOI21_X1 U18725 ( .B1(n16209), .B2(n15492), .A(n15491), .ZN(n15493) );
  OAI211_X1 U18726 ( .C1(n16159), .C2(n16217), .A(n15494), .B(n15493), .ZN(
        P2_U3036) );
  INV_X1 U18727 ( .A(n18984), .ZN(n15501) );
  AOI21_X1 U18728 ( .B1(n15497), .B2(n15496), .A(n15495), .ZN(n15500) );
  OAI22_X1 U18729 ( .A1(n16212), .A2(n15498), .B1(n14218), .B2(n18934), .ZN(
        n15499) );
  AOI211_X1 U18730 ( .C1(n15501), .C2(n16209), .A(n15500), .B(n15499), .ZN(
        n15504) );
  NAND2_X1 U18731 ( .A1(n15502), .A2(n16227), .ZN(n15503) );
  OAI211_X1 U18732 ( .C1(n15505), .C2(n16223), .A(n15504), .B(n15503), .ZN(
        P2_U3037) );
  INV_X1 U18733 ( .A(n15506), .ZN(n15510) );
  OAI22_X1 U18734 ( .A1(n15507), .A2(n16212), .B1(n16222), .B2(n19003), .ZN(
        n15508) );
  AOI211_X1 U18735 ( .C1(n12618), .C2(n15510), .A(n15509), .B(n15508), .ZN(
        n15517) );
  AOI22_X1 U18736 ( .A1(n16227), .A2(n15512), .B1(n15511), .B2(
        P2_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n15516) );
  OAI211_X1 U18737 ( .C1(P2_INSTADDRPOINTER_REG_1__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n15514), .B(n15513), .ZN(n15515) );
  NAND3_X1 U18738 ( .A1(n15517), .A2(n15516), .A3(n15515), .ZN(P2_U3045) );
  NAND2_X1 U18739 ( .A1(n18950), .A2(n15541), .ZN(n15522) );
  INV_X1 U18740 ( .A(n15518), .ZN(n15519) );
  NOR2_X1 U18741 ( .A1(n15520), .A2(n15519), .ZN(n15533) );
  INV_X1 U18742 ( .A(n12628), .ZN(n15531) );
  MUX2_X1 U18743 ( .A(n15533), .B(n15531), .S(
        P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .Z(n15521) );
  NAND2_X1 U18744 ( .A1(n15522), .A2(n15521), .ZN(n16238) );
  INV_X1 U18745 ( .A(n15523), .ZN(n15524) );
  AOI22_X1 U18746 ( .A1(n18917), .A2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B1(
        n18942), .B2(n18929), .ZN(n15528) );
  AOI222_X1 U18747 ( .A1(n16238), .A2(n15552), .B1(n15524), .B2(n15551), .C1(
        P2_STATE2_REG_1__SCAN_IN), .C2(n15528), .ZN(n15526) );
  NAND2_X1 U18748 ( .A1(n15662), .A2(P2_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(
        n15525) );
  OAI21_X1 U18749 ( .B1(n15526), .B2(n15662), .A(n15525), .ZN(P2_U3601) );
  NOR2_X1 U18750 ( .A1(n15528), .A2(n15527), .ZN(n15549) );
  INV_X1 U18751 ( .A(n15549), .ZN(n15537) );
  OAI21_X1 U18752 ( .B1(n18929), .B2(n15530), .A(n15529), .ZN(n15550) );
  INV_X1 U18753 ( .A(n15552), .ZN(n19785) );
  OAI22_X1 U18754 ( .A1(n15533), .A2(n15532), .B1(n15531), .B2(
        P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n15534) );
  AOI22_X1 U18755 ( .A1(n15536), .A2(n15541), .B1(n15535), .B2(n15534), .ZN(
        n16240) );
  OAI222_X1 U18756 ( .A1(n16286), .A2(n19808), .B1(n15537), .B2(n15550), .C1(
        n19785), .C2(n16240), .ZN(n15538) );
  INV_X1 U18757 ( .A(n15662), .ZN(n15665) );
  MUX2_X1 U18758 ( .A(P2_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n15538), .S(
        n15665), .Z(P2_U3600) );
  NAND2_X1 U18759 ( .A1(n15540), .A2(n15539), .ZN(n15547) );
  NAND2_X1 U18760 ( .A1(n19105), .A2(n15541), .ZN(n15546) );
  NOR2_X1 U18761 ( .A1(n15542), .A2(n10546), .ZN(n15543) );
  AOI22_X1 U18762 ( .A1(n15544), .A2(n15547), .B1(n15543), .B2(n12628), .ZN(
        n15545) );
  OAI211_X1 U18763 ( .C1(n15548), .C2(n15547), .A(n15546), .B(n15545), .ZN(
        n16235) );
  AOI222_X1 U18764 ( .A1(n16235), .A2(n15552), .B1(n19804), .B2(n15551), .C1(
        n15550), .C2(n15549), .ZN(n15553) );
  MUX2_X1 U18765 ( .A(n15554), .B(n15553), .S(n15665), .Z(n15555) );
  INV_X1 U18766 ( .A(n15555), .ZN(P2_U3599) );
  AOI22_X1 U18767 ( .A1(n9846), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n15559) );
  AOI22_X1 U18768 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n15558) );
  AOI22_X1 U18769 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(
        n9842), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n15557) );
  AOI22_X1 U18770 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n15556) );
  NAND4_X1 U18771 ( .A1(n15559), .A2(n15558), .A3(n15557), .A4(n15556), .ZN(
        n15566) );
  AOI22_X1 U18772 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9812), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n15564) );
  AOI22_X1 U18773 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(n9841), .B2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n15563) );
  AOI22_X1 U18774 ( .A1(n9838), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n17068), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n15562) );
  AOI22_X1 U18775 ( .A1(n9811), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(n9815), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n15561) );
  NAND4_X1 U18776 ( .A1(n15564), .A2(n15563), .A3(n15562), .A4(n15561), .ZN(
        n15565) );
  NOR2_X1 U18777 ( .A1(n15566), .A2(n15565), .ZN(n16859) );
  AOI22_X1 U18778 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17024), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n15570) );
  AOI22_X1 U18779 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n15569) );
  AOI22_X1 U18780 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(n9816), .B2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n15568) );
  AOI22_X1 U18781 ( .A1(n15609), .A2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n15567) );
  NAND4_X1 U18782 ( .A1(n15570), .A2(n15569), .A3(n15568), .A4(n15567), .ZN(
        n15576) );
  AOI22_X1 U18783 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n15574) );
  AOI22_X1 U18784 ( .A1(n17068), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n9846), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n15573) );
  AOI22_X1 U18785 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n15572) );
  AOI22_X1 U18786 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n15571) );
  NAND4_X1 U18787 ( .A1(n15574), .A2(n15573), .A3(n15572), .A4(n15571), .ZN(
        n15575) );
  NOR2_X1 U18788 ( .A1(n15576), .A2(n15575), .ZN(n16869) );
  AOI22_X1 U18789 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9816), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n15580) );
  AOI22_X1 U18790 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n15579) );
  AOI22_X1 U18791 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n15578) );
  AOI22_X1 U18792 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9842), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n15577) );
  NAND4_X1 U18793 ( .A1(n15580), .A2(n15579), .A3(n15578), .A4(n15577), .ZN(
        n15586) );
  AOI22_X1 U18794 ( .A1(n9809), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(n9830), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n15584) );
  AOI22_X1 U18795 ( .A1(n9838), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n9846), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n15583) );
  AOI22_X1 U18796 ( .A1(n17024), .A2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n15582) );
  AOI22_X1 U18797 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9841), .B2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n15581) );
  NAND4_X1 U18798 ( .A1(n15584), .A2(n15583), .A3(n15582), .A4(n15581), .ZN(
        n15585) );
  NOR2_X1 U18799 ( .A1(n15586), .A2(n15585), .ZN(n16879) );
  AOI22_X1 U18800 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n15590) );
  AOI22_X1 U18801 ( .A1(n9809), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(n9815), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n15589) );
  AOI22_X1 U18802 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9818), .B2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n15588) );
  AOI22_X1 U18803 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n15587) );
  NAND4_X1 U18804 ( .A1(n15590), .A2(n15589), .A3(n15588), .A4(n15587), .ZN(
        n15596) );
  AOI22_X1 U18805 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n15594) );
  AOI22_X1 U18806 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n15593) );
  AOI22_X1 U18807 ( .A1(n17024), .A2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n15592) );
  AOI22_X1 U18808 ( .A1(n9811), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(n9846), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n15591) );
  NAND4_X1 U18809 ( .A1(n15594), .A2(n15593), .A3(n15592), .A4(n15591), .ZN(
        n15595) );
  NOR2_X1 U18810 ( .A1(n15596), .A2(n15595), .ZN(n16880) );
  NOR2_X1 U18811 ( .A1(n16879), .A2(n16880), .ZN(n16878) );
  AOI22_X1 U18812 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9830), .B1(
        n17069), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n15608) );
  AOI22_X1 U18813 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_7__1__SCAN_IN), .B2(n9815), .ZN(n15607) );
  AOI22_X1 U18814 ( .A1(n9810), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(n9811), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n15597) );
  OAI21_X1 U18815 ( .B1(n15599), .B2(n15598), .A(n15597), .ZN(n15605) );
  AOI22_X1 U18816 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n17049), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n15609), .ZN(n15603) );
  AOI22_X1 U18817 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_12__1__SCAN_IN), .B1(
        n9846), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n15602) );
  AOI22_X1 U18818 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17048), .B1(
        n9819), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n15601) );
  AOI22_X1 U18819 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n17034), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n15600) );
  NAND4_X1 U18820 ( .A1(n15603), .A2(n15602), .A3(n15601), .A4(n15600), .ZN(
        n15604) );
  AOI211_X1 U18821 ( .C1(n9818), .C2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A(
        n15605), .B(n15604), .ZN(n15606) );
  NAND3_X1 U18822 ( .A1(n15608), .A2(n15607), .A3(n15606), .ZN(n16874) );
  NAND2_X1 U18823 ( .A1(n16878), .A2(n16874), .ZN(n16873) );
  NOR2_X1 U18824 ( .A1(n16869), .A2(n16873), .ZN(n16868) );
  AOI22_X1 U18825 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n15620) );
  AOI22_X1 U18826 ( .A1(n9841), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n17024), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n15619) );
  INV_X1 U18827 ( .A(P3_INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n20972) );
  AOI22_X1 U18828 ( .A1(n9811), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n15610) );
  OAI21_X1 U18829 ( .B1(n15611), .B2(n20972), .A(n15610), .ZN(n15617) );
  AOI22_X1 U18830 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .B1(
        n17069), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n15615) );
  AOI22_X1 U18831 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9815), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n15614) );
  AOI22_X1 U18832 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n15613) );
  AOI22_X1 U18833 ( .A1(n9846), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n15612) );
  NAND4_X1 U18834 ( .A1(n15615), .A2(n15614), .A3(n15613), .A4(n15612), .ZN(
        n15616) );
  AOI211_X1 U18835 ( .C1(n9809), .C2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A(
        n15617), .B(n15616), .ZN(n15618) );
  NAND3_X1 U18836 ( .A1(n15620), .A2(n15619), .A3(n15618), .ZN(n16864) );
  NAND2_X1 U18837 ( .A1(n16868), .A2(n16864), .ZN(n16863) );
  NOR2_X1 U18838 ( .A1(n16859), .A2(n16863), .ZN(n16858) );
  AOI22_X1 U18839 ( .A1(n9810), .A2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .B1(n9830), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15631) );
  AOI22_X1 U18840 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n15630) );
  INV_X1 U18841 ( .A(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n20969) );
  AOI22_X1 U18842 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n15621) );
  OAI21_X1 U18843 ( .B1(n15622), .B2(n20969), .A(n15621), .ZN(n15628) );
  AOI22_X1 U18844 ( .A1(n17069), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(
        n9815), .B2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n15626) );
  AOI22_X1 U18845 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n15625) );
  AOI22_X1 U18846 ( .A1(n17024), .A2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .B1(
        n9846), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15624) );
  AOI22_X1 U18847 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(
        n9842), .B2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n15623) );
  NAND4_X1 U18848 ( .A1(n15626), .A2(n15625), .A3(n15624), .A4(n15623), .ZN(
        n15627) );
  AOI211_X1 U18849 ( .C1(n9818), .C2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n15628), .B(n15627), .ZN(n15629) );
  NAND3_X1 U18850 ( .A1(n15631), .A2(n15630), .A3(n15629), .ZN(n15632) );
  NAND2_X1 U18851 ( .A1(n16858), .A2(n15632), .ZN(n16851) );
  OAI21_X1 U18852 ( .B1(n16858), .B2(n15632), .A(n16851), .ZN(n17127) );
  NAND3_X1 U18853 ( .A1(n18134), .A2(n15633), .A3(n18117), .ZN(n15635) );
  NAND2_X1 U18854 ( .A1(n15635), .A2(n15634), .ZN(n15742) );
  NOR2_X2 U18855 ( .A1(n17107), .A2(n18134), .ZN(n17101) );
  INV_X2 U18856 ( .A(n17101), .ZN(n17109) );
  INV_X1 U18857 ( .A(P3_EBX_REG_28__SCAN_IN), .ZN(n16819) );
  NAND2_X1 U18858 ( .A1(P3_EBX_REG_6__SCAN_IN), .A2(P3_EBX_REG_5__SCAN_IN), 
        .ZN(n15650) );
  INV_X1 U18859 ( .A(n15650), .ZN(n17077) );
  INV_X1 U18860 ( .A(P3_EBX_REG_0__SCAN_IN), .ZN(n17105) );
  INV_X1 U18861 ( .A(P3_EBX_REG_1__SCAN_IN), .ZN(n17103) );
  NOR2_X1 U18862 ( .A1(n17105), .A2(n17103), .ZN(n17097) );
  AND2_X1 U18863 ( .A1(P3_EBX_REG_2__SCAN_IN), .A2(n17097), .ZN(n17090) );
  NAND3_X1 U18864 ( .A1(P3_EBX_REG_4__SCAN_IN), .A2(P3_EBX_REG_3__SCAN_IN), 
        .A3(n17090), .ZN(n17086) );
  NAND2_X1 U18865 ( .A1(P3_EBX_REG_13__SCAN_IN), .A2(P3_EBX_REG_12__SCAN_IN), 
        .ZN(n15652) );
  NAND2_X1 U18866 ( .A1(P3_EBX_REG_15__SCAN_IN), .A2(P3_EBX_REG_14__SCAN_IN), 
        .ZN(n16974) );
  NAND4_X1 U18867 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(P3_EBX_REG_11__SCAN_IN), 
        .A3(P3_EBX_REG_10__SCAN_IN), .A4(P3_EBX_REG_9__SCAN_IN), .ZN(n15636)
         );
  NOR4_X1 U18868 ( .A1(n17086), .A2(n15652), .A3(n16974), .A4(n15636), .ZN(
        n15637) );
  NAND4_X1 U18869 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .A3(n17077), .A4(n15637), .ZN(n16975) );
  NOR2_X1 U18870 ( .A1(n17107), .A2(n16975), .ZN(n16961) );
  NAND2_X1 U18871 ( .A1(P3_EBX_REG_17__SCAN_IN), .A2(n16961), .ZN(n16960) );
  NAND2_X1 U18872 ( .A1(P3_EBX_REG_19__SCAN_IN), .A2(n16949), .ZN(n16935) );
  NOR2_X1 U18873 ( .A1(n17153), .A2(n16935), .ZN(n16923) );
  NAND2_X1 U18874 ( .A1(P3_EBX_REG_20__SCAN_IN), .A2(n16923), .ZN(n16911) );
  NOR2_X1 U18875 ( .A1(n16562), .A2(n16911), .ZN(n16884) );
  NAND2_X1 U18876 ( .A1(P3_EBX_REG_22__SCAN_IN), .A2(n16884), .ZN(n16877) );
  NAND2_X1 U18877 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(n16883), .ZN(n16867) );
  NOR2_X1 U18878 ( .A1(n16520), .A2(n16867), .ZN(n16872) );
  NAND2_X1 U18879 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(n16872), .ZN(n16857) );
  NOR3_X1 U18880 ( .A1(n16819), .A2(n16818), .A3(n16857), .ZN(n16853) );
  NOR2_X1 U18881 ( .A1(n17101), .A2(n16853), .ZN(n16849) );
  NOR2_X1 U18882 ( .A1(n16818), .A2(n16857), .ZN(n16862) );
  AOI22_X1 U18883 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16849), .B1(n16862), 
        .B2(n16819), .ZN(n15638) );
  OAI21_X1 U18884 ( .B1(n17127), .B2(n17109), .A(n15638), .ZN(P3_U2675) );
  AOI22_X1 U18885 ( .A1(n17024), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n15649) );
  AOI22_X1 U18886 ( .A1(n17069), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n9845), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n15648) );
  AOI22_X1 U18887 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(n9815), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n15639) );
  OAI21_X1 U18888 ( .B1(n11658), .B2(n20969), .A(n15639), .ZN(n15646) );
  AOI22_X1 U18889 ( .A1(n9809), .A2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .B1(n9819), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n15644) );
  AOI22_X1 U18890 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(n9830), .B2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n15643) );
  AOI22_X1 U18891 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n15642) );
  AOI22_X1 U18892 ( .A1(n15609), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n15641) );
  NAND4_X1 U18893 ( .A1(n15644), .A2(n15643), .A3(n15642), .A4(n15641), .ZN(
        n15645) );
  AOI211_X1 U18894 ( .C1(n9813), .C2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A(
        n15646), .B(n15645), .ZN(n15647) );
  NAND3_X1 U18895 ( .A1(n15649), .A2(n15648), .A3(n15647), .ZN(n17201) );
  INV_X1 U18896 ( .A(n17201), .ZN(n15654) );
  NOR3_X1 U18897 ( .A1(n17107), .A2(n17086), .A3(n15650), .ZN(n17084) );
  NAND3_X1 U18898 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(P3_EBX_REG_7__SCAN_IN), 
        .A3(n17084), .ZN(n17060) );
  NOR2_X1 U18899 ( .A1(n16701), .A2(n17060), .ZN(n17062) );
  NAND2_X1 U18900 ( .A1(P3_EBX_REG_10__SCAN_IN), .A2(n17062), .ZN(n17046) );
  NOR2_X1 U18901 ( .A1(n16679), .A2(n17046), .ZN(n17033) );
  INV_X1 U18902 ( .A(n17033), .ZN(n15651) );
  NOR2_X1 U18903 ( .A1(n15652), .A2(n15651), .ZN(n17002) );
  INV_X1 U18904 ( .A(n17002), .ZN(n16973) );
  OAI221_X1 U18905 ( .B1(P3_EBX_REG_13__SCAN_IN), .B2(P3_EBX_REG_12__SCAN_IN), 
        .C1(P3_EBX_REG_13__SCAN_IN), .C2(n17033), .A(n16973), .ZN(n15653) );
  AOI22_X1 U18906 ( .A1(n17101), .A2(n15654), .B1(n15653), .B2(n17109), .ZN(
        P3_U2690) );
  NAND2_X1 U18907 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n18323) );
  AOI221_X1 U18908 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18323), .C1(n15656), 
        .C2(n18323), .A(n15655), .ZN(n18086) );
  NOR2_X1 U18909 ( .A1(n15657), .A2(n20944), .ZN(n15658) );
  OAI21_X1 U18910 ( .B1(n15658), .B2(n16306), .A(n18087), .ZN(n18084) );
  AOI22_X1 U18911 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n18086), .B1(
        n18084), .B2(n18576), .ZN(P3_U2865) );
  NOR2_X1 U18912 ( .A1(n12562), .A2(n15660), .ZN(n15661) );
  NAND2_X1 U18913 ( .A1(n15659), .A2(n15661), .ZN(n16262) );
  OR3_X1 U18914 ( .A1(n15662), .A2(n19785), .A3(n16262), .ZN(n15663) );
  OAI21_X1 U18915 ( .B1(n15665), .B2(n15664), .A(n15663), .ZN(P2_U3595) );
  INV_X1 U18916 ( .A(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n16329) );
  NOR2_X1 U18917 ( .A1(n17649), .A2(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(
        n15666) );
  NOR3_X2 U18918 ( .A1(n15668), .A2(n17375), .A3(n17604), .ZN(n15727) );
  INV_X1 U18919 ( .A(n15727), .ZN(n15669) );
  NAND2_X1 U18920 ( .A1(n15726), .A2(n15669), .ZN(n15670) );
  XOR2_X1 U18921 ( .A(n16329), .B(n15670), .Z(n16344) );
  NAND2_X1 U18922 ( .A1(n17375), .A2(n16345), .ZN(n15672) );
  NAND2_X1 U18923 ( .A1(n15677), .A2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(
        n16349) );
  NOR2_X1 U18924 ( .A1(n17374), .A2(n16349), .ZN(n16328) );
  NAND2_X1 U18925 ( .A1(n16315), .A2(n18066), .ZN(n17791) );
  NOR2_X1 U18926 ( .A1(n17762), .A2(n16349), .ZN(n16339) );
  NAND2_X1 U18927 ( .A1(n18052), .A2(n18073), .ZN(n18079) );
  OAI22_X1 U18928 ( .A1(n16328), .A2(n17791), .B1(n16339), .B2(n18079), .ZN(
        n15671) );
  NOR2_X1 U18929 ( .A1(n18055), .A2(n15671), .ZN(n15731) );
  OAI221_X1 U18930 ( .B1(n18061), .B2(n15673), .C1(n18061), .C2(n15672), .A(
        n15731), .ZN(n15674) );
  AOI22_X1 U18931 ( .A1(n9820), .A2(P3_REIP_REG_29__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n15674), .ZN(n15679) );
  NAND3_X1 U18932 ( .A1(n18073), .A2(n15675), .A3(n17779), .ZN(n16347) );
  INV_X1 U18933 ( .A(n17791), .ZN(n17995) );
  NAND2_X1 U18934 ( .A1(n17760), .A2(n17995), .ZN(n15676) );
  OAI211_X1 U18935 ( .C1(n18079), .C2(n17762), .A(n16347), .B(n15676), .ZN(
        n15733) );
  NAND3_X1 U18936 ( .A1(n15677), .A2(n16329), .A3(n15733), .ZN(n15678) );
  OAI211_X1 U18937 ( .C1(n16344), .C2(n17909), .A(n15679), .B(n15678), .ZN(
        P3_U2833) );
  AOI22_X1 U18938 ( .A1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n18958), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n18885), .ZN(n15691) );
  OAI22_X1 U18939 ( .A1(n15680), .A2(n18947), .B1(n18840), .B2(n15003), .ZN(
        n15681) );
  INV_X1 U18940 ( .A(n15681), .ZN(n15690) );
  OAI22_X1 U18941 ( .A1(n15682), .A2(n18937), .B1(n16106), .B2(n18945), .ZN(
        n15683) );
  INV_X1 U18942 ( .A(n15683), .ZN(n15689) );
  OAI21_X1 U18943 ( .B1(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n9908), .A(
        n15686), .ZN(n16131) );
  NAND2_X1 U18944 ( .A1(n15687), .A2(n16131), .ZN(n16006) );
  OAI211_X1 U18945 ( .C1(n15687), .C2(n16131), .A(n18890), .B(n16006), .ZN(
        n15688) );
  NAND4_X1 U18946 ( .A1(n15691), .A2(n15690), .A3(n15689), .A4(n15688), .ZN(
        P2_U2833) );
  NOR4_X1 U18947 ( .A1(n15693), .A2(P1_STATEBS16_REG_SCAN_IN), .A3(n15692), 
        .A4(n20122), .ZN(n15694) );
  AOI221_X1 U18948 ( .B1(n15695), .B2(n20689), .C1(n15993), .C2(n20689), .A(
        n15694), .ZN(n15996) );
  AOI211_X1 U18949 ( .C1(P1_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .C2(n15697), .A(
        n20551), .B(n15696), .ZN(n15698) );
  INV_X1 U18950 ( .A(n15698), .ZN(n15702) );
  OAI22_X1 U18951 ( .A1(n15700), .A2(n15699), .B1(n15698), .B2(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n15701) );
  OAI21_X1 U18952 ( .B1(n20440), .B2(n15702), .A(n15701), .ZN(n15705) );
  INV_X1 U18953 ( .A(n15703), .ZN(n15704) );
  AOI222_X1 U18954 ( .A1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n15705), 
        .B1(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n15704), .C1(n15705), 
        .C2(n15704), .ZN(n15707) );
  AND2_X1 U18955 ( .A1(n15708), .A2(n15707), .ZN(n15706) );
  OAI221_X1 U18956 ( .B1(n15708), .B2(n15707), .C1(n20184), .C2(n15706), .A(
        n20100), .ZN(n15715) );
  NOR2_X1 U18957 ( .A1(n15710), .A2(n15709), .ZN(n15713) );
  OAI21_X1 U18958 ( .B1(P1_FLUSH_REG_SCAN_IN), .B2(P1_MORE_REG_SCAN_IN), .A(
        n15711), .ZN(n15712) );
  NAND4_X1 U18959 ( .A1(n15715), .A2(n15714), .A3(n15713), .A4(n15712), .ZN(
        n15716) );
  OAI21_X1 U18960 ( .B1(n15717), .B2(n15716), .A(n16000), .ZN(n15720) );
  AOI21_X1 U18961 ( .B1(n15996), .B2(n15720), .A(n11192), .ZN(n20692) );
  OAI211_X1 U18962 ( .C1(P1_STATE2_REG_2__SCAN_IN), .C2(n15993), .A(n20692), 
        .B(n15718), .ZN(n15999) );
  OAI21_X1 U18963 ( .B1(n20691), .B2(n15720), .A(n15719), .ZN(n15721) );
  OAI22_X1 U18964 ( .A1(n15723), .A2(n15722), .B1(n15999), .B2(n15721), .ZN(
        n15724) );
  AOI21_X1 U18965 ( .B1(n15725), .B2(n15996), .A(n15724), .ZN(P1_U3161) );
  INV_X1 U18966 ( .A(n16298), .ZN(n15728) );
  NAND2_X1 U18967 ( .A1(n15728), .A2(n16299), .ZN(n15729) );
  NAND2_X1 U18968 ( .A1(n15729), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16301) );
  OAI21_X1 U18969 ( .B1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n15729), .A(
        n16301), .ZN(n16327) );
  NOR2_X1 U18970 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16349), .ZN(
        n16323) );
  OAI211_X1 U18971 ( .C1(n15730), .C2(n16349), .A(n16345), .B(n18073), .ZN(
        n16346) );
  INV_X1 U18972 ( .A(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n16348) );
  AOI21_X1 U18973 ( .B1(n15731), .B2(n16346), .A(n16348), .ZN(n15732) );
  AOI21_X1 U18974 ( .B1(n16323), .B2(n15733), .A(n15732), .ZN(n15734) );
  NAND2_X1 U18975 ( .A1(n9820), .A2(P3_REIP_REG_30__SCAN_IN), .ZN(n16319) );
  OAI211_X1 U18976 ( .C1(n17909), .C2(n16327), .A(n15734), .B(n16319), .ZN(
        P3_U2832) );
  INV_X1 U18977 ( .A(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n20960) );
  NOR2_X1 U18978 ( .A1(n20699), .A2(n20960), .ZN(n15735) );
  INV_X1 U18979 ( .A(HOLD), .ZN(n20700) );
  OAI222_X1 U18980 ( .A1(n15735), .A2(P1_STATE_REG_1__SCAN_IN), .B1(n15735), 
        .B2(HOLD), .C1(n20700), .C2(n11119), .ZN(n15737) );
  NAND2_X1 U18981 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(n20791), .ZN(n20698) );
  NAND3_X1 U18982 ( .A1(n15737), .A2(n15736), .A3(n20698), .ZN(P1_U3195) );
  AND2_X1 U18983 ( .A1(n19978), .A2(P1_DATAO_REG_31__SCAN_IN), .ZN(P1_U2905)
         );
  NOR2_X1 U18984 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n15740) );
  NOR2_X1 U18985 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(P2_STATE2_REG_1__SCAN_IN), .ZN(n15739) );
  NAND2_X1 U18986 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19842), .ZN(n19710) );
  OAI21_X1 U18987 ( .B1(n19710), .B2(n19849), .A(n16295), .ZN(n15738) );
  AOI211_X1 U18988 ( .C1(n15740), .C2(n19836), .A(n15739), .B(n15738), .ZN(
        P2_U3178) );
  INV_X1 U18989 ( .A(n19830), .ZN(n16278) );
  OAI221_X1 U18990 ( .B1(n15741), .B2(n16295), .C1(n16278), .C2(n16295), .A(
        n19613), .ZN(n19822) );
  NOR2_X1 U18991 ( .A1(n20934), .A2(n19822), .ZN(P2_U3047) );
  NAND3_X1 U18992 ( .A1(n18094), .A2(n18100), .A3(n15742), .ZN(n15743) );
  NAND2_X1 U18993 ( .A1(n18134), .A2(n17111), .ZN(n17155) );
  INV_X1 U18994 ( .A(P3_EAX_REG_0__SCAN_IN), .ZN(n17310) );
  NAND2_X1 U18995 ( .A1(n15745), .A2(n17111), .ZN(n17243) );
  AOI22_X1 U18996 ( .A1(n17255), .A2(BUF2_REG_0__SCAN_IN), .B1(n17245), .B2(
        n15746), .ZN(n15747) );
  OAI221_X1 U18997 ( .B1(P3_EAX_REG_0__SCAN_IN), .B2(n17155), .C1(n17310), 
        .C2(n17111), .A(n15747), .ZN(P3_U2735) );
  INV_X1 U18998 ( .A(P1_REIP_REG_25__SCAN_IN), .ZN(n15752) );
  AOI21_X1 U18999 ( .B1(n15781), .B2(n15761), .A(n15780), .ZN(n15778) );
  OAI21_X1 U19000 ( .B1(P1_REIP_REG_24__SCAN_IN), .B2(n19892), .A(n15778), 
        .ZN(n15751) );
  OAI22_X1 U19001 ( .A1(n19934), .A2(n15749), .B1(n19954), .B2(n15748), .ZN(
        n15750) );
  AOI221_X1 U19002 ( .B1(n15753), .B2(n15752), .C1(n15751), .C2(
        P1_REIP_REG_25__SCAN_IN), .A(n15750), .ZN(n15759) );
  INV_X1 U19003 ( .A(n15754), .ZN(n15755) );
  OAI22_X1 U19004 ( .A1(n15756), .A2(n15796), .B1(n15755), .B2(n19953), .ZN(
        n15757) );
  INV_X1 U19005 ( .A(n15757), .ZN(n15758) );
  OAI211_X1 U19006 ( .C1(n15760), .C2(n19937), .A(n15759), .B(n15758), .ZN(
        P1_U2815) );
  OAI22_X1 U19007 ( .A1(n19954), .A2(n12344), .B1(n15778), .B2(n20739), .ZN(
        n15763) );
  NOR3_X1 U19008 ( .A1(n19892), .A2(P1_REIP_REG_24__SCAN_IN), .A3(n15761), 
        .ZN(n15762) );
  AOI211_X1 U19009 ( .C1(P1_EBX_REG_24__SCAN_IN), .C2(n19955), .A(n15763), .B(
        n15762), .ZN(n15768) );
  INV_X1 U19010 ( .A(n15764), .ZN(n15765) );
  AOI22_X1 U19011 ( .A1(n15766), .A2(n19908), .B1(n15765), .B2(n19951), .ZN(
        n15767) );
  OAI211_X1 U19012 ( .C1(n15769), .C2(n19953), .A(n15768), .B(n15767), .ZN(
        P1_U2816) );
  AND2_X1 U19013 ( .A1(n15781), .A2(n15779), .ZN(n15803) );
  AOI21_X1 U19014 ( .B1(n15770), .B2(n15803), .A(P1_REIP_REG_23__SCAN_IN), 
        .ZN(n15777) );
  AOI22_X1 U19015 ( .A1(n19955), .A2(P1_EBX_REG_23__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n19932), .ZN(n15776) );
  OAI22_X1 U19016 ( .A1(n15772), .A2(n15796), .B1(n19937), .B2(n15771), .ZN(
        n15773) );
  AOI21_X1 U19017 ( .B1(n15774), .B2(n19941), .A(n15773), .ZN(n15775) );
  OAI211_X1 U19018 ( .C1(n15778), .C2(n15777), .A(n15776), .B(n15775), .ZN(
        P1_U2817) );
  NAND2_X1 U19019 ( .A1(n15779), .A2(P1_REIP_REG_20__SCAN_IN), .ZN(n15792) );
  OAI21_X1 U19020 ( .B1(n15780), .B2(n15792), .A(n19952), .ZN(n15804) );
  INV_X1 U19021 ( .A(P1_REIP_REG_21__SCAN_IN), .ZN(n15793) );
  NAND2_X1 U19022 ( .A1(n15781), .A2(n15793), .ZN(n15791) );
  AOI21_X1 U19023 ( .B1(n15804), .B2(n15791), .A(n20736), .ZN(n15788) );
  NAND2_X1 U19024 ( .A1(n15803), .A2(n20736), .ZN(n15783) );
  NOR2_X1 U19025 ( .A1(n15783), .A2(n15782), .ZN(n15787) );
  INV_X1 U19026 ( .A(P1_EBX_REG_22__SCAN_IN), .ZN(n15785) );
  INV_X1 U19027 ( .A(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n15784) );
  OAI22_X1 U19028 ( .A1(n19934), .A2(n15785), .B1(n15784), .B2(n19954), .ZN(
        n15786) );
  NOR3_X1 U19029 ( .A1(n15788), .A2(n15787), .A3(n15786), .ZN(n15790) );
  AOI22_X1 U19030 ( .A1(n15862), .A2(n19908), .B1(n19951), .B2(n15927), .ZN(
        n15789) );
  OAI211_X1 U19031 ( .C1(n15865), .C2(n19953), .A(n15790), .B(n15789), .ZN(
        P1_U2818) );
  OAI22_X1 U19032 ( .A1(n15804), .A2(n15793), .B1(n15792), .B2(n15791), .ZN(
        n15794) );
  AOI21_X1 U19033 ( .B1(n19955), .B2(P1_EBX_REG_21__SCAN_IN), .A(n15794), .ZN(
        n15801) );
  OAI22_X1 U19034 ( .A1(n15797), .A2(n15796), .B1(n19937), .B2(n15795), .ZN(
        n15798) );
  AOI21_X1 U19035 ( .B1(n15799), .B2(n19941), .A(n15798), .ZN(n15800) );
  OAI211_X1 U19036 ( .C1(n15802), .C2(n19954), .A(n15801), .B(n15800), .ZN(
        P1_U2819) );
  NOR2_X1 U19037 ( .A1(P1_REIP_REG_20__SCAN_IN), .A2(n15803), .ZN(n15805) );
  OAI22_X1 U19038 ( .A1(n15805), .A2(n15804), .B1(n15854), .B2(n19934), .ZN(
        n15806) );
  AOI21_X1 U19039 ( .B1(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n19932), .A(
        n15806), .ZN(n15809) );
  INV_X1 U19040 ( .A(n15807), .ZN(n15852) );
  AOI22_X1 U19041 ( .A1(n15868), .A2(n19908), .B1(n19951), .B2(n15852), .ZN(
        n15808) );
  OAI211_X1 U19042 ( .C1(n15866), .C2(n19953), .A(n15809), .B(n15808), .ZN(
        P1_U2820) );
  OAI22_X1 U19043 ( .A1(n19934), .A2(n15811), .B1(n19954), .B2(n15810), .ZN(
        n15812) );
  AOI211_X1 U19044 ( .C1(n19941), .C2(n15813), .A(n15986), .B(n15812), .ZN(
        n15819) );
  OAI21_X1 U19045 ( .B1(n15814), .B2(n15827), .A(n14656), .ZN(n15815) );
  AOI22_X1 U19046 ( .A1(n15817), .A2(n19908), .B1(n15816), .B2(n15815), .ZN(
        n15818) );
  OAI211_X1 U19047 ( .C1(n19937), .C2(n15820), .A(n15819), .B(n15818), .ZN(
        P1_U2823) );
  INV_X1 U19048 ( .A(P1_REIP_REG_16__SCAN_IN), .ZN(n15944) );
  NAND2_X1 U19049 ( .A1(P1_REIP_REG_15__SCAN_IN), .A2(n15944), .ZN(n15826) );
  AOI22_X1 U19050 ( .A1(n15934), .A2(n19951), .B1(n19955), .B2(
        P1_EBX_REG_16__SCAN_IN), .ZN(n15821) );
  OAI21_X1 U19051 ( .B1(n15879), .B2(n19953), .A(n15821), .ZN(n15822) );
  AOI211_X1 U19052 ( .C1(n19932), .C2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .A(
        n15986), .B(n15822), .ZN(n15825) );
  OAI21_X1 U19053 ( .B1(P1_REIP_REG_15__SCAN_IN), .B2(n15827), .A(n15837), 
        .ZN(n15823) );
  AOI22_X1 U19054 ( .A1(n15876), .A2(n19908), .B1(P1_REIP_REG_16__SCAN_IN), 
        .B2(n15823), .ZN(n15824) );
  OAI211_X1 U19055 ( .C1(n15827), .C2(n15826), .A(n15825), .B(n15824), .ZN(
        P1_U2824) );
  INV_X1 U19056 ( .A(P1_REIP_REG_13__SCAN_IN), .ZN(n21083) );
  NOR2_X1 U19057 ( .A1(n21083), .A2(n15828), .ZN(n15829) );
  AOI21_X1 U19058 ( .B1(n15829), .B2(n15849), .A(P1_REIP_REG_14__SCAN_IN), 
        .ZN(n15836) );
  OAI21_X1 U19059 ( .B1(n19954), .B2(n15830), .A(n20046), .ZN(n15833) );
  NOR2_X1 U19060 ( .A1(n19937), .A2(n15831), .ZN(n15832) );
  AOI211_X1 U19061 ( .C1(P1_EBX_REG_14__SCAN_IN), .C2(n19955), .A(n15833), .B(
        n15832), .ZN(n15835) );
  AOI22_X1 U19062 ( .A1(n15881), .A2(n19908), .B1(n19941), .B2(n15880), .ZN(
        n15834) );
  OAI211_X1 U19063 ( .C1(n15837), .C2(n15836), .A(n15835), .B(n15834), .ZN(
        P1_U2826) );
  AOI22_X1 U19064 ( .A1(n19955), .A2(P1_EBX_REG_12__SCAN_IN), .B1(
        P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n19932), .ZN(n15843) );
  AOI21_X1 U19065 ( .B1(n15855), .B2(n19951), .A(n15986), .ZN(n15842) );
  INV_X1 U19066 ( .A(n15838), .ZN(n15885) );
  AOI22_X1 U19067 ( .A1(n15886), .A2(n19941), .B1(n19908), .B2(n15885), .ZN(
        n15841) );
  OAI221_X1 U19068 ( .B1(P1_REIP_REG_12__SCAN_IN), .B2(P1_REIP_REG_11__SCAN_IN), .C1(P1_REIP_REG_12__SCAN_IN), .C2(n15849), .A(n15839), .ZN(n15840) );
  NAND4_X1 U19069 ( .A1(n15843), .A2(n15842), .A3(n15841), .A4(n15840), .ZN(
        P1_U2828) );
  INV_X1 U19070 ( .A(P1_REIP_REG_11__SCAN_IN), .ZN(n15848) );
  INV_X1 U19071 ( .A(n15844), .ZN(n15945) );
  AOI22_X1 U19072 ( .A1(n19955), .A2(P1_EBX_REG_11__SCAN_IN), .B1(n19951), 
        .B2(n15945), .ZN(n15845) );
  OAI21_X1 U19073 ( .B1(n15846), .B2(n15848), .A(n15845), .ZN(n15847) );
  AOI211_X1 U19074 ( .C1(n19932), .C2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n15986), .B(n15847), .ZN(n15851) );
  AOI22_X1 U19075 ( .A1(n15894), .A2(n19908), .B1(n15849), .B2(n15848), .ZN(
        n15850) );
  OAI211_X1 U19076 ( .C1(n15897), .C2(n19953), .A(n15851), .B(n15850), .ZN(
        P1_U2829) );
  AOI22_X1 U19077 ( .A1(n15868), .A2(n19964), .B1(n15856), .B2(n15852), .ZN(
        n15853) );
  OAI21_X1 U19078 ( .B1(n19968), .B2(n15854), .A(n15853), .ZN(P1_U2852) );
  AOI22_X1 U19079 ( .A1(n15885), .A2(n19964), .B1(n15856), .B2(n15855), .ZN(
        n15857) );
  OAI21_X1 U19080 ( .B1(n19968), .B2(n15858), .A(n15857), .ZN(P1_U2860) );
  AOI22_X1 U19081 ( .A1(n20038), .A2(P1_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        n15986), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15864) );
  NAND2_X1 U19082 ( .A1(n15860), .A2(n15859), .ZN(n15861) );
  XNOR2_X1 U19083 ( .A(n15861), .B(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(
        n15928) );
  AOI22_X1 U19084 ( .A1(n15862), .A2(n20101), .B1(n20043), .B2(n15928), .ZN(
        n15863) );
  OAI211_X1 U19085 ( .C1(n15909), .C2(n15865), .A(n15864), .B(n15863), .ZN(
        P1_U2977) );
  AOI22_X1 U19086 ( .A1(n20038), .A2(P1_PHYADDRPOINTER_REG_20__SCAN_IN), .B1(
        n15986), .B2(P1_REIP_REG_20__SCAN_IN), .ZN(n15870) );
  INV_X1 U19087 ( .A(n15866), .ZN(n15867) );
  AOI22_X1 U19088 ( .A1(n15868), .A2(n20101), .B1(n15867), .B2(n15911), .ZN(
        n15869) );
  OAI211_X1 U19089 ( .C1(n15871), .C2(n19863), .A(n15870), .B(n15869), .ZN(
        P1_U2979) );
  AOI22_X1 U19090 ( .A1(n20038), .A2(P1_PHYADDRPOINTER_REG_16__SCAN_IN), .B1(
        n15986), .B2(P1_REIP_REG_16__SCAN_IN), .ZN(n15878) );
  OAI22_X1 U19091 ( .A1(n15873), .A2(n15872), .B1(n14636), .B2(
        P1_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n15874) );
  XOR2_X1 U19092 ( .A(n15875), .B(n15874), .Z(n15935) );
  AOI22_X1 U19093 ( .A1(n15935), .A2(n20043), .B1(n20101), .B2(n15876), .ZN(
        n15877) );
  OAI211_X1 U19094 ( .C1(n15909), .C2(n15879), .A(n15878), .B(n15877), .ZN(
        P1_U2983) );
  AOI22_X1 U19095 ( .A1(n20038), .A2(P1_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        n15986), .B2(P1_REIP_REG_14__SCAN_IN), .ZN(n15883) );
  AOI22_X1 U19096 ( .A1(n15881), .A2(n20101), .B1(n15911), .B2(n15880), .ZN(
        n15882) );
  OAI211_X1 U19097 ( .C1(n15884), .C2(n19863), .A(n15883), .B(n15882), .ZN(
        P1_U2985) );
  AOI22_X1 U19098 ( .A1(n20038), .A2(P1_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        n15986), .B2(P1_REIP_REG_12__SCAN_IN), .ZN(n15888) );
  AOI22_X1 U19099 ( .A1(n15911), .A2(n15886), .B1(n20101), .B2(n15885), .ZN(
        n15887) );
  OAI211_X1 U19100 ( .C1(n15889), .C2(n19863), .A(n15888), .B(n15887), .ZN(
        P1_U2987) );
  AOI22_X1 U19101 ( .A1(n20038), .A2(P1_PHYADDRPOINTER_REG_11__SCAN_IN), .B1(
        n15986), .B2(P1_REIP_REG_11__SCAN_IN), .ZN(n15896) );
  NAND3_X1 U19102 ( .A1(n15890), .A2(n14688), .A3(
        P1_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n15892) );
  NAND2_X1 U19103 ( .A1(n15892), .A2(n15891), .ZN(n15893) );
  XOR2_X1 U19104 ( .A(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B(n15893), .Z(
        n15947) );
  AOI22_X1 U19105 ( .A1(n20043), .A2(n15947), .B1(n20101), .B2(n15894), .ZN(
        n15895) );
  OAI211_X1 U19106 ( .C1(n15909), .C2(n15897), .A(n15896), .B(n15895), .ZN(
        P1_U2988) );
  AOI22_X1 U19107 ( .A1(n20038), .A2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .B1(
        n15986), .B2(P1_REIP_REG_7__SCAN_IN), .ZN(n15902) );
  XNOR2_X1 U19108 ( .A(n15899), .B(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(
        n15900) );
  XNOR2_X1 U19109 ( .A(n15898), .B(n15900), .ZN(n15977) );
  AOI22_X1 U19110 ( .A1(n15977), .A2(n20043), .B1(n20101), .B2(n19897), .ZN(
        n15901) );
  OAI211_X1 U19111 ( .C1(n15909), .C2(n19901), .A(n15902), .B(n15901), .ZN(
        P1_U2992) );
  AOI22_X1 U19112 ( .A1(n20038), .A2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        n15986), .B2(P1_REIP_REG_6__SCAN_IN), .ZN(n15908) );
  NAND2_X1 U19113 ( .A1(n15904), .A2(n15903), .ZN(n15905) );
  XNOR2_X1 U19114 ( .A(n15906), .B(n15905), .ZN(n15989) );
  AOI22_X1 U19115 ( .A1(n15989), .A2(n20043), .B1(n20101), .B2(n19965), .ZN(
        n15907) );
  OAI211_X1 U19116 ( .C1(n15909), .C2(n19906), .A(n15908), .B(n15907), .ZN(
        P1_U2993) );
  AOI222_X1 U19117 ( .A1(n15912), .A2(n15911), .B1(n20101), .B2(n19918), .C1(
        n20043), .C2(n15910), .ZN(n15914) );
  OAI211_X1 U19118 ( .C1(n15916), .C2(n15915), .A(n15914), .B(n15913), .ZN(
        P1_U2994) );
  INV_X1 U19119 ( .A(n15917), .ZN(n15919) );
  AOI22_X1 U19120 ( .A1(n15919), .A2(n20077), .B1(n20089), .B2(n15918), .ZN(
        n15924) );
  OAI22_X1 U19121 ( .A1(P1_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n15922), .B1(
        n15921), .B2(n15920), .ZN(n15923) );
  OAI211_X1 U19122 ( .C1(n15925), .C2(n20046), .A(n15924), .B(n15923), .ZN(
        P1_U3005) );
  AOI22_X1 U19123 ( .A1(P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n15926), .B1(
        n15986), .B2(P1_REIP_REG_22__SCAN_IN), .ZN(n15933) );
  AOI22_X1 U19124 ( .A1(n15928), .A2(n20077), .B1(n20089), .B2(n15927), .ZN(
        n15932) );
  OAI211_X1 U19125 ( .C1(P1_INSTADDRPOINTER_REG_21__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_22__SCAN_IN), .A(n15930), .B(n15929), .ZN(
        n15931) );
  NAND3_X1 U19126 ( .A1(n15933), .A2(n15932), .A3(n15931), .ZN(P1_U3009) );
  AOI22_X1 U19127 ( .A1(n15935), .A2(n20077), .B1(n20089), .B2(n15934), .ZN(
        n15943) );
  INV_X1 U19128 ( .A(n15936), .ZN(n15940) );
  OAI22_X1 U19129 ( .A1(n15940), .A2(n15939), .B1(n15938), .B2(n15937), .ZN(
        n15941) );
  OAI21_X1 U19130 ( .B1(P1_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(
        P1_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n15941), .ZN(n15942) );
  OAI211_X1 U19131 ( .C1(n15944), .C2(n20046), .A(n15943), .B(n15942), .ZN(
        P1_U3015) );
  AOI22_X1 U19132 ( .A1(n15945), .A2(n20089), .B1(n15986), .B2(
        P1_REIP_REG_11__SCAN_IN), .ZN(n15949) );
  AOI22_X1 U19133 ( .A1(n15947), .A2(n20077), .B1(
        P1_INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n15946), .ZN(n15948) );
  OAI211_X1 U19134 ( .C1(P1_INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n15950), .A(
        n15949), .B(n15948), .ZN(P1_U3020) );
  AOI21_X1 U19135 ( .B1(n20089), .B2(n15952), .A(n15951), .ZN(n15959) );
  AOI21_X1 U19136 ( .B1(n15960), .B2(n15954), .A(n15953), .ZN(n15956) );
  AOI22_X1 U19137 ( .A1(n15957), .A2(n20077), .B1(n15956), .B2(n15955), .ZN(
        n15958) );
  OAI211_X1 U19138 ( .C1(n15961), .C2(n15960), .A(n15959), .B(n15958), .ZN(
        P1_U3021) );
  INV_X1 U19139 ( .A(n15962), .ZN(n15964) );
  OAI21_X1 U19140 ( .B1(n14738), .B2(n15964), .A(n15963), .ZN(n15988) );
  AOI21_X1 U19141 ( .B1(n15974), .B2(n20076), .A(n15988), .ZN(n15979) );
  INV_X1 U19142 ( .A(n15965), .ZN(n15966) );
  AOI21_X1 U19143 ( .B1(n20089), .B2(n15967), .A(n15966), .ZN(n15972) );
  NAND2_X1 U19144 ( .A1(P1_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        P1_INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n15969) );
  AOI211_X1 U19145 ( .C1(n15973), .C2(n15980), .A(n15974), .B(n15992), .ZN(
        n15968) );
  AOI22_X1 U19146 ( .A1(n15970), .A2(n20077), .B1(n15969), .B2(n15968), .ZN(
        n15971) );
  OAI211_X1 U19147 ( .C1(n15979), .C2(n15973), .A(n15972), .B(n15971), .ZN(
        P1_U3023) );
  OR2_X1 U19148 ( .A1(n15974), .A2(n15992), .ZN(n15981) );
  OAI22_X1 U19149 ( .A1(n15975), .A2(n19895), .B1(n20717), .B2(n20046), .ZN(
        n15976) );
  AOI21_X1 U19150 ( .B1(n15977), .B2(n20077), .A(n15976), .ZN(n15978) );
  OAI221_X1 U19151 ( .B1(P1_INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n15981), .C1(
        n15980), .C2(n15979), .A(n15978), .ZN(P1_U3024) );
  OR2_X1 U19152 ( .A1(n15983), .A2(n15982), .ZN(n15984) );
  NAND2_X1 U19153 ( .A1(n15985), .A2(n15984), .ZN(n19961) );
  INV_X1 U19154 ( .A(n19961), .ZN(n15987) );
  AOI22_X1 U19155 ( .A1(n20089), .A2(n15987), .B1(n15986), .B2(
        P1_REIP_REG_6__SCAN_IN), .ZN(n15991) );
  AOI22_X1 U19156 ( .A1(n15989), .A2(n20077), .B1(
        P1_INSTADDRPOINTER_REG_6__SCAN_IN), .B2(n15988), .ZN(n15990) );
  OAI211_X1 U19157 ( .C1(P1_INSTADDRPOINTER_REG_6__SCAN_IN), .C2(n15992), .A(
        n15991), .B(n15990), .ZN(P1_U3025) );
  NAND4_X1 U19158 ( .A1(P1_STATE2_REG_0__SCAN_IN), .A2(
        P1_STATE2_REG_1__SCAN_IN), .A3(n20691), .A4(n15993), .ZN(n15994) );
  AND2_X1 U19159 ( .A1(n15995), .A2(n15994), .ZN(n20690) );
  AOI21_X1 U19160 ( .B1(n20690), .B2(n15997), .A(n15996), .ZN(n15998) );
  AOI21_X1 U19161 ( .B1(n16000), .B2(n15999), .A(n15998), .ZN(P1_U3162) );
  OAI21_X1 U19162 ( .B1(n20692), .B2(n20388), .A(n16001), .ZN(P1_U3466) );
  INV_X1 U19163 ( .A(n16002), .ZN(n16032) );
  INV_X1 U19164 ( .A(n16003), .ZN(n16057) );
  INV_X1 U19165 ( .A(n16004), .ZN(n16078) );
  INV_X1 U19166 ( .A(n16005), .ZN(n16100) );
  NAND2_X1 U19167 ( .A1(n18929), .A2(n16006), .ZN(n16099) );
  NAND2_X1 U19168 ( .A1(n16100), .A2(n16099), .ZN(n16098) );
  NAND2_X1 U19169 ( .A1(n18929), .A2(n16098), .ZN(n16088) );
  NAND2_X1 U19170 ( .A1(n16089), .A2(n16088), .ZN(n16087) );
  NAND2_X1 U19171 ( .A1(n18929), .A2(n16087), .ZN(n16077) );
  NAND2_X1 U19172 ( .A1(n16078), .A2(n16077), .ZN(n16076) );
  NAND2_X1 U19173 ( .A1(n18929), .A2(n16076), .ZN(n16067) );
  NAND2_X1 U19174 ( .A1(n16068), .A2(n16067), .ZN(n16066) );
  NAND2_X1 U19175 ( .A1(n18929), .A2(n16066), .ZN(n16056) );
  NAND2_X1 U19176 ( .A1(n16057), .A2(n16056), .ZN(n16055) );
  NAND2_X1 U19177 ( .A1(n18929), .A2(n16055), .ZN(n16043) );
  NAND2_X1 U19178 ( .A1(n16044), .A2(n16043), .ZN(n16042) );
  NAND2_X1 U19179 ( .A1(n18929), .A2(n16042), .ZN(n16031) );
  NAND2_X1 U19180 ( .A1(n16032), .A2(n16031), .ZN(n16030) );
  NAND2_X1 U19181 ( .A1(n18929), .A2(n16030), .ZN(n16020) );
  NAND2_X1 U19182 ( .A1(n16021), .A2(n16020), .ZN(n16019) );
  AOI22_X1 U19183 ( .A1(P2_PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n18958), .B1(
        P2_REIP_REG_31__SCAN_IN), .B2(n18885), .ZN(n16009) );
  NAND3_X1 U19184 ( .A1(n19081), .A2(P2_EBX_REG_31__SCAN_IN), .A3(n16007), 
        .ZN(n16008) );
  OAI211_X1 U19185 ( .C1(n16010), .C2(n18947), .A(n16009), .B(n16008), .ZN(
        n16011) );
  INV_X1 U19186 ( .A(n16011), .ZN(n16015) );
  INV_X1 U19187 ( .A(n16012), .ZN(n18961) );
  AOI22_X1 U19188 ( .A1(n16013), .A2(n18949), .B1(n18877), .B2(n18961), .ZN(
        n16014) );
  OAI211_X1 U19189 ( .C1(n18852), .C2(n16019), .A(n16015), .B(n16014), .ZN(
        P2_U2824) );
  AOI22_X1 U19190 ( .A1(P2_PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n18958), .B1(
        P2_REIP_REG_30__SCAN_IN), .B2(n18885), .ZN(n16025) );
  AOI22_X1 U19191 ( .A1(n16016), .A2(n18933), .B1(P2_EBX_REG_30__SCAN_IN), 
        .B2(n18951), .ZN(n16024) );
  AOI22_X1 U19192 ( .A1(n16018), .A2(n18949), .B1(n18877), .B2(n16017), .ZN(
        n16023) );
  OAI211_X1 U19193 ( .C1(n16021), .C2(n16020), .A(n18890), .B(n16019), .ZN(
        n16022) );
  NAND4_X1 U19194 ( .A1(n16025), .A2(n16024), .A3(n16023), .A4(n16022), .ZN(
        P2_U2825) );
  AOI22_X1 U19195 ( .A1(P2_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n18958), .B1(
        P2_REIP_REG_29__SCAN_IN), .B2(n18885), .ZN(n16036) );
  AOI22_X1 U19196 ( .A1(n16026), .A2(n18933), .B1(P2_EBX_REG_29__SCAN_IN), 
        .B2(n18951), .ZN(n16035) );
  OAI22_X1 U19197 ( .A1(n16028), .A2(n18937), .B1(n16027), .B2(n18945), .ZN(
        n16029) );
  INV_X1 U19198 ( .A(n16029), .ZN(n16034) );
  OAI211_X1 U19199 ( .C1(n16032), .C2(n16031), .A(n18890), .B(n16030), .ZN(
        n16033) );
  NAND4_X1 U19200 ( .A1(n16036), .A2(n16035), .A3(n16034), .A4(n16033), .ZN(
        P2_U2826) );
  AOI22_X1 U19201 ( .A1(P2_PHYADDRPOINTER_REG_28__SCAN_IN), .A2(n18958), .B1(
        P2_REIP_REG_28__SCAN_IN), .B2(n18885), .ZN(n16038) );
  NAND2_X1 U19202 ( .A1(n18951), .A2(P2_EBX_REG_28__SCAN_IN), .ZN(n16037) );
  OAI211_X1 U19203 ( .C1(n16039), .C2(n18947), .A(n16038), .B(n16037), .ZN(
        n16040) );
  AOI21_X1 U19204 ( .B1(n16041), .B2(n18949), .A(n16040), .ZN(n16046) );
  OAI211_X1 U19205 ( .C1(n16044), .C2(n16043), .A(n18890), .B(n16042), .ZN(
        n16045) );
  OAI211_X1 U19206 ( .C1(n18945), .C2(n16047), .A(n16046), .B(n16045), .ZN(
        P2_U2827) );
  INV_X1 U19207 ( .A(n16048), .ZN(n16054) );
  OAI22_X1 U19208 ( .A1(n16049), .A2(n18831), .B1(n19767), .B2(n18954), .ZN(
        n16050) );
  AOI21_X1 U19209 ( .B1(n18951), .B2(P2_EBX_REG_27__SCAN_IN), .A(n16050), .ZN(
        n16051) );
  OAI21_X1 U19210 ( .B1(n16052), .B2(n18947), .A(n16051), .ZN(n16053) );
  AOI21_X1 U19211 ( .B1(n16054), .B2(n18949), .A(n16053), .ZN(n16059) );
  OAI211_X1 U19212 ( .C1(n16057), .C2(n16056), .A(n18890), .B(n16055), .ZN(
        n16058) );
  OAI211_X1 U19213 ( .C1(n18945), .C2(n16060), .A(n16059), .B(n16058), .ZN(
        P2_U2828) );
  AOI22_X1 U19214 ( .A1(P2_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n18958), .B1(
        P2_REIP_REG_26__SCAN_IN), .B2(n18885), .ZN(n16072) );
  INV_X1 U19215 ( .A(P2_EBX_REG_26__SCAN_IN), .ZN(n16061) );
  OAI22_X1 U19216 ( .A1(n16062), .A2(n18947), .B1(n18840), .B2(n16061), .ZN(
        n16063) );
  INV_X1 U19217 ( .A(n16063), .ZN(n16071) );
  AOI22_X1 U19218 ( .A1(n16065), .A2(n18949), .B1(n16064), .B2(n18877), .ZN(
        n16070) );
  OAI211_X1 U19219 ( .C1(n16068), .C2(n16067), .A(n18890), .B(n16066), .ZN(
        n16069) );
  NAND4_X1 U19220 ( .A1(n16072), .A2(n16071), .A3(n16070), .A4(n16069), .ZN(
        P2_U2829) );
  AOI22_X1 U19221 ( .A1(P2_PHYADDRPOINTER_REG_25__SCAN_IN), .A2(n18958), .B1(
        P2_REIP_REG_25__SCAN_IN), .B2(n18885), .ZN(n16082) );
  AOI22_X1 U19222 ( .A1(n16073), .A2(n18933), .B1(P2_EBX_REG_25__SCAN_IN), 
        .B2(n18951), .ZN(n16081) );
  AOI22_X1 U19223 ( .A1(n16075), .A2(n18949), .B1(n18877), .B2(n16074), .ZN(
        n16080) );
  OAI211_X1 U19224 ( .C1(n16078), .C2(n16077), .A(n18890), .B(n16076), .ZN(
        n16079) );
  NAND4_X1 U19225 ( .A1(n16082), .A2(n16081), .A3(n16080), .A4(n16079), .ZN(
        P2_U2830) );
  AOI22_X1 U19226 ( .A1(P2_PHYADDRPOINTER_REG_24__SCAN_IN), .A2(n18958), .B1(
        P2_REIP_REG_24__SCAN_IN), .B2(n18885), .ZN(n16093) );
  AOI22_X1 U19227 ( .A1(n16083), .A2(n18933), .B1(P2_EBX_REG_24__SCAN_IN), 
        .B2(n18951), .ZN(n16092) );
  OAI22_X1 U19228 ( .A1(n16085), .A2(n18937), .B1(n16084), .B2(n18945), .ZN(
        n16086) );
  INV_X1 U19229 ( .A(n16086), .ZN(n16091) );
  OAI211_X1 U19230 ( .C1(n16089), .C2(n16088), .A(n18890), .B(n16087), .ZN(
        n16090) );
  NAND4_X1 U19231 ( .A1(n16093), .A2(n16092), .A3(n16091), .A4(n16090), .ZN(
        P2_U2831) );
  AOI22_X1 U19232 ( .A1(P2_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n18958), .B1(
        P2_REIP_REG_23__SCAN_IN), .B2(n18885), .ZN(n16104) );
  AOI22_X1 U19233 ( .A1(n16094), .A2(n18933), .B1(P2_EBX_REG_23__SCAN_IN), 
        .B2(n18951), .ZN(n16103) );
  INV_X1 U19234 ( .A(n16095), .ZN(n16097) );
  AOI22_X1 U19235 ( .A1(n16097), .A2(n18949), .B1(n16096), .B2(n18877), .ZN(
        n16102) );
  OAI211_X1 U19236 ( .C1(n16100), .C2(n16099), .A(n18890), .B(n16098), .ZN(
        n16101) );
  NAND4_X1 U19237 ( .A1(n16104), .A2(n16103), .A3(n16102), .A4(n16101), .ZN(
        P2_U2832) );
  INV_X1 U19238 ( .A(n19140), .ZN(n16105) );
  AOI22_X1 U19239 ( .A1(n18965), .A2(n16105), .B1(n19004), .B2(
        P2_EAX_REG_22__SCAN_IN), .ZN(n16111) );
  AOI22_X1 U19240 ( .A1(n18967), .A2(BUF1_REG_22__SCAN_IN), .B1(n18966), .B2(
        BUF2_REG_22__SCAN_IN), .ZN(n16110) );
  OAI22_X1 U19241 ( .A1(n16107), .A2(n19009), .B1(n18969), .B2(n16106), .ZN(
        n16108) );
  INV_X1 U19242 ( .A(n16108), .ZN(n16109) );
  NAND3_X1 U19243 ( .A1(n16111), .A2(n16110), .A3(n16109), .ZN(P2_U2897) );
  AOI22_X1 U19244 ( .A1(n18965), .A2(n16112), .B1(P2_EAX_REG_20__SCAN_IN), 
        .B2(n19004), .ZN(n16117) );
  AOI22_X1 U19245 ( .A1(n18967), .A2(BUF1_REG_20__SCAN_IN), .B1(n18966), .B2(
        BUF2_REG_20__SCAN_IN), .ZN(n16116) );
  AOI22_X1 U19246 ( .A1(n16114), .A2(n16121), .B1(n19005), .B2(n16113), .ZN(
        n16115) );
  NAND3_X1 U19247 ( .A1(n16117), .A2(n16116), .A3(n16115), .ZN(P2_U2899) );
  AOI22_X1 U19248 ( .A1(n18965), .A2(n16118), .B1(P2_EAX_REG_18__SCAN_IN), 
        .B2(n19004), .ZN(n16125) );
  AOI22_X1 U19249 ( .A1(n18967), .A2(BUF1_REG_18__SCAN_IN), .B1(n18966), .B2(
        BUF2_REG_18__SCAN_IN), .ZN(n16124) );
  INV_X1 U19250 ( .A(n16119), .ZN(n16122) );
  INV_X1 U19251 ( .A(n18810), .ZN(n16120) );
  AOI22_X1 U19252 ( .A1(n16122), .A2(n16121), .B1(n19005), .B2(n16120), .ZN(
        n16123) );
  NAND3_X1 U19253 ( .A1(n16125), .A2(n16124), .A3(n16123), .ZN(P2_U2901) );
  AOI22_X1 U19254 ( .A1(n19086), .A2(P2_PHYADDRPOINTER_REG_22__SCAN_IN), .B1(
        P2_REIP_REG_22__SCAN_IN), .B2(n19085), .ZN(n16130) );
  AOI222_X1 U19255 ( .A1(n16128), .A2(n19087), .B1(n19104), .B2(n16127), .C1(
        n19102), .C2(n16126), .ZN(n16129) );
  OAI211_X1 U19256 ( .C1(n19098), .C2(n16131), .A(n16130), .B(n16129), .ZN(
        P2_U2992) );
  AOI22_X1 U19257 ( .A1(n19086), .A2(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B1(
        P2_REIP_REG_14__SCAN_IN), .B2(n19085), .ZN(n16137) );
  AOI21_X1 U19258 ( .B1(n16196), .B2(n15440), .A(n15247), .ZN(n16195) );
  NAND2_X1 U19259 ( .A1(n16133), .A2(n16132), .ZN(n16135) );
  XOR2_X1 U19260 ( .A(n16135), .B(n16134), .Z(n16194) );
  AOI222_X1 U19261 ( .A1(n16195), .A2(n19102), .B1(n19087), .B2(n16194), .C1(
        n19104), .C2(n16193), .ZN(n16136) );
  OAI211_X1 U19262 ( .C1(n19098), .C2(n16138), .A(n16137), .B(n16136), .ZN(
        P2_U3000) );
  AOI22_X1 U19263 ( .A1(P2_REIP_REG_13__SCAN_IN), .A2(n19085), .B1(n19101), 
        .B2(n18863), .ZN(n16143) );
  OAI22_X1 U19264 ( .A1(n16140), .A2(n19092), .B1(n19108), .B2(n16139), .ZN(
        n16141) );
  AOI21_X1 U19265 ( .B1(n19104), .B2(n18862), .A(n16141), .ZN(n16142) );
  OAI211_X1 U19266 ( .C1(n19113), .C2(n16144), .A(n16143), .B(n16142), .ZN(
        P2_U3001) );
  AOI22_X1 U19267 ( .A1(n19086), .A2(P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B1(
        P2_REIP_REG_12__SCAN_IN), .B2(n19085), .ZN(n16151) );
  NOR2_X1 U19268 ( .A1(n16174), .A2(n18874), .ZN(n16148) );
  NOR3_X1 U19269 ( .A1(n16146), .A2(n16145), .A3(n19092), .ZN(n16147) );
  AOI211_X1 U19270 ( .C1(n19087), .C2(n16149), .A(n16148), .B(n16147), .ZN(
        n16150) );
  OAI211_X1 U19271 ( .C1(n19098), .C2(n18869), .A(n16151), .B(n16150), .ZN(
        P2_U3002) );
  AOI22_X1 U19272 ( .A1(P2_REIP_REG_11__SCAN_IN), .A2(n19085), .B1(n19101), 
        .B2(n18888), .ZN(n16156) );
  OAI22_X1 U19273 ( .A1(n16153), .A2(n19092), .B1(n16152), .B2(n19108), .ZN(
        n16154) );
  AOI21_X1 U19274 ( .B1(n19104), .B2(n18889), .A(n16154), .ZN(n16155) );
  OAI211_X1 U19275 ( .C1(n19113), .C2(n16157), .A(n16156), .B(n16155), .ZN(
        P2_U3003) );
  AOI22_X1 U19276 ( .A1(n19086), .A2(P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B1(
        P2_REIP_REG_10__SCAN_IN), .B2(n19085), .ZN(n16163) );
  NOR3_X1 U19277 ( .A1(n16158), .A2(n9848), .A3(n19092), .ZN(n16161) );
  OAI22_X1 U19278 ( .A1(n16159), .A2(n19108), .B1(n16174), .B2(n18900), .ZN(
        n16160) );
  NOR2_X1 U19279 ( .A1(n16161), .A2(n16160), .ZN(n16162) );
  OAI211_X1 U19280 ( .C1(n19098), .C2(n18897), .A(n16163), .B(n16162), .ZN(
        P2_U3004) );
  AOI22_X1 U19281 ( .A1(n19086), .A2(P2_PHYADDRPOINTER_REG_8__SCAN_IN), .B1(
        P2_REIP_REG_8__SCAN_IN), .B2(n19085), .ZN(n16177) );
  INV_X1 U19282 ( .A(n16164), .ZN(n16165) );
  AOI21_X1 U19283 ( .B1(n14080), .B2(n16166), .A(n16165), .ZN(n16170) );
  NAND2_X1 U19284 ( .A1(n16168), .A2(n16167), .ZN(n16169) );
  XNOR2_X1 U19285 ( .A(n16170), .B(n16169), .ZN(n16218) );
  OAI21_X1 U19286 ( .B1(n16173), .B2(n16172), .A(n16171), .ZN(n16213) );
  OAI222_X1 U19287 ( .A1(n16211), .A2(n16174), .B1(n19108), .B2(n16218), .C1(
        n19092), .C2(n16213), .ZN(n16175) );
  INV_X1 U19288 ( .A(n16175), .ZN(n16176) );
  OAI211_X1 U19289 ( .C1(n19098), .C2(n16178), .A(n16177), .B(n16176), .ZN(
        P2_U3006) );
  AOI22_X1 U19290 ( .A1(n19086), .A2(P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B1(
        P2_REIP_REG_6__SCAN_IN), .B2(n19085), .ZN(n16184) );
  INV_X1 U19291 ( .A(n16179), .ZN(n16182) );
  AOI222_X1 U19292 ( .A1(n16182), .A2(n19102), .B1(n19087), .B2(n16181), .C1(
        n19104), .C2(n16180), .ZN(n16183) );
  OAI211_X1 U19293 ( .C1(n19098), .C2(n18919), .A(n16184), .B(n16183), .ZN(
        P2_U3008) );
  AOI22_X1 U19294 ( .A1(P2_REIP_REG_5__SCAN_IN), .A2(n19085), .B1(n19101), 
        .B2(n18930), .ZN(n16190) );
  OAI22_X1 U19295 ( .A1(n16186), .A2(n19092), .B1(n19108), .B2(n16185), .ZN(
        n16187) );
  AOI21_X1 U19296 ( .B1(n19104), .B2(n16188), .A(n16187), .ZN(n16189) );
  OAI211_X1 U19297 ( .C1(n19113), .C2(n16191), .A(n16190), .B(n16189), .ZN(
        P2_U3009) );
  AOI22_X1 U19298 ( .A1(n16192), .A2(P2_INSTADDRPOINTER_REG_14__SCAN_IN), .B1(
        n16209), .B2(n18975), .ZN(n16201) );
  AOI222_X1 U19299 ( .A1(n16195), .A2(n12618), .B1(n16227), .B2(n16194), .C1(
        n16219), .C2(n16193), .ZN(n16200) );
  NAND2_X1 U19300 ( .A1(P2_REIP_REG_14__SCAN_IN), .A2(n19085), .ZN(n16199) );
  NAND4_X1 U19301 ( .A1(P2_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        P2_INSTADDRPOINTER_REG_13__SCAN_IN), .A3(n16197), .A4(n16196), .ZN(
        n16198) );
  NAND4_X1 U19302 ( .A1(n16201), .A2(n16200), .A3(n16199), .A4(n16198), .ZN(
        P2_U3032) );
  NAND2_X1 U19303 ( .A1(P2_REIP_REG_8__SCAN_IN), .A2(n19085), .ZN(n16205) );
  OAI211_X1 U19304 ( .C1(P2_INSTADDRPOINTER_REG_8__SCAN_IN), .C2(
        P2_INSTADDRPOINTER_REG_7__SCAN_IN), .A(n16203), .B(n16202), .ZN(n16204) );
  OAI211_X1 U19305 ( .C1(n16207), .C2(n16206), .A(n16205), .B(n16204), .ZN(
        n16208) );
  AOI21_X1 U19306 ( .B1(n16210), .B2(n16209), .A(n16208), .ZN(n16216) );
  OAI22_X1 U19307 ( .A1(n16213), .A2(n16223), .B1(n16212), .B2(n16211), .ZN(
        n16214) );
  INV_X1 U19308 ( .A(n16214), .ZN(n16215) );
  OAI211_X1 U19309 ( .C1(n16218), .C2(n16217), .A(n16216), .B(n16215), .ZN(
        P2_U3038) );
  OAI211_X1 U19310 ( .C1(n18996), .C2(n16222), .A(n16221), .B(n16220), .ZN(
        n16226) );
  NOR2_X1 U19311 ( .A1(n16224), .A2(n16223), .ZN(n16225) );
  AOI211_X1 U19312 ( .C1(n16228), .C2(n16227), .A(n16226), .B(n16225), .ZN(
        n16229) );
  OAI221_X1 U19313 ( .B1(n16231), .B2(n10009), .C1(n16231), .C2(n16230), .A(
        n16229), .ZN(P2_U3043) );
  OR2_X1 U19314 ( .A1(n16245), .A2(n16268), .ZN(n16234) );
  NAND2_X1 U19315 ( .A1(n16268), .A2(n16232), .ZN(n16233) );
  NAND2_X1 U19316 ( .A1(n16234), .A2(n16233), .ZN(n16269) );
  INV_X1 U19317 ( .A(n16268), .ZN(n16243) );
  INV_X1 U19318 ( .A(n16238), .ZN(n16237) );
  MUX2_X1 U19319 ( .A(n16235), .B(P2_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(
        n16268), .Z(n16270) );
  INV_X1 U19320 ( .A(n16270), .ZN(n16236) );
  OR2_X1 U19321 ( .A1(n16236), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n16246) );
  AOI22_X1 U19322 ( .A1(n16237), .A2(n19470), .B1(
        P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n16246), .ZN(n16242) );
  OAI21_X1 U19323 ( .B1(n16238), .B2(n19823), .A(n19814), .ZN(n16239) );
  NAND2_X1 U19324 ( .A1(n16240), .A2(n16239), .ZN(n16241) );
  AND3_X1 U19325 ( .A1(n16243), .A2(n16242), .A3(n16241), .ZN(n16244) );
  OAI21_X1 U19326 ( .B1(n16245), .B2(n19796), .A(n16244), .ZN(n16250) );
  INV_X1 U19327 ( .A(n16246), .ZN(n16247) );
  NAND2_X1 U19328 ( .A1(n16248), .A2(n16247), .ZN(n16249) );
  OAI211_X1 U19329 ( .C1(n16269), .C2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n16250), .B(n16249), .ZN(n16251) );
  NAND2_X1 U19330 ( .A1(n16251), .A2(n20934), .ZN(n16274) );
  OR2_X1 U19331 ( .A1(n16257), .A2(n16252), .ZN(n16260) );
  INV_X1 U19332 ( .A(n16253), .ZN(n16254) );
  NAND2_X1 U19333 ( .A1(n16255), .A2(n16254), .ZN(n16259) );
  NAND2_X1 U19334 ( .A1(n16257), .A2(n16256), .ZN(n16258) );
  AND3_X1 U19335 ( .A1(n16260), .A2(n16259), .A3(n16258), .ZN(n19832) );
  INV_X1 U19336 ( .A(P2_MORE_REG_SCAN_IN), .ZN(n16261) );
  NAND2_X1 U19337 ( .A1(n15741), .A2(n16261), .ZN(n16264) );
  OAI21_X1 U19338 ( .B1(n10842), .B2(n19838), .A(n16262), .ZN(n16263) );
  AOI21_X1 U19339 ( .B1(n16265), .B2(n16264), .A(n16263), .ZN(n16266) );
  NAND2_X1 U19340 ( .A1(n19832), .A2(n16266), .ZN(n16267) );
  AOI21_X1 U19341 ( .B1(n16268), .B2(P2_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A(
        n16267), .ZN(n16273) );
  INV_X1 U19342 ( .A(n16269), .ZN(n16271) );
  NAND2_X1 U19343 ( .A1(n16271), .A2(n16270), .ZN(n16272) );
  NOR2_X1 U19344 ( .A1(n19849), .A2(n19710), .ZN(n16275) );
  AOI211_X1 U19345 ( .C1(n16278), .C2(n16277), .A(n16276), .B(n16275), .ZN(
        n16291) );
  NAND2_X1 U19346 ( .A1(n16293), .A2(n15527), .ZN(n16279) );
  NAND2_X1 U19347 ( .A1(n16279), .A2(P2_STATE2_REG_0__SCAN_IN), .ZN(n16285) );
  NAND2_X1 U19348 ( .A1(n16281), .A2(n16280), .ZN(n16282) );
  OR2_X1 U19349 ( .A1(n12660), .A2(n16282), .ZN(n16284) );
  AND2_X1 U19350 ( .A1(n19846), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n16283) );
  AND2_X1 U19351 ( .A1(n16284), .A2(n16283), .ZN(n16288) );
  NAND2_X1 U19352 ( .A1(n10983), .A2(n16286), .ZN(n16287) );
  AOI22_X1 U19353 ( .A1(n16288), .A2(n19843), .B1(n16287), .B2(n19841), .ZN(
        n16289) );
  AOI21_X1 U19354 ( .B1(n16294), .B2(P2_STATE2_REG_0__SCAN_IN), .A(n16289), 
        .ZN(n16290) );
  OAI211_X1 U19355 ( .C1(n16293), .C2(n16292), .A(n16291), .B(n16290), .ZN(
        P2_U3176) );
  INV_X1 U19356 ( .A(n16294), .ZN(n19713) );
  OAI221_X1 U19357 ( .B1(n19798), .B2(P2_STATE2_REG_0__SCAN_IN), .C1(n19798), 
        .C2(n19713), .A(n16295), .ZN(P2_U3593) );
  INV_X1 U19358 ( .A(n18531), .ZN(n16296) );
  NAND3_X1 U19359 ( .A1(n16313), .A2(n18586), .A3(n18741), .ZN(n17754) );
  INV_X1 U19360 ( .A(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n18707) );
  AOI22_X1 U19361 ( .A1(n17649), .A2(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        n18707), .B2(n17604), .ZN(n16305) );
  NOR2_X1 U19362 ( .A1(n17649), .A2(n16298), .ZN(n16303) );
  OAI21_X1 U19363 ( .B1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n16348), .A(
        n16299), .ZN(n16300) );
  OAI22_X1 U19364 ( .A1(n16303), .A2(n16300), .B1(
        P3_INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n18707), .ZN(n16304) );
  NAND2_X1 U19365 ( .A1(n16301), .A2(n16305), .ZN(n16302) );
  OAI22_X1 U19366 ( .A1(n16305), .A2(n16304), .B1(n16303), .B2(n16302), .ZN(
        n16357) );
  NOR2_X1 U19367 ( .A1(n18074), .A2(n18684), .ZN(n16351) );
  INV_X1 U19368 ( .A(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n17398) );
  NOR2_X1 U19369 ( .A1(n17442), .A2(n17410), .ZN(n17411) );
  NAND3_X1 U19370 ( .A1(n17411), .A2(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n17397) );
  NOR2_X1 U19371 ( .A1(n17398), .A2(n17397), .ZN(n17368) );
  NAND3_X1 U19372 ( .A1(n17368), .A2(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A3(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n16334) );
  NOR2_X1 U19373 ( .A1(n16479), .A2(n16334), .ZN(n16308) );
  NAND2_X1 U19374 ( .A1(n18604), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17533) );
  AOI21_X1 U19375 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n17452), .A(
        n18476), .ZN(n17582) );
  NAND2_X1 U19376 ( .A1(n16308), .A2(n17531), .ZN(n16321) );
  XNOR2_X1 U19377 ( .A(P3_PHYADDRPOINTER_REG_31__SCAN_IN), .B(
        P3_PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n16311) );
  NOR2_X1 U19378 ( .A1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .A2(n17483), .ZN(
        n16331) );
  INV_X1 U19379 ( .A(n16307), .ZN(n16309) );
  INV_X2 U19380 ( .A(n18476), .ZN(n18348) );
  OR2_X1 U19381 ( .A1(n18348), .A2(n16308), .ZN(n16335) );
  OAI211_X1 U19382 ( .C1(n16309), .C2(n17533), .A(n17750), .B(n16335), .ZN(
        n16338) );
  NOR2_X1 U19383 ( .A1(n16331), .A2(n16338), .ZN(n16320) );
  OAI22_X1 U19384 ( .A1(n16321), .A2(n16311), .B1(n16320), .B2(n16310), .ZN(
        n16312) );
  AOI211_X1 U19385 ( .C1(n17575), .C2(n16797), .A(n16351), .B(n16312), .ZN(
        n16318) );
  NAND2_X1 U19386 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16339), .ZN(
        n16314) );
  XOR2_X1 U19387 ( .A(n16314), .B(n18707), .Z(n16354) );
  NAND2_X1 U19388 ( .A1(n16328), .A2(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(
        n16316) );
  XOR2_X1 U19389 ( .A(n16316), .B(n18707), .Z(n16353) );
  AOI22_X1 U19390 ( .A1(n17742), .A2(n16354), .B1(n17579), .B2(n16353), .ZN(
        n16317) );
  OAI221_X1 U19391 ( .B1(P3_PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n16321), .C1(
        n16469), .C2(n16320), .A(n16319), .ZN(n16322) );
  AOI21_X1 U19392 ( .B1(n17575), .B2(n16468), .A(n16322), .ZN(n16326) );
  OAI22_X1 U19393 ( .A1(n16339), .A2(n17755), .B1(n16328), .B2(n17652), .ZN(
        n16324) );
  AOI22_X1 U19394 ( .A1(n17606), .A2(n17742), .B1(n17579), .B2(n17647), .ZN(
        n17643) );
  NOR2_X2 U19395 ( .A1(n17870), .A2(n17643), .ZN(n17540) );
  INV_X1 U19396 ( .A(n17540), .ZN(n17459) );
  NOR2_X1 U19397 ( .A1(n17756), .A2(n17459), .ZN(n17392) );
  AOI22_X1 U19398 ( .A1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .A2(n16324), .B1(
        n16323), .B2(n17392), .ZN(n16325) );
  OAI211_X1 U19399 ( .C1(n17555), .C2(n16327), .A(n16326), .B(n16325), .ZN(
        P3_U2800) );
  AOI211_X1 U19400 ( .C1(n16330), .C2(n16329), .A(n16328), .B(n17652), .ZN(
        n16337) );
  NAND2_X1 U19401 ( .A1(n9820), .A2(P3_REIP_REG_29__SCAN_IN), .ZN(n16333) );
  OAI21_X1 U19402 ( .B1(n16331), .B2(n17575), .A(n16478), .ZN(n16332) );
  OAI211_X1 U19403 ( .C1(n16335), .C2(n16334), .A(n16333), .B(n16332), .ZN(
        n16336) );
  AOI211_X1 U19404 ( .C1(P3_PHYADDRPOINTER_REG_29__SCAN_IN), .C2(n16338), .A(
        n16337), .B(n16336), .ZN(n16343) );
  NOR2_X1 U19405 ( .A1(n16339), .A2(n17755), .ZN(n16340) );
  OAI21_X1 U19406 ( .B1(n16341), .B2(P3_INSTADDRPOINTER_REG_29__SCAN_IN), .A(
        n16340), .ZN(n16342) );
  OAI211_X1 U19407 ( .C1(n16344), .C2(n17555), .A(n16343), .B(n16342), .ZN(
        P3_U2801) );
  INV_X1 U19408 ( .A(n16345), .ZN(n17887) );
  NOR2_X1 U19409 ( .A1(n18061), .A2(n17887), .ZN(n18068) );
  INV_X1 U19410 ( .A(n18068), .ZN(n18011) );
  OAI211_X1 U19411 ( .C1(P3_INSTADDRPOINTER_REG_30__SCAN_IN), .C2(n18011), .A(
        n18062), .B(n16346), .ZN(n16352) );
  NOR4_X1 U19412 ( .A1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .A2(n16349), .A3(
        n16348), .A4(n16347), .ZN(n16350) );
  AOI211_X1 U19413 ( .C1(P3_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(n16352), .A(
        n16351), .B(n16350), .ZN(n16356) );
  AOI22_X1 U19414 ( .A1(n16354), .A2(n18037), .B1(n16353), .B2(n17995), .ZN(
        n16355) );
  NOR3_X1 U19415 ( .A1(P3_W_R_N_REG_SCAN_IN), .A2(P3_BE_N_REG_0__SCAN_IN), 
        .A3(P3_BE_N_REG_1__SCAN_IN), .ZN(n16359) );
  NOR4_X1 U19416 ( .A1(P3_BE_N_REG_2__SCAN_IN), .A2(P3_BE_N_REG_3__SCAN_IN), 
        .A3(P3_D_C_N_REG_SCAN_IN), .A4(P3_ADS_N_REG_SCAN_IN), .ZN(n16358) );
  NAND4_X1 U19417 ( .A1(P3_M_IO_N_REG_SCAN_IN), .A2(n16359), .A3(n16358), .A4(
        U215), .ZN(U213) );
  INV_X1 U19418 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n19017) );
  INV_X2 U19419 ( .A(U214), .ZN(n16405) );
  NOR2_X1 U19420 ( .A1(n16405), .A2(n16360), .ZN(n16393) );
  INV_X2 U19421 ( .A(n16393), .ZN(n16407) );
  INV_X1 U19422 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n16440) );
  OAI222_X1 U19423 ( .A1(U212), .A2(n19017), .B1(n16407), .B2(n19147), .C1(
        U214), .C2(n16440), .ZN(U216) );
  AOI22_X1 U19424 ( .A1(P1_DATAO_REG_30__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n16404), .ZN(n16361) );
  OAI21_X1 U19425 ( .B1(n14508), .B2(n16407), .A(n16361), .ZN(U217) );
  AOI22_X1 U19426 ( .A1(P1_DATAO_REG_29__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_29__SCAN_IN), .B2(n16404), .ZN(n16362) );
  OAI21_X1 U19427 ( .B1(n14307), .B2(n16407), .A(n16362), .ZN(U218) );
  AOI22_X1 U19428 ( .A1(P1_DATAO_REG_28__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_28__SCAN_IN), .B2(n16404), .ZN(n16363) );
  OAI21_X1 U19429 ( .B1(n16364), .B2(n16407), .A(n16363), .ZN(U219) );
  INV_X1 U19430 ( .A(BUF1_REG_27__SCAN_IN), .ZN(n16366) );
  AOI22_X1 U19431 ( .A1(P1_DATAO_REG_27__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_27__SCAN_IN), .B2(n16404), .ZN(n16365) );
  OAI21_X1 U19432 ( .B1(n16366), .B2(n16407), .A(n16365), .ZN(U220) );
  INV_X1 U19433 ( .A(BUF1_REG_26__SCAN_IN), .ZN(n16368) );
  AOI22_X1 U19434 ( .A1(P1_DATAO_REG_26__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_26__SCAN_IN), .B2(n16404), .ZN(n16367) );
  OAI21_X1 U19435 ( .B1(n16368), .B2(n16407), .A(n16367), .ZN(U221) );
  INV_X1 U19436 ( .A(BUF1_REG_25__SCAN_IN), .ZN(n20121) );
  AOI22_X1 U19437 ( .A1(P1_DATAO_REG_25__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_25__SCAN_IN), .B2(n16404), .ZN(n16369) );
  OAI21_X1 U19438 ( .B1(n20121), .B2(n16407), .A(n16369), .ZN(U222) );
  INV_X1 U19439 ( .A(BUF1_REG_24__SCAN_IN), .ZN(n16371) );
  AOI22_X1 U19440 ( .A1(P1_DATAO_REG_24__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_24__SCAN_IN), .B2(n16404), .ZN(n16370) );
  OAI21_X1 U19441 ( .B1(n16371), .B2(n16407), .A(n16370), .ZN(U223) );
  AOI22_X1 U19442 ( .A1(P1_DATAO_REG_23__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_23__SCAN_IN), .B2(n16404), .ZN(n16372) );
  OAI21_X1 U19443 ( .B1(n15068), .B2(n16407), .A(n16372), .ZN(U224) );
  AOI22_X1 U19444 ( .A1(P1_DATAO_REG_22__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_22__SCAN_IN), .B2(n16404), .ZN(n16373) );
  OAI21_X1 U19445 ( .B1(n14540), .B2(n16407), .A(n16373), .ZN(U225) );
  INV_X1 U19446 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n16428) );
  INV_X1 U19447 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n20876) );
  OAI222_X1 U19448 ( .A1(U212), .A2(n16428), .B1(n16407), .B2(n15074), .C1(
        U214), .C2(n20876), .ZN(U226) );
  AOI22_X1 U19449 ( .A1(P1_DATAO_REG_20__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_20__SCAN_IN), .B2(n16404), .ZN(n16374) );
  OAI21_X1 U19450 ( .B1(n16375), .B2(n16407), .A(n16374), .ZN(U227) );
  AOI22_X1 U19451 ( .A1(P1_DATAO_REG_19__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_19__SCAN_IN), .B2(n16404), .ZN(n16376) );
  OAI21_X1 U19452 ( .B1(n15085), .B2(n16407), .A(n16376), .ZN(U228) );
  AOI22_X1 U19453 ( .A1(P1_DATAO_REG_18__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_18__SCAN_IN), .B2(n16404), .ZN(n16377) );
  OAI21_X1 U19454 ( .B1(n14561), .B2(n16407), .A(n16377), .ZN(U229) );
  AOI22_X1 U19455 ( .A1(P1_DATAO_REG_17__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_17__SCAN_IN), .B2(n16404), .ZN(n16378) );
  OAI21_X1 U19456 ( .B1(n14208), .B2(n16407), .A(n16378), .ZN(U230) );
  AOI22_X1 U19457 ( .A1(P1_DATAO_REG_16__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n16404), .ZN(n16379) );
  OAI21_X1 U19458 ( .B1(n14176), .B2(n16407), .A(n16379), .ZN(U231) );
  AOI22_X1 U19459 ( .A1(P1_DATAO_REG_15__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_15__SCAN_IN), .B2(n16404), .ZN(n16380) );
  OAI21_X1 U19460 ( .B1(n13285), .B2(n16407), .A(n16380), .ZN(U232) );
  AOI222_X1 U19461 ( .A1(n16404), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n16393), 
        .B2(BUF1_REG_14__SCAN_IN), .C1(n16405), .C2(P1_DATAO_REG_14__SCAN_IN), 
        .ZN(n16381) );
  INV_X1 U19462 ( .A(n16381), .ZN(U233) );
  INV_X1 U19463 ( .A(BUF1_REG_13__SCAN_IN), .ZN(n16383) );
  AOI22_X1 U19464 ( .A1(P1_DATAO_REG_13__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n16404), .ZN(n16382) );
  OAI21_X1 U19465 ( .B1(n16383), .B2(n16407), .A(n16382), .ZN(U234) );
  AOI22_X1 U19466 ( .A1(P1_DATAO_REG_12__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n16404), .ZN(n16384) );
  OAI21_X1 U19467 ( .B1(n14136), .B2(n16407), .A(n16384), .ZN(U235) );
  AOI22_X1 U19468 ( .A1(P1_DATAO_REG_11__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_11__SCAN_IN), .B2(n16404), .ZN(n16385) );
  OAI21_X1 U19469 ( .B1(n14125), .B2(n16407), .A(n16385), .ZN(U236) );
  AOI222_X1 U19470 ( .A1(n16404), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n16393), 
        .B2(BUF1_REG_10__SCAN_IN), .C1(n16405), .C2(P1_DATAO_REG_10__SCAN_IN), 
        .ZN(n16386) );
  INV_X1 U19471 ( .A(n16386), .ZN(U237) );
  AOI22_X1 U19472 ( .A1(P1_DATAO_REG_9__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_9__SCAN_IN), .B2(n16404), .ZN(n16387) );
  OAI21_X1 U19473 ( .B1(n16388), .B2(n16407), .A(n16387), .ZN(U238) );
  AOI22_X1 U19474 ( .A1(P1_DATAO_REG_8__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n16404), .ZN(n16389) );
  OAI21_X1 U19475 ( .B1(n16390), .B2(n16407), .A(n16389), .ZN(U239) );
  INV_X1 U19476 ( .A(BUF1_REG_7__SCAN_IN), .ZN(n16392) );
  AOI22_X1 U19477 ( .A1(P1_DATAO_REG_7__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_7__SCAN_IN), .B2(n16404), .ZN(n16391) );
  OAI21_X1 U19478 ( .B1(n16392), .B2(n16407), .A(n16391), .ZN(U240) );
  AOI222_X1 U19479 ( .A1(n16404), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n16393), 
        .B2(BUF1_REG_6__SCAN_IN), .C1(n16405), .C2(P1_DATAO_REG_6__SCAN_IN), 
        .ZN(n16394) );
  INV_X1 U19480 ( .A(n16394), .ZN(U241) );
  INV_X1 U19481 ( .A(BUF1_REG_5__SCAN_IN), .ZN(n16396) );
  AOI22_X1 U19482 ( .A1(P1_DATAO_REG_5__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_5__SCAN_IN), .B2(n16404), .ZN(n16395) );
  OAI21_X1 U19483 ( .B1(n16396), .B2(n16407), .A(n16395), .ZN(U242) );
  INV_X1 U19484 ( .A(BUF1_REG_4__SCAN_IN), .ZN(n16398) );
  AOI22_X1 U19485 ( .A1(P1_DATAO_REG_4__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_4__SCAN_IN), .B2(n16404), .ZN(n16397) );
  OAI21_X1 U19486 ( .B1(n16398), .B2(n16407), .A(n16397), .ZN(U243) );
  INV_X1 U19487 ( .A(BUF1_REG_3__SCAN_IN), .ZN(n16400) );
  AOI22_X1 U19488 ( .A1(P1_DATAO_REG_3__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_3__SCAN_IN), .B2(n16404), .ZN(n16399) );
  OAI21_X1 U19489 ( .B1(n16400), .B2(n16407), .A(n16399), .ZN(U244) );
  INV_X1 U19490 ( .A(BUF1_REG_2__SCAN_IN), .ZN(n16402) );
  AOI22_X1 U19491 ( .A1(P1_DATAO_REG_2__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_2__SCAN_IN), .B2(n16404), .ZN(n16401) );
  OAI21_X1 U19492 ( .B1(n16402), .B2(n16407), .A(n16401), .ZN(U245) );
  INV_X1 U19493 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n20937) );
  INV_X1 U19494 ( .A(BUF1_REG_1__SCAN_IN), .ZN(n20916) );
  INV_X1 U19495 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n16403) );
  OAI222_X1 U19496 ( .A1(U212), .A2(n20937), .B1(n16407), .B2(n20916), .C1(
        U214), .C2(n16403), .ZN(U246) );
  INV_X1 U19497 ( .A(BUF1_REG_0__SCAN_IN), .ZN(n16408) );
  AOI22_X1 U19498 ( .A1(P1_DATAO_REG_0__SCAN_IN), .A2(n16405), .B1(
        P2_DATAO_REG_0__SCAN_IN), .B2(n16404), .ZN(n16406) );
  OAI21_X1 U19499 ( .B1(n16408), .B2(n16407), .A(n16406), .ZN(U247) );
  OAI22_X1 U19500 ( .A1(U215), .A2(P2_DATAO_REG_0__SCAN_IN), .B1(
        BUF2_REG_0__SCAN_IN), .B2(n16438), .ZN(n16409) );
  INV_X1 U19501 ( .A(n16409), .ZN(U251) );
  INV_X1 U19502 ( .A(BUF2_REG_1__SCAN_IN), .ZN(n18099) );
  AOI22_X1 U19503 ( .A1(n16438), .A2(n20937), .B1(n18099), .B2(U215), .ZN(U252) );
  OAI22_X1 U19504 ( .A1(U215), .A2(P2_DATAO_REG_2__SCAN_IN), .B1(
        BUF2_REG_2__SCAN_IN), .B2(n16422), .ZN(n16410) );
  INV_X1 U19505 ( .A(n16410), .ZN(U253) );
  OAI22_X1 U19506 ( .A1(U215), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(
        BUF2_REG_3__SCAN_IN), .B2(n16422), .ZN(n16411) );
  INV_X1 U19507 ( .A(n16411), .ZN(U254) );
  OAI22_X1 U19508 ( .A1(U215), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(
        BUF2_REG_4__SCAN_IN), .B2(n16422), .ZN(n16412) );
  INV_X1 U19509 ( .A(n16412), .ZN(U255) );
  OAI22_X1 U19510 ( .A1(U215), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(
        BUF2_REG_5__SCAN_IN), .B2(n16422), .ZN(n16413) );
  INV_X1 U19511 ( .A(n16413), .ZN(U256) );
  INV_X1 U19512 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n21037) );
  INV_X1 U19513 ( .A(BUF2_REG_6__SCAN_IN), .ZN(n18127) );
  AOI22_X1 U19514 ( .A1(n16438), .A2(n21037), .B1(n18127), .B2(U215), .ZN(U257) );
  OAI22_X1 U19515 ( .A1(U215), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(
        BUF2_REG_7__SCAN_IN), .B2(n16422), .ZN(n16414) );
  INV_X1 U19516 ( .A(n16414), .ZN(U258) );
  OAI22_X1 U19517 ( .A1(U215), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(
        BUF2_REG_8__SCAN_IN), .B2(n16422), .ZN(n16415) );
  INV_X1 U19518 ( .A(n16415), .ZN(U259) );
  OAI22_X1 U19519 ( .A1(U215), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(
        BUF2_REG_9__SCAN_IN), .B2(n16422), .ZN(n16416) );
  INV_X1 U19520 ( .A(n16416), .ZN(U260) );
  INV_X1 U19521 ( .A(P2_DATAO_REG_10__SCAN_IN), .ZN(n20945) );
  INV_X1 U19522 ( .A(BUF2_REG_10__SCAN_IN), .ZN(n17353) );
  AOI22_X1 U19523 ( .A1(n16438), .A2(n20945), .B1(n17353), .B2(U215), .ZN(U261) );
  OAI22_X1 U19524 ( .A1(U215), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(
        BUF2_REG_11__SCAN_IN), .B2(n16438), .ZN(n16417) );
  INV_X1 U19525 ( .A(n16417), .ZN(U262) );
  OAI22_X1 U19526 ( .A1(U215), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(
        BUF2_REG_12__SCAN_IN), .B2(n16422), .ZN(n16418) );
  INV_X1 U19527 ( .A(n16418), .ZN(U263) );
  OAI22_X1 U19528 ( .A1(U215), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(
        BUF2_REG_13__SCAN_IN), .B2(n16438), .ZN(n16419) );
  INV_X1 U19529 ( .A(n16419), .ZN(U264) );
  OAI22_X1 U19530 ( .A1(U215), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(
        BUF2_REG_14__SCAN_IN), .B2(n16422), .ZN(n16420) );
  INV_X1 U19531 ( .A(n16420), .ZN(U265) );
  OAI22_X1 U19532 ( .A1(U215), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(
        BUF2_REG_15__SCAN_IN), .B2(n16438), .ZN(n16421) );
  INV_X1 U19533 ( .A(n16421), .ZN(U266) );
  OAI22_X1 U19534 ( .A1(U215), .A2(P2_DATAO_REG_16__SCAN_IN), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n16422), .ZN(n16423) );
  INV_X1 U19535 ( .A(n16423), .ZN(U267) );
  OAI22_X1 U19536 ( .A1(U215), .A2(P2_DATAO_REG_17__SCAN_IN), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n16438), .ZN(n16424) );
  INV_X1 U19537 ( .A(n16424), .ZN(U268) );
  OAI22_X1 U19538 ( .A1(U215), .A2(P2_DATAO_REG_18__SCAN_IN), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n16438), .ZN(n16425) );
  INV_X1 U19539 ( .A(n16425), .ZN(U269) );
  OAI22_X1 U19540 ( .A1(U215), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n16438), .ZN(n16426) );
  INV_X1 U19541 ( .A(n16426), .ZN(U270) );
  OAI22_X1 U19542 ( .A1(U215), .A2(P2_DATAO_REG_20__SCAN_IN), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n16438), .ZN(n16427) );
  INV_X1 U19543 ( .A(n16427), .ZN(U271) );
  AOI22_X1 U19544 ( .A1(n16438), .A2(n16428), .B1(n15075), .B2(U215), .ZN(U272) );
  OAI22_X1 U19545 ( .A1(U215), .A2(P2_DATAO_REG_22__SCAN_IN), .B1(
        BUF2_REG_22__SCAN_IN), .B2(n16438), .ZN(n16429) );
  INV_X1 U19546 ( .A(n16429), .ZN(U273) );
  OAI22_X1 U19547 ( .A1(U215), .A2(P2_DATAO_REG_23__SCAN_IN), .B1(
        BUF2_REG_23__SCAN_IN), .B2(n16438), .ZN(n16430) );
  INV_X1 U19548 ( .A(n16430), .ZN(U274) );
  OAI22_X1 U19549 ( .A1(U215), .A2(P2_DATAO_REG_24__SCAN_IN), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n16438), .ZN(n16431) );
  INV_X1 U19550 ( .A(n16431), .ZN(U275) );
  OAI22_X1 U19551 ( .A1(U215), .A2(P2_DATAO_REG_25__SCAN_IN), .B1(
        BUF2_REG_25__SCAN_IN), .B2(n16438), .ZN(n16432) );
  INV_X1 U19552 ( .A(n16432), .ZN(U276) );
  OAI22_X1 U19553 ( .A1(U215), .A2(P2_DATAO_REG_26__SCAN_IN), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n16438), .ZN(n16433) );
  INV_X1 U19554 ( .A(n16433), .ZN(U277) );
  OAI22_X1 U19555 ( .A1(U215), .A2(P2_DATAO_REG_27__SCAN_IN), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n16438), .ZN(n16434) );
  INV_X1 U19556 ( .A(n16434), .ZN(U278) );
  OAI22_X1 U19557 ( .A1(U215), .A2(P2_DATAO_REG_28__SCAN_IN), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n16438), .ZN(n16435) );
  INV_X1 U19558 ( .A(n16435), .ZN(U279) );
  OAI22_X1 U19559 ( .A1(U215), .A2(P2_DATAO_REG_29__SCAN_IN), .B1(
        BUF2_REG_29__SCAN_IN), .B2(n16438), .ZN(n16436) );
  INV_X1 U19560 ( .A(n16436), .ZN(U280) );
  OAI22_X1 U19561 ( .A1(U215), .A2(P2_DATAO_REG_30__SCAN_IN), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n16438), .ZN(n16437) );
  INV_X1 U19562 ( .A(n16437), .ZN(U281) );
  INV_X1 U19563 ( .A(BUF2_REG_31__SCAN_IN), .ZN(n19145) );
  AOI22_X1 U19564 ( .A1(n16438), .A2(n19017), .B1(n19145), .B2(U215), .ZN(U282) );
  INV_X1 U19565 ( .A(P3_DATAO_REG_31__SCAN_IN), .ZN(n16439) );
  AOI222_X1 U19566 ( .A1(n16440), .A2(P1_DATAO_REG_30__SCAN_IN), .B1(n19017), 
        .B2(P2_DATAO_REG_30__SCAN_IN), .C1(n16439), .C2(
        P3_DATAO_REG_30__SCAN_IN), .ZN(n16441) );
  INV_X2 U19567 ( .A(n16443), .ZN(n16442) );
  INV_X1 U19568 ( .A(P3_ADDRESS_REG_9__SCAN_IN), .ZN(n18642) );
  INV_X1 U19569 ( .A(P2_ADDRESS_REG_9__SCAN_IN), .ZN(n19743) );
  AOI22_X1 U19570 ( .A1(n16442), .A2(n18642), .B1(n19743), .B2(n16443), .ZN(
        U347) );
  INV_X1 U19571 ( .A(P3_ADDRESS_REG_8__SCAN_IN), .ZN(n21104) );
  INV_X1 U19572 ( .A(P2_ADDRESS_REG_8__SCAN_IN), .ZN(n19742) );
  AOI22_X1 U19573 ( .A1(n16442), .A2(n21104), .B1(n19742), .B2(n16443), .ZN(
        U348) );
  INV_X1 U19574 ( .A(P3_ADDRESS_REG_7__SCAN_IN), .ZN(n18639) );
  INV_X1 U19575 ( .A(P2_ADDRESS_REG_7__SCAN_IN), .ZN(n19741) );
  AOI22_X1 U19576 ( .A1(n16442), .A2(n18639), .B1(n19741), .B2(n16443), .ZN(
        U349) );
  INV_X1 U19577 ( .A(P3_ADDRESS_REG_6__SCAN_IN), .ZN(n18637) );
  INV_X1 U19578 ( .A(P2_ADDRESS_REG_6__SCAN_IN), .ZN(n19740) );
  AOI22_X1 U19579 ( .A1(n16442), .A2(n18637), .B1(n19740), .B2(n16443), .ZN(
        U350) );
  INV_X1 U19580 ( .A(P3_ADDRESS_REG_5__SCAN_IN), .ZN(n18635) );
  INV_X1 U19581 ( .A(P2_ADDRESS_REG_5__SCAN_IN), .ZN(n20893) );
  AOI22_X1 U19582 ( .A1(n16442), .A2(n18635), .B1(n20893), .B2(n16443), .ZN(
        U351) );
  INV_X1 U19583 ( .A(P3_ADDRESS_REG_4__SCAN_IN), .ZN(n18633) );
  INV_X1 U19584 ( .A(P2_ADDRESS_REG_4__SCAN_IN), .ZN(n19739) );
  AOI22_X1 U19585 ( .A1(n16442), .A2(n18633), .B1(n19739), .B2(n16443), .ZN(
        U352) );
  INV_X1 U19586 ( .A(P3_ADDRESS_REG_3__SCAN_IN), .ZN(n18632) );
  INV_X1 U19587 ( .A(P2_ADDRESS_REG_3__SCAN_IN), .ZN(n21095) );
  AOI22_X1 U19588 ( .A1(n16442), .A2(n18632), .B1(n21095), .B2(n16443), .ZN(
        U353) );
  INV_X1 U19589 ( .A(P3_ADDRESS_REG_2__SCAN_IN), .ZN(n18630) );
  AOI22_X1 U19590 ( .A1(n16442), .A2(n18630), .B1(n19738), .B2(n16443), .ZN(
        U354) );
  INV_X1 U19591 ( .A(P3_ADDRESS_REG_29__SCAN_IN), .ZN(n18683) );
  INV_X1 U19592 ( .A(P2_ADDRESS_REG_29__SCAN_IN), .ZN(n19773) );
  AOI22_X1 U19593 ( .A1(n16442), .A2(n18683), .B1(n19773), .B2(n16443), .ZN(
        U355) );
  INV_X1 U19594 ( .A(P3_ADDRESS_REG_28__SCAN_IN), .ZN(n18679) );
  INV_X1 U19595 ( .A(P2_ADDRESS_REG_28__SCAN_IN), .ZN(n19771) );
  AOI22_X1 U19596 ( .A1(n16442), .A2(n18679), .B1(n19771), .B2(n16443), .ZN(
        U356) );
  INV_X1 U19597 ( .A(P3_ADDRESS_REG_26__SCAN_IN), .ZN(n18674) );
  INV_X1 U19598 ( .A(P2_ADDRESS_REG_26__SCAN_IN), .ZN(n19766) );
  AOI22_X1 U19599 ( .A1(n16442), .A2(n18674), .B1(n19766), .B2(n16443), .ZN(
        U358) );
  INV_X1 U19600 ( .A(P3_ADDRESS_REG_25__SCAN_IN), .ZN(n18673) );
  INV_X1 U19601 ( .A(P2_ADDRESS_REG_25__SCAN_IN), .ZN(n19765) );
  AOI22_X1 U19602 ( .A1(n16442), .A2(n18673), .B1(n19765), .B2(n16443), .ZN(
        U359) );
  INV_X1 U19603 ( .A(P3_ADDRESS_REG_24__SCAN_IN), .ZN(n18671) );
  INV_X1 U19604 ( .A(P2_ADDRESS_REG_24__SCAN_IN), .ZN(n19764) );
  AOI22_X1 U19605 ( .A1(n16442), .A2(n18671), .B1(n19764), .B2(n16443), .ZN(
        U360) );
  INV_X1 U19606 ( .A(P3_ADDRESS_REG_23__SCAN_IN), .ZN(n18668) );
  INV_X1 U19607 ( .A(P2_ADDRESS_REG_23__SCAN_IN), .ZN(n19762) );
  AOI22_X1 U19608 ( .A1(n16442), .A2(n18668), .B1(n19762), .B2(n16443), .ZN(
        U361) );
  INV_X1 U19609 ( .A(P3_ADDRESS_REG_22__SCAN_IN), .ZN(n18667) );
  INV_X1 U19610 ( .A(P2_ADDRESS_REG_22__SCAN_IN), .ZN(n19761) );
  AOI22_X1 U19611 ( .A1(n16442), .A2(n18667), .B1(n19761), .B2(n16443), .ZN(
        U362) );
  INV_X1 U19612 ( .A(P3_ADDRESS_REG_21__SCAN_IN), .ZN(n18666) );
  INV_X1 U19613 ( .A(P2_ADDRESS_REG_21__SCAN_IN), .ZN(n19760) );
  AOI22_X1 U19614 ( .A1(n16442), .A2(n18666), .B1(n19760), .B2(n16443), .ZN(
        U363) );
  INV_X1 U19615 ( .A(P3_ADDRESS_REG_20__SCAN_IN), .ZN(n18664) );
  INV_X1 U19616 ( .A(P2_ADDRESS_REG_20__SCAN_IN), .ZN(n19759) );
  AOI22_X1 U19617 ( .A1(n16442), .A2(n18664), .B1(n19759), .B2(n16443), .ZN(
        U364) );
  INV_X1 U19618 ( .A(P3_ADDRESS_REG_1__SCAN_IN), .ZN(n18628) );
  INV_X1 U19619 ( .A(P2_ADDRESS_REG_1__SCAN_IN), .ZN(n19737) );
  AOI22_X1 U19620 ( .A1(n16442), .A2(n18628), .B1(n19737), .B2(n16443), .ZN(
        U365) );
  INV_X1 U19621 ( .A(P3_ADDRESS_REG_19__SCAN_IN), .ZN(n18662) );
  INV_X1 U19622 ( .A(P2_ADDRESS_REG_19__SCAN_IN), .ZN(n19757) );
  AOI22_X1 U19623 ( .A1(n16442), .A2(n18662), .B1(n19757), .B2(n16443), .ZN(
        U366) );
  INV_X1 U19624 ( .A(P3_ADDRESS_REG_18__SCAN_IN), .ZN(n18660) );
  INV_X1 U19625 ( .A(P2_ADDRESS_REG_18__SCAN_IN), .ZN(n19755) );
  AOI22_X1 U19626 ( .A1(n16442), .A2(n18660), .B1(n19755), .B2(n16443), .ZN(
        U367) );
  INV_X1 U19627 ( .A(P3_ADDRESS_REG_17__SCAN_IN), .ZN(n18658) );
  INV_X1 U19628 ( .A(P2_ADDRESS_REG_17__SCAN_IN), .ZN(n19753) );
  AOI22_X1 U19629 ( .A1(n16442), .A2(n18658), .B1(n19753), .B2(n16443), .ZN(
        U368) );
  INV_X1 U19630 ( .A(P3_ADDRESS_REG_16__SCAN_IN), .ZN(n18656) );
  INV_X1 U19631 ( .A(P2_ADDRESS_REG_16__SCAN_IN), .ZN(n19751) );
  AOI22_X1 U19632 ( .A1(n16442), .A2(n18656), .B1(n19751), .B2(n16443), .ZN(
        U369) );
  INV_X1 U19633 ( .A(P3_ADDRESS_REG_15__SCAN_IN), .ZN(n18654) );
  INV_X1 U19634 ( .A(P2_ADDRESS_REG_15__SCAN_IN), .ZN(n19749) );
  AOI22_X1 U19635 ( .A1(n16442), .A2(n18654), .B1(n19749), .B2(n16443), .ZN(
        U370) );
  INV_X1 U19636 ( .A(P3_ADDRESS_REG_14__SCAN_IN), .ZN(n18652) );
  INV_X1 U19637 ( .A(P2_ADDRESS_REG_14__SCAN_IN), .ZN(n19748) );
  AOI22_X1 U19638 ( .A1(n16442), .A2(n18652), .B1(n19748), .B2(n16443), .ZN(
        U371) );
  INV_X1 U19639 ( .A(P3_ADDRESS_REG_13__SCAN_IN), .ZN(n18650) );
  INV_X1 U19640 ( .A(P2_ADDRESS_REG_13__SCAN_IN), .ZN(n19746) );
  AOI22_X1 U19641 ( .A1(n16442), .A2(n18650), .B1(n19746), .B2(n16443), .ZN(
        U372) );
  INV_X1 U19642 ( .A(P3_ADDRESS_REG_12__SCAN_IN), .ZN(n18648) );
  INV_X1 U19643 ( .A(P2_ADDRESS_REG_12__SCAN_IN), .ZN(n19745) );
  AOI22_X1 U19644 ( .A1(n16442), .A2(n18648), .B1(n19745), .B2(n16443), .ZN(
        U373) );
  INV_X1 U19645 ( .A(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n18646) );
  INV_X1 U19646 ( .A(P2_ADDRESS_REG_11__SCAN_IN), .ZN(n19744) );
  AOI22_X1 U19647 ( .A1(n16442), .A2(n18646), .B1(n19744), .B2(n16443), .ZN(
        U374) );
  INV_X1 U19648 ( .A(P3_ADDRESS_REG_10__SCAN_IN), .ZN(n18644) );
  INV_X1 U19649 ( .A(P2_ADDRESS_REG_10__SCAN_IN), .ZN(n21030) );
  AOI22_X1 U19650 ( .A1(n16442), .A2(n18644), .B1(n21030), .B2(n16443), .ZN(
        U375) );
  INV_X1 U19651 ( .A(P3_ADDRESS_REG_0__SCAN_IN), .ZN(n18626) );
  INV_X1 U19652 ( .A(P2_ADDRESS_REG_0__SCAN_IN), .ZN(n19736) );
  AOI22_X1 U19653 ( .A1(n16442), .A2(n18626), .B1(n19736), .B2(n16443), .ZN(
        U376) );
  INV_X1 U19654 ( .A(P3_STATE_REG_2__SCAN_IN), .ZN(n18625) );
  NAND2_X1 U19655 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(n18625), .ZN(n18612) );
  AOI22_X1 U19656 ( .A1(P3_STATE_REG_0__SCAN_IN), .A2(n18612), .B1(
        P3_STATE_REG_1__SCAN_IN), .B2(n18623), .ZN(n18693) );
  AOI21_X1 U19657 ( .B1(P3_STATE_REG_0__SCAN_IN), .B2(P3_ADS_N_REG_SCAN_IN), 
        .A(n18693), .ZN(n16444) );
  INV_X1 U19658 ( .A(n16444), .ZN(P3_U2633) );
  INV_X1 U19659 ( .A(n17751), .ZN(n18598) );
  OAI21_X1 U19660 ( .B1(n16449), .B2(n17313), .A(P3_CODEFETCH_REG_SCAN_IN), 
        .ZN(n16445) );
  OAI21_X1 U19661 ( .B1(n16446), .B2(n18598), .A(n16445), .ZN(P3_U2634) );
  AOI21_X1 U19662 ( .B1(n18623), .B2(n18625), .A(P3_D_C_N_REG_SCAN_IN), .ZN(
        n16447) );
  AOI22_X1 U19663 ( .A1(n18682), .A2(P3_CODEFETCH_REG_SCAN_IN), .B1(n16447), 
        .B2(n18755), .ZN(P3_U2635) );
  OAI21_X1 U19664 ( .B1(n18609), .B2(BS16), .A(n18693), .ZN(n18691) );
  OAI21_X1 U19665 ( .B1(n18693), .B2(n18745), .A(n18691), .ZN(P3_U2636) );
  NOR3_X1 U19666 ( .A1(n16449), .A2(n16448), .A3(n18530), .ZN(n18536) );
  NOR2_X1 U19667 ( .A1(n18536), .A2(n18595), .ZN(n18738) );
  OAI21_X1 U19668 ( .B1(n18738), .B2(n18082), .A(n16450), .ZN(P3_U2637) );
  NOR4_X1 U19669 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_20__SCAN_IN), .A3(P3_DATAWIDTH_REG_21__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_22__SCAN_IN), .ZN(n16454) );
  NOR4_X1 U19670 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_16__SCAN_IN), .A3(P3_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_18__SCAN_IN), .ZN(n16453) );
  NOR4_X1 U19671 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_29__SCAN_IN), .A3(P3_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_31__SCAN_IN), .ZN(n16452) );
  NOR4_X1 U19672 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_24__SCAN_IN), .A3(P3_DATAWIDTH_REG_25__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_27__SCAN_IN), .ZN(n16451) );
  NAND4_X1 U19673 ( .A1(n16454), .A2(n16453), .A3(n16452), .A4(n16451), .ZN(
        n16460) );
  NOR4_X1 U19674 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_4__SCAN_IN), .A3(P3_DATAWIDTH_REG_5__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_6__SCAN_IN), .ZN(n16458) );
  AOI211_X1 U19675 ( .C1(P3_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_3__SCAN_IN), .B(
        P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n16457) );
  NOR4_X1 U19676 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_12__SCAN_IN), .A3(P3_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_14__SCAN_IN), .ZN(n16456) );
  NOR4_X1 U19677 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_8__SCAN_IN), .A3(P3_DATAWIDTH_REG_9__SCAN_IN), .A4(
        P3_DATAWIDTH_REG_10__SCAN_IN), .ZN(n16455) );
  NAND4_X1 U19678 ( .A1(n16458), .A2(n16457), .A3(n16456), .A4(n16455), .ZN(
        n16459) );
  NOR2_X1 U19679 ( .A1(n16460), .A2(n16459), .ZN(n18736) );
  INV_X1 U19680 ( .A(P3_BYTEENABLE_REG_1__SCAN_IN), .ZN(n16462) );
  NOR3_X1 U19681 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(
        P3_DATAWIDTH_REG_1__SCAN_IN), .A3(P3_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n16463) );
  OAI21_X1 U19682 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(n16463), .A(n18736), .ZN(
        n16461) );
  OAI21_X1 U19683 ( .B1(n18736), .B2(n16462), .A(n16461), .ZN(P3_U2638) );
  INV_X1 U19684 ( .A(P3_REIP_REG_1__SCAN_IN), .ZN(n18729) );
  INV_X1 U19685 ( .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(n18692) );
  AOI21_X1 U19686 ( .B1(n18729), .B2(n18692), .A(n16463), .ZN(n16465) );
  INV_X1 U19687 ( .A(P3_BYTEENABLE_REG_3__SCAN_IN), .ZN(n16464) );
  INV_X1 U19688 ( .A(n18736), .ZN(n18731) );
  AOI22_X1 U19689 ( .A1(n18736), .A2(n16465), .B1(n16464), .B2(n18731), .ZN(
        P3_U2639) );
  NAND2_X1 U19690 ( .A1(n16811), .A2(n16466), .ZN(n16485) );
  XOR2_X1 U19691 ( .A(n16468), .B(n16467), .Z(n16472) );
  OAI22_X1 U19692 ( .A1(n16480), .A2(n18681), .B1(n16469), .B2(n16798), .ZN(
        n16470) );
  OAI21_X1 U19693 ( .B1(n16812), .B2(n16473), .A(P3_EBX_REG_30__SCAN_IN), .ZN(
        n16474) );
  OAI211_X1 U19694 ( .C1(P3_EBX_REG_30__SCAN_IN), .C2(n16485), .A(n16475), .B(
        n16474), .ZN(P3_U2641) );
  NOR2_X1 U19695 ( .A1(n16489), .A2(n16856), .ZN(n16486) );
  AOI211_X1 U19696 ( .C1(n16478), .C2(n16477), .A(n16476), .B(n18602), .ZN(
        n16482) );
  INV_X1 U19697 ( .A(P3_REIP_REG_29__SCAN_IN), .ZN(n18678) );
  OAI22_X1 U19698 ( .A1(n16480), .A2(n18678), .B1(n16479), .B2(n16798), .ZN(
        n16481) );
  AOI211_X1 U19699 ( .C1(P3_EBX_REG_29__SCAN_IN), .C2(n16812), .A(n16482), .B(
        n16481), .ZN(n16484) );
  NAND3_X1 U19700 ( .A1(P3_REIP_REG_28__SCAN_IN), .A2(n16487), .A3(n18678), 
        .ZN(n16483) );
  OAI211_X1 U19701 ( .C1(n16486), .C2(n16485), .A(n16484), .B(n16483), .ZN(
        P3_U2642) );
  INV_X1 U19702 ( .A(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n17369) );
  INV_X1 U19703 ( .A(P3_REIP_REG_28__SCAN_IN), .ZN(n18676) );
  AOI22_X1 U19704 ( .A1(P3_EBX_REG_28__SCAN_IN), .A2(n16812), .B1(n16487), 
        .B2(n18676), .ZN(n16497) );
  INV_X1 U19705 ( .A(n16488), .ZN(n16512) );
  OAI21_X1 U19706 ( .B1(P3_REIP_REG_27__SCAN_IN), .B2(n16500), .A(n16512), 
        .ZN(n16495) );
  AOI211_X1 U19707 ( .C1(P3_EBX_REG_28__SCAN_IN), .C2(n16503), .A(n16489), .B(
        n16779), .ZN(n16494) );
  AOI211_X1 U19708 ( .C1(n16492), .C2(n16491), .A(n16490), .B(n18602), .ZN(
        n16493) );
  AOI211_X1 U19709 ( .C1(P3_REIP_REG_28__SCAN_IN), .C2(n16495), .A(n16494), 
        .B(n16493), .ZN(n16496) );
  OAI211_X1 U19710 ( .C1(n17369), .C2(n16798), .A(n16497), .B(n16496), .ZN(
        P3_U2643) );
  AOI211_X1 U19711 ( .C1(n17384), .C2(n16499), .A(n16498), .B(n18602), .ZN(
        n16502) );
  OAI22_X1 U19712 ( .A1(P3_REIP_REG_27__SCAN_IN), .A2(n16500), .B1(n17389), 
        .B2(n16798), .ZN(n16501) );
  AOI211_X1 U19713 ( .C1(P3_EBX_REG_27__SCAN_IN), .C2(n16812), .A(n16502), .B(
        n16501), .ZN(n16505) );
  OAI211_X1 U19714 ( .C1(n16507), .C2(n16818), .A(n16811), .B(n16503), .ZN(
        n16504) );
  OAI211_X1 U19715 ( .C1(n16512), .C2(n18675), .A(n16505), .B(n16504), .ZN(
        P3_U2644) );
  AOI21_X1 U19716 ( .B1(n16518), .B2(P3_REIP_REG_25__SCAN_IN), .A(
        P3_REIP_REG_26__SCAN_IN), .ZN(n16513) );
  AOI22_X1 U19717 ( .A1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n16754), .B1(
        n16812), .B2(P3_EBX_REG_26__SCAN_IN), .ZN(n16511) );
  NOR2_X1 U19718 ( .A1(n16514), .A2(n16770), .ZN(n16506) );
  XNOR2_X1 U19719 ( .A(n17399), .B(n16506), .ZN(n16509) );
  AOI211_X1 U19720 ( .C1(P3_EBX_REG_26__SCAN_IN), .C2(n16519), .A(n16507), .B(
        n16779), .ZN(n16508) );
  AOI21_X1 U19721 ( .B1(n16509), .B2(n16788), .A(n16508), .ZN(n16510) );
  OAI211_X1 U19722 ( .C1(n16513), .C2(n16512), .A(n16511), .B(n16510), .ZN(
        P3_U2645) );
  AOI21_X1 U19723 ( .B1(n16536), .B2(n16782), .A(n16796), .ZN(n16545) );
  INV_X1 U19724 ( .A(n16545), .ZN(n16531) );
  AOI21_X1 U19725 ( .B1(n16782), .B2(n18669), .A(n16531), .ZN(n16523) );
  AOI211_X1 U19726 ( .C1(n17416), .C2(n16515), .A(n16514), .B(n18602), .ZN(
        n16517) );
  OAI22_X1 U19727 ( .A1(n17414), .A2(n16798), .B1(n16801), .B2(n16520), .ZN(
        n16516) );
  AOI211_X1 U19728 ( .C1(n16518), .C2(n18670), .A(n16517), .B(n16516), .ZN(
        n16522) );
  OAI211_X1 U19729 ( .C1(n16526), .C2(n16520), .A(n16811), .B(n16519), .ZN(
        n16521) );
  OAI211_X1 U19730 ( .C1(n16523), .C2(n18670), .A(n16522), .B(n16521), .ZN(
        P3_U2646) );
  NOR2_X1 U19731 ( .A1(P3_REIP_REG_24__SCAN_IN), .A2(n16802), .ZN(n16524) );
  AOI22_X1 U19732 ( .A1(n16812), .A2(P3_EBX_REG_24__SCAN_IN), .B1(n16525), 
        .B2(n16524), .ZN(n16533) );
  AOI211_X1 U19733 ( .C1(P3_EBX_REG_24__SCAN_IN), .C2(n16541), .A(n16526), .B(
        n16779), .ZN(n16530) );
  AOI211_X1 U19734 ( .C1(n17431), .C2(n16528), .A(n16527), .B(n18602), .ZN(
        n16529) );
  AOI211_X1 U19735 ( .C1(P3_REIP_REG_24__SCAN_IN), .C2(n16531), .A(n16530), 
        .B(n16529), .ZN(n16532) );
  OAI211_X1 U19736 ( .C1(n17424), .C2(n16798), .A(n16533), .B(n16532), .ZN(
        P3_U2647) );
  AOI211_X1 U19737 ( .C1(n17439), .C2(n16535), .A(n16534), .B(n18602), .ZN(
        n16540) );
  NAND2_X1 U19738 ( .A1(n16782), .A2(n16536), .ZN(n16537) );
  OAI22_X1 U19739 ( .A1(n16801), .A2(n16542), .B1(n16538), .B2(n16537), .ZN(
        n16539) );
  AOI211_X1 U19740 ( .C1(n16754), .C2(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A(
        n16540), .B(n16539), .ZN(n16544) );
  OAI211_X1 U19741 ( .C1(n16548), .C2(n16542), .A(n16811), .B(n16541), .ZN(
        n16543) );
  OAI211_X1 U19742 ( .C1(n16545), .C2(n20919), .A(n16544), .B(n16543), .ZN(
        P3_U2648) );
  NOR2_X1 U19743 ( .A1(P3_REIP_REG_22__SCAN_IN), .A2(n16802), .ZN(n16546) );
  AOI22_X1 U19744 ( .A1(n16812), .A2(P3_EBX_REG_22__SCAN_IN), .B1(n16547), 
        .B2(n16546), .ZN(n16555) );
  AOI21_X1 U19745 ( .B1(n16782), .B2(n16565), .A(n16796), .ZN(n16556) );
  OAI21_X1 U19746 ( .B1(P3_REIP_REG_21__SCAN_IN), .B2(n16802), .A(n16556), 
        .ZN(n16553) );
  AOI211_X1 U19747 ( .C1(P3_EBX_REG_22__SCAN_IN), .C2(n16561), .A(n16548), .B(
        n16779), .ZN(n16552) );
  AOI211_X1 U19748 ( .C1(n17455), .C2(n16550), .A(n16549), .B(n18602), .ZN(
        n16551) );
  AOI211_X1 U19749 ( .C1(P3_REIP_REG_22__SCAN_IN), .C2(n16553), .A(n16552), 
        .B(n16551), .ZN(n16554) );
  OAI211_X1 U19750 ( .C1(n17465), .C2(n16798), .A(n16555), .B(n16554), .ZN(
        P3_U2649) );
  NAND2_X1 U19751 ( .A1(n16782), .A2(n18663), .ZN(n16566) );
  INV_X1 U19752 ( .A(n16556), .ZN(n16573) );
  AOI211_X1 U19753 ( .C1(n17470), .C2(n16558), .A(n16557), .B(n18602), .ZN(
        n16560) );
  INV_X1 U19754 ( .A(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n17467) );
  OAI22_X1 U19755 ( .A1(n17467), .A2(n16798), .B1(n16801), .B2(n16562), .ZN(
        n16559) );
  AOI211_X1 U19756 ( .C1(n16573), .C2(P3_REIP_REG_21__SCAN_IN), .A(n16560), 
        .B(n16559), .ZN(n16564) );
  OAI211_X1 U19757 ( .C1(n16570), .C2(n16562), .A(n16811), .B(n16561), .ZN(
        n16563) );
  OAI211_X1 U19758 ( .C1(n16566), .C2(n16565), .A(n16564), .B(n16563), .ZN(
        P3_U2650) );
  INV_X1 U19759 ( .A(P3_EBX_REG_20__SCAN_IN), .ZN(n16816) );
  INV_X1 U19760 ( .A(n16567), .ZN(n16568) );
  AOI211_X1 U19761 ( .C1(n17487), .C2(n16569), .A(n16568), .B(n18602), .ZN(
        n16572) );
  AOI211_X1 U19762 ( .C1(P3_EBX_REG_20__SCAN_IN), .C2(n16579), .A(n16570), .B(
        n16779), .ZN(n16571) );
  AOI211_X1 U19763 ( .C1(n16754), .C2(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .A(
        n16572), .B(n16571), .ZN(n16576) );
  OAI221_X1 U19764 ( .B1(P3_REIP_REG_20__SCAN_IN), .B2(n16782), .C1(
        P3_REIP_REG_20__SCAN_IN), .C2(n16574), .A(n16573), .ZN(n16575) );
  OAI211_X1 U19765 ( .C1(n16816), .C2(n16801), .A(n16576), .B(n16575), .ZN(
        P3_U2651) );
  INV_X1 U19766 ( .A(n16578), .ZN(n16577) );
  AOI21_X1 U19767 ( .B1(n16782), .B2(n16577), .A(n16796), .ZN(n16603) );
  INV_X1 U19768 ( .A(P3_REIP_REG_18__SCAN_IN), .ZN(n18657) );
  NAND3_X1 U19769 ( .A1(n16782), .A2(n16578), .A3(n18657), .ZN(n16588) );
  INV_X1 U19770 ( .A(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n17509) );
  NOR2_X1 U19771 ( .A1(n17509), .A2(n16601), .ZN(n16590) );
  OAI21_X1 U19772 ( .B1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n16590), .A(
        n17449), .ZN(n17496) );
  AOI21_X1 U19773 ( .B1(n16593), .B2(n16590), .A(n16770), .ZN(n16592) );
  XNOR2_X1 U19774 ( .A(n17496), .B(n16592), .ZN(n16586) );
  INV_X1 U19775 ( .A(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n17494) );
  OAI22_X1 U19776 ( .A1(n17494), .A2(n16798), .B1(n16801), .B2(n16580), .ZN(
        n16585) );
  NAND2_X1 U19777 ( .A1(n16782), .A2(n18659), .ZN(n16582) );
  OAI211_X1 U19778 ( .C1(n16596), .C2(n16580), .A(n16811), .B(n16579), .ZN(
        n16581) );
  OAI211_X1 U19779 ( .C1(n16583), .C2(n16582), .A(n18074), .B(n16581), .ZN(
        n16584) );
  AOI211_X1 U19780 ( .C1(n16788), .C2(n16586), .A(n16585), .B(n16584), .ZN(
        n16587) );
  OAI221_X1 U19781 ( .B1(n18659), .B2(n16603), .C1(n18659), .C2(n16588), .A(
        n16587), .ZN(P3_U2652) );
  INV_X1 U19782 ( .A(n16588), .ZN(n16589) );
  AOI211_X1 U19783 ( .C1(n16812), .C2(P3_EBX_REG_18__SCAN_IN), .A(n9820), .B(
        n16589), .ZN(n16600) );
  INV_X1 U19784 ( .A(n16590), .ZN(n16591) );
  OAI21_X1 U19785 ( .B1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n17493), .A(
        n16591), .ZN(n17506) );
  INV_X1 U19786 ( .A(n16592), .ZN(n16595) );
  NAND2_X1 U19787 ( .A1(n16770), .A2(n16788), .ZN(n16792) );
  OAI221_X1 U19788 ( .B1(n17506), .B2(n16593), .C1(n17506), .C2(n17509), .A(
        n16788), .ZN(n16594) );
  AOI22_X1 U19789 ( .A1(n17506), .A2(n16595), .B1(n16792), .B2(n16594), .ZN(
        n16598) );
  AOI211_X1 U19790 ( .C1(P3_EBX_REG_18__SCAN_IN), .C2(n16605), .A(n16596), .B(
        n16779), .ZN(n16597) );
  AOI211_X1 U19791 ( .C1(n16754), .C2(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(
        n16598), .B(n16597), .ZN(n16599) );
  OAI211_X1 U19792 ( .C1(n16603), .C2(n18657), .A(n16600), .B(n16599), .ZN(
        P3_U2653) );
  NOR2_X1 U19793 ( .A1(n17745), .A2(n17517), .ZN(n16616) );
  OAI21_X1 U19794 ( .B1(P3_PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n16616), .A(
        n16601), .ZN(n17523) );
  NOR2_X1 U19795 ( .A1(n17745), .A2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n16789) );
  INV_X1 U19796 ( .A(n16789), .ZN(n16757) );
  OAI21_X1 U19797 ( .B1(n17517), .B2(n16757), .A(n16797), .ZN(n16602) );
  XOR2_X1 U19798 ( .A(n17523), .B(n16602), .Z(n16610) );
  AOI221_X1 U19799 ( .B1(n16802), .B2(n18655), .C1(n16604), .C2(n18655), .A(
        n16603), .ZN(n16609) );
  OAI211_X1 U19800 ( .C1(n16619), .C2(n16612), .A(n16811), .B(n16605), .ZN(
        n16606) );
  OAI21_X1 U19801 ( .B1(n16798), .B2(n16607), .A(n16606), .ZN(n16608) );
  AOI211_X1 U19802 ( .C1(n16788), .C2(n16610), .A(n16609), .B(n16608), .ZN(
        n16611) );
  OAI211_X1 U19803 ( .C1(n16801), .C2(n16612), .A(n16611), .B(n18074), .ZN(
        P3_U2654) );
  NOR2_X1 U19804 ( .A1(P3_REIP_REG_16__SCAN_IN), .A2(n16802), .ZN(n16613) );
  AOI22_X1 U19805 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n16754), .B1(
        n16614), .B2(n16613), .ZN(n16626) );
  INV_X1 U19806 ( .A(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n16617) );
  AOI21_X1 U19807 ( .B1(n16617), .B2(n16627), .A(n16616), .ZN(n17535) );
  INV_X1 U19808 ( .A(n17535), .ZN(n16618) );
  AOI221_X1 U19809 ( .B1(n16615), .B2(n17535), .C1(n10184), .C2(n16618), .A(
        n18602), .ZN(n16621) );
  AOI211_X1 U19810 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16631), .A(n16619), .B(
        n16779), .ZN(n16620) );
  AOI211_X1 U19811 ( .C1(P3_EBX_REG_16__SCAN_IN), .C2(n16812), .A(n16621), .B(
        n16620), .ZN(n16625) );
  INV_X1 U19812 ( .A(n16622), .ZN(n16639) );
  OAI21_X1 U19813 ( .B1(n16639), .B2(n16802), .A(n16810), .ZN(n16641) );
  NAND3_X1 U19814 ( .A1(n18651), .A2(n16782), .A3(n16639), .ZN(n16634) );
  INV_X1 U19815 ( .A(n16634), .ZN(n16623) );
  OAI21_X1 U19816 ( .B1(n16641), .B2(n16623), .A(P3_REIP_REG_16__SCAN_IN), 
        .ZN(n16624) );
  NAND4_X1 U19817 ( .A1(n16626), .A2(n16625), .A3(n18074), .A4(n16624), .ZN(
        P3_U2655) );
  OAI21_X1 U19818 ( .B1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .B2(n17534), .A(
        n16627), .ZN(n17545) );
  INV_X1 U19819 ( .A(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n17548) );
  INV_X1 U19820 ( .A(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n16800) );
  OAI221_X1 U19821 ( .B1(n17545), .B2(n17548), .C1(n17545), .C2(n16800), .A(
        n16788), .ZN(n16628) );
  AOI22_X1 U19822 ( .A1(n10184), .A2(n17545), .B1(n16792), .B2(n16628), .ZN(
        n16630) );
  OAI22_X1 U19823 ( .A1(n17548), .A2(n16798), .B1(n16801), .B2(n16632), .ZN(
        n16629) );
  AOI211_X1 U19824 ( .C1(n16641), .C2(P3_REIP_REG_15__SCAN_IN), .A(n16630), 
        .B(n16629), .ZN(n16635) );
  OAI211_X1 U19825 ( .C1(n16636), .C2(n16632), .A(n16811), .B(n16631), .ZN(
        n16633) );
  NAND4_X1 U19826 ( .A1(n16635), .A2(n18074), .A3(n16634), .A4(n16633), .ZN(
        P3_U2656) );
  AOI211_X1 U19827 ( .C1(P3_EBX_REG_14__SCAN_IN), .C2(n16653), .A(n16636), .B(
        n16779), .ZN(n16637) );
  AOI21_X1 U19828 ( .B1(n16754), .B2(P3_PHYADDRPOINTER_REG_14__SCAN_IN), .A(
        n16637), .ZN(n16645) );
  NAND2_X1 U19829 ( .A1(n16782), .A2(n16638), .ZN(n16649) );
  NOR2_X1 U19830 ( .A1(n16639), .A2(n16649), .ZN(n16640) );
  AOI22_X1 U19831 ( .A1(n16812), .A2(P3_EBX_REG_14__SCAN_IN), .B1(
        P3_REIP_REG_13__SCAN_IN), .B2(n16640), .ZN(n16644) );
  AOI21_X1 U19832 ( .B1(n17561), .B2(n16646), .A(n17534), .ZN(n17563) );
  NAND2_X1 U19833 ( .A1(n17558), .A2(n16789), .ZN(n16710) );
  INV_X1 U19834 ( .A(n16710), .ZN(n16696) );
  NAND2_X1 U19835 ( .A1(n17559), .A2(n16696), .ZN(n16660) );
  OAI21_X1 U19836 ( .B1(n17583), .B2(n16660), .A(n16797), .ZN(n16647) );
  XNOR2_X1 U19837 ( .A(n17563), .B(n16647), .ZN(n16642) );
  AOI22_X1 U19838 ( .A1(n16788), .A2(n16642), .B1(P3_REIP_REG_14__SCAN_IN), 
        .B2(n16641), .ZN(n16643) );
  NAND4_X1 U19839 ( .A1(n16645), .A2(n16644), .A3(n16643), .A4(n18074), .ZN(
        P3_U2657) );
  INV_X1 U19840 ( .A(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n16657) );
  AOI21_X1 U19841 ( .B1(n16782), .B2(n16665), .A(n16796), .ZN(n16675) );
  NAND2_X1 U19842 ( .A1(n16782), .A2(n18645), .ZN(n16666) );
  INV_X1 U19843 ( .A(P3_REIP_REG_13__SCAN_IN), .ZN(n18647) );
  AOI21_X1 U19844 ( .B1(n16675), .B2(n16666), .A(n18647), .ZN(n16652) );
  INV_X1 U19845 ( .A(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n17594) );
  NOR2_X1 U19846 ( .A1(n17594), .A2(n17571), .ZN(n16659) );
  OAI21_X1 U19847 ( .B1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n16659), .A(
        n16646), .ZN(n16648) );
  INV_X1 U19848 ( .A(n16648), .ZN(n17574) );
  AOI21_X1 U19849 ( .B1(n16659), .B2(n16800), .A(n16770), .ZN(n16661) );
  AOI221_X1 U19850 ( .B1(n17574), .B2(n16661), .C1(n16648), .C2(n16647), .A(
        n18602), .ZN(n16651) );
  OAI22_X1 U19851 ( .A1(P3_REIP_REG_13__SCAN_IN), .A2(n16649), .B1(n16801), 
        .B2(n16654), .ZN(n16650) );
  NOR4_X1 U19852 ( .A1(n9820), .A2(n16652), .A3(n16651), .A4(n16650), .ZN(
        n16656) );
  OAI211_X1 U19853 ( .C1(n16658), .C2(n16654), .A(n16811), .B(n16653), .ZN(
        n16655) );
  OAI211_X1 U19854 ( .C1(n16798), .C2(n16657), .A(n16656), .B(n16655), .ZN(
        P3_U2658) );
  AOI211_X1 U19855 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16678), .A(n16658), .B(
        n16779), .ZN(n16668) );
  AOI21_X1 U19856 ( .B1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n16754), .A(
        n9820), .ZN(n16664) );
  INV_X1 U19857 ( .A(n16792), .ZN(n16756) );
  AOI21_X1 U19858 ( .B1(n17594), .B2(n17571), .A(n16659), .ZN(n17592) );
  AOI21_X1 U19859 ( .B1(n17592), .B2(n16660), .A(n18602), .ZN(n16662) );
  OAI22_X1 U19860 ( .A1(n16756), .A2(n16662), .B1(n17592), .B2(n16661), .ZN(
        n16663) );
  OAI211_X1 U19861 ( .C1(n16666), .C2(n16665), .A(n16664), .B(n16663), .ZN(
        n16667) );
  AOI211_X1 U19862 ( .C1(P3_EBX_REG_12__SCAN_IN), .C2(n16812), .A(n16668), .B(
        n16667), .ZN(n16669) );
  OAI21_X1 U19863 ( .B1(n16675), .B2(n18645), .A(n16669), .ZN(P3_U2659) );
  INV_X1 U19864 ( .A(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n16682) );
  NOR2_X1 U19865 ( .A1(n16802), .A2(n16670), .ZN(n16740) );
  NAND2_X1 U19866 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16740), .ZN(n16686) );
  INV_X1 U19867 ( .A(n16686), .ZN(n16725) );
  AOI21_X1 U19868 ( .B1(n16671), .B2(n16725), .A(P3_REIP_REG_11__SCAN_IN), 
        .ZN(n16676) );
  NAND2_X1 U19869 ( .A1(n17609), .A2(n16718), .ZN(n16694) );
  NOR2_X1 U19870 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n16694), .ZN(
        n16672) );
  AOI21_X1 U19871 ( .B1(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n16672), .A(
        n16770), .ZN(n16673) );
  INV_X1 U19872 ( .A(P3_PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n17618) );
  NOR2_X1 U19873 ( .A1(n17618), .A2(n16694), .ZN(n16685) );
  OAI21_X1 U19874 ( .B1(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n16685), .A(
        n17571), .ZN(n17613) );
  XOR2_X1 U19875 ( .A(n16673), .B(n17613), .Z(n16674) );
  OAI22_X1 U19876 ( .A1(n16676), .A2(n16675), .B1(n18602), .B2(n16674), .ZN(
        n16677) );
  AOI211_X1 U19877 ( .C1(n16812), .C2(P3_EBX_REG_11__SCAN_IN), .A(n9820), .B(
        n16677), .ZN(n16681) );
  OAI211_X1 U19878 ( .C1(n16683), .C2(n16679), .A(n16811), .B(n16678), .ZN(
        n16680) );
  OAI211_X1 U19879 ( .C1(n16798), .C2(n16682), .A(n16681), .B(n16680), .ZN(
        P3_U2660) );
  AOI211_X1 U19880 ( .C1(P3_EBX_REG_10__SCAN_IN), .C2(n16699), .A(n16683), .B(
        n16779), .ZN(n16684) );
  AOI211_X1 U19881 ( .C1(n16812), .C2(P3_EBX_REG_10__SCAN_IN), .A(n9820), .B(
        n16684), .ZN(n16693) );
  AOI21_X1 U19882 ( .B1(n17618), .B2(n16694), .A(n16685), .ZN(n17621) );
  OAI21_X1 U19883 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16694), .A(
        n16797), .ZN(n16698) );
  XNOR2_X1 U19884 ( .A(n17621), .B(n16698), .ZN(n16691) );
  INV_X1 U19885 ( .A(P3_REIP_REG_6__SCAN_IN), .ZN(n21078) );
  INV_X1 U19886 ( .A(P3_REIP_REG_7__SCAN_IN), .ZN(n18636) );
  NOR3_X1 U19887 ( .A1(n21078), .A2(n18636), .A3(n16686), .ZN(n16714) );
  NAND2_X1 U19888 ( .A1(P3_REIP_REG_8__SCAN_IN), .A2(n16714), .ZN(n16705) );
  XOR2_X1 U19889 ( .A(P3_REIP_REG_10__SCAN_IN), .B(n18640), .Z(n16689) );
  NAND2_X1 U19890 ( .A1(n16687), .A2(n16810), .ZN(n16720) );
  NAND2_X1 U19891 ( .A1(n16802), .A2(n16810), .ZN(n16809) );
  OAI21_X1 U19892 ( .B1(n16688), .B2(n16720), .A(n16809), .ZN(n16708) );
  OAI22_X1 U19893 ( .A1(n16705), .A2(n16689), .B1(n18641), .B2(n16708), .ZN(
        n16690) );
  AOI21_X1 U19894 ( .B1(n16788), .B2(n16691), .A(n16690), .ZN(n16692) );
  OAI211_X1 U19895 ( .C1(n17618), .C2(n16798), .A(n16693), .B(n16692), .ZN(
        P3_U2661) );
  INV_X1 U19896 ( .A(n16718), .ZN(n16709) );
  NOR2_X1 U19897 ( .A1(n21012), .A2(n16709), .ZN(n16695) );
  OAI21_X1 U19898 ( .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n16695), .A(
        n16694), .ZN(n17636) );
  OAI221_X1 U19899 ( .B1(n17636), .B2(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .C1(
        n17636), .C2(n16696), .A(n16788), .ZN(n16697) );
  OAI22_X1 U19900 ( .A1(n17636), .A2(n16792), .B1(n16698), .B2(n16697), .ZN(
        n16703) );
  OAI211_X1 U19901 ( .C1(n16706), .C2(n16701), .A(n16811), .B(n16699), .ZN(
        n16700) );
  OAI211_X1 U19902 ( .C1(n16801), .C2(n16701), .A(n18074), .B(n16700), .ZN(
        n16702) );
  AOI211_X1 U19903 ( .C1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .C2(n16754), .A(
        n16703), .B(n16702), .ZN(n16704) );
  OAI221_X1 U19904 ( .B1(P3_REIP_REG_9__SCAN_IN), .B2(n16705), .C1(n18640), 
        .C2(n16708), .A(n16704), .ZN(P3_U2662) );
  AOI211_X1 U19905 ( .C1(P3_EBX_REG_8__SCAN_IN), .C2(n16721), .A(n16706), .B(
        n16779), .ZN(n16707) );
  AOI211_X1 U19906 ( .C1(n16812), .C2(P3_EBX_REG_8__SCAN_IN), .A(n9820), .B(
        n16707), .ZN(n16717) );
  INV_X1 U19907 ( .A(n16708), .ZN(n16715) );
  INV_X1 U19908 ( .A(P3_REIP_REG_8__SCAN_IN), .ZN(n18638) );
  AOI22_X1 U19909 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(n16709), .B1(
        n16718), .B2(n21012), .ZN(n17658) );
  NAND2_X1 U19910 ( .A1(n16797), .A2(n16710), .ZN(n16712) );
  OAI21_X1 U19911 ( .B1(n17658), .B2(n16712), .A(n16788), .ZN(n16711) );
  AOI21_X1 U19912 ( .B1(n17658), .B2(n16712), .A(n16711), .ZN(n16713) );
  AOI221_X1 U19913 ( .B1(n16715), .B2(P3_REIP_REG_8__SCAN_IN), .C1(n16714), 
        .C2(n18638), .A(n16713), .ZN(n16716) );
  OAI211_X1 U19914 ( .C1(n21012), .C2(n16798), .A(n16717), .B(n16716), .ZN(
        P3_U2663) );
  AOI21_X1 U19915 ( .B1(n17665), .B2(n16731), .A(n16718), .ZN(n17670) );
  OAI21_X1 U19916 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16731), .A(
        n16797), .ZN(n16719) );
  XOR2_X1 U19917 ( .A(n17670), .B(n16719), .Z(n16728) );
  NAND2_X1 U19918 ( .A1(n16809), .A2(n16720), .ZN(n16744) );
  NAND2_X1 U19919 ( .A1(n16725), .A2(n21078), .ZN(n16737) );
  AOI21_X1 U19920 ( .B1(n16744), .B2(n16737), .A(n18636), .ZN(n16724) );
  OAI211_X1 U19921 ( .C1(n16730), .C2(n17080), .A(n16811), .B(n16721), .ZN(
        n16722) );
  OAI211_X1 U19922 ( .C1(n16801), .C2(n17080), .A(n18074), .B(n16722), .ZN(
        n16723) );
  AOI211_X1 U19923 ( .C1(n16754), .C2(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n16724), .B(n16723), .ZN(n16727) );
  NAND3_X1 U19924 ( .A1(P3_REIP_REG_6__SCAN_IN), .A2(n16725), .A3(n18636), 
        .ZN(n16726) );
  OAI211_X1 U19925 ( .C1(n16728), .C2(n18602), .A(n16727), .B(n16726), .ZN(
        P3_U2664) );
  NAND2_X1 U19926 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n16729) );
  NOR2_X1 U19927 ( .A1(n17745), .A2(n16729), .ZN(n16769) );
  NAND2_X1 U19928 ( .A1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A2(n16769), .ZN(
        n16755) );
  NOR2_X1 U19929 ( .A1(n17693), .A2(n16755), .ZN(n16741) );
  OAI21_X1 U19930 ( .B1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n16741), .A(
        n16731), .ZN(n17687) );
  OAI221_X1 U19931 ( .B1(n16770), .B2(n16741), .C1(n16770), .C2(n16800), .A(
        n16788), .ZN(n16739) );
  AOI211_X1 U19932 ( .C1(P3_EBX_REG_6__SCAN_IN), .C2(n16747), .A(n16730), .B(
        n16779), .ZN(n16736) );
  OAI21_X1 U19933 ( .B1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n16731), .A(
        n17687), .ZN(n16732) );
  OAI22_X1 U19934 ( .A1(n21078), .A2(n16744), .B1(n16799), .B2(n16732), .ZN(
        n16735) );
  AOI22_X1 U19935 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n16754), .B1(
        n16812), .B2(P3_EBX_REG_6__SCAN_IN), .ZN(n16733) );
  INV_X1 U19936 ( .A(n16733), .ZN(n16734) );
  NOR4_X1 U19937 ( .A1(n9820), .A2(n16736), .A3(n16735), .A4(n16734), .ZN(
        n16738) );
  OAI211_X1 U19938 ( .C1(n17687), .C2(n16739), .A(n16738), .B(n16737), .ZN(
        P3_U2665) );
  NOR2_X1 U19939 ( .A1(P3_REIP_REG_5__SCAN_IN), .A2(n16740), .ZN(n16745) );
  AOI21_X1 U19940 ( .B1(n17693), .B2(n16755), .A(n16741), .ZN(n16742) );
  INV_X1 U19941 ( .A(n16742), .ZN(n17699) );
  OAI21_X1 U19942 ( .B1(n17694), .B2(n16757), .A(n16797), .ZN(n16758) );
  XNOR2_X1 U19943 ( .A(n17699), .B(n16758), .ZN(n16743) );
  OAI22_X1 U19944 ( .A1(n16745), .A2(n16744), .B1(n18602), .B2(n16743), .ZN(
        n16746) );
  AOI211_X1 U19945 ( .C1(n16812), .C2(P3_EBX_REG_5__SCAN_IN), .A(n9820), .B(
        n16746), .ZN(n16750) );
  OAI211_X1 U19946 ( .C1(n16751), .C2(n16748), .A(n16811), .B(n16747), .ZN(
        n16749) );
  OAI211_X1 U19947 ( .C1(n16798), .C2(n17693), .A(n16750), .B(n16749), .ZN(
        P3_U2666) );
  AOI211_X1 U19948 ( .C1(P3_EBX_REG_4__SCAN_IN), .C2(n16775), .A(n16751), .B(
        n16779), .ZN(n16753) );
  NOR2_X1 U19949 ( .A1(n18746), .A2(n18759), .ZN(n16808) );
  INV_X1 U19950 ( .A(n16808), .ZN(n18761) );
  OAI221_X1 U19951 ( .B1(n18761), .B2(n11658), .C1(n18761), .C2(n18539), .A(
        n18074), .ZN(n16752) );
  AOI211_X1 U19952 ( .C1(n16754), .C2(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .A(
        n16753), .B(n16752), .ZN(n16764) );
  OAI21_X1 U19953 ( .B1(P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n16769), .A(
        n16755), .ZN(n17711) );
  INV_X1 U19954 ( .A(n17711), .ZN(n16759) );
  AOI22_X1 U19955 ( .A1(n16812), .A2(P3_EBX_REG_4__SCAN_IN), .B1(n16759), .B2(
        n16756), .ZN(n16763) );
  INV_X1 U19956 ( .A(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n17720) );
  INV_X1 U19957 ( .A(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n21053) );
  OR3_X1 U19958 ( .A1(n17720), .A2(n21053), .A3(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n17703) );
  OAI22_X1 U19959 ( .A1(n16759), .A2(n16758), .B1(n16757), .B2(n17703), .ZN(
        n16760) );
  OAI21_X1 U19960 ( .B1(n16766), .B2(n16802), .A(n16810), .ZN(n16768) );
  AOI22_X1 U19961 ( .A1(n16788), .A2(n16760), .B1(P3_REIP_REG_4__SCAN_IN), 
        .B2(n16768), .ZN(n16762) );
  INV_X1 U19962 ( .A(P3_REIP_REG_4__SCAN_IN), .ZN(n18631) );
  NAND3_X1 U19963 ( .A1(n16782), .A2(n16766), .A3(n18631), .ZN(n16761) );
  NAND4_X1 U19964 ( .A1(n16764), .A2(n16763), .A3(n16762), .A4(n16761), .ZN(
        P3_U2667) );
  NOR2_X1 U19965 ( .A1(n18727), .A2(n18557), .ZN(n18547) );
  INV_X1 U19966 ( .A(n18547), .ZN(n16765) );
  AOI21_X1 U19967 ( .B1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n16765), .A(
        n17019), .ZN(n18697) );
  OR2_X1 U19968 ( .A1(n16802), .A2(n16766), .ZN(n16767) );
  OAI22_X1 U19969 ( .A1(n18697), .A2(n18761), .B1(n16781), .B2(n16767), .ZN(
        n16774) );
  INV_X1 U19970 ( .A(n16768), .ZN(n16772) );
  NAND2_X1 U19971 ( .A1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n16778) );
  AOI21_X1 U19972 ( .B1(n17720), .B2(n16778), .A(n16769), .ZN(n17718) );
  AOI21_X1 U19973 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(n16789), .A(
        n16770), .ZN(n16787) );
  XNOR2_X1 U19974 ( .A(n17718), .B(n16787), .ZN(n16771) );
  OAI22_X1 U19975 ( .A1(n16772), .A2(n18629), .B1(n18602), .B2(n16771), .ZN(
        n16773) );
  AOI211_X1 U19976 ( .C1(n16812), .C2(P3_EBX_REG_3__SCAN_IN), .A(n16774), .B(
        n16773), .ZN(n16777) );
  OAI211_X1 U19977 ( .C1(n16780), .C2(n17091), .A(n16811), .B(n16775), .ZN(
        n16776) );
  OAI211_X1 U19978 ( .C1(n16798), .C2(n17720), .A(n16777), .B(n16776), .ZN(
        P3_U2668) );
  OAI21_X1 U19979 ( .B1(P3_PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A(n16778), .ZN(n17735) );
  NAND2_X1 U19980 ( .A1(n17105), .A2(n17103), .ZN(n16794) );
  AOI211_X1 U19981 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16794), .A(n16780), .B(
        n16779), .ZN(n16786) );
  AOI21_X1 U19982 ( .B1(n18713), .B2(n18563), .A(n18547), .ZN(n18709) );
  AOI22_X1 U19983 ( .A1(P3_REIP_REG_2__SCAN_IN), .A2(n16796), .B1(n18709), 
        .B2(n16808), .ZN(n16784) );
  OAI211_X1 U19984 ( .C1(P3_REIP_REG_1__SCAN_IN), .C2(P3_REIP_REG_2__SCAN_IN), 
        .A(n16782), .B(n16781), .ZN(n16783) );
  OAI211_X1 U19985 ( .C1(n16798), .C2(n21053), .A(n16784), .B(n16783), .ZN(
        n16785) );
  AOI211_X1 U19986 ( .C1(P3_EBX_REG_2__SCAN_IN), .C2(n16812), .A(n16786), .B(
        n16785), .ZN(n16791) );
  OAI211_X1 U19987 ( .C1(n16789), .C2(n17735), .A(n16788), .B(n16787), .ZN(
        n16790) );
  OAI211_X1 U19988 ( .C1(n16792), .C2(n17735), .A(n16791), .B(n16790), .ZN(
        P3_U2669) );
  NAND2_X1 U19989 ( .A1(n18563), .A2(n16793), .ZN(n18714) );
  INV_X1 U19990 ( .A(n16794), .ZN(n16795) );
  NOR2_X1 U19991 ( .A1(n16795), .A2(n17097), .ZN(n17100) );
  AOI22_X1 U19992 ( .A1(n16811), .A2(n17100), .B1(P3_REIP_REG_1__SCAN_IN), 
        .B2(n16796), .ZN(n16807) );
  AOI21_X1 U19993 ( .B1(n16797), .B2(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A(
        n18602), .ZN(n16805) );
  OAI21_X1 U19994 ( .B1(n16800), .B2(n16799), .A(n16798), .ZN(n16804) );
  OAI22_X1 U19995 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(n16802), .B1(n16801), 
        .B2(n17103), .ZN(n16803) );
  AOI221_X1 U19996 ( .B1(n16805), .B2(n17745), .C1(n16804), .C2(
        P3_PHYADDRPOINTER_REG_1__SCAN_IN), .A(n16803), .ZN(n16806) );
  OAI211_X1 U19997 ( .C1(n18714), .C2(n18761), .A(n16807), .B(n16806), .ZN(
        P3_U2670) );
  AOI22_X1 U19998 ( .A1(P3_REIP_REG_0__SCAN_IN), .A2(n16809), .B1(n16808), 
        .B2(n18727), .ZN(n16815) );
  NAND3_X1 U19999 ( .A1(P3_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18757), .A3(
        n16810), .ZN(n16814) );
  OAI21_X1 U20000 ( .B1(n16812), .B2(n16811), .A(P3_EBX_REG_0__SCAN_IN), .ZN(
        n16813) );
  NAND3_X1 U20001 ( .A1(n16815), .A2(n16814), .A3(n16813), .ZN(P3_U2671) );
  NOR2_X1 U20002 ( .A1(n16816), .A2(n16935), .ZN(n16898) );
  NAND4_X1 U20003 ( .A1(P3_EBX_REG_24__SCAN_IN), .A2(P3_EBX_REG_23__SCAN_IN), 
        .A3(P3_EBX_REG_22__SCAN_IN), .A4(P3_EBX_REG_21__SCAN_IN), .ZN(n16817)
         );
  NOR4_X1 U20004 ( .A1(n16856), .A2(n16819), .A3(n16818), .A4(n16817), .ZN(
        n16820) );
  NAND4_X1 U20005 ( .A1(P3_EBX_REG_26__SCAN_IN), .A2(P3_EBX_REG_25__SCAN_IN), 
        .A3(n16898), .A4(n16820), .ZN(n16845) );
  NOR2_X1 U20006 ( .A1(n16846), .A2(n16845), .ZN(n16844) );
  NAND2_X1 U20007 ( .A1(n17109), .A2(P3_EBX_REG_31__SCAN_IN), .ZN(n16822) );
  NAND2_X1 U20008 ( .A1(n16844), .A2(n18134), .ZN(n16821) );
  OAI22_X1 U20009 ( .A1(n16844), .A2(n16822), .B1(P3_EBX_REG_31__SCAN_IN), 
        .B2(n16821), .ZN(P3_U2672) );
  AOI22_X1 U20010 ( .A1(n9841), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(n9815), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16826) );
  AOI22_X1 U20011 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n16825) );
  AOI22_X1 U20012 ( .A1(n9810), .A2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .B1(n9819), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16824) );
  AOI22_X1 U20013 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16823) );
  NAND4_X1 U20014 ( .A1(n16826), .A2(n16825), .A3(n16824), .A4(n16823), .ZN(
        n16832) );
  AOI22_X1 U20015 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n16830) );
  AOI22_X1 U20016 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n9845), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16829) );
  AOI22_X1 U20017 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n16828) );
  AOI22_X1 U20018 ( .A1(n17048), .A2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .B1(
        n9842), .B2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n16827) );
  NAND4_X1 U20019 ( .A1(n16830), .A2(n16829), .A3(n16828), .A4(n16827), .ZN(
        n16831) );
  NOR2_X1 U20020 ( .A1(n16832), .A2(n16831), .ZN(n16843) );
  AOI22_X1 U20021 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n16836) );
  AOI22_X1 U20022 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .B1(
        n9819), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16835) );
  AOI22_X1 U20023 ( .A1(n9816), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16834) );
  AOI22_X1 U20024 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n16833) );
  NAND4_X1 U20025 ( .A1(n16836), .A2(n16835), .A3(n16834), .A4(n16833), .ZN(
        n16842) );
  AOI22_X1 U20026 ( .A1(n9841), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n9811), .B2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n16840) );
  AOI22_X1 U20027 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n17024), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16839) );
  AOI22_X1 U20028 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16838) );
  AOI22_X1 U20029 ( .A1(n11857), .A2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .B1(
        n9846), .B2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n16837) );
  NAND4_X1 U20030 ( .A1(n16840), .A2(n16839), .A3(n16838), .A4(n16837), .ZN(
        n16841) );
  NOR2_X1 U20031 ( .A1(n16842), .A2(n16841), .ZN(n16852) );
  NOR2_X1 U20032 ( .A1(n16852), .A2(n16851), .ZN(n16850) );
  XNOR2_X1 U20033 ( .A(n16843), .B(n16850), .ZN(n17114) );
  AOI211_X1 U20034 ( .C1(n16846), .C2(n16845), .A(n16844), .B(n17101), .ZN(
        n16847) );
  AOI21_X1 U20035 ( .B1(n17101), .B2(n17114), .A(n16847), .ZN(n16848) );
  INV_X1 U20036 ( .A(n16848), .ZN(P3_U2673) );
  INV_X1 U20037 ( .A(n16849), .ZN(n16855) );
  AOI21_X1 U20038 ( .B1(n16852), .B2(n16851), .A(n16850), .ZN(n17119) );
  AOI22_X1 U20039 ( .A1(n17101), .A2(n17119), .B1(n16853), .B2(n16856), .ZN(
        n16854) );
  OAI21_X1 U20040 ( .B1(n16856), .B2(n16855), .A(n16854), .ZN(P3_U2674) );
  INV_X1 U20041 ( .A(n16857), .ZN(n16866) );
  AOI21_X1 U20042 ( .B1(P3_EBX_REG_27__SCAN_IN), .B2(n17109), .A(n16866), .ZN(
        n16861) );
  AOI21_X1 U20043 ( .B1(n16859), .B2(n16863), .A(n16858), .ZN(n17128) );
  INV_X1 U20044 ( .A(n17128), .ZN(n16860) );
  OAI22_X1 U20045 ( .A1(n16862), .A2(n16861), .B1(n16860), .B2(n17109), .ZN(
        P3_U2676) );
  AOI21_X1 U20046 ( .B1(P3_EBX_REG_26__SCAN_IN), .B2(n17109), .A(n16872), .ZN(
        n16865) );
  OAI21_X1 U20047 ( .B1(n16868), .B2(n16864), .A(n16863), .ZN(n17137) );
  OAI22_X1 U20048 ( .A1(n16866), .A2(n16865), .B1(n17137), .B2(n17109), .ZN(
        P3_U2677) );
  INV_X1 U20049 ( .A(n16867), .ZN(n16876) );
  AOI21_X1 U20050 ( .B1(P3_EBX_REG_25__SCAN_IN), .B2(n17109), .A(n16876), .ZN(
        n16871) );
  AOI21_X1 U20051 ( .B1(n16869), .B2(n16873), .A(n16868), .ZN(n17138) );
  INV_X1 U20052 ( .A(n17138), .ZN(n16870) );
  OAI22_X1 U20053 ( .A1(n16872), .A2(n16871), .B1(n16870), .B2(n17109), .ZN(
        P3_U2678) );
  AOI21_X1 U20054 ( .B1(P3_EBX_REG_24__SCAN_IN), .B2(n17109), .A(n16883), .ZN(
        n16875) );
  OAI21_X1 U20055 ( .B1(n16878), .B2(n16874), .A(n16873), .ZN(n17147) );
  OAI22_X1 U20056 ( .A1(n16876), .A2(n16875), .B1(n17147), .B2(n17109), .ZN(
        P3_U2679) );
  INV_X1 U20057 ( .A(n16877), .ZN(n16897) );
  AOI21_X1 U20058 ( .B1(P3_EBX_REG_23__SCAN_IN), .B2(n17109), .A(n16897), .ZN(
        n16882) );
  AOI21_X1 U20059 ( .B1(n16880), .B2(n16879), .A(n16878), .ZN(n17148) );
  INV_X1 U20060 ( .A(n17148), .ZN(n16881) );
  OAI22_X1 U20061 ( .A1(n16883), .A2(n16882), .B1(n16881), .B2(n17109), .ZN(
        P3_U2680) );
  AOI21_X1 U20062 ( .B1(P3_EBX_REG_22__SCAN_IN), .B2(n17109), .A(n16884), .ZN(
        n16896) );
  AOI22_X1 U20063 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n16894) );
  AOI22_X1 U20064 ( .A1(n9838), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(n9829), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16893) );
  AOI22_X1 U20065 ( .A1(n9822), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9842), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16885) );
  OAI21_X1 U20066 ( .B1(n11658), .B2(n20918), .A(n16885), .ZN(n16891) );
  AOI22_X1 U20067 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n16889) );
  AOI22_X1 U20068 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16888) );
  AOI22_X1 U20069 ( .A1(n9845), .A2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        n9816), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16887) );
  AOI22_X1 U20070 ( .A1(n15640), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16886) );
  NAND4_X1 U20071 ( .A1(n16889), .A2(n16888), .A3(n16887), .A4(n16886), .ZN(
        n16890) );
  AOI211_X1 U20072 ( .C1(n17019), .C2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A(
        n16891), .B(n16890), .ZN(n16892) );
  NAND3_X1 U20073 ( .A1(n16894), .A2(n16893), .A3(n16892), .ZN(n17154) );
  INV_X1 U20074 ( .A(n17154), .ZN(n16895) );
  OAI22_X1 U20075 ( .A1(n16897), .A2(n16896), .B1(n16895), .B2(n17109), .ZN(
        P3_U2681) );
  NOR2_X1 U20076 ( .A1(n17101), .A2(n16898), .ZN(n16922) );
  AOI22_X1 U20077 ( .A1(n9809), .A2(P3_INSTQUEUE_REG_4__5__SCAN_IN), .B1(n9832), .B2(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n16902) );
  AOI22_X1 U20078 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_14__5__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n16901) );
  AOI22_X1 U20079 ( .A1(n9811), .A2(P3_INSTQUEUE_REG_2__5__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n16900) );
  AOI22_X1 U20080 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_7__5__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n16899) );
  NAND4_X1 U20081 ( .A1(n16902), .A2(n16901), .A3(n16900), .A4(n16899), .ZN(
        n16908) );
  AOI22_X1 U20082 ( .A1(n9841), .A2(P3_INSTQUEUE_REG_8__5__SCAN_IN), .B1(n9815), .B2(P3_INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n16906) );
  AOI22_X1 U20083 ( .A1(n9838), .A2(P3_INSTQUEUE_REG_9__5__SCAN_IN), .B1(n9812), .B2(P3_INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n16905) );
  AOI22_X1 U20084 ( .A1(n17048), .A2(P3_INSTQUEUE_REG_15__5__SCAN_IN), .B1(
        n9846), .B2(P3_INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n16904) );
  AOI22_X1 U20085 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_10__5__SCAN_IN), .B1(
        n17069), .B2(P3_INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n16903) );
  NAND4_X1 U20086 ( .A1(n16906), .A2(n16905), .A3(n16904), .A4(n16903), .ZN(
        n16907) );
  NOR2_X1 U20087 ( .A1(n16908), .A2(n16907), .ZN(n17162) );
  INV_X1 U20088 ( .A(n17162), .ZN(n16909) );
  AOI22_X1 U20089 ( .A1(P3_EBX_REG_21__SCAN_IN), .A2(n16922), .B1(n17101), 
        .B2(n16909), .ZN(n16910) );
  OAI21_X1 U20090 ( .B1(P3_EBX_REG_21__SCAN_IN), .B2(n16911), .A(n16910), .ZN(
        P3_U2682) );
  AOI22_X1 U20091 ( .A1(n17048), .A2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n16915) );
  AOI22_X1 U20092 ( .A1(n9838), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n16914) );
  AOI22_X1 U20093 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .B1(
        n9816), .B2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n16913) );
  AOI22_X1 U20094 ( .A1(n11857), .A2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n16912) );
  NAND4_X1 U20095 ( .A1(n16915), .A2(n16914), .A3(n16913), .A4(n16912), .ZN(
        n16921) );
  AOI22_X1 U20096 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .B1(n9846), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n16919) );
  AOI22_X1 U20097 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .B1(
        n9819), .B2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n16918) );
  AOI22_X1 U20098 ( .A1(n9841), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(n9811), .B2(P3_INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n16917) );
  AOI22_X1 U20099 ( .A1(n17069), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(
        n9832), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n16916) );
  NAND4_X1 U20100 ( .A1(n16919), .A2(n16918), .A3(n16917), .A4(n16916), .ZN(
        n16920) );
  NOR2_X1 U20101 ( .A1(n16921), .A2(n16920), .ZN(n17169) );
  OAI21_X1 U20102 ( .B1(P3_EBX_REG_20__SCAN_IN), .B2(n16923), .A(n16922), .ZN(
        n16924) );
  OAI21_X1 U20103 ( .B1(n17169), .B2(n17109), .A(n16924), .ZN(P3_U2683) );
  AOI22_X1 U20104 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n9846), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n16928) );
  AOI22_X1 U20105 ( .A1(n9841), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(n9816), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n16927) );
  AOI22_X1 U20106 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n16926) );
  AOI22_X1 U20107 ( .A1(n17048), .A2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n16925) );
  NAND4_X1 U20108 ( .A1(n16928), .A2(n16927), .A3(n16926), .A4(n16925), .ZN(
        n16934) );
  AOI22_X1 U20109 ( .A1(n17049), .A2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .B1(
        n9832), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n16932) );
  AOI22_X1 U20110 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(n9830), .B2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n16931) );
  AOI22_X1 U20111 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(
        n9819), .B2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n16930) );
  AOI22_X1 U20112 ( .A1(n9809), .A2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n16929) );
  NAND4_X1 U20113 ( .A1(n16932), .A2(n16931), .A3(n16930), .A4(n16929), .ZN(
        n16933) );
  NOR2_X1 U20114 ( .A1(n16934), .A2(n16933), .ZN(n17174) );
  OAI21_X1 U20115 ( .B1(P3_EBX_REG_19__SCAN_IN), .B2(n16949), .A(n16935), .ZN(
        n16936) );
  AOI22_X1 U20116 ( .A1(n17101), .A2(n17174), .B1(n16936), .B2(n17109), .ZN(
        P3_U2684) );
  OAI21_X1 U20117 ( .B1(P3_EBX_REG_18__SCAN_IN), .B2(n16937), .A(n17109), .ZN(
        n16948) );
  AOI22_X1 U20118 ( .A1(n9811), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(n9832), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n16941) );
  AOI22_X1 U20119 ( .A1(n9829), .A2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n16940) );
  AOI22_X1 U20120 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n11827), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n16939) );
  AOI22_X1 U20121 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n16938) );
  NAND4_X1 U20122 ( .A1(n16941), .A2(n16940), .A3(n16939), .A4(n16938), .ZN(
        n16947) );
  AOI22_X1 U20123 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n17069), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n16945) );
  AOI22_X1 U20124 ( .A1(n11857), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(
        n17024), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n16944) );
  AOI22_X1 U20125 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n16943) );
  AOI22_X1 U20126 ( .A1(n9845), .A2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .B1(
        n9815), .B2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n16942) );
  NAND4_X1 U20127 ( .A1(n16945), .A2(n16944), .A3(n16943), .A4(n16942), .ZN(
        n16946) );
  NOR2_X1 U20128 ( .A1(n16947), .A2(n16946), .ZN(n17178) );
  OAI22_X1 U20129 ( .A1(n16949), .A2(n16948), .B1(n17178), .B2(n17109), .ZN(
        P3_U2685) );
  AOI22_X1 U20130 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(n9810), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n16953) );
  AOI22_X1 U20131 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_11__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n9846), .ZN(n16952) );
  AOI22_X1 U20132 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_2__1__SCAN_IN), .B2(n9811), .ZN(n16951) );
  AOI22_X1 U20133 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n9822), .B1(
        P3_INSTQUEUE_REG_1__1__SCAN_IN), .B2(n17034), .ZN(n16950) );
  NAND4_X1 U20134 ( .A1(n16953), .A2(n16952), .A3(n16951), .A4(n16950), .ZN(
        n16959) );
  AOI22_X1 U20135 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n17049), .B1(
        n9819), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n16957) );
  AOI22_X1 U20136 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n9815), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n15609), .ZN(n16956) );
  AOI22_X1 U20137 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n16955) );
  AOI22_X1 U20138 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_5__1__SCAN_IN), .B1(
        n17024), .B2(P3_INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n16954) );
  NAND4_X1 U20139 ( .A1(n16957), .A2(n16956), .A3(n16955), .A4(n16954), .ZN(
        n16958) );
  NOR2_X1 U20140 ( .A1(n16959), .A2(n16958), .ZN(n17184) );
  OAI21_X1 U20141 ( .B1(P3_EBX_REG_17__SCAN_IN), .B2(n16961), .A(n16960), .ZN(
        n16962) );
  AOI22_X1 U20142 ( .A1(n17101), .A2(n17184), .B1(n16962), .B2(n17109), .ZN(
        P3_U2686) );
  AOI22_X1 U20143 ( .A1(n11857), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(
        n9822), .B2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n16966) );
  AOI22_X1 U20144 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n16965) );
  AOI22_X1 U20145 ( .A1(n9812), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n9815), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n16964) );
  AOI22_X1 U20146 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n16963) );
  NAND4_X1 U20147 ( .A1(n16966), .A2(n16965), .A3(n16964), .A4(n16963), .ZN(
        n16972) );
  AOI22_X1 U20148 ( .A1(n17024), .A2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n16970) );
  AOI22_X1 U20149 ( .A1(n11827), .A2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .B1(
        n9846), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n16969) );
  AOI22_X1 U20150 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n16968) );
  AOI22_X1 U20151 ( .A1(n9838), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n16967) );
  NAND4_X1 U20152 ( .A1(n16970), .A2(n16969), .A3(n16968), .A4(n16967), .ZN(
        n16971) );
  NOR2_X1 U20153 ( .A1(n16972), .A2(n16971), .ZN(n17190) );
  NOR2_X1 U20154 ( .A1(n16974), .A2(n16973), .ZN(n16976) );
  NOR2_X1 U20155 ( .A1(n17101), .A2(n16976), .ZN(n16990) );
  NAND2_X1 U20156 ( .A1(P3_EBX_REG_16__SCAN_IN), .A2(n16990), .ZN(n16978) );
  NAND3_X1 U20157 ( .A1(n18134), .A2(n16976), .A3(n16975), .ZN(n16977) );
  OAI211_X1 U20158 ( .C1(n17190), .C2(n17109), .A(n16978), .B(n16977), .ZN(
        P3_U2687) );
  AOI22_X1 U20159 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_4__7__SCAN_IN), .B1(n9822), .B2(P3_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n16982) );
  AOI22_X1 U20160 ( .A1(n9811), .A2(P3_INSTQUEUE_REG_1__7__SCAN_IN), .B1(n9815), .B2(P3_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n16981) );
  AOI22_X1 U20161 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_8__7__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n16980) );
  AOI22_X1 U20162 ( .A1(n11857), .A2(P3_INSTQUEUE_REG_3__7__SCAN_IN), .B1(
        n9842), .B2(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n16979) );
  NAND4_X1 U20163 ( .A1(n16982), .A2(n16981), .A3(n16980), .A4(n16979), .ZN(
        n16989) );
  AOI22_X1 U20164 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_2__7__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n16987) );
  AOI22_X1 U20165 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_10__7__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n16986) );
  AOI22_X1 U20166 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_9__7__SCAN_IN), .B1(
        n9819), .B2(P3_INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n16985) );
  AOI22_X1 U20167 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_6__7__SCAN_IN), .B1(
        n9846), .B2(P3_INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n16984) );
  NAND4_X1 U20168 ( .A1(n16987), .A2(n16986), .A3(n16985), .A4(n16984), .ZN(
        n16988) );
  NOR2_X1 U20169 ( .A1(n16989), .A2(n16988), .ZN(n17194) );
  AND2_X1 U20170 ( .A1(P3_EBX_REG_14__SCAN_IN), .A2(n17002), .ZN(n17004) );
  OAI21_X1 U20171 ( .B1(P3_EBX_REG_15__SCAN_IN), .B2(n17004), .A(n16990), .ZN(
        n16991) );
  OAI21_X1 U20172 ( .B1(n17194), .B2(n17109), .A(n16991), .ZN(P3_U2688) );
  AOI22_X1 U20173 ( .A1(n9845), .A2(P3_INSTQUEUE_REG_11__6__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n16995) );
  AOI22_X1 U20174 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_9__6__SCAN_IN), .B1(
        n17024), .B2(P3_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n16994) );
  AOI22_X1 U20175 ( .A1(n11857), .A2(P3_INSTQUEUE_REG_3__6__SCAN_IN), .B1(
        n9815), .B2(P3_INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n16993) );
  AOI22_X1 U20176 ( .A1(n15609), .A2(P3_INSTQUEUE_REG_15__6__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n16992) );
  NAND4_X1 U20177 ( .A1(n16995), .A2(n16994), .A3(n16993), .A4(n16992), .ZN(
        n17001) );
  AOI22_X1 U20178 ( .A1(n17069), .A2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n16999) );
  AOI22_X1 U20179 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_13__6__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n16998) );
  AOI22_X1 U20180 ( .A1(n9841), .A2(P3_INSTQUEUE_REG_7__6__SCAN_IN), .B1(n9811), .B2(P3_INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n16997) );
  AOI22_X1 U20181 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_8__6__SCAN_IN), .B1(n9812), .B2(P3_INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n16996) );
  NAND4_X1 U20182 ( .A1(n16999), .A2(n16998), .A3(n16997), .A4(n16996), .ZN(
        n17000) );
  NOR2_X1 U20183 ( .A1(n17001), .A2(n17000), .ZN(n17200) );
  OAI21_X1 U20184 ( .B1(P3_EBX_REG_14__SCAN_IN), .B2(n17002), .A(n17109), .ZN(
        n17003) );
  OAI22_X1 U20185 ( .A1(n17200), .A2(n17109), .B1(n17004), .B2(n17003), .ZN(
        P3_U2689) );
  NAND2_X1 U20186 ( .A1(n18134), .A2(n17033), .ZN(n17018) );
  AOI22_X1 U20187 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_8__4__SCAN_IN), .B1(n9830), .B2(P3_INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n17015) );
  AOI22_X1 U20188 ( .A1(n9810), .A2(P3_INSTQUEUE_REG_3__4__SCAN_IN), .B1(n9841), .B2(P3_INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n17014) );
  AOI22_X1 U20189 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_6__4__SCAN_IN), .B1(
        n9846), .B2(P3_INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n17005) );
  OAI21_X1 U20190 ( .B1(n17006), .B2(n20907), .A(n17005), .ZN(n17012) );
  AOI22_X1 U20191 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_9__4__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n17010) );
  AOI22_X1 U20192 ( .A1(n17024), .A2(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B1(
        n9815), .B2(P3_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n17009) );
  AOI22_X1 U20193 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_13__4__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n17008) );
  AOI22_X1 U20194 ( .A1(n9811), .A2(P3_INSTQUEUE_REG_1__4__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n17007) );
  NAND4_X1 U20195 ( .A1(n17010), .A2(n17009), .A3(n17008), .A4(n17007), .ZN(
        n17011) );
  AOI211_X1 U20196 ( .C1(n9813), .C2(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A(
        n17012), .B(n17011), .ZN(n17013) );
  NAND3_X1 U20197 ( .A1(n17015), .A2(n17014), .A3(n17013), .ZN(n17205) );
  INV_X1 U20198 ( .A(n17205), .ZN(n17017) );
  NAND3_X1 U20199 ( .A1(n17018), .A2(P3_EBX_REG_12__SCAN_IN), .A3(n17109), 
        .ZN(n17016) );
  OAI221_X1 U20200 ( .B1(n17018), .B2(P3_EBX_REG_12__SCAN_IN), .C1(n17109), 
        .C2(n17017), .A(n17016), .ZN(P3_U2691) );
  AOI22_X1 U20201 ( .A1(n11806), .A2(P3_INSTQUEUE_REG_10__3__SCAN_IN), .B1(
        n17069), .B2(P3_INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n17023) );
  AOI22_X1 U20202 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_9__3__SCAN_IN), .B1(
        n9832), .B2(P3_INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n17022) );
  AOI22_X1 U20203 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_13__3__SCAN_IN), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n17021) );
  AOI22_X1 U20204 ( .A1(n9816), .A2(P3_INSTQUEUE_REG_5__3__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n17020) );
  NAND4_X1 U20205 ( .A1(n17023), .A2(n17022), .A3(n17021), .A4(n17020), .ZN(
        n17030) );
  AOI22_X1 U20206 ( .A1(n17024), .A2(P3_INSTQUEUE_REG_14__3__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n17028) );
  AOI22_X1 U20207 ( .A1(n9811), .A2(P3_INSTQUEUE_REG_1__3__SCAN_IN), .B1(n9845), .B2(P3_INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n17027) );
  AOI22_X1 U20208 ( .A1(n9809), .A2(P3_INSTQUEUE_REG_3__3__SCAN_IN), .B1(n9822), .B2(P3_INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n17026) );
  AOI22_X1 U20209 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n17025) );
  NAND4_X1 U20210 ( .A1(n17028), .A2(n17027), .A3(n17026), .A4(n17025), .ZN(
        n17029) );
  NOR2_X1 U20211 ( .A1(n17030), .A2(n17029), .ZN(n17211) );
  INV_X1 U20212 ( .A(n17046), .ZN(n17031) );
  OAI21_X1 U20213 ( .B1(P3_EBX_REG_11__SCAN_IN), .B2(n17031), .A(n17109), .ZN(
        n17032) );
  OAI22_X1 U20214 ( .A1(n17211), .A2(n17109), .B1(n17033), .B2(n17032), .ZN(
        P3_U2692) );
  AOI22_X1 U20215 ( .A1(n9841), .A2(P3_INSTQUEUE_REG_7__2__SCAN_IN), .B1(n9811), .B2(P3_INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n17039) );
  AOI22_X1 U20216 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_2__2__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n17038) );
  AOI22_X1 U20217 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_10__2__SCAN_IN), .B1(
        n9810), .B2(P3_INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n17037) );
  AOI22_X1 U20218 ( .A1(n17035), .A2(P3_INSTQUEUE_REG_6__2__SCAN_IN), .B1(
        n17034), .B2(P3_INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n17036) );
  NAND4_X1 U20219 ( .A1(n17039), .A2(n17038), .A3(n17037), .A4(n17036), .ZN(
        n17045) );
  AOI22_X1 U20220 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_8__2__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n17043) );
  AOI22_X1 U20221 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_13__2__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n17042) );
  AOI22_X1 U20222 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_9__2__SCAN_IN), .B1(
        n9846), .B2(P3_INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n17041) );
  AOI22_X1 U20223 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_4__2__SCAN_IN), .B1(n9815), .B2(P3_INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n17040) );
  NAND4_X1 U20224 ( .A1(n17043), .A2(n17042), .A3(n17041), .A4(n17040), .ZN(
        n17044) );
  NOR2_X1 U20225 ( .A1(n17045), .A2(n17044), .ZN(n17215) );
  OAI21_X1 U20226 ( .B1(P3_EBX_REG_10__SCAN_IN), .B2(n17062), .A(n17046), .ZN(
        n17047) );
  AOI22_X1 U20227 ( .A1(n17101), .A2(n17215), .B1(n17047), .B2(n17109), .ZN(
        P3_U2693) );
  AOI22_X1 U20228 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n17049), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n17053) );
  AOI22_X1 U20229 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n9811), .B1(
        P3_INSTQUEUE_REG_15__1__SCAN_IN), .B2(n15609), .ZN(n17052) );
  AOI22_X1 U20230 ( .A1(n16983), .A2(P3_INSTQUEUE_REG_2__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_0__1__SCAN_IN), .B2(n9842), .ZN(n17051) );
  AOI22_X1 U20231 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n9846), .B1(
        n9830), .B2(P3_INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n17050) );
  NAND4_X1 U20232 ( .A1(n17053), .A2(n17052), .A3(n17051), .A4(n17050), .ZN(
        n17059) );
  AOI22_X1 U20233 ( .A1(n9819), .A2(P3_INSTQUEUE_REG_13__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_5__1__SCAN_IN), .B2(n9816), .ZN(n17057) );
  AOI22_X1 U20234 ( .A1(n17019), .A2(P3_INSTQUEUE_REG_9__1__SCAN_IN), .B1(
        n9812), .B2(P3_INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n17056) );
  AOI22_X1 U20235 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_8__1__SCAN_IN), .B1(
        P3_INSTQUEUE_REG_12__1__SCAN_IN), .B2(n15640), .ZN(n17055) );
  AOI22_X1 U20236 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n9822), .B1(n9809), .B2(P3_INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n17054) );
  NAND4_X1 U20237 ( .A1(n17057), .A2(n17056), .A3(n17055), .A4(n17054), .ZN(
        n17058) );
  NOR2_X1 U20238 ( .A1(n17059), .A2(n17058), .ZN(n17218) );
  INV_X1 U20239 ( .A(n17060), .ZN(n17079) );
  OAI21_X1 U20240 ( .B1(P3_EBX_REG_9__SCAN_IN), .B2(n17079), .A(n17109), .ZN(
        n17061) );
  OAI22_X1 U20241 ( .A1(n17218), .A2(n17109), .B1(n17062), .B2(n17061), .ZN(
        P3_U2694) );
  AOI22_X1 U20242 ( .A1(n9815), .A2(P3_INSTQUEUE_REG_5__0__SCAN_IN), .B1(
        n15640), .B2(P3_INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n17067) );
  AOI22_X1 U20243 ( .A1(n9818), .A2(P3_INSTQUEUE_REG_8__0__SCAN_IN), .B1(
        n17035), .B2(P3_INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n17066) );
  AOI22_X1 U20244 ( .A1(n9846), .A2(P3_INSTQUEUE_REG_11__0__SCAN_IN), .B1(
        n15609), .B2(P3_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n17065) );
  AOI22_X1 U20245 ( .A1(n17063), .A2(P3_INSTQUEUE_REG_9__0__SCAN_IN), .B1(
        n9842), .B2(P3_INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n17064) );
  NAND4_X1 U20246 ( .A1(n17067), .A2(n17066), .A3(n17065), .A4(n17064), .ZN(
        n17075) );
  AOI22_X1 U20247 ( .A1(n9830), .A2(P3_INSTQUEUE_REG_4__0__SCAN_IN), .B1(n9841), .B2(P3_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n17073) );
  AOI22_X1 U20248 ( .A1(n11827), .A2(P3_INSTQUEUE_REG_13__0__SCAN_IN), .B1(
        n9811), .B2(P3_INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n17072) );
  AOI22_X1 U20249 ( .A1(n9809), .A2(P3_INSTQUEUE_REG_3__0__SCAN_IN), .B1(
        n17048), .B2(P3_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n17071) );
  AOI22_X1 U20250 ( .A1(n9813), .A2(P3_INSTQUEUE_REG_10__0__SCAN_IN), .B1(
        n17069), .B2(P3_INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n17070) );
  NAND4_X1 U20251 ( .A1(n17073), .A2(n17072), .A3(n17071), .A4(n17070), .ZN(
        n17074) );
  NOR2_X1 U20252 ( .A1(n17075), .A2(n17074), .ZN(n17225) );
  NOR2_X1 U20253 ( .A1(n17153), .A2(n17107), .ZN(n17106) );
  INV_X1 U20254 ( .A(n17106), .ZN(n17076) );
  NOR2_X1 U20255 ( .A1(n17086), .A2(n17076), .ZN(n17093) );
  AND2_X1 U20256 ( .A1(n17077), .A2(n17093), .ZN(n17081) );
  AOI22_X1 U20257 ( .A1(P3_EBX_REG_8__SCAN_IN), .A2(n17109), .B1(
        P3_EBX_REG_7__SCAN_IN), .B2(n17081), .ZN(n17078) );
  OAI22_X1 U20258 ( .A1(n17225), .A2(n17109), .B1(n17079), .B2(n17078), .ZN(
        P3_U2695) );
  NAND2_X1 U20259 ( .A1(n17109), .A2(P3_EBX_REG_7__SCAN_IN), .ZN(n17083) );
  AOI22_X1 U20260 ( .A1(P3_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n17101), .B1(
        n17081), .B2(n17080), .ZN(n17082) );
  OAI21_X1 U20261 ( .B1(n17084), .B2(n17083), .A(n17082), .ZN(P3_U2696) );
  NAND2_X1 U20262 ( .A1(P3_EBX_REG_5__SCAN_IN), .A2(n17093), .ZN(n17087) );
  INV_X1 U20263 ( .A(P3_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n18131) );
  NAND3_X1 U20264 ( .A1(n17087), .A2(P3_EBX_REG_6__SCAN_IN), .A3(n17109), .ZN(
        n17085) );
  OAI221_X1 U20265 ( .B1(n17087), .B2(P3_EBX_REG_6__SCAN_IN), .C1(n17109), 
        .C2(n18131), .A(n17085), .ZN(P3_U2697) );
  INV_X1 U20266 ( .A(P3_INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n18126) );
  NOR2_X1 U20267 ( .A1(n17107), .A2(n17086), .ZN(n17088) );
  OAI211_X1 U20268 ( .C1(P3_EBX_REG_5__SCAN_IN), .C2(n17088), .A(n17087), .B(
        n17109), .ZN(n17089) );
  OAI21_X1 U20269 ( .B1(n17109), .B2(n18126), .A(n17089), .ZN(P3_U2698) );
  NAND2_X1 U20270 ( .A1(n17090), .A2(n17106), .ZN(n17094) );
  NOR2_X1 U20271 ( .A1(n17091), .A2(n17094), .ZN(n17096) );
  AOI21_X1 U20272 ( .B1(P3_EBX_REG_4__SCAN_IN), .B2(n17109), .A(n17096), .ZN(
        n17092) );
  INV_X1 U20273 ( .A(P3_INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n18121) );
  OAI22_X1 U20274 ( .A1(n17093), .A2(n17092), .B1(n18121), .B2(n17109), .ZN(
        P3_U2699) );
  INV_X1 U20275 ( .A(n17094), .ZN(n17098) );
  AOI21_X1 U20276 ( .B1(P3_EBX_REG_3__SCAN_IN), .B2(n17109), .A(n17098), .ZN(
        n17095) );
  INV_X1 U20277 ( .A(P3_INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n18115) );
  OAI22_X1 U20278 ( .A1(n17096), .A2(n17095), .B1(n18115), .B2(n17109), .ZN(
        P3_U2700) );
  INV_X1 U20279 ( .A(n17107), .ZN(n17104) );
  AOI21_X1 U20280 ( .B1(n17104), .B2(n17097), .A(P3_EBX_REG_2__SCAN_IN), .ZN(
        n17099) );
  AOI221_X1 U20281 ( .B1(n17099), .B2(n17109), .C1(n18110), .C2(n17101), .A(
        n17098), .ZN(P3_U2701) );
  AOI22_X1 U20282 ( .A1(P3_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n17101), .B1(
        n17100), .B2(n17106), .ZN(n17102) );
  OAI21_X1 U20283 ( .B1(n17104), .B2(n17103), .A(n17102), .ZN(P3_U2702) );
  AOI22_X1 U20284 ( .A1(P3_EBX_REG_0__SCAN_IN), .A2(n17107), .B1(n17106), .B2(
        n17105), .ZN(n17108) );
  OAI21_X1 U20285 ( .B1(n18098), .B2(n17109), .A(n17108), .ZN(P3_U2703) );
  INV_X1 U20286 ( .A(P3_EAX_REG_29__SCAN_IN), .ZN(n17332) );
  INV_X1 U20287 ( .A(P3_EAX_REG_26__SCAN_IN), .ZN(n17266) );
  INV_X1 U20288 ( .A(P3_EAX_REG_22__SCAN_IN), .ZN(n17273) );
  INV_X1 U20289 ( .A(P3_EAX_REG_17__SCAN_IN), .ZN(n17316) );
  INV_X1 U20290 ( .A(P3_EAX_REG_15__SCAN_IN), .ZN(n17365) );
  INV_X1 U20291 ( .A(P3_EAX_REG_8__SCAN_IN), .ZN(n17296) );
  INV_X1 U20292 ( .A(P3_EAX_REG_1__SCAN_IN), .ZN(n17337) );
  INV_X1 U20293 ( .A(P3_EAX_REG_7__SCAN_IN), .ZN(n17344) );
  INV_X1 U20294 ( .A(P3_EAX_REG_2__SCAN_IN), .ZN(n17305) );
  NAND4_X1 U20295 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(P3_EAX_REG_6__SCAN_IN), 
        .A3(P3_EAX_REG_4__SCAN_IN), .A4(P3_EAX_REG_3__SCAN_IN), .ZN(n17226) );
  NOR3_X1 U20296 ( .A1(n17344), .A2(n17305), .A3(n17226), .ZN(n17228) );
  INV_X1 U20297 ( .A(P3_EAX_REG_13__SCAN_IN), .ZN(n17358) );
  NAND4_X1 U20298 ( .A1(P3_EAX_REG_11__SCAN_IN), .A2(P3_EAX_REG_10__SCAN_IN), 
        .A3(P3_EAX_REG_9__SCAN_IN), .A4(P3_EAX_REG_12__SCAN_IN), .ZN(n17110)
         );
  NOR2_X1 U20299 ( .A1(n17358), .A2(n17110), .ZN(n17196) );
  NAND4_X1 U20300 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(P3_EAX_REG_20__SCAN_IN), 
        .A3(P3_EAX_REG_19__SCAN_IN), .A4(P3_EAX_REG_18__SCAN_IN), .ZN(n17160)
         );
  NAND2_X1 U20301 ( .A1(n17120), .A2(P3_EAX_REG_30__SCAN_IN), .ZN(n17113) );
  NAND2_X1 U20302 ( .A1(n17112), .A2(n17252), .ZN(n17161) );
  INV_X1 U20303 ( .A(P3_EAX_REG_30__SCAN_IN), .ZN(n17334) );
  AOI22_X1 U20304 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n17185), .B1(n17245), .B2(
        n17114), .ZN(n17117) );
  NOR2_X2 U20305 ( .A1(n17115), .A2(n17247), .ZN(n17186) );
  AOI22_X1 U20306 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17186), .B1(n17120), .B2(
        n17334), .ZN(n17116) );
  OAI211_X1 U20307 ( .C1(n17118), .C2(n17334), .A(n17117), .B(n17116), .ZN(
        P3_U2705) );
  INV_X1 U20308 ( .A(BUF2_REG_29__SCAN_IN), .ZN(n20974) );
  AOI22_X1 U20309 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17186), .B1(n17245), .B2(
        n17119), .ZN(n17123) );
  AOI211_X1 U20310 ( .C1(n17332), .C2(n17124), .A(n17120), .B(n17252), .ZN(
        n17121) );
  INV_X1 U20311 ( .A(n17121), .ZN(n17122) );
  OAI211_X1 U20312 ( .C1(n17161), .C2(n20974), .A(n17123), .B(n17122), .ZN(
        P3_U2706) );
  AOI22_X1 U20313 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17186), .B1(
        BUF2_REG_28__SCAN_IN), .B2(n17185), .ZN(n17126) );
  OAI211_X1 U20314 ( .C1(n17132), .C2(P3_EAX_REG_28__SCAN_IN), .A(n17247), .B(
        n17124), .ZN(n17125) );
  OAI211_X1 U20315 ( .C1(n17127), .C2(n17257), .A(n17126), .B(n17125), .ZN(
        P3_U2707) );
  AOI21_X1 U20316 ( .B1(P3_EAX_REG_27__SCAN_IN), .B2(n17247), .A(n17133), .ZN(
        n17131) );
  AOI22_X1 U20317 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n17185), .B1(n17245), .B2(
        n17128), .ZN(n17130) );
  NAND2_X1 U20318 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17186), .ZN(n17129) );
  OAI211_X1 U20319 ( .C1(n17132), .C2(n17131), .A(n17130), .B(n17129), .ZN(
        P3_U2708) );
  AOI22_X1 U20320 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17186), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n17185), .ZN(n17136) );
  AOI211_X1 U20321 ( .C1(n17266), .C2(n17139), .A(n17133), .B(n17252), .ZN(
        n17134) );
  INV_X1 U20322 ( .A(n17134), .ZN(n17135) );
  OAI211_X1 U20323 ( .C1(n17137), .C2(n17257), .A(n17136), .B(n17135), .ZN(
        P3_U2709) );
  INV_X1 U20324 ( .A(BUF2_REG_25__SCAN_IN), .ZN(n18101) );
  AOI22_X1 U20325 ( .A1(BUF2_REG_9__SCAN_IN), .A2(n17186), .B1(n17245), .B2(
        n17138), .ZN(n17142) );
  OAI211_X1 U20326 ( .C1(n17140), .C2(P3_EAX_REG_25__SCAN_IN), .A(n17247), .B(
        n17139), .ZN(n17141) );
  OAI211_X1 U20327 ( .C1(n17161), .C2(n18101), .A(n17142), .B(n17141), .ZN(
        P3_U2710) );
  AOI22_X1 U20328 ( .A1(BUF2_REG_8__SCAN_IN), .A2(n17186), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n17185), .ZN(n17146) );
  OAI211_X1 U20329 ( .C1(n17144), .C2(P3_EAX_REG_24__SCAN_IN), .A(n17247), .B(
        n17143), .ZN(n17145) );
  OAI211_X1 U20330 ( .C1(n17147), .C2(n17257), .A(n17146), .B(n17145), .ZN(
        P3_U2711) );
  AOI22_X1 U20331 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17186), .B1(n17245), .B2(
        n17148), .ZN(n17152) );
  OAI211_X1 U20332 ( .C1(P3_EAX_REG_23__SCAN_IN), .C2(n17150), .A(n17247), .B(
        n17149), .ZN(n17151) );
  OAI211_X1 U20333 ( .C1(n17161), .C2(n15069), .A(n17152), .B(n17151), .ZN(
        P3_U2712) );
  NAND2_X1 U20334 ( .A1(n17179), .A2(n17273), .ZN(n17159) );
  AOI22_X1 U20335 ( .A1(BUF2_REG_22__SCAN_IN), .A2(n17185), .B1(n17245), .B2(
        n17154), .ZN(n17158) );
  INV_X1 U20336 ( .A(P3_EAX_REG_19__SCAN_IN), .ZN(n17280) );
  NAND2_X1 U20337 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17179), .ZN(n17175) );
  NAND2_X1 U20338 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17170), .ZN(n17166) );
  NAND2_X1 U20339 ( .A1(n17247), .A2(n17166), .ZN(n17165) );
  OAI21_X1 U20340 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17155), .A(n17165), .ZN(
        n17156) );
  AOI22_X1 U20341 ( .A1(BUF2_REG_6__SCAN_IN), .A2(n17186), .B1(
        P3_EAX_REG_22__SCAN_IN), .B2(n17156), .ZN(n17157) );
  OAI211_X1 U20342 ( .C1(n17160), .C2(n17159), .A(n17158), .B(n17157), .ZN(
        P3_U2713) );
  INV_X1 U20343 ( .A(P3_EAX_REG_21__SCAN_IN), .ZN(n17275) );
  OAI22_X1 U20344 ( .A1(n17162), .A2(n17257), .B1(n15075), .B2(n17161), .ZN(
        n17163) );
  AOI21_X1 U20345 ( .B1(BUF2_REG_5__SCAN_IN), .B2(n17186), .A(n17163), .ZN(
        n17164) );
  OAI221_X1 U20346 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(n17166), .C1(n17275), 
        .C2(n17165), .A(n17164), .ZN(P3_U2714) );
  AOI22_X1 U20347 ( .A1(BUF2_REG_4__SCAN_IN), .A2(n17186), .B1(
        BUF2_REG_20__SCAN_IN), .B2(n17185), .ZN(n17168) );
  OAI211_X1 U20348 ( .C1(n17170), .C2(P3_EAX_REG_20__SCAN_IN), .A(n17247), .B(
        n17166), .ZN(n17167) );
  OAI211_X1 U20349 ( .C1(n17169), .C2(n17257), .A(n17168), .B(n17167), .ZN(
        P3_U2715) );
  AOI22_X1 U20350 ( .A1(BUF2_REG_3__SCAN_IN), .A2(n17186), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n17185), .ZN(n17173) );
  AOI211_X1 U20351 ( .C1(n17280), .C2(n17175), .A(n17170), .B(n17252), .ZN(
        n17171) );
  INV_X1 U20352 ( .A(n17171), .ZN(n17172) );
  OAI211_X1 U20353 ( .C1(n17174), .C2(n17257), .A(n17173), .B(n17172), .ZN(
        P3_U2716) );
  AOI22_X1 U20354 ( .A1(BUF2_REG_2__SCAN_IN), .A2(n17186), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n17185), .ZN(n17177) );
  OAI211_X1 U20355 ( .C1(n17179), .C2(P3_EAX_REG_18__SCAN_IN), .A(n17247), .B(
        n17175), .ZN(n17176) );
  OAI211_X1 U20356 ( .C1(n17178), .C2(n17257), .A(n17177), .B(n17176), .ZN(
        P3_U2717) );
  AOI22_X1 U20357 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17186), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n17185), .ZN(n17183) );
  INV_X1 U20358 ( .A(n17187), .ZN(n17181) );
  INV_X1 U20359 ( .A(n17179), .ZN(n17180) );
  OAI211_X1 U20360 ( .C1(n17181), .C2(P3_EAX_REG_17__SCAN_IN), .A(n17247), .B(
        n17180), .ZN(n17182) );
  OAI211_X1 U20361 ( .C1(n17184), .C2(n17257), .A(n17183), .B(n17182), .ZN(
        P3_U2718) );
  AOI22_X1 U20362 ( .A1(BUF2_REG_0__SCAN_IN), .A2(n17186), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n17185), .ZN(n17189) );
  OAI211_X1 U20363 ( .C1(P3_EAX_REG_16__SCAN_IN), .C2(n17191), .A(n17247), .B(
        n17187), .ZN(n17188) );
  OAI211_X1 U20364 ( .C1(n17190), .C2(n17257), .A(n17189), .B(n17188), .ZN(
        P3_U2719) );
  AOI211_X1 U20365 ( .C1(n17365), .C2(n17197), .A(n17252), .B(n17191), .ZN(
        n17192) );
  AOI21_X1 U20366 ( .B1(n17255), .B2(BUF2_REG_15__SCAN_IN), .A(n17192), .ZN(
        n17193) );
  OAI21_X1 U20367 ( .B1(n17194), .B2(n17257), .A(n17193), .ZN(P3_U2720) );
  NAND2_X1 U20368 ( .A1(n18134), .A2(n17221), .ZN(n17216) );
  NOR2_X1 U20369 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17216), .ZN(n17195) );
  AOI22_X1 U20370 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17255), .B1(n17196), .B2(
        n17195), .ZN(n17199) );
  NAND3_X1 U20371 ( .A1(P3_EAX_REG_14__SCAN_IN), .A2(n17247), .A3(n17197), 
        .ZN(n17198) );
  OAI211_X1 U20372 ( .C1(n17200), .C2(n17257), .A(n17199), .B(n17198), .ZN(
        P3_U2721) );
  INV_X1 U20373 ( .A(P3_EAX_REG_11__SCAN_IN), .ZN(n17355) );
  INV_X1 U20374 ( .A(P3_EAX_REG_9__SCAN_IN), .ZN(n20947) );
  NOR2_X1 U20375 ( .A1(n20947), .A2(n17216), .ZN(n17220) );
  NAND2_X1 U20376 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17220), .ZN(n17212) );
  NOR2_X1 U20377 ( .A1(n17355), .A2(n17212), .ZN(n17204) );
  NAND2_X1 U20378 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(n17204), .ZN(n17203) );
  NAND2_X1 U20379 ( .A1(n17247), .A2(n17203), .ZN(n17207) );
  AOI22_X1 U20380 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17255), .B1(n17245), .B2(
        n17201), .ZN(n17202) );
  OAI221_X1 U20381 ( .B1(P3_EAX_REG_13__SCAN_IN), .B2(n17203), .C1(n17358), 
        .C2(n17207), .A(n17202), .ZN(P3_U2722) );
  INV_X1 U20382 ( .A(n17204), .ZN(n17209) );
  INV_X1 U20383 ( .A(P3_EAX_REG_12__SCAN_IN), .ZN(n21063) );
  AOI22_X1 U20384 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17255), .B1(n17245), .B2(
        n17205), .ZN(n17206) );
  OAI221_X1 U20385 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(n17209), .C1(n21063), 
        .C2(n17207), .A(n17206), .ZN(P3_U2723) );
  OAI21_X1 U20386 ( .B1(n17252), .B2(n17355), .A(n17212), .ZN(n17208) );
  AOI22_X1 U20387 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17255), .B1(n17209), .B2(
        n17208), .ZN(n17210) );
  OAI21_X1 U20388 ( .B1(n17211), .B2(n17257), .A(n17210), .ZN(P3_U2724) );
  NAND2_X1 U20389 ( .A1(BUF2_REG_10__SCAN_IN), .A2(n17255), .ZN(n17214) );
  OAI211_X1 U20390 ( .C1(P3_EAX_REG_10__SCAN_IN), .C2(n17220), .A(n17247), .B(
        n17212), .ZN(n17213) );
  OAI211_X1 U20391 ( .C1(n17215), .C2(n17257), .A(n17214), .B(n17213), .ZN(
        P3_U2725) );
  INV_X1 U20392 ( .A(BUF2_REG_9__SCAN_IN), .ZN(n17348) );
  OAI21_X1 U20393 ( .B1(n20947), .B2(n17252), .A(n17216), .ZN(n17217) );
  INV_X1 U20394 ( .A(n17217), .ZN(n17219) );
  OAI222_X1 U20395 ( .A1(n17243), .A2(n17348), .B1(n17220), .B2(n17219), .C1(
        n17257), .C2(n17218), .ZN(P3_U2726) );
  AOI211_X1 U20396 ( .C1(n17296), .C2(n17222), .A(n17252), .B(n17221), .ZN(
        n17223) );
  AOI21_X1 U20397 ( .B1(n17255), .B2(BUF2_REG_8__SCAN_IN), .A(n17223), .ZN(
        n17224) );
  OAI21_X1 U20398 ( .B1(n17225), .B2(n17257), .A(n17224), .ZN(P3_U2727) );
  NAND3_X1 U20399 ( .A1(n18134), .A2(n17251), .A3(P3_EAX_REG_2__SCAN_IN), .ZN(
        n17246) );
  NOR2_X1 U20400 ( .A1(n17226), .A2(n17246), .ZN(n17230) );
  AOI21_X1 U20401 ( .B1(P3_EAX_REG_7__SCAN_IN), .B2(n17247), .A(n17230), .ZN(
        n17229) );
  AOI22_X1 U20402 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17255), .B1(n17245), .B2(
        n11904), .ZN(n17227) );
  OAI221_X1 U20403 ( .B1(n17229), .B2(n17228), .C1(n17229), .C2(n17251), .A(
        n17227), .ZN(P3_U2728) );
  INV_X1 U20404 ( .A(P3_EAX_REG_5__SCAN_IN), .ZN(n21002) );
  INV_X1 U20405 ( .A(P3_EAX_REG_3__SCAN_IN), .ZN(n17303) );
  NOR2_X1 U20406 ( .A1(n17303), .A2(n17246), .ZN(n17242) );
  NAND2_X1 U20407 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17242), .ZN(n17232) );
  NOR2_X1 U20408 ( .A1(n21002), .A2(n17232), .ZN(n17234) );
  AOI21_X1 U20409 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(n17247), .A(n17234), .ZN(
        n17231) );
  OAI222_X1 U20410 ( .A1(n17243), .A2(n18127), .B1(n17231), .B2(n17230), .C1(
        n17257), .C2(n17681), .ZN(P3_U2729) );
  INV_X1 U20411 ( .A(BUF2_REG_5__SCAN_IN), .ZN(n18122) );
  INV_X1 U20412 ( .A(n17232), .ZN(n17238) );
  AOI21_X1 U20413 ( .B1(P3_EAX_REG_5__SCAN_IN), .B2(n17247), .A(n17238), .ZN(
        n17235) );
  OAI222_X1 U20414 ( .A1(n17243), .A2(n18122), .B1(n17235), .B2(n17234), .C1(
        n17257), .C2(n17233), .ZN(P3_U2730) );
  INV_X1 U20415 ( .A(BUF2_REG_4__SCAN_IN), .ZN(n18116) );
  AOI21_X1 U20416 ( .B1(P3_EAX_REG_4__SCAN_IN), .B2(n17247), .A(n17242), .ZN(
        n17237) );
  OAI222_X1 U20417 ( .A1(n18116), .A2(n17243), .B1(n17238), .B2(n17237), .C1(
        n17257), .C2(n17236), .ZN(P3_U2731) );
  INV_X1 U20418 ( .A(BUF2_REG_3__SCAN_IN), .ZN(n18111) );
  INV_X1 U20419 ( .A(n17246), .ZN(n17239) );
  AOI21_X1 U20420 ( .B1(P3_EAX_REG_3__SCAN_IN), .B2(n17247), .A(n17239), .ZN(
        n17241) );
  OAI222_X1 U20421 ( .A1(n18111), .A2(n17243), .B1(n17242), .B2(n17241), .C1(
        n17257), .C2(n17240), .ZN(P3_U2732) );
  AOI22_X1 U20422 ( .A1(n17255), .A2(BUF2_REG_2__SCAN_IN), .B1(n17245), .B2(
        n17244), .ZN(n17249) );
  OAI211_X1 U20423 ( .C1(n17251), .C2(P3_EAX_REG_2__SCAN_IN), .A(n17247), .B(
        n17246), .ZN(n17248) );
  NAND2_X1 U20424 ( .A1(n17249), .A2(n17248), .ZN(P3_U2733) );
  INV_X1 U20425 ( .A(n17250), .ZN(n17258) );
  AOI211_X1 U20426 ( .C1(n17337), .C2(n17253), .A(n17252), .B(n17251), .ZN(
        n17254) );
  AOI21_X1 U20427 ( .B1(n17255), .B2(BUF2_REG_1__SCAN_IN), .A(n17254), .ZN(
        n17256) );
  OAI21_X1 U20428 ( .B1(n17258), .B2(n17257), .A(n17256), .ZN(P3_U2734) );
  NOR2_X2 U20429 ( .A1(n18706), .A2(n17533), .ZN(n18743) );
  INV_X1 U20430 ( .A(n17313), .ZN(n17311) );
  NOR2_X4 U20431 ( .A1(n18743), .A2(n17260), .ZN(n17278) );
  AND2_X1 U20432 ( .A1(n17278), .A2(P3_DATAO_REG_31__SCAN_IN), .ZN(P3_U2736)
         );
  NAND2_X1 U20433 ( .A1(n17260), .A2(n18746), .ZN(n17285) );
  AOI22_X1 U20434 ( .A1(n18743), .A2(P3_UWORD_REG_14__SCAN_IN), .B1(
        P3_DATAO_REG_30__SCAN_IN), .B2(n17278), .ZN(n17261) );
  OAI21_X1 U20435 ( .B1(n17334), .B2(n17285), .A(n17261), .ZN(P3_U2737) );
  AOI22_X1 U20436 ( .A1(n18743), .A2(P3_UWORD_REG_13__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_29__SCAN_IN), .ZN(n17262) );
  OAI21_X1 U20437 ( .B1(n17332), .B2(n17285), .A(n17262), .ZN(P3_U2738) );
  INV_X1 U20438 ( .A(P3_EAX_REG_28__SCAN_IN), .ZN(n17330) );
  AOI22_X1 U20439 ( .A1(n18743), .A2(P3_UWORD_REG_12__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_28__SCAN_IN), .ZN(n17263) );
  OAI21_X1 U20440 ( .B1(n17330), .B2(n17285), .A(n17263), .ZN(P3_U2739) );
  INV_X1 U20441 ( .A(P3_EAX_REG_27__SCAN_IN), .ZN(n17328) );
  AOI22_X1 U20442 ( .A1(n18743), .A2(P3_UWORD_REG_11__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_27__SCAN_IN), .ZN(n17264) );
  OAI21_X1 U20443 ( .B1(n17328), .B2(n17285), .A(n17264), .ZN(P3_U2740) );
  AOI22_X1 U20444 ( .A1(n18743), .A2(P3_UWORD_REG_10__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_26__SCAN_IN), .ZN(n17265) );
  OAI21_X1 U20445 ( .B1(n17266), .B2(n17285), .A(n17265), .ZN(P3_U2741) );
  INV_X1 U20446 ( .A(P3_EAX_REG_25__SCAN_IN), .ZN(n17268) );
  AOI22_X1 U20447 ( .A1(n18743), .A2(P3_UWORD_REG_9__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_25__SCAN_IN), .ZN(n17267) );
  OAI21_X1 U20448 ( .B1(n17268), .B2(n17285), .A(n17267), .ZN(P3_U2742) );
  INV_X1 U20449 ( .A(P3_EAX_REG_24__SCAN_IN), .ZN(n17270) );
  AOI22_X1 U20450 ( .A1(n18743), .A2(P3_UWORD_REG_8__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_24__SCAN_IN), .ZN(n17269) );
  OAI21_X1 U20451 ( .B1(n17270), .B2(n17285), .A(n17269), .ZN(P3_U2743) );
  INV_X1 U20452 ( .A(P3_EAX_REG_23__SCAN_IN), .ZN(n17323) );
  CLKBUF_X1 U20453 ( .A(n18743), .Z(n17307) );
  AOI22_X1 U20454 ( .A1(n17307), .A2(P3_UWORD_REG_7__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_23__SCAN_IN), .ZN(n17271) );
  OAI21_X1 U20455 ( .B1(n17323), .B2(n17285), .A(n17271), .ZN(P3_U2744) );
  AOI22_X1 U20456 ( .A1(n17307), .A2(P3_UWORD_REG_6__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_22__SCAN_IN), .ZN(n17272) );
  OAI21_X1 U20457 ( .B1(n17273), .B2(n17285), .A(n17272), .ZN(P3_U2745) );
  AOI22_X1 U20458 ( .A1(n17307), .A2(P3_UWORD_REG_5__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_21__SCAN_IN), .ZN(n17274) );
  OAI21_X1 U20459 ( .B1(n17275), .B2(n17285), .A(n17274), .ZN(P3_U2746) );
  INV_X1 U20460 ( .A(P3_EAX_REG_20__SCAN_IN), .ZN(n17277) );
  AOI22_X1 U20461 ( .A1(n17307), .A2(P3_UWORD_REG_4__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_20__SCAN_IN), .ZN(n17276) );
  OAI21_X1 U20462 ( .B1(n17277), .B2(n17285), .A(n17276), .ZN(P3_U2747) );
  AOI22_X1 U20463 ( .A1(n17307), .A2(P3_UWORD_REG_3__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_19__SCAN_IN), .ZN(n17279) );
  OAI21_X1 U20464 ( .B1(n17280), .B2(n17285), .A(n17279), .ZN(P3_U2748) );
  INV_X1 U20465 ( .A(P3_EAX_REG_18__SCAN_IN), .ZN(n17282) );
  AOI22_X1 U20466 ( .A1(n17307), .A2(P3_UWORD_REG_2__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_18__SCAN_IN), .ZN(n17281) );
  OAI21_X1 U20467 ( .B1(n17282), .B2(n17285), .A(n17281), .ZN(P3_U2749) );
  AOI22_X1 U20468 ( .A1(n17307), .A2(P3_UWORD_REG_1__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_17__SCAN_IN), .ZN(n17283) );
  OAI21_X1 U20469 ( .B1(n17316), .B2(n17285), .A(n17283), .ZN(P3_U2750) );
  INV_X1 U20470 ( .A(P3_EAX_REG_16__SCAN_IN), .ZN(n17286) );
  AOI22_X1 U20471 ( .A1(n17307), .A2(P3_UWORD_REG_0__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_16__SCAN_IN), .ZN(n17284) );
  OAI21_X1 U20472 ( .B1(n17286), .B2(n17285), .A(n17284), .ZN(P3_U2751) );
  AOI22_X1 U20473 ( .A1(n17307), .A2(P3_LWORD_REG_15__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_15__SCAN_IN), .ZN(n17287) );
  OAI21_X1 U20474 ( .B1(n17365), .B2(n17309), .A(n17287), .ZN(P3_U2752) );
  INV_X1 U20475 ( .A(P3_EAX_REG_14__SCAN_IN), .ZN(n17360) );
  AOI22_X1 U20476 ( .A1(n17307), .A2(P3_LWORD_REG_14__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_14__SCAN_IN), .ZN(n17288) );
  OAI21_X1 U20477 ( .B1(n17360), .B2(n17309), .A(n17288), .ZN(P3_U2753) );
  AOI22_X1 U20478 ( .A1(n17307), .A2(P3_LWORD_REG_13__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_13__SCAN_IN), .ZN(n17289) );
  OAI21_X1 U20479 ( .B1(n17358), .B2(n17309), .A(n17289), .ZN(P3_U2754) );
  AOI22_X1 U20480 ( .A1(n17307), .A2(P3_LWORD_REG_12__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_12__SCAN_IN), .ZN(n17290) );
  OAI21_X1 U20481 ( .B1(n21063), .B2(n17309), .A(n17290), .ZN(P3_U2755) );
  AOI22_X1 U20482 ( .A1(n17307), .A2(P3_LWORD_REG_11__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_11__SCAN_IN), .ZN(n17291) );
  OAI21_X1 U20483 ( .B1(n17355), .B2(n17309), .A(n17291), .ZN(P3_U2756) );
  INV_X1 U20484 ( .A(P3_EAX_REG_10__SCAN_IN), .ZN(n17293) );
  AOI22_X1 U20485 ( .A1(n17307), .A2(P3_LWORD_REG_10__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_10__SCAN_IN), .ZN(n17292) );
  OAI21_X1 U20486 ( .B1(n17293), .B2(n17309), .A(n17292), .ZN(P3_U2757) );
  AOI22_X1 U20487 ( .A1(n17307), .A2(P3_LWORD_REG_9__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_9__SCAN_IN), .ZN(n17294) );
  OAI21_X1 U20488 ( .B1(n20947), .B2(n17309), .A(n17294), .ZN(P3_U2758) );
  AOI22_X1 U20489 ( .A1(n17307), .A2(P3_LWORD_REG_8__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_8__SCAN_IN), .ZN(n17295) );
  OAI21_X1 U20490 ( .B1(n17296), .B2(n17309), .A(n17295), .ZN(P3_U2759) );
  AOI22_X1 U20491 ( .A1(n17307), .A2(P3_LWORD_REG_7__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_7__SCAN_IN), .ZN(n17297) );
  OAI21_X1 U20492 ( .B1(n17344), .B2(n17309), .A(n17297), .ZN(P3_U2760) );
  INV_X1 U20493 ( .A(P3_EAX_REG_6__SCAN_IN), .ZN(n21047) );
  AOI22_X1 U20494 ( .A1(n17307), .A2(P3_LWORD_REG_6__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_6__SCAN_IN), .ZN(n17298) );
  OAI21_X1 U20495 ( .B1(n21047), .B2(n17309), .A(n17298), .ZN(P3_U2761) );
  AOI22_X1 U20496 ( .A1(n17307), .A2(P3_LWORD_REG_5__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_5__SCAN_IN), .ZN(n17299) );
  OAI21_X1 U20497 ( .B1(n21002), .B2(n17309), .A(n17299), .ZN(P3_U2762) );
  INV_X1 U20498 ( .A(P3_EAX_REG_4__SCAN_IN), .ZN(n17301) );
  AOI22_X1 U20499 ( .A1(n17307), .A2(P3_LWORD_REG_4__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_4__SCAN_IN), .ZN(n17300) );
  OAI21_X1 U20500 ( .B1(n17301), .B2(n17309), .A(n17300), .ZN(P3_U2763) );
  AOI22_X1 U20501 ( .A1(n17307), .A2(P3_LWORD_REG_3__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_3__SCAN_IN), .ZN(n17302) );
  OAI21_X1 U20502 ( .B1(n17303), .B2(n17309), .A(n17302), .ZN(P3_U2764) );
  AOI22_X1 U20503 ( .A1(n17307), .A2(P3_LWORD_REG_2__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n17304) );
  OAI21_X1 U20504 ( .B1(n17305), .B2(n17309), .A(n17304), .ZN(P3_U2765) );
  AOI22_X1 U20505 ( .A1(n17307), .A2(P3_LWORD_REG_1__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_1__SCAN_IN), .ZN(n17306) );
  OAI21_X1 U20506 ( .B1(n17337), .B2(n17309), .A(n17306), .ZN(P3_U2766) );
  AOI22_X1 U20507 ( .A1(n17307), .A2(P3_LWORD_REG_0__SCAN_IN), .B1(n17278), 
        .B2(P3_DATAO_REG_0__SCAN_IN), .ZN(n17308) );
  OAI21_X1 U20508 ( .B1(n17310), .B2(n17309), .A(n17308), .ZN(P3_U2767) );
  INV_X1 U20509 ( .A(BUF2_REG_0__SCAN_IN), .ZN(n18091) );
  OAI211_X1 U20510 ( .C1(n18747), .C2(n18100), .A(n17312), .B(n17311), .ZN(
        n17361) );
  NOR2_X2 U20511 ( .A1(n17349), .A2(n18100), .ZN(n17362) );
  NOR2_X2 U20512 ( .A1(n17313), .A2(n18589), .ZN(n17350) );
  AOI22_X1 U20513 ( .A1(P3_EAX_REG_16__SCAN_IN), .A2(n17350), .B1(
        P3_UWORD_REG_0__SCAN_IN), .B2(n17349), .ZN(n17314) );
  OAI21_X1 U20514 ( .B1(n18091), .B2(n17352), .A(n17314), .ZN(P3_U2768) );
  AOI22_X1 U20515 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17362), .B1(
        P3_UWORD_REG_1__SCAN_IN), .B2(n17349), .ZN(n17315) );
  OAI21_X1 U20516 ( .B1(n17316), .B2(n17364), .A(n17315), .ZN(P3_U2769) );
  INV_X1 U20517 ( .A(BUF2_REG_2__SCAN_IN), .ZN(n18105) );
  AOI22_X1 U20518 ( .A1(P3_EAX_REG_18__SCAN_IN), .A2(n17350), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(n17349), .ZN(n17317) );
  OAI21_X1 U20519 ( .B1(n18105), .B2(n17352), .A(n17317), .ZN(P3_U2770) );
  AOI22_X1 U20520 ( .A1(P3_EAX_REG_19__SCAN_IN), .A2(n17350), .B1(
        P3_UWORD_REG_3__SCAN_IN), .B2(n17349), .ZN(n17318) );
  OAI21_X1 U20521 ( .B1(n18111), .B2(n17352), .A(n17318), .ZN(P3_U2771) );
  AOI22_X1 U20522 ( .A1(P3_EAX_REG_20__SCAN_IN), .A2(n17350), .B1(
        P3_UWORD_REG_4__SCAN_IN), .B2(n17349), .ZN(n17319) );
  OAI21_X1 U20523 ( .B1(n18116), .B2(n17352), .A(n17319), .ZN(P3_U2772) );
  AOI22_X1 U20524 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(n17350), .B1(
        P3_UWORD_REG_5__SCAN_IN), .B2(n17349), .ZN(n17320) );
  OAI21_X1 U20525 ( .B1(n18122), .B2(n17352), .A(n17320), .ZN(P3_U2773) );
  AOI22_X1 U20526 ( .A1(P3_EAX_REG_22__SCAN_IN), .A2(n17350), .B1(
        P3_UWORD_REG_6__SCAN_IN), .B2(n17349), .ZN(n17321) );
  OAI21_X1 U20527 ( .B1(n18127), .B2(n17352), .A(n17321), .ZN(P3_U2774) );
  AOI22_X1 U20528 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17362), .B1(
        P3_UWORD_REG_7__SCAN_IN), .B2(n17349), .ZN(n17322) );
  OAI21_X1 U20529 ( .B1(n17323), .B2(n17364), .A(n17322), .ZN(P3_U2775) );
  INV_X1 U20530 ( .A(BUF2_REG_8__SCAN_IN), .ZN(n17346) );
  AOI22_X1 U20531 ( .A1(P3_EAX_REG_24__SCAN_IN), .A2(n17350), .B1(
        P3_UWORD_REG_8__SCAN_IN), .B2(n17349), .ZN(n17324) );
  OAI21_X1 U20532 ( .B1(n17346), .B2(n17352), .A(n17324), .ZN(P3_U2776) );
  AOI22_X1 U20533 ( .A1(P3_EAX_REG_25__SCAN_IN), .A2(n17350), .B1(
        P3_UWORD_REG_9__SCAN_IN), .B2(n17349), .ZN(n17325) );
  OAI21_X1 U20534 ( .B1(n17348), .B2(n17352), .A(n17325), .ZN(P3_U2777) );
  AOI22_X1 U20535 ( .A1(P3_EAX_REG_26__SCAN_IN), .A2(n17350), .B1(
        P3_UWORD_REG_10__SCAN_IN), .B2(n17349), .ZN(n17326) );
  OAI21_X1 U20536 ( .B1(n17353), .B2(n17352), .A(n17326), .ZN(P3_U2778) );
  AOI22_X1 U20537 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17362), .B1(
        P3_UWORD_REG_11__SCAN_IN), .B2(n17349), .ZN(n17327) );
  OAI21_X1 U20538 ( .B1(n17328), .B2(n17364), .A(n17327), .ZN(P3_U2779) );
  AOI22_X1 U20539 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17362), .B1(
        P3_UWORD_REG_12__SCAN_IN), .B2(n17349), .ZN(n17329) );
  OAI21_X1 U20540 ( .B1(n17330), .B2(n17364), .A(n17329), .ZN(P3_U2780) );
  AOI22_X1 U20541 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17362), .B1(
        P3_UWORD_REG_13__SCAN_IN), .B2(n17349), .ZN(n17331) );
  OAI21_X1 U20542 ( .B1(n17332), .B2(n17364), .A(n17331), .ZN(P3_U2781) );
  AOI22_X1 U20543 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17362), .B1(
        P3_UWORD_REG_14__SCAN_IN), .B2(n17349), .ZN(n17333) );
  OAI21_X1 U20544 ( .B1(n17334), .B2(n17364), .A(n17333), .ZN(P3_U2782) );
  AOI22_X1 U20545 ( .A1(P3_EAX_REG_0__SCAN_IN), .A2(n17350), .B1(
        P3_LWORD_REG_0__SCAN_IN), .B2(n17349), .ZN(n17335) );
  OAI21_X1 U20546 ( .B1(n18091), .B2(n17352), .A(n17335), .ZN(P3_U2783) );
  AOI22_X1 U20547 ( .A1(BUF2_REG_1__SCAN_IN), .A2(n17362), .B1(
        P3_LWORD_REG_1__SCAN_IN), .B2(n17349), .ZN(n17336) );
  OAI21_X1 U20548 ( .B1(n17337), .B2(n17364), .A(n17336), .ZN(P3_U2784) );
  AOI22_X1 U20549 ( .A1(P3_EAX_REG_2__SCAN_IN), .A2(n17350), .B1(
        P3_LWORD_REG_2__SCAN_IN), .B2(n17349), .ZN(n17338) );
  OAI21_X1 U20550 ( .B1(n18105), .B2(n17352), .A(n17338), .ZN(P3_U2785) );
  AOI22_X1 U20551 ( .A1(P3_EAX_REG_3__SCAN_IN), .A2(n17350), .B1(
        P3_LWORD_REG_3__SCAN_IN), .B2(n17361), .ZN(n17339) );
  OAI21_X1 U20552 ( .B1(n18111), .B2(n17352), .A(n17339), .ZN(P3_U2786) );
  AOI22_X1 U20553 ( .A1(P3_EAX_REG_4__SCAN_IN), .A2(n17350), .B1(
        P3_LWORD_REG_4__SCAN_IN), .B2(n17361), .ZN(n17340) );
  OAI21_X1 U20554 ( .B1(n18116), .B2(n17352), .A(n17340), .ZN(P3_U2787) );
  AOI22_X1 U20555 ( .A1(P3_EAX_REG_5__SCAN_IN), .A2(n17350), .B1(
        P3_LWORD_REG_5__SCAN_IN), .B2(n17361), .ZN(n17341) );
  OAI21_X1 U20556 ( .B1(n18122), .B2(n17352), .A(n17341), .ZN(P3_U2788) );
  AOI22_X1 U20557 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(n17350), .B1(
        P3_LWORD_REG_6__SCAN_IN), .B2(n17361), .ZN(n17342) );
  OAI21_X1 U20558 ( .B1(n18127), .B2(n17352), .A(n17342), .ZN(P3_U2789) );
  AOI22_X1 U20559 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n17362), .B1(
        P3_LWORD_REG_7__SCAN_IN), .B2(n17361), .ZN(n17343) );
  OAI21_X1 U20560 ( .B1(n17344), .B2(n17364), .A(n17343), .ZN(P3_U2790) );
  AOI22_X1 U20561 ( .A1(P3_EAX_REG_8__SCAN_IN), .A2(n17350), .B1(
        P3_LWORD_REG_8__SCAN_IN), .B2(n17349), .ZN(n17345) );
  OAI21_X1 U20562 ( .B1(n17346), .B2(n17352), .A(n17345), .ZN(P3_U2791) );
  AOI22_X1 U20563 ( .A1(P3_EAX_REG_9__SCAN_IN), .A2(n17350), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(n17349), .ZN(n17347) );
  OAI21_X1 U20564 ( .B1(n17348), .B2(n17352), .A(n17347), .ZN(P3_U2792) );
  AOI22_X1 U20565 ( .A1(P3_EAX_REG_10__SCAN_IN), .A2(n17350), .B1(
        P3_LWORD_REG_10__SCAN_IN), .B2(n17349), .ZN(n17351) );
  OAI21_X1 U20566 ( .B1(n17353), .B2(n17352), .A(n17351), .ZN(P3_U2793) );
  AOI22_X1 U20567 ( .A1(BUF2_REG_11__SCAN_IN), .A2(n17362), .B1(
        P3_LWORD_REG_11__SCAN_IN), .B2(n17361), .ZN(n17354) );
  OAI21_X1 U20568 ( .B1(n17355), .B2(n17364), .A(n17354), .ZN(P3_U2794) );
  AOI22_X1 U20569 ( .A1(BUF2_REG_12__SCAN_IN), .A2(n17362), .B1(
        P3_LWORD_REG_12__SCAN_IN), .B2(n17361), .ZN(n17356) );
  OAI21_X1 U20570 ( .B1(n21063), .B2(n17364), .A(n17356), .ZN(P3_U2795) );
  AOI22_X1 U20571 ( .A1(BUF2_REG_13__SCAN_IN), .A2(n17362), .B1(
        P3_LWORD_REG_13__SCAN_IN), .B2(n17361), .ZN(n17357) );
  OAI21_X1 U20572 ( .B1(n17358), .B2(n17364), .A(n17357), .ZN(P3_U2796) );
  AOI22_X1 U20573 ( .A1(BUF2_REG_14__SCAN_IN), .A2(n17362), .B1(
        P3_LWORD_REG_14__SCAN_IN), .B2(n17361), .ZN(n17359) );
  OAI21_X1 U20574 ( .B1(n17360), .B2(n17364), .A(n17359), .ZN(P3_U2797) );
  AOI22_X1 U20575 ( .A1(BUF2_REG_15__SCAN_IN), .A2(n17362), .B1(
        P3_LWORD_REG_15__SCAN_IN), .B2(n17361), .ZN(n17363) );
  OAI21_X1 U20576 ( .B1(n17365), .B2(n17364), .A(n17363), .ZN(P3_U2798) );
  INV_X1 U20577 ( .A(n17721), .ZN(n17451) );
  OAI22_X1 U20578 ( .A1(n17368), .A2(n17451), .B1(n17366), .B2(n17533), .ZN(
        n17367) );
  NOR2_X1 U20579 ( .A1(n17708), .A2(n17367), .ZN(n17396) );
  OAI21_X1 U20580 ( .B1(P3_PHYADDRPOINTER_REG_26__SCAN_IN), .B2(n17483), .A(
        n17396), .ZN(n17385) );
  NAND2_X1 U20581 ( .A1(n17368), .A2(n17531), .ZN(n17388) );
  AOI221_X1 U20582 ( .B1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C1(n17389), .C2(n17369), .A(
        n17388), .ZN(n17373) );
  OAI21_X1 U20583 ( .B1(n17598), .B2(n17371), .A(n17370), .ZN(n17372) );
  AOI211_X1 U20584 ( .C1(P3_PHYADDRPOINTER_REG_28__SCAN_IN), .C2(n17385), .A(
        n17373), .B(n17372), .ZN(n17383) );
  NAND2_X1 U20585 ( .A1(n17755), .A2(n17652), .ZN(n17481) );
  AOI22_X1 U20586 ( .A1(n17579), .A2(n17374), .B1(n17742), .B2(n17762), .ZN(
        n17402) );
  NAND2_X1 U20587 ( .A1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n17402), .ZN(
        n17391) );
  NAND3_X1 U20588 ( .A1(P3_INSTADDRPOINTER_REG_28__SCAN_IN), .A2(n17481), .A3(
        n17391), .ZN(n17382) );
  INV_X1 U20589 ( .A(n17480), .ZN(n17821) );
  NAND2_X1 U20590 ( .A1(n17821), .A2(n17540), .ZN(n17489) );
  NAND3_X1 U20591 ( .A1(n17376), .A2(n17502), .A3(n17375), .ZN(n17381) );
  OAI211_X1 U20592 ( .C1(n17379), .C2(n17378), .A(n17655), .B(n17377), .ZN(
        n17380) );
  NAND4_X1 U20593 ( .A1(n17383), .A2(n17382), .A3(n17381), .A4(n17380), .ZN(
        P3_U2802) );
  AOI22_X1 U20594 ( .A1(P3_PHYADDRPOINTER_REG_27__SCAN_IN), .A2(n17385), .B1(
        n17575), .B2(n17384), .ZN(n17395) );
  OAI21_X1 U20595 ( .B1(n17649), .B2(n17387), .A(n17386), .ZN(n17765) );
  INV_X1 U20596 ( .A(n17388), .ZN(n17390) );
  AOI22_X1 U20597 ( .A1(n17655), .A2(n17765), .B1(n17390), .B2(n17389), .ZN(
        n17394) );
  OAI21_X1 U20598 ( .B1(P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n17392), .A(
        n17391), .ZN(n17393) );
  NAND2_X1 U20599 ( .A1(n9820), .A2(P3_REIP_REG_27__SCAN_IN), .ZN(n17766) );
  NAND4_X1 U20600 ( .A1(n17395), .A2(n17394), .A3(n17393), .A4(n17766), .ZN(
        P3_U2803) );
  INV_X1 U20601 ( .A(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n17771) );
  NAND3_X1 U20602 ( .A1(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A3(n17771), .ZN(n17770) );
  NAND3_X1 U20603 ( .A1(n17433), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        n17502), .ZN(n17428) );
  NAND2_X1 U20604 ( .A1(n9820), .A2(P3_REIP_REG_26__SCAN_IN), .ZN(n17774) );
  INV_X1 U20605 ( .A(n17774), .ZN(n17406) );
  AOI221_X1 U20606 ( .B1(n18348), .B2(n17398), .C1(n17397), .C2(n17398), .A(
        n17396), .ZN(n17405) );
  AOI21_X1 U20607 ( .B1(n17598), .B2(n17483), .A(n17399), .ZN(n17404) );
  AOI21_X1 U20608 ( .B1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n17401), .A(
        n17400), .ZN(n17776) );
  OAI22_X1 U20609 ( .A1(n17402), .A2(n17771), .B1(n17776), .B2(n17555), .ZN(
        n17403) );
  NOR4_X1 U20610 ( .A1(n17406), .A2(n17405), .A3(n17404), .A4(n17403), .ZN(
        n17407) );
  OAI21_X1 U20611 ( .B1(n17770), .B2(n17428), .A(n17407), .ZN(P3_U2804) );
  NAND3_X1 U20612 ( .A1(n17792), .A2(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17778) );
  INV_X1 U20613 ( .A(n17778), .ZN(n17780) );
  NAND2_X1 U20614 ( .A1(n17780), .A2(n17896), .ZN(n17408) );
  XOR2_X1 U20615 ( .A(n17408), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17790) );
  NOR2_X1 U20616 ( .A1(n18074), .A2(n18670), .ZN(n17785) );
  OR2_X1 U20617 ( .A1(n18348), .A2(n17411), .ZN(n17443) );
  OAI211_X1 U20618 ( .C1(n17409), .C2(n17533), .A(n17750), .B(n17443), .ZN(
        n17440) );
  AOI21_X1 U20619 ( .B1(n17452), .B2(n17410), .A(n17440), .ZN(n17423) );
  NAND2_X1 U20620 ( .A1(n17411), .A2(n17531), .ZN(n17425) );
  OAI21_X1 U20621 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_25__SCAN_IN), .A(n17412), .ZN(n17413) );
  OAI22_X1 U20622 ( .A1(n17423), .A2(n17414), .B1(n17425), .B2(n17413), .ZN(
        n17415) );
  AOI211_X1 U20623 ( .C1(n17416), .C2(n17575), .A(n17785), .B(n17415), .ZN(
        n17422) );
  NAND3_X1 U20624 ( .A1(n17902), .A2(n17769), .A3(
        P3_INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n17417) );
  XOR2_X1 U20625 ( .A(n17417), .B(n17781), .Z(n17786) );
  AOI21_X1 U20626 ( .B1(n17419), .B2(n17604), .A(n17418), .ZN(n17420) );
  XOR2_X1 U20627 ( .A(n17420), .B(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .Z(
        n17787) );
  AOI22_X1 U20628 ( .A1(n17742), .A2(n17786), .B1(n17655), .B2(n17787), .ZN(
        n17421) );
  OAI211_X1 U20629 ( .C1(n17652), .C2(n17790), .A(n17422), .B(n17421), .ZN(
        P3_U2805) );
  NAND2_X1 U20630 ( .A1(n17902), .A2(n17769), .ZN(n17793) );
  NAND2_X1 U20631 ( .A1(n17896), .A2(n17769), .ZN(n17796) );
  AOI22_X1 U20632 ( .A1(n17742), .A2(n17793), .B1(n17579), .B2(n17796), .ZN(
        n17447) );
  NAND2_X1 U20633 ( .A1(n9820), .A2(P3_REIP_REG_24__SCAN_IN), .ZN(n17804) );
  OAI221_X1 U20634 ( .B1(P3_PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n17425), .C1(
        n17424), .C2(n17423), .A(n17804), .ZN(n17430) );
  AOI21_X1 U20635 ( .B1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n17427), .A(
        n17426), .ZN(n17806) );
  OAI22_X1 U20636 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n17428), .B1(
        n17806), .B2(n17555), .ZN(n17429) );
  AOI211_X1 U20637 ( .C1(n17575), .C2(n17431), .A(n17430), .B(n17429), .ZN(
        n17432) );
  OAI21_X1 U20638 ( .B1(n17447), .B2(n10167), .A(n17432), .ZN(P3_U2806) );
  NAND2_X1 U20639 ( .A1(n17433), .A2(n17502), .ZN(n17448) );
  AOI22_X1 U20640 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n17604), .B1(
        n17435), .B2(n17457), .ZN(n17436) );
  NAND2_X1 U20641 ( .A1(n17434), .A2(n17436), .ZN(n17437) );
  XOR2_X1 U20642 ( .A(n17437), .B(n17798), .Z(n17807) );
  NOR3_X1 U20643 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17483), .A3(
        n17438), .ZN(n17445) );
  AOI22_X1 U20644 ( .A1(P3_PHYADDRPOINTER_REG_23__SCAN_IN), .A2(n17440), .B1(
        n17575), .B2(n17439), .ZN(n17441) );
  NAND2_X1 U20645 ( .A1(n9820), .A2(P3_REIP_REG_23__SCAN_IN), .ZN(n17813) );
  OAI211_X1 U20646 ( .C1(n17443), .C2(n17442), .A(n17441), .B(n17813), .ZN(
        n17444) );
  AOI211_X1 U20647 ( .C1(n17807), .C2(n17655), .A(n17445), .B(n17444), .ZN(
        n17446) );
  OAI221_X1 U20648 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17448), 
        .C1(n17798), .C2(n17447), .A(n17446), .ZN(P3_U2807) );
  INV_X1 U20649 ( .A(n17533), .ZN(n17572) );
  AOI21_X1 U20650 ( .B1(n17572), .B2(n17449), .A(n17708), .ZN(n17450) );
  OAI21_X1 U20651 ( .B1(n17453), .B2(n17451), .A(n17450), .ZN(n17486) );
  AOI21_X1 U20652 ( .B1(n17452), .B2(n21050), .A(n17486), .ZN(n17466) );
  INV_X1 U20653 ( .A(P3_REIP_REG_22__SCAN_IN), .ZN(n18665) );
  NOR2_X1 U20654 ( .A1(n18074), .A2(n18665), .ZN(n17827) );
  NAND2_X1 U20655 ( .A1(n17453), .A2(n17531), .ZN(n17468) );
  AOI221_X1 U20656 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(
        P3_PHYADDRPOINTER_REG_21__SCAN_IN), .C1(n17465), .C2(n17467), .A(
        n17468), .ZN(n17454) );
  AOI211_X1 U20657 ( .C1(n17455), .C2(n17575), .A(n17827), .B(n17454), .ZN(
        n17464) );
  NAND2_X1 U20658 ( .A1(n17821), .A2(n17815), .ZN(n17822) );
  INV_X1 U20659 ( .A(n17434), .ZN(n17456) );
  AOI221_X1 U20660 ( .B1(n17529), .B2(n17457), .C1(n17822), .C2(n17457), .A(
        n17456), .ZN(n17458) );
  XOR2_X1 U20661 ( .A(n17458), .B(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(
        n17826) );
  NOR2_X1 U20662 ( .A1(n17459), .A2(n17822), .ZN(n17461) );
  OAI22_X1 U20663 ( .A1(n17896), .A2(n17652), .B1(n17902), .B2(n17755), .ZN(
        n17539) );
  AOI21_X1 U20664 ( .B1(n17481), .B2(n17822), .A(n17539), .ZN(n17479) );
  INV_X1 U20665 ( .A(n17479), .ZN(n17460) );
  MUX2_X1 U20666 ( .A(n17461), .B(n17460), .S(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .Z(n17462) );
  AOI21_X1 U20667 ( .B1(n17655), .B2(n17826), .A(n17462), .ZN(n17463) );
  OAI211_X1 U20668 ( .C1(n17466), .C2(n17465), .A(n17464), .B(n17463), .ZN(
        P3_U2808) );
  NAND2_X1 U20669 ( .A1(n9820), .A2(P3_REIP_REG_21__SCAN_IN), .ZN(n17838) );
  OAI221_X1 U20670 ( .B1(P3_PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n17468), .C1(
        n17467), .C2(n17466), .A(n17838), .ZN(n17469) );
  AOI21_X1 U20671 ( .B1(n17575), .B2(n17470), .A(n17469), .ZN(n17477) );
  INV_X1 U20672 ( .A(n17475), .ZN(n17834) );
  INV_X1 U20673 ( .A(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17516) );
  NOR3_X1 U20674 ( .A1(n17516), .A2(n17604), .A3(n17471), .ZN(n17500) );
  INV_X1 U20675 ( .A(n17472), .ZN(n17512) );
  AOI22_X1 U20676 ( .A1(n17834), .A2(n17500), .B1(n17512), .B2(n17473), .ZN(
        n17474) );
  XOR2_X1 U20677 ( .A(n17478), .B(n17474), .Z(n17832) );
  NOR2_X1 U20678 ( .A1(P3_INSTADDRPOINTER_REG_21__SCAN_IN), .A2(n17475), .ZN(
        n17833) );
  AOI22_X1 U20679 ( .A1(n17655), .A2(n17832), .B1(n17502), .B2(n17833), .ZN(
        n17476) );
  OAI211_X1 U20680 ( .C1(n17479), .C2(n17478), .A(n17477), .B(n17476), .ZN(
        P3_U2809) );
  NOR2_X1 U20681 ( .A1(n17480), .A2(n17855), .ZN(n17842) );
  INV_X1 U20682 ( .A(n17842), .ZN(n17817) );
  AOI21_X1 U20683 ( .B1(n17481), .B2(n17817), .A(n17539), .ZN(n17505) );
  INV_X1 U20684 ( .A(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n17492) );
  OAI221_X1 U20685 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17511), 
        .C1(n17855), .C2(n17500), .A(n17434), .ZN(n17482) );
  XOR2_X1 U20686 ( .A(n17492), .B(n17482), .Z(n17846) );
  NAND2_X1 U20687 ( .A1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .A2(n17492), .ZN(
        n17850) );
  NAND2_X1 U20688 ( .A1(n17598), .A2(n17483), .ZN(n17741) );
  OAI21_X1 U20689 ( .B1(n18348), .B2(n17484), .A(n21050), .ZN(n17485) );
  AOI22_X1 U20690 ( .A1(n17487), .A2(n17741), .B1(n17486), .B2(n17485), .ZN(
        n17488) );
  NAND2_X1 U20691 ( .A1(n9820), .A2(P3_REIP_REG_20__SCAN_IN), .ZN(n17848) );
  OAI211_X1 U20692 ( .C1(n17489), .C2(n17850), .A(n17488), .B(n17848), .ZN(
        n17490) );
  AOI21_X1 U20693 ( .B1(n17655), .B2(n17846), .A(n17490), .ZN(n17491) );
  OAI21_X1 U20694 ( .B1(n17505), .B2(n17492), .A(n17491), .ZN(P3_U2810) );
  AOI21_X1 U20695 ( .B1(n17721), .B2(n10181), .A(n17708), .ZN(n17527) );
  OAI21_X1 U20696 ( .B1(n17493), .B2(n17533), .A(n17527), .ZN(n17508) );
  NOR2_X1 U20697 ( .A1(n18074), .A2(n18659), .ZN(n17851) );
  NOR2_X1 U20698 ( .A1(n17509), .A2(n17494), .ZN(n17498) );
  OAI211_X1 U20699 ( .C1(P3_PHYADDRPOINTER_REG_18__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_19__SCAN_IN), .A(n17495), .B(n17531), .ZN(n17497) );
  OAI22_X1 U20700 ( .A1(n17498), .A2(n17497), .B1(n17496), .B2(n17598), .ZN(
        n17499) );
  AOI211_X1 U20701 ( .C1(P3_PHYADDRPOINTER_REG_19__SCAN_IN), .C2(n17508), .A(
        n17851), .B(n17499), .ZN(n17504) );
  AOI21_X1 U20702 ( .B1(n17511), .B2(n17512), .A(n17500), .ZN(n17501) );
  XOR2_X1 U20703 ( .A(n17855), .B(n17501), .Z(n17852) );
  AOI22_X1 U20704 ( .A1(n17655), .A2(n17852), .B1(n17502), .B2(n17855), .ZN(
        n17503) );
  OAI211_X1 U20705 ( .C1(n17505), .C2(n17855), .A(n17504), .B(n17503), .ZN(
        P3_U2811) );
  INV_X1 U20706 ( .A(n17865), .ZN(n17862) );
  AOI21_X1 U20707 ( .B1(n17540), .B2(n17862), .A(n17539), .ZN(n17522) );
  NOR2_X1 U20708 ( .A1(n17582), .A2(n10181), .ZN(n17510) );
  OAI22_X1 U20709 ( .A1(n18074), .A2(n18657), .B1(n17598), .B2(n17506), .ZN(
        n17507) );
  AOI221_X1 U20710 ( .B1(n17510), .B2(n17509), .C1(n17508), .C2(
        P3_PHYADDRPOINTER_REG_18__SCAN_IN), .A(n17507), .ZN(n17515) );
  AOI21_X1 U20711 ( .B1(n17649), .B2(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A(
        n17511), .ZN(n17513) );
  XOR2_X1 U20712 ( .A(n17513), .B(n17512), .Z(n17872) );
  NOR2_X1 U20713 ( .A1(P3_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n17862), .ZN(
        n17871) );
  AOI22_X1 U20714 ( .A1(n17655), .A2(n17872), .B1(n17540), .B2(n17871), .ZN(
        n17514) );
  OAI211_X1 U20715 ( .C1(n17522), .C2(n17516), .A(n17515), .B(n17514), .ZN(
        P3_U2812) );
  INV_X1 U20716 ( .A(n17517), .ZN(n17518) );
  AOI21_X1 U20717 ( .B1(n17518), .B2(n18476), .A(
        P3_PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n17526) );
  OAI21_X1 U20718 ( .B1(n17520), .B2(n17866), .A(n17519), .ZN(n17876) );
  AOI21_X1 U20719 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17540), .A(
        P3_INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n17521) );
  OAI22_X1 U20720 ( .A1(n17736), .A2(n17523), .B1(n17522), .B2(n17521), .ZN(
        n17524) );
  AOI21_X1 U20721 ( .B1(n17655), .B2(n17876), .A(n17524), .ZN(n17525) );
  NAND2_X1 U20722 ( .A1(n9820), .A2(P3_REIP_REG_17__SCAN_IN), .ZN(n17879) );
  OAI211_X1 U20723 ( .C1(n17527), .C2(n17526), .A(n17525), .B(n17879), .ZN(
        P3_U2813) );
  AOI21_X1 U20724 ( .B1(n17649), .B2(n17529), .A(n17528), .ZN(n17530) );
  XOR2_X1 U20725 ( .A(n17888), .B(n17530), .Z(n17893) );
  OAI211_X1 U20726 ( .C1(P3_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A(n17532), .B(n17531), .ZN(n17537) );
  INV_X1 U20727 ( .A(n17532), .ZN(n17544) );
  AOI21_X1 U20728 ( .B1(n17721), .B2(n17544), .A(n17708), .ZN(n17560) );
  OAI21_X1 U20729 ( .B1(n17534), .B2(n17533), .A(n17560), .ZN(n17547) );
  AOI22_X1 U20730 ( .A1(P3_PHYADDRPOINTER_REG_16__SCAN_IN), .A2(n17547), .B1(
        n17575), .B2(n17535), .ZN(n17536) );
  NAND2_X1 U20731 ( .A1(n9820), .A2(P3_REIP_REG_16__SCAN_IN), .ZN(n17891) );
  OAI211_X1 U20732 ( .C1(n10297), .C2(n17537), .A(n17536), .B(n17891), .ZN(
        n17538) );
  AOI221_X1 U20733 ( .B1(n17540), .B2(n17888), .C1(n17539), .C2(
        P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A(n17538), .ZN(n17541) );
  OAI21_X1 U20734 ( .B1(n17555), .B2(n17893), .A(n17541), .ZN(P3_U2814) );
  AND2_X1 U20735 ( .A1(n17542), .A2(n17604), .ZN(n17566) );
  NAND2_X1 U20736 ( .A1(n17941), .A2(n17647), .ZN(n17929) );
  NOR2_X1 U20737 ( .A1(n17604), .A2(n17929), .ZN(n17567) );
  NAND2_X1 U20738 ( .A1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .A2(n17934), .ZN(
        n17940) );
  OAI221_X1 U20739 ( .B1(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n17566), 
        .C1(n17910), .C2(n17567), .A(n17940), .ZN(n17543) );
  XOR2_X1 U20740 ( .A(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B(n17543), .Z(
        n17908) );
  NOR2_X1 U20741 ( .A1(n17582), .A2(n17544), .ZN(n17549) );
  OAI22_X1 U20742 ( .A1(n18074), .A2(n18651), .B1(n17598), .B2(n17545), .ZN(
        n17546) );
  AOI221_X1 U20743 ( .B1(n17549), .B2(n17548), .C1(n17547), .C2(
        P3_PHYADDRPOINTER_REG_15__SCAN_IN), .A(n17546), .ZN(n17554) );
  NOR2_X1 U20744 ( .A1(n17896), .A2(n17652), .ZN(n17552) );
  NAND2_X1 U20745 ( .A1(n17550), .A2(n17564), .ZN(n17895) );
  NOR2_X1 U20746 ( .A1(n17902), .A2(n17755), .ZN(n17551) );
  NAND2_X1 U20747 ( .A1(n17556), .A2(n17550), .ZN(n17903) );
  AOI22_X1 U20748 ( .A1(n17552), .A2(n17895), .B1(n17551), .B2(n17903), .ZN(
        n17553) );
  OAI211_X1 U20749 ( .C1(n17555), .C2(n17908), .A(n17554), .B(n17553), .ZN(
        P3_U2815) );
  OAI21_X1 U20750 ( .B1(n17557), .B2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17556), .ZN(n17925) );
  AND2_X1 U20751 ( .A1(n18476), .A2(n17558), .ZN(n17645) );
  NAND2_X1 U20752 ( .A1(n17559), .A2(n17645), .ZN(n17610) );
  AOI221_X1 U20753 ( .B1(n17583), .B2(n17561), .C1(n17610), .C2(n17561), .A(
        n17560), .ZN(n17562) );
  INV_X1 U20754 ( .A(P3_REIP_REG_14__SCAN_IN), .ZN(n18649) );
  NOR2_X1 U20755 ( .A1(n18074), .A2(n18649), .ZN(n17920) );
  AOI211_X1 U20756 ( .C1(n17563), .C2(n17741), .A(n17562), .B(n17920), .ZN(
        n17570) );
  INV_X1 U20757 ( .A(n17564), .ZN(n17565) );
  AOI221_X1 U20758 ( .B1(n17576), .B2(n17910), .C1(n17914), .C2(n17910), .A(
        n17565), .ZN(n17921) );
  OAI21_X1 U20759 ( .B1(n17567), .B2(n17566), .A(n17940), .ZN(n17568) );
  XOR2_X1 U20760 ( .A(n17568), .B(n17910), .Z(n17922) );
  AOI22_X1 U20761 ( .A1(n17579), .A2(n17921), .B1(n17655), .B2(n17922), .ZN(
        n17569) );
  OAI211_X1 U20762 ( .C1(n17755), .C2(n17925), .A(n17570), .B(n17569), .ZN(
        P3_U2816) );
  AOI22_X1 U20763 ( .A1(n17572), .A2(n17571), .B1(n17721), .B2(n17581), .ZN(
        n17573) );
  NAND2_X1 U20764 ( .A1(n17573), .A2(n17750), .ZN(n17593) );
  AOI22_X1 U20765 ( .A1(P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A2(n17593), .B1(
        n17575), .B2(n17574), .ZN(n17586) );
  INV_X1 U20766 ( .A(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17951) );
  AOI22_X1 U20767 ( .A1(n17941), .A2(n17647), .B1(n17951), .B2(n17604), .ZN(
        n17577) );
  AOI21_X1 U20768 ( .B1(n17587), .B2(n17604), .A(n17577), .ZN(n17578) );
  XOR2_X1 U20769 ( .A(n17578), .B(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .Z(
        n17937) );
  AOI22_X1 U20770 ( .A1(n17579), .A2(n17929), .B1(n17742), .B2(n17930), .ZN(
        n17601) );
  INV_X1 U20771 ( .A(n17643), .ZN(n17607) );
  NAND2_X1 U20772 ( .A1(n17926), .A2(n17607), .ZN(n17602) );
  OAI22_X1 U20773 ( .A1(n17601), .A2(n17934), .B1(n17940), .B2(n17602), .ZN(
        n17580) );
  AOI21_X1 U20774 ( .B1(n17655), .B2(n17937), .A(n17580), .ZN(n17585) );
  NAND2_X1 U20775 ( .A1(n9820), .A2(P3_REIP_REG_13__SCAN_IN), .ZN(n17938) );
  NOR2_X1 U20776 ( .A1(n17582), .A2(n17581), .ZN(n17595) );
  OAI211_X1 U20777 ( .C1(P3_PHYADDRPOINTER_REG_12__SCAN_IN), .C2(
        P3_PHYADDRPOINTER_REG_13__SCAN_IN), .A(n17595), .B(n17583), .ZN(n17584) );
  NAND4_X1 U20778 ( .A1(n17586), .A2(n17585), .A3(n17938), .A4(n17584), .ZN(
        P3_U2817) );
  INV_X1 U20779 ( .A(n17587), .ZN(n17590) );
  INV_X1 U20780 ( .A(n17926), .ZN(n17588) );
  NOR2_X1 U20781 ( .A1(n17588), .A2(n17576), .ZN(n17589) );
  MUX2_X1 U20782 ( .A(n17590), .B(n17589), .S(n17649), .Z(n17591) );
  XOR2_X1 U20783 ( .A(n17591), .B(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .Z(
        n17949) );
  INV_X1 U20784 ( .A(n17592), .ZN(n17597) );
  NOR2_X1 U20785 ( .A1(n18074), .A2(n18645), .ZN(n17948) );
  AOI221_X1 U20786 ( .B1(n17595), .B2(n17594), .C1(n17593), .C2(
        P3_PHYADDRPOINTER_REG_12__SCAN_IN), .A(n17948), .ZN(n17596) );
  OAI21_X1 U20787 ( .B1(n17598), .B2(n17597), .A(n17596), .ZN(n17599) );
  AOI21_X1 U20788 ( .B1(n17655), .B2(n17949), .A(n17599), .ZN(n17600) );
  OAI221_X1 U20789 ( .B1(P3_INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n17602), 
        .C1(n17951), .C2(n17601), .A(n17600), .ZN(P3_U2818) );
  INV_X1 U20790 ( .A(n17959), .ZN(n17927) );
  NAND2_X1 U20791 ( .A1(n17927), .A2(n17608), .ZN(n17965) );
  NAND2_X1 U20792 ( .A1(n17604), .A2(n17646), .ZN(n17632) );
  INV_X1 U20793 ( .A(n17632), .ZN(n17622) );
  OR4_X1 U20794 ( .A1(n17988), .A2(n18009), .A3(n17604), .A4(n17603), .ZN(
        n17631) );
  NOR2_X1 U20795 ( .A1(n17959), .A2(n17631), .ZN(n17625) );
  AOI21_X1 U20796 ( .B1(n17630), .B2(n17622), .A(n17625), .ZN(n17605) );
  XOR2_X1 U20797 ( .A(n17608), .B(n17605), .Z(n17952) );
  OAI22_X1 U20798 ( .A1(n17606), .A2(n17755), .B1(n17652), .B2(n17647), .ZN(
        n17626) );
  INV_X1 U20799 ( .A(n17626), .ZN(n17642) );
  NAND2_X1 U20800 ( .A1(n17959), .A2(n17607), .ZN(n17629) );
  AOI21_X1 U20801 ( .B1(n17642), .B2(n17629), .A(n17608), .ZN(n17615) );
  NAND2_X1 U20802 ( .A1(n17609), .A2(n17645), .ZN(n17634) );
  NOR2_X1 U20803 ( .A1(n17618), .A2(n17634), .ZN(n17617) );
  INV_X1 U20804 ( .A(n17746), .ZN(n17635) );
  OAI211_X1 U20805 ( .C1(n17617), .C2(P3_PHYADDRPOINTER_REG_11__SCAN_IN), .A(
        n17635), .B(n17610), .ZN(n17612) );
  NAND2_X1 U20806 ( .A1(n9820), .A2(P3_REIP_REG_11__SCAN_IN), .ZN(n17611) );
  OAI211_X1 U20807 ( .C1(n17736), .C2(n17613), .A(n17612), .B(n17611), .ZN(
        n17614) );
  AOI211_X1 U20808 ( .C1(n17655), .C2(n17952), .A(n17615), .B(n17614), .ZN(
        n17616) );
  OAI21_X1 U20809 ( .B1(n17643), .B2(n17965), .A(n17616), .ZN(P3_U2819) );
  AOI211_X1 U20810 ( .C1(n17634), .C2(n17618), .A(n17746), .B(n17617), .ZN(
        n17620) );
  NOR2_X1 U20811 ( .A1(n18074), .A2(n18641), .ZN(n17619) );
  AOI211_X1 U20812 ( .C1(n17621), .C2(n17741), .A(n17620), .B(n17619), .ZN(
        n17628) );
  INV_X1 U20813 ( .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17979) );
  NOR2_X1 U20814 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17979), .ZN(
        n17970) );
  INV_X1 U20815 ( .A(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17623) );
  AOI221_X1 U20816 ( .B1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .B2(n17632), 
        .C1(n17623), .C2(n17622), .A(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(
        n17624) );
  AOI211_X1 U20817 ( .C1(n17970), .C2(n17631), .A(n17625), .B(n17624), .ZN(
        n17971) );
  AOI22_X1 U20818 ( .A1(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n17626), .B1(
        n17655), .B2(n17971), .ZN(n17627) );
  OAI211_X1 U20819 ( .C1(n17630), .C2(n17629), .A(n17628), .B(n17627), .ZN(
        P3_U2820) );
  NAND2_X1 U20820 ( .A1(n17632), .A2(n17631), .ZN(n17633) );
  XOR2_X1 U20821 ( .A(n17633), .B(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .Z(
        n17981) );
  NOR2_X1 U20822 ( .A1(n18074), .A2(n18640), .ZN(n17640) );
  INV_X1 U20823 ( .A(n17634), .ZN(n17638) );
  AOI22_X1 U20824 ( .A1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A2(n17635), .B1(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(n17645), .ZN(n17637) );
  OAI22_X1 U20825 ( .A1(n17638), .A2(n17637), .B1(n17736), .B2(n17636), .ZN(
        n17639) );
  AOI211_X1 U20826 ( .C1(n17655), .C2(n17981), .A(n17640), .B(n17639), .ZN(
        n17641) );
  OAI221_X1 U20827 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17643), .C1(
        n17979), .C2(n17642), .A(n17641), .ZN(P3_U2821) );
  AOI21_X1 U20828 ( .B1(n17721), .B2(n17664), .A(n17708), .ZN(n17666) );
  OAI21_X1 U20829 ( .B1(P3_PHYADDRPOINTER_REG_7__SCAN_IN), .B2(n18348), .A(
        n17666), .ZN(n17644) );
  NOR2_X1 U20830 ( .A1(n18074), .A2(n18638), .ZN(n17989) );
  AOI221_X1 U20831 ( .B1(n17645), .B2(n21012), .C1(n17644), .C2(
        P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A(n17989), .ZN(n17657) );
  INV_X1 U20832 ( .A(n17646), .ZN(n17648) );
  AND2_X1 U20833 ( .A1(n17648), .A2(n17576), .ZN(n17996) );
  AOI21_X1 U20834 ( .B1(n17649), .B2(n17653), .A(n10292), .ZN(n17993) );
  OAI21_X1 U20835 ( .B1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .B2(n17651), .A(
        n17650), .ZN(n17999) );
  OAI22_X1 U20836 ( .A1(n17653), .A2(n17652), .B1(n17755), .B2(n17999), .ZN(
        n17654) );
  AOI21_X1 U20837 ( .B1(n17655), .B2(n17993), .A(n17654), .ZN(n17656) );
  OAI211_X1 U20838 ( .C1(n17736), .C2(n17658), .A(n17657), .B(n17656), .ZN(
        P3_U2822) );
  NOR2_X1 U20839 ( .A1(n17659), .A2(n17661), .ZN(n17662) );
  OAI22_X1 U20840 ( .A1(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .A2(n17662), .B1(
        n17661), .B2(n17660), .ZN(n18003) );
  NAND2_X1 U20841 ( .A1(n18476), .A2(n17665), .ZN(n17663) );
  OAI22_X1 U20842 ( .A1(n17666), .A2(n17665), .B1(n17664), .B2(n17663), .ZN(
        n17667) );
  AOI21_X1 U20843 ( .B1(n9820), .B2(P3_REIP_REG_7__SCAN_IN), .A(n17667), .ZN(
        n17672) );
  AOI21_X1 U20844 ( .B1(n18009), .B2(n17669), .A(n17668), .ZN(n18005) );
  AOI22_X1 U20845 ( .A1(n17738), .A2(n18005), .B1(n17670), .B2(n17741), .ZN(
        n17671) );
  OAI211_X1 U20846 ( .C1(n17755), .C2(n18003), .A(n17672), .B(n17671), .ZN(
        P3_U2823) );
  AOI21_X1 U20847 ( .B1(n9928), .B2(n17674), .A(n17673), .ZN(n18016) );
  NAND2_X1 U20848 ( .A1(n18476), .A2(n17684), .ZN(n17675) );
  OAI22_X1 U20849 ( .A1(P3_PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n17675), .B1(
        n18074), .B2(n21078), .ZN(n17676) );
  AOI21_X1 U20850 ( .B1(n17738), .B2(n18016), .A(n17676), .ZN(n17686) );
  AOI22_X1 U20851 ( .A1(n17679), .A2(n17690), .B1(n17678), .B2(n17677), .ZN(
        n17683) );
  AOI22_X1 U20852 ( .A1(n17681), .A2(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .B1(
        n18019), .B2(n17680), .ZN(n17682) );
  XNOR2_X1 U20853 ( .A(n17683), .B(n17682), .ZN(n18015) );
  AOI21_X1 U20854 ( .B1(n17684), .B2(n18476), .A(n17746), .ZN(n17696) );
  AOI22_X1 U20855 ( .A1(n17742), .A2(n18015), .B1(
        P3_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n17696), .ZN(n17685) );
  OAI211_X1 U20856 ( .C1(n17736), .C2(n17687), .A(n17686), .B(n17685), .ZN(
        P3_U2824) );
  AOI21_X1 U20857 ( .B1(n18026), .B2(n17689), .A(n17688), .ZN(n18023) );
  AOI22_X1 U20858 ( .A1(n9820), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n17738), .B2(
        n18023), .ZN(n17698) );
  AOI21_X1 U20859 ( .B1(n17692), .B2(n17691), .A(n17690), .ZN(n18020) );
  OAI21_X1 U20860 ( .B1(n17708), .B2(n17694), .A(n17693), .ZN(n17695) );
  AOI22_X1 U20861 ( .A1(n17742), .A2(n18020), .B1(n17696), .B2(n17695), .ZN(
        n17697) );
  OAI211_X1 U20862 ( .C1(n17736), .C2(n17699), .A(n17698), .B(n17697), .ZN(
        P3_U2825) );
  AOI21_X1 U20863 ( .B1(n17702), .B2(n17701), .A(n17700), .ZN(n18028) );
  OAI22_X1 U20864 ( .A1(n18074), .A2(n18631), .B1(n18348), .B2(n17703), .ZN(
        n17704) );
  AOI21_X1 U20865 ( .B1(n17738), .B2(n18028), .A(n17704), .ZN(n17710) );
  AOI21_X1 U20866 ( .B1(n17707), .B2(n17706), .A(n17705), .ZN(n18029) );
  NOR2_X1 U20867 ( .A1(n17708), .A2(n21053), .ZN(n17731) );
  AOI21_X1 U20868 ( .B1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .B2(n17731), .A(
        n17746), .ZN(n17719) );
  AOI22_X1 U20869 ( .A1(n17742), .A2(n18029), .B1(
        P3_PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n17719), .ZN(n17709) );
  OAI211_X1 U20870 ( .C1(n17736), .C2(n17711), .A(n17710), .B(n17709), .ZN(
        P3_U2826) );
  AOI21_X1 U20871 ( .B1(n17714), .B2(n17713), .A(n17712), .ZN(n18036) );
  AOI21_X1 U20872 ( .B1(n17717), .B2(n17716), .A(n17715), .ZN(n18038) );
  AOI22_X1 U20873 ( .A1(n17742), .A2(n18036), .B1(n17738), .B2(n18038), .ZN(
        n17724) );
  AOI22_X1 U20874 ( .A1(P3_PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n17719), .B1(
        n17718), .B2(n17741), .ZN(n17723) );
  NAND3_X1 U20875 ( .A1(n17721), .A2(n17731), .A3(n17720), .ZN(n17722) );
  NAND2_X1 U20876 ( .A1(n9820), .A2(P3_REIP_REG_3__SCAN_IN), .ZN(n18039) );
  NAND4_X1 U20877 ( .A1(n17724), .A2(n17723), .A3(n17722), .A4(n18039), .ZN(
        P3_U2827) );
  AOI21_X1 U20878 ( .B1(n17727), .B2(n17726), .A(n17725), .ZN(n18054) );
  AOI22_X1 U20879 ( .A1(n9820), .A2(P3_REIP_REG_2__SCAN_IN), .B1(n17738), .B2(
        n18054), .ZN(n17734) );
  AOI21_X1 U20880 ( .B1(n17730), .B2(n17729), .A(n17728), .ZN(n18053) );
  AOI21_X1 U20881 ( .B1(n18348), .B2(n21053), .A(n17731), .ZN(n17732) );
  AOI21_X1 U20882 ( .B1(n18053), .B2(n17742), .A(n17732), .ZN(n17733) );
  OAI211_X1 U20883 ( .C1(n17736), .C2(n17735), .A(n17734), .B(n17733), .ZN(
        P3_U2828) );
  AOI21_X1 U20884 ( .B1(n17740), .B2(n17747), .A(n17737), .ZN(n18065) );
  AOI22_X1 U20885 ( .A1(n9820), .A2(P3_REIP_REG_1__SCAN_IN), .B1(n17738), .B2(
        n18065), .ZN(n17744) );
  OAI21_X1 U20886 ( .B1(n17749), .B2(n17740), .A(n17739), .ZN(n18059) );
  AOI22_X1 U20887 ( .A1(n17742), .A2(n18059), .B1(n17745), .B2(n17741), .ZN(
        n17743) );
  OAI211_X1 U20888 ( .C1(n17746), .C2(n17745), .A(n17744), .B(n17743), .ZN(
        P3_U2829) );
  INV_X1 U20889 ( .A(n17747), .ZN(n17748) );
  NOR2_X1 U20890 ( .A1(n17749), .A2(n17748), .ZN(n18080) );
  INV_X1 U20891 ( .A(n18080), .ZN(n18078) );
  NAND2_X1 U20892 ( .A1(n18706), .A2(n18603), .ZN(n18607) );
  INV_X1 U20893 ( .A(n18607), .ZN(n18749) );
  OAI21_X1 U20894 ( .B1(n17751), .B2(n18749), .A(n17750), .ZN(n17752) );
  AOI22_X1 U20895 ( .A1(n9820), .A2(P3_REIP_REG_0__SCAN_IN), .B1(
        P3_PHYADDRPOINTER_REG_0__SCAN_IN), .B2(n17752), .ZN(n17753) );
  OAI221_X1 U20896 ( .B1(n18080), .B2(n17755), .C1(n18078), .C2(n17754), .A(
        n17753), .ZN(P3_U2830) );
  AOI221_X1 U20897 ( .B1(n17809), .B2(n17768), .C1(n17756), .C2(n17768), .A(
        n18061), .ZN(n17764) );
  NOR2_X1 U20898 ( .A1(n18554), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n18046) );
  NOR2_X1 U20899 ( .A1(n18046), .A2(n17818), .ZN(n17859) );
  AOI21_X1 U20900 ( .B1(n17859), .B2(n17780), .A(n17858), .ZN(n17777) );
  AOI22_X1 U20901 ( .A1(n18549), .A2(n17781), .B1(n18566), .B2(n17757), .ZN(
        n17759) );
  OAI211_X1 U20902 ( .C1(n17760), .C2(n17897), .A(n17759), .B(n17758), .ZN(
        n17761) );
  AOI211_X1 U20903 ( .C1(n18052), .C2(n17762), .A(n17777), .B(n17761), .ZN(
        n17772) );
  OAI211_X1 U20904 ( .C1(n18568), .C2(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_27__SCAN_IN), .B(n17772), .ZN(n17763) );
  AOI22_X1 U20905 ( .A1(n17994), .A2(n17765), .B1(n17764), .B2(n17763), .ZN(
        n17767) );
  OAI211_X1 U20906 ( .C1(n18062), .C2(n17768), .A(n17767), .B(n17766), .ZN(
        P3_U2835) );
  INV_X1 U20907 ( .A(n17769), .ZN(n17797) );
  OR2_X1 U20908 ( .A1(n17797), .A2(n17809), .ZN(n17801) );
  OAI22_X1 U20909 ( .A1(n17772), .A2(n17771), .B1(n17770), .B2(n17801), .ZN(
        n17773) );
  AOI22_X1 U20910 ( .A1(P3_INSTADDRPOINTER_REG_26__SCAN_IN), .A2(n18055), .B1(
        n18073), .B2(n17773), .ZN(n17775) );
  OAI211_X1 U20911 ( .C1(n17776), .C2(n17909), .A(n17775), .B(n17774), .ZN(
        P3_U2836) );
  AOI221_X1 U20912 ( .B1(n17861), .B2(n18540), .C1(n17778), .C2(n18540), .A(
        n17777), .ZN(n17783) );
  NAND2_X1 U20913 ( .A1(n17780), .A2(n17779), .ZN(n17782) );
  AOI221_X1 U20914 ( .B1(n17783), .B2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), 
        .C1(n17782), .C2(n17781), .A(n18061), .ZN(n17784) );
  AOI211_X1 U20915 ( .C1(n18055), .C2(P3_INSTADDRPOINTER_REG_25__SCAN_IN), .A(
        n17785), .B(n17784), .ZN(n17789) );
  AOI22_X1 U20916 ( .A1(n17994), .A2(n17787), .B1(n18037), .B2(n17786), .ZN(
        n17788) );
  OAI211_X1 U20917 ( .C1(n17791), .C2(n17790), .A(n17789), .B(n17788), .ZN(
        P3_U2837) );
  INV_X1 U20918 ( .A(n17897), .ZN(n17953) );
  AND2_X1 U20919 ( .A1(n17792), .A2(n17859), .ZN(n17816) );
  INV_X1 U20920 ( .A(n17793), .ZN(n17794) );
  OAI22_X1 U20921 ( .A1(n17858), .A2(n17816), .B1(n17794), .B2(n18534), .ZN(
        n17795) );
  AOI211_X1 U20922 ( .C1(n17953), .C2(n17796), .A(n18055), .B(n17795), .ZN(
        n17800) );
  AOI21_X1 U20923 ( .B1(n17887), .B2(n17800), .A(n10167), .ZN(n17803) );
  OAI22_X1 U20924 ( .A1(n18540), .A2(n17798), .B1(n17861), .B2(n17797), .ZN(
        n17799) );
  AOI21_X1 U20925 ( .B1(n17800), .B2(n17799), .A(n9820), .ZN(n17810) );
  NOR3_X1 U20926 ( .A1(P3_INSTADDRPOINTER_REG_24__SCAN_IN), .A2(n18061), .A3(
        n17801), .ZN(n17802) );
  AOI21_X1 U20927 ( .B1(n17803), .B2(n17810), .A(n17802), .ZN(n17805) );
  OAI211_X1 U20928 ( .C1(n17806), .C2(n17909), .A(n17805), .B(n17804), .ZN(
        P3_U2838) );
  INV_X1 U20929 ( .A(n17807), .ZN(n17814) );
  NOR3_X1 U20930 ( .A1(n18055), .A2(n17809), .A3(n17808), .ZN(n17811) );
  OAI21_X1 U20931 ( .B1(P3_INSTADDRPOINTER_REG_23__SCAN_IN), .B2(n17811), .A(
        n17810), .ZN(n17812) );
  OAI211_X1 U20932 ( .C1(n17814), .C2(n17909), .A(n17813), .B(n17812), .ZN(
        P3_U2839) );
  AOI22_X1 U20933 ( .A1(n17815), .A2(n17840), .B1(
        P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18073), .ZN(n17831) );
  INV_X1 U20934 ( .A(n17815), .ZN(n17825) );
  AOI21_X1 U20935 ( .B1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n18554), .A(
        n17816), .ZN(n17824) );
  NOR2_X1 U20936 ( .A1(n18052), .A2(n17953), .ZN(n17864) );
  INV_X1 U20937 ( .A(n17864), .ZN(n17958) );
  OAI22_X1 U20938 ( .A1(n17902), .A2(n18534), .B1(n17896), .B2(n17897), .ZN(
        n17857) );
  AOI221_X1 U20939 ( .B1(n17818), .B2(n18549), .C1(n17817), .C2(n18549), .A(
        n17857), .ZN(n17819) );
  OAI221_X1 U20940 ( .B1(n18561), .B2(n17821), .C1(n18561), .C2(n17820), .A(
        n17819), .ZN(n17844) );
  AOI21_X1 U20941 ( .B1(n17822), .B2(n17958), .A(n17844), .ZN(n17823) );
  OAI21_X1 U20942 ( .B1(n18568), .B2(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A(
        n17823), .ZN(n17836) );
  AOI211_X1 U20943 ( .C1(n17933), .C2(n17825), .A(n17824), .B(n17836), .ZN(
        n17830) );
  AOI22_X1 U20944 ( .A1(P3_INSTADDRPOINTER_REG_22__SCAN_IN), .A2(n18055), .B1(
        n17994), .B2(n17826), .ZN(n17829) );
  INV_X1 U20945 ( .A(n17827), .ZN(n17828) );
  OAI211_X1 U20946 ( .C1(n17831), .C2(n17830), .A(n17829), .B(n17828), .ZN(
        P3_U2840) );
  AOI22_X1 U20947 ( .A1(n17840), .A2(n17833), .B1(n17994), .B2(n17832), .ZN(
        n17839) );
  NOR2_X1 U20948 ( .A1(n18540), .A2(n18566), .ZN(n18060) );
  OAI211_X1 U20949 ( .C1(n17834), .C2(n18060), .A(n18073), .B(n17841), .ZN(
        n17835) );
  OAI211_X1 U20950 ( .C1(n17836), .C2(n17835), .A(
        P3_INSTADDRPOINTER_REG_21__SCAN_IN), .B(n18074), .ZN(n17837) );
  NAND3_X1 U20951 ( .A1(n17839), .A2(n17838), .A3(n17837), .ZN(P3_U2841) );
  INV_X1 U20952 ( .A(n17840), .ZN(n17856) );
  NAND2_X1 U20953 ( .A1(n17855), .A2(P3_STATE2_REG_2__SCAN_IN), .ZN(n17845) );
  OAI211_X1 U20954 ( .C1(n17842), .C2(n17864), .A(n18073), .B(n17841), .ZN(
        n17843) );
  OAI21_X1 U20955 ( .B1(n17844), .B2(n17843), .A(n18074), .ZN(n17854) );
  OAI21_X1 U20956 ( .B1(n18060), .B2(n17845), .A(n17854), .ZN(n17847) );
  AOI22_X1 U20957 ( .A1(P3_INSTADDRPOINTER_REG_20__SCAN_IN), .A2(n17847), .B1(
        n17994), .B2(n17846), .ZN(n17849) );
  OAI211_X1 U20958 ( .C1(n17856), .C2(n17850), .A(n17849), .B(n17848), .ZN(
        P3_U2842) );
  AOI21_X1 U20959 ( .B1(n17994), .B2(n17852), .A(n17851), .ZN(n17853) );
  OAI221_X1 U20960 ( .B1(P3_INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n17856), 
        .C1(n17855), .C2(n17854), .A(n17853), .ZN(P3_U2843) );
  NOR2_X1 U20961 ( .A1(n18061), .A2(n17857), .ZN(n17886) );
  AOI21_X1 U20962 ( .B1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .B2(n17859), .A(
        n17858), .ZN(n17860) );
  AOI221_X1 U20963 ( .B1(n17862), .B2(n18540), .C1(n17861), .C2(n18540), .A(
        n17860), .ZN(n17863) );
  OAI211_X1 U20964 ( .C1(n17865), .C2(n17864), .A(n17886), .B(n17863), .ZN(
        n17877) );
  OAI221_X1 U20965 ( .B1(n17877), .B2(n17866), .C1(n17877), .C2(n18045), .A(
        P3_INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n17874) );
  OAI22_X1 U20966 ( .A1(n18561), .A2(n17984), .B1(n17985), .B2(n18044), .ZN(
        n17867) );
  NOR2_X1 U20967 ( .A1(n18035), .A2(n17868), .ZN(n17915) );
  OAI21_X1 U20968 ( .B1(n17915), .B2(n17869), .A(n18073), .ZN(n17964) );
  NOR2_X1 U20969 ( .A1(n17870), .A2(n17964), .ZN(n17889) );
  AOI22_X1 U20970 ( .A1(n17994), .A2(n17872), .B1(n17889), .B2(n17871), .ZN(
        n17873) );
  OAI221_X1 U20971 ( .B1(n9820), .B2(n17874), .C1(n18074), .C2(n18657), .A(
        n17873), .ZN(P3_U2844) );
  NOR2_X1 U20972 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n17888), .ZN(
        n17875) );
  AOI22_X1 U20973 ( .A1(n17994), .A2(n17876), .B1(n17889), .B2(n17875), .ZN(
        n17880) );
  NAND3_X1 U20974 ( .A1(P3_INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n18074), .A3(
        n17877), .ZN(n17878) );
  NAND3_X1 U20975 ( .A1(n17880), .A2(n17879), .A3(n17878), .ZN(P3_U2845) );
  NAND2_X1 U20976 ( .A1(n18554), .A2(P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(
        n17884) );
  NAND2_X1 U20977 ( .A1(n18540), .A2(n17881), .ZN(n17955) );
  AOI21_X1 U20978 ( .B1(n17894), .B2(n17955), .A(n17967), .ZN(n17883) );
  NOR2_X1 U20979 ( .A1(n18568), .A2(n17882), .ZN(n17969) );
  AOI211_X1 U20980 ( .C1(n17885), .C2(n17884), .A(n17883), .B(n17969), .ZN(
        n17901) );
  AOI221_X1 U20981 ( .B1(n17887), .B2(n17886), .C1(n17901), .C2(n17886), .A(
        n9820), .ZN(n17890) );
  AOI22_X1 U20982 ( .A1(P3_INSTADDRPOINTER_REG_16__SCAN_IN), .A2(n17890), .B1(
        n17889), .B2(n17888), .ZN(n17892) );
  OAI211_X1 U20983 ( .C1(n17893), .C2(n17909), .A(n17892), .B(n17891), .ZN(
        P3_U2846) );
  AOI22_X1 U20984 ( .A1(n9820), .A2(P3_REIP_REG_15__SCAN_IN), .B1(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .B2(n18055), .ZN(n17907) );
  AOI21_X1 U20985 ( .B1(n17894), .B2(n17915), .A(
        P3_INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n17900) );
  INV_X1 U20986 ( .A(n17895), .ZN(n17899) );
  OR2_X1 U20987 ( .A1(n17897), .A2(n17896), .ZN(n17898) );
  OAI22_X1 U20988 ( .A1(n17901), .A2(n17900), .B1(n17899), .B2(n17898), .ZN(
        n17905) );
  NOR2_X1 U20989 ( .A1(n17902), .A2(n18079), .ZN(n17904) );
  AOI22_X1 U20990 ( .A1(n18073), .A2(n17905), .B1(n17904), .B2(n17903), .ZN(
        n17906) );
  OAI211_X1 U20991 ( .C1(n17909), .C2(n17908), .A(n17907), .B(n17906), .ZN(
        P3_U2847) );
  AOI21_X1 U20992 ( .B1(n17941), .B2(n17974), .A(n18554), .ZN(n17932) );
  AOI211_X1 U20993 ( .C1(n18540), .C2(n17911), .A(n17969), .B(n17910), .ZN(
        n17912) );
  OAI211_X1 U20994 ( .C1(P3_INSTADDRPOINTER_REG_13__SCAN_IN), .C2(n18060), .A(
        n17912), .B(n17955), .ZN(n17913) );
  AOI211_X1 U20995 ( .C1(n18549), .C2(n17914), .A(n17932), .B(n17913), .ZN(
        n17918) );
  AOI21_X1 U20996 ( .B1(n17916), .B2(n17915), .A(
        P3_INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n17917) );
  NOR3_X1 U20997 ( .A1(n17918), .A2(n17917), .A3(n18061), .ZN(n17919) );
  AOI211_X1 U20998 ( .C1(n18055), .C2(P3_INSTADDRPOINTER_REG_14__SCAN_IN), .A(
        n17920), .B(n17919), .ZN(n17924) );
  AOI22_X1 U20999 ( .A1(n17994), .A2(n17922), .B1(n17995), .B2(n17921), .ZN(
        n17923) );
  OAI211_X1 U21000 ( .C1(n18079), .C2(n17925), .A(n17924), .B(n17923), .ZN(
        P3_U2848) );
  INV_X1 U21001 ( .A(n17964), .ZN(n17980) );
  NAND2_X1 U21002 ( .A1(n17926), .A2(n17980), .ZN(n17946) );
  OAI21_X1 U21003 ( .B1(n18568), .B2(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A(
        P3_INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n17942) );
  OAI22_X1 U21004 ( .A1(n18568), .A2(n17927), .B1(n17926), .B2(n18561), .ZN(
        n17928) );
  NOR2_X1 U21005 ( .A1(n17969), .A2(n17928), .ZN(n17960) );
  AOI22_X1 U21006 ( .A1(n18052), .A2(n17930), .B1(n17953), .B2(n17929), .ZN(
        n17931) );
  NAND3_X1 U21007 ( .A1(n17960), .A2(n17931), .A3(n17955), .ZN(n17943) );
  AOI211_X1 U21008 ( .C1(n17933), .C2(n17942), .A(n17932), .B(n17943), .ZN(
        n17935) );
  AOI211_X1 U21009 ( .C1(n18073), .C2(n17935), .A(n9820), .B(n17934), .ZN(
        n17936) );
  AOI21_X1 U21010 ( .B1(n17937), .B2(n17994), .A(n17936), .ZN(n17939) );
  OAI211_X1 U21011 ( .C1(n17940), .C2(n17946), .A(n17939), .B(n17938), .ZN(
        P3_U2849) );
  NAND2_X1 U21012 ( .A1(n17941), .A2(n17974), .ZN(n17944) );
  AOI211_X1 U21013 ( .C1(n17944), .C2(n18566), .A(n17943), .B(n17942), .ZN(
        n17945) );
  AOI211_X1 U21014 ( .C1(n17946), .C2(n17951), .A(n18061), .B(n17945), .ZN(
        n17947) );
  AOI211_X1 U21015 ( .C1(n17994), .C2(n17949), .A(n17948), .B(n17947), .ZN(
        n17950) );
  OAI21_X1 U21016 ( .B1(n17951), .B2(n18062), .A(n17950), .ZN(P3_U2850) );
  AOI22_X1 U21017 ( .A1(n9820), .A2(P3_REIP_REG_11__SCAN_IN), .B1(n17994), 
        .B2(n17952), .ZN(n17963) );
  AOI21_X1 U21018 ( .B1(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n17974), .A(
        n18554), .ZN(n17957) );
  AOI22_X1 U21019 ( .A1(n18052), .A2(n17954), .B1(n17953), .B2(n17576), .ZN(
        n17956) );
  NAND3_X1 U21020 ( .A1(n17956), .A2(n18062), .A3(n17955), .ZN(n17978) );
  AOI211_X1 U21021 ( .C1(n17959), .C2(n17958), .A(n17957), .B(n17978), .ZN(
        n17966) );
  OAI211_X1 U21022 ( .C1(n18554), .C2(P3_INSTADDRPOINTER_REG_10__SCAN_IN), .A(
        n17960), .B(n17966), .ZN(n17961) );
  NAND3_X1 U21023 ( .A1(P3_INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n18074), .A3(
        n17961), .ZN(n17962) );
  OAI211_X1 U21024 ( .C1(n17965), .C2(n17964), .A(n17963), .B(n17962), .ZN(
        P3_U2851) );
  OAI21_X1 U21025 ( .B1(n17967), .B2(P3_INSTADDRPOINTER_REG_9__SCAN_IN), .A(
        n17966), .ZN(n17968) );
  OAI21_X1 U21026 ( .B1(n17969), .B2(n17968), .A(
        P3_INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n17973) );
  AOI22_X1 U21027 ( .A1(n17994), .A2(n17971), .B1(n17980), .B2(n17970), .ZN(
        n17972) );
  OAI221_X1 U21028 ( .B1(n9820), .B2(n17973), .C1(n18074), .C2(n18641), .A(
        n17972), .ZN(P3_U2852) );
  INV_X1 U21029 ( .A(n17992), .ZN(n17987) );
  AOI221_X1 U21030 ( .B1(n18554), .B2(n18568), .C1(n18554), .C2(
        P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A(n17974), .ZN(n17975) );
  AOI221_X1 U21031 ( .B1(n18549), .B2(n17987), .C1(n18549), .C2(n17985), .A(
        n17975), .ZN(n17976) );
  INV_X1 U21032 ( .A(n17976), .ZN(n17977) );
  OAI21_X1 U21033 ( .B1(n17978), .B2(n17977), .A(
        P3_INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n17983) );
  AOI22_X1 U21034 ( .A1(n17994), .A2(n17981), .B1(n17980), .B2(n17979), .ZN(
        n17982) );
  OAI221_X1 U21035 ( .B1(n9820), .B2(n17983), .C1(n18074), .C2(n18640), .A(
        n17982), .ZN(P3_U2853) );
  NOR3_X1 U21036 ( .A1(P3_INSTADDRPOINTER_REG_8__SCAN_IN), .A2(n18035), .A3(
        n18061), .ZN(n17991) );
  INV_X1 U21037 ( .A(n17984), .ZN(n18048) );
  OAI21_X1 U21038 ( .B1(n18046), .B2(n17985), .A(n18045), .ZN(n17986) );
  OAI21_X1 U21039 ( .B1(n18048), .B2(n18561), .A(n17986), .ZN(n18010) );
  OAI21_X1 U21040 ( .B1(n17987), .B2(n18010), .A(n18068), .ZN(n18008) );
  AOI21_X1 U21041 ( .B1(n18062), .B2(n18008), .A(n17988), .ZN(n17990) );
  AOI211_X1 U21042 ( .C1(n17992), .C2(n17991), .A(n17990), .B(n17989), .ZN(
        n17998) );
  AOI22_X1 U21043 ( .A1(n17996), .A2(n17995), .B1(n17994), .B2(n17993), .ZN(
        n17997) );
  OAI211_X1 U21044 ( .C1(n18079), .C2(n17999), .A(n17998), .B(n17997), .ZN(
        P3_U2854) );
  NOR3_X1 U21045 ( .A1(n18035), .A2(n18000), .A3(n18061), .ZN(n18002) );
  NOR2_X1 U21046 ( .A1(n18074), .A2(n18636), .ZN(n18001) );
  AOI221_X1 U21047 ( .B1(n18055), .B2(P3_INSTADDRPOINTER_REG_7__SCAN_IN), .C1(
        n18002), .C2(n18009), .A(n18001), .ZN(n18007) );
  INV_X1 U21048 ( .A(n18003), .ZN(n18004) );
  AOI22_X1 U21049 ( .A1(n18066), .A2(n18005), .B1(n18037), .B2(n18004), .ZN(
        n18006) );
  OAI211_X1 U21050 ( .C1(n18009), .C2(n18008), .A(n18007), .B(n18006), .ZN(
        P3_U2855) );
  NAND2_X1 U21051 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        P3_INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n18013) );
  NOR2_X1 U21052 ( .A1(n18041), .A2(n18010), .ZN(n18034) );
  OAI21_X1 U21053 ( .B1(n18034), .B2(n18011), .A(n18062), .ZN(n18030) );
  AOI21_X1 U21054 ( .B1(n18068), .B2(n18013), .A(n18030), .ZN(n18027) );
  NOR2_X1 U21055 ( .A1(n18035), .A2(n18061), .ZN(n18012) );
  NAND2_X1 U21056 ( .A1(P3_INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n18012), .ZN(
        n18033) );
  NOR3_X1 U21057 ( .A1(P3_INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n18013), .A3(
        n18033), .ZN(n18014) );
  AOI21_X1 U21058 ( .B1(P3_REIP_REG_6__SCAN_IN), .B2(n9820), .A(n18014), .ZN(
        n18018) );
  AOI22_X1 U21059 ( .A1(n18066), .A2(n18016), .B1(n18037), .B2(n18015), .ZN(
        n18017) );
  OAI211_X1 U21060 ( .C1(n18027), .C2(n18019), .A(n18018), .B(n18017), .ZN(
        P3_U2856) );
  AOI22_X1 U21061 ( .A1(n9820), .A2(P3_REIP_REG_5__SCAN_IN), .B1(n18037), .B2(
        n18020), .ZN(n18025) );
  NOR3_X1 U21062 ( .A1(P3_INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n18021), .A3(
        n18033), .ZN(n18022) );
  AOI21_X1 U21063 ( .B1(n18023), .B2(n18066), .A(n18022), .ZN(n18024) );
  OAI211_X1 U21064 ( .C1(n18027), .C2(n18026), .A(n18025), .B(n18024), .ZN(
        P3_U2857) );
  AOI22_X1 U21065 ( .A1(n9820), .A2(P3_REIP_REG_4__SCAN_IN), .B1(n18066), .B2(
        n18028), .ZN(n18032) );
  AOI22_X1 U21066 ( .A1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .A2(n18030), .B1(
        n18037), .B2(n18029), .ZN(n18031) );
  OAI211_X1 U21067 ( .C1(P3_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n18033), .A(
        n18032), .B(n18031), .ZN(P3_U2858) );
  AOI211_X1 U21068 ( .C1(n18035), .C2(n18041), .A(n18034), .B(n18061), .ZN(
        n18043) );
  AOI22_X1 U21069 ( .A1(n18066), .A2(n18038), .B1(n18037), .B2(n18036), .ZN(
        n18040) );
  OAI211_X1 U21070 ( .C1(n18062), .C2(n18041), .A(n18040), .B(n18039), .ZN(
        n18042) );
  OR2_X1 U21071 ( .A1(n18043), .A2(n18042), .ZN(P3_U2859) );
  NOR3_X1 U21072 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18708), .A3(
        n18044), .ZN(n18051) );
  OAI211_X1 U21073 ( .C1(n18046), .C2(n18708), .A(
        P3_INSTADDRPOINTER_REG_2__SCAN_IN), .B(n18045), .ZN(n18047) );
  OAI221_X1 U21074 ( .B1(n18561), .B2(n18049), .C1(n18561), .C2(n18048), .A(
        n18047), .ZN(n18050) );
  AOI211_X1 U21075 ( .C1(n18053), .C2(n18052), .A(n18051), .B(n18050), .ZN(
        n18058) );
  AOI22_X1 U21076 ( .A1(P3_INSTADDRPOINTER_REG_2__SCAN_IN), .A2(n18055), .B1(
        n18066), .B2(n18054), .ZN(n18057) );
  NAND2_X1 U21077 ( .A1(n9820), .A2(P3_REIP_REG_2__SCAN_IN), .ZN(n18056) );
  OAI211_X1 U21078 ( .C1(n18058), .C2(n18061), .A(n18057), .B(n18056), .ZN(
        P3_U2860) );
  INV_X1 U21079 ( .A(n18059), .ZN(n18071) );
  NOR2_X1 U21080 ( .A1(n18074), .A2(n18729), .ZN(n18064) );
  OR3_X1 U21081 ( .A1(n18061), .A2(P3_INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        n18060), .ZN(n18072) );
  AOI21_X1 U21082 ( .B1(n18062), .B2(n18072), .A(n18708), .ZN(n18063) );
  AOI211_X1 U21083 ( .C1(n18066), .C2(n18065), .A(n18064), .B(n18063), .ZN(
        n18070) );
  NAND3_X1 U21084 ( .A1(n18068), .A2(n18708), .A3(n18067), .ZN(n18069) );
  OAI211_X1 U21085 ( .C1(n18071), .C2(n18079), .A(n18070), .B(n18069), .ZN(
        P3_U2861) );
  OAI221_X1 U21086 ( .B1(n18724), .B2(n18568), .C1(n18724), .C2(n18073), .A(
        n18072), .ZN(n18075) );
  AOI22_X1 U21087 ( .A1(n9820), .A2(P3_REIP_REG_0__SCAN_IN), .B1(n18075), .B2(
        n18074), .ZN(n18076) );
  OAI221_X1 U21088 ( .B1(n18080), .B2(n18079), .C1(n18078), .C2(n18077), .A(
        n18076), .ZN(P3_U2862) );
  AOI211_X1 U21089 ( .C1(n18082), .C2(n18081), .A(n18603), .B(n18706), .ZN(
        n18590) );
  OAI21_X1 U21090 ( .B1(n18590), .B2(n18140), .A(n18087), .ZN(n18083) );
  OAI221_X1 U21091 ( .B1(n18088), .B2(n18740), .C1(n18088), .C2(n18087), .A(
        n18083), .ZN(P3_U2863) );
  INV_X1 U21092 ( .A(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18579) );
  NAND2_X1 U21093 ( .A1(n18579), .A2(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(
        n18277) );
  INV_X1 U21094 ( .A(n18277), .ZN(n18278) );
  NAND2_X1 U21095 ( .A1(n18576), .A2(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n18371) );
  NOR2_X1 U21096 ( .A1(n18444), .A2(n18371), .ZN(n18397) );
  NOR2_X1 U21097 ( .A1(n18278), .A2(n18397), .ZN(n18085) );
  OAI22_X1 U21098 ( .A1(n18086), .A2(n18579), .B1(n18085), .B2(n18084), .ZN(
        P3_U2866) );
  NOR2_X1 U21099 ( .A1(n18580), .A2(n18087), .ZN(P3_U2867) );
  NAND2_X1 U21100 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n18571) );
  NOR2_X1 U21101 ( .A1(n18576), .A2(n18579), .ZN(n18421) );
  INV_X1 U21102 ( .A(n18421), .ZN(n18090) );
  NOR2_X2 U21103 ( .A1(n18571), .A2(n18090), .ZN(n18469) );
  NAND2_X1 U21104 ( .A1(n20944), .A2(n18088), .ZN(n18572) );
  NOR2_X1 U21105 ( .A1(P3_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n18189) );
  INV_X1 U21106 ( .A(n18189), .ZN(n18233) );
  NOR2_X1 U21107 ( .A1(n18572), .A2(n18233), .ZN(n18196) );
  NOR2_X1 U21108 ( .A1(n18469), .A2(n18206), .ZN(n18167) );
  INV_X1 U21109 ( .A(n18394), .ZN(n18447) );
  OAI21_X1 U21110 ( .B1(n18696), .B2(n18088), .A(n18447), .ZN(n18089) );
  NOR2_X1 U21111 ( .A1(n20944), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18345) );
  NOR2_X1 U21112 ( .A1(n18088), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18322) );
  OR2_X1 U21113 ( .A1(n18345), .A2(n18322), .ZN(n18396) );
  NAND2_X1 U21114 ( .A1(n18421), .A2(n18396), .ZN(n18443) );
  OAI22_X1 U21115 ( .A1(n18167), .A2(n18089), .B1(n18348), .B2(n18443), .ZN(
        n18137) );
  NOR2_X1 U21116 ( .A1(n18090), .A2(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n18475) );
  NAND2_X1 U21117 ( .A1(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n18475), .ZN(
        n18442) );
  INV_X1 U21118 ( .A(n18442), .ZN(n18522) );
  AND2_X1 U21119 ( .A1(BUF2_REG_24__SCAN_IN), .A2(n18476), .ZN(n18472) );
  NOR2_X2 U21120 ( .A1(n18394), .A2(n18091), .ZN(n18471) );
  NOR2_X1 U21121 ( .A1(n9805), .A2(n18167), .ZN(n18132) );
  AOI22_X1 U21122 ( .A1(n18522), .A2(n18472), .B1(n18471), .B2(n18132), .ZN(
        n18097) );
  NAND2_X1 U21123 ( .A1(n18093), .A2(n18092), .ZN(n18133) );
  NOR2_X1 U21124 ( .A1(n18094), .A2(n18133), .ZN(n18139) );
  INV_X1 U21125 ( .A(BUF2_REG_16__SCAN_IN), .ZN(n18095) );
  NOR2_X2 U21126 ( .A1(n18348), .A2(n18095), .ZN(n18477) );
  NAND2_X1 U21127 ( .A1(n18421), .A2(n18345), .ZN(n18468) );
  INV_X1 U21128 ( .A(n18468), .ZN(n18448) );
  AOI22_X1 U21129 ( .A1(n18206), .A2(n18139), .B1(n18477), .B2(n18448), .ZN(
        n18096) );
  OAI211_X1 U21130 ( .C1(n18098), .C2(n18137), .A(n18097), .B(n18096), .ZN(
        P3_U2868) );
  INV_X1 U21131 ( .A(P3_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n18104) );
  AND2_X1 U21132 ( .A1(n18476), .A2(BUF2_REG_17__SCAN_IN), .ZN(n18483) );
  NOR2_X2 U21133 ( .A1(n18394), .A2(n18099), .ZN(n18481) );
  AOI22_X1 U21134 ( .A1(n18448), .A2(n18483), .B1(n18132), .B2(n18481), .ZN(
        n18103) );
  NOR2_X1 U21135 ( .A1(n18100), .A2(n18133), .ZN(n18143) );
  NOR2_X2 U21136 ( .A1(n18101), .A2(n18348), .ZN(n18482) );
  AOI22_X1 U21137 ( .A1(n18206), .A2(n18143), .B1(n18522), .B2(n18482), .ZN(
        n18102) );
  OAI211_X1 U21138 ( .C1(n18104), .C2(n18137), .A(n18103), .B(n18102), .ZN(
        P3_U2869) );
  AND2_X1 U21139 ( .A1(n18476), .A2(BUF2_REG_18__SCAN_IN), .ZN(n18489) );
  NOR2_X2 U21140 ( .A1(n18394), .A2(n18105), .ZN(n18487) );
  AOI22_X1 U21141 ( .A1(n18448), .A2(n18489), .B1(n18132), .B2(n18487), .ZN(
        n18109) );
  NOR2_X1 U21142 ( .A1(n18106), .A2(n18133), .ZN(n18146) );
  INV_X1 U21143 ( .A(BUF2_REG_26__SCAN_IN), .ZN(n18107) );
  NOR2_X2 U21144 ( .A1(n18107), .A2(n18348), .ZN(n18488) );
  AOI22_X1 U21145 ( .A1(n18196), .A2(n18146), .B1(n18522), .B2(n18488), .ZN(
        n18108) );
  OAI211_X1 U21146 ( .C1(n18110), .C2(n18137), .A(n18109), .B(n18108), .ZN(
        P3_U2870) );
  AND2_X1 U21147 ( .A1(BUF2_REG_27__SCAN_IN), .A2(n18476), .ZN(n18494) );
  NOR2_X2 U21148 ( .A1(n18394), .A2(n18111), .ZN(n18493) );
  AOI22_X1 U21149 ( .A1(n18522), .A2(n18494), .B1(n18132), .B2(n18493), .ZN(
        n18114) );
  NOR2_X1 U21150 ( .A1(n18112), .A2(n18133), .ZN(n18149) );
  NOR2_X2 U21151 ( .A1(n18348), .A2(n15087), .ZN(n18495) );
  AOI22_X1 U21152 ( .A1(n18196), .A2(n18149), .B1(n18448), .B2(n18495), .ZN(
        n18113) );
  OAI211_X1 U21153 ( .C1(n18115), .C2(n18137), .A(n18114), .B(n18113), .ZN(
        P3_U2871) );
  AND2_X1 U21154 ( .A1(BUF2_REG_20__SCAN_IN), .A2(n18476), .ZN(n18501) );
  NOR2_X2 U21155 ( .A1(n18116), .A2(n18394), .ZN(n18499) );
  AOI22_X1 U21156 ( .A1(n18448), .A2(n18501), .B1(n18132), .B2(n18499), .ZN(
        n18120) );
  NOR2_X1 U21157 ( .A1(n18117), .A2(n18133), .ZN(n18152) );
  NOR2_X2 U21158 ( .A1(n18118), .A2(n18348), .ZN(n18500) );
  AOI22_X1 U21159 ( .A1(n18196), .A2(n18152), .B1(n18522), .B2(n18500), .ZN(
        n18119) );
  OAI211_X1 U21160 ( .C1(n18121), .C2(n18137), .A(n18120), .B(n18119), .ZN(
        P3_U2872) );
  NOR2_X2 U21161 ( .A1(n15075), .A2(n18348), .ZN(n18506) );
  NOR2_X2 U21162 ( .A1(n18122), .A2(n18394), .ZN(n18505) );
  AOI22_X1 U21163 ( .A1(n18448), .A2(n18506), .B1(n18132), .B2(n18505), .ZN(
        n18125) );
  NOR2_X1 U21164 ( .A1(n18123), .A2(n18133), .ZN(n18155) );
  NOR2_X2 U21165 ( .A1(n20974), .A2(n18348), .ZN(n18507) );
  AOI22_X1 U21166 ( .A1(n18206), .A2(n18155), .B1(n18522), .B2(n18507), .ZN(
        n18124) );
  OAI211_X1 U21167 ( .C1(n18126), .C2(n18137), .A(n18125), .B(n18124), .ZN(
        P3_U2873) );
  AND2_X1 U21168 ( .A1(BUF2_REG_30__SCAN_IN), .A2(n18476), .ZN(n18512) );
  NOR2_X2 U21169 ( .A1(n18127), .A2(n18394), .ZN(n18511) );
  AOI22_X1 U21170 ( .A1(n18522), .A2(n18512), .B1(n18132), .B2(n18511), .ZN(
        n18130) );
  NOR2_X1 U21171 ( .A1(n18128), .A2(n18133), .ZN(n18158) );
  INV_X1 U21172 ( .A(BUF2_REG_22__SCAN_IN), .ZN(n20905) );
  NOR2_X2 U21173 ( .A1(n20905), .A2(n18348), .ZN(n18513) );
  AOI22_X1 U21174 ( .A1(n18196), .A2(n18158), .B1(n18448), .B2(n18513), .ZN(
        n18129) );
  OAI211_X1 U21175 ( .C1(n18131), .C2(n18137), .A(n18130), .B(n18129), .ZN(
        P3_U2874) );
  INV_X1 U21176 ( .A(P3_INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n18138) );
  NOR2_X2 U21177 ( .A1(n15069), .A2(n18348), .ZN(n18521) );
  AND2_X1 U21178 ( .A1(BUF2_REG_7__SCAN_IN), .A2(n18447), .ZN(n18518) );
  AOI22_X1 U21179 ( .A1(n18448), .A2(n18521), .B1(n18132), .B2(n18518), .ZN(
        n18136) );
  NOR2_X1 U21180 ( .A1(n18134), .A2(n18133), .ZN(n18161) );
  NOR2_X2 U21181 ( .A1(n19145), .A2(n18348), .ZN(n18520) );
  AOI22_X1 U21182 ( .A1(n18206), .A2(n18161), .B1(n18522), .B2(n18520), .ZN(
        n18135) );
  OAI211_X1 U21183 ( .C1(n18138), .C2(n18137), .A(n18136), .B(n18135), .ZN(
        P3_U2875) );
  NAND2_X1 U21184 ( .A1(n18322), .A2(n18189), .ZN(n18166) );
  AOI22_X1 U21185 ( .A1(n18448), .A2(n18472), .B1(n18471), .B2(n18162), .ZN(
        n18142) );
  NOR2_X1 U21186 ( .A1(n18579), .A2(n18323), .ZN(n18473) );
  NOR2_X1 U21187 ( .A1(n18394), .A2(n18140), .ZN(n18474) );
  INV_X1 U21188 ( .A(n18474), .ZN(n18188) );
  NOR2_X1 U21189 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18188), .ZN(
        n18420) );
  AOI22_X1 U21190 ( .A1(n18476), .A2(n18473), .B1(n18189), .B2(n18420), .ZN(
        n18163) );
  AOI22_X1 U21191 ( .A1(P3_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n18163), .B1(
        n18469), .B2(n18477), .ZN(n18141) );
  OAI211_X1 U21192 ( .C1(n18480), .C2(n18166), .A(n18142), .B(n18141), .ZN(
        P3_U2876) );
  INV_X1 U21193 ( .A(n18143), .ZN(n18486) );
  AOI22_X1 U21194 ( .A1(n18448), .A2(n18482), .B1(n18481), .B2(n18162), .ZN(
        n18145) );
  AOI22_X1 U21195 ( .A1(P3_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n18163), .B1(
        n18469), .B2(n18483), .ZN(n18144) );
  OAI211_X1 U21196 ( .C1(n18486), .C2(n18166), .A(n18145), .B(n18144), .ZN(
        P3_U2877) );
  INV_X1 U21197 ( .A(n18146), .ZN(n18492) );
  AOI22_X1 U21198 ( .A1(n18469), .A2(n18489), .B1(n18487), .B2(n18162), .ZN(
        n18148) );
  AOI22_X1 U21199 ( .A1(P3_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n18163), .B1(
        n18448), .B2(n18488), .ZN(n18147) );
  OAI211_X1 U21200 ( .C1(n18492), .C2(n18166), .A(n18148), .B(n18147), .ZN(
        P3_U2878) );
  INV_X1 U21201 ( .A(n18149), .ZN(n18498) );
  AOI22_X1 U21202 ( .A1(n18448), .A2(n18494), .B1(n18493), .B2(n18162), .ZN(
        n18151) );
  AOI22_X1 U21203 ( .A1(P3_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n18163), .B1(
        n18469), .B2(n18495), .ZN(n18150) );
  OAI211_X1 U21204 ( .C1(n18498), .C2(n18166), .A(n18151), .B(n18150), .ZN(
        P3_U2879) );
  INV_X1 U21205 ( .A(n18152), .ZN(n18504) );
  AOI22_X1 U21206 ( .A1(n18448), .A2(n18500), .B1(n18499), .B2(n18162), .ZN(
        n18154) );
  AOI22_X1 U21207 ( .A1(P3_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n18163), .B1(
        n18469), .B2(n18501), .ZN(n18153) );
  OAI211_X1 U21208 ( .C1(n18504), .C2(n18166), .A(n18154), .B(n18153), .ZN(
        P3_U2880) );
  AOI22_X1 U21209 ( .A1(n18469), .A2(n18506), .B1(n18505), .B2(n18162), .ZN(
        n18157) );
  AOI22_X1 U21210 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n18163), .B1(
        n18448), .B2(n18507), .ZN(n18156) );
  OAI211_X1 U21211 ( .C1(n18510), .C2(n18166), .A(n18157), .B(n18156), .ZN(
        P3_U2881) );
  INV_X1 U21212 ( .A(n18158), .ZN(n18516) );
  AOI22_X1 U21213 ( .A1(n18469), .A2(n18513), .B1(n18511), .B2(n18162), .ZN(
        n18160) );
  AOI22_X1 U21214 ( .A1(P3_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n18163), .B1(
        n18448), .B2(n18512), .ZN(n18159) );
  OAI211_X1 U21215 ( .C1(n18516), .C2(n18166), .A(n18160), .B(n18159), .ZN(
        P3_U2882) );
  INV_X1 U21216 ( .A(n18161), .ZN(n18526) );
  AOI22_X1 U21217 ( .A1(n18469), .A2(n18521), .B1(n18518), .B2(n18162), .ZN(
        n18165) );
  AOI22_X1 U21218 ( .A1(P3_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n18163), .B1(
        n18448), .B2(n18520), .ZN(n18164) );
  OAI211_X1 U21219 ( .C1(n18526), .C2(n18166), .A(n18165), .B(n18164), .ZN(
        P3_U2883) );
  NAND2_X1 U21220 ( .A1(n18345), .A2(n18189), .ZN(n18187) );
  INV_X1 U21221 ( .A(n18166), .ZN(n18228) );
  INV_X1 U21222 ( .A(n18187), .ZN(n18250) );
  NOR2_X1 U21223 ( .A1(n18228), .A2(n18250), .ZN(n18211) );
  NOR2_X1 U21224 ( .A1(n9805), .A2(n18211), .ZN(n18183) );
  AOI22_X1 U21225 ( .A1(n18469), .A2(n18472), .B1(n18471), .B2(n18183), .ZN(
        n18170) );
  OAI22_X1 U21226 ( .A1(n18167), .A2(n18348), .B1(n18211), .B2(n18394), .ZN(
        n18168) );
  OAI21_X1 U21227 ( .B1(n18250), .B2(n18696), .A(n18168), .ZN(n18184) );
  AOI22_X1 U21228 ( .A1(P3_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n18184), .B1(
        n18196), .B2(n18477), .ZN(n18169) );
  OAI211_X1 U21229 ( .C1(n18480), .C2(n18187), .A(n18170), .B(n18169), .ZN(
        P3_U2884) );
  AOI22_X1 U21230 ( .A1(n18469), .A2(n18482), .B1(n18481), .B2(n18183), .ZN(
        n18172) );
  AOI22_X1 U21231 ( .A1(P3_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n18184), .B1(
        n18196), .B2(n18483), .ZN(n18171) );
  OAI211_X1 U21232 ( .C1(n18486), .C2(n18187), .A(n18172), .B(n18171), .ZN(
        P3_U2885) );
  AOI22_X1 U21233 ( .A1(n18206), .A2(n18489), .B1(n18487), .B2(n18183), .ZN(
        n18174) );
  AOI22_X1 U21234 ( .A1(P3_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n18184), .B1(
        n18469), .B2(n18488), .ZN(n18173) );
  OAI211_X1 U21235 ( .C1(n18492), .C2(n18187), .A(n18174), .B(n18173), .ZN(
        P3_U2886) );
  AOI22_X1 U21236 ( .A1(n18469), .A2(n18494), .B1(n18493), .B2(n18183), .ZN(
        n18176) );
  AOI22_X1 U21237 ( .A1(P3_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n18184), .B1(
        n18196), .B2(n18495), .ZN(n18175) );
  OAI211_X1 U21238 ( .C1(n18498), .C2(n18187), .A(n18176), .B(n18175), .ZN(
        P3_U2887) );
  AOI22_X1 U21239 ( .A1(n18206), .A2(n18501), .B1(n18499), .B2(n18183), .ZN(
        n18178) );
  AOI22_X1 U21240 ( .A1(P3_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n18184), .B1(
        n18469), .B2(n18500), .ZN(n18177) );
  OAI211_X1 U21241 ( .C1(n18504), .C2(n18187), .A(n18178), .B(n18177), .ZN(
        P3_U2888) );
  AOI22_X1 U21242 ( .A1(n18469), .A2(n18507), .B1(n18505), .B2(n18183), .ZN(
        n18180) );
  AOI22_X1 U21243 ( .A1(P3_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n18184), .B1(
        n18196), .B2(n18506), .ZN(n18179) );
  OAI211_X1 U21244 ( .C1(n18510), .C2(n18187), .A(n18180), .B(n18179), .ZN(
        P3_U2889) );
  AOI22_X1 U21245 ( .A1(n18206), .A2(n18513), .B1(n18511), .B2(n18183), .ZN(
        n18182) );
  AOI22_X1 U21246 ( .A1(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n18184), .B1(
        n18469), .B2(n18512), .ZN(n18181) );
  OAI211_X1 U21247 ( .C1(n18516), .C2(n18187), .A(n18182), .B(n18181), .ZN(
        P3_U2890) );
  AOI22_X1 U21248 ( .A1(n18206), .A2(n18521), .B1(n18518), .B2(n18183), .ZN(
        n18186) );
  AOI22_X1 U21249 ( .A1(P3_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n18184), .B1(
        n18469), .B2(n18520), .ZN(n18185) );
  OAI211_X1 U21250 ( .C1(n18526), .C2(n18187), .A(n18186), .B(n18185), .ZN(
        P3_U2891) );
  NOR2_X2 U21251 ( .A1(n18571), .A2(n18233), .ZN(n18272) );
  INV_X1 U21252 ( .A(n18272), .ZN(n18210) );
  AOI22_X1 U21253 ( .A1(n18477), .A2(n18228), .B1(n18471), .B2(n18205), .ZN(
        n18191) );
  AOI21_X1 U21254 ( .B1(n20944), .B2(n18444), .A(n18188), .ZN(n18279) );
  NAND2_X1 U21255 ( .A1(n18189), .A2(n18279), .ZN(n18207) );
  AOI22_X1 U21256 ( .A1(P3_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n18207), .B1(
        n18206), .B2(n18472), .ZN(n18190) );
  OAI211_X1 U21257 ( .C1(n18480), .C2(n18210), .A(n18191), .B(n18190), .ZN(
        P3_U2892) );
  AOI22_X1 U21258 ( .A1(n18206), .A2(n18482), .B1(n18481), .B2(n18205), .ZN(
        n18193) );
  AOI22_X1 U21259 ( .A1(P3_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n18207), .B1(
        n18483), .B2(n18228), .ZN(n18192) );
  OAI211_X1 U21260 ( .C1(n18486), .C2(n18210), .A(n18193), .B(n18192), .ZN(
        P3_U2893) );
  AOI22_X1 U21261 ( .A1(n18206), .A2(n18488), .B1(n18487), .B2(n18205), .ZN(
        n18195) );
  AOI22_X1 U21262 ( .A1(P3_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n18207), .B1(
        n18489), .B2(n18228), .ZN(n18194) );
  OAI211_X1 U21263 ( .C1(n18492), .C2(n18210), .A(n18195), .B(n18194), .ZN(
        P3_U2894) );
  AOI22_X1 U21264 ( .A1(n18495), .A2(n18228), .B1(n18493), .B2(n18205), .ZN(
        n18198) );
  AOI22_X1 U21265 ( .A1(P3_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n18207), .B1(
        n18196), .B2(n18494), .ZN(n18197) );
  OAI211_X1 U21266 ( .C1(n18498), .C2(n18210), .A(n18198), .B(n18197), .ZN(
        P3_U2895) );
  AOI22_X1 U21267 ( .A1(n18206), .A2(n18500), .B1(n18499), .B2(n18205), .ZN(
        n18200) );
  AOI22_X1 U21268 ( .A1(P3_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n18207), .B1(
        n18501), .B2(n18228), .ZN(n18199) );
  OAI211_X1 U21269 ( .C1(n18504), .C2(n18210), .A(n18200), .B(n18199), .ZN(
        P3_U2896) );
  AOI22_X1 U21270 ( .A1(n18506), .A2(n18228), .B1(n18505), .B2(n18205), .ZN(
        n18202) );
  AOI22_X1 U21271 ( .A1(P3_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n18207), .B1(
        n18206), .B2(n18507), .ZN(n18201) );
  OAI211_X1 U21272 ( .C1(n18510), .C2(n18210), .A(n18202), .B(n18201), .ZN(
        P3_U2897) );
  AOI22_X1 U21273 ( .A1(n18513), .A2(n18228), .B1(n18511), .B2(n18205), .ZN(
        n18204) );
  AOI22_X1 U21274 ( .A1(P3_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n18207), .B1(
        n18206), .B2(n18512), .ZN(n18203) );
  OAI211_X1 U21275 ( .C1(n18516), .C2(n18210), .A(n18204), .B(n18203), .ZN(
        P3_U2898) );
  AOI22_X1 U21276 ( .A1(n18521), .A2(n18228), .B1(n18518), .B2(n18205), .ZN(
        n18209) );
  AOI22_X1 U21277 ( .A1(P3_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n18207), .B1(
        n18206), .B2(n18520), .ZN(n18208) );
  OAI211_X1 U21278 ( .C1(n18526), .C2(n18210), .A(n18209), .B(n18208), .ZN(
        P3_U2899) );
  NOR2_X2 U21279 ( .A1(n18572), .A2(n18277), .ZN(n18295) );
  INV_X1 U21280 ( .A(n18295), .ZN(n18232) );
  NOR2_X1 U21281 ( .A1(n18272), .A2(n18295), .ZN(n18255) );
  NOR2_X1 U21282 ( .A1(n9805), .A2(n18255), .ZN(n18227) );
  AOI22_X1 U21283 ( .A1(n18472), .A2(n18228), .B1(n18471), .B2(n18227), .ZN(
        n18214) );
  OAI22_X1 U21284 ( .A1(n18211), .A2(n18348), .B1(n18255), .B2(n18394), .ZN(
        n18212) );
  OAI21_X1 U21285 ( .B1(n18295), .B2(n18696), .A(n18212), .ZN(n18229) );
  AOI22_X1 U21286 ( .A1(P3_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n18229), .B1(
        n18477), .B2(n18250), .ZN(n18213) );
  OAI211_X1 U21287 ( .C1(n18480), .C2(n18232), .A(n18214), .B(n18213), .ZN(
        P3_U2900) );
  AOI22_X1 U21288 ( .A1(n18482), .A2(n18228), .B1(n18481), .B2(n18227), .ZN(
        n18216) );
  AOI22_X1 U21289 ( .A1(P3_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n18229), .B1(
        n18483), .B2(n18250), .ZN(n18215) );
  OAI211_X1 U21290 ( .C1(n18486), .C2(n18232), .A(n18216), .B(n18215), .ZN(
        P3_U2901) );
  AOI22_X1 U21291 ( .A1(n18489), .A2(n18250), .B1(n18487), .B2(n18227), .ZN(
        n18218) );
  AOI22_X1 U21292 ( .A1(P3_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n18229), .B1(
        n18488), .B2(n18228), .ZN(n18217) );
  OAI211_X1 U21293 ( .C1(n18492), .C2(n18232), .A(n18218), .B(n18217), .ZN(
        P3_U2902) );
  AOI22_X1 U21294 ( .A1(n18495), .A2(n18250), .B1(n18493), .B2(n18227), .ZN(
        n18220) );
  AOI22_X1 U21295 ( .A1(P3_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n18229), .B1(
        n18494), .B2(n18228), .ZN(n18219) );
  OAI211_X1 U21296 ( .C1(n18498), .C2(n18232), .A(n18220), .B(n18219), .ZN(
        P3_U2903) );
  AOI22_X1 U21297 ( .A1(n18500), .A2(n18228), .B1(n18499), .B2(n18227), .ZN(
        n18222) );
  AOI22_X1 U21298 ( .A1(P3_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n18229), .B1(
        n18501), .B2(n18250), .ZN(n18221) );
  OAI211_X1 U21299 ( .C1(n18504), .C2(n18232), .A(n18222), .B(n18221), .ZN(
        P3_U2904) );
  AOI22_X1 U21300 ( .A1(n18506), .A2(n18250), .B1(n18505), .B2(n18227), .ZN(
        n18224) );
  AOI22_X1 U21301 ( .A1(P3_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n18229), .B1(
        n18507), .B2(n18228), .ZN(n18223) );
  OAI211_X1 U21302 ( .C1(n18510), .C2(n18232), .A(n18224), .B(n18223), .ZN(
        P3_U2905) );
  AOI22_X1 U21303 ( .A1(n18512), .A2(n18228), .B1(n18511), .B2(n18227), .ZN(
        n18226) );
  AOI22_X1 U21304 ( .A1(P3_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n18229), .B1(
        n18513), .B2(n18250), .ZN(n18225) );
  OAI211_X1 U21305 ( .C1(n18516), .C2(n18232), .A(n18226), .B(n18225), .ZN(
        P3_U2906) );
  AOI22_X1 U21306 ( .A1(n18521), .A2(n18250), .B1(n18518), .B2(n18227), .ZN(
        n18231) );
  AOI22_X1 U21307 ( .A1(P3_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n18229), .B1(
        n18520), .B2(n18228), .ZN(n18230) );
  OAI211_X1 U21308 ( .C1(n18526), .C2(n18232), .A(n18231), .B(n18230), .ZN(
        P3_U2907) );
  NAND2_X1 U21309 ( .A1(n18322), .A2(n18278), .ZN(n18254) );
  AOI22_X1 U21310 ( .A1(n18472), .A2(n18250), .B1(n18471), .B2(n18249), .ZN(
        n18236) );
  NOR2_X1 U21311 ( .A1(n20944), .A2(n18233), .ZN(n18234) );
  AOI22_X1 U21312 ( .A1(n18476), .A2(n18234), .B1(n18420), .B2(n18278), .ZN(
        n18251) );
  AOI22_X1 U21313 ( .A1(P3_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n18251), .B1(
        n18477), .B2(n18272), .ZN(n18235) );
  OAI211_X1 U21314 ( .C1(n18480), .C2(n18254), .A(n18236), .B(n18235), .ZN(
        P3_U2908) );
  AOI22_X1 U21315 ( .A1(n18482), .A2(n18250), .B1(n18481), .B2(n18249), .ZN(
        n18238) );
  AOI22_X1 U21316 ( .A1(P3_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n18251), .B1(
        n18483), .B2(n18272), .ZN(n18237) );
  OAI211_X1 U21317 ( .C1(n18486), .C2(n18254), .A(n18238), .B(n18237), .ZN(
        P3_U2909) );
  AOI22_X1 U21318 ( .A1(n18488), .A2(n18250), .B1(n18487), .B2(n18249), .ZN(
        n18240) );
  AOI22_X1 U21319 ( .A1(P3_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n18251), .B1(
        n18489), .B2(n18272), .ZN(n18239) );
  OAI211_X1 U21320 ( .C1(n18492), .C2(n18254), .A(n18240), .B(n18239), .ZN(
        P3_U2910) );
  AOI22_X1 U21321 ( .A1(n18494), .A2(n18250), .B1(n18493), .B2(n18249), .ZN(
        n18242) );
  AOI22_X1 U21322 ( .A1(P3_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n18251), .B1(
        n18495), .B2(n18272), .ZN(n18241) );
  OAI211_X1 U21323 ( .C1(n18498), .C2(n18254), .A(n18242), .B(n18241), .ZN(
        P3_U2911) );
  AOI22_X1 U21324 ( .A1(n18500), .A2(n18250), .B1(n18499), .B2(n18249), .ZN(
        n18244) );
  AOI22_X1 U21325 ( .A1(P3_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n18251), .B1(
        n18501), .B2(n18272), .ZN(n18243) );
  OAI211_X1 U21326 ( .C1(n18504), .C2(n18254), .A(n18244), .B(n18243), .ZN(
        P3_U2912) );
  AOI22_X1 U21327 ( .A1(n18506), .A2(n18272), .B1(n18505), .B2(n18249), .ZN(
        n18246) );
  AOI22_X1 U21328 ( .A1(P3_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n18251), .B1(
        n18507), .B2(n18250), .ZN(n18245) );
  OAI211_X1 U21329 ( .C1(n18510), .C2(n18254), .A(n18246), .B(n18245), .ZN(
        P3_U2913) );
  AOI22_X1 U21330 ( .A1(n18513), .A2(n18272), .B1(n18511), .B2(n18249), .ZN(
        n18248) );
  AOI22_X1 U21331 ( .A1(P3_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n18251), .B1(
        n18512), .B2(n18250), .ZN(n18247) );
  OAI211_X1 U21332 ( .C1(n18516), .C2(n18254), .A(n18248), .B(n18247), .ZN(
        P3_U2914) );
  AOI22_X1 U21333 ( .A1(n18521), .A2(n18272), .B1(n18518), .B2(n18249), .ZN(
        n18253) );
  AOI22_X1 U21334 ( .A1(P3_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n18251), .B1(
        n18520), .B2(n18250), .ZN(n18252) );
  OAI211_X1 U21335 ( .C1(n18526), .C2(n18254), .A(n18253), .B(n18252), .ZN(
        P3_U2915) );
  NAND2_X1 U21336 ( .A1(n18345), .A2(n18278), .ZN(n18276) );
  INV_X1 U21337 ( .A(n18254), .ZN(n18317) );
  INV_X1 U21338 ( .A(n18276), .ZN(n18341) );
  NOR2_X1 U21339 ( .A1(n18317), .A2(n18341), .ZN(n18300) );
  NOR2_X1 U21340 ( .A1(n9805), .A2(n18300), .ZN(n18271) );
  AOI22_X1 U21341 ( .A1(n18477), .A2(n18295), .B1(n18471), .B2(n18271), .ZN(
        n18258) );
  OAI21_X1 U21342 ( .B1(n18255), .B2(n18444), .A(n18300), .ZN(n18256) );
  OAI211_X1 U21343 ( .C1(n18341), .C2(n18696), .A(n18447), .B(n18256), .ZN(
        n18273) );
  AOI22_X1 U21344 ( .A1(P3_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n18273), .B1(
        n18472), .B2(n18272), .ZN(n18257) );
  OAI211_X1 U21345 ( .C1(n18480), .C2(n18276), .A(n18258), .B(n18257), .ZN(
        P3_U2916) );
  AOI22_X1 U21346 ( .A1(P3_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n18273), .B1(
        n18481), .B2(n18271), .ZN(n18260) );
  AOI22_X1 U21347 ( .A1(n18482), .A2(n18272), .B1(n18483), .B2(n18295), .ZN(
        n18259) );
  OAI211_X1 U21348 ( .C1(n18486), .C2(n18276), .A(n18260), .B(n18259), .ZN(
        P3_U2917) );
  AOI22_X1 U21349 ( .A1(P3_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n18273), .B1(
        n18487), .B2(n18271), .ZN(n18262) );
  AOI22_X1 U21350 ( .A1(n18488), .A2(n18272), .B1(n18489), .B2(n18295), .ZN(
        n18261) );
  OAI211_X1 U21351 ( .C1(n18492), .C2(n18276), .A(n18262), .B(n18261), .ZN(
        P3_U2918) );
  AOI22_X1 U21352 ( .A1(n18494), .A2(n18272), .B1(n18493), .B2(n18271), .ZN(
        n18264) );
  AOI22_X1 U21353 ( .A1(P3_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n18273), .B1(
        n18495), .B2(n18295), .ZN(n18263) );
  OAI211_X1 U21354 ( .C1(n18498), .C2(n18276), .A(n18264), .B(n18263), .ZN(
        P3_U2919) );
  AOI22_X1 U21355 ( .A1(P3_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n18273), .B1(
        n18499), .B2(n18271), .ZN(n18266) );
  AOI22_X1 U21356 ( .A1(n18500), .A2(n18272), .B1(n18501), .B2(n18295), .ZN(
        n18265) );
  OAI211_X1 U21357 ( .C1(n18504), .C2(n18276), .A(n18266), .B(n18265), .ZN(
        P3_U2920) );
  AOI22_X1 U21358 ( .A1(n18506), .A2(n18295), .B1(n18505), .B2(n18271), .ZN(
        n18268) );
  AOI22_X1 U21359 ( .A1(P3_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n18273), .B1(
        n18507), .B2(n18272), .ZN(n18267) );
  OAI211_X1 U21360 ( .C1(n18510), .C2(n18276), .A(n18268), .B(n18267), .ZN(
        P3_U2921) );
  AOI22_X1 U21361 ( .A1(P3_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n18273), .B1(
        n18511), .B2(n18271), .ZN(n18270) );
  AOI22_X1 U21362 ( .A1(n18513), .A2(n18295), .B1(n18512), .B2(n18272), .ZN(
        n18269) );
  OAI211_X1 U21363 ( .C1(n18516), .C2(n18276), .A(n18270), .B(n18269), .ZN(
        P3_U2922) );
  AOI22_X1 U21364 ( .A1(n18521), .A2(n18295), .B1(n18518), .B2(n18271), .ZN(
        n18275) );
  AOI22_X1 U21365 ( .A1(P3_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n18273), .B1(
        n18520), .B2(n18272), .ZN(n18274) );
  OAI211_X1 U21366 ( .C1(n18526), .C2(n18276), .A(n18275), .B(n18274), .ZN(
        P3_U2923) );
  NOR2_X2 U21367 ( .A1(n18571), .A2(n18277), .ZN(n18366) );
  INV_X1 U21368 ( .A(n18366), .ZN(n18299) );
  AOI22_X1 U21369 ( .A1(n18472), .A2(n18295), .B1(n18471), .B2(n18294), .ZN(
        n18281) );
  NAND2_X1 U21370 ( .A1(n18279), .A2(n18278), .ZN(n18296) );
  AOI22_X1 U21371 ( .A1(P3_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n18296), .B1(
        n18477), .B2(n18317), .ZN(n18280) );
  OAI211_X1 U21372 ( .C1(n18480), .C2(n18299), .A(n18281), .B(n18280), .ZN(
        P3_U2924) );
  AOI22_X1 U21373 ( .A1(n18482), .A2(n18295), .B1(n18481), .B2(n18294), .ZN(
        n18283) );
  AOI22_X1 U21374 ( .A1(P3_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n18296), .B1(
        n18483), .B2(n18317), .ZN(n18282) );
  OAI211_X1 U21375 ( .C1(n18486), .C2(n18299), .A(n18283), .B(n18282), .ZN(
        P3_U2925) );
  AOI22_X1 U21376 ( .A1(n18489), .A2(n18317), .B1(n18487), .B2(n18294), .ZN(
        n18285) );
  AOI22_X1 U21377 ( .A1(P3_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n18296), .B1(
        n18488), .B2(n18295), .ZN(n18284) );
  OAI211_X1 U21378 ( .C1(n18492), .C2(n18299), .A(n18285), .B(n18284), .ZN(
        P3_U2926) );
  AOI22_X1 U21379 ( .A1(n18494), .A2(n18295), .B1(n18493), .B2(n18294), .ZN(
        n18287) );
  AOI22_X1 U21380 ( .A1(P3_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n18296), .B1(
        n18495), .B2(n18317), .ZN(n18286) );
  OAI211_X1 U21381 ( .C1(n18498), .C2(n18299), .A(n18287), .B(n18286), .ZN(
        P3_U2927) );
  AOI22_X1 U21382 ( .A1(n18499), .A2(n18294), .B1(n18501), .B2(n18317), .ZN(
        n18289) );
  AOI22_X1 U21383 ( .A1(P3_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n18296), .B1(
        n18500), .B2(n18295), .ZN(n18288) );
  OAI211_X1 U21384 ( .C1(n18504), .C2(n18299), .A(n18289), .B(n18288), .ZN(
        P3_U2928) );
  AOI22_X1 U21385 ( .A1(n18506), .A2(n18317), .B1(n18505), .B2(n18294), .ZN(
        n18291) );
  AOI22_X1 U21386 ( .A1(P3_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n18296), .B1(
        n18507), .B2(n18295), .ZN(n18290) );
  OAI211_X1 U21387 ( .C1(n18510), .C2(n18299), .A(n18291), .B(n18290), .ZN(
        P3_U2929) );
  AOI22_X1 U21388 ( .A1(n18513), .A2(n18317), .B1(n18511), .B2(n18294), .ZN(
        n18293) );
  AOI22_X1 U21389 ( .A1(P3_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n18296), .B1(
        n18512), .B2(n18295), .ZN(n18292) );
  OAI211_X1 U21390 ( .C1(n18516), .C2(n18299), .A(n18293), .B(n18292), .ZN(
        P3_U2930) );
  AOI22_X1 U21391 ( .A1(n18520), .A2(n18295), .B1(n18518), .B2(n18294), .ZN(
        n18298) );
  AOI22_X1 U21392 ( .A1(P3_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n18296), .B1(
        n18521), .B2(n18317), .ZN(n18297) );
  OAI211_X1 U21393 ( .C1(n18526), .C2(n18299), .A(n18298), .B(n18297), .ZN(
        P3_U2931) );
  NOR2_X2 U21394 ( .A1(n18572), .A2(n18371), .ZN(n18389) );
  INV_X1 U21395 ( .A(n18389), .ZN(n18321) );
  NOR2_X1 U21396 ( .A1(n18366), .A2(n18389), .ZN(n18349) );
  NOR2_X1 U21397 ( .A1(n9805), .A2(n18349), .ZN(n18316) );
  AOI22_X1 U21398 ( .A1(n18477), .A2(n18341), .B1(n18471), .B2(n18316), .ZN(
        n18303) );
  OAI21_X1 U21399 ( .B1(n18300), .B2(n18444), .A(n18349), .ZN(n18301) );
  OAI211_X1 U21400 ( .C1(n18389), .C2(n18696), .A(n18447), .B(n18301), .ZN(
        n18318) );
  AOI22_X1 U21401 ( .A1(P3_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n18318), .B1(
        n18472), .B2(n18317), .ZN(n18302) );
  OAI211_X1 U21402 ( .C1(n18480), .C2(n18321), .A(n18303), .B(n18302), .ZN(
        P3_U2932) );
  AOI22_X1 U21403 ( .A1(n18483), .A2(n18341), .B1(n18481), .B2(n18316), .ZN(
        n18305) );
  AOI22_X1 U21404 ( .A1(P3_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n18318), .B1(
        n18482), .B2(n18317), .ZN(n18304) );
  OAI211_X1 U21405 ( .C1(n18486), .C2(n18321), .A(n18305), .B(n18304), .ZN(
        P3_U2933) );
  AOI22_X1 U21406 ( .A1(n18489), .A2(n18341), .B1(n18487), .B2(n18316), .ZN(
        n18307) );
  AOI22_X1 U21407 ( .A1(P3_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n18318), .B1(
        n18488), .B2(n18317), .ZN(n18306) );
  OAI211_X1 U21408 ( .C1(n18492), .C2(n18321), .A(n18307), .B(n18306), .ZN(
        P3_U2934) );
  AOI22_X1 U21409 ( .A1(n18494), .A2(n18317), .B1(n18493), .B2(n18316), .ZN(
        n18309) );
  AOI22_X1 U21410 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n18318), .B1(
        n18495), .B2(n18341), .ZN(n18308) );
  OAI211_X1 U21411 ( .C1(n18498), .C2(n18321), .A(n18309), .B(n18308), .ZN(
        P3_U2935) );
  AOI22_X1 U21412 ( .A1(n18499), .A2(n18316), .B1(n18501), .B2(n18341), .ZN(
        n18311) );
  AOI22_X1 U21413 ( .A1(P3_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n18318), .B1(
        n18500), .B2(n18317), .ZN(n18310) );
  OAI211_X1 U21414 ( .C1(n18504), .C2(n18321), .A(n18311), .B(n18310), .ZN(
        P3_U2936) );
  AOI22_X1 U21415 ( .A1(n18506), .A2(n18341), .B1(n18505), .B2(n18316), .ZN(
        n18313) );
  AOI22_X1 U21416 ( .A1(P3_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n18318), .B1(
        n18507), .B2(n18317), .ZN(n18312) );
  OAI211_X1 U21417 ( .C1(n18510), .C2(n18321), .A(n18313), .B(n18312), .ZN(
        P3_U2937) );
  AOI22_X1 U21418 ( .A1(P3_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n18318), .B1(
        n18511), .B2(n18316), .ZN(n18315) );
  AOI22_X1 U21419 ( .A1(n18513), .A2(n18341), .B1(n18512), .B2(n18317), .ZN(
        n18314) );
  OAI211_X1 U21420 ( .C1(n18516), .C2(n18321), .A(n18315), .B(n18314), .ZN(
        P3_U2938) );
  AOI22_X1 U21421 ( .A1(n18521), .A2(n18341), .B1(n18518), .B2(n18316), .ZN(
        n18320) );
  AOI22_X1 U21422 ( .A1(P3_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n18318), .B1(
        n18520), .B2(n18317), .ZN(n18319) );
  OAI211_X1 U21423 ( .C1(n18526), .C2(n18321), .A(n18320), .B(n18319), .ZN(
        P3_U2939) );
  INV_X1 U21424 ( .A(n18371), .ZN(n18373) );
  NAND2_X1 U21425 ( .A1(n18322), .A2(n18373), .ZN(n18346) );
  AOI22_X1 U21426 ( .A1(n18477), .A2(n18366), .B1(n18471), .B2(n18340), .ZN(
        n18327) );
  NOR2_X1 U21427 ( .A1(P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n18323), .ZN(
        n18325) );
  NOR2_X1 U21428 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(n18371), .ZN(
        n18324) );
  AOI22_X1 U21429 ( .A1(n18476), .A2(n18325), .B1(n18474), .B2(n18324), .ZN(
        n18342) );
  AOI22_X1 U21430 ( .A1(P3_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n18342), .B1(
        n18472), .B2(n18341), .ZN(n18326) );
  OAI211_X1 U21431 ( .C1(n18480), .C2(n18346), .A(n18327), .B(n18326), .ZN(
        P3_U2940) );
  AOI22_X1 U21432 ( .A1(n18482), .A2(n18341), .B1(n18481), .B2(n18340), .ZN(
        n18329) );
  AOI22_X1 U21433 ( .A1(P3_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n18342), .B1(
        n18483), .B2(n18366), .ZN(n18328) );
  OAI211_X1 U21434 ( .C1(n18486), .C2(n18346), .A(n18329), .B(n18328), .ZN(
        P3_U2941) );
  AOI22_X1 U21435 ( .A1(n18488), .A2(n18341), .B1(n18487), .B2(n18340), .ZN(
        n18331) );
  AOI22_X1 U21436 ( .A1(P3_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n18342), .B1(
        n18489), .B2(n18366), .ZN(n18330) );
  OAI211_X1 U21437 ( .C1(n18492), .C2(n18346), .A(n18331), .B(n18330), .ZN(
        P3_U2942) );
  AOI22_X1 U21438 ( .A1(n18494), .A2(n18341), .B1(n18493), .B2(n18340), .ZN(
        n18333) );
  AOI22_X1 U21439 ( .A1(P3_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n18342), .B1(
        n18495), .B2(n18366), .ZN(n18332) );
  OAI211_X1 U21440 ( .C1(n18498), .C2(n18346), .A(n18333), .B(n18332), .ZN(
        P3_U2943) );
  AOI22_X1 U21441 ( .A1(n18500), .A2(n18341), .B1(n18499), .B2(n18340), .ZN(
        n18335) );
  AOI22_X1 U21442 ( .A1(P3_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n18342), .B1(
        n18501), .B2(n18366), .ZN(n18334) );
  OAI211_X1 U21443 ( .C1(n18504), .C2(n18346), .A(n18335), .B(n18334), .ZN(
        P3_U2944) );
  AOI22_X1 U21444 ( .A1(n18507), .A2(n18341), .B1(n18505), .B2(n18340), .ZN(
        n18337) );
  AOI22_X1 U21445 ( .A1(P3_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n18342), .B1(
        n18506), .B2(n18366), .ZN(n18336) );
  OAI211_X1 U21446 ( .C1(n18510), .C2(n18346), .A(n18337), .B(n18336), .ZN(
        P3_U2945) );
  AOI22_X1 U21447 ( .A1(n18513), .A2(n18366), .B1(n18511), .B2(n18340), .ZN(
        n18339) );
  AOI22_X1 U21448 ( .A1(P3_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n18342), .B1(
        n18512), .B2(n18341), .ZN(n18338) );
  OAI211_X1 U21449 ( .C1(n18516), .C2(n18346), .A(n18339), .B(n18338), .ZN(
        P3_U2946) );
  AOI22_X1 U21450 ( .A1(n18520), .A2(n18341), .B1(n18518), .B2(n18340), .ZN(
        n18344) );
  AOI22_X1 U21451 ( .A1(P3_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n18342), .B1(
        n18521), .B2(n18366), .ZN(n18343) );
  OAI211_X1 U21452 ( .C1(n18526), .C2(n18346), .A(n18344), .B(n18343), .ZN(
        P3_U2947) );
  NAND2_X1 U21453 ( .A1(n18345), .A2(n18373), .ZN(n18370) );
  AOI21_X1 U21454 ( .B1(n18346), .B2(n18370), .A(n9805), .ZN(n18365) );
  AOI22_X1 U21455 ( .A1(n18477), .A2(n18389), .B1(n18471), .B2(n18365), .ZN(
        n18352) );
  INV_X1 U21456 ( .A(n18370), .ZN(n18438) );
  INV_X1 U21457 ( .A(n18346), .ZN(n18414) );
  NOR2_X1 U21458 ( .A1(n18414), .A2(n18438), .ZN(n18347) );
  OAI22_X1 U21459 ( .A1(n18349), .A2(n18348), .B1(n18347), .B2(n18394), .ZN(
        n18350) );
  OAI21_X1 U21460 ( .B1(n18438), .B2(n18696), .A(n18350), .ZN(n18367) );
  AOI22_X1 U21461 ( .A1(P3_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n18367), .B1(
        n18472), .B2(n18366), .ZN(n18351) );
  OAI211_X1 U21462 ( .C1(n18480), .C2(n18370), .A(n18352), .B(n18351), .ZN(
        P3_U2948) );
  AOI22_X1 U21463 ( .A1(n18483), .A2(n18389), .B1(n18481), .B2(n18365), .ZN(
        n18354) );
  AOI22_X1 U21464 ( .A1(P3_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n18367), .B1(
        n18482), .B2(n18366), .ZN(n18353) );
  OAI211_X1 U21465 ( .C1(n18486), .C2(n18370), .A(n18354), .B(n18353), .ZN(
        P3_U2949) );
  AOI22_X1 U21466 ( .A1(n18489), .A2(n18389), .B1(n18487), .B2(n18365), .ZN(
        n18356) );
  AOI22_X1 U21467 ( .A1(P3_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n18367), .B1(
        n18488), .B2(n18366), .ZN(n18355) );
  OAI211_X1 U21468 ( .C1(n18492), .C2(n18370), .A(n18356), .B(n18355), .ZN(
        P3_U2950) );
  AOI22_X1 U21469 ( .A1(n18494), .A2(n18366), .B1(n18493), .B2(n18365), .ZN(
        n18358) );
  AOI22_X1 U21470 ( .A1(P3_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n18367), .B1(
        n18495), .B2(n18389), .ZN(n18357) );
  OAI211_X1 U21471 ( .C1(n18498), .C2(n18370), .A(n18358), .B(n18357), .ZN(
        P3_U2951) );
  AOI22_X1 U21472 ( .A1(n18499), .A2(n18365), .B1(n18501), .B2(n18389), .ZN(
        n18360) );
  AOI22_X1 U21473 ( .A1(P3_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n18367), .B1(
        n18500), .B2(n18366), .ZN(n18359) );
  OAI211_X1 U21474 ( .C1(n18504), .C2(n18370), .A(n18360), .B(n18359), .ZN(
        P3_U2952) );
  AOI22_X1 U21475 ( .A1(n18507), .A2(n18366), .B1(n18505), .B2(n18365), .ZN(
        n18362) );
  AOI22_X1 U21476 ( .A1(P3_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n18367), .B1(
        n18506), .B2(n18389), .ZN(n18361) );
  OAI211_X1 U21477 ( .C1(n18510), .C2(n18370), .A(n18362), .B(n18361), .ZN(
        P3_U2953) );
  AOI22_X1 U21478 ( .A1(n18512), .A2(n18366), .B1(n18511), .B2(n18365), .ZN(
        n18364) );
  AOI22_X1 U21479 ( .A1(P3_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n18367), .B1(
        n18513), .B2(n18389), .ZN(n18363) );
  OAI211_X1 U21480 ( .C1(n18516), .C2(n18370), .A(n18364), .B(n18363), .ZN(
        P3_U2954) );
  AOI22_X1 U21481 ( .A1(n18521), .A2(n18389), .B1(n18518), .B2(n18365), .ZN(
        n18369) );
  AOI22_X1 U21482 ( .A1(P3_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n18367), .B1(
        n18520), .B2(n18366), .ZN(n18368) );
  OAI211_X1 U21483 ( .C1(n18526), .C2(n18370), .A(n18369), .B(n18368), .ZN(
        P3_U2955) );
  NOR2_X2 U21484 ( .A1(n18571), .A2(n18371), .ZN(n18464) );
  INV_X1 U21485 ( .A(n18464), .ZN(n18393) );
  NOR2_X1 U21486 ( .A1(n20944), .A2(n18371), .ZN(n18422) );
  INV_X1 U21487 ( .A(n18422), .ZN(n18372) );
  NOR2_X1 U21488 ( .A1(n9805), .A2(n18372), .ZN(n18388) );
  AOI22_X1 U21489 ( .A1(n18477), .A2(n18414), .B1(n18471), .B2(n18388), .ZN(
        n18375) );
  OAI211_X1 U21490 ( .C1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .C2(n18476), .A(
        n18474), .B(n18373), .ZN(n18390) );
  AOI22_X1 U21491 ( .A1(P3_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n18390), .B1(
        n18472), .B2(n18389), .ZN(n18374) );
  OAI211_X1 U21492 ( .C1(n18480), .C2(n18393), .A(n18375), .B(n18374), .ZN(
        P3_U2956) );
  AOI22_X1 U21493 ( .A1(n18483), .A2(n18414), .B1(n18481), .B2(n18388), .ZN(
        n18377) );
  AOI22_X1 U21494 ( .A1(P3_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n18390), .B1(
        n18482), .B2(n18389), .ZN(n18376) );
  OAI211_X1 U21495 ( .C1(n18486), .C2(n18393), .A(n18377), .B(n18376), .ZN(
        P3_U2957) );
  AOI22_X1 U21496 ( .A1(n18489), .A2(n18414), .B1(n18487), .B2(n18388), .ZN(
        n18379) );
  AOI22_X1 U21497 ( .A1(P3_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n18390), .B1(
        n18488), .B2(n18389), .ZN(n18378) );
  OAI211_X1 U21498 ( .C1(n18492), .C2(n18393), .A(n18379), .B(n18378), .ZN(
        P3_U2958) );
  AOI22_X1 U21499 ( .A1(n18494), .A2(n18389), .B1(n18493), .B2(n18388), .ZN(
        n18381) );
  AOI22_X1 U21500 ( .A1(P3_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n18390), .B1(
        n18495), .B2(n18414), .ZN(n18380) );
  OAI211_X1 U21501 ( .C1(n18498), .C2(n18393), .A(n18381), .B(n18380), .ZN(
        P3_U2959) );
  AOI22_X1 U21502 ( .A1(n18499), .A2(n18388), .B1(n18501), .B2(n18414), .ZN(
        n18383) );
  AOI22_X1 U21503 ( .A1(P3_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n18390), .B1(
        n18500), .B2(n18389), .ZN(n18382) );
  OAI211_X1 U21504 ( .C1(n18504), .C2(n18393), .A(n18383), .B(n18382), .ZN(
        P3_U2960) );
  AOI22_X1 U21505 ( .A1(n18507), .A2(n18389), .B1(n18505), .B2(n18388), .ZN(
        n18385) );
  AOI22_X1 U21506 ( .A1(P3_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n18390), .B1(
        n18506), .B2(n18414), .ZN(n18384) );
  OAI211_X1 U21507 ( .C1(n18510), .C2(n18393), .A(n18385), .B(n18384), .ZN(
        P3_U2961) );
  AOI22_X1 U21508 ( .A1(n18513), .A2(n18414), .B1(n18511), .B2(n18388), .ZN(
        n18387) );
  AOI22_X1 U21509 ( .A1(P3_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n18390), .B1(
        n18512), .B2(n18389), .ZN(n18386) );
  OAI211_X1 U21510 ( .C1(n18516), .C2(n18393), .A(n18387), .B(n18386), .ZN(
        P3_U2962) );
  AOI22_X1 U21511 ( .A1(n18521), .A2(n18414), .B1(n18518), .B2(n18388), .ZN(
        n18392) );
  AOI22_X1 U21512 ( .A1(P3_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n18390), .B1(
        n18520), .B2(n18389), .ZN(n18391) );
  OAI211_X1 U21513 ( .C1(n18526), .C2(n18393), .A(n18392), .B(n18391), .ZN(
        P3_U2963) );
  INV_X1 U21514 ( .A(n18475), .ZN(n18419) );
  NOR2_X2 U21515 ( .A1(n18419), .A2(P3_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(
        n18519) );
  INV_X1 U21516 ( .A(n18519), .ZN(n18418) );
  NAND2_X1 U21517 ( .A1(n18393), .A2(n18418), .ZN(n18398) );
  INV_X1 U21518 ( .A(n18398), .ZN(n18445) );
  NOR2_X1 U21519 ( .A1(n9805), .A2(n18445), .ZN(n18413) );
  AOI22_X1 U21520 ( .A1(n18477), .A2(n18438), .B1(n18471), .B2(n18413), .ZN(
        n18400) );
  AOI21_X1 U21521 ( .B1(P3_STATE2_REG_3__SCAN_IN), .B2(n18418), .A(n18394), 
        .ZN(n18395) );
  OAI221_X1 U21522 ( .B1(n18398), .B2(n18397), .C1(n18398), .C2(n18396), .A(
        n18395), .ZN(n18415) );
  AOI22_X1 U21523 ( .A1(P3_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n18415), .B1(
        n18472), .B2(n18414), .ZN(n18399) );
  OAI211_X1 U21524 ( .C1(n18480), .C2(n18418), .A(n18400), .B(n18399), .ZN(
        P3_U2964) );
  AOI22_X1 U21525 ( .A1(P3_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n18415), .B1(
        n18481), .B2(n18413), .ZN(n18402) );
  AOI22_X1 U21526 ( .A1(n18482), .A2(n18414), .B1(n18483), .B2(n18438), .ZN(
        n18401) );
  OAI211_X1 U21527 ( .C1(n18486), .C2(n18418), .A(n18402), .B(n18401), .ZN(
        P3_U2965) );
  AOI22_X1 U21528 ( .A1(n18488), .A2(n18414), .B1(n18487), .B2(n18413), .ZN(
        n18404) );
  AOI22_X1 U21529 ( .A1(P3_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n18415), .B1(
        n18489), .B2(n18438), .ZN(n18403) );
  OAI211_X1 U21530 ( .C1(n18492), .C2(n18418), .A(n18404), .B(n18403), .ZN(
        P3_U2966) );
  AOI22_X1 U21531 ( .A1(P3_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n18415), .B1(
        n18493), .B2(n18413), .ZN(n18406) );
  AOI22_X1 U21532 ( .A1(n18495), .A2(n18438), .B1(n18494), .B2(n18414), .ZN(
        n18405) );
  OAI211_X1 U21533 ( .C1(n18498), .C2(n18418), .A(n18406), .B(n18405), .ZN(
        P3_U2967) );
  AOI22_X1 U21534 ( .A1(P3_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n18415), .B1(
        n18499), .B2(n18413), .ZN(n18408) );
  AOI22_X1 U21535 ( .A1(n18500), .A2(n18414), .B1(n18501), .B2(n18438), .ZN(
        n18407) );
  OAI211_X1 U21536 ( .C1(n18504), .C2(n18418), .A(n18408), .B(n18407), .ZN(
        P3_U2968) );
  AOI22_X1 U21537 ( .A1(n18507), .A2(n18414), .B1(n18505), .B2(n18413), .ZN(
        n18410) );
  AOI22_X1 U21538 ( .A1(P3_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n18415), .B1(
        n18506), .B2(n18438), .ZN(n18409) );
  OAI211_X1 U21539 ( .C1(n18510), .C2(n18418), .A(n18410), .B(n18409), .ZN(
        P3_U2969) );
  AOI22_X1 U21540 ( .A1(P3_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n18415), .B1(
        n18511), .B2(n18413), .ZN(n18412) );
  AOI22_X1 U21541 ( .A1(n18513), .A2(n18438), .B1(n18512), .B2(n18414), .ZN(
        n18411) );
  OAI211_X1 U21542 ( .C1(n18516), .C2(n18418), .A(n18412), .B(n18411), .ZN(
        P3_U2970) );
  AOI22_X1 U21543 ( .A1(n18520), .A2(n18414), .B1(n18518), .B2(n18413), .ZN(
        n18417) );
  AOI22_X1 U21544 ( .A1(P3_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n18415), .B1(
        n18521), .B2(n18438), .ZN(n18416) );
  OAI211_X1 U21545 ( .C1(n18526), .C2(n18418), .A(n18417), .B(n18416), .ZN(
        P3_U2971) );
  NOR2_X1 U21546 ( .A1(n9805), .A2(n18419), .ZN(n18437) );
  AOI22_X1 U21547 ( .A1(n18472), .A2(n18438), .B1(n18471), .B2(n18437), .ZN(
        n18424) );
  AOI22_X1 U21548 ( .A1(n18476), .A2(n18422), .B1(n18421), .B2(n18420), .ZN(
        n18439) );
  AOI22_X1 U21549 ( .A1(P3_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n18439), .B1(
        n18477), .B2(n18464), .ZN(n18423) );
  OAI211_X1 U21550 ( .C1(n18480), .C2(n18442), .A(n18424), .B(n18423), .ZN(
        P3_U2972) );
  AOI22_X1 U21551 ( .A1(n18482), .A2(n18438), .B1(n18481), .B2(n18437), .ZN(
        n18426) );
  AOI22_X1 U21552 ( .A1(P3_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n18439), .B1(
        n18483), .B2(n18464), .ZN(n18425) );
  OAI211_X1 U21553 ( .C1(n18442), .C2(n18486), .A(n18426), .B(n18425), .ZN(
        P3_U2973) );
  AOI22_X1 U21554 ( .A1(n18489), .A2(n18464), .B1(n18487), .B2(n18437), .ZN(
        n18428) );
  AOI22_X1 U21555 ( .A1(P3_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n18439), .B1(
        n18488), .B2(n18438), .ZN(n18427) );
  OAI211_X1 U21556 ( .C1(n18442), .C2(n18492), .A(n18428), .B(n18427), .ZN(
        P3_U2974) );
  AOI22_X1 U21557 ( .A1(n18495), .A2(n18464), .B1(n18493), .B2(n18437), .ZN(
        n18430) );
  AOI22_X1 U21558 ( .A1(P3_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n18439), .B1(
        n18494), .B2(n18438), .ZN(n18429) );
  OAI211_X1 U21559 ( .C1(n18442), .C2(n18498), .A(n18430), .B(n18429), .ZN(
        P3_U2975) );
  AOI22_X1 U21560 ( .A1(n18500), .A2(n18438), .B1(n18499), .B2(n18437), .ZN(
        n18432) );
  AOI22_X1 U21561 ( .A1(P3_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n18439), .B1(
        n18501), .B2(n18464), .ZN(n18431) );
  OAI211_X1 U21562 ( .C1(n18442), .C2(n18504), .A(n18432), .B(n18431), .ZN(
        P3_U2976) );
  AOI22_X1 U21563 ( .A1(n18507), .A2(n18438), .B1(n18505), .B2(n18437), .ZN(
        n18434) );
  AOI22_X1 U21564 ( .A1(P3_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n18439), .B1(
        n18506), .B2(n18464), .ZN(n18433) );
  OAI211_X1 U21565 ( .C1(n18442), .C2(n18510), .A(n18434), .B(n18433), .ZN(
        P3_U2977) );
  AOI22_X1 U21566 ( .A1(n18513), .A2(n18464), .B1(n18511), .B2(n18437), .ZN(
        n18436) );
  AOI22_X1 U21567 ( .A1(P3_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n18439), .B1(
        n18512), .B2(n18438), .ZN(n18435) );
  OAI211_X1 U21568 ( .C1(n18442), .C2(n18516), .A(n18436), .B(n18435), .ZN(
        P3_U2978) );
  AOI22_X1 U21569 ( .A1(n18520), .A2(n18438), .B1(n18518), .B2(n18437), .ZN(
        n18441) );
  AOI22_X1 U21570 ( .A1(P3_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n18439), .B1(
        n18521), .B2(n18464), .ZN(n18440) );
  OAI211_X1 U21571 ( .C1(n18442), .C2(n18526), .A(n18441), .B(n18440), .ZN(
        P3_U2979) );
  NOR2_X1 U21572 ( .A1(n9805), .A2(n18443), .ZN(n18463) );
  AOI22_X1 U21573 ( .A1(n18472), .A2(n18464), .B1(n18471), .B2(n18463), .ZN(
        n18450) );
  OAI21_X1 U21574 ( .B1(n18445), .B2(n18444), .A(n18443), .ZN(n18446) );
  OAI211_X1 U21575 ( .C1(n18448), .C2(n18696), .A(n18447), .B(n18446), .ZN(
        n18465) );
  AOI22_X1 U21576 ( .A1(P3_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n18465), .B1(
        n18477), .B2(n18519), .ZN(n18449) );
  OAI211_X1 U21577 ( .C1(n18468), .C2(n18480), .A(n18450), .B(n18449), .ZN(
        P3_U2980) );
  AOI22_X1 U21578 ( .A1(n18482), .A2(n18464), .B1(n18481), .B2(n18463), .ZN(
        n18452) );
  AOI22_X1 U21579 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n18465), .B1(
        n18483), .B2(n18519), .ZN(n18451) );
  OAI211_X1 U21580 ( .C1(n18468), .C2(n18486), .A(n18452), .B(n18451), .ZN(
        P3_U2981) );
  AOI22_X1 U21581 ( .A1(n18488), .A2(n18464), .B1(n18487), .B2(n18463), .ZN(
        n18454) );
  AOI22_X1 U21582 ( .A1(P3_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n18465), .B1(
        n18489), .B2(n18519), .ZN(n18453) );
  OAI211_X1 U21583 ( .C1(n18468), .C2(n18492), .A(n18454), .B(n18453), .ZN(
        P3_U2982) );
  AOI22_X1 U21584 ( .A1(n18495), .A2(n18519), .B1(n18493), .B2(n18463), .ZN(
        n18456) );
  AOI22_X1 U21585 ( .A1(P3_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n18465), .B1(
        n18494), .B2(n18464), .ZN(n18455) );
  OAI211_X1 U21586 ( .C1(n18468), .C2(n18498), .A(n18456), .B(n18455), .ZN(
        P3_U2983) );
  AOI22_X1 U21587 ( .A1(n18499), .A2(n18463), .B1(n18501), .B2(n18519), .ZN(
        n18458) );
  AOI22_X1 U21588 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n18465), .B1(
        n18500), .B2(n18464), .ZN(n18457) );
  OAI211_X1 U21589 ( .C1(n18468), .C2(n18504), .A(n18458), .B(n18457), .ZN(
        P3_U2984) );
  AOI22_X1 U21590 ( .A1(n18506), .A2(n18519), .B1(n18505), .B2(n18463), .ZN(
        n18460) );
  AOI22_X1 U21591 ( .A1(P3_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n18465), .B1(
        n18507), .B2(n18464), .ZN(n18459) );
  OAI211_X1 U21592 ( .C1(n18468), .C2(n18510), .A(n18460), .B(n18459), .ZN(
        P3_U2985) );
  AOI22_X1 U21593 ( .A1(n18513), .A2(n18519), .B1(n18511), .B2(n18463), .ZN(
        n18462) );
  AOI22_X1 U21594 ( .A1(P3_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n18465), .B1(
        n18512), .B2(n18464), .ZN(n18461) );
  OAI211_X1 U21595 ( .C1(n18468), .C2(n18516), .A(n18462), .B(n18461), .ZN(
        P3_U2986) );
  AOI22_X1 U21596 ( .A1(n18521), .A2(n18519), .B1(n18518), .B2(n18463), .ZN(
        n18467) );
  AOI22_X1 U21597 ( .A1(P3_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n18465), .B1(
        n18520), .B2(n18464), .ZN(n18466) );
  OAI211_X1 U21598 ( .C1(n18468), .C2(n18526), .A(n18467), .B(n18466), .ZN(
        P3_U2987) );
  INV_X1 U21599 ( .A(n18469), .ZN(n18527) );
  INV_X1 U21600 ( .A(n18473), .ZN(n18470) );
  NOR2_X1 U21601 ( .A1(n9805), .A2(n18470), .ZN(n18517) );
  AOI22_X1 U21602 ( .A1(n18472), .A2(n18519), .B1(n18471), .B2(n18517), .ZN(
        n18479) );
  AOI22_X1 U21603 ( .A1(n18476), .A2(n18475), .B1(n18474), .B2(n18473), .ZN(
        n18523) );
  AOI22_X1 U21604 ( .A1(P3_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n18523), .B1(
        n18477), .B2(n18522), .ZN(n18478) );
  OAI211_X1 U21605 ( .C1(n18527), .C2(n18480), .A(n18479), .B(n18478), .ZN(
        P3_U2988) );
  AOI22_X1 U21606 ( .A1(n18482), .A2(n18519), .B1(n18481), .B2(n18517), .ZN(
        n18485) );
  AOI22_X1 U21607 ( .A1(P3_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n18523), .B1(
        n18522), .B2(n18483), .ZN(n18484) );
  OAI211_X1 U21608 ( .C1(n18527), .C2(n18486), .A(n18485), .B(n18484), .ZN(
        P3_U2989) );
  AOI22_X1 U21609 ( .A1(n18488), .A2(n18519), .B1(n18487), .B2(n18517), .ZN(
        n18491) );
  AOI22_X1 U21610 ( .A1(P3_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n18523), .B1(
        n18522), .B2(n18489), .ZN(n18490) );
  OAI211_X1 U21611 ( .C1(n18527), .C2(n18492), .A(n18491), .B(n18490), .ZN(
        P3_U2990) );
  AOI22_X1 U21612 ( .A1(n18494), .A2(n18519), .B1(n18493), .B2(n18517), .ZN(
        n18497) );
  AOI22_X1 U21613 ( .A1(P3_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n18523), .B1(
        n18522), .B2(n18495), .ZN(n18496) );
  OAI211_X1 U21614 ( .C1(n18527), .C2(n18498), .A(n18497), .B(n18496), .ZN(
        P3_U2991) );
  AOI22_X1 U21615 ( .A1(n18500), .A2(n18519), .B1(n18499), .B2(n18517), .ZN(
        n18503) );
  AOI22_X1 U21616 ( .A1(P3_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n18523), .B1(
        n18522), .B2(n18501), .ZN(n18502) );
  OAI211_X1 U21617 ( .C1(n18527), .C2(n18504), .A(n18503), .B(n18502), .ZN(
        P3_U2992) );
  AOI22_X1 U21618 ( .A1(n18522), .A2(n18506), .B1(n18505), .B2(n18517), .ZN(
        n18509) );
  AOI22_X1 U21619 ( .A1(P3_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n18523), .B1(
        n18507), .B2(n18519), .ZN(n18508) );
  OAI211_X1 U21620 ( .C1(n18527), .C2(n18510), .A(n18509), .B(n18508), .ZN(
        P3_U2993) );
  AOI22_X1 U21621 ( .A1(n18512), .A2(n18519), .B1(n18511), .B2(n18517), .ZN(
        n18515) );
  AOI22_X1 U21622 ( .A1(P3_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n18523), .B1(
        n18522), .B2(n18513), .ZN(n18514) );
  OAI211_X1 U21623 ( .C1(n18527), .C2(n18516), .A(n18515), .B(n18514), .ZN(
        P3_U2994) );
  AOI22_X1 U21624 ( .A1(n18520), .A2(n18519), .B1(n18518), .B2(n18517), .ZN(
        n18525) );
  AOI22_X1 U21625 ( .A1(P3_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n18523), .B1(
        n18522), .B2(n18521), .ZN(n18524) );
  OAI211_X1 U21626 ( .C1(n18527), .C2(n18526), .A(n18525), .B(n18524), .ZN(
        P3_U2995) );
  NAND2_X1 U21627 ( .A1(n9878), .A2(n18528), .ZN(n18529) );
  AOI22_X1 U21628 ( .A1(n18532), .A2(n18531), .B1(n18530), .B2(n18529), .ZN(
        n18533) );
  OAI221_X1 U21629 ( .B1(n18535), .B2(n18561), .C1(n18535), .C2(n18534), .A(
        n18533), .ZN(n18739) );
  OAI21_X1 U21630 ( .B1(P3_MORE_REG_SCAN_IN), .B2(P3_FLUSH_REG_SCAN_IN), .A(
        n18536), .ZN(n18538) );
  OAI211_X1 U21631 ( .C1(n18565), .C2(n18539), .A(n18538), .B(n18537), .ZN(
        n18585) );
  NOR2_X1 U21632 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18549), .ZN(
        n18569) );
  INV_X1 U21633 ( .A(n18569), .ZN(n18541) );
  NAND2_X1 U21634 ( .A1(n18713), .A2(n18563), .ZN(n18546) );
  AOI22_X1 U21635 ( .A1(n18542), .A2(n18541), .B1(n18540), .B2(n18546), .ZN(
        n18698) );
  NOR2_X1 U21636 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18698), .ZN(
        n18551) );
  AOI21_X1 U21637 ( .B1(n18545), .B2(n18544), .A(n18543), .ZN(n18553) );
  OAI21_X1 U21638 ( .B1(n18553), .B2(n18547), .A(n18546), .ZN(n18548) );
  AOI21_X1 U21639 ( .B1(n18557), .B2(n18549), .A(n18548), .ZN(n18701) );
  NAND2_X1 U21640 ( .A1(n18565), .A2(n18701), .ZN(n18550) );
  AOI22_X1 U21641 ( .A1(n18565), .A2(n18551), .B1(
        P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n18550), .ZN(n18583) );
  INV_X1 U21642 ( .A(n18565), .ZN(n18574) );
  AOI221_X1 U21643 ( .B1(P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18553), 
        .C1(n18552), .C2(n18553), .A(n18713), .ZN(n18564) );
  NOR2_X1 U21644 ( .A1(n18554), .A2(n18727), .ZN(n18556) );
  OAI211_X1 U21645 ( .C1(n18556), .C2(n18555), .A(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(n18713), .ZN(n18560) );
  OAI211_X1 U21646 ( .C1(P3_INSTQUEUERD_ADDR_REG_2__SCAN_IN), .C2(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n18558), .B(n18557), .ZN(
        n18559) );
  OAI211_X1 U21647 ( .C1(n18709), .C2(n18561), .A(n18560), .B(n18559), .ZN(
        n18562) );
  AOI21_X1 U21648 ( .B1(n18564), .B2(n18563), .A(n18562), .ZN(n18705) );
  AOI22_X1 U21649 ( .A1(n18574), .A2(n18713), .B1(n18705), .B2(n18565), .ZN(
        n18578) );
  NOR2_X1 U21650 ( .A1(n18567), .A2(n18566), .ZN(n18570) );
  AOI22_X1 U21651 ( .A1(P3_INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n18568), .B1(
        n18570), .B2(n18727), .ZN(n18722) );
  OAI22_X1 U21652 ( .A1(n18570), .A2(n18714), .B1(
        P3_INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B2(n18569), .ZN(n18718) );
  AOI222_X1 U21653 ( .A1(n18722), .A2(n18718), .B1(n18722), .B2(n20944), .C1(
        n18718), .C2(n18571), .ZN(n18573) );
  OAI21_X1 U21654 ( .B1(n18574), .B2(n18573), .A(n18572), .ZN(n18577) );
  AND2_X1 U21655 ( .A1(n18578), .A2(n18577), .ZN(n18575) );
  OAI221_X1 U21656 ( .B1(n18578), .B2(n18577), .C1(n18576), .C2(n18575), .A(
        n18580), .ZN(n18582) );
  AOI21_X1 U21657 ( .B1(n18580), .B2(n18579), .A(n18578), .ZN(n18581) );
  AOI222_X1 U21658 ( .A1(n18583), .A2(n18582), .B1(n18583), .B2(
        P3_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C1(n18582), .C2(n18581), .ZN(
        n18584) );
  NOR4_X1 U21659 ( .A1(n18586), .A2(n18739), .A3(n18585), .A4(n18584), .ZN(
        n18596) );
  AOI22_X1 U21660 ( .A1(n18615), .A2(n18743), .B1(n18721), .B2(n18749), .ZN(
        n18587) );
  INV_X1 U21661 ( .A(n18587), .ZN(n18592) );
  OAI211_X1 U21662 ( .C1(n18589), .C2(n18588), .A(n18741), .B(n18596), .ZN(
        n18695) );
  OAI21_X1 U21663 ( .B1(P3_STATE2_REG_2__SCAN_IN), .B2(n18747), .A(n18695), 
        .ZN(n18597) );
  NOR2_X1 U21664 ( .A1(n18590), .A2(n18597), .ZN(n18591) );
  MUX2_X1 U21665 ( .A(n18592), .B(n18591), .S(P3_STATE2_REG_0__SCAN_IN), .Z(
        n18594) );
  OAI211_X1 U21666 ( .C1(n18596), .C2(n18595), .A(n18594), .B(n18593), .ZN(
        P3_U2996) );
  NAND2_X1 U21667 ( .A1(n18615), .A2(n18743), .ZN(n18601) );
  NAND4_X1 U21668 ( .A1(P3_STATE2_REG_0__SCAN_IN), .A2(
        P3_STATE2_REG_1__SCAN_IN), .A3(n18615), .A4(n18603), .ZN(n18605) );
  OR3_X1 U21669 ( .A1(n9805), .A2(n18598), .A3(n18597), .ZN(n18600) );
  NAND4_X1 U21670 ( .A1(n18602), .A2(n18601), .A3(n18605), .A4(n18600), .ZN(
        P3_U2997) );
  NAND3_X1 U21671 ( .A1(n18604), .A2(n18603), .A3(n18745), .ZN(n18606) );
  AND4_X1 U21672 ( .A1(n18607), .A2(n18606), .A3(n18605), .A4(n18694), .ZN(
        P3_U2998) );
  INV_X1 U21673 ( .A(n18693), .ZN(n18608) );
  AND2_X1 U21674 ( .A1(P3_DATAWIDTH_REG_31__SCAN_IN), .A2(n18608), .ZN(
        P3_U2999) );
  AND2_X1 U21675 ( .A1(P3_DATAWIDTH_REG_30__SCAN_IN), .A2(n18608), .ZN(
        P3_U3000) );
  AND2_X1 U21676 ( .A1(P3_DATAWIDTH_REG_29__SCAN_IN), .A2(n18608), .ZN(
        P3_U3001) );
  AND2_X1 U21677 ( .A1(P3_DATAWIDTH_REG_28__SCAN_IN), .A2(n18608), .ZN(
        P3_U3002) );
  AND2_X1 U21678 ( .A1(P3_DATAWIDTH_REG_27__SCAN_IN), .A2(n18608), .ZN(
        P3_U3003) );
  AND2_X1 U21679 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(n18608), .ZN(
        P3_U3004) );
  AND2_X1 U21680 ( .A1(P3_DATAWIDTH_REG_25__SCAN_IN), .A2(n18608), .ZN(
        P3_U3005) );
  AND2_X1 U21681 ( .A1(P3_DATAWIDTH_REG_24__SCAN_IN), .A2(n18608), .ZN(
        P3_U3006) );
  AND2_X1 U21682 ( .A1(P3_DATAWIDTH_REG_23__SCAN_IN), .A2(n18608), .ZN(
        P3_U3007) );
  AND2_X1 U21683 ( .A1(P3_DATAWIDTH_REG_22__SCAN_IN), .A2(n18608), .ZN(
        P3_U3008) );
  AND2_X1 U21684 ( .A1(P3_DATAWIDTH_REG_21__SCAN_IN), .A2(n18608), .ZN(
        P3_U3009) );
  AND2_X1 U21685 ( .A1(P3_DATAWIDTH_REG_20__SCAN_IN), .A2(n18608), .ZN(
        P3_U3010) );
  AND2_X1 U21686 ( .A1(P3_DATAWIDTH_REG_19__SCAN_IN), .A2(n18608), .ZN(
        P3_U3011) );
  AND2_X1 U21687 ( .A1(P3_DATAWIDTH_REG_18__SCAN_IN), .A2(n18608), .ZN(
        P3_U3012) );
  AND2_X1 U21688 ( .A1(P3_DATAWIDTH_REG_17__SCAN_IN), .A2(n18608), .ZN(
        P3_U3013) );
  AND2_X1 U21689 ( .A1(P3_DATAWIDTH_REG_16__SCAN_IN), .A2(n18608), .ZN(
        P3_U3014) );
  AND2_X1 U21690 ( .A1(P3_DATAWIDTH_REG_15__SCAN_IN), .A2(n18608), .ZN(
        P3_U3015) );
  AND2_X1 U21691 ( .A1(P3_DATAWIDTH_REG_14__SCAN_IN), .A2(n18608), .ZN(
        P3_U3016) );
  AND2_X1 U21692 ( .A1(P3_DATAWIDTH_REG_13__SCAN_IN), .A2(n18608), .ZN(
        P3_U3017) );
  AND2_X1 U21693 ( .A1(P3_DATAWIDTH_REG_12__SCAN_IN), .A2(n18608), .ZN(
        P3_U3018) );
  AND2_X1 U21694 ( .A1(P3_DATAWIDTH_REG_11__SCAN_IN), .A2(n18608), .ZN(
        P3_U3019) );
  AND2_X1 U21695 ( .A1(P3_DATAWIDTH_REG_10__SCAN_IN), .A2(n18608), .ZN(
        P3_U3020) );
  AND2_X1 U21696 ( .A1(P3_DATAWIDTH_REG_9__SCAN_IN), .A2(n18608), .ZN(P3_U3021) );
  AND2_X1 U21697 ( .A1(P3_DATAWIDTH_REG_8__SCAN_IN), .A2(n18608), .ZN(P3_U3022) );
  AND2_X1 U21698 ( .A1(P3_DATAWIDTH_REG_7__SCAN_IN), .A2(n18608), .ZN(P3_U3023) );
  AND2_X1 U21699 ( .A1(P3_DATAWIDTH_REG_6__SCAN_IN), .A2(n18608), .ZN(P3_U3024) );
  AND2_X1 U21700 ( .A1(P3_DATAWIDTH_REG_5__SCAN_IN), .A2(n18608), .ZN(P3_U3025) );
  AND2_X1 U21701 ( .A1(P3_DATAWIDTH_REG_4__SCAN_IN), .A2(n18608), .ZN(P3_U3026) );
  AND2_X1 U21702 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(n18608), .ZN(P3_U3027) );
  AND2_X1 U21703 ( .A1(P3_DATAWIDTH_REG_2__SCAN_IN), .A2(n18608), .ZN(P3_U3028) );
  OAI21_X1 U21704 ( .B1(n18609), .B2(n20700), .A(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(n18610) );
  AOI22_X1 U21705 ( .A1(n18623), .A2(n18625), .B1(n18755), .B2(n18610), .ZN(
        n18611) );
  NAND3_X1 U21706 ( .A1(NA), .A2(n18623), .A3(n20880), .ZN(n18618) );
  OAI211_X1 U21707 ( .C1(n18747), .C2(n18612), .A(n18611), .B(n18618), .ZN(
        P3_U3029) );
  NOR2_X1 U21708 ( .A1(n18625), .A2(n20700), .ZN(n18621) );
  INV_X1 U21709 ( .A(n18621), .ZN(n18614) );
  INV_X1 U21710 ( .A(n18612), .ZN(n18613) );
  AOI22_X1 U21711 ( .A1(P3_REQUESTPENDING_REG_SCAN_IN), .A2(n18614), .B1(HOLD), 
        .B2(n18613), .ZN(n18616) );
  NAND2_X1 U21712 ( .A1(n18615), .A2(P3_STATE_REG_1__SCAN_IN), .ZN(n18619) );
  OAI211_X1 U21713 ( .C1(n18616), .C2(n18623), .A(n18619), .B(n18744), .ZN(
        P3_U3030) );
  INV_X1 U21714 ( .A(n18619), .ZN(n18617) );
  AOI21_X1 U21715 ( .B1(n18623), .B2(n18618), .A(n18617), .ZN(n18624) );
  OAI22_X1 U21716 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(
        P3_REQUESTPENDING_REG_SCAN_IN), .B1(NA), .B2(n18619), .ZN(n18620) );
  OAI22_X1 U21717 ( .A1(n18621), .A2(n18620), .B1(
        P3_REQUESTPENDING_REG_SCAN_IN), .B2(HOLD), .ZN(n18622) );
  OAI22_X1 U21718 ( .A1(n18624), .A2(n18625), .B1(n18623), .B2(n18622), .ZN(
        P3_U3031) );
  INV_X1 U21719 ( .A(n18755), .ZN(n18754) );
  INV_X1 U21720 ( .A(P3_REIP_REG_2__SCAN_IN), .ZN(n18627) );
  OAI222_X1 U21721 ( .A1(n18729), .A2(n18680), .B1(n18626), .B2(n18754), .C1(
        n18627), .C2(n18685), .ZN(P3_U3032) );
  OAI222_X1 U21722 ( .A1(n18685), .A2(n18629), .B1(n18628), .B2(n18682), .C1(
        n18627), .C2(n18680), .ZN(P3_U3033) );
  OAI222_X1 U21723 ( .A1(n18685), .A2(n18631), .B1(n18630), .B2(n18754), .C1(
        n18629), .C2(n18680), .ZN(P3_U3034) );
  OAI222_X1 U21724 ( .A1(n18685), .A2(n18634), .B1(n18632), .B2(n18682), .C1(
        n18631), .C2(n18680), .ZN(P3_U3035) );
  OAI222_X1 U21725 ( .A1(n18634), .A2(n18680), .B1(n18633), .B2(n18754), .C1(
        n21078), .C2(n18685), .ZN(P3_U3036) );
  OAI222_X1 U21726 ( .A1(n21078), .A2(n18680), .B1(n18635), .B2(n18754), .C1(
        n18636), .C2(n18685), .ZN(P3_U3037) );
  OAI222_X1 U21727 ( .A1(n18685), .A2(n18638), .B1(n18637), .B2(n18682), .C1(
        n18636), .C2(n18680), .ZN(P3_U3038) );
  OAI222_X1 U21728 ( .A1(n18685), .A2(n18640), .B1(n18639), .B2(n18754), .C1(
        n18638), .C2(n18680), .ZN(P3_U3039) );
  OAI222_X1 U21729 ( .A1(n18685), .A2(n18641), .B1(n21104), .B2(n18754), .C1(
        n18640), .C2(n18680), .ZN(P3_U3040) );
  INV_X1 U21730 ( .A(P3_REIP_REG_11__SCAN_IN), .ZN(n18643) );
  OAI222_X1 U21731 ( .A1(n18685), .A2(n18643), .B1(n18642), .B2(n18754), .C1(
        n18641), .C2(n18680), .ZN(P3_U3041) );
  OAI222_X1 U21732 ( .A1(n18685), .A2(n18645), .B1(n18644), .B2(n18754), .C1(
        n18643), .C2(n18680), .ZN(P3_U3042) );
  OAI222_X1 U21733 ( .A1(n18685), .A2(n18647), .B1(n18646), .B2(n18754), .C1(
        n18645), .C2(n18680), .ZN(P3_U3043) );
  OAI222_X1 U21734 ( .A1(n18685), .A2(n18649), .B1(n18648), .B2(n18754), .C1(
        n18647), .C2(n18680), .ZN(P3_U3044) );
  OAI222_X1 U21735 ( .A1(n18685), .A2(n18651), .B1(n18650), .B2(n18754), .C1(
        n18649), .C2(n18680), .ZN(P3_U3045) );
  INV_X1 U21736 ( .A(P3_REIP_REG_16__SCAN_IN), .ZN(n18653) );
  OAI222_X1 U21737 ( .A1(n18685), .A2(n18653), .B1(n18652), .B2(n18754), .C1(
        n18651), .C2(n18680), .ZN(P3_U3046) );
  OAI222_X1 U21738 ( .A1(n18685), .A2(n18655), .B1(n18654), .B2(n18754), .C1(
        n18653), .C2(n18680), .ZN(P3_U3047) );
  OAI222_X1 U21739 ( .A1(n18685), .A2(n18657), .B1(n18656), .B2(n18754), .C1(
        n18655), .C2(n18680), .ZN(P3_U3048) );
  OAI222_X1 U21740 ( .A1(n18685), .A2(n18659), .B1(n18658), .B2(n18754), .C1(
        n18657), .C2(n18680), .ZN(P3_U3049) );
  INV_X1 U21741 ( .A(P3_REIP_REG_20__SCAN_IN), .ZN(n18661) );
  OAI222_X1 U21742 ( .A1(n18685), .A2(n18661), .B1(n18660), .B2(n18754), .C1(
        n18659), .C2(n18680), .ZN(P3_U3050) );
  OAI222_X1 U21743 ( .A1(n18685), .A2(n18663), .B1(n18662), .B2(n18754), .C1(
        n18661), .C2(n18680), .ZN(P3_U3051) );
  OAI222_X1 U21744 ( .A1(n18685), .A2(n18665), .B1(n18664), .B2(n18754), .C1(
        n18663), .C2(n18680), .ZN(P3_U3052) );
  OAI222_X1 U21745 ( .A1(n18685), .A2(n20919), .B1(n18666), .B2(n18754), .C1(
        n18665), .C2(n18680), .ZN(P3_U3053) );
  OAI222_X1 U21746 ( .A1(n18685), .A2(n18669), .B1(n18667), .B2(n18682), .C1(
        n20919), .C2(n18680), .ZN(P3_U3054) );
  OAI222_X1 U21747 ( .A1(n18669), .A2(n18680), .B1(n18668), .B2(n18682), .C1(
        n18670), .C2(n18685), .ZN(P3_U3055) );
  OAI222_X1 U21748 ( .A1(n18685), .A2(n18672), .B1(n18671), .B2(n18682), .C1(
        n18670), .C2(n18680), .ZN(P3_U3056) );
  OAI222_X1 U21749 ( .A1(n18685), .A2(n18675), .B1(n18673), .B2(n18682), .C1(
        n18672), .C2(n18680), .ZN(P3_U3057) );
  OAI222_X1 U21750 ( .A1(n18680), .A2(n18675), .B1(n18674), .B2(n18682), .C1(
        n18676), .C2(n18685), .ZN(P3_U3058) );
  INV_X1 U21751 ( .A(P3_ADDRESS_REG_27__SCAN_IN), .ZN(n18677) );
  OAI222_X1 U21752 ( .A1(n18685), .A2(n18678), .B1(n18677), .B2(n18682), .C1(
        n18676), .C2(n18680), .ZN(P3_U3059) );
  OAI222_X1 U21753 ( .A1(n18685), .A2(n18681), .B1(n18679), .B2(n18682), .C1(
        n18678), .C2(n18680), .ZN(P3_U3060) );
  OAI222_X1 U21754 ( .A1(n18685), .A2(n18684), .B1(n18683), .B2(n18682), .C1(
        n18681), .C2(n18680), .ZN(P3_U3061) );
  OAI22_X1 U21755 ( .A1(n18755), .A2(P3_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P3_BE_N_REG_3__SCAN_IN), .B2(n18754), .ZN(n18686) );
  INV_X1 U21756 ( .A(n18686), .ZN(P3_U3274) );
  OAI22_X1 U21757 ( .A1(n18755), .A2(P3_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P3_BE_N_REG_2__SCAN_IN), .B2(n18754), .ZN(n18687) );
  INV_X1 U21758 ( .A(n18687), .ZN(P3_U3275) );
  OAI22_X1 U21759 ( .A1(n18755), .A2(P3_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P3_BE_N_REG_1__SCAN_IN), .B2(n18754), .ZN(n18688) );
  INV_X1 U21760 ( .A(n18688), .ZN(P3_U3276) );
  OAI22_X1 U21761 ( .A1(n18755), .A2(P3_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P3_BE_N_REG_0__SCAN_IN), .B2(n18682), .ZN(n18689) );
  INV_X1 U21762 ( .A(n18689), .ZN(P3_U3277) );
  OAI21_X1 U21763 ( .B1(n18693), .B2(P3_DATAWIDTH_REG_0__SCAN_IN), .A(n18691), 
        .ZN(n18690) );
  INV_X1 U21764 ( .A(n18690), .ZN(P3_U3280) );
  OAI21_X1 U21765 ( .B1(n18693), .B2(n18692), .A(n18691), .ZN(P3_U3281) );
  OAI221_X1 U21766 ( .B1(n18696), .B2(P3_STATE2_REG_0__SCAN_IN), .C1(n18696), 
        .C2(n18695), .A(n18694), .ZN(P3_U3282) );
  INV_X1 U21767 ( .A(n18697), .ZN(n18700) );
  NOR3_X1 U21768 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18698), .A3(
        n18757), .ZN(n18699) );
  AOI21_X1 U21769 ( .B1(n18721), .B2(n18700), .A(n18699), .ZN(n18704) );
  INV_X1 U21770 ( .A(n18728), .ZN(n18725) );
  OAI21_X1 U21771 ( .B1(n18757), .B2(n18701), .A(n18725), .ZN(n18702) );
  INV_X1 U21772 ( .A(n18702), .ZN(n18703) );
  OAI22_X1 U21773 ( .A1(n18728), .A2(n18704), .B1(n18703), .B2(n11640), .ZN(
        P3_U3285) );
  INV_X1 U21774 ( .A(n18705), .ZN(n18711) );
  NOR2_X1 U21775 ( .A1(n18706), .A2(n18724), .ZN(n18715) );
  OAI22_X1 U21776 ( .A1(n18708), .A2(n18707), .B1(
        P3_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(
        P3_INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n18716) );
  INV_X1 U21777 ( .A(n18716), .ZN(n18710) );
  AOI222_X1 U21778 ( .A1(n18711), .A2(n18723), .B1(n18715), .B2(n18710), .C1(
        n18721), .C2(n18709), .ZN(n18712) );
  AOI22_X1 U21779 ( .A1(n18728), .A2(n18713), .B1(n18712), .B2(n18725), .ZN(
        P3_U3288) );
  INV_X1 U21780 ( .A(n18714), .ZN(n18717) );
  AOI222_X1 U21781 ( .A1(n18718), .A2(n18723), .B1(n18721), .B2(n18717), .C1(
        n18716), .C2(n18715), .ZN(n18719) );
  AOI22_X1 U21782 ( .A1(n18728), .A2(n18720), .B1(n18719), .B2(n18725), .ZN(
        P3_U3289) );
  AOI222_X1 U21783 ( .A1(n18724), .A2(P3_STATE2_REG_1__SCAN_IN), .B1(n18723), 
        .B2(n18722), .C1(n18727), .C2(n18721), .ZN(n18726) );
  AOI22_X1 U21784 ( .A1(n18728), .A2(n18727), .B1(n18726), .B2(n18725), .ZN(
        P3_U3290) );
  AOI21_X1 U21785 ( .B1(P3_REIP_REG_0__SCAN_IN), .B2(
        P3_DATAWIDTH_REG_0__SCAN_IN), .A(P3_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n18730) );
  AOI22_X1 U21786 ( .A1(P3_REIP_REG_1__SCAN_IN), .A2(P3_REIP_REG_0__SCAN_IN), 
        .B1(n18730), .B2(n18729), .ZN(n18733) );
  INV_X1 U21787 ( .A(P3_BYTEENABLE_REG_2__SCAN_IN), .ZN(n18732) );
  AOI22_X1 U21788 ( .A1(n18736), .A2(n18733), .B1(n18732), .B2(n18731), .ZN(
        P3_U3292) );
  INV_X1 U21789 ( .A(P3_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18735) );
  OAI21_X1 U21790 ( .B1(P3_REIP_REG_1__SCAN_IN), .B2(P3_REIP_REG_0__SCAN_IN), 
        .A(n18736), .ZN(n18734) );
  OAI21_X1 U21791 ( .B1(n18736), .B2(n18735), .A(n18734), .ZN(P3_U3293) );
  INV_X1 U21792 ( .A(P3_W_R_N_REG_SCAN_IN), .ZN(n18737) );
  AOI22_X1 U21793 ( .A1(n18754), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18737), 
        .B2(n18755), .ZN(P3_U3294) );
  MUX2_X1 U21794 ( .A(P3_MORE_REG_SCAN_IN), .B(n18739), .S(n18738), .Z(
        P3_U3295) );
  OAI21_X1 U21795 ( .B1(n18741), .B2(n18740), .A(n18759), .ZN(n18742) );
  AOI21_X1 U21796 ( .B1(n18743), .B2(n18747), .A(n18742), .ZN(n18753) );
  AOI21_X1 U21797 ( .B1(n18746), .B2(n18745), .A(n18744), .ZN(n18748) );
  OAI211_X1 U21798 ( .C1(n18758), .C2(n18748), .A(P3_STATE2_REG_2__SCAN_IN), 
        .B(n18747), .ZN(n18750) );
  AOI21_X1 U21799 ( .B1(P3_STATE2_REG_0__SCAN_IN), .B2(n18750), .A(n18749), 
        .ZN(n18752) );
  NAND2_X1 U21800 ( .A1(n18753), .A2(P3_REQUESTPENDING_REG_SCAN_IN), .ZN(
        n18751) );
  OAI21_X1 U21801 ( .B1(n18753), .B2(n18752), .A(n18751), .ZN(P3_U3296) );
  OAI22_X1 U21802 ( .A1(n18755), .A2(P3_MEMORYFETCH_REG_SCAN_IN), .B1(
        P3_M_IO_N_REG_SCAN_IN), .B2(n18754), .ZN(n18756) );
  INV_X1 U21803 ( .A(n18756), .ZN(P3_U3297) );
  OAI21_X1 U21804 ( .B1(n18757), .B2(P3_STATE2_REG_2__SCAN_IN), .A(n18759), 
        .ZN(n18762) );
  OAI22_X1 U21805 ( .A1(n18762), .A2(P3_READREQUEST_REG_SCAN_IN), .B1(n18759), 
        .B2(n18758), .ZN(n18760) );
  INV_X1 U21806 ( .A(n18760), .ZN(P3_U3298) );
  OAI21_X1 U21807 ( .B1(n18762), .B2(P3_MEMORYFETCH_REG_SCAN_IN), .A(n18761), 
        .ZN(n18763) );
  INV_X1 U21808 ( .A(n18763), .ZN(P3_U3299) );
  INV_X1 U21809 ( .A(P2_STATE_REG_0__SCAN_IN), .ZN(n18768) );
  NAND2_X1 U21810 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19735), .ZN(n19725) );
  NAND2_X1 U21811 ( .A1(n18768), .A2(n18764), .ZN(n19722) );
  OAI21_X1 U21812 ( .B1(n18768), .B2(n19725), .A(n19722), .ZN(n19783) );
  AOI21_X1 U21813 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(P2_ADS_N_REG_SCAN_IN), 
        .A(n19783), .ZN(n18765) );
  INV_X1 U21814 ( .A(n18765), .ZN(P2_U2815) );
  INV_X1 U21815 ( .A(P2_CODEFETCH_REG_SCAN_IN), .ZN(n18767) );
  OAI22_X1 U21816 ( .A1(n19847), .A2(n18767), .B1(n10983), .B2(n18766), .ZN(
        P2_U2816) );
  NAND2_X1 U21817 ( .A1(n18768), .A2(P2_STATE_REG_1__SCAN_IN), .ZN(n19854) );
  AOI21_X1 U21818 ( .B1(n18768), .B2(n19735), .A(P2_D_C_N_REG_SCAN_IN), .ZN(
        n18769) );
  AOI22_X1 U21819 ( .A1(n19853), .A2(P2_CODEFETCH_REG_SCAN_IN), .B1(n18769), 
        .B2(n19854), .ZN(P2_U2817) );
  OAI21_X1 U21820 ( .B1(n19728), .B2(BS16), .A(n19783), .ZN(n19781) );
  OAI21_X1 U21821 ( .B1(n19783), .B2(n19836), .A(n19781), .ZN(P2_U2818) );
  NOR4_X1 U21822 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_9__SCAN_IN), .A3(P2_DATAWIDTH_REG_10__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_11__SCAN_IN), .ZN(n18779) );
  NOR4_X1 U21823 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_5__SCAN_IN), .A3(P2_DATAWIDTH_REG_6__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_7__SCAN_IN), .ZN(n18778) );
  AOI211_X1 U21824 ( .C1(P2_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P2_DATAWIDTH_REG_0__SCAN_IN), .A(P2_DATAWIDTH_REG_24__SCAN_IN), .B(
        P2_DATAWIDTH_REG_2__SCAN_IN), .ZN(n18770) );
  INV_X1 U21825 ( .A(P2_DATAWIDTH_REG_4__SCAN_IN), .ZN(n20921) );
  INV_X1 U21826 ( .A(P2_DATAWIDTH_REG_18__SCAN_IN), .ZN(n21068) );
  NAND3_X1 U21827 ( .A1(n18770), .A2(n20921), .A3(n21068), .ZN(n18776) );
  NOR4_X1 U21828 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_19__SCAN_IN), .A3(P2_DATAWIDTH_REG_20__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_22__SCAN_IN), .ZN(n18774) );
  NOR4_X1 U21829 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_13__SCAN_IN), .A3(P2_DATAWIDTH_REG_15__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_16__SCAN_IN), .ZN(n18773) );
  NOR4_X1 U21830 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_29__SCAN_IN), .A3(P2_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_31__SCAN_IN), .ZN(n18772) );
  NOR4_X1 U21831 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_25__SCAN_IN), .A3(P2_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P2_DATAWIDTH_REG_27__SCAN_IN), .ZN(n18771) );
  NAND4_X1 U21832 ( .A1(n18774), .A2(n18773), .A3(n18772), .A4(n18771), .ZN(
        n18775) );
  NOR4_X1 U21833 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(
        P2_DATAWIDTH_REG_21__SCAN_IN), .A3(n18776), .A4(n18775), .ZN(n18777)
         );
  NAND3_X1 U21834 ( .A1(n18779), .A2(n18778), .A3(n18777), .ZN(n18787) );
  NOR2_X1 U21835 ( .A1(P2_REIP_REG_1__SCAN_IN), .A2(n18787), .ZN(n18782) );
  INV_X1 U21836 ( .A(P2_BYTEENABLE_REG_0__SCAN_IN), .ZN(n18780) );
  AOI22_X1 U21837 ( .A1(n18782), .A2(n18955), .B1(n18787), .B2(n18780), .ZN(
        P2_U2820) );
  OR3_X1 U21838 ( .A1(P2_REIP_REG_0__SCAN_IN), .A2(P2_DATAWIDTH_REG_1__SCAN_IN), .A3(P2_DATAWIDTH_REG_0__SCAN_IN), .ZN(n18786) );
  INV_X1 U21839 ( .A(P2_BYTEENABLE_REG_1__SCAN_IN), .ZN(n18781) );
  AOI22_X1 U21840 ( .A1(n18782), .A2(n18786), .B1(n18787), .B2(n18781), .ZN(
        P2_U2821) );
  INV_X1 U21841 ( .A(P2_DATAWIDTH_REG_1__SCAN_IN), .ZN(n19782) );
  NAND2_X1 U21842 ( .A1(n18782), .A2(n19782), .ZN(n18785) );
  INV_X1 U21843 ( .A(n18787), .ZN(n18789) );
  OAI21_X1 U21844 ( .B1(n10425), .B2(n18955), .A(n18789), .ZN(n18783) );
  OAI21_X1 U21845 ( .B1(P2_BYTEENABLE_REG_2__SCAN_IN), .B2(n18789), .A(n18783), 
        .ZN(n18784) );
  OAI221_X1 U21846 ( .B1(n18785), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .C1(n18785), .C2(P2_REIP_REG_0__SCAN_IN), .A(n18784), .ZN(P2_U2822) );
  INV_X1 U21847 ( .A(P2_BYTEENABLE_REG_3__SCAN_IN), .ZN(n18788) );
  OAI221_X1 U21848 ( .B1(n18789), .B2(n18788), .C1(n18787), .C2(n18786), .A(
        n18785), .ZN(P2_U2823) );
  NAND2_X1 U21849 ( .A1(n18929), .A2(n18790), .ZN(n18791) );
  XOR2_X1 U21850 ( .A(n18792), .B(n18791), .Z(n18803) );
  OAI21_X1 U21851 ( .B1(n19754), .B2(n18954), .A(n18934), .ZN(n18796) );
  OAI22_X1 U21852 ( .A1(n18794), .A2(n18947), .B1(n18831), .B2(n18793), .ZN(
        n18795) );
  AOI211_X1 U21853 ( .C1(P2_EBX_REG_19__SCAN_IN), .C2(n18951), .A(n18796), .B(
        n18795), .ZN(n18802) );
  INV_X1 U21854 ( .A(n18797), .ZN(n18798) );
  OAI22_X1 U21855 ( .A1(n18799), .A2(n18937), .B1(n18798), .B2(n18945), .ZN(
        n18800) );
  INV_X1 U21856 ( .A(n18800), .ZN(n18801) );
  OAI211_X1 U21857 ( .C1(n19714), .C2(n18803), .A(n18802), .B(n18801), .ZN(
        P2_U2836) );
  NOR2_X1 U21858 ( .A1(n18917), .A2(n18804), .ZN(n18806) );
  XOR2_X1 U21859 ( .A(n18806), .B(n18805), .Z(n18815) );
  AOI22_X1 U21860 ( .A1(n18951), .A2(P2_EBX_REG_18__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n18958), .ZN(n18807) );
  OAI21_X1 U21861 ( .B1(n18808), .B2(n18947), .A(n18807), .ZN(n18809) );
  AOI211_X1 U21862 ( .C1(P2_REIP_REG_18__SCAN_IN), .C2(n18885), .A(n19085), 
        .B(n18809), .ZN(n18814) );
  OAI22_X1 U21863 ( .A1(n18811), .A2(n18937), .B1(n18810), .B2(n18945), .ZN(
        n18812) );
  INV_X1 U21864 ( .A(n18812), .ZN(n18813) );
  OAI211_X1 U21865 ( .C1(n19714), .C2(n18815), .A(n18814), .B(n18813), .ZN(
        P2_U2837) );
  NAND2_X1 U21866 ( .A1(n18929), .A2(n18816), .ZN(n18817) );
  XOR2_X1 U21867 ( .A(n18818), .B(n18817), .Z(n18827) );
  OAI21_X1 U21868 ( .B1(n19750), .B2(n18954), .A(n18934), .ZN(n18822) );
  OAI22_X1 U21869 ( .A1(n18820), .A2(n18947), .B1(n18831), .B2(n18819), .ZN(
        n18821) );
  AOI211_X1 U21870 ( .C1(P2_EBX_REG_17__SCAN_IN), .C2(n18951), .A(n18822), .B(
        n18821), .ZN(n18826) );
  AOI22_X1 U21871 ( .A1(n18824), .A2(n18949), .B1(n18823), .B2(n18877), .ZN(
        n18825) );
  OAI211_X1 U21872 ( .C1(n19714), .C2(n18827), .A(n18826), .B(n18825), .ZN(
        P2_U2838) );
  NOR2_X1 U21873 ( .A1(n18917), .A2(n18828), .ZN(n18830) );
  XOR2_X1 U21874 ( .A(n18830), .B(n18829), .Z(n18839) );
  OAI21_X1 U21875 ( .B1(n15415), .B2(n18954), .A(n18934), .ZN(n18834) );
  OAI22_X1 U21876 ( .A1(n18832), .A2(n18947), .B1(n18831), .B2(n10090), .ZN(
        n18833) );
  AOI211_X1 U21877 ( .C1(P2_EBX_REG_16__SCAN_IN), .C2(n18951), .A(n18834), .B(
        n18833), .ZN(n18838) );
  OAI22_X1 U21878 ( .A1(n18835), .A2(n18937), .B1(n18968), .B2(n18945), .ZN(
        n18836) );
  INV_X1 U21879 ( .A(n18836), .ZN(n18837) );
  OAI211_X1 U21880 ( .C1(n19714), .C2(n18839), .A(n18838), .B(n18837), .ZN(
        P2_U2839) );
  OAI21_X1 U21881 ( .B1(n19747), .B2(n18954), .A(n18934), .ZN(n18843) );
  OAI22_X1 U21882 ( .A1(n18841), .A2(n18947), .B1(n18840), .B2(n21015), .ZN(
        n18842) );
  AOI211_X1 U21883 ( .C1(P2_PHYADDRPOINTER_REG_15__SCAN_IN), .C2(n18958), .A(
        n18843), .B(n18842), .ZN(n18850) );
  NAND2_X1 U21884 ( .A1(n18929), .A2(n18844), .ZN(n18845) );
  XOR2_X1 U21885 ( .A(n18846), .B(n18845), .Z(n18848) );
  AOI22_X1 U21886 ( .A1(n18848), .A2(n18890), .B1(n18847), .B2(n18949), .ZN(
        n18849) );
  OAI211_X1 U21887 ( .C1(n18851), .C2(n18945), .A(n18850), .B(n18849), .ZN(
        P2_U2840) );
  AOI211_X1 U21888 ( .C1(n18863), .C2(n18854), .A(n18853), .B(n18852), .ZN(
        n18861) );
  NAND2_X1 U21889 ( .A1(n18855), .A2(n18933), .ZN(n18859) );
  AOI22_X1 U21890 ( .A1(P2_EBX_REG_13__SCAN_IN), .A2(n18951), .B1(
        P2_PHYADDRPOINTER_REG_13__SCAN_IN), .B2(n18958), .ZN(n18856) );
  OAI211_X1 U21891 ( .C1(n18954), .C2(n12793), .A(n18856), .B(n18934), .ZN(
        n18857) );
  INV_X1 U21892 ( .A(n18857), .ZN(n18858) );
  NAND2_X1 U21893 ( .A1(n18859), .A2(n18858), .ZN(n18860) );
  NOR2_X1 U21894 ( .A1(n18861), .A2(n18860), .ZN(n18866) );
  AOI22_X1 U21895 ( .A1(n18864), .A2(n18863), .B1(n18862), .B2(n18949), .ZN(
        n18865) );
  OAI211_X1 U21896 ( .C1(n18867), .C2(n18945), .A(n18866), .B(n18865), .ZN(
        P2_U2842) );
  NOR2_X1 U21897 ( .A1(n18917), .A2(n18868), .ZN(n18870) );
  XOR2_X1 U21898 ( .A(n18870), .B(n18869), .Z(n18881) );
  AOI22_X1 U21899 ( .A1(n18951), .A2(P2_EBX_REG_12__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_12__SCAN_IN), .B2(n18958), .ZN(n18871) );
  OAI21_X1 U21900 ( .B1(n18872), .B2(n18947), .A(n18871), .ZN(n18873) );
  AOI211_X1 U21901 ( .C1(P2_REIP_REG_12__SCAN_IN), .C2(n18885), .A(n19085), 
        .B(n18873), .ZN(n18880) );
  INV_X1 U21902 ( .A(n18874), .ZN(n18878) );
  INV_X1 U21903 ( .A(n18875), .ZN(n18876) );
  AOI22_X1 U21904 ( .A1(n18878), .A2(n18949), .B1(n18877), .B2(n18876), .ZN(
        n18879) );
  OAI211_X1 U21905 ( .C1(n19714), .C2(n18881), .A(n18880), .B(n18879), .ZN(
        P2_U2843) );
  AOI22_X1 U21906 ( .A1(n18951), .A2(P2_EBX_REG_11__SCAN_IN), .B1(
        P2_PHYADDRPOINTER_REG_11__SCAN_IN), .B2(n18958), .ZN(n18882) );
  OAI21_X1 U21907 ( .B1(n18883), .B2(n18947), .A(n18882), .ZN(n18884) );
  AOI211_X1 U21908 ( .C1(P2_REIP_REG_11__SCAN_IN), .C2(n18885), .A(n19085), 
        .B(n18884), .ZN(n18893) );
  NAND2_X1 U21909 ( .A1(n18929), .A2(n18886), .ZN(n18887) );
  XNOR2_X1 U21910 ( .A(n18888), .B(n18887), .ZN(n18891) );
  AOI22_X1 U21911 ( .A1(n18891), .A2(n18890), .B1(n18889), .B2(n18949), .ZN(
        n18892) );
  OAI211_X1 U21912 ( .C1(n18894), .C2(n18945), .A(n18893), .B(n18892), .ZN(
        P2_U2844) );
  NOR2_X1 U21913 ( .A1(n18917), .A2(n18895), .ZN(n18896) );
  XOR2_X1 U21914 ( .A(n18897), .B(n18896), .Z(n18904) );
  AOI22_X1 U21915 ( .A1(n18898), .A2(n18933), .B1(
        P2_PHYADDRPOINTER_REG_10__SCAN_IN), .B2(n18958), .ZN(n18899) );
  OAI211_X1 U21916 ( .C1(n12751), .C2(n18954), .A(n18899), .B(n18934), .ZN(
        n18902) );
  OAI22_X1 U21917 ( .A1(n18981), .A2(n18945), .B1(n18900), .B2(n18937), .ZN(
        n18901) );
  AOI211_X1 U21918 ( .C1(P2_EBX_REG_10__SCAN_IN), .C2(n18951), .A(n18902), .B(
        n18901), .ZN(n18903) );
  OAI21_X1 U21919 ( .B1(n19714), .B2(n18904), .A(n18903), .ZN(P2_U2845) );
  NAND2_X1 U21920 ( .A1(n18929), .A2(n18905), .ZN(n18907) );
  XOR2_X1 U21921 ( .A(n18907), .B(n18906), .Z(n18915) );
  AOI22_X1 U21922 ( .A1(n18908), .A2(n18933), .B1(P2_EBX_REG_7__SCAN_IN), .B2(
        n18951), .ZN(n18909) );
  OAI211_X1 U21923 ( .C1(n10916), .C2(n18954), .A(n18909), .B(n18934), .ZN(
        n18913) );
  OAI22_X1 U21924 ( .A1(n18911), .A2(n18945), .B1(n18910), .B2(n18937), .ZN(
        n18912) );
  AOI211_X1 U21925 ( .C1(P2_PHYADDRPOINTER_REG_7__SCAN_IN), .C2(n18958), .A(
        n18913), .B(n18912), .ZN(n18914) );
  OAI21_X1 U21926 ( .B1(n18915), .B2(n19714), .A(n18914), .ZN(P2_U2848) );
  NOR2_X1 U21927 ( .A1(n18917), .A2(n18916), .ZN(n18918) );
  XOR2_X1 U21928 ( .A(n18919), .B(n18918), .Z(n18927) );
  AOI22_X1 U21929 ( .A1(n18920), .A2(n18933), .B1(
        P2_PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n18958), .ZN(n18921) );
  OAI211_X1 U21930 ( .C1(n10912), .C2(n18954), .A(n18921), .B(n18934), .ZN(
        n18925) );
  OAI22_X1 U21931 ( .A1(n18923), .A2(n18945), .B1(n18922), .B2(n18937), .ZN(
        n18924) );
  AOI211_X1 U21932 ( .C1(P2_EBX_REG_6__SCAN_IN), .C2(n18951), .A(n18925), .B(
        n18924), .ZN(n18926) );
  OAI21_X1 U21933 ( .B1(n19714), .B2(n18927), .A(n18926), .ZN(P2_U2849) );
  NAND2_X1 U21934 ( .A1(n18929), .A2(n18928), .ZN(n18931) );
  XOR2_X1 U21935 ( .A(n18931), .B(n18930), .Z(n18941) );
  AOI22_X1 U21936 ( .A1(n18933), .A2(n18932), .B1(n18951), .B2(
        P2_EBX_REG_5__SCAN_IN), .ZN(n18935) );
  OAI211_X1 U21937 ( .C1(n10904), .C2(n18954), .A(n18935), .B(n18934), .ZN(
        n18939) );
  OAI22_X1 U21938 ( .A1(n18994), .A2(n18945), .B1(n18937), .B2(n18936), .ZN(
        n18938) );
  AOI211_X1 U21939 ( .C1(P2_PHYADDRPOINTER_REG_5__SCAN_IN), .C2(n18958), .A(
        n18939), .B(n18938), .ZN(n18940) );
  OAI21_X1 U21940 ( .B1(n18941), .B2(n19714), .A(n18940), .ZN(P2_U2850) );
  INV_X1 U21941 ( .A(n18943), .ZN(n18946) );
  OAI22_X1 U21942 ( .A1(n18947), .A2(n18946), .B1(n18945), .B2(n18944), .ZN(
        n18948) );
  AOI21_X1 U21943 ( .B1(n18950), .B2(n18949), .A(n18948), .ZN(n18953) );
  NAND2_X1 U21944 ( .A1(n18951), .A2(P2_EBX_REG_0__SCAN_IN), .ZN(n18952) );
  OAI211_X1 U21945 ( .C1(n18955), .C2(n18954), .A(n18953), .B(n18952), .ZN(
        n18956) );
  AOI21_X1 U21946 ( .B1(n18957), .B2(n19158), .A(n18956), .ZN(n18960) );
  NAND2_X1 U21947 ( .A1(P2_PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n18958), .ZN(
        n18959) );
  OAI211_X1 U21948 ( .C1(n14927), .C2(n19714), .A(n18960), .B(n18959), .ZN(
        P2_U2855) );
  AOI22_X1 U21949 ( .A1(n18966), .A2(BUF2_REG_31__SCAN_IN), .B1(n19005), .B2(
        n18961), .ZN(n18963) );
  AOI22_X1 U21950 ( .A1(n18967), .A2(BUF1_REG_31__SCAN_IN), .B1(
        P2_EAX_REG_31__SCAN_IN), .B2(n19004), .ZN(n18962) );
  NAND2_X1 U21951 ( .A1(n18963), .A2(n18962), .ZN(P2_U2888) );
  INV_X1 U21952 ( .A(n19115), .ZN(n18964) );
  AOI22_X1 U21953 ( .A1(n18965), .A2(n18964), .B1(P2_EAX_REG_16__SCAN_IN), 
        .B2(n19004), .ZN(n18974) );
  AOI22_X1 U21954 ( .A1(n18967), .A2(BUF1_REG_16__SCAN_IN), .B1(n18966), .B2(
        BUF2_REG_16__SCAN_IN), .ZN(n18973) );
  OAI22_X1 U21955 ( .A1(n18970), .A2(n19009), .B1(n18969), .B2(n18968), .ZN(
        n18971) );
  INV_X1 U21956 ( .A(n18971), .ZN(n18972) );
  NAND3_X1 U21957 ( .A1(n18974), .A2(n18973), .A3(n18972), .ZN(P2_U2903) );
  INV_X1 U21958 ( .A(n18975), .ZN(n18978) );
  AOI22_X1 U21959 ( .A1(n18989), .A2(n18976), .B1(P2_EAX_REG_14__SCAN_IN), 
        .B2(n19004), .ZN(n18977) );
  OAI21_X1 U21960 ( .B1(n18995), .B2(n18978), .A(n18977), .ZN(P2_U2905) );
  AOI22_X1 U21961 ( .A1(n18989), .A2(n18979), .B1(P2_EAX_REG_10__SCAN_IN), 
        .B2(n19004), .ZN(n18980) );
  OAI21_X1 U21962 ( .B1(n18995), .B2(n18981), .A(n18980), .ZN(P2_U2909) );
  AOI22_X1 U21963 ( .A1(n18989), .A2(n18982), .B1(P2_EAX_REG_9__SCAN_IN), .B2(
        n19004), .ZN(n18983) );
  OAI21_X1 U21964 ( .B1(n18995), .B2(n18984), .A(n18983), .ZN(P2_U2910) );
  AOI22_X1 U21965 ( .A1(n18989), .A2(n18985), .B1(P2_EAX_REG_8__SCAN_IN), .B2(
        n19004), .ZN(n18986) );
  OAI21_X1 U21966 ( .B1(n18995), .B2(n18987), .A(n18986), .ZN(P2_U2911) );
  INV_X1 U21967 ( .A(n19135), .ZN(n18988) );
  AOI22_X1 U21968 ( .A1(n18989), .A2(n18988), .B1(P2_EAX_REG_5__SCAN_IN), .B2(
        n19004), .ZN(n18993) );
  OR3_X1 U21969 ( .A1(n18991), .A2(n18990), .A3(n19009), .ZN(n18992) );
  OAI211_X1 U21970 ( .C1(n18995), .C2(n18994), .A(n18993), .B(n18992), .ZN(
        P2_U2914) );
  INV_X1 U21971 ( .A(n18996), .ZN(n19794) );
  AOI22_X1 U21972 ( .A1(n19794), .A2(n19005), .B1(P2_EAX_REG_3__SCAN_IN), .B2(
        n19004), .ZN(n19002) );
  AOI21_X1 U21973 ( .B1(n18999), .B2(n18998), .A(n18997), .ZN(n19000) );
  OR2_X1 U21974 ( .A1(n19000), .A2(n19009), .ZN(n19001) );
  OAI211_X1 U21975 ( .C1(n19130), .C2(n19013), .A(n19002), .B(n19001), .ZN(
        P2_U2916) );
  INV_X1 U21976 ( .A(n19003), .ZN(n19812) );
  AOI22_X1 U21977 ( .A1(n19005), .A2(n19812), .B1(n19004), .B2(
        P2_EAX_REG_1__SCAN_IN), .ZN(n19012) );
  AOI21_X1 U21978 ( .B1(n19008), .B2(n19007), .A(n19006), .ZN(n19010) );
  OR2_X1 U21979 ( .A1(n19010), .A2(n19009), .ZN(n19011) );
  OAI211_X1 U21980 ( .C1(n19119), .C2(n19013), .A(n19012), .B(n19011), .ZN(
        P2_U2918) );
  OAI21_X1 U21981 ( .B1(n19015), .B2(n19014), .A(n13452), .ZN(n19016) );
  NOR2_X1 U21982 ( .A1(P2_STATE2_REG_0__SCAN_IN), .A2(n19815), .ZN(n19056) );
  CLKBUF_X1 U21983 ( .A(n19056), .Z(n19850) );
  NOR2_X1 U21984 ( .A1(n19059), .A2(n19017), .ZN(P2_U2920) );
  NAND2_X1 U21985 ( .A1(n19057), .A2(n19835), .ZN(n19046) );
  AOI22_X1 U21986 ( .A1(n19850), .A2(P2_UWORD_REG_14__SCAN_IN), .B1(
        P2_DATAO_REG_30__SCAN_IN), .B2(n19076), .ZN(n19018) );
  OAI21_X1 U21987 ( .B1(n19019), .B2(n19046), .A(n19018), .ZN(P2_U2921) );
  AOI22_X1 U21988 ( .A1(n19056), .A2(P2_UWORD_REG_13__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_29__SCAN_IN), .ZN(n19020) );
  OAI21_X1 U21989 ( .B1(n19021), .B2(n19046), .A(n19020), .ZN(P2_U2922) );
  AOI22_X1 U21990 ( .A1(n19056), .A2(P2_UWORD_REG_12__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_28__SCAN_IN), .ZN(n19022) );
  OAI21_X1 U21991 ( .B1(n19023), .B2(n19046), .A(n19022), .ZN(P2_U2923) );
  AOI22_X1 U21992 ( .A1(n19056), .A2(P2_UWORD_REG_11__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_27__SCAN_IN), .ZN(n19024) );
  OAI21_X1 U21993 ( .B1(n19025), .B2(n19046), .A(n19024), .ZN(P2_U2924) );
  AOI22_X1 U21994 ( .A1(n19056), .A2(P2_UWORD_REG_10__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_26__SCAN_IN), .ZN(n19026) );
  OAI21_X1 U21995 ( .B1(n19027), .B2(n19046), .A(n19026), .ZN(P2_U2925) );
  AOI22_X1 U21996 ( .A1(n19056), .A2(P2_UWORD_REG_9__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_25__SCAN_IN), .ZN(n19028) );
  OAI21_X1 U21997 ( .B1(n19029), .B2(n19046), .A(n19028), .ZN(P2_U2926) );
  AOI22_X1 U21998 ( .A1(n19056), .A2(P2_UWORD_REG_8__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_24__SCAN_IN), .ZN(n19030) );
  OAI21_X1 U21999 ( .B1(n19031), .B2(n19046), .A(n19030), .ZN(P2_U2927) );
  AOI22_X1 U22000 ( .A1(n19056), .A2(P2_UWORD_REG_7__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_23__SCAN_IN), .ZN(n19032) );
  OAI21_X1 U22001 ( .B1(n21103), .B2(n19046), .A(n19032), .ZN(P2_U2928) );
  INV_X1 U22002 ( .A(P2_EAX_REG_22__SCAN_IN), .ZN(n19034) );
  AOI22_X1 U22003 ( .A1(n19056), .A2(P2_UWORD_REG_6__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_22__SCAN_IN), .ZN(n19033) );
  OAI21_X1 U22004 ( .B1(n19034), .B2(n19046), .A(n19033), .ZN(P2_U2929) );
  AOI22_X1 U22005 ( .A1(n19850), .A2(P2_UWORD_REG_5__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_21__SCAN_IN), .ZN(n19035) );
  OAI21_X1 U22006 ( .B1(n19036), .B2(n19046), .A(n19035), .ZN(P2_U2930) );
  INV_X1 U22007 ( .A(P2_EAX_REG_20__SCAN_IN), .ZN(n19038) );
  AOI22_X1 U22008 ( .A1(n19056), .A2(P2_UWORD_REG_4__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_20__SCAN_IN), .ZN(n19037) );
  OAI21_X1 U22009 ( .B1(n19038), .B2(n19046), .A(n19037), .ZN(P2_U2931) );
  AOI22_X1 U22010 ( .A1(n19850), .A2(P2_UWORD_REG_3__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_19__SCAN_IN), .ZN(n19039) );
  OAI21_X1 U22011 ( .B1(n19040), .B2(n19046), .A(n19039), .ZN(P2_U2932) );
  INV_X1 U22012 ( .A(P2_EAX_REG_18__SCAN_IN), .ZN(n19042) );
  INV_X2 U22013 ( .A(n19059), .ZN(n19076) );
  AOI22_X1 U22014 ( .A1(n19850), .A2(P2_UWORD_REG_2__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_18__SCAN_IN), .ZN(n19041) );
  OAI21_X1 U22015 ( .B1(n19042), .B2(n19046), .A(n19041), .ZN(P2_U2933) );
  AOI22_X1 U22016 ( .A1(n19850), .A2(P2_UWORD_REG_1__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_17__SCAN_IN), .ZN(n19043) );
  OAI21_X1 U22017 ( .B1(n19044), .B2(n19046), .A(n19043), .ZN(P2_U2934) );
  AOI22_X1 U22018 ( .A1(n19850), .A2(P2_UWORD_REG_0__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_16__SCAN_IN), .ZN(n19045) );
  OAI21_X1 U22019 ( .B1(n19047), .B2(n19046), .A(n19045), .ZN(P2_U2935) );
  AOI22_X1 U22020 ( .A1(n19850), .A2(P2_LWORD_REG_15__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_15__SCAN_IN), .ZN(n19048) );
  OAI21_X1 U22021 ( .B1(n13355), .B2(n19078), .A(n19048), .ZN(P2_U2936) );
  INV_X1 U22022 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n20998) );
  AOI22_X1 U22023 ( .A1(P2_EAX_REG_14__SCAN_IN), .A2(n19057), .B1(n19056), 
        .B2(P2_LWORD_REG_14__SCAN_IN), .ZN(n19049) );
  OAI21_X1 U22024 ( .B1(n19059), .B2(n20998), .A(n19049), .ZN(P2_U2937) );
  AOI22_X1 U22025 ( .A1(n19850), .A2(P2_LWORD_REG_13__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_13__SCAN_IN), .ZN(n19050) );
  OAI21_X1 U22026 ( .B1(n19051), .B2(n19078), .A(n19050), .ZN(P2_U2938) );
  AOI22_X1 U22027 ( .A1(n19850), .A2(P2_LWORD_REG_12__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_12__SCAN_IN), .ZN(n19052) );
  OAI21_X1 U22028 ( .B1(n19053), .B2(n19078), .A(n19052), .ZN(P2_U2939) );
  AOI22_X1 U22029 ( .A1(n19850), .A2(P2_LWORD_REG_11__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_11__SCAN_IN), .ZN(n19054) );
  OAI21_X1 U22030 ( .B1(n19055), .B2(n19078), .A(n19054), .ZN(P2_U2940) );
  AOI22_X1 U22031 ( .A1(P2_EAX_REG_10__SCAN_IN), .A2(n19057), .B1(n19056), 
        .B2(P2_LWORD_REG_10__SCAN_IN), .ZN(n19058) );
  OAI21_X1 U22032 ( .B1(n19059), .B2(n20945), .A(n19058), .ZN(P2_U2941) );
  AOI22_X1 U22033 ( .A1(n19850), .A2(P2_LWORD_REG_9__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_9__SCAN_IN), .ZN(n19060) );
  OAI21_X1 U22034 ( .B1(n19061), .B2(n19078), .A(n19060), .ZN(P2_U2942) );
  AOI22_X1 U22035 ( .A1(n19850), .A2(P2_LWORD_REG_8__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_8__SCAN_IN), .ZN(n19062) );
  OAI21_X1 U22036 ( .B1(n19063), .B2(n19078), .A(n19062), .ZN(P2_U2943) );
  AOI22_X1 U22037 ( .A1(n19850), .A2(P2_LWORD_REG_7__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_7__SCAN_IN), .ZN(n19064) );
  OAI21_X1 U22038 ( .B1(n19065), .B2(n19078), .A(n19064), .ZN(P2_U2944) );
  AOI22_X1 U22039 ( .A1(n19850), .A2(P2_LWORD_REG_6__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_6__SCAN_IN), .ZN(n19066) );
  OAI21_X1 U22040 ( .B1(n19067), .B2(n19078), .A(n19066), .ZN(P2_U2945) );
  INV_X1 U22041 ( .A(P2_EAX_REG_5__SCAN_IN), .ZN(n21093) );
  AOI22_X1 U22042 ( .A1(n19850), .A2(P2_LWORD_REG_5__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_5__SCAN_IN), .ZN(n19068) );
  OAI21_X1 U22043 ( .B1(n21093), .B2(n19078), .A(n19068), .ZN(P2_U2946) );
  INV_X1 U22044 ( .A(P2_EAX_REG_4__SCAN_IN), .ZN(n19070) );
  AOI22_X1 U22045 ( .A1(n19850), .A2(P2_LWORD_REG_4__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_4__SCAN_IN), .ZN(n19069) );
  OAI21_X1 U22046 ( .B1(n19070), .B2(n19078), .A(n19069), .ZN(P2_U2947) );
  INV_X1 U22047 ( .A(P2_EAX_REG_3__SCAN_IN), .ZN(n19072) );
  AOI22_X1 U22048 ( .A1(n19850), .A2(P2_LWORD_REG_3__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_3__SCAN_IN), .ZN(n19071) );
  OAI21_X1 U22049 ( .B1(n19072), .B2(n19078), .A(n19071), .ZN(P2_U2948) );
  AOI22_X1 U22050 ( .A1(n19850), .A2(P2_LWORD_REG_2__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_2__SCAN_IN), .ZN(n19073) );
  OAI21_X1 U22051 ( .B1(n20879), .B2(n19078), .A(n19073), .ZN(P2_U2949) );
  INV_X1 U22052 ( .A(P2_EAX_REG_1__SCAN_IN), .ZN(n19075) );
  AOI22_X1 U22053 ( .A1(n19850), .A2(P2_LWORD_REG_1__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_1__SCAN_IN), .ZN(n19074) );
  OAI21_X1 U22054 ( .B1(n19075), .B2(n19078), .A(n19074), .ZN(P2_U2950) );
  AOI22_X1 U22055 ( .A1(n19850), .A2(P2_LWORD_REG_0__SCAN_IN), .B1(n19076), 
        .B2(P2_DATAO_REG_0__SCAN_IN), .ZN(n19077) );
  OAI21_X1 U22056 ( .B1(n13358), .B2(n19078), .A(n19077), .ZN(P2_U2951) );
  AOI22_X1 U22057 ( .A1(n19082), .A2(P2_LWORD_REG_10__SCAN_IN), .B1(
        P2_EAX_REG_10__SCAN_IN), .B2(n19081), .ZN(n19080) );
  NAND2_X1 U22058 ( .A1(n19080), .A2(n19079), .ZN(P2_U2977) );
  AOI22_X1 U22059 ( .A1(n19082), .A2(P2_LWORD_REG_14__SCAN_IN), .B1(n19081), 
        .B2(P2_EAX_REG_14__SCAN_IN), .ZN(n19084) );
  NAND2_X1 U22060 ( .A1(n19084), .A2(n19083), .ZN(P2_U2981) );
  AOI22_X1 U22061 ( .A1(n19086), .A2(P2_PHYADDRPOINTER_REG_4__SCAN_IN), .B1(
        P2_REIP_REG_4__SCAN_IN), .B2(n19085), .ZN(n19096) );
  NAND2_X1 U22062 ( .A1(n19088), .A2(n19087), .ZN(n19091) );
  NAND2_X1 U22063 ( .A1(n19089), .A2(n19104), .ZN(n19090) );
  OAI211_X1 U22064 ( .C1(n19093), .C2(n19092), .A(n19091), .B(n19090), .ZN(
        n19094) );
  INV_X1 U22065 ( .A(n19094), .ZN(n19095) );
  OAI211_X1 U22066 ( .C1(n19098), .C2(n19097), .A(n19096), .B(n19095), .ZN(
        P2_U3010) );
  INV_X1 U22067 ( .A(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n20950) );
  INV_X1 U22068 ( .A(n19099), .ZN(n19103) );
  AOI22_X1 U22069 ( .A1(n19103), .A2(n19102), .B1(n19101), .B2(n19100), .ZN(
        n19107) );
  NAND2_X1 U22070 ( .A1(n19105), .A2(n19104), .ZN(n19106) );
  OAI211_X1 U22071 ( .C1(n19109), .C2(n19108), .A(n19107), .B(n19106), .ZN(
        n19110) );
  INV_X1 U22072 ( .A(n19110), .ZN(n19112) );
  OAI211_X1 U22073 ( .C1(n19113), .C2(n20950), .A(n19112), .B(n19111), .ZN(
        P2_U3012) );
  AOI22_X1 U22074 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n19151), .B1(
        BUF2_REG_24__SCAN_IN), .B2(n19152), .ZN(n19559) );
  INV_X1 U22075 ( .A(n19559), .ZN(n19657) );
  AND2_X1 U22076 ( .A1(n19114), .A2(n19148), .ZN(n19656) );
  AOI22_X1 U22077 ( .A1(n19657), .A2(n19702), .B1(n19149), .B2(n19656), .ZN(
        n19118) );
  AOI22_X1 U22078 ( .A1(BUF1_REG_16__SCAN_IN), .A2(n19151), .B1(
        BUF2_REG_16__SCAN_IN), .B2(n19152), .ZN(n19484) );
  AOI22_X1 U22079 ( .A1(n19116), .A2(n19153), .B1(n19182), .B2(n19658), .ZN(
        n19117) );
  OAI211_X1 U22080 ( .C1(n19157), .C2(n20891), .A(n19118), .B(n19117), .ZN(
        P2_U3048) );
  INV_X1 U22081 ( .A(P2_INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n19123) );
  AOI22_X1 U22082 ( .A1(BUF2_REG_25__SCAN_IN), .A2(n19152), .B1(
        BUF1_REG_25__SCAN_IN), .B2(n19151), .ZN(n19565) );
  AOI22_X1 U22083 ( .A1(n19663), .A2(n19702), .B1(n19149), .B2(n19661), .ZN(
        n19122) );
  AOI22_X1 U22084 ( .A1(BUF1_REG_17__SCAN_IN), .A2(n19151), .B1(
        BUF2_REG_17__SCAN_IN), .B2(n19152), .ZN(n19450) );
  INV_X1 U22085 ( .A(n19450), .ZN(n19662) );
  AOI22_X1 U22086 ( .A1(n19120), .A2(n19153), .B1(n19182), .B2(n19662), .ZN(
        n19121) );
  OAI211_X1 U22087 ( .C1(n19157), .C2(n19123), .A(n19122), .B(n19121), .ZN(
        P2_U3049) );
  AOI22_X1 U22088 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n19151), .B1(
        BUF2_REG_26__SCAN_IN), .B2(n19152), .ZN(n19571) );
  AOI22_X1 U22089 ( .A1(n19668), .A2(n19702), .B1(n19149), .B2(n19666), .ZN(
        n19128) );
  AOI22_X1 U22090 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n19151), .B1(
        BUF2_REG_18__SCAN_IN), .B2(n19152), .ZN(n19491) );
  INV_X1 U22091 ( .A(n19491), .ZN(n19667) );
  AOI22_X1 U22092 ( .A1(n19126), .A2(n19153), .B1(n19182), .B2(n19667), .ZN(
        n19127) );
  OAI211_X1 U22093 ( .C1(n19157), .C2(n12872), .A(n19128), .B(n19127), .ZN(
        P2_U3050) );
  AOI22_X1 U22094 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n19151), .B1(
        BUF2_REG_27__SCAN_IN), .B2(n19152), .ZN(n19577) );
  INV_X1 U22095 ( .A(n19577), .ZN(n19673) );
  AOI22_X1 U22096 ( .A1(n19673), .A2(n19702), .B1(n19149), .B2(n19671), .ZN(
        n19132) );
  NOR2_X2 U22097 ( .A1(n19130), .A2(n19613), .ZN(n19672) );
  AOI22_X1 U22098 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n19151), .B1(
        BUF2_REG_19__SCAN_IN), .B2(n19152), .ZN(n19363) );
  AOI22_X1 U22099 ( .A1(n19672), .A2(n19153), .B1(n19182), .B2(n19674), .ZN(
        n19131) );
  OAI211_X1 U22100 ( .C1(n19157), .C2(n19133), .A(n19132), .B(n19131), .ZN(
        P2_U3051) );
  OAI22_X2 U22101 ( .A1(n20974), .A2(n19144), .B1(n14307), .B2(n19146), .ZN(
        n19686) );
  NOR2_X2 U22102 ( .A1(n19134), .A2(n19139), .ZN(n19683) );
  AOI22_X1 U22103 ( .A1(n19686), .A2(n19702), .B1(n19149), .B2(n19683), .ZN(
        n19137) );
  NOR2_X2 U22104 ( .A1(n19135), .A2(n19613), .ZN(n19684) );
  OAI22_X1 U22105 ( .A1(n15074), .A2(n19146), .B1(n15075), .B2(n19144), .ZN(
        n19685) );
  AOI22_X1 U22106 ( .A1(n19684), .A2(n19153), .B1(n19182), .B2(n19685), .ZN(
        n19136) );
  OAI211_X1 U22107 ( .C1(n19157), .C2(n19138), .A(n19137), .B(n19136), .ZN(
        P2_U3053) );
  INV_X1 U22108 ( .A(P2_INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n19143) );
  AOI22_X2 U22109 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n19151), .B1(
        BUF2_REG_30__SCAN_IN), .B2(n19152), .ZN(n19596) );
  INV_X1 U22110 ( .A(n19596), .ZN(n19691) );
  AOI22_X1 U22111 ( .A1(n19691), .A2(n19702), .B1(n19149), .B2(n9807), .ZN(
        n19142) );
  NOR2_X2 U22112 ( .A1(n19140), .A2(n19613), .ZN(n19690) );
  OAI22_X2 U22113 ( .A1(n14540), .A2(n19146), .B1(n20905), .B2(n19144), .ZN(
        n19692) );
  AOI22_X1 U22114 ( .A1(n19690), .A2(n19153), .B1(n19182), .B2(n19692), .ZN(
        n19141) );
  OAI211_X1 U22115 ( .C1(n19157), .C2(n19143), .A(n19142), .B(n19141), .ZN(
        P2_U3054) );
  OAI22_X1 U22116 ( .A1(n19147), .A2(n19146), .B1(n19145), .B2(n19144), .ZN(
        n19699) );
  AND2_X1 U22117 ( .A1(n10443), .A2(n19148), .ZN(n19696) );
  AOI22_X1 U22118 ( .A1(n19699), .A2(n19702), .B1(n19149), .B2(n19696), .ZN(
        n19155) );
  NOR2_X2 U22119 ( .A1(n19150), .A2(n19613), .ZN(n19697) );
  AOI22_X1 U22120 ( .A1(BUF2_REG_23__SCAN_IN), .A2(n19152), .B1(
        BUF1_REG_23__SCAN_IN), .B2(n19151), .ZN(n19436) );
  AOI22_X1 U22121 ( .A1(n19697), .A2(n19153), .B1(n19182), .B2(n19701), .ZN(
        n19154) );
  OAI211_X1 U22122 ( .C1(n19157), .C2(n19156), .A(n19155), .B(n19154), .ZN(
        P2_U3055) );
  NOR2_X1 U22123 ( .A1(n19406), .A2(n19219), .ZN(n19180) );
  NOR3_X1 U22124 ( .A1(n19159), .A2(n19180), .A3(n19842), .ZN(n19161) );
  AOI211_X2 U22125 ( .C1(n19162), .C2(n19842), .A(n19708), .B(n19161), .ZN(
        n19181) );
  AOI22_X1 U22126 ( .A1(n19181), .A2(n19116), .B1(n19656), .B2(n19180), .ZN(
        n19166) );
  NAND2_X1 U22127 ( .A1(n19788), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19791) );
  INV_X1 U22128 ( .A(n19791), .ZN(n19350) );
  NAND2_X1 U22129 ( .A1(n19350), .A2(n19160), .ZN(n19163) );
  AOI21_X1 U22130 ( .B1(n19163), .B2(n19162), .A(n19161), .ZN(n19164) );
  OAI211_X1 U22131 ( .C1(n19180), .C2(n19798), .A(n19164), .B(n19648), .ZN(
        n19183) );
  AOI22_X1 U22132 ( .A1(P2_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n19183), .B1(
        n19182), .B2(n19657), .ZN(n19165) );
  OAI211_X1 U22133 ( .C1(n19484), .C2(n19217), .A(n19166), .B(n19165), .ZN(
        P2_U3056) );
  AOI22_X1 U22134 ( .A1(n19181), .A2(n19120), .B1(n19661), .B2(n19180), .ZN(
        n19168) );
  AOI22_X1 U22135 ( .A1(P2_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n19183), .B1(
        n19182), .B2(n19663), .ZN(n19167) );
  OAI211_X1 U22136 ( .C1(n19450), .C2(n19217), .A(n19168), .B(n19167), .ZN(
        P2_U3057) );
  AOI22_X1 U22137 ( .A1(n19181), .A2(n19126), .B1(n19666), .B2(n19180), .ZN(
        n19170) );
  AOI22_X1 U22138 ( .A1(P2_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n19183), .B1(
        n19182), .B2(n19668), .ZN(n19169) );
  OAI211_X1 U22139 ( .C1(n19491), .C2(n19217), .A(n19170), .B(n19169), .ZN(
        P2_U3058) );
  AOI22_X1 U22140 ( .A1(n19181), .A2(n19672), .B1(n19671), .B2(n19180), .ZN(
        n19172) );
  AOI22_X1 U22141 ( .A1(P2_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n19183), .B1(
        n19182), .B2(n19673), .ZN(n19171) );
  OAI211_X1 U22142 ( .C1(n19363), .C2(n19217), .A(n19172), .B(n19171), .ZN(
        P2_U3059) );
  AOI22_X1 U22143 ( .A1(n19181), .A2(n19678), .B1(n19677), .B2(n19180), .ZN(
        n19174) );
  AOI22_X1 U22144 ( .A1(P2_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n19183), .B1(
        n19182), .B2(n19680), .ZN(n19173) );
  OAI211_X1 U22145 ( .C1(n19583), .C2(n19217), .A(n19174), .B(n19173), .ZN(
        P2_U3060) );
  AOI22_X1 U22146 ( .A1(n19181), .A2(n19684), .B1(n19683), .B2(n19180), .ZN(
        n19176) );
  AOI22_X1 U22147 ( .A1(P2_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n19183), .B1(
        n19182), .B2(n19686), .ZN(n19175) );
  OAI211_X1 U22148 ( .C1(n19590), .C2(n19217), .A(n19176), .B(n19175), .ZN(
        P2_U3061) );
  AOI22_X1 U22149 ( .A1(n19181), .A2(n19690), .B1(n9807), .B2(n19180), .ZN(
        n19178) );
  AOI22_X1 U22150 ( .A1(P2_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n19183), .B1(
        n19207), .B2(n19692), .ZN(n19177) );
  OAI211_X1 U22151 ( .C1(n19596), .C2(n19179), .A(n19178), .B(n19177), .ZN(
        P2_U3062) );
  AOI22_X1 U22152 ( .A1(n19181), .A2(n19697), .B1(n19696), .B2(n19180), .ZN(
        n19185) );
  AOI22_X1 U22153 ( .A1(P2_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n19183), .B1(
        n19182), .B2(n19699), .ZN(n19184) );
  OAI211_X1 U22154 ( .C1(n19436), .C2(n19217), .A(n19185), .B(n19184), .ZN(
        P2_U3063) );
  NOR2_X1 U22155 ( .A1(n19437), .A2(n19219), .ZN(n19212) );
  OAI21_X1 U22156 ( .B1(n19186), .B2(n19212), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19189) );
  INV_X1 U22157 ( .A(n19440), .ZN(n19188) );
  INV_X1 U22158 ( .A(n19219), .ZN(n19187) );
  NAND2_X1 U22159 ( .A1(n19188), .A2(n19187), .ZN(n19192) );
  NAND2_X1 U22160 ( .A1(n19189), .A2(n19192), .ZN(n19213) );
  AOI22_X1 U22161 ( .A1(n19213), .A2(n19116), .B1(n19656), .B2(n19212), .ZN(
        n19198) );
  INV_X1 U22162 ( .A(n19212), .ZN(n19191) );
  OAI21_X1 U22163 ( .B1(n19190), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19191), 
        .ZN(n19195) );
  INV_X1 U22164 ( .A(n19468), .ZN(n19784) );
  NOR2_X1 U22165 ( .A1(n19238), .A2(n19207), .ZN(n19193) );
  OAI21_X1 U22166 ( .B1(n19193), .B2(n19836), .A(n19192), .ZN(n19194) );
  MUX2_X1 U22167 ( .A(n19195), .B(n19194), .S(n19612), .Z(n19196) );
  NAND2_X1 U22168 ( .A1(n19196), .A2(n19648), .ZN(n19214) );
  AOI22_X1 U22169 ( .A1(P2_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n19214), .B1(
        n19238), .B2(n19658), .ZN(n19197) );
  OAI211_X1 U22170 ( .C1(n19559), .C2(n19217), .A(n19198), .B(n19197), .ZN(
        P2_U3064) );
  AOI22_X1 U22171 ( .A1(n19213), .A2(n19120), .B1(n19661), .B2(n19212), .ZN(
        n19200) );
  AOI22_X1 U22172 ( .A1(P2_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n19214), .B1(
        n19207), .B2(n19663), .ZN(n19199) );
  OAI211_X1 U22173 ( .C1(n19450), .C2(n19248), .A(n19200), .B(n19199), .ZN(
        P2_U3065) );
  AOI22_X1 U22174 ( .A1(n19213), .A2(n19126), .B1(n19666), .B2(n19212), .ZN(
        n19202) );
  AOI22_X1 U22175 ( .A1(P2_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n19214), .B1(
        n19207), .B2(n19668), .ZN(n19201) );
  OAI211_X1 U22176 ( .C1(n19491), .C2(n19248), .A(n19202), .B(n19201), .ZN(
        P2_U3066) );
  AOI22_X1 U22177 ( .A1(n19213), .A2(n19672), .B1(n19671), .B2(n19212), .ZN(
        n19204) );
  AOI22_X1 U22178 ( .A1(P2_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n19214), .B1(
        n19238), .B2(n19674), .ZN(n19203) );
  OAI211_X1 U22179 ( .C1(n19577), .C2(n19217), .A(n19204), .B(n19203), .ZN(
        P2_U3067) );
  AOI22_X1 U22180 ( .A1(n19213), .A2(n19678), .B1(n19677), .B2(n19212), .ZN(
        n19206) );
  AOI22_X1 U22181 ( .A1(P2_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n19214), .B1(
        n19207), .B2(n19680), .ZN(n19205) );
  OAI211_X1 U22182 ( .C1(n19583), .C2(n19248), .A(n19206), .B(n19205), .ZN(
        P2_U3068) );
  AOI22_X1 U22183 ( .A1(n19213), .A2(n19684), .B1(n19683), .B2(n19212), .ZN(
        n19209) );
  AOI22_X1 U22184 ( .A1(P2_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n19214), .B1(
        n19207), .B2(n19686), .ZN(n19208) );
  OAI211_X1 U22185 ( .C1(n19590), .C2(n19248), .A(n19209), .B(n19208), .ZN(
        P2_U3069) );
  AOI22_X1 U22186 ( .A1(n19213), .A2(n19690), .B1(n9807), .B2(n19212), .ZN(
        n19211) );
  AOI22_X1 U22187 ( .A1(P2_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n19214), .B1(
        n19238), .B2(n19692), .ZN(n19210) );
  OAI211_X1 U22188 ( .C1(n19596), .C2(n19217), .A(n19211), .B(n19210), .ZN(
        P2_U3070) );
  AOI22_X1 U22189 ( .A1(n19213), .A2(n19697), .B1(n19696), .B2(n19212), .ZN(
        n19216) );
  AOI22_X1 U22190 ( .A1(P2_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n19214), .B1(
        n19238), .B2(n19701), .ZN(n19215) );
  OAI211_X1 U22191 ( .C1(n19606), .C2(n19217), .A(n19216), .B(n19215), .ZN(
        P2_U3071) );
  INV_X1 U22192 ( .A(n19470), .ZN(n19218) );
  NOR2_X1 U22193 ( .A1(n19218), .A2(n19219), .ZN(n19243) );
  AOI22_X1 U22194 ( .A1(n19658), .A2(n19268), .B1(n19243), .B2(n19656), .ZN(
        n19229) );
  OAI21_X1 U22195 ( .B1(n19791), .B2(n19468), .A(n19612), .ZN(n19227) );
  NOR2_X1 U22196 ( .A1(n19814), .A2(n19219), .ZN(n19223) );
  INV_X1 U22197 ( .A(n19224), .ZN(n19221) );
  INV_X1 U22198 ( .A(n19243), .ZN(n19220) );
  OAI211_X1 U22199 ( .C1(n19221), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19220), 
        .B(n19790), .ZN(n19222) );
  OAI211_X1 U22200 ( .C1(n19227), .C2(n19223), .A(n19648), .B(n19222), .ZN(
        n19245) );
  INV_X1 U22201 ( .A(n19223), .ZN(n19226) );
  OAI21_X1 U22202 ( .B1(n19224), .B2(n19243), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19225) );
  OAI21_X1 U22203 ( .B1(n19227), .B2(n19226), .A(n19225), .ZN(n19244) );
  AOI22_X1 U22204 ( .A1(P2_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n19245), .B1(
        n19116), .B2(n19244), .ZN(n19228) );
  OAI211_X1 U22205 ( .C1(n19559), .C2(n19248), .A(n19229), .B(n19228), .ZN(
        P2_U3072) );
  AOI22_X1 U22206 ( .A1(n19662), .A2(n19268), .B1(n19243), .B2(n19661), .ZN(
        n19231) );
  AOI22_X1 U22207 ( .A1(P2_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n19245), .B1(
        n19120), .B2(n19244), .ZN(n19230) );
  OAI211_X1 U22208 ( .C1(n19565), .C2(n19248), .A(n19231), .B(n19230), .ZN(
        P2_U3073) );
  AOI22_X1 U22209 ( .A1(n19668), .A2(n19238), .B1(n19243), .B2(n19666), .ZN(
        n19233) );
  AOI22_X1 U22210 ( .A1(P2_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n19245), .B1(
        n19126), .B2(n19244), .ZN(n19232) );
  OAI211_X1 U22211 ( .C1(n19491), .C2(n19278), .A(n19233), .B(n19232), .ZN(
        P2_U3074) );
  AOI22_X1 U22212 ( .A1(n19673), .A2(n19238), .B1(n19243), .B2(n19671), .ZN(
        n19235) );
  AOI22_X1 U22213 ( .A1(P2_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n19245), .B1(
        n19672), .B2(n19244), .ZN(n19234) );
  OAI211_X1 U22214 ( .C1(n19363), .C2(n19278), .A(n19235), .B(n19234), .ZN(
        P2_U3075) );
  AOI22_X1 U22215 ( .A1(n19680), .A2(n19238), .B1(n19677), .B2(n19243), .ZN(
        n19237) );
  AOI22_X1 U22216 ( .A1(P2_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n19245), .B1(
        n19678), .B2(n19244), .ZN(n19236) );
  OAI211_X1 U22217 ( .C1(n19583), .C2(n19278), .A(n19237), .B(n19236), .ZN(
        P2_U3076) );
  AOI22_X1 U22218 ( .A1(n19686), .A2(n19238), .B1(n19243), .B2(n19683), .ZN(
        n19240) );
  AOI22_X1 U22219 ( .A1(P2_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n19245), .B1(
        n19684), .B2(n19244), .ZN(n19239) );
  OAI211_X1 U22220 ( .C1(n19590), .C2(n19278), .A(n19240), .B(n19239), .ZN(
        P2_U3077) );
  AOI22_X1 U22221 ( .A1(n19692), .A2(n19268), .B1(n19243), .B2(n9807), .ZN(
        n19242) );
  AOI22_X1 U22222 ( .A1(P2_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n19245), .B1(
        n19690), .B2(n19244), .ZN(n19241) );
  OAI211_X1 U22223 ( .C1(n19596), .C2(n19248), .A(n19242), .B(n19241), .ZN(
        P2_U3078) );
  AOI22_X1 U22224 ( .A1(n19701), .A2(n19268), .B1(n19243), .B2(n19696), .ZN(
        n19247) );
  AOI22_X1 U22225 ( .A1(P2_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n19245), .B1(
        n19697), .B2(n19244), .ZN(n19246) );
  OAI211_X1 U22226 ( .C1(n19606), .C2(n19248), .A(n19247), .B(n19246), .ZN(
        P2_U3079) );
  OR2_X1 U22227 ( .A1(n19249), .A2(n19320), .ZN(n19515) );
  INV_X1 U22228 ( .A(n19515), .ZN(n19518) );
  NAND2_X1 U22229 ( .A1(n19518), .A2(n19796), .ZN(n19255) );
  INV_X1 U22230 ( .A(n19319), .ZN(n19317) );
  NOR3_X2 U22231 ( .A1(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n19317), .ZN(n19273) );
  OAI21_X1 U22232 ( .B1(n19250), .B2(n19273), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19251) );
  OAI21_X1 U22233 ( .B1(n19255), .B2(n19790), .A(n19251), .ZN(n19274) );
  AOI22_X1 U22234 ( .A1(n19274), .A2(n19116), .B1(n19656), .B2(n19273), .ZN(
        n19259) );
  AOI21_X1 U22235 ( .B1(n19252), .B2(P2_STATE2_REG_2__SCAN_IN), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19257) );
  OAI21_X1 U22236 ( .B1(n19268), .B2(n19303), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19254) );
  AOI21_X1 U22237 ( .B1(n19255), .B2(n19254), .A(n19613), .ZN(n19256) );
  AOI22_X1 U22238 ( .A1(P2_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n19275), .B1(
        n19303), .B2(n19658), .ZN(n19258) );
  OAI211_X1 U22239 ( .C1(n19559), .C2(n19278), .A(n19259), .B(n19258), .ZN(
        P2_U3080) );
  AOI22_X1 U22240 ( .A1(n19274), .A2(n19120), .B1(n19661), .B2(n19273), .ZN(
        n19261) );
  AOI22_X1 U22241 ( .A1(P2_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n19275), .B1(
        n19268), .B2(n19663), .ZN(n19260) );
  OAI211_X1 U22242 ( .C1(n19450), .C2(n19315), .A(n19261), .B(n19260), .ZN(
        P2_U3081) );
  AOI22_X1 U22243 ( .A1(n19274), .A2(n19126), .B1(n19666), .B2(n19273), .ZN(
        n19263) );
  AOI22_X1 U22244 ( .A1(P2_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n19275), .B1(
        n19268), .B2(n19668), .ZN(n19262) );
  OAI211_X1 U22245 ( .C1(n19491), .C2(n19315), .A(n19263), .B(n19262), .ZN(
        P2_U3082) );
  AOI22_X1 U22246 ( .A1(n19274), .A2(n19672), .B1(n19671), .B2(n19273), .ZN(
        n19265) );
  AOI22_X1 U22247 ( .A1(P2_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n19275), .B1(
        n19268), .B2(n19673), .ZN(n19264) );
  OAI211_X1 U22248 ( .C1(n19363), .C2(n19315), .A(n19265), .B(n19264), .ZN(
        P2_U3083) );
  AOI22_X1 U22249 ( .A1(n19274), .A2(n19678), .B1(n19677), .B2(n19273), .ZN(
        n19267) );
  AOI22_X1 U22250 ( .A1(P2_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n19275), .B1(
        n19268), .B2(n19680), .ZN(n19266) );
  OAI211_X1 U22251 ( .C1(n19583), .C2(n19315), .A(n19267), .B(n19266), .ZN(
        P2_U3084) );
  AOI22_X1 U22252 ( .A1(n19274), .A2(n19684), .B1(n19683), .B2(n19273), .ZN(
        n19270) );
  AOI22_X1 U22253 ( .A1(P2_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n19275), .B1(
        n19268), .B2(n19686), .ZN(n19269) );
  OAI211_X1 U22254 ( .C1(n19590), .C2(n19315), .A(n19270), .B(n19269), .ZN(
        P2_U3085) );
  AOI22_X1 U22255 ( .A1(n19274), .A2(n19690), .B1(n9807), .B2(n19273), .ZN(
        n19272) );
  AOI22_X1 U22256 ( .A1(P2_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n19275), .B1(
        n19303), .B2(n19692), .ZN(n19271) );
  OAI211_X1 U22257 ( .C1(n19596), .C2(n19278), .A(n19272), .B(n19271), .ZN(
        P2_U3086) );
  AOI22_X1 U22258 ( .A1(n19274), .A2(n19697), .B1(n19696), .B2(n19273), .ZN(
        n19277) );
  AOI22_X1 U22259 ( .A1(P2_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n19275), .B1(
        n19303), .B2(n19701), .ZN(n19276) );
  OAI211_X1 U22260 ( .C1(n19606), .C2(n19278), .A(n19277), .B(n19276), .ZN(
        P2_U3087) );
  OAI21_X1 U22261 ( .B1(n19791), .B2(n19555), .A(n19612), .ZN(n19287) );
  NAND2_X1 U22262 ( .A1(n19319), .A2(n19814), .ZN(n19286) );
  INV_X1 U22263 ( .A(n19286), .ZN(n19279) );
  OR2_X1 U22264 ( .A1(n19287), .A2(n19279), .ZN(n19283) );
  NAND2_X1 U22265 ( .A1(n19284), .A2(n19798), .ZN(n19281) );
  NOR2_X1 U22266 ( .A1(n19317), .A2(n19406), .ZN(n19310) );
  NOR2_X1 U22267 ( .A1(n19310), .A2(n19612), .ZN(n19280) );
  AOI21_X1 U22268 ( .B1(n19281), .B2(n19280), .A(n19613), .ZN(n19282) );
  INV_X1 U22269 ( .A(P2_INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n19290) );
  NOR2_X2 U22270 ( .A1(n19347), .A2(n19555), .ZN(n19336) );
  AOI22_X1 U22271 ( .A1(n19658), .A2(n19336), .B1(n19656), .B2(n19310), .ZN(
        n19289) );
  OAI21_X1 U22272 ( .B1(n19284), .B2(n19310), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19285) );
  OAI21_X1 U22273 ( .B1(n19287), .B2(n19286), .A(n19285), .ZN(n19311) );
  AOI22_X1 U22274 ( .A1(n19116), .A2(n19311), .B1(n19303), .B2(n19657), .ZN(
        n19288) );
  OAI211_X1 U22275 ( .C1(n19307), .C2(n19290), .A(n19289), .B(n19288), .ZN(
        P2_U3088) );
  INV_X1 U22276 ( .A(P2_INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n19293) );
  AOI22_X1 U22277 ( .A1(n19663), .A2(n19303), .B1(n19661), .B2(n19310), .ZN(
        n19292) );
  AOI22_X1 U22278 ( .A1(n19120), .A2(n19311), .B1(n19336), .B2(n19662), .ZN(
        n19291) );
  OAI211_X1 U22279 ( .C1(n19307), .C2(n19293), .A(n19292), .B(n19291), .ZN(
        P2_U3089) );
  AOI22_X1 U22280 ( .A1(n19667), .A2(n19336), .B1(n19666), .B2(n19310), .ZN(
        n19295) );
  AOI22_X1 U22281 ( .A1(n19126), .A2(n19311), .B1(n19303), .B2(n19668), .ZN(
        n19294) );
  OAI211_X1 U22282 ( .C1(n19307), .C2(n19296), .A(n19295), .B(n19294), .ZN(
        P2_U3090) );
  INV_X1 U22283 ( .A(P2_INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n19299) );
  AOI22_X1 U22284 ( .A1(n19673), .A2(n19303), .B1(n19310), .B2(n19671), .ZN(
        n19298) );
  AOI22_X1 U22285 ( .A1(n19672), .A2(n19311), .B1(n19336), .B2(n19674), .ZN(
        n19297) );
  OAI211_X1 U22286 ( .C1(n19307), .C2(n19299), .A(n19298), .B(n19297), .ZN(
        P2_U3091) );
  INV_X1 U22287 ( .A(P2_INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n19302) );
  AOI22_X1 U22288 ( .A1(n19680), .A2(n19303), .B1(n19677), .B2(n19310), .ZN(
        n19301) );
  INV_X1 U22289 ( .A(n19583), .ZN(n19679) );
  AOI22_X1 U22290 ( .A1(n19678), .A2(n19311), .B1(n19336), .B2(n19679), .ZN(
        n19300) );
  OAI211_X1 U22291 ( .C1(n19307), .C2(n19302), .A(n19301), .B(n19300), .ZN(
        P2_U3092) );
  INV_X1 U22292 ( .A(P2_INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n19306) );
  AOI22_X1 U22293 ( .A1(n19686), .A2(n19303), .B1(n19683), .B2(n19310), .ZN(
        n19305) );
  AOI22_X1 U22294 ( .A1(n19684), .A2(n19311), .B1(n19336), .B2(n19685), .ZN(
        n19304) );
  OAI211_X1 U22295 ( .C1(n19307), .C2(n19306), .A(n19305), .B(n19304), .ZN(
        P2_U3093) );
  AOI22_X1 U22296 ( .A1(n19692), .A2(n19336), .B1(n9807), .B2(n19310), .ZN(
        n19309) );
  INV_X1 U22297 ( .A(n19307), .ZN(n19312) );
  AOI22_X1 U22298 ( .A1(P2_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n19312), .B1(
        n19690), .B2(n19311), .ZN(n19308) );
  OAI211_X1 U22299 ( .C1(n19596), .C2(n19315), .A(n19309), .B(n19308), .ZN(
        P2_U3094) );
  AOI22_X1 U22300 ( .A1(n19701), .A2(n19336), .B1(n19696), .B2(n19310), .ZN(
        n19314) );
  AOI22_X1 U22301 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n19312), .B1(
        n19697), .B2(n19311), .ZN(n19313) );
  OAI211_X1 U22302 ( .C1(n19606), .C2(n19315), .A(n19314), .B(n19313), .ZN(
        P2_U3095) );
  INV_X1 U22303 ( .A(n19336), .ZN(n19346) );
  NOR2_X1 U22304 ( .A1(n19317), .A2(n19437), .ZN(n19341) );
  OAI21_X1 U22305 ( .B1(n19321), .B2(n19341), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19316) );
  OAI21_X1 U22306 ( .B1(n19440), .B2(n19317), .A(n19316), .ZN(n19342) );
  AOI22_X1 U22307 ( .A1(n19342), .A2(n19116), .B1(n19656), .B2(n19341), .ZN(
        n19327) );
  OAI21_X1 U22308 ( .B1(n19336), .B2(n19372), .A(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19324) );
  NAND2_X1 U22309 ( .A1(n19320), .A2(n19319), .ZN(n19323) );
  AOI211_X1 U22310 ( .C1(n19321), .C2(n19798), .A(n19341), .B(n19612), .ZN(
        n19322) );
  AOI211_X1 U22311 ( .C1(n19324), .C2(n19323), .A(n19322), .B(n19613), .ZN(
        n19325) );
  AOI22_X1 U22312 ( .A1(P2_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n19343), .B1(
        n19372), .B2(n19658), .ZN(n19326) );
  OAI211_X1 U22313 ( .C1(n19559), .C2(n19346), .A(n19327), .B(n19326), .ZN(
        P2_U3096) );
  AOI22_X1 U22314 ( .A1(n19342), .A2(n19120), .B1(n19661), .B2(n19341), .ZN(
        n19329) );
  AOI22_X1 U22315 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n19343), .B1(
        n19336), .B2(n19663), .ZN(n19328) );
  OAI211_X1 U22316 ( .C1(n19450), .C2(n19370), .A(n19329), .B(n19328), .ZN(
        P2_U3097) );
  AOI22_X1 U22317 ( .A1(n19342), .A2(n19126), .B1(n19666), .B2(n19341), .ZN(
        n19331) );
  AOI22_X1 U22318 ( .A1(P2_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n19343), .B1(
        n19336), .B2(n19668), .ZN(n19330) );
  OAI211_X1 U22319 ( .C1(n19491), .C2(n19370), .A(n19331), .B(n19330), .ZN(
        P2_U3098) );
  AOI22_X1 U22320 ( .A1(n19342), .A2(n19672), .B1(n19671), .B2(n19341), .ZN(
        n19333) );
  AOI22_X1 U22321 ( .A1(P2_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n19343), .B1(
        n19372), .B2(n19674), .ZN(n19332) );
  OAI211_X1 U22322 ( .C1(n19577), .C2(n19346), .A(n19333), .B(n19332), .ZN(
        P2_U3099) );
  AOI22_X1 U22323 ( .A1(n19342), .A2(n19678), .B1(n19677), .B2(n19341), .ZN(
        n19335) );
  AOI22_X1 U22324 ( .A1(P2_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n19343), .B1(
        n19336), .B2(n19680), .ZN(n19334) );
  OAI211_X1 U22325 ( .C1(n19583), .C2(n19370), .A(n19335), .B(n19334), .ZN(
        P2_U3100) );
  AOI22_X1 U22326 ( .A1(n19342), .A2(n19684), .B1(n19683), .B2(n19341), .ZN(
        n19338) );
  AOI22_X1 U22327 ( .A1(P2_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n19343), .B1(
        n19336), .B2(n19686), .ZN(n19337) );
  OAI211_X1 U22328 ( .C1(n19590), .C2(n19370), .A(n19338), .B(n19337), .ZN(
        P2_U3101) );
  AOI22_X1 U22329 ( .A1(n19342), .A2(n19690), .B1(n9807), .B2(n19341), .ZN(
        n19340) );
  AOI22_X1 U22330 ( .A1(P2_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n19343), .B1(
        n19372), .B2(n19692), .ZN(n19339) );
  OAI211_X1 U22331 ( .C1(n19596), .C2(n19346), .A(n19340), .B(n19339), .ZN(
        P2_U3102) );
  AOI22_X1 U22332 ( .A1(n19342), .A2(n19697), .B1(n19696), .B2(n19341), .ZN(
        n19345) );
  AOI22_X1 U22333 ( .A1(P2_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n19343), .B1(
        n19372), .B2(n19701), .ZN(n19344) );
  OAI211_X1 U22334 ( .C1(n19606), .C2(n19346), .A(n19345), .B(n19344), .ZN(
        P2_U3103) );
  NAND2_X1 U22335 ( .A1(n19610), .A2(n19796), .ZN(n19352) );
  NOR3_X1 U22336 ( .A1(n19348), .A2(n19382), .A3(n19842), .ZN(n19351) );
  AOI211_X2 U22337 ( .C1(n19352), .C2(n19842), .A(n19708), .B(n19351), .ZN(
        n19371) );
  AOI22_X1 U22338 ( .A1(n19371), .A2(n19116), .B1(n19382), .B2(n19656), .ZN(
        n19356) );
  INV_X1 U22339 ( .A(n19789), .ZN(n19349) );
  NAND2_X1 U22340 ( .A1(n19350), .A2(n19349), .ZN(n19353) );
  AOI211_X1 U22341 ( .C1(n19353), .C2(n19352), .A(n19351), .B(n19613), .ZN(
        n19354) );
  OAI21_X1 U22342 ( .B1(n19382), .B2(n19798), .A(n19354), .ZN(n19373) );
  AOI22_X1 U22343 ( .A1(P2_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n19373), .B1(
        n19372), .B2(n19657), .ZN(n19355) );
  OAI211_X1 U22344 ( .C1(n19484), .C2(n19405), .A(n19356), .B(n19355), .ZN(
        P2_U3104) );
  AOI22_X1 U22345 ( .A1(n19371), .A2(n19120), .B1(n19382), .B2(n19661), .ZN(
        n19358) );
  AOI22_X1 U22346 ( .A1(P2_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n19373), .B1(
        n19372), .B2(n19663), .ZN(n19357) );
  OAI211_X1 U22347 ( .C1(n19450), .C2(n19405), .A(n19358), .B(n19357), .ZN(
        P2_U3105) );
  AOI22_X1 U22348 ( .A1(n19371), .A2(n19126), .B1(n19382), .B2(n19666), .ZN(
        n19360) );
  AOI22_X1 U22349 ( .A1(P2_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n19373), .B1(
        n19395), .B2(n19667), .ZN(n19359) );
  OAI211_X1 U22350 ( .C1(n19571), .C2(n19370), .A(n19360), .B(n19359), .ZN(
        P2_U3106) );
  AOI22_X1 U22351 ( .A1(n19371), .A2(n19672), .B1(n19382), .B2(n19671), .ZN(
        n19362) );
  AOI22_X1 U22352 ( .A1(P2_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n19373), .B1(
        n19372), .B2(n19673), .ZN(n19361) );
  OAI211_X1 U22353 ( .C1(n19363), .C2(n19405), .A(n19362), .B(n19361), .ZN(
        P2_U3107) );
  AOI22_X1 U22354 ( .A1(n19371), .A2(n19678), .B1(n19382), .B2(n19677), .ZN(
        n19365) );
  AOI22_X1 U22355 ( .A1(P2_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n19373), .B1(
        n19372), .B2(n19680), .ZN(n19364) );
  OAI211_X1 U22356 ( .C1(n19583), .C2(n19405), .A(n19365), .B(n19364), .ZN(
        P2_U3108) );
  AOI22_X1 U22357 ( .A1(n19371), .A2(n19684), .B1(n19382), .B2(n19683), .ZN(
        n19367) );
  AOI22_X1 U22358 ( .A1(P2_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n19373), .B1(
        n19372), .B2(n19686), .ZN(n19366) );
  OAI211_X1 U22359 ( .C1(n19590), .C2(n19405), .A(n19367), .B(n19366), .ZN(
        P2_U3109) );
  AOI22_X1 U22360 ( .A1(n19371), .A2(n19690), .B1(n19382), .B2(n9807), .ZN(
        n19369) );
  AOI22_X1 U22361 ( .A1(P2_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n19373), .B1(
        n19395), .B2(n19692), .ZN(n19368) );
  OAI211_X1 U22362 ( .C1(n19596), .C2(n19370), .A(n19369), .B(n19368), .ZN(
        P2_U3110) );
  AOI22_X1 U22363 ( .A1(n19371), .A2(n19697), .B1(n19382), .B2(n19696), .ZN(
        n19375) );
  AOI22_X1 U22364 ( .A1(P2_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n19373), .B1(
        n19372), .B2(n19699), .ZN(n19374) );
  OAI211_X1 U22365 ( .C1(n19436), .C2(n19405), .A(n19375), .B(n19374), .ZN(
        P2_U3111) );
  NAND2_X1 U22366 ( .A1(n16248), .A2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(
        n19473) );
  NOR2_X1 U22367 ( .A1(n19473), .A2(P2_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(
        n19411) );
  INV_X1 U22368 ( .A(n19411), .ZN(n19414) );
  NOR2_X1 U22369 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19414), .ZN(
        n19400) );
  AOI22_X1 U22370 ( .A1(n19658), .A2(n19431), .B1(n19656), .B2(n19400), .ZN(
        n19386) );
  AOI21_X1 U22371 ( .B1(n19405), .B2(n19430), .A(n19836), .ZN(n19376) );
  NOR2_X1 U22372 ( .A1(n19376), .A2(n19790), .ZN(n19381) );
  OAI21_X1 U22373 ( .B1(n19377), .B2(n19842), .A(n19798), .ZN(n19378) );
  AOI21_X1 U22374 ( .B1(n19381), .B2(n19379), .A(n19378), .ZN(n19380) );
  OAI21_X1 U22375 ( .B1(n19400), .B2(n19380), .A(n19648), .ZN(n19402) );
  OAI21_X1 U22376 ( .B1(n19382), .B2(n19400), .A(n19381), .ZN(n19384) );
  OAI21_X1 U22377 ( .B1(n19377), .B2(n19400), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19383) );
  NAND2_X1 U22378 ( .A1(n19384), .A2(n19383), .ZN(n19401) );
  AOI22_X1 U22379 ( .A1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n19402), .B1(
        n19116), .B2(n19401), .ZN(n19385) );
  OAI211_X1 U22380 ( .C1(n19559), .C2(n19405), .A(n19386), .B(n19385), .ZN(
        P2_U3112) );
  AOI22_X1 U22381 ( .A1(n19663), .A2(n19395), .B1(n19661), .B2(n19400), .ZN(
        n19388) );
  AOI22_X1 U22382 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n19402), .B1(
        n19401), .B2(n19120), .ZN(n19387) );
  OAI211_X1 U22383 ( .C1(n19450), .C2(n19430), .A(n19388), .B(n19387), .ZN(
        P2_U3113) );
  AOI22_X1 U22384 ( .A1(n19668), .A2(n19395), .B1(n19400), .B2(n19666), .ZN(
        n19390) );
  AOI22_X1 U22385 ( .A1(P2_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n19402), .B1(
        n19401), .B2(n19126), .ZN(n19389) );
  OAI211_X1 U22386 ( .C1(n19491), .C2(n19430), .A(n19390), .B(n19389), .ZN(
        P2_U3114) );
  AOI22_X1 U22387 ( .A1(n19674), .A2(n19431), .B1(n19400), .B2(n19671), .ZN(
        n19392) );
  AOI22_X1 U22388 ( .A1(P2_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n19402), .B1(
        n19401), .B2(n19672), .ZN(n19391) );
  OAI211_X1 U22389 ( .C1(n19577), .C2(n19405), .A(n19392), .B(n19391), .ZN(
        P2_U3115) );
  AOI22_X1 U22390 ( .A1(n19680), .A2(n19395), .B1(n19677), .B2(n19400), .ZN(
        n19394) );
  AOI22_X1 U22391 ( .A1(P2_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n19402), .B1(
        n19401), .B2(n19678), .ZN(n19393) );
  OAI211_X1 U22392 ( .C1(n19583), .C2(n19430), .A(n19394), .B(n19393), .ZN(
        P2_U3116) );
  AOI22_X1 U22393 ( .A1(n19686), .A2(n19395), .B1(n19683), .B2(n19400), .ZN(
        n19397) );
  AOI22_X1 U22394 ( .A1(P2_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n19402), .B1(
        n19401), .B2(n19684), .ZN(n19396) );
  OAI211_X1 U22395 ( .C1(n19590), .C2(n19430), .A(n19397), .B(n19396), .ZN(
        P2_U3117) );
  AOI22_X1 U22396 ( .A1(n19692), .A2(n19431), .B1(n9807), .B2(n19400), .ZN(
        n19399) );
  AOI22_X1 U22397 ( .A1(P2_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n19402), .B1(
        n19401), .B2(n19690), .ZN(n19398) );
  OAI211_X1 U22398 ( .C1(n19596), .C2(n19405), .A(n19399), .B(n19398), .ZN(
        P2_U3118) );
  AOI22_X1 U22399 ( .A1(n19701), .A2(n19431), .B1(n19696), .B2(n19400), .ZN(
        n19404) );
  AOI22_X1 U22400 ( .A1(P2_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n19402), .B1(
        n19401), .B2(n19697), .ZN(n19403) );
  OAI211_X1 U22401 ( .C1(n19606), .C2(n19405), .A(n19404), .B(n19403), .ZN(
        P2_U3119) );
  NOR2_X1 U22402 ( .A1(n19406), .A2(n19473), .ZN(n19441) );
  AOI22_X1 U22403 ( .A1(n19657), .A2(n19431), .B1(n19656), .B2(n19441), .ZN(
        n19417) );
  NAND2_X1 U22404 ( .A1(n19407), .A2(P2_STATEBS16_REG_SCAN_IN), .ZN(n19651) );
  OAI21_X1 U22405 ( .B1(n19651), .B2(n19408), .A(n19612), .ZN(n19415) );
  INV_X1 U22406 ( .A(n19441), .ZN(n19409) );
  OAI211_X1 U22407 ( .C1(n10514), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19409), 
        .B(n19790), .ZN(n19410) );
  OAI211_X1 U22408 ( .C1(n19415), .C2(n19411), .A(n19648), .B(n19410), .ZN(
        n19433) );
  OAI21_X1 U22409 ( .B1(n19412), .B2(n19441), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19413) );
  OAI21_X1 U22410 ( .B1(n19415), .B2(n19414), .A(n19413), .ZN(n19432) );
  AOI22_X1 U22411 ( .A1(P2_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n19433), .B1(
        n19116), .B2(n19432), .ZN(n19416) );
  OAI211_X1 U22412 ( .C1(n19484), .C2(n19467), .A(n19417), .B(n19416), .ZN(
        P2_U3120) );
  AOI22_X1 U22413 ( .A1(n19663), .A2(n19431), .B1(n19661), .B2(n19441), .ZN(
        n19419) );
  AOI22_X1 U22414 ( .A1(P2_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n19433), .B1(
        n19120), .B2(n19432), .ZN(n19418) );
  OAI211_X1 U22415 ( .C1(n19450), .C2(n19467), .A(n19419), .B(n19418), .ZN(
        P2_U3121) );
  AOI22_X1 U22416 ( .A1(n19667), .A2(n19457), .B1(n19666), .B2(n19441), .ZN(
        n19421) );
  AOI22_X1 U22417 ( .A1(P2_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n19433), .B1(
        n19126), .B2(n19432), .ZN(n19420) );
  OAI211_X1 U22418 ( .C1(n19571), .C2(n19430), .A(n19421), .B(n19420), .ZN(
        P2_U3122) );
  AOI22_X1 U22419 ( .A1(n19674), .A2(n19457), .B1(n19671), .B2(n19441), .ZN(
        n19423) );
  AOI22_X1 U22420 ( .A1(P2_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n19433), .B1(
        n19672), .B2(n19432), .ZN(n19422) );
  OAI211_X1 U22421 ( .C1(n19577), .C2(n19430), .A(n19423), .B(n19422), .ZN(
        P2_U3123) );
  AOI22_X1 U22422 ( .A1(n19680), .A2(n19431), .B1(n19677), .B2(n19441), .ZN(
        n19425) );
  AOI22_X1 U22423 ( .A1(P2_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n19433), .B1(
        n19678), .B2(n19432), .ZN(n19424) );
  OAI211_X1 U22424 ( .C1(n19583), .C2(n19467), .A(n19425), .B(n19424), .ZN(
        P2_U3124) );
  AOI22_X1 U22425 ( .A1(n19686), .A2(n19431), .B1(n19683), .B2(n19441), .ZN(
        n19427) );
  AOI22_X1 U22426 ( .A1(P2_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n19433), .B1(
        n19684), .B2(n19432), .ZN(n19426) );
  OAI211_X1 U22427 ( .C1(n19590), .C2(n19467), .A(n19427), .B(n19426), .ZN(
        P2_U3125) );
  AOI22_X1 U22428 ( .A1(n19692), .A2(n19457), .B1(n9807), .B2(n19441), .ZN(
        n19429) );
  AOI22_X1 U22429 ( .A1(P2_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n19433), .B1(
        n19690), .B2(n19432), .ZN(n19428) );
  OAI211_X1 U22430 ( .C1(n19596), .C2(n19430), .A(n19429), .B(n19428), .ZN(
        P2_U3126) );
  AOI22_X1 U22431 ( .A1(n19699), .A2(n19431), .B1(n19696), .B2(n19441), .ZN(
        n19435) );
  AOI22_X1 U22432 ( .A1(P2_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n19433), .B1(
        n19697), .B2(n19432), .ZN(n19434) );
  OAI211_X1 U22433 ( .C1(n19436), .C2(n19467), .A(n19435), .B(n19434), .ZN(
        P2_U3127) );
  NOR2_X1 U22434 ( .A1(n19437), .A2(n19473), .ZN(n19462) );
  OAI21_X1 U22435 ( .B1(n19438), .B2(n19462), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19439) );
  OAI21_X1 U22436 ( .B1(n19473), .B2(n19440), .A(n19439), .ZN(n19463) );
  AOI22_X1 U22437 ( .A1(n19463), .A2(n19116), .B1(n19656), .B2(n19462), .ZN(
        n19447) );
  AOI221_X1 U22438 ( .B1(n19499), .B2(P2_STATEBS16_REG_SCAN_IN), .C1(n19457), 
        .C2(P2_STATEBS16_REG_SCAN_IN), .A(n19441), .ZN(n19443) );
  MUX2_X1 U22439 ( .A(n19443), .B(n19442), .S(P2_STATE2_REG_2__SCAN_IN), .Z(
        n19444) );
  NOR2_X1 U22440 ( .A1(n19444), .A2(P2_STATE2_REG_3__SCAN_IN), .ZN(n19445) );
  AOI22_X1 U22441 ( .A1(P2_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n19464), .B1(
        n19499), .B2(n19658), .ZN(n19446) );
  OAI211_X1 U22442 ( .C1(n19559), .C2(n19467), .A(n19447), .B(n19446), .ZN(
        P2_U3128) );
  AOI22_X1 U22443 ( .A1(n19463), .A2(n19120), .B1(n19661), .B2(n19462), .ZN(
        n19449) );
  AOI22_X1 U22444 ( .A1(P2_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n19464), .B1(
        n19457), .B2(n19663), .ZN(n19448) );
  OAI211_X1 U22445 ( .C1(n19450), .C2(n19511), .A(n19449), .B(n19448), .ZN(
        P2_U3129) );
  AOI22_X1 U22446 ( .A1(n19463), .A2(n19126), .B1(n19666), .B2(n19462), .ZN(
        n19452) );
  AOI22_X1 U22447 ( .A1(P2_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n19464), .B1(
        n19457), .B2(n19668), .ZN(n19451) );
  OAI211_X1 U22448 ( .C1(n19491), .C2(n19511), .A(n19452), .B(n19451), .ZN(
        P2_U3130) );
  AOI22_X1 U22449 ( .A1(n19463), .A2(n19672), .B1(n19671), .B2(n19462), .ZN(
        n19454) );
  AOI22_X1 U22450 ( .A1(P2_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n19464), .B1(
        n19499), .B2(n19674), .ZN(n19453) );
  OAI211_X1 U22451 ( .C1(n19577), .C2(n19467), .A(n19454), .B(n19453), .ZN(
        P2_U3131) );
  AOI22_X1 U22452 ( .A1(n19463), .A2(n19678), .B1(n19677), .B2(n19462), .ZN(
        n19456) );
  AOI22_X1 U22453 ( .A1(P2_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n19464), .B1(
        n19457), .B2(n19680), .ZN(n19455) );
  OAI211_X1 U22454 ( .C1(n19583), .C2(n19511), .A(n19456), .B(n19455), .ZN(
        P2_U3132) );
  AOI22_X1 U22455 ( .A1(n19463), .A2(n19684), .B1(n19683), .B2(n19462), .ZN(
        n19459) );
  AOI22_X1 U22456 ( .A1(P2_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n19464), .B1(
        n19457), .B2(n19686), .ZN(n19458) );
  OAI211_X1 U22457 ( .C1(n19590), .C2(n19511), .A(n19459), .B(n19458), .ZN(
        P2_U3133) );
  AOI22_X1 U22458 ( .A1(n19463), .A2(n19690), .B1(n9807), .B2(n19462), .ZN(
        n19461) );
  AOI22_X1 U22459 ( .A1(P2_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n19464), .B1(
        n19499), .B2(n19692), .ZN(n19460) );
  OAI211_X1 U22460 ( .C1(n19596), .C2(n19467), .A(n19461), .B(n19460), .ZN(
        P2_U3134) );
  AOI22_X1 U22461 ( .A1(n19463), .A2(n19697), .B1(n19696), .B2(n19462), .ZN(
        n19466) );
  AOI22_X1 U22462 ( .A1(P2_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n19464), .B1(
        n19499), .B2(n19701), .ZN(n19465) );
  OAI211_X1 U22463 ( .C1(n19606), .C2(n19467), .A(n19466), .B(n19465), .ZN(
        P2_U3135) );
  INV_X1 U22464 ( .A(n19473), .ZN(n19469) );
  AND2_X1 U22465 ( .A1(n19470), .A2(n19469), .ZN(n19481) );
  INV_X1 U22466 ( .A(n19481), .ZN(n19505) );
  NAND2_X1 U22467 ( .A1(n19505), .A2(P2_STATE2_REG_2__SCAN_IN), .ZN(n19471) );
  NOR2_X1 U22468 ( .A1(n19472), .A2(n19471), .ZN(n19477) );
  OR2_X1 U22469 ( .A1(n19814), .A2(n19473), .ZN(n19478) );
  INV_X1 U22470 ( .A(n19478), .ZN(n19474) );
  AOI21_X1 U22471 ( .B1(n19798), .B2(n19474), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19475) );
  OR2_X1 U22472 ( .A1(n19477), .A2(n19475), .ZN(n19506) );
  INV_X1 U22473 ( .A(n19116), .ZN(n19547) );
  INV_X1 U22474 ( .A(n19656), .ZN(n19546) );
  OAI22_X1 U22475 ( .A1(n19506), .A2(n19547), .B1(n19546), .B2(n19505), .ZN(
        n19476) );
  INV_X1 U22476 ( .A(n19476), .ZN(n19483) );
  INV_X1 U22477 ( .A(n19651), .ZN(n19550) );
  NAND2_X1 U22478 ( .A1(n19550), .A2(n19784), .ZN(n19479) );
  AOI21_X1 U22479 ( .B1(n19479), .B2(n19478), .A(n19477), .ZN(n19480) );
  OAI211_X1 U22480 ( .C1(n19481), .C2(n19798), .A(n19480), .B(n19648), .ZN(
        n19508) );
  AOI22_X1 U22481 ( .A1(P2_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n19508), .B1(
        n19499), .B2(n19657), .ZN(n19482) );
  OAI211_X1 U22482 ( .C1(n19484), .C2(n19541), .A(n19483), .B(n19482), .ZN(
        P2_U3136) );
  INV_X1 U22483 ( .A(n19120), .ZN(n19561) );
  INV_X1 U22484 ( .A(n19661), .ZN(n19560) );
  OAI22_X1 U22485 ( .A1(n19506), .A2(n19561), .B1(n19560), .B2(n19505), .ZN(
        n19485) );
  INV_X1 U22486 ( .A(n19485), .ZN(n19487) );
  AOI22_X1 U22487 ( .A1(P2_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n19508), .B1(
        n19531), .B2(n19662), .ZN(n19486) );
  OAI211_X1 U22488 ( .C1(n19565), .C2(n19511), .A(n19487), .B(n19486), .ZN(
        P2_U3137) );
  INV_X1 U22489 ( .A(n19126), .ZN(n19567) );
  INV_X1 U22490 ( .A(n19666), .ZN(n19566) );
  OAI22_X1 U22491 ( .A1(n19506), .A2(n19567), .B1(n19566), .B2(n19505), .ZN(
        n19488) );
  INV_X1 U22492 ( .A(n19488), .ZN(n19490) );
  AOI22_X1 U22493 ( .A1(P2_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n19508), .B1(
        n19499), .B2(n19668), .ZN(n19489) );
  OAI211_X1 U22494 ( .C1(n19491), .C2(n19541), .A(n19490), .B(n19489), .ZN(
        P2_U3138) );
  INV_X1 U22495 ( .A(n19672), .ZN(n19573) );
  INV_X1 U22496 ( .A(n19671), .ZN(n19572) );
  OAI22_X1 U22497 ( .A1(n19506), .A2(n19573), .B1(n19572), .B2(n19505), .ZN(
        n19492) );
  INV_X1 U22498 ( .A(n19492), .ZN(n19494) );
  AOI22_X1 U22499 ( .A1(P2_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n19508), .B1(
        n19531), .B2(n19674), .ZN(n19493) );
  OAI211_X1 U22500 ( .C1(n19577), .C2(n19511), .A(n19494), .B(n19493), .ZN(
        P2_U3139) );
  INV_X1 U22501 ( .A(n19678), .ZN(n19579) );
  OAI22_X1 U22502 ( .A1(n19506), .A2(n19579), .B1(n19578), .B2(n19505), .ZN(
        n19495) );
  INV_X1 U22503 ( .A(n19495), .ZN(n19497) );
  AOI22_X1 U22504 ( .A1(P2_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n19508), .B1(
        n19499), .B2(n19680), .ZN(n19496) );
  OAI211_X1 U22505 ( .C1(n19583), .C2(n19541), .A(n19497), .B(n19496), .ZN(
        P2_U3140) );
  INV_X1 U22506 ( .A(n19684), .ZN(n19585) );
  INV_X1 U22507 ( .A(n19683), .ZN(n19584) );
  OAI22_X1 U22508 ( .A1(n19506), .A2(n19585), .B1(n19584), .B2(n19505), .ZN(
        n19498) );
  INV_X1 U22509 ( .A(n19498), .ZN(n19501) );
  AOI22_X1 U22510 ( .A1(P2_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n19508), .B1(
        n19499), .B2(n19686), .ZN(n19500) );
  OAI211_X1 U22511 ( .C1(n19590), .C2(n19541), .A(n19501), .B(n19500), .ZN(
        P2_U3141) );
  INV_X1 U22512 ( .A(n19690), .ZN(n19592) );
  OAI22_X1 U22514 ( .A1(n19506), .A2(n19592), .B1(n21192), .B2(n19505), .ZN(
        n19502) );
  INV_X1 U22515 ( .A(n19502), .ZN(n19504) );
  AOI22_X1 U22516 ( .A1(P2_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n19508), .B1(
        n19531), .B2(n19692), .ZN(n19503) );
  OAI211_X1 U22517 ( .C1(n19596), .C2(n19511), .A(n19504), .B(n19503), .ZN(
        P2_U3142) );
  INV_X1 U22518 ( .A(n19697), .ZN(n19599) );
  INV_X1 U22519 ( .A(n19696), .ZN(n19598) );
  OAI22_X1 U22520 ( .A1(n19506), .A2(n19599), .B1(n19598), .B2(n19505), .ZN(
        n19507) );
  INV_X1 U22521 ( .A(n19507), .ZN(n19510) );
  AOI22_X1 U22522 ( .A1(P2_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n19508), .B1(
        n19531), .B2(n19701), .ZN(n19509) );
  OAI211_X1 U22523 ( .C1(n19606), .C2(n19511), .A(n19510), .B(n19509), .ZN(
        P2_U3143) );
  INV_X1 U22524 ( .A(n19512), .ZN(n19516) );
  NAND3_X1 U22525 ( .A1(P2_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n19814), .ZN(n19552) );
  NOR2_X1 U22526 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19552), .ZN(
        n19536) );
  OAI21_X1 U22527 ( .B1(n19513), .B2(n19536), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19514) );
  OAI21_X1 U22528 ( .B1(n19516), .B2(n19515), .A(n19514), .ZN(n19537) );
  AOI22_X1 U22529 ( .A1(n19537), .A2(n19116), .B1(n19656), .B2(n19536), .ZN(
        n19522) );
  AOI21_X1 U22530 ( .B1(n19541), .B2(n19605), .A(n19836), .ZN(n19517) );
  AOI21_X1 U22531 ( .B1(n19518), .B2(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A(
        n19517), .ZN(n19520) );
  AOI211_X1 U22532 ( .C1(n19513), .C2(n19798), .A(n19536), .B(n19612), .ZN(
        n19519) );
  AOI22_X1 U22533 ( .A1(P2_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n19538), .B1(
        n19587), .B2(n19658), .ZN(n19521) );
  OAI211_X1 U22534 ( .C1(n19559), .C2(n19541), .A(n19522), .B(n19521), .ZN(
        P2_U3144) );
  AOI22_X1 U22535 ( .A1(n19537), .A2(n19120), .B1(n19661), .B2(n19536), .ZN(
        n19524) );
  AOI22_X1 U22536 ( .A1(P2_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n19538), .B1(
        n19587), .B2(n19662), .ZN(n19523) );
  OAI211_X1 U22537 ( .C1(n19565), .C2(n19541), .A(n19524), .B(n19523), .ZN(
        P2_U3145) );
  AOI22_X1 U22538 ( .A1(n19537), .A2(n19126), .B1(n19666), .B2(n19536), .ZN(
        n19526) );
  AOI22_X1 U22539 ( .A1(P2_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n19538), .B1(
        n19587), .B2(n19667), .ZN(n19525) );
  OAI211_X1 U22540 ( .C1(n19571), .C2(n19541), .A(n19526), .B(n19525), .ZN(
        P2_U3146) );
  AOI22_X1 U22541 ( .A1(n19537), .A2(n19672), .B1(n19671), .B2(n19536), .ZN(
        n19528) );
  AOI22_X1 U22542 ( .A1(P2_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n19538), .B1(
        n19587), .B2(n19674), .ZN(n19527) );
  OAI211_X1 U22543 ( .C1(n19577), .C2(n19541), .A(n19528), .B(n19527), .ZN(
        P2_U3147) );
  AOI22_X1 U22544 ( .A1(n19537), .A2(n19678), .B1(n19677), .B2(n19536), .ZN(
        n19530) );
  AOI22_X1 U22545 ( .A1(P2_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n19538), .B1(
        n19531), .B2(n19680), .ZN(n19529) );
  OAI211_X1 U22546 ( .C1(n19583), .C2(n19605), .A(n19530), .B(n19529), .ZN(
        P2_U3148) );
  AOI22_X1 U22547 ( .A1(n19537), .A2(n19684), .B1(n19683), .B2(n19536), .ZN(
        n19533) );
  AOI22_X1 U22548 ( .A1(P2_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n19538), .B1(
        n19531), .B2(n19686), .ZN(n19532) );
  OAI211_X1 U22549 ( .C1(n19590), .C2(n19605), .A(n19533), .B(n19532), .ZN(
        P2_U3149) );
  AOI22_X1 U22550 ( .A1(n19537), .A2(n19690), .B1(n9807), .B2(n19536), .ZN(
        n19535) );
  AOI22_X1 U22551 ( .A1(P2_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n19538), .B1(
        n19587), .B2(n19692), .ZN(n19534) );
  OAI211_X1 U22552 ( .C1(n19596), .C2(n19541), .A(n19535), .B(n19534), .ZN(
        P2_U3150) );
  AOI22_X1 U22553 ( .A1(n19537), .A2(n19697), .B1(n19696), .B2(n19536), .ZN(
        n19540) );
  AOI22_X1 U22554 ( .A1(P2_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n19538), .B1(
        n19587), .B2(n19701), .ZN(n19539) );
  OAI211_X1 U22555 ( .C1(n19606), .C2(n19541), .A(n19540), .B(n19539), .ZN(
        P2_U3151) );
  NOR2_X1 U22556 ( .A1(n19823), .A2(n19552), .ZN(n19611) );
  INV_X1 U22557 ( .A(n19611), .ZN(n19597) );
  NAND2_X1 U22558 ( .A1(P2_STATE2_REG_2__SCAN_IN), .A2(n19597), .ZN(n19542) );
  NOR2_X1 U22559 ( .A1(n19543), .A2(n19542), .ZN(n19551) );
  INV_X1 U22560 ( .A(n19552), .ZN(n19544) );
  AOI21_X1 U22561 ( .B1(n19798), .B2(n19544), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19545) );
  OR2_X1 U22562 ( .A1(n19551), .A2(n19545), .ZN(n19600) );
  OAI22_X1 U22563 ( .A1(n19600), .A2(n19547), .B1(n19546), .B2(n19597), .ZN(
        n19548) );
  INV_X1 U22564 ( .A(n19548), .ZN(n19558) );
  INV_X1 U22565 ( .A(n19555), .ZN(n19549) );
  NAND2_X1 U22566 ( .A1(n19550), .A2(n19549), .ZN(n19553) );
  AOI21_X1 U22567 ( .B1(n19553), .B2(n19552), .A(n19551), .ZN(n19554) );
  OAI211_X1 U22568 ( .C1(n19611), .C2(n19798), .A(n19554), .B(n19648), .ZN(
        n19602) );
  AOI22_X1 U22569 ( .A1(P2_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n19602), .B1(
        n19641), .B2(n19658), .ZN(n19557) );
  OAI211_X1 U22570 ( .C1(n19559), .C2(n19605), .A(n19558), .B(n19557), .ZN(
        P2_U3152) );
  OAI22_X1 U22571 ( .A1(n19600), .A2(n19561), .B1(n19560), .B2(n19597), .ZN(
        n19562) );
  INV_X1 U22572 ( .A(n19562), .ZN(n19564) );
  AOI22_X1 U22573 ( .A1(P2_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n19602), .B1(
        n19641), .B2(n19662), .ZN(n19563) );
  OAI211_X1 U22574 ( .C1(n19565), .C2(n19605), .A(n19564), .B(n19563), .ZN(
        P2_U3153) );
  OAI22_X1 U22575 ( .A1(n19600), .A2(n19567), .B1(n19566), .B2(n19597), .ZN(
        n19568) );
  INV_X1 U22576 ( .A(n19568), .ZN(n19570) );
  AOI22_X1 U22577 ( .A1(P2_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n19602), .B1(
        n19641), .B2(n19667), .ZN(n19569) );
  OAI211_X1 U22578 ( .C1(n19571), .C2(n19605), .A(n19570), .B(n19569), .ZN(
        P2_U3154) );
  OAI22_X1 U22579 ( .A1(n19600), .A2(n19573), .B1(n19572), .B2(n19597), .ZN(
        n19574) );
  INV_X1 U22580 ( .A(n19574), .ZN(n19576) );
  AOI22_X1 U22581 ( .A1(P2_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n19602), .B1(
        n19641), .B2(n19674), .ZN(n19575) );
  OAI211_X1 U22582 ( .C1(n19577), .C2(n19605), .A(n19576), .B(n19575), .ZN(
        P2_U3155) );
  OAI22_X1 U22583 ( .A1(n19600), .A2(n19579), .B1(n19578), .B2(n19597), .ZN(
        n19580) );
  INV_X1 U22584 ( .A(n19580), .ZN(n19582) );
  AOI22_X1 U22585 ( .A1(P2_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n19602), .B1(
        n19587), .B2(n19680), .ZN(n19581) );
  OAI211_X1 U22586 ( .C1(n19583), .C2(n19608), .A(n19582), .B(n19581), .ZN(
        P2_U3156) );
  OAI22_X1 U22587 ( .A1(n19600), .A2(n19585), .B1(n19584), .B2(n19597), .ZN(
        n19586) );
  INV_X1 U22588 ( .A(n19586), .ZN(n19589) );
  AOI22_X1 U22589 ( .A1(P2_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n19602), .B1(
        n19587), .B2(n19686), .ZN(n19588) );
  OAI211_X1 U22590 ( .C1(n19590), .C2(n19608), .A(n19589), .B(n19588), .ZN(
        P2_U3157) );
  OAI22_X1 U22591 ( .A1(n19600), .A2(n19592), .B1(n21192), .B2(n19597), .ZN(
        n19593) );
  INV_X1 U22592 ( .A(n19593), .ZN(n19595) );
  AOI22_X1 U22593 ( .A1(P2_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n19602), .B1(
        n19641), .B2(n19692), .ZN(n19594) );
  OAI211_X1 U22594 ( .C1(n19596), .C2(n19605), .A(n19595), .B(n19594), .ZN(
        P2_U3158) );
  OAI22_X1 U22595 ( .A1(n19600), .A2(n19599), .B1(n19598), .B2(n19597), .ZN(
        n19601) );
  INV_X1 U22596 ( .A(n19601), .ZN(n19604) );
  AOI22_X1 U22597 ( .A1(P2_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n19602), .B1(
        n19641), .B2(n19701), .ZN(n19603) );
  OAI211_X1 U22598 ( .C1(n19606), .C2(n19605), .A(n19604), .B(n19603), .ZN(
        P2_U3159) );
  NAND2_X1 U22599 ( .A1(n19615), .A2(n19608), .ZN(n19609) );
  AOI21_X1 U22600 ( .B1(n19609), .B2(P2_STATEBS16_REG_SCAN_IN), .A(n19790), 
        .ZN(n19616) );
  NAND2_X1 U22601 ( .A1(P2_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n19610), .ZN(
        n19652) );
  NOR2_X1 U22602 ( .A1(P2_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n19652), .ZN(
        n19640) );
  NOR2_X1 U22603 ( .A1(n19640), .A2(n19611), .ZN(n19619) );
  AOI211_X1 U22604 ( .C1(n19617), .C2(n19798), .A(n19640), .B(n19612), .ZN(
        n19614) );
  INV_X1 U22605 ( .A(P2_INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n19623) );
  AOI22_X1 U22606 ( .A1(n19658), .A2(n19700), .B1(n19640), .B2(n19656), .ZN(
        n19622) );
  INV_X1 U22607 ( .A(n19616), .ZN(n19620) );
  OAI21_X1 U22608 ( .B1(n19617), .B2(n19640), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19618) );
  AOI22_X1 U22609 ( .A1(n19116), .A2(n19642), .B1(n19641), .B2(n19657), .ZN(
        n19621) );
  OAI211_X1 U22610 ( .C1(n19646), .C2(n19623), .A(n19622), .B(n19621), .ZN(
        P2_U3160) );
  AOI22_X1 U22611 ( .A1(n19663), .A2(n19641), .B1(n19640), .B2(n19661), .ZN(
        n19625) );
  AOI22_X1 U22612 ( .A1(n19120), .A2(n19642), .B1(n19700), .B2(n19662), .ZN(
        n19624) );
  OAI211_X1 U22613 ( .C1(n19646), .C2(n10529), .A(n19625), .B(n19624), .ZN(
        P2_U3161) );
  INV_X1 U22614 ( .A(P2_INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n19628) );
  AOI22_X1 U22615 ( .A1(n19668), .A2(n19641), .B1(n19640), .B2(n19666), .ZN(
        n19627) );
  AOI22_X1 U22616 ( .A1(n19126), .A2(n19642), .B1(n19700), .B2(n19667), .ZN(
        n19626) );
  OAI211_X1 U22617 ( .C1(n19646), .C2(n19628), .A(n19627), .B(n19626), .ZN(
        P2_U3162) );
  INV_X1 U22618 ( .A(P2_INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n19631) );
  AOI22_X1 U22619 ( .A1(n19674), .A2(n19700), .B1(n19640), .B2(n19671), .ZN(
        n19630) );
  AOI22_X1 U22620 ( .A1(n19672), .A2(n19642), .B1(n19641), .B2(n19673), .ZN(
        n19629) );
  OAI211_X1 U22621 ( .C1(n19646), .C2(n19631), .A(n19630), .B(n19629), .ZN(
        P2_U3163) );
  INV_X1 U22622 ( .A(P2_INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n20902) );
  AOI22_X1 U22623 ( .A1(n19679), .A2(n19700), .B1(n19677), .B2(n19640), .ZN(
        n19633) );
  AOI22_X1 U22624 ( .A1(n19678), .A2(n19642), .B1(n19641), .B2(n19680), .ZN(
        n19632) );
  OAI211_X1 U22625 ( .C1(n19646), .C2(n20902), .A(n19633), .B(n19632), .ZN(
        P2_U3164) );
  INV_X1 U22626 ( .A(P2_INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n19636) );
  AOI22_X1 U22627 ( .A1(n19685), .A2(n19700), .B1(n19640), .B2(n19683), .ZN(
        n19635) );
  AOI22_X1 U22628 ( .A1(n19684), .A2(n19642), .B1(n19641), .B2(n19686), .ZN(
        n19634) );
  OAI211_X1 U22629 ( .C1(n19646), .C2(n19636), .A(n19635), .B(n19634), .ZN(
        P2_U3165) );
  INV_X1 U22630 ( .A(P2_INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n19639) );
  AOI22_X1 U22631 ( .A1(n19692), .A2(n19700), .B1(n19640), .B2(n9807), .ZN(
        n19638) );
  AOI22_X1 U22632 ( .A1(n19690), .A2(n19642), .B1(n19641), .B2(n19691), .ZN(
        n19637) );
  OAI211_X1 U22633 ( .C1(n19646), .C2(n19639), .A(n19638), .B(n19637), .ZN(
        P2_U3166) );
  INV_X1 U22634 ( .A(P2_INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n19645) );
  AOI22_X1 U22635 ( .A1(n19701), .A2(n19700), .B1(n19640), .B2(n19696), .ZN(
        n19644) );
  AOI22_X1 U22636 ( .A1(n19697), .A2(n19642), .B1(n19641), .B2(n19699), .ZN(
        n19643) );
  OAI211_X1 U22637 ( .C1(n19646), .C2(n19645), .A(n19644), .B(n19643), .ZN(
        P2_U3167) );
  NOR3_X1 U22638 ( .A1(n19647), .A2(n19695), .A3(n19842), .ZN(n19655) );
  INV_X1 U22639 ( .A(n19655), .ZN(n19649) );
  OAI211_X1 U22640 ( .C1(n19695), .C2(n19798), .A(n19649), .B(n19648), .ZN(
        n19650) );
  AOI221_X2 U22641 ( .B1(n19789), .B2(n19652), .C1(n19651), .C2(n19652), .A(
        n19650), .ZN(n19706) );
  INV_X1 U22642 ( .A(P2_INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n21028) );
  INV_X1 U22643 ( .A(n19652), .ZN(n19653) );
  AOI21_X1 U22644 ( .B1(n19798), .B2(n19653), .A(P2_STATE2_REG_2__SCAN_IN), 
        .ZN(n19654) );
  NOR2_X1 U22645 ( .A1(n19655), .A2(n19654), .ZN(n19698) );
  AOI22_X1 U22646 ( .A1(n19698), .A2(n19116), .B1(n19656), .B2(n19695), .ZN(
        n19660) );
  AOI22_X1 U22647 ( .A1(n19702), .A2(n19658), .B1(n19700), .B2(n19657), .ZN(
        n19659) );
  OAI211_X1 U22648 ( .C1(n19706), .C2(n21028), .A(n19660), .B(n19659), .ZN(
        P2_U3168) );
  AOI22_X1 U22649 ( .A1(n19698), .A2(n19120), .B1(n19661), .B2(n19695), .ZN(
        n19665) );
  AOI22_X1 U22650 ( .A1(n19700), .A2(n19663), .B1(n19702), .B2(n19662), .ZN(
        n19664) );
  OAI211_X1 U22651 ( .C1(n19706), .C2(n13013), .A(n19665), .B(n19664), .ZN(
        P2_U3169) );
  AOI22_X1 U22652 ( .A1(n19698), .A2(n19126), .B1(n19666), .B2(n19695), .ZN(
        n19670) );
  AOI22_X1 U22653 ( .A1(n19700), .A2(n19668), .B1(n19702), .B2(n19667), .ZN(
        n19669) );
  OAI211_X1 U22654 ( .C1(n19706), .C2(n13042), .A(n19670), .B(n19669), .ZN(
        P2_U3170) );
  AOI22_X1 U22655 ( .A1(n19698), .A2(n19672), .B1(n19671), .B2(n19695), .ZN(
        n19676) );
  AOI22_X1 U22656 ( .A1(n19702), .A2(n19674), .B1(n19700), .B2(n19673), .ZN(
        n19675) );
  OAI211_X1 U22657 ( .C1(n19706), .C2(n13069), .A(n19676), .B(n19675), .ZN(
        P2_U3171) );
  AOI22_X1 U22658 ( .A1(n19698), .A2(n19678), .B1(n19677), .B2(n19695), .ZN(
        n19682) );
  AOI22_X1 U22659 ( .A1(n19700), .A2(n19680), .B1(n19702), .B2(n19679), .ZN(
        n19681) );
  OAI211_X1 U22660 ( .C1(n19706), .C2(n13093), .A(n19682), .B(n19681), .ZN(
        P2_U3172) );
  AOI22_X1 U22661 ( .A1(n19698), .A2(n19684), .B1(n19683), .B2(n19695), .ZN(
        n19688) );
  AOI22_X1 U22662 ( .A1(n19700), .A2(n19686), .B1(n19702), .B2(n19685), .ZN(
        n19687) );
  OAI211_X1 U22663 ( .C1(n19706), .C2(n13124), .A(n19688), .B(n19687), .ZN(
        P2_U3173) );
  AOI22_X1 U22664 ( .A1(n19698), .A2(n19690), .B1(n9807), .B2(n19695), .ZN(
        n19694) );
  AOI22_X1 U22665 ( .A1(n19702), .A2(n19692), .B1(n19700), .B2(n19691), .ZN(
        n19693) );
  OAI211_X1 U22666 ( .C1(n19706), .C2(n13151), .A(n19694), .B(n19693), .ZN(
        P2_U3174) );
  INV_X1 U22667 ( .A(P2_INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n19705) );
  AOI22_X1 U22668 ( .A1(n19698), .A2(n19697), .B1(n19696), .B2(n19695), .ZN(
        n19704) );
  AOI22_X1 U22669 ( .A1(n19702), .A2(n19701), .B1(n19700), .B2(n19699), .ZN(
        n19703) );
  OAI211_X1 U22670 ( .C1(n19706), .C2(n19705), .A(n19704), .B(n19703), .ZN(
        P2_U3175) );
  AOI211_X1 U22671 ( .C1(n19843), .C2(n19842), .A(n19708), .B(n19707), .ZN(
        n19712) );
  NAND2_X1 U22672 ( .A1(P2_STATE2_REG_1__SCAN_IN), .A2(n19843), .ZN(n19709) );
  AOI21_X1 U22673 ( .B1(n19710), .B2(n19713), .A(n19709), .ZN(n19711) );
  AOI21_X1 U22674 ( .B1(n19713), .B2(n19712), .A(n19711), .ZN(n19715) );
  NAND2_X1 U22675 ( .A1(n19715), .A2(n19714), .ZN(P2_U3177) );
  AND2_X1 U22676 ( .A1(P2_DATAWIDTH_REG_31__SCAN_IN), .A2(n19716), .ZN(
        P2_U3179) );
  AND2_X1 U22677 ( .A1(P2_DATAWIDTH_REG_30__SCAN_IN), .A2(n19716), .ZN(
        P2_U3180) );
  AND2_X1 U22678 ( .A1(P2_DATAWIDTH_REG_29__SCAN_IN), .A2(n19716), .ZN(
        P2_U3181) );
  AND2_X1 U22679 ( .A1(P2_DATAWIDTH_REG_28__SCAN_IN), .A2(n19716), .ZN(
        P2_U3182) );
  AND2_X1 U22680 ( .A1(P2_DATAWIDTH_REG_27__SCAN_IN), .A2(n19716), .ZN(
        P2_U3183) );
  AND2_X1 U22681 ( .A1(P2_DATAWIDTH_REG_26__SCAN_IN), .A2(n19716), .ZN(
        P2_U3184) );
  AND2_X1 U22682 ( .A1(P2_DATAWIDTH_REG_25__SCAN_IN), .A2(n19716), .ZN(
        P2_U3185) );
  INV_X1 U22683 ( .A(P2_DATAWIDTH_REG_24__SCAN_IN), .ZN(n21081) );
  NOR2_X1 U22684 ( .A1(n21081), .A2(n19783), .ZN(P2_U3186) );
  AND2_X1 U22685 ( .A1(P2_DATAWIDTH_REG_23__SCAN_IN), .A2(n19716), .ZN(
        P2_U3187) );
  AND2_X1 U22686 ( .A1(P2_DATAWIDTH_REG_22__SCAN_IN), .A2(n19716), .ZN(
        P2_U3188) );
  INV_X1 U22687 ( .A(P2_DATAWIDTH_REG_21__SCAN_IN), .ZN(n20931) );
  NOR2_X1 U22688 ( .A1(n20931), .A2(n19783), .ZN(P2_U3189) );
  AND2_X1 U22689 ( .A1(P2_DATAWIDTH_REG_20__SCAN_IN), .A2(n19716), .ZN(
        P2_U3190) );
  AND2_X1 U22690 ( .A1(P2_DATAWIDTH_REG_19__SCAN_IN), .A2(n19716), .ZN(
        P2_U3191) );
  NOR2_X1 U22691 ( .A1(n21068), .A2(n19783), .ZN(P2_U3192) );
  AND2_X1 U22692 ( .A1(P2_DATAWIDTH_REG_17__SCAN_IN), .A2(n19716), .ZN(
        P2_U3193) );
  AND2_X1 U22693 ( .A1(P2_DATAWIDTH_REG_16__SCAN_IN), .A2(n19716), .ZN(
        P2_U3194) );
  AND2_X1 U22694 ( .A1(P2_DATAWIDTH_REG_15__SCAN_IN), .A2(n19716), .ZN(
        P2_U3195) );
  AND2_X1 U22695 ( .A1(P2_DATAWIDTH_REG_14__SCAN_IN), .A2(n19716), .ZN(
        P2_U3196) );
  AND2_X1 U22696 ( .A1(P2_DATAWIDTH_REG_13__SCAN_IN), .A2(n19716), .ZN(
        P2_U3197) );
  AND2_X1 U22697 ( .A1(P2_DATAWIDTH_REG_12__SCAN_IN), .A2(n19716), .ZN(
        P2_U3198) );
  AND2_X1 U22698 ( .A1(P2_DATAWIDTH_REG_11__SCAN_IN), .A2(n19716), .ZN(
        P2_U3199) );
  AND2_X1 U22699 ( .A1(P2_DATAWIDTH_REG_10__SCAN_IN), .A2(n19716), .ZN(
        P2_U3200) );
  AND2_X1 U22700 ( .A1(P2_DATAWIDTH_REG_9__SCAN_IN), .A2(n19716), .ZN(P2_U3201) );
  AND2_X1 U22701 ( .A1(P2_DATAWIDTH_REG_8__SCAN_IN), .A2(n19716), .ZN(P2_U3202) );
  AND2_X1 U22702 ( .A1(P2_DATAWIDTH_REG_7__SCAN_IN), .A2(n19716), .ZN(P2_U3203) );
  AND2_X1 U22703 ( .A1(P2_DATAWIDTH_REG_6__SCAN_IN), .A2(n19716), .ZN(P2_U3204) );
  AND2_X1 U22704 ( .A1(P2_DATAWIDTH_REG_5__SCAN_IN), .A2(n19716), .ZN(P2_U3205) );
  NOR2_X1 U22705 ( .A1(n20921), .A2(n19783), .ZN(P2_U3206) );
  AND2_X1 U22706 ( .A1(P2_DATAWIDTH_REG_3__SCAN_IN), .A2(n19716), .ZN(P2_U3207) );
  AND2_X1 U22707 ( .A1(P2_DATAWIDTH_REG_2__SCAN_IN), .A2(n19716), .ZN(P2_U3208) );
  NAND2_X1 U22708 ( .A1(P2_STATE_REG_1__SCAN_IN), .A2(n19843), .ZN(n19729) );
  NAND3_X1 U22709 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(
        P2_STATE_REG_0__SCAN_IN), .A3(n19729), .ZN(n19718) );
  AOI211_X1 U22710 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(n20700), .A(
        n19728), .B(n19853), .ZN(n19717) );
  INV_X1 U22711 ( .A(NA), .ZN(n20705) );
  NOR2_X1 U22712 ( .A1(n20705), .A2(n19722), .ZN(n19734) );
  AOI211_X1 U22713 ( .C1(n19735), .C2(n19718), .A(n19717), .B(n19734), .ZN(
        n19719) );
  INV_X1 U22714 ( .A(n19719), .ZN(P2_U3209) );
  INV_X1 U22715 ( .A(P2_REQUESTPENDING_REG_SCAN_IN), .ZN(n19720) );
  AOI21_X1 U22716 ( .B1(P2_STATE_REG_0__SCAN_IN), .B2(n20700), .A(n19735), 
        .ZN(n19726) );
  NOR2_X1 U22717 ( .A1(n19720), .A2(n19726), .ZN(n19723) );
  AOI21_X1 U22718 ( .B1(n19723), .B2(n19722), .A(n19721), .ZN(n19724) );
  OAI211_X1 U22719 ( .C1(n20700), .C2(n19725), .A(n19724), .B(n19729), .ZN(
        P2_U3210) );
  AOI21_X1 U22720 ( .B1(n19843), .B2(n19727), .A(n19726), .ZN(n19733) );
  INV_X1 U22721 ( .A(n19728), .ZN(n19730) );
  OAI22_X1 U22722 ( .A1(P2_REQUESTPENDING_REG_SCAN_IN), .A2(n19730), .B1(NA), 
        .B2(n19729), .ZN(n19731) );
  OAI211_X1 U22723 ( .C1(P2_REQUESTPENDING_REG_SCAN_IN), .C2(HOLD), .A(
        P2_STATE_REG_0__SCAN_IN), .B(n19731), .ZN(n19732) );
  OAI21_X1 U22724 ( .B1(n19734), .B2(n19733), .A(n19732), .ZN(P2_U3211) );
  OAI222_X1 U22725 ( .A1(n19775), .A2(n10480), .B1(n19736), .B2(n19853), .C1(
        n10425), .C2(n19772), .ZN(P2_U3212) );
  OAI222_X1 U22726 ( .A1(n19775), .A2(n12690), .B1(n19737), .B2(n19853), .C1(
        n10480), .C2(n19772), .ZN(P2_U3213) );
  OAI222_X1 U22727 ( .A1(n19775), .A2(n12700), .B1(n19738), .B2(n19853), .C1(
        n12690), .C2(n19772), .ZN(P2_U3214) );
  OAI222_X1 U22728 ( .A1(n19775), .A2(n10904), .B1(n21095), .B2(n19853), .C1(
        n12700), .C2(n19772), .ZN(P2_U3215) );
  OAI222_X1 U22729 ( .A1(n19775), .A2(n10912), .B1(n19739), .B2(n19853), .C1(
        n10904), .C2(n19772), .ZN(P2_U3216) );
  OAI222_X1 U22730 ( .A1(n19775), .A2(n10916), .B1(n20893), .B2(n19853), .C1(
        n10912), .C2(n19772), .ZN(P2_U3217) );
  OAI222_X1 U22731 ( .A1(n19775), .A2(n14050), .B1(n19740), .B2(n19853), .C1(
        n10916), .C2(n19772), .ZN(P2_U3218) );
  OAI222_X1 U22732 ( .A1(n19775), .A2(n14218), .B1(n19741), .B2(n19853), .C1(
        n14050), .C2(n19772), .ZN(P2_U3219) );
  OAI222_X1 U22733 ( .A1(n19775), .A2(n12751), .B1(n19742), .B2(n19853), .C1(
        n14218), .C2(n19772), .ZN(P2_U3220) );
  OAI222_X1 U22734 ( .A1(n19775), .A2(n12765), .B1(n19743), .B2(n19853), .C1(
        n12751), .C2(n19772), .ZN(P2_U3221) );
  OAI222_X1 U22735 ( .A1(n19775), .A2(n12779), .B1(n21030), .B2(n19853), .C1(
        n12765), .C2(n19772), .ZN(P2_U3222) );
  OAI222_X1 U22736 ( .A1(n19775), .A2(n12793), .B1(n19744), .B2(n19853), .C1(
        n12779), .C2(n19772), .ZN(P2_U3223) );
  OAI222_X1 U22737 ( .A1(n19775), .A2(n14023), .B1(n19745), .B2(n19853), .C1(
        n12793), .C2(n19772), .ZN(P2_U3224) );
  OAI222_X1 U22738 ( .A1(n19775), .A2(n19747), .B1(n19746), .B2(n19853), .C1(
        n14023), .C2(n19772), .ZN(P2_U3225) );
  OAI222_X1 U22739 ( .A1(n19775), .A2(n15415), .B1(n19748), .B2(n19853), .C1(
        n19747), .C2(n19772), .ZN(P2_U3226) );
  OAI222_X1 U22740 ( .A1(n19775), .A2(n19750), .B1(n19749), .B2(n19853), .C1(
        n15415), .C2(n19772), .ZN(P2_U3227) );
  OAI222_X1 U22741 ( .A1(n19775), .A2(n19752), .B1(n19751), .B2(n19853), .C1(
        n19750), .C2(n19772), .ZN(P2_U3228) );
  OAI222_X1 U22742 ( .A1(n19775), .A2(n19754), .B1(n19753), .B2(n19853), .C1(
        n19752), .C2(n19772), .ZN(P2_U3229) );
  OAI222_X1 U22743 ( .A1(n19775), .A2(n19756), .B1(n19755), .B2(n19853), .C1(
        n19754), .C2(n19772), .ZN(P2_U3230) );
  OAI222_X1 U22744 ( .A1(n19775), .A2(n19758), .B1(n19757), .B2(n19853), .C1(
        n19756), .C2(n19772), .ZN(P2_U3231) );
  OAI222_X1 U22745 ( .A1(n19775), .A2(n12830), .B1(n19759), .B2(n19853), .C1(
        n19758), .C2(n19772), .ZN(P2_U3232) );
  OAI222_X1 U22746 ( .A1(n19775), .A2(n10960), .B1(n19760), .B2(n19853), .C1(
        n12830), .C2(n19772), .ZN(P2_U3233) );
  OAI222_X1 U22747 ( .A1(n19775), .A2(n10963), .B1(n19761), .B2(n19853), .C1(
        n10960), .C2(n19772), .ZN(P2_U3234) );
  OAI222_X1 U22748 ( .A1(n19775), .A2(n19763), .B1(n19762), .B2(n19853), .C1(
        n10963), .C2(n19772), .ZN(P2_U3235) );
  OAI222_X1 U22749 ( .A1(n19775), .A2(n21017), .B1(n19764), .B2(n19853), .C1(
        n19763), .C2(n19772), .ZN(P2_U3236) );
  OAI222_X1 U22750 ( .A1(n19775), .A2(n19767), .B1(n19765), .B2(n19853), .C1(
        n21017), .C2(n19772), .ZN(P2_U3237) );
  OAI222_X1 U22751 ( .A1(n19772), .A2(n19767), .B1(n19766), .B2(n19853), .C1(
        n19768), .C2(n19775), .ZN(P2_U3238) );
  INV_X1 U22752 ( .A(P2_ADDRESS_REG_27__SCAN_IN), .ZN(n19769) );
  OAI222_X1 U22753 ( .A1(n19775), .A2(n19770), .B1(n19769), .B2(n19853), .C1(
        n19768), .C2(n19772), .ZN(P2_U3239) );
  OAI222_X1 U22754 ( .A1(n19775), .A2(n12844), .B1(n19771), .B2(n19853), .C1(
        n19770), .C2(n19772), .ZN(P2_U3240) );
  INV_X1 U22755 ( .A(P2_REIP_REG_31__SCAN_IN), .ZN(n19774) );
  OAI222_X1 U22756 ( .A1(n19775), .A2(n19774), .B1(n19773), .B2(n19853), .C1(
        n12844), .C2(n19772), .ZN(P2_U3241) );
  OAI22_X1 U22757 ( .A1(n19854), .A2(P2_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P2_BE_N_REG_3__SCAN_IN), .B2(n19853), .ZN(n19776) );
  INV_X1 U22758 ( .A(n19776), .ZN(P2_U3585) );
  OAI22_X1 U22759 ( .A1(n19854), .A2(P2_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P2_BE_N_REG_2__SCAN_IN), .B2(n19853), .ZN(n19777) );
  INV_X1 U22760 ( .A(n19777), .ZN(P2_U3586) );
  OAI22_X1 U22761 ( .A1(n19854), .A2(P2_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P2_BE_N_REG_1__SCAN_IN), .B2(n19853), .ZN(n19778) );
  INV_X1 U22762 ( .A(n19778), .ZN(P2_U3587) );
  OAI22_X1 U22763 ( .A1(n19854), .A2(P2_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P2_BE_N_REG_0__SCAN_IN), .B2(n19853), .ZN(n19779) );
  INV_X1 U22764 ( .A(n19779), .ZN(P2_U3588) );
  OAI21_X1 U22765 ( .B1(n19783), .B2(P2_DATAWIDTH_REG_0__SCAN_IN), .A(n19781), 
        .ZN(n19780) );
  INV_X1 U22766 ( .A(n19780), .ZN(P2_U3591) );
  OAI21_X1 U22767 ( .B1(n19783), .B2(n19782), .A(n19781), .ZN(P2_U3592) );
  INV_X1 U22768 ( .A(n19822), .ZN(n19821) );
  NOR2_X1 U22769 ( .A1(n19790), .A2(n19836), .ZN(n19809) );
  NAND2_X1 U22770 ( .A1(n19784), .A2(n19809), .ZN(n19800) );
  NAND3_X1 U22771 ( .A1(n19786), .A2(n19785), .A3(P2_STATEBS16_REG_SCAN_IN), 
        .ZN(n19787) );
  NAND2_X1 U22772 ( .A1(n19787), .A2(n19806), .ZN(n19797) );
  AOI21_X1 U22773 ( .B1(n19800), .B2(n19797), .A(n19788), .ZN(n19793) );
  NOR3_X1 U22774 ( .A1(n19791), .A2(n19790), .A3(n19789), .ZN(n19792) );
  AOI211_X1 U22775 ( .C1(n19794), .C2(P2_STATE2_REG_3__SCAN_IN), .A(n19793), 
        .B(n19792), .ZN(n19795) );
  AOI22_X1 U22776 ( .A1(n19821), .A2(n19796), .B1(n19795), .B2(n19822), .ZN(
        P2_U3602) );
  INV_X1 U22777 ( .A(n19797), .ZN(n19803) );
  NOR2_X1 U22778 ( .A1(n19799), .A2(n19798), .ZN(n19802) );
  INV_X1 U22779 ( .A(n19800), .ZN(n19801) );
  AOI211_X1 U22780 ( .C1(n19804), .C2(n19803), .A(n19802), .B(n19801), .ZN(
        n19805) );
  AOI22_X1 U22781 ( .A1(n19821), .A2(n16248), .B1(n19805), .B2(n19822), .ZN(
        P2_U3603) );
  INV_X1 U22782 ( .A(n19806), .ZN(n19817) );
  NOR2_X1 U22783 ( .A1(n19817), .A2(n19807), .ZN(n19810) );
  MUX2_X1 U22784 ( .A(n19810), .B(n19809), .S(n19808), .Z(n19811) );
  AOI21_X1 U22785 ( .B1(P2_STATE2_REG_3__SCAN_IN), .B2(n19812), .A(n19811), 
        .ZN(n19813) );
  AOI22_X1 U22786 ( .A1(n19821), .A2(n19814), .B1(n19813), .B2(n19822), .ZN(
        P2_U3604) );
  OAI22_X1 U22787 ( .A1(n19818), .A2(n19817), .B1(n19816), .B2(n19815), .ZN(
        n19819) );
  AOI21_X1 U22788 ( .B1(n19823), .B2(P2_STATE2_REG_3__SCAN_IN), .A(n19819), 
        .ZN(n19820) );
  OAI22_X1 U22789 ( .A1(n19823), .A2(n19822), .B1(n19821), .B2(n19820), .ZN(
        P2_U3605) );
  INV_X1 U22790 ( .A(P2_W_R_N_REG_SCAN_IN), .ZN(n19824) );
  AOI22_X1 U22791 ( .A1(n19853), .A2(P2_READREQUEST_REG_SCAN_IN), .B1(n19824), 
        .B2(n19854), .ZN(P2_U3608) );
  INV_X1 U22792 ( .A(n19825), .ZN(n19829) );
  INV_X1 U22793 ( .A(n19826), .ZN(n19828) );
  AOI22_X1 U22794 ( .A1(n19830), .A2(n19829), .B1(n19828), .B2(n19827), .ZN(
        n19831) );
  NAND2_X1 U22795 ( .A1(n19832), .A2(n19831), .ZN(n19834) );
  MUX2_X1 U22796 ( .A(P2_MORE_REG_SCAN_IN), .B(n19834), .S(n19833), .Z(
        P2_U3609) );
  OAI21_X1 U22797 ( .B1(n19836), .B2(n19837), .A(n19835), .ZN(n19840) );
  NAND3_X1 U22798 ( .A1(n19838), .A2(P2_STATE2_REG_0__SCAN_IN), .A3(n19837), 
        .ZN(n19839) );
  MUX2_X1 U22799 ( .A(n19840), .B(n19839), .S(n12668), .Z(n19845) );
  OAI21_X1 U22800 ( .B1(n19843), .B2(n19842), .A(n19841), .ZN(n19844) );
  NAND2_X1 U22801 ( .A1(n19845), .A2(n19844), .ZN(n19852) );
  AOI21_X1 U22802 ( .B1(P2_STATE2_REG_2__SCAN_IN), .B2(n19846), .A(
        P2_STATE2_REG_3__SCAN_IN), .ZN(n19848) );
  AOI211_X1 U22803 ( .C1(n19850), .C2(n19849), .A(n19848), .B(n19847), .ZN(
        n19851) );
  MUX2_X1 U22804 ( .A(n19852), .B(P2_REQUESTPENDING_REG_SCAN_IN), .S(n19851), 
        .Z(P2_U3610) );
  OAI22_X1 U22805 ( .A1(n19854), .A2(P2_MEMORYFETCH_REG_SCAN_IN), .B1(
        P2_M_IO_N_REG_SCAN_IN), .B2(n19853), .ZN(n19855) );
  INV_X1 U22806 ( .A(n19855), .ZN(P2_U3611) );
  AOI21_X1 U22807 ( .B1(P1_STATE_REG_1__SCAN_IN), .B2(n11119), .A(n20699), 
        .ZN(n20701) );
  INV_X1 U22808 ( .A(P1_ADS_N_REG_SCAN_IN), .ZN(n19856) );
  AND2_X1 U22809 ( .A1(n20699), .A2(P1_STATE_REG_1__SCAN_IN), .ZN(n20786) );
  AOI21_X1 U22810 ( .B1(n20701), .B2(n19856), .A(n20786), .ZN(P1_U2802) );
  OAI21_X1 U22811 ( .B1(n19858), .B2(n19857), .A(P1_CODEFETCH_REG_SCAN_IN), 
        .ZN(n19859) );
  OAI21_X1 U22812 ( .B1(n19860), .B2(n11192), .A(n19859), .ZN(P1_U2803) );
  INV_X1 U22813 ( .A(n20786), .ZN(n20784) );
  NOR2_X1 U22814 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(P1_STATE_REG_0__SCAN_IN), 
        .ZN(n19862) );
  INV_X1 U22815 ( .A(n20786), .ZN(n20798) );
  OAI21_X1 U22816 ( .B1(n19862), .B2(P1_D_C_N_REG_SCAN_IN), .A(n20798), .ZN(
        n19861) );
  OAI21_X1 U22817 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(n20784), .A(n19861), 
        .ZN(P1_U2804) );
  NOR2_X1 U22818 ( .A1(n20701), .A2(n20786), .ZN(n20756) );
  OAI21_X1 U22819 ( .B1(BS16), .B2(n19862), .A(n20756), .ZN(n20754) );
  OAI21_X1 U22820 ( .B1(n20756), .B2(n20765), .A(n20754), .ZN(P1_U2805) );
  OAI21_X1 U22821 ( .B1(n19865), .B2(n19864), .A(n19863), .ZN(P1_U2806) );
  NOR4_X1 U22822 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_20__SCAN_IN), .A3(P1_DATAWIDTH_REG_22__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_23__SCAN_IN), .ZN(n19869) );
  NOR4_X1 U22823 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_16__SCAN_IN), .A3(P1_DATAWIDTH_REG_17__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_18__SCAN_IN), .ZN(n19868) );
  NOR4_X1 U22824 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_29__SCAN_IN), .A3(P1_DATAWIDTH_REG_30__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_31__SCAN_IN), .ZN(n19867) );
  NOR4_X1 U22825 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_25__SCAN_IN), .A3(P1_DATAWIDTH_REG_26__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_27__SCAN_IN), .ZN(n19866) );
  NAND4_X1 U22826 ( .A1(n19869), .A2(n19868), .A3(n19867), .A4(n19866), .ZN(
        n19875) );
  NOR4_X1 U22827 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_3__SCAN_IN), .A3(P1_DATAWIDTH_REG_4__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_5__SCAN_IN), .ZN(n19873) );
  AOI211_X1 U22828 ( .C1(P1_DATAWIDTH_REG_1__SCAN_IN), .C2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_21__SCAN_IN), .B(
        P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n19872) );
  NOR4_X1 U22829 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_12__SCAN_IN), .A3(P1_DATAWIDTH_REG_13__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_14__SCAN_IN), .ZN(n19871) );
  NOR4_X1 U22830 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_7__SCAN_IN), .A3(P1_DATAWIDTH_REG_8__SCAN_IN), .A4(
        P1_DATAWIDTH_REG_10__SCAN_IN), .ZN(n19870) );
  NAND4_X1 U22831 ( .A1(n19873), .A2(n19872), .A3(n19871), .A4(n19870), .ZN(
        n19874) );
  NOR2_X1 U22832 ( .A1(n19875), .A2(n19874), .ZN(n20783) );
  INV_X1 U22833 ( .A(P1_BYTEENABLE_REG_1__SCAN_IN), .ZN(n19877) );
  NOR3_X1 U22834 ( .A1(P1_REIP_REG_0__SCAN_IN), .A2(
        P1_DATAWIDTH_REG_1__SCAN_IN), .A3(P1_DATAWIDTH_REG_0__SCAN_IN), .ZN(
        n19878) );
  OAI21_X1 U22835 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(n19878), .A(n20783), .ZN(
        n19876) );
  OAI21_X1 U22836 ( .B1(n20783), .B2(n19877), .A(n19876), .ZN(P1_U2807) );
  INV_X1 U22837 ( .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(n20755) );
  AOI21_X1 U22838 ( .B1(n20776), .B2(n20755), .A(n19878), .ZN(n19880) );
  INV_X1 U22839 ( .A(P1_BYTEENABLE_REG_3__SCAN_IN), .ZN(n19879) );
  INV_X1 U22840 ( .A(n20783), .ZN(n20778) );
  AOI22_X1 U22841 ( .A1(n20783), .A2(n19880), .B1(n19879), .B2(n20778), .ZN(
        P1_U2808) );
  AOI22_X1 U22842 ( .A1(n19881), .A2(P1_REIP_REG_9__SCAN_IN), .B1(n19955), 
        .B2(P1_EBX_REG_9__SCAN_IN), .ZN(n19882) );
  OAI21_X1 U22843 ( .B1(n19937), .B2(n19883), .A(n19882), .ZN(n19884) );
  AOI211_X1 U22844 ( .C1(n19932), .C2(P1_PHYADDRPOINTER_REG_9__SCAN_IN), .A(
        n15986), .B(n19884), .ZN(n19889) );
  INV_X1 U22845 ( .A(n19885), .ZN(n19887) );
  AOI22_X1 U22846 ( .A1(n19887), .A2(n19908), .B1(n19941), .B2(n19886), .ZN(
        n19888) );
  OAI211_X1 U22847 ( .C1(P1_REIP_REG_9__SCAN_IN), .C2(n19890), .A(n19889), .B(
        n19888), .ZN(P1_U2831) );
  NOR2_X1 U22848 ( .A1(n19891), .A2(n13858), .ZN(n19893) );
  OAI21_X1 U22849 ( .B1(n19893), .B2(n19892), .A(n19931), .ZN(n19903) );
  AOI22_X1 U22850 ( .A1(n19903), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_EBX_REG_7__SCAN_IN), .B2(n19955), .ZN(n19894) );
  OAI21_X1 U22851 ( .B1(n19937), .B2(n19895), .A(n19894), .ZN(n19896) );
  AOI211_X1 U22852 ( .C1(n19932), .C2(P1_PHYADDRPOINTER_REG_7__SCAN_IN), .A(
        n15986), .B(n19896), .ZN(n19900) );
  AOI22_X1 U22853 ( .A1(n20717), .A2(n19898), .B1(n19897), .B2(n19908), .ZN(
        n19899) );
  OAI211_X1 U22854 ( .C1(n19901), .C2(n19953), .A(n19900), .B(n19899), .ZN(
        P1_U2833) );
  OAI22_X1 U22855 ( .A1(n19937), .A2(n19961), .B1(n19967), .B2(n19934), .ZN(
        n19902) );
  AOI21_X1 U22856 ( .B1(n19903), .B2(P1_REIP_REG_6__SCAN_IN), .A(n19902), .ZN(
        n19904) );
  INV_X1 U22857 ( .A(n19904), .ZN(n19905) );
  AOI211_X1 U22858 ( .C1(n19932), .C2(P1_PHYADDRPOINTER_REG_6__SCAN_IN), .A(
        n15986), .B(n19905), .ZN(n19910) );
  INV_X1 U22859 ( .A(n19906), .ZN(n19907) );
  AOI22_X1 U22860 ( .A1(n19965), .A2(n19908), .B1(n19941), .B2(n19907), .ZN(
        n19909) );
  OAI211_X1 U22861 ( .C1(P1_REIP_REG_6__SCAN_IN), .C2(n19911), .A(n19910), .B(
        n19909), .ZN(P1_U2834) );
  INV_X1 U22862 ( .A(n19931), .ZN(n19913) );
  AOI22_X1 U22863 ( .A1(P1_REIP_REG_5__SCAN_IN), .A2(n19913), .B1(n19912), 
        .B2(n13858), .ZN(n19920) );
  INV_X1 U22864 ( .A(n19960), .ZN(n19943) );
  AOI21_X1 U22865 ( .B1(n19932), .B2(P1_PHYADDRPOINTER_REG_5__SCAN_IN), .A(
        n15986), .ZN(n19915) );
  NAND2_X1 U22866 ( .A1(n19955), .A2(P1_EBX_REG_5__SCAN_IN), .ZN(n19914) );
  OAI211_X1 U22867 ( .C1(n19937), .C2(n19916), .A(n19915), .B(n19914), .ZN(
        n19917) );
  AOI21_X1 U22868 ( .B1(n19918), .B2(n19943), .A(n19917), .ZN(n19919) );
  OAI211_X1 U22869 ( .C1(n19921), .C2(n19953), .A(n19920), .B(n19919), .ZN(
        P1_U2835) );
  AOI22_X1 U22870 ( .A1(n19951), .A2(n20051), .B1(n19922), .B2(n19956), .ZN(
        n19930) );
  INV_X1 U22871 ( .A(P1_REIP_REG_3__SCAN_IN), .ZN(n20712) );
  OR4_X1 U22872 ( .A1(n20712), .A2(n13734), .A3(n19933), .A4(
        P1_REIP_REG_4__SCAN_IN), .ZN(n19923) );
  OAI211_X1 U22873 ( .C1(n19924), .C2(n19934), .A(n19923), .B(n20046), .ZN(
        n19928) );
  OAI22_X1 U22874 ( .A1(n19926), .A2(n19960), .B1(n19925), .B2(n19953), .ZN(
        n19927) );
  AOI211_X1 U22875 ( .C1(P1_PHYADDRPOINTER_REG_4__SCAN_IN), .C2(n19932), .A(
        n19928), .B(n19927), .ZN(n19929) );
  OAI211_X1 U22876 ( .C1(n19931), .C2(n20710), .A(n19930), .B(n19929), .ZN(
        P1_U2836) );
  AOI22_X1 U22877 ( .A1(n19956), .A2(n20771), .B1(n19932), .B2(
        P1_PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n19950) );
  NOR2_X1 U22878 ( .A1(n19933), .A2(P1_REIP_REG_3__SCAN_IN), .ZN(n19939) );
  OAI22_X1 U22879 ( .A1(n19937), .A2(n19936), .B1(n19935), .B2(n19934), .ZN(
        n19938) );
  AOI21_X1 U22880 ( .B1(n19939), .B2(P1_REIP_REG_2__SCAN_IN), .A(n19938), .ZN(
        n19949) );
  INV_X1 U22881 ( .A(n19940), .ZN(n19942) );
  AOI22_X1 U22882 ( .A1(n19944), .A2(n19943), .B1(n19942), .B2(n19941), .ZN(
        n19948) );
  OAI21_X1 U22883 ( .B1(n19946), .B2(n19945), .A(P1_REIP_REG_3__SCAN_IN), .ZN(
        n19947) );
  NAND4_X1 U22884 ( .A1(n19950), .A2(n19949), .A3(n19948), .A4(n19947), .ZN(
        P1_U2837) );
  AOI22_X1 U22885 ( .A1(n19952), .A2(P1_REIP_REG_0__SCAN_IN), .B1(n19951), 
        .B2(n20088), .ZN(n19959) );
  NAND2_X1 U22886 ( .A1(n19954), .A2(n19953), .ZN(n19957) );
  AOI222_X1 U22887 ( .A1(n19957), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n19956), .B2(n20217), .C1(P1_EBX_REG_0__SCAN_IN), .C2(n19955), .ZN(
        n19958) );
  OAI211_X1 U22888 ( .C1(n19960), .C2(n20049), .A(n19959), .B(n19958), .ZN(
        P1_U2840) );
  NOR2_X1 U22889 ( .A1(n19962), .A2(n19961), .ZN(n19963) );
  AOI21_X1 U22890 ( .B1(n19965), .B2(n19964), .A(n19963), .ZN(n19966) );
  OAI21_X1 U22891 ( .B1(n19968), .B2(n19967), .A(n19966), .ZN(P1_U2866) );
  AOI22_X1 U22892 ( .A1(n19993), .A2(P1_LWORD_REG_15__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_15__SCAN_IN), .ZN(n19970) );
  OAI21_X1 U22893 ( .B1(n19971), .B2(n19995), .A(n19970), .ZN(P1_U2921) );
  INV_X1 U22894 ( .A(P1_EAX_REG_14__SCAN_IN), .ZN(n20036) );
  AOI22_X1 U22895 ( .A1(n19993), .A2(P1_LWORD_REG_14__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_14__SCAN_IN), .ZN(n19972) );
  OAI21_X1 U22896 ( .B1(n20036), .B2(n19995), .A(n19972), .ZN(P1_U2922) );
  INV_X1 U22897 ( .A(P1_EAX_REG_13__SCAN_IN), .ZN(n20032) );
  AOI22_X1 U22898 ( .A1(n19993), .A2(P1_LWORD_REG_13__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_13__SCAN_IN), .ZN(n19973) );
  OAI21_X1 U22899 ( .B1(n20032), .B2(n19995), .A(n19973), .ZN(P1_U2923) );
  AOI22_X1 U22900 ( .A1(n19993), .A2(P1_LWORD_REG_12__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_12__SCAN_IN), .ZN(n19974) );
  OAI21_X1 U22901 ( .B1(n14138), .B2(n19995), .A(n19974), .ZN(P1_U2924) );
  AOI22_X1 U22902 ( .A1(n19993), .A2(P1_LWORD_REG_11__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_11__SCAN_IN), .ZN(n19975) );
  OAI21_X1 U22903 ( .B1(n14127), .B2(n19995), .A(n19975), .ZN(P1_U2925) );
  AOI22_X1 U22904 ( .A1(n19993), .A2(P1_LWORD_REG_10__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_10__SCAN_IN), .ZN(n19976) );
  OAI21_X1 U22905 ( .B1(n14064), .B2(n19995), .A(n19976), .ZN(P1_U2926) );
  AOI22_X1 U22906 ( .A1(n19993), .A2(P1_LWORD_REG_9__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_9__SCAN_IN), .ZN(n19977) );
  OAI21_X1 U22907 ( .B1(n13980), .B2(n19995), .A(n19977), .ZN(P1_U2927) );
  AOI22_X1 U22908 ( .A1(n19993), .A2(P1_LWORD_REG_8__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_8__SCAN_IN), .ZN(n19979) );
  OAI21_X1 U22909 ( .B1(n13906), .B2(n19995), .A(n19979), .ZN(P1_U2928) );
  AOI22_X1 U22910 ( .A1(n19993), .A2(P1_LWORD_REG_7__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_7__SCAN_IN), .ZN(n19980) );
  OAI21_X1 U22911 ( .B1(n19981), .B2(n19995), .A(n19980), .ZN(P1_U2929) );
  AOI22_X1 U22912 ( .A1(n19993), .A2(P1_LWORD_REG_6__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_6__SCAN_IN), .ZN(n19982) );
  OAI21_X1 U22913 ( .B1(n12032), .B2(n19995), .A(n19982), .ZN(P1_U2930) );
  INV_X1 U22914 ( .A(P1_EAX_REG_5__SCAN_IN), .ZN(n19984) );
  AOI22_X1 U22915 ( .A1(n19993), .A2(P1_LWORD_REG_5__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_5__SCAN_IN), .ZN(n19983) );
  OAI21_X1 U22916 ( .B1(n19984), .B2(n19995), .A(n19983), .ZN(P1_U2931) );
  AOI22_X1 U22917 ( .A1(n19993), .A2(P1_LWORD_REG_4__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_4__SCAN_IN), .ZN(n19985) );
  OAI21_X1 U22918 ( .B1(n19986), .B2(n19995), .A(n19985), .ZN(P1_U2932) );
  AOI22_X1 U22919 ( .A1(n19993), .A2(P1_LWORD_REG_3__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_3__SCAN_IN), .ZN(n19987) );
  OAI21_X1 U22920 ( .B1(n19988), .B2(n19995), .A(n19987), .ZN(P1_U2933) );
  AOI22_X1 U22921 ( .A1(n19993), .A2(P1_LWORD_REG_2__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_2__SCAN_IN), .ZN(n19989) );
  OAI21_X1 U22922 ( .B1(n19990), .B2(n19995), .A(n19989), .ZN(P1_U2934) );
  AOI22_X1 U22923 ( .A1(n19993), .A2(P1_LWORD_REG_1__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_1__SCAN_IN), .ZN(n19991) );
  OAI21_X1 U22924 ( .B1(n19992), .B2(n19995), .A(n19991), .ZN(P1_U2935) );
  AOI22_X1 U22925 ( .A1(n19993), .A2(P1_LWORD_REG_0__SCAN_IN), .B1(n19978), 
        .B2(P1_DATAO_REG_0__SCAN_IN), .ZN(n19994) );
  OAI21_X1 U22926 ( .B1(n19996), .B2(n19995), .A(n19994), .ZN(P1_U2936) );
  NOR2_X1 U22927 ( .A1(n20016), .A2(n19997), .ZN(n20019) );
  AOI21_X1 U22928 ( .B1(P1_UWORD_REG_8__SCAN_IN), .B2(n20026), .A(n20019), 
        .ZN(n19998) );
  OAI21_X1 U22929 ( .B1(n19999), .B2(n20035), .A(n19998), .ZN(P1_U2945) );
  NOR2_X1 U22930 ( .A1(n20016), .A2(n20000), .ZN(n20021) );
  AOI21_X1 U22931 ( .B1(P1_UWORD_REG_9__SCAN_IN), .B2(n20026), .A(n20021), 
        .ZN(n20001) );
  OAI21_X1 U22932 ( .B1(n20002), .B2(n20035), .A(n20001), .ZN(P1_U2946) );
  NOR2_X1 U22933 ( .A1(n20016), .A2(n20003), .ZN(n20023) );
  AOI21_X1 U22934 ( .B1(P1_UWORD_REG_10__SCAN_IN), .B2(n20026), .A(n20023), 
        .ZN(n20004) );
  OAI21_X1 U22935 ( .B1(n14521), .B2(n20035), .A(n20004), .ZN(P1_U2947) );
  NOR2_X1 U22936 ( .A1(n20016), .A2(n20005), .ZN(n20025) );
  AOI21_X1 U22937 ( .B1(P1_UWORD_REG_11__SCAN_IN), .B2(n20026), .A(n20025), 
        .ZN(n20006) );
  OAI21_X1 U22938 ( .B1(n20007), .B2(n20035), .A(n20006), .ZN(P1_U2948) );
  NOR2_X1 U22939 ( .A1(n20016), .A2(n20008), .ZN(n20028) );
  AOI21_X1 U22940 ( .B1(P1_UWORD_REG_12__SCAN_IN), .B2(n20026), .A(n20028), 
        .ZN(n20009) );
  OAI21_X1 U22941 ( .B1(n14512), .B2(n20035), .A(n20009), .ZN(P1_U2949) );
  INV_X1 U22942 ( .A(n20010), .ZN(n20011) );
  NOR2_X1 U22943 ( .A1(n20016), .A2(n20011), .ZN(n20030) );
  AOI21_X1 U22944 ( .B1(P1_UWORD_REG_13__SCAN_IN), .B2(n20026), .A(n20030), 
        .ZN(n20012) );
  OAI21_X1 U22945 ( .B1(n20013), .B2(n20035), .A(n20012), .ZN(P1_U2950) );
  INV_X1 U22946 ( .A(n20014), .ZN(n20015) );
  NOR2_X1 U22947 ( .A1(n20016), .A2(n20015), .ZN(n20033) );
  AOI21_X1 U22948 ( .B1(P1_UWORD_REG_14__SCAN_IN), .B2(n20026), .A(n20033), 
        .ZN(n20017) );
  OAI21_X1 U22949 ( .B1(n20018), .B2(n20035), .A(n20017), .ZN(P1_U2951) );
  AOI21_X1 U22950 ( .B1(P1_LWORD_REG_8__SCAN_IN), .B2(n20026), .A(n20019), 
        .ZN(n20020) );
  OAI21_X1 U22951 ( .B1(n13906), .B2(n20035), .A(n20020), .ZN(P1_U2960) );
  AOI21_X1 U22952 ( .B1(P1_LWORD_REG_9__SCAN_IN), .B2(n20026), .A(n20021), 
        .ZN(n20022) );
  OAI21_X1 U22953 ( .B1(n13980), .B2(n20035), .A(n20022), .ZN(P1_U2961) );
  AOI21_X1 U22954 ( .B1(P1_LWORD_REG_10__SCAN_IN), .B2(n20026), .A(n20023), 
        .ZN(n20024) );
  OAI21_X1 U22955 ( .B1(n14064), .B2(n20035), .A(n20024), .ZN(P1_U2962) );
  AOI21_X1 U22956 ( .B1(P1_LWORD_REG_11__SCAN_IN), .B2(n20026), .A(n20025), 
        .ZN(n20027) );
  OAI21_X1 U22957 ( .B1(n14127), .B2(n20035), .A(n20027), .ZN(P1_U2963) );
  AOI21_X1 U22958 ( .B1(P1_LWORD_REG_12__SCAN_IN), .B2(n20026), .A(n20028), 
        .ZN(n20029) );
  OAI21_X1 U22959 ( .B1(n14138), .B2(n20035), .A(n20029), .ZN(P1_U2964) );
  AOI21_X1 U22960 ( .B1(P1_LWORD_REG_13__SCAN_IN), .B2(n20026), .A(n20030), 
        .ZN(n20031) );
  OAI21_X1 U22961 ( .B1(n20032), .B2(n20035), .A(n20031), .ZN(P1_U2965) );
  AOI21_X1 U22962 ( .B1(P1_LWORD_REG_14__SCAN_IN), .B2(n20026), .A(n20033), 
        .ZN(n20034) );
  OAI21_X1 U22963 ( .B1(n20036), .B2(n20035), .A(n20034), .ZN(P1_U2966) );
  OR2_X1 U22964 ( .A1(n20038), .A2(n20037), .ZN(n20044) );
  OR2_X1 U22965 ( .A1(n20039), .A2(P1_INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(
        n20040) );
  NAND2_X1 U22966 ( .A1(n20041), .A2(n20040), .ZN(n20094) );
  INV_X1 U22967 ( .A(n20094), .ZN(n20042) );
  AOI22_X1 U22968 ( .A1(n20044), .A2(P1_PHYADDRPOINTER_REG_0__SCAN_IN), .B1(
        n20043), .B2(n20042), .ZN(n20047) );
  INV_X1 U22969 ( .A(P1_REIP_REG_0__SCAN_IN), .ZN(n20045) );
  OR2_X1 U22970 ( .A1(n20046), .A2(n20045), .ZN(n20091) );
  OAI211_X1 U22971 ( .C1(n20049), .C2(n20048), .A(n20047), .B(n20091), .ZN(
        P1_U2999) );
  AOI21_X1 U22972 ( .B1(n20089), .B2(n20051), .A(n20050), .ZN(n20052) );
  OAI21_X1 U22973 ( .B1(n20053), .B2(n11321), .A(n20052), .ZN(n20054) );
  AOI21_X1 U22974 ( .B1(n20055), .B2(n20077), .A(n20054), .ZN(n20059) );
  OAI211_X1 U22975 ( .C1(P1_INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        P1_INSTADDRPOINTER_REG_3__SCAN_IN), .A(n20057), .B(n20056), .ZN(n20058) );
  NAND2_X1 U22976 ( .A1(n20059), .A2(n20058), .ZN(P1_U3027) );
  AOI21_X1 U22977 ( .B1(n20089), .B2(n20061), .A(n20060), .ZN(n20074) );
  NOR2_X1 U22978 ( .A1(n10100), .A2(n20087), .ZN(n20063) );
  OAI221_X1 U22979 ( .B1(n20064), .B2(P1_INSTADDRPOINTER_REG_2__SCAN_IN), .C1(
        n20064), .C2(n20063), .A(n20062), .ZN(n20073) );
  OAI21_X1 U22980 ( .B1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .B2(n20066), .A(
        n20065), .ZN(n20067) );
  AOI22_X1 U22981 ( .A1(n20068), .A2(n20077), .B1(
        P1_INSTADDRPOINTER_REG_2__SCAN_IN), .B2(n20067), .ZN(n20072) );
  NAND3_X1 U22982 ( .A1(P1_INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n20070), .A3(
        n20069), .ZN(n20071) );
  NAND4_X1 U22983 ( .A1(n20074), .A2(n20073), .A3(n20072), .A4(n20071), .ZN(
        P1_U3029) );
  NAND2_X1 U22984 ( .A1(n10100), .A2(n20075), .ZN(n20090) );
  NAND2_X1 U22985 ( .A1(n20087), .A2(n20076), .ZN(n20083) );
  NAND2_X1 U22986 ( .A1(n20078), .A2(n20077), .ZN(n20082) );
  AOI21_X1 U22987 ( .B1(n20089), .B2(n20080), .A(n20079), .ZN(n20081) );
  OAI211_X1 U22988 ( .C1(n20084), .C2(n20083), .A(n20082), .B(n20081), .ZN(
        n20085) );
  INV_X1 U22989 ( .A(n20085), .ZN(n20086) );
  OAI221_X1 U22990 ( .B1(n20087), .B2(n20098), .C1(n20087), .C2(n20090), .A(
        n20086), .ZN(P1_U3030) );
  NAND2_X1 U22991 ( .A1(n20089), .A2(n20088), .ZN(n20093) );
  AND2_X1 U22992 ( .A1(n20091), .A2(n20090), .ZN(n20092) );
  OAI211_X1 U22993 ( .C1(n20095), .C2(n20094), .A(n20093), .B(n20092), .ZN(
        n20096) );
  INV_X1 U22994 ( .A(n20096), .ZN(n20097) );
  OAI221_X1 U22995 ( .B1(n10100), .B2(n20099), .C1(n10100), .C2(n20098), .A(
        n20097), .ZN(P1_U3031) );
  NOR2_X1 U22996 ( .A1(n20100), .A2(n20773), .ZN(P1_U3032) );
  NAND2_X1 U22997 ( .A1(n20101), .A2(n14173), .ZN(n20120) );
  NAND2_X1 U22998 ( .A1(n20102), .A2(n20101), .ZN(n20119) );
  INV_X1 U22999 ( .A(n20766), .ZN(n20103) );
  AOI22_X1 U23000 ( .A1(BUF1_REG_24__SCAN_IN), .A2(n20142), .B1(DATAI_24_), 
        .B2(n20143), .ZN(n20642) );
  INV_X1 U23001 ( .A(n20642), .ZN(n20592) );
  NAND2_X1 U23002 ( .A1(n11501), .A2(n20144), .ZN(n20441) );
  NOR3_X1 U23003 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20157) );
  INV_X1 U23004 ( .A(n20157), .ZN(n20154) );
  NOR2_X1 U23005 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20154), .ZN(
        n20146) );
  AOI22_X1 U23006 ( .A1(n20683), .A2(n20592), .B1(n20632), .B2(n20146), .ZN(
        n20118) );
  INV_X1 U23007 ( .A(n20114), .ZN(n20106) );
  NOR2_X1 U23008 ( .A1(n20106), .A2(n20691), .ZN(n20513) );
  INV_X1 U23009 ( .A(n20683), .ZN(n20107) );
  NAND3_X1 U23010 ( .A1(n20107), .A2(n20169), .A3(n20581), .ZN(n20108) );
  NAND2_X1 U23011 ( .A1(n20581), .A2(n20765), .ZN(n20510) );
  NAND2_X1 U23012 ( .A1(n20108), .A2(n20510), .ZN(n20113) );
  INV_X1 U23013 ( .A(n13655), .ZN(n20109) );
  NAND2_X1 U23014 ( .A1(n9926), .A2(n20380), .ZN(n20115) );
  INV_X1 U23015 ( .A(n20381), .ZN(n20110) );
  NAND2_X1 U23016 ( .A1(n20437), .A2(n20110), .ZN(n20259) );
  AOI22_X1 U23017 ( .A1(n20113), .A2(n20115), .B1(P1_STATE2_REG_2__SCAN_IN), 
        .B2(n20259), .ZN(n20111) );
  OAI211_X1 U23018 ( .C1(n20146), .C2(n20388), .A(n20447), .B(n20111), .ZN(
        n20150) );
  NAND2_X1 U23019 ( .A1(n20112), .A2(n20147), .ZN(n20523) );
  INV_X1 U23020 ( .A(n20113), .ZN(n20116) );
  NOR2_X1 U23021 ( .A1(n20114), .A2(n20691), .ZN(n20438) );
  INV_X1 U23022 ( .A(n20438), .ZN(n20383) );
  AOI22_X1 U23023 ( .A1(P1_INSTQUEUE_REG_0__0__SCAN_IN), .A2(n20150), .B1(
        n20633), .B2(n20149), .ZN(n20117) );
  OAI211_X1 U23024 ( .C1(n20595), .C2(n20169), .A(n20118), .B(n20117), .ZN(
        P1_U3033) );
  INV_X1 U23025 ( .A(DATAI_25_), .ZN(n21054) );
  NAND2_X1 U23026 ( .A1(n20122), .A2(n20144), .ZN(n20450) );
  AOI22_X1 U23027 ( .A1(n20683), .A2(n20596), .B1(n20643), .B2(n20146), .ZN(
        n20125) );
  NAND2_X1 U23028 ( .A1(n20123), .A2(n20147), .ZN(n20526) );
  AOI22_X1 U23029 ( .A1(P1_INSTQUEUE_REG_0__1__SCAN_IN), .A2(n20150), .B1(
        n20644), .B2(n20149), .ZN(n20124) );
  OAI211_X1 U23030 ( .C1(n20599), .C2(n20169), .A(n20125), .B(n20124), .ZN(
        P1_U3034) );
  AOI22_X1 U23031 ( .A1(BUF1_REG_18__SCAN_IN), .A2(n20142), .B1(DATAI_18_), 
        .B2(n20143), .ZN(n20603) );
  AOI22_X1 U23032 ( .A1(BUF1_REG_26__SCAN_IN), .A2(n20142), .B1(DATAI_26_), 
        .B2(n20143), .ZN(n20654) );
  INV_X1 U23033 ( .A(n20654), .ZN(n20600) );
  NAND2_X1 U23034 ( .A1(n11108), .A2(n20144), .ZN(n20454) );
  AOI22_X1 U23035 ( .A1(n20683), .A2(n20600), .B1(n20649), .B2(n20146), .ZN(
        n20128) );
  NAND2_X1 U23036 ( .A1(n20126), .A2(n20147), .ZN(n20529) );
  AOI22_X1 U23037 ( .A1(P1_INSTQUEUE_REG_0__2__SCAN_IN), .A2(n20150), .B1(
        n20650), .B2(n20149), .ZN(n20127) );
  OAI211_X1 U23038 ( .C1(n20603), .C2(n20169), .A(n20128), .B(n20127), .ZN(
        P1_U3035) );
  AOI22_X1 U23039 ( .A1(BUF1_REG_19__SCAN_IN), .A2(n20142), .B1(DATAI_19_), 
        .B2(n20143), .ZN(n20607) );
  AOI22_X1 U23040 ( .A1(BUF1_REG_27__SCAN_IN), .A2(n20142), .B1(DATAI_27_), 
        .B2(n20143), .ZN(n20660) );
  INV_X1 U23041 ( .A(n20660), .ZN(n20604) );
  NAND2_X1 U23042 ( .A1(n20129), .A2(n20144), .ZN(n20458) );
  AOI22_X1 U23043 ( .A1(n20683), .A2(n20604), .B1(n20655), .B2(n20146), .ZN(
        n20132) );
  NAND2_X1 U23044 ( .A1(n20130), .A2(n20147), .ZN(n20532) );
  AOI22_X1 U23045 ( .A1(P1_INSTQUEUE_REG_0__3__SCAN_IN), .A2(n20150), .B1(
        n20656), .B2(n20149), .ZN(n20131) );
  OAI211_X1 U23046 ( .C1(n20607), .C2(n20169), .A(n20132), .B(n20131), .ZN(
        P1_U3036) );
  AOI22_X1 U23047 ( .A1(BUF1_REG_20__SCAN_IN), .A2(n20142), .B1(DATAI_20_), 
        .B2(n20143), .ZN(n20611) );
  AOI22_X1 U23048 ( .A1(BUF1_REG_28__SCAN_IN), .A2(n20142), .B1(DATAI_28_), 
        .B2(n20143), .ZN(n20666) );
  INV_X1 U23049 ( .A(n20666), .ZN(n20608) );
  NAND2_X1 U23050 ( .A1(n11127), .A2(n20144), .ZN(n20462) );
  AOI22_X1 U23051 ( .A1(n20683), .A2(n20608), .B1(n20661), .B2(n20146), .ZN(
        n20135) );
  NAND2_X1 U23052 ( .A1(n20133), .A2(n20147), .ZN(n20535) );
  AOI22_X1 U23053 ( .A1(P1_INSTQUEUE_REG_0__4__SCAN_IN), .A2(n20150), .B1(
        n20662), .B2(n20149), .ZN(n20134) );
  OAI211_X1 U23054 ( .C1(n20611), .C2(n20169), .A(n20135), .B(n20134), .ZN(
        P1_U3037) );
  AOI22_X1 U23055 ( .A1(BUF1_REG_21__SCAN_IN), .A2(n20142), .B1(DATAI_21_), 
        .B2(n20143), .ZN(n20615) );
  AOI22_X1 U23056 ( .A1(BUF1_REG_29__SCAN_IN), .A2(n20142), .B1(DATAI_29_), 
        .B2(n20143), .ZN(n20672) );
  INV_X1 U23057 ( .A(n20672), .ZN(n20612) );
  NAND2_X1 U23058 ( .A1(n11180), .A2(n20144), .ZN(n20333) );
  AOI22_X1 U23059 ( .A1(n20683), .A2(n20612), .B1(n20667), .B2(n20146), .ZN(
        n20138) );
  NAND2_X1 U23060 ( .A1(n20136), .A2(n20147), .ZN(n20538) );
  AOI22_X1 U23061 ( .A1(P1_INSTQUEUE_REG_0__5__SCAN_IN), .A2(n20150), .B1(
        n20668), .B2(n20149), .ZN(n20137) );
  OAI211_X1 U23062 ( .C1(n20615), .C2(n20169), .A(n20138), .B(n20137), .ZN(
        P1_U3038) );
  AOI22_X1 U23063 ( .A1(BUF1_REG_22__SCAN_IN), .A2(n20142), .B1(DATAI_22_), 
        .B2(n20143), .ZN(n20619) );
  AOI22_X1 U23064 ( .A1(BUF1_REG_30__SCAN_IN), .A2(n20142), .B1(DATAI_30_), 
        .B2(n20143), .ZN(n20678) );
  INV_X1 U23065 ( .A(n20678), .ZN(n20616) );
  NAND2_X1 U23066 ( .A1(n11120), .A2(n20144), .ZN(n20337) );
  AOI22_X1 U23067 ( .A1(n20683), .A2(n20616), .B1(n20673), .B2(n20146), .ZN(
        n20141) );
  NAND2_X1 U23068 ( .A1(n20139), .A2(n20147), .ZN(n20541) );
  AOI22_X1 U23069 ( .A1(P1_INSTQUEUE_REG_0__6__SCAN_IN), .A2(n20150), .B1(
        n20674), .B2(n20149), .ZN(n20140) );
  OAI211_X1 U23070 ( .C1(n20619), .C2(n20169), .A(n20141), .B(n20140), .ZN(
        P1_U3039) );
  AOI22_X1 U23071 ( .A1(BUF1_REG_23__SCAN_IN), .A2(n20142), .B1(DATAI_23_), 
        .B2(n20143), .ZN(n20627) );
  AOI22_X1 U23072 ( .A1(DATAI_31_), .A2(n20143), .B1(BUF1_REG_31__SCAN_IN), 
        .B2(n20142), .ZN(n20688) );
  INV_X1 U23073 ( .A(n20688), .ZN(n20622) );
  NAND2_X1 U23074 ( .A1(n20145), .A2(n20144), .ZN(n20472) );
  AOI22_X1 U23075 ( .A1(n20683), .A2(n20622), .B1(n20679), .B2(n20146), .ZN(
        n20152) );
  NAND2_X1 U23076 ( .A1(n20148), .A2(n20147), .ZN(n20547) );
  AOI22_X1 U23077 ( .A1(P1_INSTQUEUE_REG_0__7__SCAN_IN), .A2(n20150), .B1(
        n20680), .B2(n20149), .ZN(n20151) );
  OAI211_X1 U23078 ( .C1(n20627), .C2(n20169), .A(n20152), .B(n20151), .ZN(
        P1_U3040) );
  INV_X1 U23079 ( .A(n20153), .ZN(n20552) );
  NOR2_X1 U23080 ( .A1(n20551), .A2(n20154), .ZN(n20174) );
  AOI21_X1 U23081 ( .B1(n9926), .B2(n20552), .A(n20174), .ZN(n20155) );
  OAI22_X1 U23082 ( .A1(n20155), .A2(n20767), .B1(n20154), .B2(n20691), .ZN(
        n20175) );
  AOI22_X1 U23083 ( .A1(n20175), .A2(n20633), .B1(n20632), .B2(n20174), .ZN(
        n20159) );
  OAI211_X1 U23084 ( .C1(n20221), .C2(n20554), .A(n20581), .B(n20155), .ZN(
        n20156) );
  OAI211_X1 U23085 ( .C1(n20581), .C2(n20157), .A(n20636), .B(n20156), .ZN(
        n20177) );
  AOI22_X1 U23086 ( .A1(P1_INSTQUEUE_REG_1__0__SCAN_IN), .A2(n20177), .B1(
        n20176), .B2(n20592), .ZN(n20158) );
  OAI211_X1 U23087 ( .C1(n20595), .C2(n20209), .A(n20159), .B(n20158), .ZN(
        P1_U3041) );
  AOI22_X1 U23088 ( .A1(n20175), .A2(n20644), .B1(n20643), .B2(n20174), .ZN(
        n20161) );
  AOI22_X1 U23089 ( .A1(P1_INSTQUEUE_REG_1__1__SCAN_IN), .A2(n20177), .B1(
        n20176), .B2(n20596), .ZN(n20160) );
  OAI211_X1 U23090 ( .C1(n20599), .C2(n20209), .A(n20161), .B(n20160), .ZN(
        P1_U3042) );
  AOI22_X1 U23091 ( .A1(n20175), .A2(n20650), .B1(n20649), .B2(n20174), .ZN(
        n20163) );
  AOI22_X1 U23092 ( .A1(P1_INSTQUEUE_REG_1__2__SCAN_IN), .A2(n20177), .B1(
        n20176), .B2(n20600), .ZN(n20162) );
  OAI211_X1 U23093 ( .C1(n20603), .C2(n20209), .A(n20163), .B(n20162), .ZN(
        P1_U3043) );
  AOI22_X1 U23094 ( .A1(n20175), .A2(n20656), .B1(n20655), .B2(n20174), .ZN(
        n20165) );
  AOI22_X1 U23095 ( .A1(P1_INSTQUEUE_REG_1__3__SCAN_IN), .A2(n20177), .B1(
        n20176), .B2(n20604), .ZN(n20164) );
  OAI211_X1 U23096 ( .C1(n20607), .C2(n20209), .A(n20165), .B(n20164), .ZN(
        P1_U3044) );
  AOI22_X1 U23097 ( .A1(n20175), .A2(n20662), .B1(n20661), .B2(n20174), .ZN(
        n20168) );
  INV_X1 U23098 ( .A(n20209), .ZN(n20166) );
  INV_X1 U23099 ( .A(n20611), .ZN(n20663) );
  AOI22_X1 U23100 ( .A1(P1_INSTQUEUE_REG_1__4__SCAN_IN), .A2(n20177), .B1(
        n20166), .B2(n20663), .ZN(n20167) );
  OAI211_X1 U23101 ( .C1(n20666), .C2(n20169), .A(n20168), .B(n20167), .ZN(
        P1_U3045) );
  AOI22_X1 U23102 ( .A1(n20175), .A2(n20668), .B1(n20667), .B2(n20174), .ZN(
        n20171) );
  AOI22_X1 U23103 ( .A1(P1_INSTQUEUE_REG_1__5__SCAN_IN), .A2(n20177), .B1(
        n20176), .B2(n20612), .ZN(n20170) );
  OAI211_X1 U23104 ( .C1(n20615), .C2(n20209), .A(n20171), .B(n20170), .ZN(
        P1_U3046) );
  AOI22_X1 U23105 ( .A1(n20175), .A2(n20674), .B1(n20673), .B2(n20174), .ZN(
        n20173) );
  AOI22_X1 U23106 ( .A1(P1_INSTQUEUE_REG_1__6__SCAN_IN), .A2(n20177), .B1(
        n20176), .B2(n20616), .ZN(n20172) );
  OAI211_X1 U23107 ( .C1(n20619), .C2(n20209), .A(n20173), .B(n20172), .ZN(
        P1_U3047) );
  AOI22_X1 U23108 ( .A1(n20175), .A2(n20680), .B1(n20679), .B2(n20174), .ZN(
        n20179) );
  AOI22_X1 U23109 ( .A1(P1_INSTQUEUE_REG_1__7__SCAN_IN), .A2(n20177), .B1(
        n20176), .B2(n20622), .ZN(n20178) );
  OAI211_X1 U23110 ( .C1(n20627), .C2(n20209), .A(n20179), .B(n20178), .ZN(
        P1_U3048) );
  NAND2_X1 U23111 ( .A1(n13700), .A2(n9828), .ZN(n20434) );
  NOR3_X1 U23112 ( .A1(n20440), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20215) );
  NAND2_X1 U23113 ( .A1(n20551), .A2(n20215), .ZN(n20208) );
  OAI22_X1 U23114 ( .A1(n20209), .A2(n20642), .B1(n20441), .B2(n20208), .ZN(
        n20180) );
  INV_X1 U23115 ( .A(n20180), .ZN(n20189) );
  NAND2_X1 U23116 ( .A1(n20250), .A2(n20209), .ZN(n20181) );
  AOI21_X1 U23117 ( .B1(n20181), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20767), 
        .ZN(n20183) );
  NAND2_X1 U23118 ( .A1(n9926), .A2(n20586), .ZN(n20186) );
  AOI22_X1 U23119 ( .A1(n20183), .A2(n20186), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20208), .ZN(n20182) );
  OAI21_X1 U23120 ( .B1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B2(n20437), .A(
        P1_STATE2_REG_2__SCAN_IN), .ZN(n20313) );
  NAND3_X1 U23121 ( .A1(n20447), .A2(n20182), .A3(n20313), .ZN(n20212) );
  INV_X1 U23122 ( .A(n20183), .ZN(n20187) );
  INV_X1 U23123 ( .A(n20437), .ZN(n20185) );
  INV_X1 U23124 ( .A(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n20184) );
  NAND2_X1 U23125 ( .A1(n20185), .A2(n20184), .ZN(n20316) );
  AOI22_X1 U23126 ( .A1(P1_INSTQUEUE_REG_2__0__SCAN_IN), .A2(n20212), .B1(
        n20633), .B2(n20211), .ZN(n20188) );
  OAI211_X1 U23127 ( .C1(n20595), .C2(n20250), .A(n20189), .B(n20188), .ZN(
        P1_U3049) );
  INV_X1 U23128 ( .A(n20596), .ZN(n20648) );
  OAI22_X1 U23129 ( .A1(n20250), .A2(n20599), .B1(n20450), .B2(n20208), .ZN(
        n20190) );
  INV_X1 U23130 ( .A(n20190), .ZN(n20192) );
  AOI22_X1 U23131 ( .A1(P1_INSTQUEUE_REG_2__1__SCAN_IN), .A2(n20212), .B1(
        n20644), .B2(n20211), .ZN(n20191) );
  OAI211_X1 U23132 ( .C1(n20648), .C2(n20209), .A(n20192), .B(n20191), .ZN(
        P1_U3050) );
  OAI22_X1 U23133 ( .A1(n20250), .A2(n20603), .B1(n20454), .B2(n20208), .ZN(
        n20193) );
  INV_X1 U23134 ( .A(n20193), .ZN(n20195) );
  AOI22_X1 U23135 ( .A1(P1_INSTQUEUE_REG_2__2__SCAN_IN), .A2(n20212), .B1(
        n20650), .B2(n20211), .ZN(n20194) );
  OAI211_X1 U23136 ( .C1(n20654), .C2(n20209), .A(n20195), .B(n20194), .ZN(
        P1_U3051) );
  OAI22_X1 U23137 ( .A1(n20209), .A2(n20660), .B1(n20458), .B2(n20208), .ZN(
        n20196) );
  INV_X1 U23138 ( .A(n20196), .ZN(n20198) );
  AOI22_X1 U23139 ( .A1(P1_INSTQUEUE_REG_2__3__SCAN_IN), .A2(n20212), .B1(
        n20656), .B2(n20211), .ZN(n20197) );
  OAI211_X1 U23140 ( .C1(n20607), .C2(n20250), .A(n20198), .B(n20197), .ZN(
        P1_U3052) );
  OAI22_X1 U23141 ( .A1(n20209), .A2(n20666), .B1(n20462), .B2(n20208), .ZN(
        n20199) );
  INV_X1 U23142 ( .A(n20199), .ZN(n20201) );
  AOI22_X1 U23143 ( .A1(P1_INSTQUEUE_REG_2__4__SCAN_IN), .A2(n20212), .B1(
        n20662), .B2(n20211), .ZN(n20200) );
  OAI211_X1 U23144 ( .C1(n20611), .C2(n20250), .A(n20201), .B(n20200), .ZN(
        P1_U3053) );
  OAI22_X1 U23145 ( .A1(n20209), .A2(n20672), .B1(n20333), .B2(n20208), .ZN(
        n20202) );
  INV_X1 U23146 ( .A(n20202), .ZN(n20204) );
  AOI22_X1 U23147 ( .A1(P1_INSTQUEUE_REG_2__5__SCAN_IN), .A2(n20212), .B1(
        n20668), .B2(n20211), .ZN(n20203) );
  OAI211_X1 U23148 ( .C1(n20615), .C2(n20250), .A(n20204), .B(n20203), .ZN(
        P1_U3054) );
  OAI22_X1 U23149 ( .A1(n20250), .A2(n20619), .B1(n20337), .B2(n20208), .ZN(
        n20205) );
  INV_X1 U23150 ( .A(n20205), .ZN(n20207) );
  AOI22_X1 U23151 ( .A1(P1_INSTQUEUE_REG_2__6__SCAN_IN), .A2(n20212), .B1(
        n20674), .B2(n20211), .ZN(n20206) );
  OAI211_X1 U23152 ( .C1(n20678), .C2(n20209), .A(n20207), .B(n20206), .ZN(
        P1_U3055) );
  OAI22_X1 U23153 ( .A1(n20209), .A2(n20688), .B1(n20472), .B2(n20208), .ZN(
        n20210) );
  INV_X1 U23154 ( .A(n20210), .ZN(n20214) );
  AOI22_X1 U23155 ( .A1(P1_INSTQUEUE_REG_2__7__SCAN_IN), .A2(n20212), .B1(
        n20680), .B2(n20211), .ZN(n20213) );
  OAI211_X1 U23156 ( .C1(n20627), .C2(n20250), .A(n20214), .B(n20213), .ZN(
        P1_U3056) );
  INV_X1 U23157 ( .A(n20215), .ZN(n20224) );
  OR2_X1 U23158 ( .A1(n20221), .A2(n20634), .ZN(n20216) );
  AND2_X1 U23159 ( .A1(n20216), .A2(n20581), .ZN(n20225) );
  INV_X1 U23160 ( .A(n20225), .ZN(n20219) );
  AND2_X1 U23161 ( .A1(n20218), .A2(n20217), .ZN(n20628) );
  AND2_X1 U23162 ( .A1(n20480), .A2(n20184), .ZN(n20222) );
  AOI21_X1 U23163 ( .B1(n9926), .B2(n20628), .A(n20222), .ZN(n20226) );
  OAI22_X1 U23164 ( .A1(n20691), .A2(n20224), .B1(n20219), .B2(n20226), .ZN(
        n20220) );
  INV_X1 U23165 ( .A(n20222), .ZN(n20249) );
  OAI22_X1 U23166 ( .A1(n20278), .A2(n20595), .B1(n20441), .B2(n20249), .ZN(
        n20223) );
  INV_X1 U23167 ( .A(n20223), .ZN(n20229) );
  AOI22_X1 U23168 ( .A1(n20226), .A2(n20225), .B1(n20767), .B2(n20224), .ZN(
        n20227) );
  NAND2_X1 U23169 ( .A1(n20636), .A2(n20227), .ZN(n20252) );
  INV_X1 U23170 ( .A(n20250), .ZN(n20243) );
  AOI22_X1 U23171 ( .A1(P1_INSTQUEUE_REG_3__0__SCAN_IN), .A2(n20252), .B1(
        n20243), .B2(n20592), .ZN(n20228) );
  OAI211_X1 U23172 ( .C1(n20255), .C2(n20523), .A(n20229), .B(n20228), .ZN(
        P1_U3057) );
  OAI22_X1 U23173 ( .A1(n20278), .A2(n20599), .B1(n20450), .B2(n20249), .ZN(
        n20230) );
  INV_X1 U23174 ( .A(n20230), .ZN(n20232) );
  AOI22_X1 U23175 ( .A1(P1_INSTQUEUE_REG_3__1__SCAN_IN), .A2(n20252), .B1(
        n20243), .B2(n20596), .ZN(n20231) );
  OAI211_X1 U23176 ( .C1(n20255), .C2(n20526), .A(n20232), .B(n20231), .ZN(
        P1_U3058) );
  OAI22_X1 U23177 ( .A1(n20250), .A2(n20654), .B1(n20454), .B2(n20249), .ZN(
        n20233) );
  INV_X1 U23178 ( .A(n20233), .ZN(n20235) );
  INV_X1 U23179 ( .A(n20603), .ZN(n20651) );
  AOI22_X1 U23180 ( .A1(P1_INSTQUEUE_REG_3__2__SCAN_IN), .A2(n20252), .B1(
        n20281), .B2(n20651), .ZN(n20234) );
  OAI211_X1 U23181 ( .C1(n20255), .C2(n20529), .A(n20235), .B(n20234), .ZN(
        P1_U3059) );
  OAI22_X1 U23182 ( .A1(n20250), .A2(n20660), .B1(n20458), .B2(n20249), .ZN(
        n20236) );
  INV_X1 U23183 ( .A(n20236), .ZN(n20238) );
  INV_X1 U23184 ( .A(n20607), .ZN(n20657) );
  AOI22_X1 U23185 ( .A1(P1_INSTQUEUE_REG_3__3__SCAN_IN), .A2(n20252), .B1(
        n20281), .B2(n20657), .ZN(n20237) );
  OAI211_X1 U23186 ( .C1(n20255), .C2(n20532), .A(n20238), .B(n20237), .ZN(
        P1_U3060) );
  OAI22_X1 U23187 ( .A1(n20250), .A2(n20666), .B1(n20462), .B2(n20249), .ZN(
        n20239) );
  INV_X1 U23188 ( .A(n20239), .ZN(n20241) );
  AOI22_X1 U23189 ( .A1(P1_INSTQUEUE_REG_3__4__SCAN_IN), .A2(n20252), .B1(
        n20281), .B2(n20663), .ZN(n20240) );
  OAI211_X1 U23190 ( .C1(n20255), .C2(n20535), .A(n20241), .B(n20240), .ZN(
        P1_U3061) );
  OAI22_X1 U23191 ( .A1(n20278), .A2(n20615), .B1(n20333), .B2(n20249), .ZN(
        n20242) );
  INV_X1 U23192 ( .A(n20242), .ZN(n20245) );
  AOI22_X1 U23193 ( .A1(P1_INSTQUEUE_REG_3__5__SCAN_IN), .A2(n20252), .B1(
        n20243), .B2(n20612), .ZN(n20244) );
  OAI211_X1 U23194 ( .C1(n20255), .C2(n20538), .A(n20245), .B(n20244), .ZN(
        P1_U3062) );
  OAI22_X1 U23195 ( .A1(n20250), .A2(n20678), .B1(n20337), .B2(n20249), .ZN(
        n20246) );
  INV_X1 U23196 ( .A(n20246), .ZN(n20248) );
  INV_X1 U23197 ( .A(n20619), .ZN(n20675) );
  AOI22_X1 U23198 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(n20252), .B1(
        n20281), .B2(n20675), .ZN(n20247) );
  OAI211_X1 U23199 ( .C1(n20255), .C2(n20541), .A(n20248), .B(n20247), .ZN(
        P1_U3063) );
  OAI22_X1 U23200 ( .A1(n20250), .A2(n20688), .B1(n20472), .B2(n20249), .ZN(
        n20251) );
  INV_X1 U23201 ( .A(n20251), .ZN(n20254) );
  INV_X1 U23202 ( .A(n20627), .ZN(n20682) );
  AOI22_X1 U23203 ( .A1(P1_INSTQUEUE_REG_3__7__SCAN_IN), .A2(n20252), .B1(
        n20281), .B2(n20682), .ZN(n20253) );
  OAI211_X1 U23204 ( .C1(n20255), .C2(n20547), .A(n20254), .B(n20253), .ZN(
        P1_U3064) );
  INV_X1 U23205 ( .A(n20378), .ZN(n20256) );
  INV_X1 U23206 ( .A(n20513), .ZN(n20584) );
  NOR2_X1 U23207 ( .A1(n13655), .A2(n20257), .ZN(n20349) );
  NAND3_X1 U23208 ( .A1(n20349), .A2(n20581), .A3(n20380), .ZN(n20258) );
  OAI21_X1 U23209 ( .B1(n20259), .B2(n20584), .A(n20258), .ZN(n20280) );
  NOR3_X1 U23210 ( .A1(n20514), .A2(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20288) );
  INV_X1 U23211 ( .A(n20288), .ZN(n20285) );
  NOR2_X1 U23212 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20285), .ZN(
        n20279) );
  AOI22_X1 U23213 ( .A1(n20280), .A2(n20633), .B1(n20632), .B2(n20279), .ZN(
        n20265) );
  INV_X1 U23214 ( .A(n20349), .ZN(n20261) );
  OAI21_X1 U23215 ( .B1(n20281), .B2(n20307), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20260) );
  OAI21_X1 U23216 ( .B1(n20586), .B2(n20261), .A(n20260), .ZN(n20263) );
  AOI22_X1 U23217 ( .A1(P1_INSTQUEUE_REG_4__0__SCAN_IN), .A2(n20282), .B1(
        n20281), .B2(n20592), .ZN(n20264) );
  OAI211_X1 U23218 ( .C1(n20595), .C2(n20304), .A(n20265), .B(n20264), .ZN(
        P1_U3065) );
  AOI22_X1 U23219 ( .A1(n20280), .A2(n20644), .B1(n20643), .B2(n20279), .ZN(
        n20267) );
  INV_X1 U23220 ( .A(n20599), .ZN(n20645) );
  AOI22_X1 U23221 ( .A1(P1_INSTQUEUE_REG_4__1__SCAN_IN), .A2(n20282), .B1(
        n20307), .B2(n20645), .ZN(n20266) );
  OAI211_X1 U23222 ( .C1(n20648), .C2(n20278), .A(n20267), .B(n20266), .ZN(
        P1_U3066) );
  AOI22_X1 U23223 ( .A1(n20280), .A2(n20650), .B1(n20649), .B2(n20279), .ZN(
        n20269) );
  AOI22_X1 U23224 ( .A1(P1_INSTQUEUE_REG_4__2__SCAN_IN), .A2(n20282), .B1(
        n20307), .B2(n20651), .ZN(n20268) );
  OAI211_X1 U23225 ( .C1(n20654), .C2(n20278), .A(n20269), .B(n20268), .ZN(
        P1_U3067) );
  AOI22_X1 U23226 ( .A1(n20280), .A2(n20656), .B1(n20655), .B2(n20279), .ZN(
        n20271) );
  AOI22_X1 U23227 ( .A1(P1_INSTQUEUE_REG_4__3__SCAN_IN), .A2(n20282), .B1(
        n20281), .B2(n20604), .ZN(n20270) );
  OAI211_X1 U23228 ( .C1(n20607), .C2(n20304), .A(n20271), .B(n20270), .ZN(
        P1_U3068) );
  AOI22_X1 U23229 ( .A1(n20280), .A2(n20662), .B1(n20661), .B2(n20279), .ZN(
        n20273) );
  AOI22_X1 U23230 ( .A1(P1_INSTQUEUE_REG_4__4__SCAN_IN), .A2(n20282), .B1(
        n20281), .B2(n20608), .ZN(n20272) );
  OAI211_X1 U23231 ( .C1(n20611), .C2(n20304), .A(n20273), .B(n20272), .ZN(
        P1_U3069) );
  AOI22_X1 U23232 ( .A1(n20280), .A2(n20668), .B1(n20667), .B2(n20279), .ZN(
        n20275) );
  AOI22_X1 U23233 ( .A1(P1_INSTQUEUE_REG_4__5__SCAN_IN), .A2(n20282), .B1(
        n20281), .B2(n20612), .ZN(n20274) );
  OAI211_X1 U23234 ( .C1(n20615), .C2(n20304), .A(n20275), .B(n20274), .ZN(
        P1_U3070) );
  AOI22_X1 U23235 ( .A1(n20280), .A2(n20674), .B1(n20673), .B2(n20279), .ZN(
        n20277) );
  AOI22_X1 U23236 ( .A1(P1_INSTQUEUE_REG_4__6__SCAN_IN), .A2(n20282), .B1(
        n20307), .B2(n20675), .ZN(n20276) );
  OAI211_X1 U23237 ( .C1(n20678), .C2(n20278), .A(n20277), .B(n20276), .ZN(
        P1_U3071) );
  AOI22_X1 U23238 ( .A1(n20280), .A2(n20680), .B1(n20679), .B2(n20279), .ZN(
        n20284) );
  AOI22_X1 U23239 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(n20282), .B1(
        n20281), .B2(n20622), .ZN(n20283) );
  OAI211_X1 U23240 ( .C1(n20627), .C2(n20304), .A(n20284), .B(n20283), .ZN(
        P1_U3072) );
  NOR2_X1 U23241 ( .A1(n20551), .A2(n20285), .ZN(n20305) );
  AOI21_X1 U23242 ( .B1(n20349), .B2(n20552), .A(n20305), .ZN(n20286) );
  OAI22_X1 U23243 ( .A1(n20286), .A2(n20767), .B1(n20285), .B2(n20691), .ZN(
        n20306) );
  AOI22_X1 U23244 ( .A1(n20306), .A2(n20633), .B1(n20632), .B2(n20305), .ZN(
        n20290) );
  OAI21_X1 U23245 ( .B1(n20351), .B2(n20554), .A(n20286), .ZN(n20287) );
  OAI221_X1 U23246 ( .B1(n20581), .B2(n20288), .C1(n20767), .C2(n20287), .A(
        n20636), .ZN(n20308) );
  AOI22_X1 U23247 ( .A1(P1_INSTQUEUE_REG_5__0__SCAN_IN), .A2(n20308), .B1(
        n20307), .B2(n20592), .ZN(n20289) );
  OAI211_X1 U23248 ( .C1(n20595), .C2(n20342), .A(n20290), .B(n20289), .ZN(
        P1_U3073) );
  AOI22_X1 U23249 ( .A1(n20306), .A2(n20644), .B1(n20643), .B2(n20305), .ZN(
        n20292) );
  AOI22_X1 U23250 ( .A1(P1_INSTQUEUE_REG_5__1__SCAN_IN), .A2(n20308), .B1(
        n20307), .B2(n20596), .ZN(n20291) );
  OAI211_X1 U23251 ( .C1(n20599), .C2(n20342), .A(n20292), .B(n20291), .ZN(
        P1_U3074) );
  AOI22_X1 U23252 ( .A1(n20306), .A2(n20650), .B1(n20649), .B2(n20305), .ZN(
        n20294) );
  AOI22_X1 U23253 ( .A1(P1_INSTQUEUE_REG_5__2__SCAN_IN), .A2(n20308), .B1(
        n20307), .B2(n20600), .ZN(n20293) );
  OAI211_X1 U23254 ( .C1(n20603), .C2(n20342), .A(n20294), .B(n20293), .ZN(
        P1_U3075) );
  AOI22_X1 U23255 ( .A1(n20306), .A2(n20656), .B1(n20655), .B2(n20305), .ZN(
        n20296) );
  INV_X1 U23256 ( .A(n20342), .ZN(n20301) );
  AOI22_X1 U23257 ( .A1(P1_INSTQUEUE_REG_5__3__SCAN_IN), .A2(n20308), .B1(
        n20301), .B2(n20657), .ZN(n20295) );
  OAI211_X1 U23258 ( .C1(n20660), .C2(n20304), .A(n20296), .B(n20295), .ZN(
        P1_U3076) );
  AOI22_X1 U23259 ( .A1(n20306), .A2(n20662), .B1(n20661), .B2(n20305), .ZN(
        n20298) );
  AOI22_X1 U23260 ( .A1(P1_INSTQUEUE_REG_5__4__SCAN_IN), .A2(n20308), .B1(
        n20301), .B2(n20663), .ZN(n20297) );
  OAI211_X1 U23261 ( .C1(n20666), .C2(n20304), .A(n20298), .B(n20297), .ZN(
        P1_U3077) );
  AOI22_X1 U23262 ( .A1(n20306), .A2(n20668), .B1(n20667), .B2(n20305), .ZN(
        n20300) );
  AOI22_X1 U23263 ( .A1(P1_INSTQUEUE_REG_5__5__SCAN_IN), .A2(n20308), .B1(
        n20307), .B2(n20612), .ZN(n20299) );
  OAI211_X1 U23264 ( .C1(n20615), .C2(n20342), .A(n20300), .B(n20299), .ZN(
        P1_U3078) );
  AOI22_X1 U23265 ( .A1(n20306), .A2(n20674), .B1(n20673), .B2(n20305), .ZN(
        n20303) );
  AOI22_X1 U23266 ( .A1(P1_INSTQUEUE_REG_5__6__SCAN_IN), .A2(n20308), .B1(
        n20301), .B2(n20675), .ZN(n20302) );
  OAI211_X1 U23267 ( .C1(n20678), .C2(n20304), .A(n20303), .B(n20302), .ZN(
        P1_U3079) );
  AOI22_X1 U23268 ( .A1(n20306), .A2(n20680), .B1(n20679), .B2(n20305), .ZN(
        n20310) );
  AOI22_X1 U23269 ( .A1(P1_INSTQUEUE_REG_5__7__SCAN_IN), .A2(n20308), .B1(
        n20307), .B2(n20622), .ZN(n20309) );
  OAI211_X1 U23270 ( .C1(n20627), .C2(n20342), .A(n20310), .B(n20309), .ZN(
        P1_U3080) );
  INV_X1 U23271 ( .A(n20350), .ZN(n20355) );
  NAND2_X1 U23272 ( .A1(n20551), .A2(n20355), .ZN(n20341) );
  OAI22_X1 U23273 ( .A1(n20342), .A2(n20642), .B1(n20441), .B2(n20341), .ZN(
        n20311) );
  INV_X1 U23274 ( .A(n20311), .ZN(n20320) );
  NAND2_X1 U23275 ( .A1(n20377), .A2(n20342), .ZN(n20312) );
  AOI21_X1 U23276 ( .B1(n20312), .B2(P1_STATEBS16_REG_SCAN_IN), .A(n20767), 
        .ZN(n20315) );
  NAND2_X1 U23277 ( .A1(n20349), .A2(n20586), .ZN(n20317) );
  AOI22_X1 U23278 ( .A1(n20315), .A2(n20317), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20341), .ZN(n20314) );
  NAND3_X1 U23279 ( .A1(n20589), .A2(n20314), .A3(n20313), .ZN(n20345) );
  INV_X1 U23280 ( .A(n20315), .ZN(n20318) );
  AOI22_X1 U23281 ( .A1(P1_INSTQUEUE_REG_6__0__SCAN_IN), .A2(n20345), .B1(
        n20633), .B2(n20344), .ZN(n20319) );
  OAI211_X1 U23282 ( .C1(n20595), .C2(n20377), .A(n20320), .B(n20319), .ZN(
        P1_U3081) );
  OAI22_X1 U23283 ( .A1(n20377), .A2(n20599), .B1(n20341), .B2(n20450), .ZN(
        n20321) );
  INV_X1 U23284 ( .A(n20321), .ZN(n20323) );
  AOI22_X1 U23285 ( .A1(P1_INSTQUEUE_REG_6__1__SCAN_IN), .A2(n20345), .B1(
        n20644), .B2(n20344), .ZN(n20322) );
  OAI211_X1 U23286 ( .C1(n20648), .C2(n20342), .A(n20323), .B(n20322), .ZN(
        P1_U3082) );
  OAI22_X1 U23287 ( .A1(n20377), .A2(n20603), .B1(n20341), .B2(n20454), .ZN(
        n20324) );
  INV_X1 U23288 ( .A(n20324), .ZN(n20326) );
  AOI22_X1 U23289 ( .A1(P1_INSTQUEUE_REG_6__2__SCAN_IN), .A2(n20345), .B1(
        n20650), .B2(n20344), .ZN(n20325) );
  OAI211_X1 U23290 ( .C1(n20654), .C2(n20342), .A(n20326), .B(n20325), .ZN(
        P1_U3083) );
  OAI22_X1 U23291 ( .A1(n20342), .A2(n20660), .B1(n20458), .B2(n20341), .ZN(
        n20327) );
  INV_X1 U23292 ( .A(n20327), .ZN(n20329) );
  AOI22_X1 U23293 ( .A1(P1_INSTQUEUE_REG_6__3__SCAN_IN), .A2(n20345), .B1(
        n20656), .B2(n20344), .ZN(n20328) );
  OAI211_X1 U23294 ( .C1(n20607), .C2(n20377), .A(n20329), .B(n20328), .ZN(
        P1_U3084) );
  OAI22_X1 U23295 ( .A1(n20377), .A2(n20611), .B1(n20341), .B2(n20462), .ZN(
        n20330) );
  INV_X1 U23296 ( .A(n20330), .ZN(n20332) );
  AOI22_X1 U23297 ( .A1(P1_INSTQUEUE_REG_6__4__SCAN_IN), .A2(n20345), .B1(
        n20662), .B2(n20344), .ZN(n20331) );
  OAI211_X1 U23298 ( .C1(n20666), .C2(n20342), .A(n20332), .B(n20331), .ZN(
        P1_U3085) );
  OAI22_X1 U23299 ( .A1(n20377), .A2(n20615), .B1(n20333), .B2(n20341), .ZN(
        n20334) );
  INV_X1 U23300 ( .A(n20334), .ZN(n20336) );
  AOI22_X1 U23301 ( .A1(P1_INSTQUEUE_REG_6__5__SCAN_IN), .A2(n20345), .B1(
        n20668), .B2(n20344), .ZN(n20335) );
  OAI211_X1 U23302 ( .C1(n20672), .C2(n20342), .A(n20336), .B(n20335), .ZN(
        P1_U3086) );
  OAI22_X1 U23303 ( .A1(n20342), .A2(n20678), .B1(n20341), .B2(n20337), .ZN(
        n20338) );
  INV_X1 U23304 ( .A(n20338), .ZN(n20340) );
  AOI22_X1 U23305 ( .A1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .A2(n20345), .B1(
        n20674), .B2(n20344), .ZN(n20339) );
  OAI211_X1 U23306 ( .C1(n20619), .C2(n20377), .A(n20340), .B(n20339), .ZN(
        P1_U3087) );
  OAI22_X1 U23307 ( .A1(n20342), .A2(n20688), .B1(n20472), .B2(n20341), .ZN(
        n20343) );
  INV_X1 U23308 ( .A(n20343), .ZN(n20347) );
  AOI22_X1 U23309 ( .A1(P1_INSTQUEUE_REG_6__7__SCAN_IN), .A2(n20345), .B1(
        n20680), .B2(n20344), .ZN(n20346) );
  OAI211_X1 U23310 ( .C1(n20627), .C2(n20377), .A(n20347), .B(n20346), .ZN(
        P1_U3088) );
  AOI21_X1 U23311 ( .B1(n20349), .B2(n20628), .A(n20372), .ZN(n20352) );
  OAI22_X1 U23312 ( .A1(n20352), .A2(n20767), .B1(n20350), .B2(n20691), .ZN(
        n20373) );
  AOI22_X1 U23313 ( .A1(n20373), .A2(n20633), .B1(n20632), .B2(n20372), .ZN(
        n20357) );
  NOR2_X1 U23314 ( .A1(n20351), .A2(n20634), .ZN(n20764) );
  INV_X1 U23315 ( .A(n20764), .ZN(n20353) );
  NAND2_X1 U23316 ( .A1(n20353), .A2(n20352), .ZN(n20354) );
  OAI221_X1 U23317 ( .B1(n20581), .B2(n20355), .C1(n20767), .C2(n20354), .A(
        n20636), .ZN(n20374) );
  INV_X1 U23318 ( .A(n20377), .ZN(n20368) );
  AOI22_X1 U23319 ( .A1(P1_INSTQUEUE_REG_7__0__SCAN_IN), .A2(n20374), .B1(
        n20368), .B2(n20592), .ZN(n20356) );
  OAI211_X1 U23320 ( .C1(n20595), .C2(n20371), .A(n20357), .B(n20356), .ZN(
        P1_U3089) );
  AOI22_X1 U23321 ( .A1(n20373), .A2(n20644), .B1(n20643), .B2(n20372), .ZN(
        n20359) );
  AOI22_X1 U23322 ( .A1(P1_INSTQUEUE_REG_7__1__SCAN_IN), .A2(n20374), .B1(
        n20368), .B2(n20596), .ZN(n20358) );
  OAI211_X1 U23323 ( .C1(n20599), .C2(n20371), .A(n20359), .B(n20358), .ZN(
        P1_U3090) );
  AOI22_X1 U23324 ( .A1(n20373), .A2(n20650), .B1(n20649), .B2(n20372), .ZN(
        n20361) );
  AOI22_X1 U23325 ( .A1(P1_INSTQUEUE_REG_7__2__SCAN_IN), .A2(n20374), .B1(
        n20368), .B2(n20600), .ZN(n20360) );
  OAI211_X1 U23326 ( .C1(n20603), .C2(n20371), .A(n20361), .B(n20360), .ZN(
        P1_U3091) );
  AOI22_X1 U23327 ( .A1(n20373), .A2(n20656), .B1(n20655), .B2(n20372), .ZN(
        n20363) );
  AOI22_X1 U23328 ( .A1(P1_INSTQUEUE_REG_7__3__SCAN_IN), .A2(n20374), .B1(
        n20405), .B2(n20657), .ZN(n20362) );
  OAI211_X1 U23329 ( .C1(n20660), .C2(n20377), .A(n20363), .B(n20362), .ZN(
        P1_U3092) );
  AOI22_X1 U23330 ( .A1(n20373), .A2(n20662), .B1(n20661), .B2(n20372), .ZN(
        n20365) );
  AOI22_X1 U23331 ( .A1(P1_INSTQUEUE_REG_7__4__SCAN_IN), .A2(n20374), .B1(
        n20368), .B2(n20608), .ZN(n20364) );
  OAI211_X1 U23332 ( .C1(n20611), .C2(n20371), .A(n20365), .B(n20364), .ZN(
        P1_U3093) );
  AOI22_X1 U23333 ( .A1(n20373), .A2(n20668), .B1(n20667), .B2(n20372), .ZN(
        n20367) );
  INV_X1 U23334 ( .A(n20615), .ZN(n20669) );
  AOI22_X1 U23335 ( .A1(P1_INSTQUEUE_REG_7__5__SCAN_IN), .A2(n20374), .B1(
        n20405), .B2(n20669), .ZN(n20366) );
  OAI211_X1 U23336 ( .C1(n20672), .C2(n20377), .A(n20367), .B(n20366), .ZN(
        P1_U3094) );
  AOI22_X1 U23337 ( .A1(n20373), .A2(n20674), .B1(n20673), .B2(n20372), .ZN(
        n20370) );
  AOI22_X1 U23338 ( .A1(P1_INSTQUEUE_REG_7__6__SCAN_IN), .A2(n20374), .B1(
        n20368), .B2(n20616), .ZN(n20369) );
  OAI211_X1 U23339 ( .C1(n20619), .C2(n20371), .A(n20370), .B(n20369), .ZN(
        P1_U3095) );
  AOI22_X1 U23340 ( .A1(n20373), .A2(n20680), .B1(n20679), .B2(n20372), .ZN(
        n20376) );
  AOI22_X1 U23341 ( .A1(P1_INSTQUEUE_REG_7__7__SCAN_IN), .A2(n20374), .B1(
        n20405), .B2(n20682), .ZN(n20375) );
  OAI211_X1 U23342 ( .C1(n20688), .C2(n20377), .A(n20376), .B(n20375), .ZN(
        P1_U3096) );
  AND2_X1 U23343 ( .A1(n13655), .A2(n20771), .ZN(n20481) );
  NOR3_X1 U23344 ( .A1(n20184), .A2(P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20412) );
  INV_X1 U23345 ( .A(n20412), .ZN(n20409) );
  NOR2_X1 U23346 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20409), .ZN(
        n20403) );
  AOI21_X1 U23347 ( .B1(n20481), .B2(n20380), .A(n20403), .ZN(n20385) );
  AND2_X1 U23348 ( .A1(n20381), .A2(n20437), .ZN(n20520) );
  INV_X1 U23349 ( .A(n20520), .ZN(n20382) );
  OAI22_X1 U23350 ( .A1(n20385), .A2(n20767), .B1(n20383), .B2(n20382), .ZN(
        n20404) );
  AOI22_X1 U23351 ( .A1(n20404), .A2(n20633), .B1(n20632), .B2(n20403), .ZN(
        n20390) );
  INV_X1 U23352 ( .A(n20433), .ZN(n20384) );
  OAI21_X1 U23353 ( .B1(n20384), .B2(n20405), .A(P1_STATEBS16_REG_SCAN_IN), 
        .ZN(n20386) );
  NAND2_X1 U23354 ( .A1(n20386), .A2(n20385), .ZN(n20387) );
  AOI22_X1 U23355 ( .A1(P1_INSTQUEUE_REG_8__0__SCAN_IN), .A2(n20406), .B1(
        n20405), .B2(n20592), .ZN(n20389) );
  OAI211_X1 U23356 ( .C1(n20595), .C2(n20433), .A(n20390), .B(n20389), .ZN(
        P1_U3097) );
  AOI22_X1 U23357 ( .A1(n20404), .A2(n20644), .B1(n20643), .B2(n20403), .ZN(
        n20392) );
  AOI22_X1 U23358 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(n20406), .B1(
        n20405), .B2(n20596), .ZN(n20391) );
  OAI211_X1 U23359 ( .C1(n20599), .C2(n20433), .A(n20392), .B(n20391), .ZN(
        P1_U3098) );
  AOI22_X1 U23360 ( .A1(n20404), .A2(n20650), .B1(n20649), .B2(n20403), .ZN(
        n20394) );
  AOI22_X1 U23361 ( .A1(P1_INSTQUEUE_REG_8__2__SCAN_IN), .A2(n20406), .B1(
        n20405), .B2(n20600), .ZN(n20393) );
  OAI211_X1 U23362 ( .C1(n20603), .C2(n20433), .A(n20394), .B(n20393), .ZN(
        P1_U3099) );
  AOI22_X1 U23363 ( .A1(n20404), .A2(n20656), .B1(n20655), .B2(n20403), .ZN(
        n20396) );
  AOI22_X1 U23364 ( .A1(P1_INSTQUEUE_REG_8__3__SCAN_IN), .A2(n20406), .B1(
        n20405), .B2(n20604), .ZN(n20395) );
  OAI211_X1 U23365 ( .C1(n20607), .C2(n20433), .A(n20396), .B(n20395), .ZN(
        P1_U3100) );
  AOI22_X1 U23366 ( .A1(n20404), .A2(n20662), .B1(n20661), .B2(n20403), .ZN(
        n20398) );
  AOI22_X1 U23367 ( .A1(P1_INSTQUEUE_REG_8__4__SCAN_IN), .A2(n20406), .B1(
        n20405), .B2(n20608), .ZN(n20397) );
  OAI211_X1 U23368 ( .C1(n20611), .C2(n20433), .A(n20398), .B(n20397), .ZN(
        P1_U3101) );
  AOI22_X1 U23369 ( .A1(n20404), .A2(n20668), .B1(n20667), .B2(n20403), .ZN(
        n20400) );
  AOI22_X1 U23370 ( .A1(P1_INSTQUEUE_REG_8__5__SCAN_IN), .A2(n20406), .B1(
        n20405), .B2(n20612), .ZN(n20399) );
  OAI211_X1 U23371 ( .C1(n20615), .C2(n20433), .A(n20400), .B(n20399), .ZN(
        P1_U3102) );
  AOI22_X1 U23372 ( .A1(n20404), .A2(n20674), .B1(n20673), .B2(n20403), .ZN(
        n20402) );
  AOI22_X1 U23373 ( .A1(P1_INSTQUEUE_REG_8__6__SCAN_IN), .A2(n20406), .B1(
        n20405), .B2(n20616), .ZN(n20401) );
  OAI211_X1 U23374 ( .C1(n20619), .C2(n20433), .A(n20402), .B(n20401), .ZN(
        P1_U3103) );
  AOI22_X1 U23375 ( .A1(n20404), .A2(n20680), .B1(n20679), .B2(n20403), .ZN(
        n20408) );
  AOI22_X1 U23376 ( .A1(P1_INSTQUEUE_REG_8__7__SCAN_IN), .A2(n20406), .B1(
        n20405), .B2(n20622), .ZN(n20407) );
  OAI211_X1 U23377 ( .C1(n20627), .C2(n20433), .A(n20408), .B(n20407), .ZN(
        P1_U3104) );
  NOR2_X1 U23378 ( .A1(n20551), .A2(n20409), .ZN(n20428) );
  AOI21_X1 U23379 ( .B1(n20481), .B2(n20552), .A(n20428), .ZN(n20410) );
  OAI22_X1 U23380 ( .A1(n20410), .A2(n20767), .B1(n20409), .B2(n20691), .ZN(
        n20429) );
  AOI22_X1 U23381 ( .A1(n20429), .A2(n20633), .B1(n20632), .B2(n20428), .ZN(
        n20415) );
  INV_X1 U23382 ( .A(n20487), .ZN(n20768) );
  OAI211_X1 U23383 ( .C1(n20768), .C2(n20554), .A(n20581), .B(n20410), .ZN(
        n20411) );
  OAI211_X1 U23384 ( .C1(n20581), .C2(n20412), .A(n20636), .B(n20411), .ZN(
        n20430) );
  INV_X1 U23385 ( .A(n20595), .ZN(n20639) );
  AOI22_X1 U23386 ( .A1(P1_INSTQUEUE_REG_9__0__SCAN_IN), .A2(n20430), .B1(
        n20475), .B2(n20639), .ZN(n20414) );
  OAI211_X1 U23387 ( .C1(n20642), .C2(n20433), .A(n20415), .B(n20414), .ZN(
        P1_U3105) );
  AOI22_X1 U23388 ( .A1(n20429), .A2(n20644), .B1(n20643), .B2(n20428), .ZN(
        n20417) );
  AOI22_X1 U23389 ( .A1(P1_INSTQUEUE_REG_9__1__SCAN_IN), .A2(n20430), .B1(
        n20475), .B2(n20645), .ZN(n20416) );
  OAI211_X1 U23390 ( .C1(n20648), .C2(n20433), .A(n20417), .B(n20416), .ZN(
        P1_U3106) );
  AOI22_X1 U23391 ( .A1(n20429), .A2(n20650), .B1(n20649), .B2(n20428), .ZN(
        n20419) );
  AOI22_X1 U23392 ( .A1(P1_INSTQUEUE_REG_9__2__SCAN_IN), .A2(n20430), .B1(
        n20475), .B2(n20651), .ZN(n20418) );
  OAI211_X1 U23393 ( .C1(n20654), .C2(n20433), .A(n20419), .B(n20418), .ZN(
        P1_U3107) );
  AOI22_X1 U23394 ( .A1(n20429), .A2(n20656), .B1(n20655), .B2(n20428), .ZN(
        n20421) );
  AOI22_X1 U23395 ( .A1(P1_INSTQUEUE_REG_9__3__SCAN_IN), .A2(n20430), .B1(
        n20475), .B2(n20657), .ZN(n20420) );
  OAI211_X1 U23396 ( .C1(n20660), .C2(n20433), .A(n20421), .B(n20420), .ZN(
        P1_U3108) );
  AOI22_X1 U23397 ( .A1(n20429), .A2(n20662), .B1(n20661), .B2(n20428), .ZN(
        n20423) );
  AOI22_X1 U23398 ( .A1(P1_INSTQUEUE_REG_9__4__SCAN_IN), .A2(n20430), .B1(
        n20475), .B2(n20663), .ZN(n20422) );
  OAI211_X1 U23399 ( .C1(n20666), .C2(n20433), .A(n20423), .B(n20422), .ZN(
        P1_U3109) );
  AOI22_X1 U23400 ( .A1(n20429), .A2(n20668), .B1(n20667), .B2(n20428), .ZN(
        n20425) );
  AOI22_X1 U23401 ( .A1(P1_INSTQUEUE_REG_9__5__SCAN_IN), .A2(n20430), .B1(
        n20475), .B2(n20669), .ZN(n20424) );
  OAI211_X1 U23402 ( .C1(n20672), .C2(n20433), .A(n20425), .B(n20424), .ZN(
        P1_U3110) );
  AOI22_X1 U23403 ( .A1(n20429), .A2(n20674), .B1(n20673), .B2(n20428), .ZN(
        n20427) );
  AOI22_X1 U23404 ( .A1(P1_INSTQUEUE_REG_9__6__SCAN_IN), .A2(n20430), .B1(
        n20475), .B2(n20675), .ZN(n20426) );
  OAI211_X1 U23405 ( .C1(n20678), .C2(n20433), .A(n20427), .B(n20426), .ZN(
        P1_U3111) );
  AOI22_X1 U23406 ( .A1(n20429), .A2(n20680), .B1(n20679), .B2(n20428), .ZN(
        n20432) );
  AOI22_X1 U23407 ( .A1(P1_INSTQUEUE_REG_9__7__SCAN_IN), .A2(n20430), .B1(
        n20475), .B2(n20682), .ZN(n20431) );
  OAI211_X1 U23408 ( .C1(n20688), .C2(n20433), .A(n20432), .B(n20431), .ZN(
        P1_U3112) );
  INV_X1 U23409 ( .A(n20475), .ZN(n20435) );
  NAND3_X1 U23410 ( .A1(n20435), .A2(n20581), .A3(n20507), .ZN(n20436) );
  NAND2_X1 U23411 ( .A1(n20436), .A2(n20510), .ZN(n20445) );
  AND2_X1 U23412 ( .A1(n20481), .A2(n20586), .ZN(n20443) );
  OR2_X1 U23413 ( .A1(n20437), .A2(n20184), .ZN(n20583) );
  INV_X1 U23414 ( .A(n20583), .ZN(n20439) );
  NOR3_X1 U23415 ( .A1(n20184), .A2(n20440), .A3(
        P1_INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n20485) );
  NAND2_X1 U23416 ( .A1(n20551), .A2(n20485), .ZN(n20473) );
  OAI22_X1 U23417 ( .A1(n20507), .A2(n20595), .B1(n20473), .B2(n20441), .ZN(
        n20442) );
  INV_X1 U23418 ( .A(n20442), .ZN(n20449) );
  INV_X1 U23419 ( .A(n20443), .ZN(n20444) );
  AOI22_X1 U23420 ( .A1(n20445), .A2(n20444), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20473), .ZN(n20446) );
  NAND2_X1 U23421 ( .A1(P1_STATE2_REG_2__SCAN_IN), .A2(n20583), .ZN(n20588) );
  NAND3_X1 U23422 ( .A1(n20447), .A2(n20446), .A3(n20588), .ZN(n20476) );
  AOI22_X1 U23423 ( .A1(P1_INSTQUEUE_REG_10__0__SCAN_IN), .A2(n20476), .B1(
        n20475), .B2(n20592), .ZN(n20448) );
  OAI211_X1 U23424 ( .C1(n20479), .C2(n20523), .A(n20449), .B(n20448), .ZN(
        P1_U3113) );
  OAI22_X1 U23425 ( .A1(n20507), .A2(n20599), .B1(n20473), .B2(n20450), .ZN(
        n20451) );
  INV_X1 U23426 ( .A(n20451), .ZN(n20453) );
  AOI22_X1 U23427 ( .A1(P1_INSTQUEUE_REG_10__1__SCAN_IN), .A2(n20476), .B1(
        n20475), .B2(n20596), .ZN(n20452) );
  OAI211_X1 U23428 ( .C1(n20479), .C2(n20526), .A(n20453), .B(n20452), .ZN(
        P1_U3114) );
  OAI22_X1 U23429 ( .A1(n20507), .A2(n20603), .B1(n20473), .B2(n20454), .ZN(
        n20455) );
  INV_X1 U23430 ( .A(n20455), .ZN(n20457) );
  AOI22_X1 U23431 ( .A1(P1_INSTQUEUE_REG_10__2__SCAN_IN), .A2(n20476), .B1(
        n20475), .B2(n20600), .ZN(n20456) );
  OAI211_X1 U23432 ( .C1(n20479), .C2(n20529), .A(n20457), .B(n20456), .ZN(
        P1_U3115) );
  OAI22_X1 U23433 ( .A1(n20507), .A2(n20607), .B1(n20473), .B2(n20458), .ZN(
        n20459) );
  INV_X1 U23434 ( .A(n20459), .ZN(n20461) );
  AOI22_X1 U23435 ( .A1(P1_INSTQUEUE_REG_10__3__SCAN_IN), .A2(n20476), .B1(
        n20475), .B2(n20604), .ZN(n20460) );
  OAI211_X1 U23436 ( .C1(n20479), .C2(n20532), .A(n20461), .B(n20460), .ZN(
        P1_U3116) );
  OAI22_X1 U23437 ( .A1(n20507), .A2(n20611), .B1(n20473), .B2(n20462), .ZN(
        n20463) );
  INV_X1 U23438 ( .A(n20463), .ZN(n20465) );
  AOI22_X1 U23439 ( .A1(P1_INSTQUEUE_REG_10__4__SCAN_IN), .A2(n20476), .B1(
        n20475), .B2(n20608), .ZN(n20464) );
  OAI211_X1 U23440 ( .C1(n20479), .C2(n20535), .A(n20465), .B(n20464), .ZN(
        P1_U3117) );
  INV_X1 U23441 ( .A(n20473), .ZN(n20468) );
  AOI22_X1 U23442 ( .A1(n20475), .A2(n20612), .B1(n20667), .B2(n20468), .ZN(
        n20467) );
  INV_X1 U23443 ( .A(n20507), .ZN(n20469) );
  AOI22_X1 U23444 ( .A1(P1_INSTQUEUE_REG_10__5__SCAN_IN), .A2(n20476), .B1(
        n20469), .B2(n20669), .ZN(n20466) );
  OAI211_X1 U23445 ( .C1(n20479), .C2(n20538), .A(n20467), .B(n20466), .ZN(
        P1_U3118) );
  AOI22_X1 U23446 ( .A1(n20475), .A2(n20616), .B1(n20468), .B2(n20673), .ZN(
        n20471) );
  AOI22_X1 U23447 ( .A1(P1_INSTQUEUE_REG_10__6__SCAN_IN), .A2(n20476), .B1(
        n20469), .B2(n20675), .ZN(n20470) );
  OAI211_X1 U23448 ( .C1(n20479), .C2(n20541), .A(n20471), .B(n20470), .ZN(
        P1_U3119) );
  OAI22_X1 U23449 ( .A1(n20507), .A2(n20627), .B1(n20473), .B2(n20472), .ZN(
        n20474) );
  INV_X1 U23450 ( .A(n20474), .ZN(n20478) );
  AOI22_X1 U23451 ( .A1(P1_INSTQUEUE_REG_10__7__SCAN_IN), .A2(n20476), .B1(
        n20475), .B2(n20622), .ZN(n20477) );
  OAI211_X1 U23452 ( .C1(n20479), .C2(n20547), .A(n20478), .B(n20477), .ZN(
        P1_U3120) );
  AND2_X1 U23453 ( .A1(P1_INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n20480), .ZN(
        n20502) );
  AOI21_X1 U23454 ( .B1(n20481), .B2(n20628), .A(n20502), .ZN(n20483) );
  INV_X1 U23455 ( .A(n20485), .ZN(n20482) );
  OAI22_X1 U23456 ( .A1(n20483), .A2(n20767), .B1(n20482), .B2(n20691), .ZN(
        n20503) );
  AOI22_X1 U23457 ( .A1(n20503), .A2(n20633), .B1(n20632), .B2(n20502), .ZN(
        n20489) );
  OAI211_X1 U23458 ( .C1(n20768), .C2(n20634), .A(n20581), .B(n20483), .ZN(
        n20484) );
  OAI211_X1 U23459 ( .C1(n20581), .C2(n20485), .A(n20636), .B(n20484), .ZN(
        n20504) );
  AOI22_X1 U23460 ( .A1(P1_INSTQUEUE_REG_11__0__SCAN_IN), .A2(n20504), .B1(
        n20543), .B2(n20639), .ZN(n20488) );
  OAI211_X1 U23461 ( .C1(n20642), .C2(n20507), .A(n20489), .B(n20488), .ZN(
        P1_U3121) );
  AOI22_X1 U23462 ( .A1(n20503), .A2(n20644), .B1(n20643), .B2(n20502), .ZN(
        n20491) );
  AOI22_X1 U23463 ( .A1(P1_INSTQUEUE_REG_11__1__SCAN_IN), .A2(n20504), .B1(
        n20543), .B2(n20645), .ZN(n20490) );
  OAI211_X1 U23464 ( .C1(n20648), .C2(n20507), .A(n20491), .B(n20490), .ZN(
        P1_U3122) );
  AOI22_X1 U23465 ( .A1(n20503), .A2(n20650), .B1(n20649), .B2(n20502), .ZN(
        n20493) );
  AOI22_X1 U23466 ( .A1(P1_INSTQUEUE_REG_11__2__SCAN_IN), .A2(n20504), .B1(
        n20543), .B2(n20651), .ZN(n20492) );
  OAI211_X1 U23467 ( .C1(n20654), .C2(n20507), .A(n20493), .B(n20492), .ZN(
        P1_U3123) );
  AOI22_X1 U23468 ( .A1(n20503), .A2(n20656), .B1(n20655), .B2(n20502), .ZN(
        n20495) );
  AOI22_X1 U23469 ( .A1(P1_INSTQUEUE_REG_11__3__SCAN_IN), .A2(n20504), .B1(
        n20543), .B2(n20657), .ZN(n20494) );
  OAI211_X1 U23470 ( .C1(n20660), .C2(n20507), .A(n20495), .B(n20494), .ZN(
        P1_U3124) );
  AOI22_X1 U23471 ( .A1(n20503), .A2(n20662), .B1(n20661), .B2(n20502), .ZN(
        n20497) );
  AOI22_X1 U23472 ( .A1(P1_INSTQUEUE_REG_11__4__SCAN_IN), .A2(n20504), .B1(
        n20543), .B2(n20663), .ZN(n20496) );
  OAI211_X1 U23473 ( .C1(n20666), .C2(n20507), .A(n20497), .B(n20496), .ZN(
        P1_U3125) );
  AOI22_X1 U23474 ( .A1(n20503), .A2(n20668), .B1(n20667), .B2(n20502), .ZN(
        n20499) );
  AOI22_X1 U23475 ( .A1(P1_INSTQUEUE_REG_11__5__SCAN_IN), .A2(n20504), .B1(
        n20543), .B2(n20669), .ZN(n20498) );
  OAI211_X1 U23476 ( .C1(n20672), .C2(n20507), .A(n20499), .B(n20498), .ZN(
        P1_U3126) );
  AOI22_X1 U23477 ( .A1(n20503), .A2(n20674), .B1(n20673), .B2(n20502), .ZN(
        n20501) );
  AOI22_X1 U23478 ( .A1(P1_INSTQUEUE_REG_11__6__SCAN_IN), .A2(n20504), .B1(
        n20543), .B2(n20675), .ZN(n20500) );
  OAI211_X1 U23479 ( .C1(n20678), .C2(n20507), .A(n20501), .B(n20500), .ZN(
        P1_U3127) );
  AOI22_X1 U23480 ( .A1(n20503), .A2(n20680), .B1(n20679), .B2(n20502), .ZN(
        n20506) );
  AOI22_X1 U23481 ( .A1(P1_INSTQUEUE_REG_11__7__SCAN_IN), .A2(n20504), .B1(
        n20543), .B2(n20682), .ZN(n20505) );
  OAI211_X1 U23482 ( .C1(n20688), .C2(n20507), .A(n20506), .B(n20505), .ZN(
        P1_U3128) );
  INV_X1 U23483 ( .A(n20575), .ZN(n20509) );
  NAND2_X1 U23484 ( .A1(n20509), .A2(n20581), .ZN(n20511) );
  OAI21_X1 U23485 ( .B1(n20511), .B2(n20543), .A(n20510), .ZN(n20518) );
  OR2_X1 U23486 ( .A1(n13655), .A2(n20512), .ZN(n20550) );
  NOR2_X1 U23487 ( .A1(n20550), .A2(n20586), .ZN(n20515) );
  NOR3_X1 U23488 ( .A1(n20514), .A2(n20184), .A3(
        P1_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n20558) );
  NAND2_X1 U23489 ( .A1(n20551), .A2(n20558), .ZN(n20516) );
  INV_X1 U23490 ( .A(n20516), .ZN(n20542) );
  AOI22_X1 U23491 ( .A1(n20575), .A2(n20639), .B1(n20632), .B2(n20542), .ZN(
        n20522) );
  INV_X1 U23492 ( .A(n20515), .ZN(n20517) );
  AOI22_X1 U23493 ( .A1(n20518), .A2(n20517), .B1(P1_STATE2_REG_3__SCAN_IN), 
        .B2(n20516), .ZN(n20519) );
  OAI211_X1 U23494 ( .C1(n20520), .C2(n20691), .A(n20589), .B(n20519), .ZN(
        n20544) );
  AOI22_X1 U23495 ( .A1(P1_INSTQUEUE_REG_12__0__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20592), .ZN(n20521) );
  OAI211_X1 U23496 ( .C1(n20548), .C2(n20523), .A(n20522), .B(n20521), .ZN(
        P1_U3129) );
  AOI22_X1 U23497 ( .A1(n20575), .A2(n20645), .B1(n20643), .B2(n20542), .ZN(
        n20525) );
  AOI22_X1 U23498 ( .A1(P1_INSTQUEUE_REG_12__1__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20596), .ZN(n20524) );
  OAI211_X1 U23499 ( .C1(n20548), .C2(n20526), .A(n20525), .B(n20524), .ZN(
        P1_U3130) );
  AOI22_X1 U23500 ( .A1(n20575), .A2(n20651), .B1(n20649), .B2(n20542), .ZN(
        n20528) );
  AOI22_X1 U23501 ( .A1(P1_INSTQUEUE_REG_12__2__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20600), .ZN(n20527) );
  OAI211_X1 U23502 ( .C1(n20548), .C2(n20529), .A(n20528), .B(n20527), .ZN(
        P1_U3131) );
  AOI22_X1 U23503 ( .A1(n20575), .A2(n20657), .B1(n20655), .B2(n20542), .ZN(
        n20531) );
  AOI22_X1 U23504 ( .A1(P1_INSTQUEUE_REG_12__3__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20604), .ZN(n20530) );
  OAI211_X1 U23505 ( .C1(n20548), .C2(n20532), .A(n20531), .B(n20530), .ZN(
        P1_U3132) );
  AOI22_X1 U23506 ( .A1(n20575), .A2(n20663), .B1(n20661), .B2(n20542), .ZN(
        n20534) );
  AOI22_X1 U23507 ( .A1(P1_INSTQUEUE_REG_12__4__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20608), .ZN(n20533) );
  OAI211_X1 U23508 ( .C1(n20548), .C2(n20535), .A(n20534), .B(n20533), .ZN(
        P1_U3133) );
  AOI22_X1 U23509 ( .A1(n20575), .A2(n20669), .B1(n20667), .B2(n20542), .ZN(
        n20537) );
  AOI22_X1 U23510 ( .A1(P1_INSTQUEUE_REG_12__5__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20612), .ZN(n20536) );
  OAI211_X1 U23511 ( .C1(n20548), .C2(n20538), .A(n20537), .B(n20536), .ZN(
        P1_U3134) );
  AOI22_X1 U23512 ( .A1(n20575), .A2(n20675), .B1(n20673), .B2(n20542), .ZN(
        n20540) );
  AOI22_X1 U23513 ( .A1(P1_INSTQUEUE_REG_12__6__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20616), .ZN(n20539) );
  OAI211_X1 U23514 ( .C1(n20548), .C2(n20541), .A(n20540), .B(n20539), .ZN(
        P1_U3135) );
  AOI22_X1 U23515 ( .A1(n20575), .A2(n20682), .B1(n20679), .B2(n20542), .ZN(
        n20546) );
  AOI22_X1 U23516 ( .A1(P1_INSTQUEUE_REG_12__7__SCAN_IN), .A2(n20544), .B1(
        n20543), .B2(n20622), .ZN(n20545) );
  OAI211_X1 U23517 ( .C1(n20548), .C2(n20547), .A(n20546), .B(n20545), .ZN(
        P1_U3136) );
  INV_X1 U23518 ( .A(n20550), .ZN(n20629) );
  INV_X1 U23519 ( .A(n20558), .ZN(n20553) );
  NOR2_X1 U23520 ( .A1(n20551), .A2(n20553), .ZN(n20573) );
  AOI21_X1 U23521 ( .B1(n20629), .B2(n20552), .A(n20573), .ZN(n20555) );
  OAI22_X1 U23522 ( .A1(n20555), .A2(n20767), .B1(n20553), .B2(n20691), .ZN(
        n20574) );
  AOI22_X1 U23523 ( .A1(n20574), .A2(n20633), .B1(n20632), .B2(n20573), .ZN(
        n20560) );
  INV_X1 U23524 ( .A(n20580), .ZN(n20635) );
  NOR2_X1 U23525 ( .A1(n20635), .A2(n20554), .ZN(n20763) );
  INV_X1 U23526 ( .A(n20763), .ZN(n20556) );
  NAND2_X1 U23527 ( .A1(n20556), .A2(n20555), .ZN(n20557) );
  OAI221_X1 U23528 ( .B1(n20581), .B2(n20558), .C1(n20767), .C2(n20557), .A(
        n20636), .ZN(n20576) );
  AOI22_X1 U23529 ( .A1(P1_INSTQUEUE_REG_13__0__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20592), .ZN(n20559) );
  OAI211_X1 U23530 ( .C1(n20595), .C2(n20591), .A(n20560), .B(n20559), .ZN(
        P1_U3137) );
  AOI22_X1 U23531 ( .A1(n20574), .A2(n20644), .B1(n20643), .B2(n20573), .ZN(
        n20562) );
  AOI22_X1 U23532 ( .A1(P1_INSTQUEUE_REG_13__1__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20596), .ZN(n20561) );
  OAI211_X1 U23533 ( .C1(n20599), .C2(n20591), .A(n20562), .B(n20561), .ZN(
        P1_U3138) );
  AOI22_X1 U23534 ( .A1(n20574), .A2(n20650), .B1(n20649), .B2(n20573), .ZN(
        n20564) );
  AOI22_X1 U23535 ( .A1(P1_INSTQUEUE_REG_13__2__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20600), .ZN(n20563) );
  OAI211_X1 U23536 ( .C1(n20603), .C2(n20591), .A(n20564), .B(n20563), .ZN(
        P1_U3139) );
  AOI22_X1 U23537 ( .A1(n20574), .A2(n20656), .B1(n20655), .B2(n20573), .ZN(
        n20566) );
  AOI22_X1 U23538 ( .A1(P1_INSTQUEUE_REG_13__3__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20604), .ZN(n20565) );
  OAI211_X1 U23539 ( .C1(n20607), .C2(n20591), .A(n20566), .B(n20565), .ZN(
        P1_U3140) );
  AOI22_X1 U23540 ( .A1(n20574), .A2(n20662), .B1(n20661), .B2(n20573), .ZN(
        n20568) );
  AOI22_X1 U23541 ( .A1(P1_INSTQUEUE_REG_13__4__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20608), .ZN(n20567) );
  OAI211_X1 U23542 ( .C1(n20611), .C2(n20591), .A(n20568), .B(n20567), .ZN(
        P1_U3141) );
  AOI22_X1 U23543 ( .A1(n20574), .A2(n20668), .B1(n20667), .B2(n20573), .ZN(
        n20570) );
  AOI22_X1 U23544 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20612), .ZN(n20569) );
  OAI211_X1 U23545 ( .C1(n20615), .C2(n20591), .A(n20570), .B(n20569), .ZN(
        P1_U3142) );
  AOI22_X1 U23546 ( .A1(n20574), .A2(n20674), .B1(n20673), .B2(n20573), .ZN(
        n20572) );
  AOI22_X1 U23547 ( .A1(P1_INSTQUEUE_REG_13__6__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20616), .ZN(n20571) );
  OAI211_X1 U23548 ( .C1(n20619), .C2(n20591), .A(n20572), .B(n20571), .ZN(
        P1_U3143) );
  AOI22_X1 U23549 ( .A1(n20574), .A2(n20680), .B1(n20679), .B2(n20573), .ZN(
        n20578) );
  AOI22_X1 U23550 ( .A1(P1_INSTQUEUE_REG_13__7__SCAN_IN), .A2(n20576), .B1(
        n20575), .B2(n20622), .ZN(n20577) );
  OAI211_X1 U23551 ( .C1(n20627), .C2(n20591), .A(n20578), .B(n20577), .ZN(
        P1_U3144) );
  NAND3_X1 U23552 ( .A1(n20629), .A2(n20586), .A3(n20581), .ZN(n20582) );
  OAI21_X1 U23553 ( .B1(n20584), .B2(n20583), .A(n20582), .ZN(n20621) );
  NOR2_X1 U23554 ( .A1(P1_INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n20630), .ZN(
        n20620) );
  AOI22_X1 U23555 ( .A1(n20621), .A2(n20633), .B1(n20632), .B2(n20620), .ZN(
        n20594) );
  AOI21_X1 U23556 ( .B1(n20591), .B2(n20687), .A(n20765), .ZN(n20585) );
  AOI21_X1 U23557 ( .B1(n20629), .B2(n20586), .A(n20585), .ZN(n20587) );
  NOR2_X1 U23558 ( .A1(n20587), .A2(P1_STATE2_REG_3__SCAN_IN), .ZN(n20590) );
  AOI22_X1 U23559 ( .A1(P1_INSTQUEUE_REG_14__0__SCAN_IN), .A2(n20624), .B1(
        n20623), .B2(n20592), .ZN(n20593) );
  OAI211_X1 U23560 ( .C1(n20595), .C2(n20687), .A(n20594), .B(n20593), .ZN(
        P1_U3145) );
  AOI22_X1 U23561 ( .A1(n20621), .A2(n20644), .B1(n20643), .B2(n20620), .ZN(
        n20598) );
  AOI22_X1 U23562 ( .A1(P1_INSTQUEUE_REG_14__1__SCAN_IN), .A2(n20624), .B1(
        n20623), .B2(n20596), .ZN(n20597) );
  OAI211_X1 U23563 ( .C1(n20599), .C2(n20687), .A(n20598), .B(n20597), .ZN(
        P1_U3146) );
  AOI22_X1 U23564 ( .A1(n20621), .A2(n20650), .B1(n20649), .B2(n20620), .ZN(
        n20602) );
  AOI22_X1 U23565 ( .A1(P1_INSTQUEUE_REG_14__2__SCAN_IN), .A2(n20624), .B1(
        n20623), .B2(n20600), .ZN(n20601) );
  OAI211_X1 U23566 ( .C1(n20603), .C2(n20687), .A(n20602), .B(n20601), .ZN(
        P1_U3147) );
  AOI22_X1 U23567 ( .A1(n20621), .A2(n20656), .B1(n20655), .B2(n20620), .ZN(
        n20606) );
  AOI22_X1 U23568 ( .A1(P1_INSTQUEUE_REG_14__3__SCAN_IN), .A2(n20624), .B1(
        n20623), .B2(n20604), .ZN(n20605) );
  OAI211_X1 U23569 ( .C1(n20607), .C2(n20687), .A(n20606), .B(n20605), .ZN(
        P1_U3148) );
  AOI22_X1 U23570 ( .A1(n20621), .A2(n20662), .B1(n20661), .B2(n20620), .ZN(
        n20610) );
  AOI22_X1 U23571 ( .A1(P1_INSTQUEUE_REG_14__4__SCAN_IN), .A2(n20624), .B1(
        n20623), .B2(n20608), .ZN(n20609) );
  OAI211_X1 U23572 ( .C1(n20611), .C2(n20687), .A(n20610), .B(n20609), .ZN(
        P1_U3149) );
  AOI22_X1 U23573 ( .A1(n20621), .A2(n20668), .B1(n20667), .B2(n20620), .ZN(
        n20614) );
  AOI22_X1 U23574 ( .A1(P1_INSTQUEUE_REG_14__5__SCAN_IN), .A2(n20624), .B1(
        n20623), .B2(n20612), .ZN(n20613) );
  OAI211_X1 U23575 ( .C1(n20615), .C2(n20687), .A(n20614), .B(n20613), .ZN(
        P1_U3150) );
  AOI22_X1 U23576 ( .A1(n20621), .A2(n20674), .B1(n20673), .B2(n20620), .ZN(
        n20618) );
  AOI22_X1 U23577 ( .A1(P1_INSTQUEUE_REG_14__6__SCAN_IN), .A2(n20624), .B1(
        n20623), .B2(n20616), .ZN(n20617) );
  OAI211_X1 U23578 ( .C1(n20619), .C2(n20687), .A(n20618), .B(n20617), .ZN(
        P1_U3151) );
  AOI22_X1 U23579 ( .A1(n20621), .A2(n20680), .B1(n20679), .B2(n20620), .ZN(
        n20626) );
  AOI22_X1 U23580 ( .A1(P1_INSTQUEUE_REG_14__7__SCAN_IN), .A2(n20624), .B1(
        n20623), .B2(n20622), .ZN(n20625) );
  OAI211_X1 U23581 ( .C1(n20627), .C2(n20687), .A(n20626), .B(n20625), .ZN(
        P1_U3152) );
  AOI21_X1 U23582 ( .B1(n20629), .B2(n20628), .A(n11272), .ZN(n20631) );
  OAI22_X1 U23583 ( .A1(n20631), .A2(n20767), .B1(n20630), .B2(n20691), .ZN(
        n20681) );
  AOI22_X1 U23584 ( .A1(n20681), .A2(n20633), .B1(n20632), .B2(n11272), .ZN(
        n20641) );
  NOR3_X1 U23585 ( .A1(n20635), .A2(n20767), .A3(n20634), .ZN(n20637) );
  OAI21_X1 U23586 ( .B1(n20638), .B2(n20637), .A(n20636), .ZN(n20684) );
  AOI22_X1 U23587 ( .A1(P1_INSTQUEUE_REG_15__0__SCAN_IN), .A2(n20684), .B1(
        n20683), .B2(n20639), .ZN(n20640) );
  OAI211_X1 U23588 ( .C1(n20642), .C2(n20687), .A(n20641), .B(n20640), .ZN(
        P1_U3153) );
  AOI22_X1 U23589 ( .A1(n20681), .A2(n20644), .B1(n20643), .B2(n11272), .ZN(
        n20647) );
  AOI22_X1 U23590 ( .A1(P1_INSTQUEUE_REG_15__1__SCAN_IN), .A2(n20684), .B1(
        n20683), .B2(n20645), .ZN(n20646) );
  OAI211_X1 U23591 ( .C1(n20648), .C2(n20687), .A(n20647), .B(n20646), .ZN(
        P1_U3154) );
  AOI22_X1 U23592 ( .A1(n20681), .A2(n20650), .B1(n20649), .B2(n11272), .ZN(
        n20653) );
  AOI22_X1 U23593 ( .A1(P1_INSTQUEUE_REG_15__2__SCAN_IN), .A2(n20684), .B1(
        n20683), .B2(n20651), .ZN(n20652) );
  OAI211_X1 U23594 ( .C1(n20654), .C2(n20687), .A(n20653), .B(n20652), .ZN(
        P1_U3155) );
  AOI22_X1 U23595 ( .A1(n20681), .A2(n20656), .B1(n20655), .B2(n11272), .ZN(
        n20659) );
  AOI22_X1 U23596 ( .A1(P1_INSTQUEUE_REG_15__3__SCAN_IN), .A2(n20684), .B1(
        n20683), .B2(n20657), .ZN(n20658) );
  OAI211_X1 U23597 ( .C1(n20660), .C2(n20687), .A(n20659), .B(n20658), .ZN(
        P1_U3156) );
  AOI22_X1 U23598 ( .A1(n20681), .A2(n20662), .B1(n20661), .B2(n11272), .ZN(
        n20665) );
  AOI22_X1 U23599 ( .A1(P1_INSTQUEUE_REG_15__4__SCAN_IN), .A2(n20684), .B1(
        n20683), .B2(n20663), .ZN(n20664) );
  OAI211_X1 U23600 ( .C1(n20666), .C2(n20687), .A(n20665), .B(n20664), .ZN(
        P1_U3157) );
  AOI22_X1 U23601 ( .A1(n20681), .A2(n20668), .B1(n20667), .B2(n11272), .ZN(
        n20671) );
  AOI22_X1 U23602 ( .A1(P1_INSTQUEUE_REG_15__5__SCAN_IN), .A2(n20684), .B1(
        n20683), .B2(n20669), .ZN(n20670) );
  OAI211_X1 U23603 ( .C1(n20672), .C2(n20687), .A(n20671), .B(n20670), .ZN(
        P1_U3158) );
  AOI22_X1 U23604 ( .A1(n20681), .A2(n20674), .B1(n20673), .B2(n11272), .ZN(
        n20677) );
  AOI22_X1 U23605 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(n20684), .B1(
        n20683), .B2(n20675), .ZN(n20676) );
  OAI211_X1 U23606 ( .C1(n20678), .C2(n20687), .A(n20677), .B(n20676), .ZN(
        P1_U3159) );
  AOI22_X1 U23607 ( .A1(n20681), .A2(n20680), .B1(n20679), .B2(n11272), .ZN(
        n20686) );
  AOI22_X1 U23608 ( .A1(P1_INSTQUEUE_REG_15__7__SCAN_IN), .A2(n20684), .B1(
        n20683), .B2(n20682), .ZN(n20685) );
  OAI211_X1 U23609 ( .C1(n20688), .C2(n20687), .A(n20686), .B(n20685), .ZN(
        P1_U3160) );
  OAI211_X1 U23610 ( .C1(n20692), .C2(n20691), .A(n20690), .B(n20689), .ZN(
        P1_U3163) );
  AND2_X1 U23611 ( .A1(P1_DATAWIDTH_REG_31__SCAN_IN), .A2(n20693), .ZN(
        P1_U3164) );
  AND2_X1 U23612 ( .A1(P1_DATAWIDTH_REG_30__SCAN_IN), .A2(n20693), .ZN(
        P1_U3165) );
  AND2_X1 U23613 ( .A1(P1_DATAWIDTH_REG_29__SCAN_IN), .A2(n20693), .ZN(
        P1_U3166) );
  AND2_X1 U23614 ( .A1(P1_DATAWIDTH_REG_28__SCAN_IN), .A2(n20693), .ZN(
        P1_U3167) );
  AND2_X1 U23615 ( .A1(P1_DATAWIDTH_REG_27__SCAN_IN), .A2(n20693), .ZN(
        P1_U3168) );
  AND2_X1 U23616 ( .A1(P1_DATAWIDTH_REG_26__SCAN_IN), .A2(n20693), .ZN(
        P1_U3169) );
  AND2_X1 U23617 ( .A1(P1_DATAWIDTH_REG_25__SCAN_IN), .A2(n20693), .ZN(
        P1_U3170) );
  AND2_X1 U23618 ( .A1(P1_DATAWIDTH_REG_24__SCAN_IN), .A2(n20693), .ZN(
        P1_U3171) );
  AND2_X1 U23619 ( .A1(P1_DATAWIDTH_REG_23__SCAN_IN), .A2(n20693), .ZN(
        P1_U3172) );
  AND2_X1 U23620 ( .A1(P1_DATAWIDTH_REG_22__SCAN_IN), .A2(n20693), .ZN(
        P1_U3173) );
  INV_X1 U23621 ( .A(P1_DATAWIDTH_REG_21__SCAN_IN), .ZN(n20862) );
  NOR2_X1 U23622 ( .A1(n20756), .A2(n20862), .ZN(P1_U3174) );
  AND2_X1 U23623 ( .A1(P1_DATAWIDTH_REG_20__SCAN_IN), .A2(n20693), .ZN(
        P1_U3175) );
  AND2_X1 U23624 ( .A1(P1_DATAWIDTH_REG_19__SCAN_IN), .A2(n20693), .ZN(
        P1_U3176) );
  AND2_X1 U23625 ( .A1(P1_DATAWIDTH_REG_18__SCAN_IN), .A2(n20693), .ZN(
        P1_U3177) );
  AND2_X1 U23626 ( .A1(P1_DATAWIDTH_REG_17__SCAN_IN), .A2(n20693), .ZN(
        P1_U3178) );
  AND2_X1 U23627 ( .A1(P1_DATAWIDTH_REG_16__SCAN_IN), .A2(n20693), .ZN(
        P1_U3179) );
  AND2_X1 U23628 ( .A1(P1_DATAWIDTH_REG_15__SCAN_IN), .A2(n20693), .ZN(
        P1_U3180) );
  AND2_X1 U23629 ( .A1(P1_DATAWIDTH_REG_14__SCAN_IN), .A2(n20693), .ZN(
        P1_U3181) );
  AND2_X1 U23630 ( .A1(P1_DATAWIDTH_REG_13__SCAN_IN), .A2(n20693), .ZN(
        P1_U3182) );
  AND2_X1 U23631 ( .A1(P1_DATAWIDTH_REG_12__SCAN_IN), .A2(n20693), .ZN(
        P1_U3183) );
  AND2_X1 U23632 ( .A1(P1_DATAWIDTH_REG_11__SCAN_IN), .A2(n20693), .ZN(
        P1_U3184) );
  AND2_X1 U23633 ( .A1(P1_DATAWIDTH_REG_10__SCAN_IN), .A2(n20693), .ZN(
        P1_U3185) );
  INV_X1 U23634 ( .A(P1_DATAWIDTH_REG_9__SCAN_IN), .ZN(n20896) );
  NOR2_X1 U23635 ( .A1(n20756), .A2(n20896), .ZN(P1_U3186) );
  AND2_X1 U23636 ( .A1(P1_DATAWIDTH_REG_8__SCAN_IN), .A2(n20693), .ZN(P1_U3187) );
  AND2_X1 U23637 ( .A1(P1_DATAWIDTH_REG_7__SCAN_IN), .A2(n20693), .ZN(P1_U3188) );
  AND2_X1 U23638 ( .A1(P1_DATAWIDTH_REG_6__SCAN_IN), .A2(n20693), .ZN(P1_U3189) );
  AND2_X1 U23639 ( .A1(P1_DATAWIDTH_REG_5__SCAN_IN), .A2(n20693), .ZN(P1_U3190) );
  AND2_X1 U23640 ( .A1(P1_DATAWIDTH_REG_4__SCAN_IN), .A2(n20693), .ZN(P1_U3191) );
  AND2_X1 U23641 ( .A1(P1_DATAWIDTH_REG_3__SCAN_IN), .A2(n20693), .ZN(P1_U3192) );
  AND2_X1 U23642 ( .A1(P1_DATAWIDTH_REG_2__SCAN_IN), .A2(n20693), .ZN(P1_U3193) );
  NAND2_X1 U23643 ( .A1(P1_STATE_REG_0__SCAN_IN), .A2(n20698), .ZN(n20704) );
  INV_X1 U23644 ( .A(n20704), .ZN(n20697) );
  NOR2_X1 U23645 ( .A1(P1_STATE_REG_1__SCAN_IN), .A2(P1_STATE_REG_2__SCAN_IN), 
        .ZN(n20694) );
  NOR2_X1 U23646 ( .A1(n20694), .A2(n20700), .ZN(n20695) );
  AOI211_X1 U23647 ( .C1(NA), .C2(n20699), .A(n20695), .B(n20960), .ZN(n20696)
         );
  OAI22_X1 U23648 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(n20697), .B1(n20786), 
        .B2(n20696), .ZN(P1_U3194) );
  NOR3_X1 U23649 ( .A1(NA), .A2(n20699), .A3(n20698), .ZN(n20703) );
  AOI21_X1 U23650 ( .B1(P1_REQUESTPENDING_REG_SCAN_IN), .B2(n11119), .A(n20700), .ZN(n20702) );
  AOI222_X1 U23651 ( .A1(n20703), .A2(n20702), .B1(n20703), .B2(
        P1_REQUESTPENDING_REG_SCAN_IN), .C1(n20702), .C2(n20701), .ZN(n20707)
         );
  OAI211_X1 U23652 ( .C1(P1_STATE_REG_1__SCAN_IN), .C2(n20705), .A(
        P1_STATE_REG_2__SCAN_IN), .B(n20704), .ZN(n20706) );
  NAND2_X1 U23653 ( .A1(n20707), .A2(n20706), .ZN(P1_U3196) );
  INV_X1 U23654 ( .A(n20747), .ZN(n20735) );
  NAND2_X1 U23655 ( .A1(n11119), .A2(n20786), .ZN(n20738) );
  INV_X1 U23656 ( .A(n20738), .ZN(n20746) );
  AOI22_X1 U23657 ( .A1(P1_ADDRESS_REG_0__SCAN_IN), .A2(n20798), .B1(
        P1_REIP_REG_2__SCAN_IN), .B2(n20746), .ZN(n20708) );
  OAI21_X1 U23658 ( .B1(n20776), .B2(n20735), .A(n20708), .ZN(P1_U3197) );
  AOI22_X1 U23659 ( .A1(P1_ADDRESS_REG_1__SCAN_IN), .A2(n20798), .B1(
        P1_REIP_REG_3__SCAN_IN), .B2(n20746), .ZN(n20709) );
  OAI21_X1 U23660 ( .B1(n13734), .B2(n20735), .A(n20709), .ZN(P1_U3198) );
  OAI222_X1 U23661 ( .A1(n20735), .A2(n20712), .B1(n20711), .B2(n20786), .C1(
        n20710), .C2(n20738), .ZN(P1_U3199) );
  AOI222_X1 U23662 ( .A1(n20746), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_3__SCAN_IN), .B2(n20784), .C1(P1_REIP_REG_4__SCAN_IN), 
        .C2(n20747), .ZN(n20713) );
  INV_X1 U23663 ( .A(n20713), .ZN(P1_U3200) );
  AOI222_X1 U23664 ( .A1(n20747), .A2(P1_REIP_REG_5__SCAN_IN), .B1(
        P1_ADDRESS_REG_4__SCAN_IN), .B2(n20784), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20746), .ZN(n20714) );
  INV_X1 U23665 ( .A(n20714), .ZN(P1_U3201) );
  AOI222_X1 U23666 ( .A1(n20746), .A2(P1_REIP_REG_7__SCAN_IN), .B1(
        P1_ADDRESS_REG_5__SCAN_IN), .B2(n20784), .C1(P1_REIP_REG_6__SCAN_IN), 
        .C2(n20747), .ZN(n20715) );
  INV_X1 U23667 ( .A(n20715), .ZN(P1_U3202) );
  AOI22_X1 U23668 ( .A1(P1_ADDRESS_REG_6__SCAN_IN), .A2(n20798), .B1(
        P1_REIP_REG_8__SCAN_IN), .B2(n20746), .ZN(n20716) );
  OAI21_X1 U23669 ( .B1(n20717), .B2(n20735), .A(n20716), .ZN(P1_U3203) );
  INV_X1 U23670 ( .A(P1_REIP_REG_8__SCAN_IN), .ZN(n20719) );
  AOI22_X1 U23671 ( .A1(P1_ADDRESS_REG_7__SCAN_IN), .A2(n20798), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20746), .ZN(n20718) );
  OAI21_X1 U23672 ( .B1(n20719), .B2(n20735), .A(n20718), .ZN(P1_U3204) );
  AOI22_X1 U23673 ( .A1(P1_ADDRESS_REG_8__SCAN_IN), .A2(n20798), .B1(
        P1_REIP_REG_9__SCAN_IN), .B2(n20747), .ZN(n20720) );
  OAI21_X1 U23674 ( .B1(n14690), .B2(n20738), .A(n20720), .ZN(P1_U3205) );
  AOI222_X1 U23675 ( .A1(n20747), .A2(P1_REIP_REG_10__SCAN_IN), .B1(
        P1_ADDRESS_REG_9__SCAN_IN), .B2(n20784), .C1(P1_REIP_REG_11__SCAN_IN), 
        .C2(n20746), .ZN(n20721) );
  INV_X1 U23676 ( .A(n20721), .ZN(P1_U3206) );
  AOI222_X1 U23677 ( .A1(n20747), .A2(P1_REIP_REG_11__SCAN_IN), .B1(
        P1_ADDRESS_REG_10__SCAN_IN), .B2(n20784), .C1(P1_REIP_REG_12__SCAN_IN), 
        .C2(n20746), .ZN(n20722) );
  INV_X1 U23678 ( .A(n20722), .ZN(P1_U3207) );
  AOI222_X1 U23679 ( .A1(n20747), .A2(P1_REIP_REG_12__SCAN_IN), .B1(
        P1_ADDRESS_REG_11__SCAN_IN), .B2(n20784), .C1(P1_REIP_REG_13__SCAN_IN), 
        .C2(n20746), .ZN(n20723) );
  INV_X1 U23680 ( .A(n20723), .ZN(P1_U3208) );
  AOI22_X1 U23681 ( .A1(P1_ADDRESS_REG_12__SCAN_IN), .A2(n20798), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20746), .ZN(n20724) );
  OAI21_X1 U23682 ( .B1(n21083), .B2(n20735), .A(n20724), .ZN(P1_U3209) );
  AOI22_X1 U23683 ( .A1(P1_ADDRESS_REG_13__SCAN_IN), .A2(n20798), .B1(
        P1_REIP_REG_14__SCAN_IN), .B2(n20747), .ZN(n20725) );
  OAI21_X1 U23684 ( .B1(n20726), .B2(n20738), .A(n20725), .ZN(P1_U3210) );
  AOI222_X1 U23685 ( .A1(n20747), .A2(P1_REIP_REG_15__SCAN_IN), .B1(
        P1_ADDRESS_REG_14__SCAN_IN), .B2(n20784), .C1(P1_REIP_REG_16__SCAN_IN), 
        .C2(n20746), .ZN(n20727) );
  INV_X1 U23686 ( .A(n20727), .ZN(P1_U3211) );
  AOI222_X1 U23687 ( .A1(n20747), .A2(P1_REIP_REG_16__SCAN_IN), .B1(
        P1_ADDRESS_REG_15__SCAN_IN), .B2(n20784), .C1(P1_REIP_REG_17__SCAN_IN), 
        .C2(n20746), .ZN(n20728) );
  INV_X1 U23688 ( .A(n20728), .ZN(P1_U3212) );
  INV_X1 U23689 ( .A(P1_ADDRESS_REG_16__SCAN_IN), .ZN(n20962) );
  OAI222_X1 U23690 ( .A1(n20735), .A2(n14656), .B1(n20962), .B2(n20786), .C1(
        n20729), .C2(n20738), .ZN(P1_U3213) );
  AOI222_X1 U23691 ( .A1(n20747), .A2(P1_REIP_REG_18__SCAN_IN), .B1(
        P1_ADDRESS_REG_17__SCAN_IN), .B2(n20784), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20746), .ZN(n20730) );
  INV_X1 U23692 ( .A(n20730), .ZN(P1_U3214) );
  AOI222_X1 U23693 ( .A1(n20746), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_18__SCAN_IN), .B2(n20784), .C1(P1_REIP_REG_19__SCAN_IN), 
        .C2(n20747), .ZN(n20731) );
  INV_X1 U23694 ( .A(n20731), .ZN(P1_U3215) );
  AOI222_X1 U23695 ( .A1(n20747), .A2(P1_REIP_REG_20__SCAN_IN), .B1(
        P1_ADDRESS_REG_19__SCAN_IN), .B2(n20784), .C1(P1_REIP_REG_21__SCAN_IN), 
        .C2(n20746), .ZN(n20732) );
  INV_X1 U23696 ( .A(n20732), .ZN(P1_U3216) );
  AOI222_X1 U23697 ( .A1(n20747), .A2(P1_REIP_REG_21__SCAN_IN), .B1(
        P1_ADDRESS_REG_20__SCAN_IN), .B2(n20784), .C1(P1_REIP_REG_22__SCAN_IN), 
        .C2(n20746), .ZN(n20733) );
  INV_X1 U23698 ( .A(n20733), .ZN(P1_U3217) );
  AOI22_X1 U23699 ( .A1(P1_ADDRESS_REG_21__SCAN_IN), .A2(n20798), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20746), .ZN(n20734) );
  OAI21_X1 U23700 ( .B1(n20736), .B2(n20735), .A(n20734), .ZN(P1_U3218) );
  AOI22_X1 U23701 ( .A1(P1_ADDRESS_REG_22__SCAN_IN), .A2(n20798), .B1(
        P1_REIP_REG_23__SCAN_IN), .B2(n20747), .ZN(n20737) );
  OAI21_X1 U23702 ( .B1(n20739), .B2(n20738), .A(n20737), .ZN(P1_U3219) );
  AOI222_X1 U23703 ( .A1(n20747), .A2(P1_REIP_REG_24__SCAN_IN), .B1(
        P1_ADDRESS_REG_23__SCAN_IN), .B2(n20784), .C1(P1_REIP_REG_25__SCAN_IN), 
        .C2(n20746), .ZN(n20740) );
  INV_X1 U23704 ( .A(n20740), .ZN(P1_U3220) );
  AOI222_X1 U23705 ( .A1(n20747), .A2(P1_REIP_REG_25__SCAN_IN), .B1(
        P1_ADDRESS_REG_24__SCAN_IN), .B2(n20784), .C1(P1_REIP_REG_26__SCAN_IN), 
        .C2(n20746), .ZN(n20741) );
  INV_X1 U23706 ( .A(n20741), .ZN(P1_U3221) );
  AOI222_X1 U23707 ( .A1(n20747), .A2(P1_REIP_REG_26__SCAN_IN), .B1(
        P1_ADDRESS_REG_25__SCAN_IN), .B2(n20784), .C1(P1_REIP_REG_27__SCAN_IN), 
        .C2(n20746), .ZN(n20742) );
  INV_X1 U23708 ( .A(n20742), .ZN(P1_U3222) );
  AOI222_X1 U23709 ( .A1(n20747), .A2(P1_REIP_REG_27__SCAN_IN), .B1(
        P1_ADDRESS_REG_26__SCAN_IN), .B2(n20784), .C1(P1_REIP_REG_28__SCAN_IN), 
        .C2(n20746), .ZN(n20743) );
  INV_X1 U23710 ( .A(n20743), .ZN(P1_U3223) );
  AOI222_X1 U23711 ( .A1(n20747), .A2(P1_REIP_REG_28__SCAN_IN), .B1(
        P1_ADDRESS_REG_27__SCAN_IN), .B2(n20784), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20746), .ZN(n20744) );
  INV_X1 U23712 ( .A(n20744), .ZN(P1_U3224) );
  AOI222_X1 U23713 ( .A1(n20746), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_28__SCAN_IN), .B2(n20784), .C1(P1_REIP_REG_29__SCAN_IN), 
        .C2(n20747), .ZN(n20745) );
  INV_X1 U23714 ( .A(n20745), .ZN(P1_U3225) );
  AOI222_X1 U23715 ( .A1(n20747), .A2(P1_REIP_REG_30__SCAN_IN), .B1(
        P1_ADDRESS_REG_29__SCAN_IN), .B2(n20784), .C1(P1_REIP_REG_31__SCAN_IN), 
        .C2(n20746), .ZN(n20748) );
  INV_X1 U23716 ( .A(n20748), .ZN(P1_U3226) );
  OAI22_X1 U23717 ( .A1(n20798), .A2(P1_BYTEENABLE_REG_3__SCAN_IN), .B1(
        P1_BE_N_REG_3__SCAN_IN), .B2(n20786), .ZN(n20749) );
  INV_X1 U23718 ( .A(n20749), .ZN(P1_U3458) );
  OAI22_X1 U23719 ( .A1(n20798), .A2(P1_BYTEENABLE_REG_2__SCAN_IN), .B1(
        P1_BE_N_REG_2__SCAN_IN), .B2(n20786), .ZN(n20750) );
  INV_X1 U23720 ( .A(n20750), .ZN(P1_U3459) );
  OAI22_X1 U23721 ( .A1(n20784), .A2(P1_BYTEENABLE_REG_1__SCAN_IN), .B1(
        P1_BE_N_REG_1__SCAN_IN), .B2(n20786), .ZN(n20751) );
  INV_X1 U23722 ( .A(n20751), .ZN(P1_U3460) );
  OAI22_X1 U23723 ( .A1(n20784), .A2(P1_BYTEENABLE_REG_0__SCAN_IN), .B1(
        P1_BE_N_REG_0__SCAN_IN), .B2(n20786), .ZN(n20752) );
  INV_X1 U23724 ( .A(n20752), .ZN(P1_U3461) );
  OAI21_X1 U23725 ( .B1(P1_DATAWIDTH_REG_0__SCAN_IN), .B2(n20756), .A(n20754), 
        .ZN(n20753) );
  INV_X1 U23726 ( .A(n20753), .ZN(P1_U3464) );
  OAI21_X1 U23727 ( .B1(n20756), .B2(n20755), .A(n20754), .ZN(P1_U3465) );
  OAI22_X1 U23728 ( .A1(n20760), .A2(n20759), .B1(n20758), .B2(n20757), .ZN(
        n20762) );
  MUX2_X1 U23729 ( .A(P1_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n20762), .S(
        n20761), .Z(P1_U3469) );
  INV_X1 U23730 ( .A(n20773), .ZN(n20775) );
  AOI21_X1 U23731 ( .B1(n20769), .B2(n20768), .A(n20767), .ZN(n20770) );
  AOI21_X1 U23732 ( .B1(n20772), .B2(n20771), .A(n20770), .ZN(n20774) );
  AOI22_X1 U23733 ( .A1(n20775), .A2(n20184), .B1(n20774), .B2(n20773), .ZN(
        P1_U3475) );
  AOI21_X1 U23734 ( .B1(P1_REIP_REG_0__SCAN_IN), .B2(
        P1_DATAWIDTH_REG_0__SCAN_IN), .A(P1_DATAWIDTH_REG_1__SCAN_IN), .ZN(
        n20777) );
  AOI22_X1 U23735 ( .A1(P1_REIP_REG_1__SCAN_IN), .A2(P1_REIP_REG_0__SCAN_IN), 
        .B1(n20777), .B2(n20776), .ZN(n20780) );
  INV_X1 U23736 ( .A(P1_BYTEENABLE_REG_2__SCAN_IN), .ZN(n20779) );
  AOI22_X1 U23737 ( .A1(n20783), .A2(n20780), .B1(n20779), .B2(n20778), .ZN(
        P1_U3481) );
  INV_X1 U23738 ( .A(P1_BYTEENABLE_REG_0__SCAN_IN), .ZN(n20782) );
  OAI21_X1 U23739 ( .B1(P1_REIP_REG_1__SCAN_IN), .B2(P1_REIP_REG_0__SCAN_IN), 
        .A(n20783), .ZN(n20781) );
  OAI21_X1 U23740 ( .B1(n20783), .B2(n20782), .A(n20781), .ZN(P1_U3482) );
  AOI22_X1 U23741 ( .A1(n20786), .A2(P1_READREQUEST_REG_SCAN_IN), .B1(n20785), 
        .B2(n20784), .ZN(P1_U3483) );
  INV_X1 U23742 ( .A(n20787), .ZN(n20788) );
  OAI211_X1 U23743 ( .C1(n20791), .C2(n20790), .A(n20789), .B(n20788), .ZN(
        n20797) );
  OAI211_X1 U23744 ( .C1(P1_STATEBS16_REG_SCAN_IN), .C2(n20793), .A(n20792), 
        .B(P1_STATE2_REG_2__SCAN_IN), .ZN(n20794) );
  NAND3_X1 U23745 ( .A1(n20797), .A2(n20795), .A3(n20794), .ZN(n20796) );
  OAI21_X1 U23746 ( .B1(n20797), .B2(n20960), .A(n20796), .ZN(P1_U3485) );
  MUX2_X1 U23747 ( .A(P1_MEMORYFETCH_REG_SCAN_IN), .B(P1_M_IO_N_REG_SCAN_IN), 
        .S(n20798), .Z(P1_U3486) );
  AOI22_X1 U23748 ( .A1(P3_ADDRESS_REG_11__SCAN_IN), .A2(keyinput198), .B1(
        P1_DATAO_REG_14__SCAN_IN), .B2(keyinput128), .ZN(n20799) );
  OAI221_X1 U23749 ( .B1(P3_ADDRESS_REG_11__SCAN_IN), .B2(keyinput198), .C1(
        P1_DATAO_REG_14__SCAN_IN), .C2(keyinput128), .A(n20799), .ZN(n20806)
         );
  AOI22_X1 U23750 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(keyinput239), .B1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(keyinput210), .ZN(n20800) );
  OAI221_X1 U23751 ( .B1(P3_DATAWIDTH_REG_3__SCAN_IN), .B2(keyinput239), .C1(
        P3_PHYADDRPOINTER_REG_22__SCAN_IN), .C2(keyinput210), .A(n20800), .ZN(
        n20805) );
  AOI22_X1 U23752 ( .A1(DATAI_13_), .A2(keyinput155), .B1(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .B2(keyinput213), .ZN(n20801) );
  OAI221_X1 U23753 ( .B1(DATAI_13_), .B2(keyinput155), .C1(
        P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(keyinput213), .A(n20801), 
        .ZN(n20804) );
  AOI22_X1 U23754 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(keyinput251), 
        .B1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .B2(keyinput151), .ZN(n20802) );
  OAI221_X1 U23755 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(keyinput251), 
        .C1(P1_INSTQUEUE_REG_6__6__SCAN_IN), .C2(keyinput151), .A(n20802), 
        .ZN(n20803) );
  NOR4_X1 U23756 ( .A1(n20806), .A2(n20805), .A3(n20804), .A4(n20803), .ZN(
        n20834) );
  AOI22_X1 U23757 ( .A1(P3_DATAO_REG_0__SCAN_IN), .A2(keyinput237), .B1(
        P1_EAX_REG_22__SCAN_IN), .B2(keyinput171), .ZN(n20807) );
  OAI221_X1 U23758 ( .B1(P3_DATAO_REG_0__SCAN_IN), .B2(keyinput237), .C1(
        P1_EAX_REG_22__SCAN_IN), .C2(keyinput171), .A(n20807), .ZN(n20814) );
  AOI22_X1 U23759 ( .A1(P1_LWORD_REG_10__SCAN_IN), .A2(keyinput244), .B1(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(keyinput173), .ZN(n20808) );
  OAI221_X1 U23760 ( .B1(P1_LWORD_REG_10__SCAN_IN), .B2(keyinput244), .C1(
        P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .C2(keyinput173), .A(n20808), 
        .ZN(n20813) );
  AOI22_X1 U23761 ( .A1(P3_EAX_REG_21__SCAN_IN), .A2(keyinput243), .B1(
        P1_INSTQUEUE_REG_13__5__SCAN_IN), .B2(keyinput166), .ZN(n20809) );
  OAI221_X1 U23762 ( .B1(P3_EAX_REG_21__SCAN_IN), .B2(keyinput243), .C1(
        P1_INSTQUEUE_REG_13__5__SCAN_IN), .C2(keyinput166), .A(n20809), .ZN(
        n20812) );
  AOI22_X1 U23763 ( .A1(P3_EAX_REG_12__SCAN_IN), .A2(keyinput140), .B1(
        P3_REIP_REG_1__SCAN_IN), .B2(keyinput149), .ZN(n20810) );
  OAI221_X1 U23764 ( .B1(P3_EAX_REG_12__SCAN_IN), .B2(keyinput140), .C1(
        P3_REIP_REG_1__SCAN_IN), .C2(keyinput149), .A(n20810), .ZN(n20811) );
  NOR4_X1 U23765 ( .A1(n20814), .A2(n20813), .A3(n20812), .A4(n20811), .ZN(
        n20833) );
  AOI22_X1 U23766 ( .A1(BUF2_REG_19__SCAN_IN), .A2(keyinput207), .B1(
        P2_EBX_REG_2__SCAN_IN), .B2(keyinput134), .ZN(n20815) );
  OAI221_X1 U23767 ( .B1(BUF2_REG_19__SCAN_IN), .B2(keyinput207), .C1(
        P2_EBX_REG_2__SCAN_IN), .C2(keyinput134), .A(n20815), .ZN(n20822) );
  AOI22_X1 U23768 ( .A1(P3_ADDRESS_REG_14__SCAN_IN), .A2(keyinput230), .B1(
        P3_EBX_REG_12__SCAN_IN), .B2(keyinput188), .ZN(n20816) );
  OAI221_X1 U23769 ( .B1(P3_ADDRESS_REG_14__SCAN_IN), .B2(keyinput230), .C1(
        P3_EBX_REG_12__SCAN_IN), .C2(keyinput188), .A(n20816), .ZN(n20821) );
  AOI22_X1 U23770 ( .A1(BUF1_REG_6__SCAN_IN), .A2(keyinput252), .B1(
        BUF2_REG_7__SCAN_IN), .B2(keyinput167), .ZN(n20817) );
  OAI221_X1 U23771 ( .B1(BUF1_REG_6__SCAN_IN), .B2(keyinput252), .C1(
        BUF2_REG_7__SCAN_IN), .C2(keyinput167), .A(n20817), .ZN(n20820) );
  AOI22_X1 U23772 ( .A1(P1_CODEFETCH_REG_SCAN_IN), .A2(keyinput203), .B1(
        P2_INSTQUEUE_REG_15__0__SCAN_IN), .B2(keyinput163), .ZN(n20818) );
  OAI221_X1 U23773 ( .B1(P1_CODEFETCH_REG_SCAN_IN), .B2(keyinput203), .C1(
        P2_INSTQUEUE_REG_15__0__SCAN_IN), .C2(keyinput163), .A(n20818), .ZN(
        n20819) );
  NOR4_X1 U23774 ( .A1(n20822), .A2(n20821), .A3(n20820), .A4(n20819), .ZN(
        n20832) );
  AOI22_X1 U23775 ( .A1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(keyinput133), 
        .B1(P1_EAX_REG_21__SCAN_IN), .B2(keyinput250), .ZN(n20823) );
  OAI221_X1 U23776 ( .B1(P3_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(keyinput133), 
        .C1(P1_EAX_REG_21__SCAN_IN), .C2(keyinput250), .A(n20823), .ZN(n20830)
         );
  AOI22_X1 U23777 ( .A1(P3_EAX_REG_6__SCAN_IN), .A2(keyinput225), .B1(
        P2_INSTQUEUE_REG_8__0__SCAN_IN), .B2(keyinput233), .ZN(n20824) );
  OAI221_X1 U23778 ( .B1(P3_EAX_REG_6__SCAN_IN), .B2(keyinput225), .C1(
        P2_INSTQUEUE_REG_8__0__SCAN_IN), .C2(keyinput233), .A(n20824), .ZN(
        n20829) );
  AOI22_X1 U23779 ( .A1(P3_ADDRESS_REG_29__SCAN_IN), .A2(keyinput201), .B1(
        P2_DATAWIDTH_REG_14__SCAN_IN), .B2(keyinput186), .ZN(n20825) );
  OAI221_X1 U23780 ( .B1(P3_ADDRESS_REG_29__SCAN_IN), .B2(keyinput201), .C1(
        P2_DATAWIDTH_REG_14__SCAN_IN), .C2(keyinput186), .A(n20825), .ZN(
        n20828) );
  AOI22_X1 U23781 ( .A1(P3_ADDRESS_REG_8__SCAN_IN), .A2(keyinput209), .B1(
        DATAI_18_), .B2(keyinput152), .ZN(n20826) );
  OAI221_X1 U23782 ( .B1(P3_ADDRESS_REG_8__SCAN_IN), .B2(keyinput209), .C1(
        DATAI_18_), .C2(keyinput152), .A(n20826), .ZN(n20827) );
  NOR4_X1 U23783 ( .A1(n20830), .A2(n20829), .A3(n20828), .A4(n20827), .ZN(
        n20831) );
  NAND4_X1 U23784 ( .A1(n20834), .A2(n20833), .A3(n20832), .A4(n20831), .ZN(
        n20987) );
  AOI22_X1 U23785 ( .A1(P2_DATAWIDTH_REG_24__SCAN_IN), .A2(keyinput147), .B1(
        P3_UWORD_REG_2__SCAN_IN), .B2(keyinput232), .ZN(n20835) );
  OAI221_X1 U23786 ( .B1(P2_DATAWIDTH_REG_24__SCAN_IN), .B2(keyinput147), .C1(
        P3_UWORD_REG_2__SCAN_IN), .C2(keyinput232), .A(n20835), .ZN(n20842) );
  AOI22_X1 U23787 ( .A1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A2(keyinput183), 
        .B1(P2_ADDRESS_REG_10__SCAN_IN), .B2(keyinput228), .ZN(n20836) );
  OAI221_X1 U23788 ( .B1(P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(keyinput183), 
        .C1(P2_ADDRESS_REG_10__SCAN_IN), .C2(keyinput228), .A(n20836), .ZN(
        n20841) );
  AOI22_X1 U23789 ( .A1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .A2(keyinput172), 
        .B1(P2_REIP_REG_28__SCAN_IN), .B2(keyinput182), .ZN(n20837) );
  OAI221_X1 U23790 ( .B1(P1_PHYADDRPOINTER_REG_19__SCAN_IN), .B2(keyinput172), 
        .C1(P2_REIP_REG_28__SCAN_IN), .C2(keyinput182), .A(n20837), .ZN(n20840) );
  AOI22_X1 U23791 ( .A1(P2_ADDRESS_REG_3__SCAN_IN), .A2(keyinput234), .B1(
        P2_INSTQUEUE_REG_10__5__SCAN_IN), .B2(keyinput246), .ZN(n20838) );
  OAI221_X1 U23792 ( .B1(P2_ADDRESS_REG_3__SCAN_IN), .B2(keyinput234), .C1(
        P2_INSTQUEUE_REG_10__5__SCAN_IN), .C2(keyinput246), .A(n20838), .ZN(
        n20839) );
  NOR4_X1 U23793 ( .A1(n20842), .A2(n20841), .A3(n20840), .A4(n20839), .ZN(
        n20874) );
  AOI22_X1 U23794 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(keyinput187), 
        .B1(P1_EBX_REG_19__SCAN_IN), .B2(keyinput148), .ZN(n20843) );
  OAI221_X1 U23795 ( .B1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B2(keyinput187), 
        .C1(P1_EBX_REG_19__SCAN_IN), .C2(keyinput148), .A(n20843), .ZN(n20850)
         );
  AOI22_X1 U23796 ( .A1(P1_BE_N_REG_2__SCAN_IN), .A2(keyinput235), .B1(
        P1_INSTQUEUE_REG_7__2__SCAN_IN), .B2(keyinput197), .ZN(n20844) );
  OAI221_X1 U23797 ( .B1(P1_BE_N_REG_2__SCAN_IN), .B2(keyinput235), .C1(
        P1_INSTQUEUE_REG_7__2__SCAN_IN), .C2(keyinput197), .A(n20844), .ZN(
        n20849) );
  AOI22_X1 U23798 ( .A1(P3_DATAWIDTH_REG_26__SCAN_IN), .A2(keyinput215), .B1(
        P1_REIP_REG_28__SCAN_IN), .B2(keyinput178), .ZN(n20845) );
  OAI221_X1 U23799 ( .B1(P3_DATAWIDTH_REG_26__SCAN_IN), .B2(keyinput215), .C1(
        P1_REIP_REG_28__SCAN_IN), .C2(keyinput178), .A(n20845), .ZN(n20848) );
  AOI22_X1 U23800 ( .A1(P3_DATAO_REG_18__SCAN_IN), .A2(keyinput135), .B1(
        P1_EBX_REG_17__SCAN_IN), .B2(keyinput205), .ZN(n20846) );
  OAI221_X1 U23801 ( .B1(P3_DATAO_REG_18__SCAN_IN), .B2(keyinput135), .C1(
        P1_EBX_REG_17__SCAN_IN), .C2(keyinput205), .A(n20846), .ZN(n20847) );
  NOR4_X1 U23802 ( .A1(n20850), .A2(n20849), .A3(n20848), .A4(n20847), .ZN(
        n20873) );
  AOI22_X1 U23803 ( .A1(DATAI_25_), .A2(keyinput160), .B1(
        P2_EBX_REG_11__SCAN_IN), .B2(keyinput159), .ZN(n20851) );
  OAI221_X1 U23804 ( .B1(DATAI_25_), .B2(keyinput160), .C1(
        P2_EBX_REG_11__SCAN_IN), .C2(keyinput159), .A(n20851), .ZN(n20858) );
  AOI22_X1 U23805 ( .A1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .A2(keyinput141), 
        .B1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .B2(keyinput194), .ZN(n20852)
         );
  OAI221_X1 U23806 ( .B1(P3_PHYADDRPOINTER_REG_8__SCAN_IN), .B2(keyinput141), 
        .C1(P3_PHYADDRPOINTER_REG_20__SCAN_IN), .C2(keyinput194), .A(n20852), 
        .ZN(n20857) );
  AOI22_X1 U23807 ( .A1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .A2(keyinput241), 
        .B1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B2(keyinput153), .ZN(n20853) );
  OAI221_X1 U23808 ( .B1(P1_INSTQUEUE_REG_3__6__SCAN_IN), .B2(keyinput241), 
        .C1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .C2(keyinput153), .A(n20853), 
        .ZN(n20856) );
  AOI22_X1 U23809 ( .A1(P3_DATAO_REG_28__SCAN_IN), .A2(keyinput150), .B1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(keyinput136), .ZN(n20854) );
  OAI221_X1 U23810 ( .B1(P3_DATAO_REG_28__SCAN_IN), .B2(keyinput150), .C1(
        P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .C2(keyinput136), .A(n20854), 
        .ZN(n20855) );
  NOR4_X1 U23811 ( .A1(n20858), .A2(n20857), .A3(n20856), .A4(n20855), .ZN(
        n20872) );
  AOI22_X1 U23812 ( .A1(n21078), .A2(keyinput216), .B1(n20860), .B2(
        keyinput249), .ZN(n20859) );
  OAI221_X1 U23813 ( .B1(n21078), .B2(keyinput216), .C1(n20860), .C2(
        keyinput249), .A(n20859), .ZN(n20870) );
  AOI22_X1 U23814 ( .A1(n13316), .A2(keyinput212), .B1(keyinput191), .B2(
        n20862), .ZN(n20861) );
  OAI221_X1 U23815 ( .B1(n13316), .B2(keyinput212), .C1(n20862), .C2(
        keyinput191), .A(n20861), .ZN(n20869) );
  INV_X1 U23816 ( .A(P2_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n20864) );
  INV_X1 U23817 ( .A(P2_EBX_REG_17__SCAN_IN), .ZN(n20999) );
  AOI22_X1 U23818 ( .A1(n20864), .A2(keyinput176), .B1(keyinput162), .B2(
        n20999), .ZN(n20863) );
  OAI221_X1 U23819 ( .B1(n20864), .B2(keyinput176), .C1(n20999), .C2(
        keyinput162), .A(n20863), .ZN(n20868) );
  INV_X1 U23820 ( .A(P3_DATAO_REG_2__SCAN_IN), .ZN(n20866) );
  AOI22_X1 U23821 ( .A1(n20866), .A2(keyinput169), .B1(n11119), .B2(
        keyinput142), .ZN(n20865) );
  OAI221_X1 U23822 ( .B1(n20866), .B2(keyinput169), .C1(n11119), .C2(
        keyinput142), .A(n20865), .ZN(n20867) );
  NOR4_X1 U23823 ( .A1(n20870), .A2(n20869), .A3(n20868), .A4(n20867), .ZN(
        n20871) );
  NAND4_X1 U23824 ( .A1(n20874), .A2(n20873), .A3(n20872), .A4(n20871), .ZN(
        n20986) );
  AOI22_X1 U23825 ( .A1(n20876), .A2(keyinput208), .B1(n21011), .B2(
        keyinput168), .ZN(n20875) );
  OAI221_X1 U23826 ( .B1(n20876), .B2(keyinput208), .C1(n21011), .C2(
        keyinput168), .A(n20875), .ZN(n20886) );
  INV_X1 U23827 ( .A(P1_INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n21071) );
  INV_X1 U23828 ( .A(P1_INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n21094) );
  AOI22_X1 U23829 ( .A1(n21071), .A2(keyinput242), .B1(keyinput184), .B2(
        n21094), .ZN(n20877) );
  OAI221_X1 U23830 ( .B1(n21071), .B2(keyinput242), .C1(n21094), .C2(
        keyinput184), .A(n20877), .ZN(n20885) );
  AOI22_X1 U23831 ( .A1(n20880), .A2(keyinput193), .B1(n20879), .B2(
        keyinput221), .ZN(n20878) );
  OAI221_X1 U23832 ( .B1(n20880), .B2(keyinput193), .C1(n20879), .C2(
        keyinput221), .A(n20878), .ZN(n20884) );
  INV_X1 U23833 ( .A(P3_LWORD_REG_9__SCAN_IN), .ZN(n20882) );
  AOI22_X1 U23834 ( .A1(n20998), .A2(keyinput236), .B1(keyinput175), .B2(
        n20882), .ZN(n20881) );
  OAI221_X1 U23835 ( .B1(n20998), .B2(keyinput236), .C1(n20882), .C2(
        keyinput175), .A(n20881), .ZN(n20883) );
  NOR4_X1 U23836 ( .A1(n20886), .A2(n20885), .A3(n20884), .A4(n20883), .ZN(
        n20929) );
  INV_X1 U23837 ( .A(P1_INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n20888) );
  INV_X1 U23838 ( .A(P2_BYTEENABLE_REG_2__SCAN_IN), .ZN(n21087) );
  AOI22_X1 U23839 ( .A1(n20888), .A2(keyinput190), .B1(keyinput196), .B2(
        n21087), .ZN(n20887) );
  OAI221_X1 U23840 ( .B1(n20888), .B2(keyinput190), .C1(n21087), .C2(
        keyinput196), .A(n20887), .ZN(n20900) );
  INV_X1 U23841 ( .A(READY2), .ZN(n20890) );
  AOI22_X1 U23842 ( .A1(n20891), .A2(keyinput206), .B1(keyinput195), .B2(
        n20890), .ZN(n20889) );
  OAI221_X1 U23843 ( .B1(n20891), .B2(keyinput206), .C1(n20890), .C2(
        keyinput195), .A(n20889), .ZN(n20899) );
  INV_X1 U23844 ( .A(P1_INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n20894) );
  AOI22_X1 U23845 ( .A1(n20894), .A2(keyinput254), .B1(n20893), .B2(
        keyinput255), .ZN(n20892) );
  OAI221_X1 U23846 ( .B1(n20894), .B2(keyinput254), .C1(n20893), .C2(
        keyinput255), .A(n20892), .ZN(n20898) );
  AOI22_X1 U23847 ( .A1(n20896), .A2(keyinput137), .B1(n21037), .B2(
        keyinput185), .ZN(n20895) );
  OAI221_X1 U23848 ( .B1(n20896), .B2(keyinput137), .C1(n21037), .C2(
        keyinput185), .A(n20895), .ZN(n20897) );
  NOR4_X1 U23849 ( .A1(n20900), .A2(n20899), .A3(n20898), .A4(n20897), .ZN(
        n20928) );
  AOI22_X1 U23850 ( .A1(n21017), .A2(keyinput227), .B1(n20902), .B2(
        keyinput238), .ZN(n20901) );
  OAI221_X1 U23851 ( .B1(n21017), .B2(keyinput227), .C1(n20902), .C2(
        keyinput238), .A(n20901), .ZN(n20912) );
  INV_X1 U23852 ( .A(P2_INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n20904) );
  AOI22_X1 U23853 ( .A1(n20905), .A2(keyinput226), .B1(n20904), .B2(
        keyinput161), .ZN(n20903) );
  OAI221_X1 U23854 ( .B1(n20905), .B2(keyinput226), .C1(n20904), .C2(
        keyinput161), .A(n20903), .ZN(n20911) );
  AOI22_X1 U23855 ( .A1(n20907), .A2(keyinput231), .B1(n21005), .B2(
        keyinput253), .ZN(n20906) );
  OAI221_X1 U23856 ( .B1(n20907), .B2(keyinput231), .C1(n21005), .C2(
        keyinput253), .A(n20906), .ZN(n20910) );
  INV_X1 U23857 ( .A(P3_LWORD_REG_11__SCAN_IN), .ZN(n21021) );
  AOI22_X1 U23858 ( .A1(n14656), .A2(keyinput154), .B1(keyinput177), .B2(
        n21021), .ZN(n20908) );
  OAI221_X1 U23859 ( .B1(n14656), .B2(keyinput154), .C1(n21021), .C2(
        keyinput177), .A(n20908), .ZN(n20909) );
  NOR4_X1 U23860 ( .A1(n20912), .A2(n20911), .A3(n20910), .A4(n20909), .ZN(
        n20927) );
  AOI22_X1 U23861 ( .A1(n20914), .A2(keyinput200), .B1(keyinput240), .B2(
        n13545), .ZN(n20913) );
  OAI221_X1 U23862 ( .B1(n20914), .B2(keyinput200), .C1(n13545), .C2(
        keyinput240), .A(n20913), .ZN(n20925) );
  AOI22_X1 U23863 ( .A1(n20916), .A2(keyinput180), .B1(n21048), .B2(
        keyinput131), .ZN(n20915) );
  OAI221_X1 U23864 ( .B1(n20916), .B2(keyinput180), .C1(n21048), .C2(
        keyinput131), .A(n20915), .ZN(n20924) );
  AOI22_X1 U23865 ( .A1(n20919), .A2(keyinput222), .B1(n20918), .B2(
        keyinput170), .ZN(n20917) );
  OAI221_X1 U23866 ( .B1(n20919), .B2(keyinput222), .C1(n20918), .C2(
        keyinput170), .A(n20917), .ZN(n20923) );
  AOI22_X1 U23867 ( .A1(n20921), .A2(keyinput214), .B1(n21034), .B2(
        keyinput202), .ZN(n20920) );
  OAI221_X1 U23868 ( .B1(n20921), .B2(keyinput214), .C1(n21034), .C2(
        keyinput202), .A(n20920), .ZN(n20922) );
  NOR4_X1 U23869 ( .A1(n20925), .A2(n20924), .A3(n20923), .A4(n20922), .ZN(
        n20926) );
  NAND4_X1 U23870 ( .A1(n20929), .A2(n20928), .A3(n20927), .A4(n20926), .ZN(
        n20985) );
  AOI22_X1 U23871 ( .A1(n20931), .A2(keyinput144), .B1(keyinput146), .B2(
        n21068), .ZN(n20930) );
  OAI221_X1 U23872 ( .B1(n20931), .B2(keyinput144), .C1(n21068), .C2(
        keyinput146), .A(n20930), .ZN(n20942) );
  INV_X1 U23873 ( .A(P1_INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n20933) );
  AOI22_X1 U23874 ( .A1(n20934), .A2(keyinput245), .B1(keyinput189), .B2(
        n20933), .ZN(n20932) );
  OAI221_X1 U23875 ( .B1(n20934), .B2(keyinput245), .C1(n20933), .C2(
        keyinput189), .A(n20932), .ZN(n20941) );
  AOI22_X1 U23876 ( .A1(n21080), .A2(keyinput247), .B1(keyinput220), .B2(
        n21002), .ZN(n20935) );
  OAI221_X1 U23877 ( .B1(n21080), .B2(keyinput247), .C1(n21002), .C2(
        keyinput220), .A(n20935), .ZN(n20940) );
  INV_X1 U23878 ( .A(DATAI_10_), .ZN(n20938) );
  AOI22_X1 U23879 ( .A1(n20938), .A2(keyinput174), .B1(keyinput218), .B2(
        n20937), .ZN(n20936) );
  OAI221_X1 U23880 ( .B1(n20938), .B2(keyinput174), .C1(n20937), .C2(
        keyinput218), .A(n20936), .ZN(n20939) );
  NOR4_X1 U23881 ( .A1(n20942), .A2(n20941), .A3(n20940), .A4(n20939), .ZN(
        n20983) );
  AOI22_X1 U23882 ( .A1(n20945), .A2(keyinput179), .B1(n20944), .B2(
        keyinput132), .ZN(n20943) );
  OAI221_X1 U23883 ( .B1(n20945), .B2(keyinput179), .C1(n20944), .C2(
        keyinput132), .A(n20943), .ZN(n20956) );
  INV_X1 U23884 ( .A(BUF2_REG_13__SCAN_IN), .ZN(n20948) );
  AOI22_X1 U23885 ( .A1(n20948), .A2(keyinput158), .B1(keyinput139), .B2(
        n20947), .ZN(n20946) );
  OAI221_X1 U23886 ( .B1(n20948), .B2(keyinput158), .C1(n20947), .C2(
        keyinput139), .A(n20946), .ZN(n20955) );
  INV_X1 U23887 ( .A(P1_INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n21065) );
  AOI22_X1 U23888 ( .A1(n21065), .A2(keyinput229), .B1(n20950), .B2(
        keyinput165), .ZN(n20949) );
  OAI221_X1 U23889 ( .B1(n21065), .B2(keyinput229), .C1(n20950), .C2(
        keyinput165), .A(n20949), .ZN(n20954) );
  AOI22_X1 U23890 ( .A1(n20952), .A2(keyinput204), .B1(keyinput138), .B2(
        n21103), .ZN(n20951) );
  OAI221_X1 U23891 ( .B1(n20952), .B2(keyinput204), .C1(n21103), .C2(
        keyinput138), .A(n20951), .ZN(n20953) );
  NOR4_X1 U23892 ( .A1(n20956), .A2(n20955), .A3(n20954), .A4(n20953), .ZN(
        n20982) );
  AOI22_X1 U23893 ( .A1(n21084), .A2(keyinput129), .B1(keyinput181), .B2(
        n15074), .ZN(n20957) );
  OAI221_X1 U23894 ( .B1(n21084), .B2(keyinput129), .C1(n15074), .C2(
        keyinput181), .A(n20957), .ZN(n20966) );
  INV_X1 U23895 ( .A(P1_UWORD_REG_5__SCAN_IN), .ZN(n21100) );
  INV_X1 U23896 ( .A(P3_UWORD_REG_12__SCAN_IN), .ZN(n21057) );
  AOI22_X1 U23897 ( .A1(n21100), .A2(keyinput248), .B1(keyinput211), .B2(
        n21057), .ZN(n20958) );
  OAI221_X1 U23898 ( .B1(n21100), .B2(keyinput248), .C1(n21057), .C2(
        keyinput211), .A(n20958), .ZN(n20965) );
  AOI22_X1 U23899 ( .A1(n20960), .A2(keyinput143), .B1(n21083), .B2(
        keyinput145), .ZN(n20959) );
  OAI221_X1 U23900 ( .B1(n20960), .B2(keyinput143), .C1(n21083), .C2(
        keyinput145), .A(n20959), .ZN(n20964) );
  AOI22_X1 U23901 ( .A1(n21093), .A2(keyinput192), .B1(keyinput157), .B2(
        n20962), .ZN(n20961) );
  OAI221_X1 U23902 ( .B1(n21093), .B2(keyinput192), .C1(n20962), .C2(
        keyinput157), .A(n20961), .ZN(n20963) );
  NOR4_X1 U23903 ( .A1(n20966), .A2(n20965), .A3(n20964), .A4(n20963), .ZN(
        n20981) );
  INV_X1 U23904 ( .A(P1_INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n20968) );
  AOI22_X1 U23905 ( .A1(n20969), .A2(keyinput199), .B1(n20968), .B2(
        keyinput219), .ZN(n20967) );
  OAI221_X1 U23906 ( .B1(n20969), .B2(keyinput199), .C1(n20968), .C2(
        keyinput219), .A(n20967), .ZN(n20979) );
  INV_X1 U23907 ( .A(P2_INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n21077) );
  INV_X1 U23908 ( .A(P1_PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n21033) );
  AOI22_X1 U23909 ( .A1(n21077), .A2(keyinput156), .B1(keyinput164), .B2(
        n21033), .ZN(n20970) );
  OAI221_X1 U23910 ( .B1(n21077), .B2(keyinput156), .C1(n21033), .C2(
        keyinput164), .A(n20970), .ZN(n20978) );
  AOI22_X1 U23911 ( .A1(n21015), .A2(keyinput224), .B1(keyinput223), .B2(
        n20972), .ZN(n20971) );
  OAI221_X1 U23912 ( .B1(n21015), .B2(keyinput224), .C1(n20972), .C2(
        keyinput223), .A(n20971), .ZN(n20977) );
  AOI22_X1 U23913 ( .A1(n20975), .A2(keyinput130), .B1(keyinput217), .B2(
        n20974), .ZN(n20973) );
  OAI221_X1 U23914 ( .B1(n20975), .B2(keyinput130), .C1(n20974), .C2(
        keyinput217), .A(n20973), .ZN(n20976) );
  NOR4_X1 U23915 ( .A1(n20979), .A2(n20978), .A3(n20977), .A4(n20976), .ZN(
        n20980) );
  NAND4_X1 U23916 ( .A1(n20983), .A2(n20982), .A3(n20981), .A4(n20980), .ZN(
        n20984) );
  NOR4_X1 U23917 ( .A1(n20987), .A2(n20986), .A3(n20985), .A4(n20984), .ZN(
        n21189) );
  AOI22_X1 U23918 ( .A1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .A2(keyinput82), 
        .B1(BUF2_REG_7__SCAN_IN), .B2(keyinput39), .ZN(n20988) );
  OAI221_X1 U23919 ( .B1(P3_PHYADDRPOINTER_REG_22__SCAN_IN), .B2(keyinput82), 
        .C1(BUF2_REG_7__SCAN_IN), .C2(keyinput39), .A(n20988), .ZN(n20995) );
  AOI22_X1 U23920 ( .A1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .A2(keyinput95), .B1(
        P2_INSTQUEUE_REG_8__0__SCAN_IN), .B2(keyinput105), .ZN(n20989) );
  OAI221_X1 U23921 ( .B1(P3_INSTQUEUE_REG_8__3__SCAN_IN), .B2(keyinput95), 
        .C1(P2_INSTQUEUE_REG_8__0__SCAN_IN), .C2(keyinput105), .A(n20989), 
        .ZN(n20994) );
  AOI22_X1 U23922 ( .A1(P2_DATAWIDTH_REG_4__SCAN_IN), .A2(keyinput86), .B1(
        P3_INSTQUEUE_REG_2__4__SCAN_IN), .B2(keyinput103), .ZN(n20990) );
  OAI221_X1 U23923 ( .B1(P2_DATAWIDTH_REG_4__SCAN_IN), .B2(keyinput86), .C1(
        P3_INSTQUEUE_REG_2__4__SCAN_IN), .C2(keyinput103), .A(n20990), .ZN(
        n20993) );
  AOI22_X1 U23924 ( .A1(P2_DATAO_REG_1__SCAN_IN), .A2(keyinput90), .B1(
        P1_INSTQUEUE_REG_7__6__SCAN_IN), .B2(keyinput62), .ZN(n20991) );
  OAI221_X1 U23925 ( .B1(P2_DATAO_REG_1__SCAN_IN), .B2(keyinput90), .C1(
        P1_INSTQUEUE_REG_7__6__SCAN_IN), .C2(keyinput62), .A(n20991), .ZN(
        n20992) );
  NOR4_X1 U23926 ( .A1(n20995), .A2(n20994), .A3(n20993), .A4(n20992), .ZN(
        n21045) );
  AOI22_X1 U23927 ( .A1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .A2(keyinput71), .B1(
        P2_ADDRESS_REG_5__SCAN_IN), .B2(keyinput127), .ZN(n20996) );
  OAI221_X1 U23928 ( .B1(P3_INSTQUEUE_REG_1__5__SCAN_IN), .B2(keyinput71), 
        .C1(P2_ADDRESS_REG_5__SCAN_IN), .C2(keyinput127), .A(n20996), .ZN(
        n21009) );
  AOI22_X1 U23929 ( .A1(n20999), .A2(keyinput34), .B1(keyinput108), .B2(n20998), .ZN(n20997) );
  OAI221_X1 U23930 ( .B1(n20999), .B2(keyinput34), .C1(n20998), .C2(
        keyinput108), .A(n20997), .ZN(n21008) );
  INV_X1 U23931 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n21001) );
  AOI22_X1 U23932 ( .A1(n21002), .A2(keyinput92), .B1(keyinput0), .B2(n21001), 
        .ZN(n21000) );
  OAI221_X1 U23933 ( .B1(n21002), .B2(keyinput92), .C1(n21001), .C2(keyinput0), 
        .A(n21000), .ZN(n21007) );
  INV_X1 U23934 ( .A(P3_EBX_REG_12__SCAN_IN), .ZN(n21004) );
  AOI22_X1 U23935 ( .A1(n21005), .A2(keyinput125), .B1(keyinput60), .B2(n21004), .ZN(n21003) );
  OAI221_X1 U23936 ( .B1(n21005), .B2(keyinput125), .C1(n21004), .C2(
        keyinput60), .A(n21003), .ZN(n21006) );
  NOR4_X1 U23937 ( .A1(n21009), .A2(n21008), .A3(n21007), .A4(n21006), .ZN(
        n21044) );
  AOI22_X1 U23938 ( .A1(n21012), .A2(keyinput13), .B1(n21011), .B2(keyinput40), 
        .ZN(n21010) );
  OAI221_X1 U23939 ( .B1(n21012), .B2(keyinput13), .C1(n21011), .C2(keyinput40), .A(n21010), .ZN(n21025) );
  AOI22_X1 U23940 ( .A1(n21015), .A2(keyinput96), .B1(keyinput20), .B2(n21014), 
        .ZN(n21013) );
  OAI221_X1 U23941 ( .B1(n21015), .B2(keyinput96), .C1(n21014), .C2(keyinput20), .A(n21013), .ZN(n21024) );
  AOI22_X1 U23942 ( .A1(n21018), .A2(keyinput31), .B1(keyinput99), .B2(n21017), 
        .ZN(n21016) );
  OAI221_X1 U23943 ( .B1(n21018), .B2(keyinput31), .C1(n21017), .C2(keyinput99), .A(n21016), .ZN(n21023) );
  AOI22_X1 U23944 ( .A1(n21021), .A2(keyinput49), .B1(n21020), .B2(keyinput6), 
        .ZN(n21019) );
  OAI221_X1 U23945 ( .B1(n21021), .B2(keyinput49), .C1(n21020), .C2(keyinput6), 
        .A(n21019), .ZN(n21022) );
  NOR4_X1 U23946 ( .A1(n21025), .A2(n21024), .A3(n21023), .A4(n21022), .ZN(
        n21043) );
  INV_X1 U23947 ( .A(P1_INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n21027) );
  AOI22_X1 U23948 ( .A1(n21028), .A2(keyinput35), .B1(keyinput23), .B2(n21027), 
        .ZN(n21026) );
  OAI221_X1 U23949 ( .B1(n21028), .B2(keyinput35), .C1(n21027), .C2(keyinput23), .A(n21026), .ZN(n21041) );
  INV_X1 U23950 ( .A(P1_INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n21031) );
  AOI22_X1 U23951 ( .A1(n21031), .A2(keyinput69), .B1(n21030), .B2(keyinput100), .ZN(n21029) );
  OAI221_X1 U23952 ( .B1(n21031), .B2(keyinput69), .C1(n21030), .C2(
        keyinput100), .A(n21029), .ZN(n21040) );
  AOI22_X1 U23953 ( .A1(n21034), .A2(keyinput74), .B1(n21033), .B2(keyinput36), 
        .ZN(n21032) );
  OAI221_X1 U23954 ( .B1(n21034), .B2(keyinput74), .C1(n21033), .C2(keyinput36), .A(n21032), .ZN(n21039) );
  INV_X1 U23955 ( .A(P3_DATAO_REG_18__SCAN_IN), .ZN(n21036) );
  AOI22_X1 U23956 ( .A1(n21037), .A2(keyinput57), .B1(keyinput7), .B2(n21036), 
        .ZN(n21035) );
  OAI221_X1 U23957 ( .B1(n21037), .B2(keyinput57), .C1(n21036), .C2(keyinput7), 
        .A(n21035), .ZN(n21038) );
  NOR4_X1 U23958 ( .A1(n21041), .A2(n21040), .A3(n21039), .A4(n21038), .ZN(
        n21042) );
  NAND4_X1 U23959 ( .A1(n21045), .A2(n21044), .A3(n21043), .A4(n21042), .ZN(
        n21188) );
  AOI22_X1 U23960 ( .A1(n21048), .A2(keyinput3), .B1(keyinput97), .B2(n21047), 
        .ZN(n21046) );
  OAI221_X1 U23961 ( .B1(n21048), .B2(keyinput3), .C1(n21047), .C2(keyinput97), 
        .A(n21046), .ZN(n21061) );
  INV_X1 U23962 ( .A(P3_DATAO_REG_0__SCAN_IN), .ZN(n21051) );
  AOI22_X1 U23963 ( .A1(n21051), .A2(keyinput109), .B1(n21050), .B2(keyinput66), .ZN(n21049) );
  OAI221_X1 U23964 ( .B1(n21051), .B2(keyinput109), .C1(n21050), .C2(
        keyinput66), .A(n21049), .ZN(n21060) );
  AOI22_X1 U23965 ( .A1(n21054), .A2(keyinput32), .B1(keyinput5), .B2(n21053), 
        .ZN(n21052) );
  OAI221_X1 U23966 ( .B1(n21054), .B2(keyinput32), .C1(n21053), .C2(keyinput5), 
        .A(n21052), .ZN(n21059) );
  INV_X1 U23967 ( .A(DATAI_18_), .ZN(n21056) );
  AOI22_X1 U23968 ( .A1(n21057), .A2(keyinput83), .B1(n21056), .B2(keyinput24), 
        .ZN(n21055) );
  OAI221_X1 U23969 ( .B1(n21057), .B2(keyinput83), .C1(n21056), .C2(keyinput24), .A(n21055), .ZN(n21058) );
  NOR4_X1 U23970 ( .A1(n21061), .A2(n21060), .A3(n21059), .A4(n21058), .ZN(
        n21111) );
  AOI22_X1 U23971 ( .A1(n21063), .A2(keyinput12), .B1(n13545), .B2(keyinput112), .ZN(n21062) );
  OAI221_X1 U23972 ( .B1(n21063), .B2(keyinput12), .C1(n13545), .C2(
        keyinput112), .A(n21062), .ZN(n21075) );
  INV_X1 U23973 ( .A(P1_LWORD_REG_10__SCAN_IN), .ZN(n21066) );
  AOI22_X1 U23974 ( .A1(n21066), .A2(keyinput116), .B1(n21065), .B2(
        keyinput101), .ZN(n21064) );
  OAI221_X1 U23975 ( .B1(n21066), .B2(keyinput116), .C1(n21065), .C2(
        keyinput101), .A(n21064), .ZN(n21074) );
  INV_X1 U23976 ( .A(P3_DATAO_REG_28__SCAN_IN), .ZN(n21069) );
  AOI22_X1 U23977 ( .A1(n21069), .A2(keyinput22), .B1(keyinput18), .B2(n21068), 
        .ZN(n21067) );
  OAI221_X1 U23978 ( .B1(n21069), .B2(keyinput22), .C1(n21068), .C2(keyinput18), .A(n21067), .ZN(n21073) );
  AOI22_X1 U23979 ( .A1(n13126), .A2(keyinput118), .B1(keyinput114), .B2(
        n21071), .ZN(n21070) );
  OAI221_X1 U23980 ( .B1(n13126), .B2(keyinput118), .C1(n21071), .C2(
        keyinput114), .A(n21070), .ZN(n21072) );
  NOR4_X1 U23981 ( .A1(n21075), .A2(n21074), .A3(n21073), .A4(n21072), .ZN(
        n21110) );
  AOI22_X1 U23982 ( .A1(n21078), .A2(keyinput88), .B1(n21077), .B2(keyinput28), 
        .ZN(n21076) );
  OAI221_X1 U23983 ( .B1(n21078), .B2(keyinput88), .C1(n21077), .C2(keyinput28), .A(n21076), .ZN(n21091) );
  AOI22_X1 U23984 ( .A1(n21081), .A2(keyinput19), .B1(n21080), .B2(keyinput119), .ZN(n21079) );
  OAI221_X1 U23985 ( .B1(n21081), .B2(keyinput19), .C1(n21080), .C2(
        keyinput119), .A(n21079), .ZN(n21090) );
  AOI22_X1 U23986 ( .A1(n21084), .A2(keyinput1), .B1(keyinput17), .B2(n21083), 
        .ZN(n21082) );
  OAI221_X1 U23987 ( .B1(n21084), .B2(keyinput1), .C1(n21083), .C2(keyinput17), 
        .A(n21082), .ZN(n21089) );
  INV_X1 U23988 ( .A(P1_INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n21086) );
  AOI22_X1 U23989 ( .A1(n21087), .A2(keyinput68), .B1(n21086), .B2(keyinput113), .ZN(n21085) );
  OAI221_X1 U23990 ( .B1(n21087), .B2(keyinput68), .C1(n21086), .C2(
        keyinput113), .A(n21085), .ZN(n21088) );
  NOR4_X1 U23991 ( .A1(n21091), .A2(n21090), .A3(n21089), .A4(n21088), .ZN(
        n21109) );
  AOI22_X1 U23992 ( .A1(n21094), .A2(keyinput56), .B1(n21093), .B2(keyinput64), 
        .ZN(n21092) );
  OAI221_X1 U23993 ( .B1(n21094), .B2(keyinput56), .C1(n21093), .C2(keyinput64), .A(n21092), .ZN(n21098) );
  XNOR2_X1 U23994 ( .A(n16232), .B(keyinput45), .ZN(n21097) );
  XNOR2_X1 U23995 ( .A(n21095), .B(keyinput106), .ZN(n21096) );
  OR3_X1 U23996 ( .A1(n21098), .A2(n21097), .A3(n21096), .ZN(n21107) );
  AOI22_X1 U23997 ( .A1(n21104), .A2(keyinput81), .B1(n21103), .B2(keyinput10), 
        .ZN(n21102) );
  OAI221_X1 U23998 ( .B1(n21104), .B2(keyinput81), .C1(n21103), .C2(keyinput10), .A(n21102), .ZN(n21105) );
  NOR3_X1 U23999 ( .A1(n21107), .A2(n21106), .A3(n21105), .ZN(n21108) );
  NAND4_X1 U24000 ( .A1(n21111), .A2(n21110), .A3(n21109), .A4(n21108), .ZN(
        n21187) );
  OAI22_X1 U24001 ( .A1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .A2(keyinput91), .B1(
        P1_DATAWIDTH_REG_21__SCAN_IN), .B2(keyinput63), .ZN(n21112) );
  AOI221_X1 U24002 ( .B1(P1_INSTQUEUE_REG_4__7__SCAN_IN), .B2(keyinput91), 
        .C1(keyinput63), .C2(P1_DATAWIDTH_REG_21__SCAN_IN), .A(n21112), .ZN(
        n21119) );
  OAI22_X1 U24003 ( .A1(BUF2_REG_13__SCAN_IN), .A2(keyinput30), .B1(keyinput21), .B2(P3_REIP_REG_1__SCAN_IN), .ZN(n21113) );
  AOI221_X1 U24004 ( .B1(BUF2_REG_13__SCAN_IN), .B2(keyinput30), .C1(
        P3_REIP_REG_1__SCAN_IN), .C2(keyinput21), .A(n21113), .ZN(n21118) );
  OAI22_X1 U24005 ( .A1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(keyinput4), 
        .B1(BUF2_REG_19__SCAN_IN), .B2(keyinput79), .ZN(n21114) );
  AOI221_X1 U24006 ( .B1(P3_INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(keyinput4), 
        .C1(keyinput79), .C2(BUF2_REG_19__SCAN_IN), .A(n21114), .ZN(n21117) );
  OAI22_X1 U24007 ( .A1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .A2(keyinput2), 
        .B1(P1_BE_N_REG_2__SCAN_IN), .B2(keyinput107), .ZN(n21115) );
  AOI221_X1 U24008 ( .B1(P2_PHYADDRPOINTER_REG_14__SCAN_IN), .B2(keyinput2), 
        .C1(keyinput107), .C2(P1_BE_N_REG_2__SCAN_IN), .A(n21115), .ZN(n21116)
         );
  NAND4_X1 U24009 ( .A1(n21119), .A2(n21118), .A3(n21117), .A4(n21116), .ZN(
        n21147) );
  OAI22_X1 U24010 ( .A1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .A2(keyinput33), .B1(
        keyinput124), .B2(BUF1_REG_6__SCAN_IN), .ZN(n21120) );
  AOI221_X1 U24011 ( .B1(P2_INSTQUEUE_REG_5__7__SCAN_IN), .B2(keyinput33), 
        .C1(BUF1_REG_6__SCAN_IN), .C2(keyinput124), .A(n21120), .ZN(n21127) );
  OAI22_X1 U24012 ( .A1(P3_STATE_REG_1__SCAN_IN), .A2(keyinput65), .B1(
        keyinput52), .B2(BUF1_REG_1__SCAN_IN), .ZN(n21121) );
  AOI221_X1 U24013 ( .B1(P3_STATE_REG_1__SCAN_IN), .B2(keyinput65), .C1(
        BUF1_REG_1__SCAN_IN), .C2(keyinput52), .A(n21121), .ZN(n21126) );
  OAI22_X1 U24014 ( .A1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .A2(keyinput110), 
        .B1(keyinput85), .B2(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n21122)
         );
  AOI221_X1 U24015 ( .B1(P2_INSTQUEUE_REG_14__4__SCAN_IN), .B2(keyinput110), 
        .C1(P2_INSTADDRPOINTER_REG_31__SCAN_IN), .C2(keyinput85), .A(n21122), 
        .ZN(n21125) );
  OAI22_X1 U24016 ( .A1(P3_REIP_REG_23__SCAN_IN), .A2(keyinput94), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(keyinput51), .ZN(n21123) );
  AOI221_X1 U24017 ( .B1(P3_REIP_REG_23__SCAN_IN), .B2(keyinput94), .C1(
        keyinput51), .C2(P2_DATAO_REG_10__SCAN_IN), .A(n21123), .ZN(n21124) );
  NAND4_X1 U24018 ( .A1(n21127), .A2(n21126), .A3(n21125), .A4(n21124), .ZN(
        n21146) );
  OAI22_X1 U24019 ( .A1(P3_DATAWIDTH_REG_3__SCAN_IN), .A2(keyinput111), .B1(
        P2_DATAWIDTH_REG_21__SCAN_IN), .B2(keyinput16), .ZN(n21128) );
  AOI221_X1 U24020 ( .B1(P3_DATAWIDTH_REG_3__SCAN_IN), .B2(keyinput111), .C1(
        keyinput16), .C2(P2_DATAWIDTH_REG_21__SCAN_IN), .A(n21128), .ZN(n21135) );
  OAI22_X1 U24021 ( .A1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .A2(keyinput25), .B1(
        keyinput70), .B2(P3_ADDRESS_REG_11__SCAN_IN), .ZN(n21129) );
  AOI221_X1 U24022 ( .B1(P2_INSTQUEUE_REG_6__1__SCAN_IN), .B2(keyinput25), 
        .C1(P3_ADDRESS_REG_11__SCAN_IN), .C2(keyinput70), .A(n21129), .ZN(
        n21134) );
  OAI22_X1 U24023 ( .A1(DATAI_10_), .A2(keyinput46), .B1(P3_EAX_REG_9__SCAN_IN), .B2(keyinput11), .ZN(n21130) );
  AOI221_X1 U24024 ( .B1(DATAI_10_), .B2(keyinput46), .C1(keyinput11), .C2(
        P3_EAX_REG_9__SCAN_IN), .A(n21130), .ZN(n21133) );
  OAI22_X1 U24025 ( .A1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .A2(keyinput61), .B1(
        keyinput115), .B2(P3_EAX_REG_21__SCAN_IN), .ZN(n21131) );
  AOI221_X1 U24026 ( .B1(P1_INSTQUEUE_REG_8__1__SCAN_IN), .B2(keyinput61), 
        .C1(P3_EAX_REG_21__SCAN_IN), .C2(keyinput115), .A(n21131), .ZN(n21132)
         );
  NAND4_X1 U24027 ( .A1(n21135), .A2(n21134), .A3(n21133), .A4(n21132), .ZN(
        n21145) );
  OAI22_X1 U24028 ( .A1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .A2(keyinput123), 
        .B1(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .B2(keyinput121), .ZN(n21136)
         );
  AOI221_X1 U24029 ( .B1(P1_INSTADDRPOINTER_REG_18__SCAN_IN), .B2(keyinput123), 
        .C1(keyinput121), .C2(P3_PHYADDRPOINTER_REG_9__SCAN_IN), .A(n21136), 
        .ZN(n21143) );
  OAI22_X1 U24030 ( .A1(P1_STATE_REG_2__SCAN_IN), .A2(keyinput14), .B1(
        keyinput87), .B2(P3_DATAWIDTH_REG_26__SCAN_IN), .ZN(n21137) );
  AOI221_X1 U24031 ( .B1(P1_STATE_REG_2__SCAN_IN), .B2(keyinput14), .C1(
        P3_DATAWIDTH_REG_26__SCAN_IN), .C2(keyinput87), .A(n21137), .ZN(n21142) );
  OAI22_X1 U24032 ( .A1(P1_REIP_REG_28__SCAN_IN), .A2(keyinput50), .B1(
        keyinput67), .B2(READY2), .ZN(n21138) );
  AOI221_X1 U24033 ( .B1(P1_REIP_REG_28__SCAN_IN), .B2(keyinput50), .C1(READY2), .C2(keyinput67), .A(n21138), .ZN(n21141) );
  OAI22_X1 U24034 ( .A1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .A2(keyinput126), 
        .B1(keyinput53), .B2(BUF1_REG_21__SCAN_IN), .ZN(n21139) );
  AOI221_X1 U24035 ( .B1(P1_INSTQUEUE_REG_15__6__SCAN_IN), .B2(keyinput126), 
        .C1(BUF1_REG_21__SCAN_IN), .C2(keyinput53), .A(n21139), .ZN(n21140) );
  NAND4_X1 U24036 ( .A1(n21143), .A2(n21142), .A3(n21141), .A4(n21140), .ZN(
        n21144) );
  NOR4_X1 U24037 ( .A1(n21147), .A2(n21146), .A3(n21145), .A4(n21144), .ZN(
        n21185) );
  OAI22_X1 U24038 ( .A1(P1_REIP_REG_17__SCAN_IN), .A2(keyinput26), .B1(
        P3_INSTQUEUE_REG_2__6__SCAN_IN), .B2(keyinput42), .ZN(n21148) );
  AOI221_X1 U24039 ( .B1(P1_REIP_REG_17__SCAN_IN), .B2(keyinput26), .C1(
        keyinput42), .C2(P3_INSTQUEUE_REG_2__6__SCAN_IN), .A(n21148), .ZN(
        n21155) );
  OAI22_X1 U24040 ( .A1(P1_ADDRESS_REG_16__SCAN_IN), .A2(keyinput29), .B1(
        keyinput104), .B2(P3_UWORD_REG_2__SCAN_IN), .ZN(n21149) );
  AOI221_X1 U24041 ( .B1(P1_ADDRESS_REG_16__SCAN_IN), .B2(keyinput29), .C1(
        P3_UWORD_REG_2__SCAN_IN), .C2(keyinput104), .A(n21149), .ZN(n21154) );
  OAI22_X1 U24042 ( .A1(P1_EBX_REG_17__SCAN_IN), .A2(keyinput77), .B1(
        P3_INSTQUEUE_REG_14__1__SCAN_IN), .B2(keyinput55), .ZN(n21150) );
  AOI221_X1 U24043 ( .B1(P1_EBX_REG_17__SCAN_IN), .B2(keyinput77), .C1(
        keyinput55), .C2(P3_INSTQUEUE_REG_14__1__SCAN_IN), .A(n21150), .ZN(
        n21153) );
  OAI22_X1 U24044 ( .A1(BUF2_REG_29__SCAN_IN), .A2(keyinput89), .B1(keyinput75), .B2(P1_CODEFETCH_REG_SCAN_IN), .ZN(n21151) );
  AOI221_X1 U24045 ( .B1(BUF2_REG_29__SCAN_IN), .B2(keyinput89), .C1(
        P1_CODEFETCH_REG_SCAN_IN), .C2(keyinput75), .A(n21151), .ZN(n21152) );
  NAND4_X1 U24046 ( .A1(n21155), .A2(n21154), .A3(n21153), .A4(n21152), .ZN(
        n21183) );
  OAI22_X1 U24047 ( .A1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(keyinput8), 
        .B1(P1_DATAWIDTH_REG_9__SCAN_IN), .B2(keyinput9), .ZN(n21156) );
  AOI221_X1 U24048 ( .B1(P1_INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(keyinput8), 
        .C1(keyinput9), .C2(P1_DATAWIDTH_REG_9__SCAN_IN), .A(n21156), .ZN(
        n21163) );
  OAI22_X1 U24049 ( .A1(BUF2_REG_22__SCAN_IN), .A2(keyinput98), .B1(
        P3_ADDRESS_REG_29__SCAN_IN), .B2(keyinput73), .ZN(n21157) );
  AOI221_X1 U24050 ( .B1(BUF2_REG_22__SCAN_IN), .B2(keyinput98), .C1(
        keyinput73), .C2(P3_ADDRESS_REG_29__SCAN_IN), .A(n21157), .ZN(n21162)
         );
  OAI22_X1 U24051 ( .A1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .A2(keyinput59), 
        .B1(keyinput84), .B2(P2_LWORD_REG_5__SCAN_IN), .ZN(n21158) );
  AOI221_X1 U24052 ( .B1(P3_INSTQUEUE_REG_14__4__SCAN_IN), .B2(keyinput59), 
        .C1(P2_LWORD_REG_5__SCAN_IN), .C2(keyinput84), .A(n21158), .ZN(n21161)
         );
  OAI22_X1 U24053 ( .A1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .A2(keyinput48), .B1(
        P1_DATAO_REG_21__SCAN_IN), .B2(keyinput80), .ZN(n21159) );
  AOI221_X1 U24054 ( .B1(P2_INSTQUEUE_REG_8__1__SCAN_IN), .B2(keyinput48), 
        .C1(keyinput80), .C2(P1_DATAO_REG_21__SCAN_IN), .A(n21159), .ZN(n21160) );
  NAND4_X1 U24055 ( .A1(n21163), .A2(n21162), .A3(n21161), .A4(n21160), .ZN(
        n21182) );
  OAI22_X1 U24056 ( .A1(P2_EAX_REG_2__SCAN_IN), .A2(keyinput93), .B1(
        P3_LWORD_REG_9__SCAN_IN), .B2(keyinput47), .ZN(n21164) );
  AOI221_X1 U24057 ( .B1(P2_EAX_REG_2__SCAN_IN), .B2(keyinput93), .C1(
        keyinput47), .C2(P3_LWORD_REG_9__SCAN_IN), .A(n21164), .ZN(n21171) );
  OAI22_X1 U24058 ( .A1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .A2(keyinput38), 
        .B1(P3_ADDRESS_REG_14__SCAN_IN), .B2(keyinput102), .ZN(n21165) );
  AOI221_X1 U24059 ( .B1(P1_INSTQUEUE_REG_13__5__SCAN_IN), .B2(keyinput38), 
        .C1(keyinput102), .C2(P3_ADDRESS_REG_14__SCAN_IN), .A(n21165), .ZN(
        n21170) );
  OAI22_X1 U24060 ( .A1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(keyinput117), 
        .B1(DATAI_13_), .B2(keyinput27), .ZN(n21166) );
  AOI221_X1 U24061 ( .B1(P2_INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(keyinput117), 
        .C1(keyinput27), .C2(DATAI_13_), .A(n21166), .ZN(n21169) );
  OAI22_X1 U24062 ( .A1(P2_REIP_REG_28__SCAN_IN), .A2(keyinput54), .B1(
        keyinput41), .B2(P3_DATAO_REG_2__SCAN_IN), .ZN(n21167) );
  AOI221_X1 U24063 ( .B1(P2_REIP_REG_28__SCAN_IN), .B2(keyinput54), .C1(
        P3_DATAO_REG_2__SCAN_IN), .C2(keyinput41), .A(n21167), .ZN(n21168) );
  NAND4_X1 U24064 ( .A1(n21171), .A2(n21170), .A3(n21169), .A4(n21168), .ZN(
        n21181) );
  OAI22_X1 U24065 ( .A1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .A2(keyinput78), .B1(
        P2_INSTADDRPOINTER_REG_0__SCAN_IN), .B2(keyinput72), .ZN(n21172) );
  AOI221_X1 U24066 ( .B1(P2_INSTQUEUE_REG_0__0__SCAN_IN), .B2(keyinput78), 
        .C1(keyinput72), .C2(P2_INSTADDRPOINTER_REG_0__SCAN_IN), .A(n21172), 
        .ZN(n21179) );
  OAI22_X1 U24067 ( .A1(P1_EAX_REG_22__SCAN_IN), .A2(keyinput43), .B1(
        keyinput15), .B2(P1_REQUESTPENDING_REG_SCAN_IN), .ZN(n21173) );
  AOI221_X1 U24068 ( .B1(P1_EAX_REG_22__SCAN_IN), .B2(keyinput43), .C1(
        P1_REQUESTPENDING_REG_SCAN_IN), .C2(keyinput15), .A(n21173), .ZN(
        n21178) );
  OAI22_X1 U24069 ( .A1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .A2(keyinput37), 
        .B1(keyinput76), .B2(P2_EBX_REG_20__SCAN_IN), .ZN(n21174) );
  AOI221_X1 U24070 ( .B1(P2_PHYADDRPOINTER_REG_2__SCAN_IN), .B2(keyinput37), 
        .C1(P2_EBX_REG_20__SCAN_IN), .C2(keyinput76), .A(n21174), .ZN(n21177)
         );
  OAI22_X1 U24071 ( .A1(P1_EAX_REG_21__SCAN_IN), .A2(keyinput122), .B1(
        P2_DATAWIDTH_REG_14__SCAN_IN), .B2(keyinput58), .ZN(n21175) );
  AOI221_X1 U24072 ( .B1(P1_EAX_REG_21__SCAN_IN), .B2(keyinput122), .C1(
        keyinput58), .C2(P2_DATAWIDTH_REG_14__SCAN_IN), .A(n21175), .ZN(n21176) );
  NAND4_X1 U24073 ( .A1(n21179), .A2(n21178), .A3(n21177), .A4(n21176), .ZN(
        n21180) );
  NOR4_X1 U24074 ( .A1(n21183), .A2(n21182), .A3(n21181), .A4(n21180), .ZN(
        n21184) );
  NAND2_X1 U24075 ( .A1(n21185), .A2(n21184), .ZN(n21186) );
  NOR4_X1 U24076 ( .A1(n21189), .A2(n21188), .A3(n21187), .A4(n21186), .ZN(
        n21191) );
  AOI22_X1 U24077 ( .A1(n16441), .A2(P3_ADDRESS_REG_27__SCAN_IN), .B1(
        P2_ADDRESS_REG_27__SCAN_IN), .B2(n16443), .ZN(n21190) );
  XNOR2_X1 U24078 ( .A(n21191), .B(n21190), .ZN(U357) );
  AND2_X1 U13951 ( .A1(n11004), .A2(n13687), .ZN(n11299) );
  NAND2_X1 U11613 ( .A1(n12562), .A2(n12571), .ZN(n12636) );
  NAND2_X2 U11377 ( .A1(P3_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(n18713), .ZN(
        n11649) );
  NOR2_X1 U11272 ( .A1(n11645), .A2(n11649), .ZN(n11819) );
  CLKBUF_X1 U11268 ( .A(n11047), .Z(n12306) );
  INV_X1 U14695 ( .A(n17006), .ZN(n17069) );
  CLKBUF_X3 U11375 ( .A(n11827), .Z(n9819) );
  AND2_X1 U13773 ( .A1(n10884), .A2(n10873), .ZN(n10879) );
  AND2_X2 U12462 ( .A1(n9837), .A2(P2_INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(
        n10566) );
  CLKBUF_X2 U11262 ( .A(n11199), .Z(n12467) );
  AND2_X1 U11284 ( .A1(n11491), .A2(n20129), .ZN(n11600) );
  AND2_X1 U11315 ( .A1(n12592), .A2(n12636), .ZN(n12659) );
  CLKBUF_X1 U11341 ( .A(n10419), .Z(n12641) );
  CLKBUF_X1 U11358 ( .A(n10416), .Z(n19838) );
  CLKBUF_X1 U11366 ( .A(n11126), .Z(n13486) );
  CLKBUF_X1 U11368 ( .A(n11987), .Z(n20378) );
  CLKBUF_X1 U11606 ( .A(n11121), .Z(n20145) );
  CLKBUF_X1 U12270 ( .A(n15110), .Z(n15111) );
  CLKBUF_X1 U12442 ( .A(n16422), .Z(n16438) );
  OR2_X1 U12513 ( .A1(n10427), .A2(n19139), .ZN(n21192) );
endmodule

