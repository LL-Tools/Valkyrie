

module b21_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, 
        SI_30_, SI_29_, SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, 
        SI_21_, SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_, 
        SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_, 
        SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN, 
        P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN, 
        P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN, 
        P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN, 
        P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN, 
        P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN, 
        P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN, 
        P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN, 
        P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN, 
        P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN, 
        P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN, 
        P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN, 
        P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN, 
        P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN, 
        P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN, 
        P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN, 
        P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN, 
        P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN, 
        P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN, 
        P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN, 
        P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN, 
        P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN, 
        P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN, 
        P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN, 
        P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN, 
        P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN, 
        P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN, 
        P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN, 
        P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN, 
        P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN, 
        P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN, 
        P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN, 
        P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN, 
        P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN, 
        P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN, 
        P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN, 
        P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN, 
        P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN, 
        P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN, 
        P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN, 
        P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN, 
        P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN, 
        P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN, 
        P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN, 
        P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN, 
        P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN, 
        P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN, 
        P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN, 
        P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN, 
        P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN, 
        P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN, P1_REG0_REG_3__SCAN_IN, 
        P1_REG0_REG_4__SCAN_IN, P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN, 
        P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN, P1_REG0_REG_9__SCAN_IN, 
        P1_REG0_REG_10__SCAN_IN, P1_REG0_REG_11__SCAN_IN, 
        P1_REG0_REG_12__SCAN_IN, P1_REG0_REG_13__SCAN_IN, 
        P1_REG0_REG_14__SCAN_IN, P1_REG0_REG_15__SCAN_IN, 
        P1_REG0_REG_16__SCAN_IN, P1_REG0_REG_17__SCAN_IN, 
        P1_REG0_REG_18__SCAN_IN, P1_REG0_REG_19__SCAN_IN, 
        P1_REG0_REG_20__SCAN_IN, P1_REG0_REG_21__SCAN_IN, 
        P1_REG0_REG_22__SCAN_IN, P1_REG0_REG_23__SCAN_IN, 
        P1_REG0_REG_24__SCAN_IN, P1_REG0_REG_25__SCAN_IN, 
        P1_REG0_REG_26__SCAN_IN, P1_REG0_REG_27__SCAN_IN, 
        P1_REG0_REG_28__SCAN_IN, P1_REG0_REG_29__SCAN_IN, 
        P1_REG0_REG_30__SCAN_IN, P1_REG0_REG_31__SCAN_IN, 
        P1_REG1_REG_0__SCAN_IN, P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN, 
        P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN, P1_REG1_REG_5__SCAN_IN, 
        P1_REG1_REG_6__SCAN_IN, P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN, 
        P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN, 
        P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN, 
        P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN, 
        P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN, 
        P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN, 
        P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN, 
        P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN, 
        P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN, 
        P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN, 
        P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN, 
        P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN, 
        P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN, 
        P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN, P1_REG2_REG_3__SCAN_IN, 
        P1_REG2_REG_4__SCAN_IN, P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN, 
        P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN, P1_REG2_REG_9__SCAN_IN, 
        P1_REG2_REG_10__SCAN_IN, P1_REG2_REG_11__SCAN_IN, 
        P1_REG2_REG_12__SCAN_IN, P1_REG2_REG_13__SCAN_IN, 
        P1_REG2_REG_14__SCAN_IN, P1_REG2_REG_15__SCAN_IN, 
        P1_REG2_REG_16__SCAN_IN, P1_REG2_REG_17__SCAN_IN, 
        P1_REG2_REG_18__SCAN_IN, P1_REG2_REG_19__SCAN_IN, 
        P1_REG2_REG_20__SCAN_IN, P1_REG2_REG_21__SCAN_IN, 
        P1_REG2_REG_22__SCAN_IN, P1_REG2_REG_23__SCAN_IN, 
        P1_REG2_REG_24__SCAN_IN, P1_REG2_REG_25__SCAN_IN, 
        P1_REG2_REG_26__SCAN_IN, P1_REG2_REG_27__SCAN_IN, 
        P1_REG2_REG_28__SCAN_IN, P1_REG2_REG_29__SCAN_IN, 
        P1_REG2_REG_30__SCAN_IN, P1_REG2_REG_31__SCAN_IN, 
        P1_ADDR_REG_19__SCAN_IN, P1_ADDR_REG_18__SCAN_IN, 
        P1_ADDR_REG_17__SCAN_IN, P1_ADDR_REG_16__SCAN_IN, 
        P1_ADDR_REG_15__SCAN_IN, P1_ADDR_REG_14__SCAN_IN, 
        P1_ADDR_REG_13__SCAN_IN, P1_ADDR_REG_12__SCAN_IN, 
        P1_ADDR_REG_11__SCAN_IN, P1_ADDR_REG_10__SCAN_IN, 
        P1_ADDR_REG_9__SCAN_IN, P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN, 
        P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN, P1_ADDR_REG_4__SCAN_IN, 
        P1_ADDR_REG_3__SCAN_IN, P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN, 
        P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN, 
        P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN, 
        P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN, 
        P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN, 
        P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN, 
        P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN, 
        P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN, 
        P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN, 
        P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN, 
        P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN, 
        P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN, 
        P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN, 
        P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN, 
        P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN, 
        P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN, 
        P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN, 
        P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN, 
        P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN, 
        P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN, 
        P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN, 
        P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN, 
        P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN, P1_REG3_REG_4__SCAN_IN, 
        P1_REG3_REG_24__SCAN_IN, P1_REG3_REG_17__SCAN_IN, 
        P1_REG3_REG_5__SCAN_IN, P1_REG3_REG_16__SCAN_IN, 
        P1_REG3_REG_25__SCAN_IN, P1_REG3_REG_12__SCAN_IN, 
        P1_REG3_REG_21__SCAN_IN, P1_REG3_REG_1__SCAN_IN, 
        P1_REG3_REG_8__SCAN_IN, P1_REG3_REG_28__SCAN_IN, 
        P1_REG3_REG_19__SCAN_IN, P1_REG3_REG_3__SCAN_IN, 
        P1_REG3_REG_10__SCAN_IN, P1_REG3_REG_23__SCAN_IN, 
        P1_REG3_REG_14__SCAN_IN, P1_REG3_REG_27__SCAN_IN, 
        P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN, P1_RD_REG_SCAN_IN, 
        P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN, P2_IR_REG_1__SCAN_IN, 
        P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN, P2_IR_REG_4__SCAN_IN, 
        P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN, P2_IR_REG_7__SCAN_IN, 
        P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN, P2_IR_REG_10__SCAN_IN, 
        P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN, P2_IR_REG_13__SCAN_IN, 
        P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN, P2_IR_REG_16__SCAN_IN, 
        P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN, P2_IR_REG_19__SCAN_IN, 
        P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN, P2_IR_REG_22__SCAN_IN, 
        P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN, P2_IR_REG_25__SCAN_IN, 
        P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN, P2_IR_REG_28__SCAN_IN, 
        P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN, P2_IR_REG_31__SCAN_IN, 
        P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN, P2_D_REG_2__SCAN_IN, 
        P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN, P2_D_REG_5__SCAN_IN, 
        P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN, P2_D_REG_8__SCAN_IN, 
        P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN, P2_D_REG_11__SCAN_IN, 
        P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN, P2_D_REG_14__SCAN_IN, 
        P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN, P2_D_REG_17__SCAN_IN, 
        P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN, P2_D_REG_20__SCAN_IN, 
        P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN, P2_D_REG_23__SCAN_IN, 
        P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN, P2_D_REG_26__SCAN_IN, 
        P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN, P2_D_REG_29__SCAN_IN, 
        P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN, P2_REG0_REG_0__SCAN_IN, 
        P2_REG0_REG_1__SCAN_IN, P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN, 
        P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN, P2_REG0_REG_6__SCAN_IN, 
        P2_REG0_REG_7__SCAN_IN, P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN, 
        P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN, 
        P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN, 
        P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN, 
        P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN, 
        P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN, 
        P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN, 
        P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN, 
        P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN, 
        P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN, 
        P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN, 
        P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN, 
        P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN, P2_REG1_REG_2__SCAN_IN, 
        P2_REG1_REG_3__SCAN_IN, P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN, 
        P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN, P2_REG1_REG_8__SCAN_IN, 
        P2_REG1_REG_9__SCAN_IN, P2_REG1_REG_10__SCAN_IN, 
        P2_REG1_REG_11__SCAN_IN, P2_REG1_REG_12__SCAN_IN, 
        P2_REG1_REG_13__SCAN_IN, P2_REG1_REG_14__SCAN_IN, 
        P2_REG1_REG_15__SCAN_IN, P2_REG1_REG_16__SCAN_IN, 
        P2_REG1_REG_17__SCAN_IN, P2_REG1_REG_18__SCAN_IN, 
        P2_REG1_REG_19__SCAN_IN, P2_REG1_REG_20__SCAN_IN, 
        P2_REG1_REG_21__SCAN_IN, P2_REG1_REG_22__SCAN_IN, 
        P2_REG1_REG_23__SCAN_IN, P2_REG1_REG_24__SCAN_IN, 
        P2_REG1_REG_25__SCAN_IN, P2_REG1_REG_26__SCAN_IN, 
        P2_REG1_REG_27__SCAN_IN, P2_REG1_REG_28__SCAN_IN, 
        P2_REG1_REG_29__SCAN_IN, P2_REG1_REG_30__SCAN_IN, 
        P2_REG1_REG_31__SCAN_IN, P2_REG2_REG_0__SCAN_IN, 
        P2_REG2_REG_1__SCAN_IN, P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN, 
        P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN, P2_REG2_REG_6__SCAN_IN, 
        P2_REG2_REG_7__SCAN_IN, P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN, 
        P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN, 
        P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN, 
        P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN, 
        P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN, 
        P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN, 
        P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN, 
        P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN, 
        P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN, 
        P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN, 
        P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN, 
        P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN, 
        P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN, 
        P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN, 
        P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN, 
        P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN, 
        P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN, 
        P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN, P2_ADDR_REG_7__SCAN_IN, 
        P2_ADDR_REG_6__SCAN_IN, P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN, 
        P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN, P2_ADDR_REG_1__SCAN_IN, 
        P2_ADDR_REG_0__SCAN_IN, P2_DATAO_REG_0__SCAN_IN, 
        P2_DATAO_REG_1__SCAN_IN, P2_DATAO_REG_2__SCAN_IN, 
        P2_DATAO_REG_3__SCAN_IN, P2_DATAO_REG_4__SCAN_IN, 
        P2_DATAO_REG_5__SCAN_IN, ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, 
        ADD_1071_U57, ADD_1071_U58, ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, 
        ADD_1071_U62, ADD_1071_U63, ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, 
        ADD_1071_U50, ADD_1071_U51, ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, 
        ADD_1071_U5, ADD_1071_U46, U126, U123, P1_U3353, P1_U3352, P1_U3351, 
        P1_U3350, P1_U3349, P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, 
        P1_U3343, P1_U3342, P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, 
        P1_U3336, P1_U3335, P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, 
        P1_U3329, P1_U3328, P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, 
        P1_U3322, P1_U3440, P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, 
        P1_U3317, P1_U3316, P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, 
        P1_U3310, P1_U3309, P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, 
        P1_U3303, P1_U3302, P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, 
        P1_U3296, P1_U3295, P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, 
        P1_U3460, P1_U3463, P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, 
        P1_U3481, P1_U3484, P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, 
        P1_U3502, P1_U3505, P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, 
        P1_U3514, P1_U3515, P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, 
        P1_U3521, P1_U3522, P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, 
        P1_U3528, P1_U3529, P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, 
        P1_U3535, P1_U3536, P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, 
        P1_U3542, P1_U3543, P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, 
        P1_U3549, P1_U3550, P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, 
        P1_U3290, P1_U3289, P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, 
        P1_U3283, P1_U3282, P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, 
        P1_U3276, P1_U3275, P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, 
        P1_U3269, P1_U3268, P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, 
        P1_U3355, P1_U3262, P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, 
        P1_U3256, P1_U3255, P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, 
        P1_U3249, P1_U3248, P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, 
        P1_U3242, P1_U3241, P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, 
        P1_U3560, P1_U3561, P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, 
        P1_U3567, P1_U3568, P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, 
        P1_U3574, P1_U3575, P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, 
        P1_U3581, P1_U3582, P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, 
        P1_U3239, P1_U3238, P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, 
        P1_U3232, P1_U3231, P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, 
        P1_U3225, P1_U3224, P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, 
        P1_U3218, P1_U3217, P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, 
        P1_U3211, P1_U3084, P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, 
        P2_U3355, P2_U3354, P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, 
        P2_U3348, P2_U3347, P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, 
        P2_U3341, P2_U3340, P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, 
        P2_U3334, P2_U3333, P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, 
        P2_U3327, P2_U3437, P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, 
        P2_U3322, P2_U3321, P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, 
        P2_U3315, P2_U3314, P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, 
        P2_U3308, P2_U3307, P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, 
        P2_U3301, P2_U3300, P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, 
        P2_U3457, P2_U3460, P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, 
        P2_U3478, P2_U3481, P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, 
        P2_U3499, P2_U3502, P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, 
        P2_U3511, P2_U3512, P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, 
        P2_U3518, P2_U3519, P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, 
        P2_U3525, P2_U3526, P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, 
        P2_U3532, P2_U3533, P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, 
        P2_U3539, P2_U3540, P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, 
        P2_U3546, P2_U3547, P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, 
        P2_U3295, P2_U3294, P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, 
        P2_U3288, P2_U3287, P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, 
        P2_U3281, P2_U3280, P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, 
        P2_U3274, P2_U3273, P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, 
        P2_U3267, P2_U3266, P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, 
        P2_U3260, P2_U3259, P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, 
        P2_U3253, P2_U3252, P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, 
        P2_U3246, P2_U3245, P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, 
        P2_U3557, P2_U3558, P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, 
        P2_U3564, P2_U3565, P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, 
        P2_U3571, P2_U3572, P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, 
        P2_U3578, P2_U3579, P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, 
        P2_U3243, P2_U3242, P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, 
        P2_U3236, P2_U3235, P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, 
        P2_U3229, P2_U3228, P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, 
        P2_U3222, P2_U3221, P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, 
        P2_U3215, P2_U3152, P2_U3151, P2_U3966 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, P2_WR_REG_SCAN_IN, SI_31_, SI_30_, SI_29_,
         SI_28_, SI_27_, SI_26_, SI_25_, SI_24_, SI_23_, SI_22_, SI_21_,
         SI_20_, SI_19_, SI_18_, SI_17_, SI_16_, SI_15_, SI_14_, SI_13_,
         SI_12_, SI_11_, SI_10_, SI_9_, SI_8_, SI_7_, SI_6_, SI_5_, SI_4_,
         SI_3_, SI_2_, SI_1_, SI_0_, P2_RD_REG_SCAN_IN, P2_STATE_REG_SCAN_IN,
         P2_REG3_REG_7__SCAN_IN, P2_REG3_REG_27__SCAN_IN,
         P2_REG3_REG_14__SCAN_IN, P2_REG3_REG_23__SCAN_IN,
         P2_REG3_REG_10__SCAN_IN, P2_REG3_REG_3__SCAN_IN,
         P2_REG3_REG_19__SCAN_IN, P2_REG3_REG_28__SCAN_IN,
         P2_REG3_REG_8__SCAN_IN, P2_REG3_REG_1__SCAN_IN,
         P2_REG3_REG_21__SCAN_IN, P2_REG3_REG_12__SCAN_IN,
         P2_REG3_REG_25__SCAN_IN, P2_REG3_REG_16__SCAN_IN,
         P2_REG3_REG_5__SCAN_IN, P2_REG3_REG_17__SCAN_IN,
         P2_REG3_REG_24__SCAN_IN, P2_REG3_REG_4__SCAN_IN,
         P2_REG3_REG_9__SCAN_IN, P2_REG3_REG_0__SCAN_IN,
         P2_REG3_REG_20__SCAN_IN, P2_REG3_REG_13__SCAN_IN,
         P2_REG3_REG_22__SCAN_IN, P2_REG3_REG_11__SCAN_IN,
         P2_REG3_REG_2__SCAN_IN, P2_REG3_REG_18__SCAN_IN,
         P2_REG3_REG_6__SCAN_IN, P2_REG3_REG_26__SCAN_IN,
         P2_REG3_REG_15__SCAN_IN, P2_B_REG_SCAN_IN, P2_DATAO_REG_31__SCAN_IN,
         P2_DATAO_REG_30__SCAN_IN, P2_DATAO_REG_29__SCAN_IN,
         P2_DATAO_REG_28__SCAN_IN, P2_DATAO_REG_27__SCAN_IN,
         P2_DATAO_REG_26__SCAN_IN, P2_DATAO_REG_25__SCAN_IN,
         P2_DATAO_REG_24__SCAN_IN, P2_DATAO_REG_23__SCAN_IN,
         P2_DATAO_REG_22__SCAN_IN, P2_DATAO_REG_21__SCAN_IN,
         P2_DATAO_REG_20__SCAN_IN, P2_DATAO_REG_19__SCAN_IN,
         P2_DATAO_REG_18__SCAN_IN, P2_DATAO_REG_17__SCAN_IN,
         P2_DATAO_REG_16__SCAN_IN, P2_DATAO_REG_15__SCAN_IN,
         P2_DATAO_REG_14__SCAN_IN, P2_DATAO_REG_13__SCAN_IN,
         P2_DATAO_REG_12__SCAN_IN, P2_DATAO_REG_11__SCAN_IN,
         P2_DATAO_REG_10__SCAN_IN, P2_DATAO_REG_9__SCAN_IN,
         P2_DATAO_REG_8__SCAN_IN, P2_DATAO_REG_7__SCAN_IN,
         P2_DATAO_REG_6__SCAN_IN, P1_IR_REG_0__SCAN_IN, P1_IR_REG_1__SCAN_IN,
         P1_IR_REG_2__SCAN_IN, P1_IR_REG_3__SCAN_IN, P1_IR_REG_4__SCAN_IN,
         P1_IR_REG_5__SCAN_IN, P1_IR_REG_6__SCAN_IN, P1_IR_REG_7__SCAN_IN,
         P1_IR_REG_8__SCAN_IN, P1_IR_REG_9__SCAN_IN, P1_IR_REG_10__SCAN_IN,
         P1_IR_REG_11__SCAN_IN, P1_IR_REG_12__SCAN_IN, P1_IR_REG_13__SCAN_IN,
         P1_IR_REG_14__SCAN_IN, P1_IR_REG_15__SCAN_IN, P1_IR_REG_16__SCAN_IN,
         P1_IR_REG_17__SCAN_IN, P1_IR_REG_18__SCAN_IN, P1_IR_REG_19__SCAN_IN,
         P1_IR_REG_20__SCAN_IN, P1_IR_REG_21__SCAN_IN, P1_IR_REG_22__SCAN_IN,
         P1_IR_REG_23__SCAN_IN, P1_IR_REG_24__SCAN_IN, P1_IR_REG_25__SCAN_IN,
         P1_IR_REG_26__SCAN_IN, P1_IR_REG_27__SCAN_IN, P1_IR_REG_28__SCAN_IN,
         P1_IR_REG_29__SCAN_IN, P1_IR_REG_30__SCAN_IN, P1_IR_REG_31__SCAN_IN,
         P1_D_REG_0__SCAN_IN, P1_D_REG_1__SCAN_IN, P1_D_REG_2__SCAN_IN,
         P1_D_REG_3__SCAN_IN, P1_D_REG_4__SCAN_IN, P1_D_REG_5__SCAN_IN,
         P1_D_REG_6__SCAN_IN, P1_D_REG_7__SCAN_IN, P1_D_REG_8__SCAN_IN,
         P1_D_REG_9__SCAN_IN, P1_D_REG_10__SCAN_IN, P1_D_REG_11__SCAN_IN,
         P1_D_REG_12__SCAN_IN, P1_D_REG_13__SCAN_IN, P1_D_REG_14__SCAN_IN,
         P1_D_REG_15__SCAN_IN, P1_D_REG_16__SCAN_IN, P1_D_REG_17__SCAN_IN,
         P1_D_REG_18__SCAN_IN, P1_D_REG_19__SCAN_IN, P1_D_REG_20__SCAN_IN,
         P1_D_REG_21__SCAN_IN, P1_D_REG_22__SCAN_IN, P1_D_REG_23__SCAN_IN,
         P1_D_REG_24__SCAN_IN, P1_D_REG_25__SCAN_IN, P1_D_REG_26__SCAN_IN,
         P1_D_REG_27__SCAN_IN, P1_D_REG_28__SCAN_IN, P1_D_REG_29__SCAN_IN,
         P1_D_REG_30__SCAN_IN, P1_D_REG_31__SCAN_IN, P1_REG0_REG_0__SCAN_IN,
         P1_REG0_REG_1__SCAN_IN, P1_REG0_REG_2__SCAN_IN,
         P1_REG0_REG_3__SCAN_IN, P1_REG0_REG_4__SCAN_IN,
         P1_REG0_REG_5__SCAN_IN, P1_REG0_REG_6__SCAN_IN,
         P1_REG0_REG_7__SCAN_IN, P1_REG0_REG_8__SCAN_IN,
         P1_REG0_REG_9__SCAN_IN, P1_REG0_REG_10__SCAN_IN,
         P1_REG0_REG_11__SCAN_IN, P1_REG0_REG_12__SCAN_IN,
         P1_REG0_REG_13__SCAN_IN, P1_REG0_REG_14__SCAN_IN,
         P1_REG0_REG_15__SCAN_IN, P1_REG0_REG_16__SCAN_IN,
         P1_REG0_REG_17__SCAN_IN, P1_REG0_REG_18__SCAN_IN,
         P1_REG0_REG_19__SCAN_IN, P1_REG0_REG_20__SCAN_IN,
         P1_REG0_REG_21__SCAN_IN, P1_REG0_REG_22__SCAN_IN,
         P1_REG0_REG_23__SCAN_IN, P1_REG0_REG_24__SCAN_IN,
         P1_REG0_REG_25__SCAN_IN, P1_REG0_REG_26__SCAN_IN,
         P1_REG0_REG_27__SCAN_IN, P1_REG0_REG_28__SCAN_IN,
         P1_REG0_REG_29__SCAN_IN, P1_REG0_REG_30__SCAN_IN,
         P1_REG0_REG_31__SCAN_IN, P1_REG1_REG_0__SCAN_IN,
         P1_REG1_REG_1__SCAN_IN, P1_REG1_REG_2__SCAN_IN,
         P1_REG1_REG_3__SCAN_IN, P1_REG1_REG_4__SCAN_IN,
         P1_REG1_REG_5__SCAN_IN, P1_REG1_REG_6__SCAN_IN,
         P1_REG1_REG_7__SCAN_IN, P1_REG1_REG_8__SCAN_IN,
         P1_REG1_REG_9__SCAN_IN, P1_REG1_REG_10__SCAN_IN,
         P1_REG1_REG_11__SCAN_IN, P1_REG1_REG_12__SCAN_IN,
         P1_REG1_REG_13__SCAN_IN, P1_REG1_REG_14__SCAN_IN,
         P1_REG1_REG_15__SCAN_IN, P1_REG1_REG_16__SCAN_IN,
         P1_REG1_REG_17__SCAN_IN, P1_REG1_REG_18__SCAN_IN,
         P1_REG1_REG_19__SCAN_IN, P1_REG1_REG_20__SCAN_IN,
         P1_REG1_REG_21__SCAN_IN, P1_REG1_REG_22__SCAN_IN,
         P1_REG1_REG_23__SCAN_IN, P1_REG1_REG_24__SCAN_IN,
         P1_REG1_REG_25__SCAN_IN, P1_REG1_REG_26__SCAN_IN,
         P1_REG1_REG_27__SCAN_IN, P1_REG1_REG_28__SCAN_IN,
         P1_REG1_REG_29__SCAN_IN, P1_REG1_REG_30__SCAN_IN,
         P1_REG1_REG_31__SCAN_IN, P1_REG2_REG_0__SCAN_IN,
         P1_REG2_REG_1__SCAN_IN, P1_REG2_REG_2__SCAN_IN,
         P1_REG2_REG_3__SCAN_IN, P1_REG2_REG_4__SCAN_IN,
         P1_REG2_REG_5__SCAN_IN, P1_REG2_REG_6__SCAN_IN,
         P1_REG2_REG_7__SCAN_IN, P1_REG2_REG_8__SCAN_IN,
         P1_REG2_REG_9__SCAN_IN, P1_REG2_REG_10__SCAN_IN,
         P1_REG2_REG_11__SCAN_IN, P1_REG2_REG_12__SCAN_IN,
         P1_REG2_REG_13__SCAN_IN, P1_REG2_REG_14__SCAN_IN,
         P1_REG2_REG_15__SCAN_IN, P1_REG2_REG_16__SCAN_IN,
         P1_REG2_REG_17__SCAN_IN, P1_REG2_REG_18__SCAN_IN,
         P1_REG2_REG_19__SCAN_IN, P1_REG2_REG_20__SCAN_IN,
         P1_REG2_REG_21__SCAN_IN, P1_REG2_REG_22__SCAN_IN,
         P1_REG2_REG_23__SCAN_IN, P1_REG2_REG_24__SCAN_IN,
         P1_REG2_REG_25__SCAN_IN, P1_REG2_REG_26__SCAN_IN,
         P1_REG2_REG_27__SCAN_IN, P1_REG2_REG_28__SCAN_IN,
         P1_REG2_REG_29__SCAN_IN, P1_REG2_REG_30__SCAN_IN,
         P1_REG2_REG_31__SCAN_IN, P1_ADDR_REG_19__SCAN_IN,
         P1_ADDR_REG_18__SCAN_IN, P1_ADDR_REG_17__SCAN_IN,
         P1_ADDR_REG_16__SCAN_IN, P1_ADDR_REG_15__SCAN_IN,
         P1_ADDR_REG_14__SCAN_IN, P1_ADDR_REG_13__SCAN_IN,
         P1_ADDR_REG_12__SCAN_IN, P1_ADDR_REG_11__SCAN_IN,
         P1_ADDR_REG_10__SCAN_IN, P1_ADDR_REG_9__SCAN_IN,
         P1_ADDR_REG_8__SCAN_IN, P1_ADDR_REG_7__SCAN_IN,
         P1_ADDR_REG_6__SCAN_IN, P1_ADDR_REG_5__SCAN_IN,
         P1_ADDR_REG_4__SCAN_IN, P1_ADDR_REG_3__SCAN_IN,
         P1_ADDR_REG_2__SCAN_IN, P1_ADDR_REG_1__SCAN_IN,
         P1_ADDR_REG_0__SCAN_IN, P1_DATAO_REG_0__SCAN_IN,
         P1_DATAO_REG_1__SCAN_IN, P1_DATAO_REG_2__SCAN_IN,
         P1_DATAO_REG_3__SCAN_IN, P1_DATAO_REG_4__SCAN_IN,
         P1_DATAO_REG_5__SCAN_IN, P1_DATAO_REG_6__SCAN_IN,
         P1_DATAO_REG_7__SCAN_IN, P1_DATAO_REG_8__SCAN_IN,
         P1_DATAO_REG_9__SCAN_IN, P1_DATAO_REG_10__SCAN_IN,
         P1_DATAO_REG_11__SCAN_IN, P1_DATAO_REG_12__SCAN_IN,
         P1_DATAO_REG_13__SCAN_IN, P1_DATAO_REG_14__SCAN_IN,
         P1_DATAO_REG_15__SCAN_IN, P1_DATAO_REG_16__SCAN_IN,
         P1_DATAO_REG_17__SCAN_IN, P1_DATAO_REG_18__SCAN_IN,
         P1_DATAO_REG_19__SCAN_IN, P1_DATAO_REG_20__SCAN_IN,
         P1_DATAO_REG_21__SCAN_IN, P1_DATAO_REG_22__SCAN_IN,
         P1_DATAO_REG_23__SCAN_IN, P1_DATAO_REG_24__SCAN_IN,
         P1_DATAO_REG_25__SCAN_IN, P1_DATAO_REG_26__SCAN_IN,
         P1_DATAO_REG_27__SCAN_IN, P1_DATAO_REG_28__SCAN_IN,
         P1_DATAO_REG_29__SCAN_IN, P1_DATAO_REG_30__SCAN_IN,
         P1_DATAO_REG_31__SCAN_IN, P1_B_REG_SCAN_IN, P1_REG3_REG_15__SCAN_IN,
         P1_REG3_REG_26__SCAN_IN, P1_REG3_REG_6__SCAN_IN,
         P1_REG3_REG_18__SCAN_IN, P1_REG3_REG_2__SCAN_IN,
         P1_REG3_REG_11__SCAN_IN, P1_REG3_REG_22__SCAN_IN,
         P1_REG3_REG_13__SCAN_IN, P1_REG3_REG_20__SCAN_IN,
         P1_REG3_REG_0__SCAN_IN, P1_REG3_REG_9__SCAN_IN,
         P1_REG3_REG_4__SCAN_IN, P1_REG3_REG_24__SCAN_IN,
         P1_REG3_REG_17__SCAN_IN, P1_REG3_REG_5__SCAN_IN,
         P1_REG3_REG_16__SCAN_IN, P1_REG3_REG_25__SCAN_IN,
         P1_REG3_REG_12__SCAN_IN, P1_REG3_REG_21__SCAN_IN,
         P1_REG3_REG_1__SCAN_IN, P1_REG3_REG_8__SCAN_IN,
         P1_REG3_REG_28__SCAN_IN, P1_REG3_REG_19__SCAN_IN,
         P1_REG3_REG_3__SCAN_IN, P1_REG3_REG_10__SCAN_IN,
         P1_REG3_REG_23__SCAN_IN, P1_REG3_REG_14__SCAN_IN,
         P1_REG3_REG_27__SCAN_IN, P1_REG3_REG_7__SCAN_IN, P1_STATE_REG_SCAN_IN,
         P1_RD_REG_SCAN_IN, P1_WR_REG_SCAN_IN, P2_IR_REG_0__SCAN_IN,
         P2_IR_REG_1__SCAN_IN, P2_IR_REG_2__SCAN_IN, P2_IR_REG_3__SCAN_IN,
         P2_IR_REG_4__SCAN_IN, P2_IR_REG_5__SCAN_IN, P2_IR_REG_6__SCAN_IN,
         P2_IR_REG_7__SCAN_IN, P2_IR_REG_8__SCAN_IN, P2_IR_REG_9__SCAN_IN,
         P2_IR_REG_10__SCAN_IN, P2_IR_REG_11__SCAN_IN, P2_IR_REG_12__SCAN_IN,
         P2_IR_REG_13__SCAN_IN, P2_IR_REG_14__SCAN_IN, P2_IR_REG_15__SCAN_IN,
         P2_IR_REG_16__SCAN_IN, P2_IR_REG_17__SCAN_IN, P2_IR_REG_18__SCAN_IN,
         P2_IR_REG_19__SCAN_IN, P2_IR_REG_20__SCAN_IN, P2_IR_REG_21__SCAN_IN,
         P2_IR_REG_22__SCAN_IN, P2_IR_REG_23__SCAN_IN, P2_IR_REG_24__SCAN_IN,
         P2_IR_REG_25__SCAN_IN, P2_IR_REG_26__SCAN_IN, P2_IR_REG_27__SCAN_IN,
         P2_IR_REG_28__SCAN_IN, P2_IR_REG_29__SCAN_IN, P2_IR_REG_30__SCAN_IN,
         P2_IR_REG_31__SCAN_IN, P2_D_REG_0__SCAN_IN, P2_D_REG_1__SCAN_IN,
         P2_D_REG_2__SCAN_IN, P2_D_REG_3__SCAN_IN, P2_D_REG_4__SCAN_IN,
         P2_D_REG_5__SCAN_IN, P2_D_REG_6__SCAN_IN, P2_D_REG_7__SCAN_IN,
         P2_D_REG_8__SCAN_IN, P2_D_REG_9__SCAN_IN, P2_D_REG_10__SCAN_IN,
         P2_D_REG_11__SCAN_IN, P2_D_REG_12__SCAN_IN, P2_D_REG_13__SCAN_IN,
         P2_D_REG_14__SCAN_IN, P2_D_REG_15__SCAN_IN, P2_D_REG_16__SCAN_IN,
         P2_D_REG_17__SCAN_IN, P2_D_REG_18__SCAN_IN, P2_D_REG_19__SCAN_IN,
         P2_D_REG_20__SCAN_IN, P2_D_REG_21__SCAN_IN, P2_D_REG_22__SCAN_IN,
         P2_D_REG_23__SCAN_IN, P2_D_REG_24__SCAN_IN, P2_D_REG_25__SCAN_IN,
         P2_D_REG_26__SCAN_IN, P2_D_REG_27__SCAN_IN, P2_D_REG_28__SCAN_IN,
         P2_D_REG_29__SCAN_IN, P2_D_REG_30__SCAN_IN, P2_D_REG_31__SCAN_IN,
         P2_REG0_REG_0__SCAN_IN, P2_REG0_REG_1__SCAN_IN,
         P2_REG0_REG_2__SCAN_IN, P2_REG0_REG_3__SCAN_IN,
         P2_REG0_REG_4__SCAN_IN, P2_REG0_REG_5__SCAN_IN,
         P2_REG0_REG_6__SCAN_IN, P2_REG0_REG_7__SCAN_IN,
         P2_REG0_REG_8__SCAN_IN, P2_REG0_REG_9__SCAN_IN,
         P2_REG0_REG_10__SCAN_IN, P2_REG0_REG_11__SCAN_IN,
         P2_REG0_REG_12__SCAN_IN, P2_REG0_REG_13__SCAN_IN,
         P2_REG0_REG_14__SCAN_IN, P2_REG0_REG_15__SCAN_IN,
         P2_REG0_REG_16__SCAN_IN, P2_REG0_REG_17__SCAN_IN,
         P2_REG0_REG_18__SCAN_IN, P2_REG0_REG_19__SCAN_IN,
         P2_REG0_REG_20__SCAN_IN, P2_REG0_REG_21__SCAN_IN,
         P2_REG0_REG_22__SCAN_IN, P2_REG0_REG_23__SCAN_IN,
         P2_REG0_REG_24__SCAN_IN, P2_REG0_REG_25__SCAN_IN,
         P2_REG0_REG_26__SCAN_IN, P2_REG0_REG_27__SCAN_IN,
         P2_REG0_REG_28__SCAN_IN, P2_REG0_REG_29__SCAN_IN,
         P2_REG0_REG_30__SCAN_IN, P2_REG0_REG_31__SCAN_IN,
         P2_REG1_REG_0__SCAN_IN, P2_REG1_REG_1__SCAN_IN,
         P2_REG1_REG_2__SCAN_IN, P2_REG1_REG_3__SCAN_IN,
         P2_REG1_REG_4__SCAN_IN, P2_REG1_REG_5__SCAN_IN,
         P2_REG1_REG_6__SCAN_IN, P2_REG1_REG_7__SCAN_IN,
         P2_REG1_REG_8__SCAN_IN, P2_REG1_REG_9__SCAN_IN,
         P2_REG1_REG_10__SCAN_IN, P2_REG1_REG_11__SCAN_IN,
         P2_REG1_REG_12__SCAN_IN, P2_REG1_REG_13__SCAN_IN,
         P2_REG1_REG_14__SCAN_IN, P2_REG1_REG_15__SCAN_IN,
         P2_REG1_REG_16__SCAN_IN, P2_REG1_REG_17__SCAN_IN,
         P2_REG1_REG_18__SCAN_IN, P2_REG1_REG_19__SCAN_IN,
         P2_REG1_REG_20__SCAN_IN, P2_REG1_REG_21__SCAN_IN,
         P2_REG1_REG_22__SCAN_IN, P2_REG1_REG_23__SCAN_IN,
         P2_REG1_REG_24__SCAN_IN, P2_REG1_REG_25__SCAN_IN,
         P2_REG1_REG_26__SCAN_IN, P2_REG1_REG_27__SCAN_IN,
         P2_REG1_REG_28__SCAN_IN, P2_REG1_REG_29__SCAN_IN,
         P2_REG1_REG_30__SCAN_IN, P2_REG1_REG_31__SCAN_IN,
         P2_REG2_REG_0__SCAN_IN, P2_REG2_REG_1__SCAN_IN,
         P2_REG2_REG_2__SCAN_IN, P2_REG2_REG_3__SCAN_IN,
         P2_REG2_REG_4__SCAN_IN, P2_REG2_REG_5__SCAN_IN,
         P2_REG2_REG_6__SCAN_IN, P2_REG2_REG_7__SCAN_IN,
         P2_REG2_REG_8__SCAN_IN, P2_REG2_REG_9__SCAN_IN,
         P2_REG2_REG_10__SCAN_IN, P2_REG2_REG_11__SCAN_IN,
         P2_REG2_REG_12__SCAN_IN, P2_REG2_REG_13__SCAN_IN,
         P2_REG2_REG_14__SCAN_IN, P2_REG2_REG_15__SCAN_IN,
         P2_REG2_REG_16__SCAN_IN, P2_REG2_REG_17__SCAN_IN,
         P2_REG2_REG_18__SCAN_IN, P2_REG2_REG_19__SCAN_IN,
         P2_REG2_REG_20__SCAN_IN, P2_REG2_REG_21__SCAN_IN,
         P2_REG2_REG_22__SCAN_IN, P2_REG2_REG_23__SCAN_IN,
         P2_REG2_REG_24__SCAN_IN, P2_REG2_REG_25__SCAN_IN,
         P2_REG2_REG_26__SCAN_IN, P2_REG2_REG_27__SCAN_IN,
         P2_REG2_REG_28__SCAN_IN, P2_REG2_REG_29__SCAN_IN,
         P2_REG2_REG_30__SCAN_IN, P2_REG2_REG_31__SCAN_IN,
         P2_ADDR_REG_19__SCAN_IN, P2_ADDR_REG_18__SCAN_IN,
         P2_ADDR_REG_17__SCAN_IN, P2_ADDR_REG_16__SCAN_IN,
         P2_ADDR_REG_15__SCAN_IN, P2_ADDR_REG_14__SCAN_IN,
         P2_ADDR_REG_13__SCAN_IN, P2_ADDR_REG_12__SCAN_IN,
         P2_ADDR_REG_11__SCAN_IN, P2_ADDR_REG_10__SCAN_IN,
         P2_ADDR_REG_9__SCAN_IN, P2_ADDR_REG_8__SCAN_IN,
         P2_ADDR_REG_7__SCAN_IN, P2_ADDR_REG_6__SCAN_IN,
         P2_ADDR_REG_5__SCAN_IN, P2_ADDR_REG_4__SCAN_IN,
         P2_ADDR_REG_3__SCAN_IN, P2_ADDR_REG_2__SCAN_IN,
         P2_ADDR_REG_1__SCAN_IN, P2_ADDR_REG_0__SCAN_IN,
         P2_DATAO_REG_0__SCAN_IN, P2_DATAO_REG_1__SCAN_IN,
         P2_DATAO_REG_2__SCAN_IN, P2_DATAO_REG_3__SCAN_IN,
         P2_DATAO_REG_4__SCAN_IN, P2_DATAO_REG_5__SCAN_IN;
  output ADD_1071_U4, ADD_1071_U55, ADD_1071_U56, ADD_1071_U57, ADD_1071_U58,
         ADD_1071_U59, ADD_1071_U60, ADD_1071_U61, ADD_1071_U62, ADD_1071_U63,
         ADD_1071_U47, ADD_1071_U48, ADD_1071_U49, ADD_1071_U50, ADD_1071_U51,
         ADD_1071_U52, ADD_1071_U53, ADD_1071_U54, ADD_1071_U5, ADD_1071_U46,
         U126, U123, P1_U3353, P1_U3352, P1_U3351, P1_U3350, P1_U3349,
         P1_U3348, P1_U3347, P1_U3346, P1_U3345, P1_U3344, P1_U3343, P1_U3342,
         P1_U3341, P1_U3340, P1_U3339, P1_U3338, P1_U3337, P1_U3336, P1_U3335,
         P1_U3334, P1_U3333, P1_U3332, P1_U3331, P1_U3330, P1_U3329, P1_U3328,
         P1_U3327, P1_U3326, P1_U3325, P1_U3324, P1_U3323, P1_U3322, P1_U3440,
         P1_U3441, P1_U3321, P1_U3320, P1_U3319, P1_U3318, P1_U3317, P1_U3316,
         P1_U3315, P1_U3314, P1_U3313, P1_U3312, P1_U3311, P1_U3310, P1_U3309,
         P1_U3308, P1_U3307, P1_U3306, P1_U3305, P1_U3304, P1_U3303, P1_U3302,
         P1_U3301, P1_U3300, P1_U3299, P1_U3298, P1_U3297, P1_U3296, P1_U3295,
         P1_U3294, P1_U3293, P1_U3292, P1_U3454, P1_U3457, P1_U3460, P1_U3463,
         P1_U3466, P1_U3469, P1_U3472, P1_U3475, P1_U3478, P1_U3481, P1_U3484,
         P1_U3487, P1_U3490, P1_U3493, P1_U3496, P1_U3499, P1_U3502, P1_U3505,
         P1_U3508, P1_U3510, P1_U3511, P1_U3512, P1_U3513, P1_U3514, P1_U3515,
         P1_U3516, P1_U3517, P1_U3518, P1_U3519, P1_U3520, P1_U3521, P1_U3522,
         P1_U3523, P1_U3524, P1_U3525, P1_U3526, P1_U3527, P1_U3528, P1_U3529,
         P1_U3530, P1_U3531, P1_U3532, P1_U3533, P1_U3534, P1_U3535, P1_U3536,
         P1_U3537, P1_U3538, P1_U3539, P1_U3540, P1_U3541, P1_U3542, P1_U3543,
         P1_U3544, P1_U3545, P1_U3546, P1_U3547, P1_U3548, P1_U3549, P1_U3550,
         P1_U3551, P1_U3552, P1_U3553, P1_U3554, P1_U3291, P1_U3290, P1_U3289,
         P1_U3288, P1_U3287, P1_U3286, P1_U3285, P1_U3284, P1_U3283, P1_U3282,
         P1_U3281, P1_U3280, P1_U3279, P1_U3278, P1_U3277, P1_U3276, P1_U3275,
         P1_U3274, P1_U3273, P1_U3272, P1_U3271, P1_U3270, P1_U3269, P1_U3268,
         P1_U3267, P1_U3266, P1_U3265, P1_U3264, P1_U3263, P1_U3355, P1_U3262,
         P1_U3261, P1_U3260, P1_U3259, P1_U3258, P1_U3257, P1_U3256, P1_U3255,
         P1_U3254, P1_U3253, P1_U3252, P1_U3251, P1_U3250, P1_U3249, P1_U3248,
         P1_U3247, P1_U3246, P1_U3245, P1_U3244, P1_U3243, P1_U3242, P1_U3241,
         P1_U3555, P1_U3556, P1_U3557, P1_U3558, P1_U3559, P1_U3560, P1_U3561,
         P1_U3562, P1_U3563, P1_U3564, P1_U3565, P1_U3566, P1_U3567, P1_U3568,
         P1_U3569, P1_U3570, P1_U3571, P1_U3572, P1_U3573, P1_U3574, P1_U3575,
         P1_U3576, P1_U3577, P1_U3578, P1_U3579, P1_U3580, P1_U3581, P1_U3582,
         P1_U3583, P1_U3584, P1_U3585, P1_U3586, P1_U3240, P1_U3239, P1_U3238,
         P1_U3237, P1_U3236, P1_U3235, P1_U3234, P1_U3233, P1_U3232, P1_U3231,
         P1_U3230, P1_U3229, P1_U3228, P1_U3227, P1_U3226, P1_U3225, P1_U3224,
         P1_U3223, P1_U3222, P1_U3221, P1_U3220, P1_U3219, P1_U3218, P1_U3217,
         P1_U3216, P1_U3215, P1_U3214, P1_U3213, P1_U3212, P1_U3211, P1_U3084,
         P1_U3083, P1_U4006, P2_U3358, P2_U3357, P2_U3356, P2_U3355, P2_U3354,
         P2_U3353, P2_U3352, P2_U3351, P2_U3350, P2_U3349, P2_U3348, P2_U3347,
         P2_U3346, P2_U3345, P2_U3344, P2_U3343, P2_U3342, P2_U3341, P2_U3340,
         P2_U3339, P2_U3338, P2_U3337, P2_U3336, P2_U3335, P2_U3334, P2_U3333,
         P2_U3332, P2_U3331, P2_U3330, P2_U3329, P2_U3328, P2_U3327, P2_U3437,
         P2_U3438, P2_U3326, P2_U3325, P2_U3324, P2_U3323, P2_U3322, P2_U3321,
         P2_U3320, P2_U3319, P2_U3318, P2_U3317, P2_U3316, P2_U3315, P2_U3314,
         P2_U3313, P2_U3312, P2_U3311, P2_U3310, P2_U3309, P2_U3308, P2_U3307,
         P2_U3306, P2_U3305, P2_U3304, P2_U3303, P2_U3302, P2_U3301, P2_U3300,
         P2_U3299, P2_U3298, P2_U3297, P2_U3451, P2_U3454, P2_U3457, P2_U3460,
         P2_U3463, P2_U3466, P2_U3469, P2_U3472, P2_U3475, P2_U3478, P2_U3481,
         P2_U3484, P2_U3487, P2_U3490, P2_U3493, P2_U3496, P2_U3499, P2_U3502,
         P2_U3505, P2_U3507, P2_U3508, P2_U3509, P2_U3510, P2_U3511, P2_U3512,
         P2_U3513, P2_U3514, P2_U3515, P2_U3516, P2_U3517, P2_U3518, P2_U3519,
         P2_U3520, P2_U3521, P2_U3522, P2_U3523, P2_U3524, P2_U3525, P2_U3526,
         P2_U3527, P2_U3528, P2_U3529, P2_U3530, P2_U3531, P2_U3532, P2_U3533,
         P2_U3534, P2_U3535, P2_U3536, P2_U3537, P2_U3538, P2_U3539, P2_U3540,
         P2_U3541, P2_U3542, P2_U3543, P2_U3544, P2_U3545, P2_U3546, P2_U3547,
         P2_U3548, P2_U3549, P2_U3550, P2_U3551, P2_U3296, P2_U3295, P2_U3294,
         P2_U3293, P2_U3292, P2_U3291, P2_U3290, P2_U3289, P2_U3288, P2_U3287,
         P2_U3286, P2_U3285, P2_U3284, P2_U3283, P2_U3282, P2_U3281, P2_U3280,
         P2_U3279, P2_U3278, P2_U3277, P2_U3276, P2_U3275, P2_U3274, P2_U3273,
         P2_U3272, P2_U3271, P2_U3270, P2_U3269, P2_U3268, P2_U3267, P2_U3266,
         P2_U3265, P2_U3264, P2_U3263, P2_U3262, P2_U3261, P2_U3260, P2_U3259,
         P2_U3258, P2_U3257, P2_U3256, P2_U3255, P2_U3254, P2_U3253, P2_U3252,
         P2_U3251, P2_U3250, P2_U3249, P2_U3248, P2_U3247, P2_U3246, P2_U3245,
         P2_U3552, P2_U3553, P2_U3554, P2_U3555, P2_U3556, P2_U3557, P2_U3558,
         P2_U3559, P2_U3560, P2_U3561, P2_U3562, P2_U3563, P2_U3564, P2_U3565,
         P2_U3566, P2_U3567, P2_U3568, P2_U3569, P2_U3570, P2_U3571, P2_U3572,
         P2_U3573, P2_U3574, P2_U3575, P2_U3576, P2_U3577, P2_U3578, P2_U3579,
         P2_U3580, P2_U3581, P2_U3582, P2_U3583, P2_U3244, P2_U3243, P2_U3242,
         P2_U3241, P2_U3240, P2_U3239, P2_U3238, P2_U3237, P2_U3236, P2_U3235,
         P2_U3234, P2_U3233, P2_U3232, P2_U3231, P2_U3230, P2_U3229, P2_U3228,
         P2_U3227, P2_U3226, P2_U3225, P2_U3224, P2_U3223, P2_U3222, P2_U3221,
         P2_U3220, P2_U3219, P2_U3218, P2_U3217, P2_U3216, P2_U3215, P2_U3152,
         P2_U3151, P2_U3966;
  wire   n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10448, n10449, n10450, n10451, n10452, n10453, n10454,
         n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462,
         n10463, n10464, n10465, n10466, n10467, n10468, n10469, n10470,
         n10471, n10472, n10473, n10474, n10475, n10476, n10477, n10478,
         n10479, n10480, n10481, n10482, n10483, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10494,
         n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
         n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510,
         n10511, n10512, n10513, n10514, n10515, n10516, n10517, n10518,
         n10519, n10520, n10521, n10522, n10523, n10524, n10525, n10526,
         n10527, n10528, n10529, n10530, n10531, n10532, n10533, n10534,
         n10535, n10536, n10537, n10538, n10539, n10540, n10541, n10542,
         n10543, n10544, n10545, n10546, n10547, n10548, n10549, n10550,
         n10551, n10552, n10553, n10554, n10555, n10556, n10557, n10558,
         n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
         n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
         n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582,
         n10583, n10584, n10585, n10586, n10587, n10588, n10589, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10601, n10602, n10603, n10604, n10605, n10606,
         n10607, n10608, n10609, n10610, n10611, n10612, n10613, n10614,
         n10615, n10616, n10617, n10618, n10619, n10620, n10621, n10622,
         n10623, n10624, n10625, n10626, n10627, n10628, n10629, n10630,
         n10631, n10632, n10633, n10634, n10635, n10636, n10637, n10638,
         n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
         n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654,
         n10655, n10656, n10657, n10658, n10659, n10660, n10661, n10662,
         n10663, n10664, n10665, n10666, n10667, n10668, n10669, n10670,
         n10671, n10672, n10673, n10674, n10675, n10676, n10677, n10678,
         n10679, n10680, n10681, n10682, n10683, n10684, n10685, n10686,
         n10687, n10688, n10689, n10690, n10691, n10692, n10693, n10694,
         n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
         n10703, n10704;

  INV_X4 U4919 ( .A(P2_STATE_REG_SCAN_IN), .ZN(P2_U3152) );
  NAND2_X1 U4920 ( .A1(n8276), .A2(n8275), .ZN(n8291) );
  AND2_X1 U4921 ( .A1(n8134), .A2(n8133), .ZN(n9885) );
  CLKBUF_X2 U4923 ( .A(n6362), .Z(n4860) );
  XNOR2_X1 U4924 ( .A(n6444), .B(P1_IR_REG_30__SCAN_IN), .ZN(n6470) );
  NAND2_X1 U4925 ( .A1(n6597), .A2(P1_U3084), .ZN(n10039) );
  INV_X2 U4926 ( .A(n5557), .ZN(n6597) );
  INV_X2 U4927 ( .A(n8686), .ZN(n6773) );
  INV_X1 U4928 ( .A(n6115), .ZN(n5615) );
  NOR2_X1 U4929 ( .A1(n5492), .A2(n5612), .ZN(n5510) );
  AND2_X1 U4930 ( .A1(n6471), .A2(n6470), .ZN(n7140) );
  INV_X1 U4931 ( .A(n6643), .ZN(n6433) );
  INV_X1 U4934 ( .A(n6792), .ZN(n7439) );
  NAND2_X1 U4935 ( .A1(n9777), .A2(n9779), .ZN(n9761) );
  INV_X1 U4936 ( .A(n6896), .ZN(n6897) );
  NAND2_X1 U4937 ( .A1(n5296), .A2(n5295), .ZN(n5557) );
  AND4_X1 U4938 ( .A1(n6634), .A2(n6633), .A3(n6632), .A4(n6631), .ZN(n6797)
         );
  INV_X1 U4939 ( .A(n6447), .ZN(n6448) );
  INV_X2 U4940 ( .A(n6597), .ZN(n8387) );
  AOI211_X1 U4941 ( .C1(n9911), .C2(n9902), .A(n8347), .B(n8346), .ZN(n8348)
         );
  NOR2_X4 U4943 ( .A1(n7590), .A2(n7587), .ZN(n7698) );
  NAND2_X1 U4944 ( .A1(n5296), .A2(n5295), .ZN(n4854) );
  INV_X1 U4945 ( .A(n5965), .ZN(n5945) );
  XNOR2_X1 U4946 ( .A(n6247), .B(n6246), .ZN(n6578) );
  OR3_X4 U4947 ( .A1(n6394), .A2(n7808), .A3(n7964), .ZN(n6581) );
  XNOR2_X2 U4948 ( .A(n6448), .B(n4986), .ZN(n10041) );
  AND2_X4 U4950 ( .A1(n10037), .A2(n6471), .ZN(n6774) );
  BUF_X4 U4951 ( .A(n7140), .Z(n4856) );
  OR2_X1 U4952 ( .A1(n6182), .A2(n6178), .ZN(n6187) );
  AND2_X1 U4953 ( .A1(n9398), .A2(n5119), .ZN(n5118) );
  NAND2_X1 U4954 ( .A1(n5307), .A2(n4890), .ZN(n8987) );
  AND2_X1 U4955 ( .A1(n9716), .A2(n5362), .ZN(n8334) );
  AND2_X1 U4956 ( .A1(n5440), .A2(n8872), .ZN(n9171) );
  AND2_X1 U4957 ( .A1(n5213), .A2(n9397), .ZN(n5119) );
  OR2_X1 U4958 ( .A1(n9184), .A2(n9178), .ZN(n5440) );
  OR2_X1 U4959 ( .A1(n9396), .A2(n10693), .ZN(n5213) );
  NOR2_X1 U4960 ( .A1(n9119), .A2(n9151), .ZN(n9118) );
  NAND2_X1 U4961 ( .A1(n4980), .A2(n4869), .ZN(n9728) );
  NAND2_X1 U4962 ( .A1(n9208), .A2(n9207), .ZN(n9206) );
  NAND2_X1 U4963 ( .A1(n4977), .A2(n5318), .ZN(n6040) );
  NAND2_X1 U4964 ( .A1(n5960), .A2(n4975), .ZN(n4974) );
  NAND2_X1 U4965 ( .A1(n5394), .A2(n5392), .ZN(n8066) );
  NAND2_X1 U4966 ( .A1(n8047), .A2(n8506), .ZN(n8280) );
  NAND2_X1 U4967 ( .A1(n4951), .A2(n4949), .ZN(n8315) );
  NAND2_X1 U4968 ( .A1(n7717), .A2(n7716), .ZN(n7756) );
  AND2_X1 U4969 ( .A1(n7710), .A2(n7709), .ZN(n7714) );
  NAND2_X1 U4970 ( .A1(n8144), .A2(n8143), .ZN(n9873) );
  NAND2_X1 U4971 ( .A1(n7508), .A2(n5232), .ZN(n7596) );
  NAND2_X1 U4972 ( .A1(n7205), .A2(n7204), .ZN(n7508) );
  NAND2_X1 U4973 ( .A1(n7860), .A2(n7859), .ZN(n9993) );
  AND2_X1 U4974 ( .A1(n7166), .A2(n7165), .ZN(n7168) );
  INV_X2 U4975 ( .A(n9378), .ZN(n9268) );
  NAND2_X1 U4976 ( .A1(n7514), .A2(n7513), .ZN(n7640) );
  NAND2_X1 U4977 ( .A1(n5358), .A2(n5356), .ZN(n6927) );
  AND2_X1 U4978 ( .A1(n6586), .A2(n6585), .ZN(n6590) );
  INV_X2 U4979 ( .A(n8683), .ZN(n8675) );
  INV_X1 U4980 ( .A(n6259), .ZN(n5157) );
  NAND2_X1 U4981 ( .A1(n5190), .A2(n10512), .ZN(n7056) );
  CLKBUF_X1 U4982 ( .A(n6773), .Z(n8672) );
  BUF_X4 U4983 ( .A(n6780), .Z(n8678) );
  NAND3_X1 U4984 ( .A1(n5595), .A2(n5594), .A3(n5159), .ZN(n6259) );
  AND2_X2 U4985 ( .A1(n6773), .A2(n6580), .ZN(n6799) );
  NAND3_X1 U4986 ( .A1(n6796), .A2(n6795), .A3(n6794), .ZN(n8301) );
  INV_X1 U4987 ( .A(n9628), .ZN(n4989) );
  INV_X1 U4988 ( .A(n8685), .ZN(n6780) );
  NAND4_X1 U4990 ( .A1(n6808), .A2(n6807), .A3(n6806), .A4(n6805), .ZN(n9628)
         );
  OR2_X2 U4991 ( .A1(n6608), .A2(n6582), .ZN(n8685) );
  NAND4_X1 U4992 ( .A1(n6474), .A2(n6472), .A3(n6475), .A4(n6473), .ZN(n9631)
         );
  AND2_X2 U4993 ( .A1(n6279), .A2(n5522), .ZN(n6115) );
  OAI21_X1 U4994 ( .B1(n6603), .B2(P1_IR_REG_0__SCAN_IN), .A(n6469), .ZN(n6989) );
  INV_X4 U4995 ( .A(n8268), .ZN(n6775) );
  XNOR2_X1 U4996 ( .A(n5513), .B(n5493), .ZN(n8926) );
  INV_X1 U4997 ( .A(n6470), .ZN(n10037) );
  XNOR2_X1 U4998 ( .A(n6225), .B(n6224), .ZN(n6394) );
  XNOR2_X1 U4999 ( .A(n6480), .B(P1_IR_REG_19__SCAN_IN), .ZN(n9772) );
  XNOR2_X1 U5000 ( .A(n5516), .B(n5515), .ZN(n8928) );
  OAI21_X1 U5001 ( .B1(n5517), .B2(P2_IR_REG_21__SCAN_IN), .A(
        P2_IR_REG_31__SCAN_IN), .ZN(n6158) );
  NAND2_X1 U5002 ( .A1(n6240), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6477) );
  INV_X2 U5003 ( .A(n7786), .ZN(n4857) );
  CLKBUF_X3 U5004 ( .A(n5510), .Z(n4859) );
  AND2_X1 U5005 ( .A1(n5046), .A2(n6237), .ZN(n5375) );
  AND2_X1 U5006 ( .A1(n6250), .A2(n5373), .ZN(n5372) );
  AND2_X1 U5007 ( .A1(n6226), .A2(n5374), .ZN(n5373) );
  AND2_X1 U5008 ( .A1(n6228), .A2(n6224), .ZN(n6250) );
  NOR2_X1 U5009 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_IR_REG_1__SCAN_IN), .ZN(
        n5566) );
  NOR2_X1 U5010 ( .A1(P2_IR_REG_3__SCAN_IN), .A2(P2_IR_REG_2__SCAN_IN), .ZN(
        n5422) );
  INV_X1 U5011 ( .A(P1_IR_REG_17__SCAN_IN), .ZN(n6357) );
  INV_X1 U5012 ( .A(P1_IR_REG_16__SCAN_IN), .ZN(n6354) );
  NOR2_X1 U5013 ( .A1(P1_IR_REG_13__SCAN_IN), .A2(P1_IR_REG_10__SCAN_IN), .ZN(
        n6214) );
  INV_X1 U5014 ( .A(P2_IR_REG_21__SCAN_IN), .ZN(n5515) );
  INV_X1 U5015 ( .A(P2_IR_REG_22__SCAN_IN), .ZN(n6157) );
  INV_X1 U5016 ( .A(P2_IR_REG_17__SCAN_IN), .ZN(n5512) );
  INV_X1 U5017 ( .A(P2_IR_REG_9__SCAN_IN), .ZN(n5785) );
  NOR2_X1 U5018 ( .A1(P1_IR_REG_1__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6317) );
  NOR3_X1 U5019 ( .A1(P2_IR_REG_12__SCAN_IN), .A2(P2_IR_REG_13__SCAN_IN), .A3(
        P2_IR_REG_8__SCAN_IN), .ZN(n5490) );
  NOR2_X1 U5020 ( .A1(P1_IR_REG_5__SCAN_IN), .A2(P1_IR_REG_4__SCAN_IN), .ZN(
        n6219) );
  NAND2_X1 U5021 ( .A1(n6603), .A2(n8387), .ZN(n4858) );
  AOI211_X2 U5022 ( .C1(n10578), .C2(n9920), .A(n9919), .B(n9918), .ZN(n9921)
         );
  XNOR2_X2 U5023 ( .A(n5497), .B(n5496), .ZN(n6646) );
  NAND2_X2 U5024 ( .A1(n6242), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6247) );
  NAND2_X2 U5025 ( .A1(n6363), .A2(n4860), .ZN(n6603) );
  XNOR2_X2 U5026 ( .A(n5122), .B(n5526), .ZN(n6188) );
  INV_X1 U5027 ( .A(n10041), .ZN(n6471) );
  NAND2_X1 U5028 ( .A1(n8354), .A2(n8353), .ZN(n8382) );
  NAND2_X1 U5029 ( .A1(n8350), .A2(n8349), .ZN(n8354) );
  INV_X1 U5030 ( .A(P1_IR_REG_14__SCAN_IN), .ZN(n6216) );
  XNOR2_X1 U5031 ( .A(n5981), .B(n10062), .ZN(n5982) );
  AOI21_X1 U5032 ( .B1(n5274), .B2(n5276), .A(n4939), .ZN(n5273) );
  INV_X1 U5033 ( .A(n5926), .ZN(n5274) );
  OR3_X1 U5034 ( .A1(n6640), .A2(n6204), .A3(n6203), .ZN(n6265) );
  OAI21_X1 U5035 ( .B1(n9190), .B2(n9142), .A(n9141), .ZN(n9177) );
  INV_X1 U5036 ( .A(n5475), .ZN(n8270) );
  OR2_X1 U5037 ( .A1(n8553), .A2(n10376), .ZN(n9881) );
  NAND2_X1 U5038 ( .A1(n10029), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6444) );
  OR2_X1 U5039 ( .A1(n8553), .A2(n6363), .ZN(n9879) );
  NAND2_X1 U5040 ( .A1(n5039), .A2(n5038), .ZN(n8538) );
  NOR2_X1 U5041 ( .A1(n9708), .A2(n8532), .ZN(n5038) );
  NOR2_X1 U5042 ( .A1(n9411), .A2(n8991), .ZN(n8861) );
  NOR2_X1 U5043 ( .A1(n5443), .A2(n5146), .ZN(n5145) );
  INV_X1 U5044 ( .A(n8845), .ZN(n5146) );
  INV_X1 U5045 ( .A(n8614), .ZN(n5383) );
  OR2_X1 U5046 ( .A1(n9923), .A2(n8667), .ZN(n8454) );
  INV_X1 U5047 ( .A(n5807), .ZN(n4970) );
  INV_X1 U5048 ( .A(SI_10_), .ZN(n10191) );
  INV_X1 U5049 ( .A(SI_9_), .ZN(n10203) );
  OAI21_X1 U5050 ( .B1(n4854), .B2(P1_DATAO_REG_3__SCAN_IN), .A(n4962), .ZN(
        n5583) );
  NAND2_X1 U5051 ( .A1(n5557), .A2(n4963), .ZN(n4962) );
  AOI21_X1 U5052 ( .B1(n4873), .B2(n5432), .A(n4905), .ZN(n5431) );
  OR2_X1 U5053 ( .A1(n9111), .A2(n8715), .ZN(n8882) );
  OR2_X1 U5054 ( .A1(n9420), .A2(n9138), .ZN(n8856) );
  NAND2_X1 U5055 ( .A1(n5106), .A2(n5107), .ZN(n5101) );
  NOR2_X1 U5056 ( .A1(n5466), .A2(n5099), .ZN(n5104) );
  INV_X1 U5057 ( .A(n5106), .ZN(n5099) );
  OR2_X1 U5058 ( .A1(n9441), .A2(n9274), .ZN(n8840) );
  NOR2_X1 U5059 ( .A1(n9451), .A2(n5208), .ZN(n5207) );
  INV_X1 U5060 ( .A(n5209), .ZN(n5208) );
  OR2_X1 U5061 ( .A1(n9457), .A2(n9338), .ZN(n8833) );
  INV_X1 U5062 ( .A(n8799), .ZN(n5153) );
  NAND2_X1 U5063 ( .A1(n9067), .A2(n10521), .ZN(n8755) );
  NOR2_X1 U5064 ( .A1(n6165), .A2(n10051), .ZN(n6951) );
  NAND2_X1 U5065 ( .A1(n4917), .A2(n5511), .ZN(n5329) );
  NAND2_X1 U5066 ( .A1(n7452), .A2(n7451), .ZN(n7461) );
  NOR2_X1 U5067 ( .A1(n4880), .A2(n5393), .ZN(n5392) );
  INV_X1 U5068 ( .A(n7954), .ZN(n5393) );
  AND2_X1 U5069 ( .A1(n8291), .A2(n9721), .ZN(n8453) );
  INV_X1 U5070 ( .A(n8542), .ZN(n8587) );
  NAND2_X1 U5071 ( .A1(n4994), .A2(n4893), .ZN(n4993) );
  AND2_X1 U5072 ( .A1(n8469), .A2(n8470), .ZN(n9859) );
  AND2_X1 U5073 ( .A1(n8482), .A2(n7727), .ZN(n4985) );
  NAND2_X1 U5074 ( .A1(n8324), .A2(n8323), .ZN(n8350) );
  OAI21_X1 U5075 ( .B1(n6091), .B2(n6090), .A(n6089), .ZN(n6108) );
  NOR2_X1 U5076 ( .A1(n5047), .A2(n6314), .ZN(n5046) );
  NAND2_X1 U5077 ( .A1(n5249), .A2(n5250), .ZN(n5894) );
  AOI21_X1 U5078 ( .B1(n5251), .B2(n5258), .A(n4904), .ZN(n5250) );
  XNOR2_X1 U5079 ( .A(n5804), .B(SI_12_), .ZN(n5807) );
  INV_X1 U5080 ( .A(n5761), .ZN(n5282) );
  XNOR2_X1 U5081 ( .A(n5734), .B(n10203), .ZN(n5732) );
  OAI22_X2 U5082 ( .A1(n5715), .A2(n5714), .B1(SI_8_), .B2(n5713), .ZN(n5733)
         );
  XNOR2_X1 U5083 ( .A(n5713), .B(SI_8_), .ZN(n5714) );
  AOI21_X1 U5084 ( .B1(n5321), .B2(n5320), .A(n5319), .ZN(n5318) );
  NAND2_X1 U5085 ( .A1(n4974), .A2(n4972), .ZN(n4977) );
  INV_X1 U5086 ( .A(n6023), .ZN(n5319) );
  NOR2_X1 U5087 ( .A1(n4868), .A2(n8923), .ZN(n5429) );
  AND4_X1 U5088 ( .A1(n5867), .A2(n5866), .A3(n5865), .A4(n5864), .ZN(n7982)
         );
  AND2_X1 U5089 ( .A1(n10409), .A2(n6171), .ZN(n6640) );
  INV_X1 U5090 ( .A(P2_IR_REG_4__SCAN_IN), .ZN(n5491) );
  AOI21_X1 U5091 ( .B1(n5097), .B2(n9183), .A(n4908), .ZN(n5095) );
  OR2_X1 U5092 ( .A1(n9405), .A2(n9053), .ZN(n8872) );
  NAND2_X1 U5093 ( .A1(n5164), .A2(n8869), .ZN(n9184) );
  NAND2_X1 U5094 ( .A1(n9206), .A2(n5448), .ZN(n5164) );
  AND2_X1 U5095 ( .A1(n9197), .A2(n8712), .ZN(n5448) );
  AOI21_X1 U5096 ( .B1(n4867), .B2(n5089), .A(n4912), .ZN(n5087) );
  AND2_X1 U5097 ( .A1(n9441), .A2(n9131), .ZN(n9132) );
  INV_X2 U5098 ( .A(n5609), .ZN(n8726) );
  NOR2_X1 U5099 ( .A1(n9457), .A2(n9124), .ZN(n5209) );
  AOI21_X1 U5100 ( .B1(n4861), .B2(n8830), .A(n4937), .ZN(n5458) );
  AND2_X1 U5101 ( .A1(n9124), .A2(n9123), .ZN(n9125) );
  OR2_X1 U5102 ( .A1(n5203), .A2(n7914), .ZN(n5483) );
  NAND2_X1 U5103 ( .A1(n8773), .A2(n8772), .ZN(n8768) );
  XNOR2_X1 U5104 ( .A(n5525), .B(P2_IR_REG_30__SCAN_IN), .ZN(n5531) );
  NAND2_X1 U5105 ( .A1(n9485), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5525) );
  XNOR2_X1 U5106 ( .A(n5528), .B(P2_IR_REG_29__SCAN_IN), .ZN(n5530) );
  NAND2_X1 U5107 ( .A1(n5527), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5528) );
  AND2_X1 U5108 ( .A1(n4886), .A2(n5526), .ZN(n5473) );
  INV_X1 U5109 ( .A(P2_IR_REG_27__SCAN_IN), .ZN(n5496) );
  NOR2_X1 U5110 ( .A1(n8670), .A2(n8671), .ZN(n5418) );
  AOI21_X1 U5111 ( .B1(n9495), .B2(n9498), .A(n9497), .ZN(n9554) );
  NAND2_X1 U5112 ( .A1(n8394), .A2(n5242), .ZN(n5241) );
  NOR2_X1 U5113 ( .A1(n8598), .A2(n4855), .ZN(n5242) );
  AND2_X1 U5114 ( .A1(n7070), .A2(P1_REG3_REG_28__SCAN_IN), .ZN(n8331) );
  NAND2_X1 U5115 ( .A1(n5217), .A2(n5216), .ZN(n9777) );
  AOI21_X1 U5116 ( .B1(n5218), .B2(n5220), .A(n4897), .ZN(n5216) );
  NAND2_X1 U5117 ( .A1(n5196), .A2(n5195), .ZN(n8056) );
  INV_X1 U5118 ( .A(n9986), .ZN(n5195) );
  NAND2_X1 U5119 ( .A1(n5230), .A2(n5228), .ZN(n8041) );
  NOR2_X1 U5120 ( .A1(n8500), .A2(n5229), .ZN(n5228) );
  INV_X1 U5121 ( .A(n8005), .ZN(n5229) );
  INV_X2 U5122 ( .A(n8136), .ZN(n8153) );
  INV_X1 U5123 ( .A(n9879), .ZN(n10622) );
  INV_X1 U5124 ( .A(n10597), .ZN(n10617) );
  OR2_X1 U5125 ( .A1(n6394), .A2(n6396), .ZN(n10046) );
  OAI21_X1 U5126 ( .B1(n5927), .B2(n5275), .A(n5273), .ZN(n5983) );
  NAND2_X1 U5127 ( .A1(n5927), .A2(n5926), .ZN(n5944) );
  NAND2_X1 U5128 ( .A1(n5253), .A2(n5255), .ZN(n5873) );
  OAI21_X1 U5129 ( .B1(n5632), .B2(n5248), .A(n5654), .ZN(n5247) );
  NAND2_X1 U5130 ( .A1(n5629), .A2(SI_5_), .ZN(n5649) );
  AND4_X1 U5131 ( .A1(n8239), .A2(n8238), .A3(n8237), .A4(n8236), .ZN(n9768)
         );
  INV_X1 U5132 ( .A(n8290), .ZN(n5355) );
  NOR2_X1 U5133 ( .A1(n8334), .A2(n5361), .ZN(n8285) );
  AOI21_X1 U5134 ( .B1(n9716), .B2(n8534), .A(n8277), .ZN(n5361) );
  INV_X1 U5135 ( .A(n8330), .ZN(n8329) );
  NAND2_X1 U5136 ( .A1(n9730), .A2(n9729), .ZN(n9927) );
  NOR2_X1 U5137 ( .A1(n5014), .A2(n5015), .ZN(n5010) );
  INV_X1 U5138 ( .A(n8416), .ZN(n5015) );
  NAND2_X1 U5139 ( .A1(n5006), .A2(n5010), .ZN(n5005) );
  NAND2_X1 U5140 ( .A1(n8356), .A2(n8472), .ZN(n5007) );
  AOI21_X1 U5141 ( .B1(n5010), .B2(n5009), .A(n8533), .ZN(n5008) );
  INV_X1 U5142 ( .A(n4881), .ZN(n5009) );
  NAND2_X1 U5143 ( .A1(n5012), .A2(n8407), .ZN(n5004) );
  OAI211_X1 U5144 ( .C1(n8787), .C2(n5053), .A(n5051), .B(n5049), .ZN(n8797)
         );
  INV_X1 U5145 ( .A(n8829), .ZN(n5061) );
  NAND2_X1 U5146 ( .A1(n5064), .A2(n5063), .ZN(n5062) );
  NOR2_X1 U5147 ( .A1(n8827), .A2(n8828), .ZN(n5063) );
  OAI21_X1 U5148 ( .B1(n5069), .B2(n5068), .A(n5065), .ZN(n5064) );
  OAI21_X1 U5149 ( .B1(n8854), .B2(n8853), .A(n9230), .ZN(n8857) );
  NAND2_X1 U5150 ( .A1(n8529), .A2(n8528), .ZN(n5042) );
  NAND2_X1 U5151 ( .A1(n5079), .A2(n5076), .ZN(n5075) );
  AOI21_X1 U5152 ( .B1(n8880), .B2(n8881), .A(n5077), .ZN(n5076) );
  NAND2_X1 U5153 ( .A1(n8876), .A2(n8824), .ZN(n5079) );
  NOR3_X1 U5154 ( .A1(n8886), .A2(n8885), .A3(n8887), .ZN(n5074) );
  MUX2_X1 U5155 ( .A(n8884), .B(n8883), .S(n8890), .Z(n8885) );
  NAND2_X1 U5156 ( .A1(n5442), .A2(n9262), .ZN(n5441) );
  NAND2_X1 U5157 ( .A1(n8543), .A2(n8541), .ZN(n5031) );
  NOR2_X1 U5158 ( .A1(n8540), .A2(n8547), .ZN(n5267) );
  NAND2_X1 U5159 ( .A1(n8543), .A2(n8544), .ZN(n5033) );
  NOR2_X1 U5160 ( .A1(n8542), .A2(n8533), .ZN(n5266) );
  NAND2_X1 U5161 ( .A1(n8545), .A2(n9694), .ZN(n5265) );
  AND2_X1 U5162 ( .A1(n8327), .A2(n8694), .ZN(n8542) );
  AND2_X1 U5163 ( .A1(n8216), .A2(P1_REG3_REG_25__SCAN_IN), .ZN(n8230) );
  INV_X1 U5164 ( .A(n8453), .ZN(n8401) );
  OR2_X1 U5165 ( .A1(n8291), .A2(n9721), .ZN(n8447) );
  NOR2_X1 U5166 ( .A1(n5322), .A2(n4973), .ZN(n4972) );
  INV_X1 U5167 ( .A(n5304), .ZN(n5303) );
  OAI21_X1 U5168 ( .B1(n6102), .B2(n5305), .A(n8936), .ZN(n5304) );
  INV_X1 U5169 ( .A(n6106), .ZN(n5305) );
  INV_X1 U5170 ( .A(n5433), .ZN(n5432) );
  OAI21_X1 U5171 ( .B1(n8889), .B2(n9317), .A(n8931), .ZN(n5433) );
  OR2_X1 U5172 ( .A1(n9400), .A2(n9146), .ZN(n8877) );
  NAND2_X1 U5173 ( .A1(n8712), .A2(n8862), .ZN(n9140) );
  NOR2_X1 U5174 ( .A1(n9229), .A2(n5463), .ZN(n5462) );
  INV_X1 U5175 ( .A(n5476), .ZN(n5463) );
  OR2_X1 U5176 ( .A1(n9436), .A2(n9293), .ZN(n8845) );
  AOI21_X1 U5177 ( .B1(n5465), .B2(n9130), .A(n4901), .ZN(n5464) );
  INV_X1 U5178 ( .A(n9132), .ZN(n5467) );
  AOI21_X1 U5179 ( .B1(n5108), .B2(n9328), .A(n4909), .ZN(n5106) );
  INV_X1 U5180 ( .A(n5108), .ZN(n5107) );
  OR2_X1 U5181 ( .A1(n9448), .A2(n9339), .ZN(n8739) );
  INV_X1 U5182 ( .A(n5133), .ZN(n5130) );
  OR2_X1 U5183 ( .A1(n7985), .A2(n9060), .ZN(n8823) );
  AOI21_X1 U5184 ( .B1(n5471), .B2(n8915), .A(n4907), .ZN(n5469) );
  OR2_X1 U5185 ( .A1(n5843), .A2(n5842), .ZN(n5862) );
  NOR2_X1 U5186 ( .A1(n7618), .A2(n5454), .ZN(n5083) );
  NAND2_X1 U5187 ( .A1(n5121), .A2(n5120), .ZN(n8796) );
  INV_X1 U5188 ( .A(n8772), .ZN(n5124) );
  NAND2_X1 U5189 ( .A1(n8753), .A2(n7319), .ZN(n5447) );
  OR2_X1 U5190 ( .A1(n9068), .A2(n10505), .ZN(n8753) );
  NAND2_X1 U5191 ( .A1(n9223), .A2(n9226), .ZN(n9212) );
  AND2_X1 U5192 ( .A1(n7069), .A2(P1_REG3_REG_24__SCAN_IN), .ZN(n8216) );
  NOR2_X1 U5193 ( .A1(n9561), .A2(n5399), .ZN(n5398) );
  INV_X1 U5194 ( .A(n8632), .ZN(n5399) );
  NOR2_X1 U5195 ( .A1(n9516), .A2(n5176), .ZN(n5175) );
  INV_X1 U5196 ( .A(n9576), .ZN(n5176) );
  NOR2_X1 U5197 ( .A1(n4866), .A2(n5169), .ZN(n5168) );
  INV_X1 U5198 ( .A(n5398), .ZN(n5169) );
  INV_X1 U5199 ( .A(n6799), .ZN(n7033) );
  OR2_X1 U5200 ( .A1(n9928), .A2(n9768), .ZN(n8458) );
  NOR2_X1 U5201 ( .A1(n5344), .A2(n9779), .ZN(n5343) );
  NOR2_X1 U5202 ( .A1(n8283), .A2(n9798), .ZN(n5344) );
  INV_X1 U5203 ( .A(n5219), .ZN(n5218) );
  OAI21_X1 U5204 ( .B1(n8191), .B2(n5220), .A(n8207), .ZN(n5219) );
  AND2_X1 U5205 ( .A1(n8521), .A2(n8522), .ZN(n8520) );
  NOR2_X1 U5206 ( .A1(n9950), .A2(n9944), .ZN(n5185) );
  NAND2_X1 U5207 ( .A1(n4920), .A2(n4870), .ZN(n4994) );
  AND2_X1 U5208 ( .A1(n5235), .A2(n4920), .ZN(n4995) );
  AND2_X1 U5209 ( .A1(n8375), .A2(n8141), .ZN(n5235) );
  OAI21_X1 U5210 ( .B1(n8280), .B2(n5370), .A(n5368), .ZN(n9857) );
  INV_X1 U5211 ( .A(n5369), .ZN(n5368) );
  INV_X1 U5212 ( .A(n8512), .ZN(n5370) );
  AND2_X1 U5213 ( .A1(n9878), .A2(n8507), .ZN(n5371) );
  NOR2_X1 U5214 ( .A1(n9532), .A2(n8056), .ZN(n5194) );
  OR2_X1 U5215 ( .A1(n9532), .A2(n9880), .ZN(n8507) );
  OR2_X1 U5216 ( .A1(n9986), .A2(n9538), .ZN(n8502) );
  AND2_X1 U5217 ( .A1(n7946), .A2(n7855), .ZN(n8495) );
  AND2_X1 U5218 ( .A1(n7509), .A2(n7507), .ZN(n5232) );
  NOR2_X1 U5219 ( .A1(n5359), .A2(n5360), .ZN(n5357) );
  INV_X1 U5220 ( .A(n6902), .ZN(n5360) );
  XNOR2_X1 U5221 ( .A(n6925), .B(n9629), .ZN(n8358) );
  NAND2_X1 U5222 ( .A1(n8564), .A2(n8560), .ZN(n5231) );
  NOR2_X1 U5223 ( .A1(n9873), .A2(n9892), .ZN(n9868) );
  NAND2_X1 U5224 ( .A1(n6140), .A2(n6139), .ZN(n8320) );
  NAND2_X1 U5225 ( .A1(n6136), .A2(n6135), .ZN(n6140) );
  NOR2_X1 U5226 ( .A1(n5293), .A2(n5289), .ZN(n5288) );
  INV_X1 U5227 ( .A(n6006), .ZN(n5289) );
  NAND2_X1 U5228 ( .A1(n5294), .A2(n6044), .ZN(n5293) );
  INV_X1 U5229 ( .A(n6027), .ZN(n5294) );
  INV_X1 U5230 ( .A(n6026), .ZN(n5292) );
  INV_X1 U5231 ( .A(n5982), .ZN(n5271) );
  INV_X1 U5232 ( .A(P1_IR_REG_19__SCAN_IN), .ZN(n6239) );
  INV_X1 U5233 ( .A(n5943), .ZN(n5277) );
  NAND2_X1 U5234 ( .A1(n5830), .A2(SI_14_), .ZN(n5853) );
  NAND2_X1 U5235 ( .A1(n4964), .A2(n4967), .ZN(n5829) );
  NAND2_X1 U5236 ( .A1(n5733), .A2(n4968), .ZN(n4964) );
  XNOR2_X1 U5237 ( .A(n5826), .B(n5809), .ZN(n5828) );
  INV_X1 U5238 ( .A(SI_13_), .ZN(n5809) );
  NAND2_X1 U5239 ( .A1(n5760), .A2(SI_11_), .ZN(n5782) );
  NAND2_X1 U5240 ( .A1(n6235), .A2(n5405), .ZN(n5404) );
  INV_X1 U5241 ( .A(P1_IR_REG_7__SCAN_IN), .ZN(n5405) );
  INV_X1 U5242 ( .A(SI_7_), .ZN(n10210) );
  INV_X1 U5243 ( .A(n5583), .ZN(n5581) );
  NAND2_X1 U5244 ( .A1(n5585), .A2(n5584), .ZN(n5602) );
  INV_X1 U5245 ( .A(P2_ADDR_REG_19__SCAN_IN), .ZN(n5297) );
  AND2_X1 U5246 ( .A1(n4976), .A2(n8959), .ZN(n4975) );
  INV_X1 U5247 ( .A(n9025), .ZN(n4976) );
  NAND2_X1 U5248 ( .A1(n9000), .A2(n8999), .ZN(n5307) );
  NAND2_X1 U5249 ( .A1(n7160), .A2(n5695), .ZN(n5317) );
  OR2_X1 U5250 ( .A1(n6951), .A2(n6170), .ZN(n6201) );
  NAND2_X1 U5251 ( .A1(n8981), .A2(n8980), .ZN(n5324) );
  AND2_X1 U5252 ( .A1(n5623), .A2(n7420), .ZN(n5309) );
  INV_X1 U5253 ( .A(n5626), .ZN(n5312) );
  AND2_X1 U5254 ( .A1(n4948), .A2(n4888), .ZN(n5326) );
  NAND2_X1 U5255 ( .A1(n7907), .A2(n5849), .ZN(n4950) );
  OR2_X1 U5256 ( .A1(n10289), .A2(n10290), .ZN(n7897) );
  AND2_X1 U5257 ( .A1(n6101), .A2(n6100), .ZN(n8991) );
  AND4_X1 U5258 ( .A1(n5746), .A2(n5745), .A3(n5744), .A4(n5743), .ZN(n9014)
         );
  NAND2_X1 U5259 ( .A1(n5589), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n5534) );
  NOR2_X1 U5260 ( .A1(n5612), .A2(P2_IR_REG_5__SCAN_IN), .ZN(n5678) );
  NOR2_X1 U5261 ( .A1(n9212), .A2(n9417), .ZN(n9211) );
  NAND2_X1 U5262 ( .A1(n9211), .A2(n9196), .ZN(n9191) );
  AND2_X1 U5263 ( .A1(n8866), .A2(n8869), .ZN(n9197) );
  NAND2_X1 U5264 ( .A1(n5141), .A2(n5139), .ZN(n9208) );
  AOI21_X1 U5265 ( .B1(n5142), .B2(n5144), .A(n5140), .ZN(n5139) );
  INV_X1 U5266 ( .A(n8856), .ZN(n5140) );
  INV_X1 U5267 ( .A(n9140), .ZN(n9207) );
  OR2_X1 U5268 ( .A1(n9250), .A2(n9264), .ZN(n5476) );
  OR2_X1 U5269 ( .A1(n9430), .A2(n9275), .ZN(n8852) );
  NAND2_X1 U5270 ( .A1(n5105), .A2(n5106), .ZN(n9304) );
  OR2_X1 U5271 ( .A1(n9327), .A2(n5107), .ZN(n5105) );
  INV_X1 U5272 ( .A(P2_IR_REG_19__SCAN_IN), .ZN(n5518) );
  INV_X1 U5273 ( .A(n5329), .ZN(n5327) );
  NOR2_X1 U5274 ( .A1(n5482), .A2(n9320), .ZN(n5108) );
  INV_X1 U5275 ( .A(n9125), .ZN(n5460) );
  NAND2_X1 U5276 ( .A1(n5459), .A2(n5060), .ZN(n5461) );
  INV_X1 U5277 ( .A(n8088), .ZN(n5459) );
  INV_X1 U5278 ( .A(n8742), .ZN(n5138) );
  INV_X1 U5279 ( .A(n8084), .ZN(n5132) );
  AOI21_X1 U5280 ( .B1(n5137), .B2(n5135), .A(n5134), .ZN(n5133) );
  INV_X1 U5281 ( .A(n8745), .ZN(n5135) );
  INV_X1 U5282 ( .A(n8743), .ZN(n5134) );
  INV_X1 U5283 ( .A(n5461), .ZN(n9126) );
  NOR2_X1 U5284 ( .A1(n7985), .A2(n5201), .ZN(n5200) );
  INV_X1 U5285 ( .A(n5202), .ZN(n5201) );
  NOR2_X1 U5286 ( .A1(n8821), .A2(n5472), .ZN(n5471) );
  INV_X1 U5287 ( .A(n5483), .ZN(n5472) );
  NOR2_X1 U5288 ( .A1(n7842), .A2(n7841), .ZN(n7844) );
  AND4_X1 U5289 ( .A1(n5797), .A2(n5796), .A3(n5795), .A4(n5794), .ZN(n8804)
         );
  NAND2_X1 U5290 ( .A1(n7698), .A2(n4883), .ZN(n7836) );
  NAND2_X1 U5291 ( .A1(n5151), .A2(n5152), .ZN(n5148) );
  INV_X1 U5292 ( .A(n8794), .ZN(n5444) );
  OR2_X1 U5293 ( .A1(n6435), .A2(n6188), .ZN(n9371) );
  AND2_X1 U5294 ( .A1(n8768), .A2(n6271), .ZN(n5456) );
  INV_X1 U5295 ( .A(n8768), .ZN(n8903) );
  AND2_X1 U5296 ( .A1(n6269), .A2(n6268), .ZN(n9365) );
  NAND2_X1 U5297 ( .A1(n5425), .A2(n9068), .ZN(n6268) );
  NAND2_X1 U5298 ( .A1(n7352), .A2(n5423), .ZN(n6269) );
  NAND2_X1 U5299 ( .A1(n5424), .A2(n10505), .ZN(n5423) );
  AND2_X1 U5300 ( .A1(n6952), .A2(n7313), .ZN(n7352) );
  AND2_X1 U5301 ( .A1(n8895), .A2(n6256), .ZN(n9376) );
  OR2_X1 U5302 ( .A1(n6951), .A2(n6267), .ZN(n7296) );
  NAND2_X1 U5303 ( .A1(n7844), .A2(n7843), .ZN(n10678) );
  OR2_X1 U5304 ( .A1(n7025), .A2(n5609), .ZN(n5639) );
  AND3_X1 U5305 ( .A1(n5571), .A2(n5570), .A3(n5569), .ZN(n10521) );
  NAND2_X1 U5306 ( .A1(n6159), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6173) );
  OR2_X1 U5307 ( .A1(n6640), .A2(n6174), .ZN(n10050) );
  INV_X1 U5308 ( .A(P2_IR_REG_28__SCAN_IN), .ZN(n5526) );
  AND2_X1 U5309 ( .A1(n4886), .A2(n5451), .ZN(n5080) );
  NAND2_X1 U5310 ( .A1(n5385), .A2(n5388), .ZN(n8110) );
  INV_X1 U5311 ( .A(n5389), .ZN(n5388) );
  OAI21_X1 U5312 ( .B1(n5392), .B2(n5390), .A(n8071), .ZN(n5389) );
  AND2_X1 U5313 ( .A1(n7030), .A2(n7023), .ZN(n5421) );
  AND2_X1 U5314 ( .A1(n6584), .A2(n6583), .ZN(n6585) );
  NAND2_X1 U5315 ( .A1(n6799), .A2(n9631), .ZN(n6586) );
  NAND2_X1 U5316 ( .A1(n6780), .A2(n9631), .ZN(n6589) );
  INV_X1 U5317 ( .A(n9507), .ZN(n5401) );
  NAND2_X1 U5318 ( .A1(n7942), .A2(n7941), .ZN(n5394) );
  OR2_X1 U5319 ( .A1(n7740), .A2(n7739), .ZN(n7862) );
  AOI21_X1 U5320 ( .B1(n5401), .B2(n5398), .A(n5396), .ZN(n5395) );
  INV_X1 U5321 ( .A(n9562), .ZN(n5396) );
  INV_X1 U5322 ( .A(n9516), .ZN(n5172) );
  NAND2_X1 U5323 ( .A1(n7755), .A2(n7754), .ZN(n5377) );
  NAND2_X1 U5324 ( .A1(n5379), .A2(n5378), .ZN(n9588) );
  AOI21_X1 U5325 ( .B1(n4865), .B2(n5382), .A(n4931), .ZN(n5378) );
  NAND2_X1 U5326 ( .A1(n7032), .A2(n7031), .ZN(n7126) );
  INV_X1 U5327 ( .A(n8659), .ZN(n5181) );
  AND2_X1 U5328 ( .A1(n4878), .A2(n9555), .ZN(n5180) );
  NOR2_X1 U5329 ( .A1(n8452), .A2(n5237), .ZN(n5036) );
  INV_X1 U5330 ( .A(n8553), .ZN(n5237) );
  NAND2_X1 U5331 ( .A1(n5263), .A2(n8547), .ZN(n5262) );
  AND4_X1 U5332 ( .A1(n7043), .A2(n7042), .A3(n7041), .A4(n7040), .ZN(n7167)
         );
  NOR2_X1 U5333 ( .A1(n7429), .A2(n7428), .ZN(n7427) );
  AND2_X1 U5334 ( .A1(n9733), .A2(n5197), .ZN(n9703) );
  NOR2_X1 U5335 ( .A1(n8327), .A2(n5198), .ZN(n5197) );
  INV_X1 U5336 ( .A(n5199), .ZN(n5198) );
  AND2_X1 U5337 ( .A1(n7073), .A2(n7072), .ZN(n8691) );
  OR2_X1 U5338 ( .A1(n9920), .A2(n9726), .ZN(n8534) );
  INV_X1 U5339 ( .A(n9708), .ZN(n9717) );
  NAND2_X1 U5340 ( .A1(n8534), .A2(n8535), .ZN(n9708) );
  NAND2_X1 U5341 ( .A1(n9761), .A2(n8242), .ZN(n4980) );
  NAND2_X1 U5342 ( .A1(n5341), .A2(n8522), .ZN(n5340) );
  INV_X1 U5343 ( .A(n5343), .ZN(n5341) );
  NAND2_X1 U5344 ( .A1(n8462), .A2(n8522), .ZN(n5342) );
  OAI21_X1 U5345 ( .B1(n9799), .B2(n8283), .A(n5343), .ZN(n5345) );
  INV_X1 U5346 ( .A(n8520), .ZN(n9779) );
  AND2_X1 U5347 ( .A1(n8461), .A2(n8462), .ZN(n9798) );
  OAI21_X1 U5348 ( .B1(n9823), .B2(n8282), .A(n8281), .ZN(n9808) );
  INV_X1 U5349 ( .A(n4996), .ZN(n9806) );
  OAI21_X1 U5350 ( .B1(n9883), .B2(n4993), .A(n4991), .ZN(n4996) );
  INV_X1 U5351 ( .A(n4992), .ZN(n4991) );
  OAI22_X1 U5352 ( .A1(n4995), .A2(n4993), .B1(n9954), .B2(n9810), .ZN(n4992)
         );
  NAND2_X1 U5353 ( .A1(n9806), .A2(n8191), .ZN(n9805) );
  NAND2_X1 U5354 ( .A1(n5194), .A2(n5193), .ZN(n9892) );
  NAND2_X1 U5355 ( .A1(n8014), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8147) );
  AND2_X1 U5356 ( .A1(n8502), .A2(n8503), .ZN(n8500) );
  AOI21_X1 U5357 ( .B1(n5233), .B2(n4984), .A(n4903), .ZN(n4983) );
  INV_X1 U5358 ( .A(n4985), .ZN(n4984) );
  NOR2_X1 U5359 ( .A1(n5366), .A2(n5365), .ZN(n5364) );
  INV_X1 U5360 ( .A(n8479), .ZN(n5366) );
  INV_X1 U5361 ( .A(n8474), .ZN(n5365) );
  OR2_X1 U5362 ( .A1(n7523), .A2(n7522), .ZN(n7655) );
  AND2_X1 U5363 ( .A1(n8416), .A2(n8411), .ZN(n8367) );
  NAND2_X1 U5364 ( .A1(n4915), .A2(n5020), .ZN(n7173) );
  NAND2_X1 U5365 ( .A1(n6927), .A2(n5021), .ZN(n5020) );
  NOR2_X1 U5366 ( .A1(n5023), .A2(n5022), .ZN(n5021) );
  INV_X1 U5367 ( .A(n9881), .ZN(n10623) );
  AND2_X1 U5368 ( .A1(n7028), .A2(n7027), .ZN(n7111) );
  NAND2_X1 U5369 ( .A1(n5024), .A2(n4988), .ZN(n7114) );
  NAND2_X1 U5370 ( .A1(n6927), .A2(n8565), .ZN(n5024) );
  NAND2_X1 U5371 ( .A1(n5475), .A2(P1_REG0_REG_2__SCAN_IN), .ZN(n6634) );
  NAND2_X1 U5372 ( .A1(n6775), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6632) );
  AND2_X1 U5373 ( .A1(n6906), .A2(n6905), .ZN(n10626) );
  INV_X1 U5374 ( .A(n5231), .ZN(n8359) );
  AND2_X1 U5375 ( .A1(n9631), .A2(n6983), .ZN(n6987) );
  NAND2_X1 U5376 ( .A1(n8360), .A2(n6991), .ZN(n6990) );
  NOR2_X1 U5377 ( .A1(n8277), .A2(n5223), .ZN(n5222) );
  INV_X1 U5378 ( .A(n5225), .ZN(n5223) );
  INV_X1 U5379 ( .A(n9694), .ZN(n9906) );
  NAND2_X1 U5380 ( .A1(n7653), .A2(n7652), .ZN(n10003) );
  OR2_X1 U5381 ( .A1(n7650), .A2(n6792), .ZN(n7653) );
  NAND2_X1 U5382 ( .A1(n5192), .A2(n6370), .ZN(n5191) );
  OR2_X1 U5383 ( .A1(n8136), .A2(n6598), .ZN(n6601) );
  XNOR2_X1 U5384 ( .A(n8391), .B(n8390), .ZN(n8727) );
  NAND2_X1 U5385 ( .A1(n8386), .A2(n8385), .ZN(n8391) );
  XNOR2_X1 U5386 ( .A(n8382), .B(n8381), .ZN(n8718) );
  AND2_X1 U5387 ( .A1(n5375), .A2(n4928), .ZN(n6446) );
  INV_X1 U5388 ( .A(P1_IR_REG_28__SCAN_IN), .ZN(n5221) );
  NAND2_X1 U5389 ( .A1(n5375), .A2(n5373), .ZN(n6249) );
  INV_X1 U5390 ( .A(n6052), .ZN(n6050) );
  XNOR2_X1 U5391 ( .A(n6477), .B(P1_IR_REG_20__SCAN_IN), .ZN(n8595) );
  NAND2_X1 U5392 ( .A1(n5944), .A2(n5943), .ZN(n5964) );
  OAI211_X1 U5393 ( .C1(n5733), .C2(n4966), .A(n4965), .B(n5828), .ZN(n5260)
         );
  NAND2_X1 U5394 ( .A1(n4969), .A2(n4967), .ZN(n4965) );
  INV_X1 U5395 ( .A(n4967), .ZN(n4966) );
  OAI21_X1 U5396 ( .B1(n5733), .B2(n5281), .A(n5278), .ZN(n5808) );
  OAI21_X1 U5397 ( .B1(n5760), .B2(SI_11_), .A(n5782), .ZN(n5761) );
  NAND2_X1 U5398 ( .A1(n5733), .A2(n5285), .ZN(n5283) );
  NAND2_X1 U5399 ( .A1(n4863), .A2(n4894), .ZN(n5284) );
  INV_X1 U5400 ( .A(n5649), .ZN(n5248) );
  AND2_X1 U5401 ( .A1(n5669), .A2(n5653), .ZN(n5654) );
  AND2_X1 U5402 ( .A1(n5649), .A2(n5631), .ZN(n5632) );
  NAND2_X1 U5403 ( .A1(n5633), .A2(n5632), .ZN(n5650) );
  AND2_X1 U5404 ( .A1(n5627), .A2(n5605), .ZN(n5606) );
  NAND2_X1 U5405 ( .A1(n5503), .A2(n5504), .ZN(n4982) );
  INV_X1 U5406 ( .A(n5553), .ZN(n4981) );
  NAND2_X1 U5407 ( .A1(n6114), .A2(n6113), .ZN(n9405) );
  AND4_X1 U5408 ( .A1(n5821), .A2(n5820), .A3(n5819), .A4(n5818), .ZN(n7914)
         );
  AND4_X1 U5409 ( .A1(n5620), .A2(n5619), .A3(n5618), .A4(n5617), .ZN(n7217)
         );
  AOI21_X1 U5410 ( .B1(n4956), .B2(n4959), .A(n4955), .ZN(n4954) );
  NAND2_X1 U5411 ( .A1(n4974), .A2(n4971), .ZN(n8981) );
  INV_X1 U5412 ( .A(n4973), .ZN(n4971) );
  NAND2_X1 U5413 ( .A1(n5908), .A2(n5907), .ZN(n9457) );
  OR2_X1 U5414 ( .A1(n8135), .A2(n5609), .ZN(n5908) );
  NAND2_X1 U5415 ( .A1(n7224), .A2(n5623), .ZN(n7419) );
  NAND2_X1 U5416 ( .A1(n5967), .A2(n5966), .ZN(n9441) );
  NAND2_X1 U5417 ( .A1(n7357), .A2(n5547), .ZN(n7089) );
  NAND2_X1 U5418 ( .A1(n5932), .A2(n5931), .ZN(n9451) );
  OR2_X1 U5419 ( .A1(n8142), .A2(n5609), .ZN(n5932) );
  AND4_X1 U5420 ( .A1(n5885), .A2(n5884), .A3(n5883), .A4(n5882), .ZN(n9058)
         );
  NAND2_X1 U5421 ( .A1(n5860), .A2(n5859), .ZN(n8310) );
  NAND2_X1 U5422 ( .A1(n4900), .A2(n4862), .ZN(n5073) );
  INV_X1 U5423 ( .A(n7217), .ZN(n9066) );
  OAI211_X1 U5424 ( .C1(n9177), .C2(n5094), .A(n5091), .B(n5090), .ZN(n9394)
         );
  NAND2_X1 U5425 ( .A1(n5097), .A2(n9144), .ZN(n5094) );
  OAI21_X1 U5426 ( .B1(n5095), .B2(n9144), .A(n5092), .ZN(n5091) );
  NAND2_X1 U5427 ( .A1(n5769), .A2(n5768), .ZN(n7693) );
  OR2_X1 U5428 ( .A1(n10050), .A2(n6948), .ZN(n9316) );
  OAI21_X1 U5429 ( .B1(n6841), .B2(n5609), .A(n5614), .ZN(n7301) );
  INV_X1 U5430 ( .A(n10505), .ZN(n5425) );
  INV_X1 U5431 ( .A(n9316), .ZN(n9377) );
  INV_X1 U5432 ( .A(n9333), .ZN(n9366) );
  NAND2_X1 U5433 ( .A1(n7296), .A2(n9316), .ZN(n9378) );
  NOR2_X1 U5434 ( .A1(P2_IR_REG_25__SCAN_IN), .A2(P2_IR_REG_26__SCAN_IN), .ZN(
        n5450) );
  NAND2_X1 U5435 ( .A1(n5419), .A2(n5416), .ZN(n8700) );
  INV_X1 U5436 ( .A(n5418), .ZN(n5416) );
  AND2_X1 U5437 ( .A1(n8690), .A2(n5417), .ZN(n5410) );
  AND4_X1 U5438 ( .A1(n8206), .A2(n8205), .A3(n8204), .A4(n8203), .ZN(n9782)
         );
  AND4_X1 U5439 ( .A1(n8225), .A2(n8224), .A3(n8223), .A4(n8222), .ZN(n9783)
         );
  AND4_X1 U5440 ( .A1(n6702), .A2(n6701), .A3(n6700), .A4(n6699), .ZN(n9766)
         );
  NAND2_X1 U5441 ( .A1(n8246), .A2(n8245), .ZN(n9923) );
  INV_X1 U5442 ( .A(n8667), .ZN(n9755) );
  INV_X1 U5443 ( .A(n7167), .ZN(n9625) );
  NAND2_X1 U5444 ( .A1(n5475), .A2(P1_REG0_REG_1__SCAN_IN), .ZN(n6481) );
  NAND2_X1 U5445 ( .A1(n6775), .A2(P1_REG2_REG_1__SCAN_IN), .ZN(n6482) );
  AOI21_X1 U5446 ( .B1(n8345), .B2(n9891), .A(n8344), .ZN(n9913) );
  INV_X1 U5447 ( .A(n8343), .ZN(n8344) );
  AOI22_X1 U5448 ( .A1(n8342), .A2(n10622), .B1(n9696), .B2(n9611), .ZN(n8343)
         );
  AND2_X1 U5449 ( .A1(n5000), .A2(n4999), .ZN(n9926) );
  AOI21_X1 U5450 ( .B1(n9732), .B2(n9891), .A(n9731), .ZN(n4999) );
  NAND2_X1 U5451 ( .A1(n5001), .A2(n10629), .ZN(n5000) );
  OR2_X1 U5452 ( .A1(n7857), .A2(n6792), .ZN(n7860) );
  NAND2_X1 U5453 ( .A1(n9841), .A2(n4942), .ZN(n9898) );
  NAND2_X1 U5454 ( .A1(n8294), .A2(n10629), .ZN(n5352) );
  NAND2_X1 U5455 ( .A1(n10637), .A2(n10632), .ZN(n5351) );
  NAND2_X1 U5456 ( .A1(n10635), .A2(P1_REG0_REG_28__SCAN_IN), .ZN(n5354) );
  AND2_X1 U5457 ( .A1(n9916), .A2(n5355), .ZN(n5353) );
  AND2_X1 U5458 ( .A1(n6398), .A2(n6397), .ZN(n6920) );
  AND2_X1 U5459 ( .A1(n6402), .A2(n6401), .ZN(n6743) );
  INV_X1 U5460 ( .A(n5158), .ZN(n8767) );
  NAND2_X1 U5461 ( .A1(n8786), .A2(n5050), .ZN(n5049) );
  NOR2_X1 U5462 ( .A1(n5053), .A2(n5054), .ZN(n5050) );
  INV_X1 U5463 ( .A(n8782), .ZN(n5054) );
  INV_X1 U5464 ( .A(n5052), .ZN(n5051) );
  NAND2_X1 U5465 ( .A1(n8782), .A2(n8783), .ZN(n5048) );
  OAI211_X1 U5466 ( .C1(n5013), .C2(n5017), .A(n5004), .B(n8533), .ZN(n5003)
         );
  NOR2_X1 U5467 ( .A1(n8816), .A2(n8817), .ZN(n5069) );
  NOR2_X1 U5468 ( .A1(n5067), .A2(n5066), .ZN(n5065) );
  INV_X1 U5469 ( .A(n8820), .ZN(n5066) );
  NAND2_X1 U5470 ( .A1(n8815), .A2(n8915), .ZN(n5068) );
  NAND2_X1 U5471 ( .A1(n5062), .A2(n5059), .ZN(n8831) );
  NOR2_X1 U5472 ( .A1(n5061), .A2(n5060), .ZN(n5059) );
  INV_X1 U5473 ( .A(n8846), .ZN(n5057) );
  NAND2_X1 U5474 ( .A1(n5025), .A2(n4884), .ZN(n8516) );
  NAND2_X1 U5475 ( .A1(n5026), .A2(n4896), .ZN(n5025) );
  NAND2_X1 U5476 ( .A1(n5055), .A2(n9245), .ZN(n8854) );
  NAND2_X1 U5477 ( .A1(n5058), .A2(n5056), .ZN(n5055) );
  NOR2_X1 U5478 ( .A1(n5057), .A2(n9262), .ZN(n5056) );
  NAND2_X1 U5479 ( .A1(n8843), .A2(n4891), .ZN(n5058) );
  OAI21_X1 U5480 ( .B1(n8865), .B2(n9140), .A(n8864), .ZN(n8871) );
  MUX2_X1 U5481 ( .A(n8859), .B(n8858), .S(n8890), .Z(n8865) );
  NAND2_X1 U5482 ( .A1(n5041), .A2(n5040), .ZN(n5039) );
  NOR2_X1 U5483 ( .A1(n8531), .A2(n8530), .ZN(n5040) );
  NAND2_X1 U5484 ( .A1(n5042), .A2(n9753), .ZN(n5041) );
  NAND2_X1 U5485 ( .A1(n5078), .A2(n8879), .ZN(n5077) );
  AND2_X1 U5486 ( .A1(n5770), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n5791) );
  AND2_X1 U5487 ( .A1(n7693), .A2(n7694), .ZN(n8809) );
  OR2_X1 U5488 ( .A1(n9993), .A2(n8126), .ZN(n8496) );
  AND2_X1 U5489 ( .A1(n8032), .A2(n9620), .ZN(n8493) );
  INV_X1 U5490 ( .A(n8410), .ZN(n5018) );
  INV_X1 U5491 ( .A(P1_IR_REG_11__SCAN_IN), .ZN(n6212) );
  INV_X1 U5492 ( .A(P1_IR_REG_15__SCAN_IN), .ZN(n6213) );
  INV_X1 U5493 ( .A(P1_IR_REG_18__SCAN_IN), .ZN(n6215) );
  INV_X1 U5494 ( .A(n5255), .ZN(n5252) );
  OAI211_X1 U5495 ( .C1(n5557), .C2(P1_DATAO_REG_0__SCAN_IN), .A(SI_0_), .B(
        n4979), .ZN(n5502) );
  NAND2_X1 U5496 ( .A1(n4854), .A2(n6467), .ZN(n4979) );
  INV_X1 U5497 ( .A(P1_RD_REG_SCAN_IN), .ZN(n5084) );
  AND2_X1 U5498 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(P2_REG3_REG_4__SCAN_IN), 
        .ZN(n5640) );
  NOR2_X1 U5499 ( .A1(n6010), .A2(n10264), .ZN(n6031) );
  INV_X1 U5500 ( .A(n8980), .ZN(n5320) );
  AND2_X1 U5501 ( .A1(n6031), .A2(P2_REG3_REG_23__SCAN_IN), .ZN(n6056) );
  INV_X1 U5502 ( .A(n9031), .ZN(n5323) );
  NOR2_X1 U5503 ( .A1(n7994), .A2(n4961), .ZN(n4960) );
  INV_X1 U5504 ( .A(n5890), .ZN(n4961) );
  OAI21_X1 U5505 ( .B1(n8894), .B2(n8893), .A(n5481), .ZN(n8927) );
  OR2_X1 U5506 ( .A1(n8892), .A2(n8891), .ZN(n5481) );
  AND2_X1 U5507 ( .A1(n5075), .A2(n5074), .ZN(n8894) );
  OR2_X1 U5508 ( .A1(n5462), .A2(n5089), .ZN(n5088) );
  INV_X1 U5509 ( .A(n9139), .ZN(n5089) );
  AND2_X1 U5510 ( .A1(n4922), .A2(n5143), .ZN(n5142) );
  NAND2_X1 U5511 ( .A1(n5145), .A2(n9280), .ZN(n5143) );
  INV_X1 U5512 ( .A(n5145), .ZN(n5144) );
  OR2_X1 U5513 ( .A1(n8709), .A2(n9264), .ZN(n8848) );
  OR2_X1 U5514 ( .A1(n9451), .A2(n9129), .ZN(n8708) );
  OR2_X1 U5515 ( .A1(n9124), .A2(n9058), .ZN(n8742) );
  OR2_X1 U5516 ( .A1(n8310), .A2(n7982), .ZN(n8744) );
  INV_X1 U5517 ( .A(n7841), .ZN(n5113) );
  NOR2_X1 U5518 ( .A1(n8805), .A2(n7840), .ZN(n7841) );
  AND2_X1 U5519 ( .A1(n4883), .A2(n5203), .ZN(n5202) );
  NAND2_X1 U5520 ( .A1(n5791), .A2(P2_REG3_REG_12__SCAN_IN), .ZN(n5816) );
  INV_X1 U5521 ( .A(n7494), .ZN(n5455) );
  NAND2_X1 U5522 ( .A1(n5071), .A2(n6257), .ZN(n8760) );
  INV_X1 U5523 ( .A(n8928), .ZN(n8733) );
  AND2_X1 U5524 ( .A1(n8793), .A2(n8794), .ZN(n8908) );
  NAND2_X1 U5525 ( .A1(n5211), .A2(n10546), .ZN(n7332) );
  INV_X1 U5526 ( .A(n7406), .ZN(n5211) );
  OR2_X1 U5527 ( .A1(n5716), .A2(P2_IR_REG_8__SCAN_IN), .ZN(n5787) );
  OR2_X1 U5528 ( .A1(n5698), .A2(P2_IR_REG_7__SCAN_IN), .ZN(n5716) );
  NOR2_X1 U5529 ( .A1(n5390), .A2(n5387), .ZN(n5386) );
  INV_X1 U5530 ( .A(n7941), .ZN(n5387) );
  OR2_X1 U5531 ( .A1(n7455), .A2(n7454), .ZN(n7458) );
  XNOR2_X1 U5532 ( .A(n6615), .B(n8675), .ZN(n6618) );
  OR2_X1 U5533 ( .A1(n9545), .A2(n9544), .ZN(n8619) );
  OR2_X1 U5534 ( .A1(n5381), .A2(n8620), .ZN(n5380) );
  OR2_X1 U5535 ( .A1(n9535), .A2(n5383), .ZN(n5381) );
  OR2_X1 U5536 ( .A1(n8620), .A2(n5383), .ZN(n5382) );
  INV_X1 U5537 ( .A(n7021), .ZN(n7022) );
  INV_X1 U5538 ( .A(n8546), .ZN(n5263) );
  AND2_X1 U5539 ( .A1(n8546), .A2(n5265), .ZN(n5264) );
  NAND2_X1 U5540 ( .A1(n5033), .A2(n5266), .ZN(n5032) );
  NAND2_X1 U5541 ( .A1(n5031), .A2(n5267), .ZN(n5030) );
  NAND2_X1 U5542 ( .A1(n8333), .A2(n9612), .ZN(n8539) );
  NOR2_X1 U5543 ( .A1(n8291), .A2(n9920), .ZN(n5199) );
  NOR2_X1 U5544 ( .A1(n9939), .A2(n5184), .ZN(n5183) );
  INV_X1 U5545 ( .A(n5185), .ZN(n5184) );
  AND2_X1 U5546 ( .A1(n6694), .A2(P1_REG3_REG_23__SCAN_IN), .ZN(n7069) );
  INV_X1 U5547 ( .A(n8192), .ZN(n5220) );
  INV_X1 U5548 ( .A(n8496), .ZN(n5337) );
  AND2_X1 U5549 ( .A1(n8478), .A2(n8479), .ZN(n8476) );
  NAND2_X1 U5550 ( .A1(n5002), .A2(n8416), .ZN(n5012) );
  NAND2_X1 U5551 ( .A1(n8402), .A2(n4881), .ZN(n5017) );
  NOR2_X1 U5552 ( .A1(n7142), .A2(n7141), .ZN(n7188) );
  INV_X1 U5553 ( .A(n8565), .ZN(n5022) );
  NAND2_X1 U5554 ( .A1(n6990), .A2(n6902), .ZN(n8561) );
  NAND2_X1 U5555 ( .A1(n9829), .A2(n5183), .ZN(n9784) );
  NAND2_X1 U5556 ( .A1(n6112), .A2(n6111), .ZN(n6136) );
  AOI21_X1 U5557 ( .B1(n5259), .B2(n5257), .A(n5256), .ZN(n5255) );
  INV_X1 U5558 ( .A(n5853), .ZN(n5256) );
  INV_X1 U5559 ( .A(n5828), .ZN(n5257) );
  NAND2_X1 U5560 ( .A1(n5254), .A2(n5259), .ZN(n5253) );
  INV_X1 U5561 ( .A(n5829), .ZN(n5254) );
  AOI21_X1 U5562 ( .B1(n4914), .B2(n5278), .A(n4872), .ZN(n4967) );
  AOI21_X1 U5563 ( .B1(n5280), .B2(n5286), .A(n5279), .ZN(n5278) );
  INV_X1 U5564 ( .A(n5782), .ZN(n5279) );
  INV_X1 U5565 ( .A(P1_IR_REG_6__SCAN_IN), .ZN(n6235) );
  INV_X1 U5566 ( .A(SI_6_), .ZN(n10213) );
  INV_X1 U5567 ( .A(SI_4_), .ZN(n10215) );
  NOR2_X1 U5568 ( .A1(P1_IR_REG_3__SCAN_IN), .A2(P1_IR_REG_2__SCAN_IN), .ZN(
        n6319) );
  AND2_X1 U5569 ( .A1(n5081), .A2(n5601), .ZN(n5584) );
  OAI21_X1 U5570 ( .B1(n4854), .B2(n5556), .A(n5555), .ZN(n5559) );
  NAND2_X1 U5571 ( .A1(n5640), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n5685) );
  OR2_X1 U5572 ( .A1(n5720), .A2(n5719), .ZN(n5741) );
  INV_X1 U5573 ( .A(n8097), .ZN(n4955) );
  AOI21_X1 U5574 ( .B1(n5303), .B2(n5305), .A(n4936), .ZN(n5301) );
  OR2_X1 U5575 ( .A1(n7159), .A2(n7160), .ZN(n8968) );
  NOR2_X1 U5576 ( .A1(n5980), .A2(n5979), .ZN(n4973) );
  NAND2_X1 U5577 ( .A1(n5956), .A2(n5955), .ZN(n5960) );
  OR2_X1 U5578 ( .A1(n7571), .A2(n7572), .ZN(n7569) );
  OR2_X1 U5579 ( .A1(n5572), .A2(n7220), .ZN(n5576) );
  OR2_X1 U5580 ( .A1(n5912), .A2(n5911), .ZN(n5933) );
  AOI21_X1 U5581 ( .B1(n4960), .B2(n4958), .A(n4957), .ZN(n4956) );
  INV_X1 U5582 ( .A(n7995), .ZN(n4957) );
  INV_X1 U5583 ( .A(n4960), .ZN(n4959) );
  INV_X1 U5584 ( .A(n8989), .ZN(n5306) );
  XNOR2_X1 U5585 ( .A(n7985), .B(n6115), .ZN(n8311) );
  INV_X1 U5586 ( .A(n5431), .ZN(n5430) );
  NAND2_X1 U5587 ( .A1(n5431), .A2(n8923), .ZN(n5428) );
  NOR4_X1 U5588 ( .A1(n8924), .A2(n8923), .A3(n9144), .A4(n8922), .ZN(n8925)
         );
  AND2_X1 U5589 ( .A1(n6064), .A2(n6063), .ZN(n9138) );
  NAND2_X1 U5590 ( .A1(n5095), .A2(n5093), .ZN(n5092) );
  NAND2_X1 U5591 ( .A1(n5096), .A2(n5078), .ZN(n5093) );
  NAND2_X1 U5592 ( .A1(n8714), .A2(n8713), .ZN(n9111) );
  NAND2_X1 U5593 ( .A1(n5439), .A2(n5437), .ZN(n9145) );
  AOI21_X1 U5594 ( .B1(n4864), .B2(n9178), .A(n5438), .ZN(n5437) );
  NAND2_X1 U5595 ( .A1(n9185), .A2(n9241), .ZN(n5162) );
  AND2_X1 U5596 ( .A1(n6126), .A2(n6095), .ZN(n9194) );
  AND2_X1 U5597 ( .A1(n6080), .A2(n6079), .ZN(n9233) );
  NAND2_X1 U5598 ( .A1(n9261), .A2(n9255), .ZN(n9266) );
  NAND2_X1 U5599 ( .A1(n9277), .A2(n8845), .ZN(n9261) );
  INV_X1 U5600 ( .A(n5100), .ZN(n5102) );
  OAI21_X1 U5601 ( .B1(n5466), .B2(n5101), .A(n5464), .ZN(n5100) );
  OR2_X1 U5602 ( .A1(n5994), .A2(n5993), .ZN(n6010) );
  AND2_X1 U5603 ( .A1(n6017), .A2(n6016), .ZN(n9275) );
  AND2_X1 U5604 ( .A1(n5976), .A2(n5975), .ZN(n9274) );
  NAND2_X1 U5605 ( .A1(n9272), .A2(n9133), .ZN(n9277) );
  NAND2_X1 U5606 ( .A1(n8089), .A2(n5205), .ZN(n9312) );
  NOR2_X1 U5607 ( .A1(n9448), .A2(n5206), .ZN(n5205) );
  INV_X1 U5608 ( .A(n5207), .ZN(n5206) );
  AND3_X1 U5609 ( .A1(n5954), .A2(n5953), .A3(n5952), .ZN(n9339) );
  NAND2_X1 U5610 ( .A1(n5126), .A2(n5127), .ZN(n9335) );
  AOI21_X1 U5611 ( .B1(n5129), .B2(n5136), .A(n5128), .ZN(n5127) );
  INV_X1 U5612 ( .A(n8833), .ZN(n5128) );
  NAND2_X1 U5613 ( .A1(n8089), .A2(n9463), .ZN(n9351) );
  OAI21_X1 U5614 ( .B1(n8087), .B2(n8916), .A(n5114), .ZN(n8088) );
  OAI21_X1 U5615 ( .B1(n7842), .B2(n5112), .A(n5111), .ZN(n8087) );
  NAND2_X1 U5616 ( .A1(n5469), .A2(n5470), .ZN(n5111) );
  NAND2_X1 U5617 ( .A1(n5469), .A2(n5113), .ZN(n5112) );
  INV_X1 U5618 ( .A(n5471), .ZN(n5470) );
  AND4_X1 U5619 ( .A1(n5848), .A2(n5847), .A3(n5846), .A4(n5845), .ZN(n9060)
         );
  NOR2_X1 U5620 ( .A1(n8913), .A2(n8807), .ZN(n5149) );
  OR2_X1 U5621 ( .A1(n10659), .A2(n7694), .ZN(n5484) );
  AND2_X1 U5622 ( .A1(n8810), .A2(n8811), .ZN(n8801) );
  NAND2_X1 U5623 ( .A1(n8909), .A2(n5083), .ZN(n5082) );
  AND2_X1 U5624 ( .A1(n8806), .A2(n8747), .ZN(n8910) );
  NOR2_X1 U5625 ( .A1(n7614), .A2(n5156), .ZN(n5155) );
  INV_X1 U5626 ( .A(n8796), .ZN(n5156) );
  NAND2_X1 U5627 ( .A1(n7495), .A2(n8794), .ZN(n7580) );
  AND4_X1 U5628 ( .A1(n5708), .A2(n5707), .A3(n5706), .A4(n5705), .ZN(n7478)
         );
  INV_X1 U5629 ( .A(n8778), .ZN(n5125) );
  NAND2_X1 U5630 ( .A1(n8778), .A2(n5124), .ZN(n5123) );
  NAND2_X1 U5631 ( .A1(n7298), .A2(n10537), .ZN(n7406) );
  NAND2_X1 U5632 ( .A1(n8760), .A2(n8755), .ZN(n8754) );
  INV_X1 U5633 ( .A(n9370), .ZN(n9241) );
  INV_X1 U5634 ( .A(n9371), .ZN(n9239) );
  OR2_X1 U5635 ( .A1(n6435), .A2(n6673), .ZN(n9370) );
  NAND2_X1 U5636 ( .A1(n8729), .A2(n8728), .ZN(n9386) );
  NAND2_X1 U5637 ( .A1(n6142), .A2(n6141), .ZN(n9400) );
  NAND2_X1 U5638 ( .A1(n6093), .A2(n6092), .ZN(n9411) );
  OR2_X1 U5639 ( .A1(n8212), .A2(n5609), .ZN(n6055) );
  NAND2_X1 U5640 ( .A1(n6009), .A2(n6008), .ZN(n9430) );
  NAND2_X1 U5641 ( .A1(n5992), .A2(n5991), .ZN(n9436) );
  OR2_X1 U5642 ( .A1(n8179), .A2(n5609), .ZN(n5992) );
  INV_X1 U5643 ( .A(n9458), .ZN(n10691) );
  NOR2_X1 U5644 ( .A1(n5329), .A2(n5514), .ZN(n5328) );
  NAND2_X1 U5645 ( .A1(n5903), .A2(n5512), .ZN(n5929) );
  AND2_X1 U5646 ( .A1(n4859), .A2(n5511), .ZN(n5903) );
  INV_X1 U5647 ( .A(n5414), .ZN(n5413) );
  OAI21_X1 U5648 ( .B1(n5420), .B2(n5415), .A(n8681), .ZN(n5414) );
  INV_X1 U5649 ( .A(n9600), .ZN(n5420) );
  NAND2_X1 U5650 ( .A1(n9554), .A2(n9555), .ZN(n9553) );
  INV_X1 U5651 ( .A(n7561), .ZN(n5402) );
  NAND2_X1 U5652 ( .A1(n7557), .A2(n7556), .ZN(n5403) );
  OR2_X1 U5653 ( .A1(n5174), .A2(n4866), .ZN(n5167) );
  AND2_X1 U5654 ( .A1(n5395), .A2(n5175), .ZN(n5174) );
  NAND2_X1 U5655 ( .A1(n8066), .A2(n4892), .ZN(n8111) );
  NAND2_X1 U5656 ( .A1(n8122), .A2(n8124), .ZN(n8121) );
  AND4_X1 U5657 ( .A1(n8256), .A2(n8255), .A3(n8254), .A4(n8253), .ZN(n8667)
         );
  AND2_X1 U5658 ( .A1(n8178), .A2(n8177), .ZN(n9848) );
  NAND2_X1 U5659 ( .A1(n9640), .A2(n9641), .ZN(n9639) );
  NOR2_X1 U5660 ( .A1(n6561), .A2(n6560), .ZN(n6559) );
  NAND2_X1 U5661 ( .A1(n6341), .A2(n6815), .ZN(n6881) );
  NOR2_X1 U5662 ( .A1(n7270), .A2(n7269), .ZN(n7268) );
  OR2_X1 U5663 ( .A1(n6291), .A2(P1_IR_REG_14__SCAN_IN), .ZN(n6349) );
  NOR2_X1 U5664 ( .A1(n6352), .A2(n7777), .ZN(n9649) );
  AOI21_X1 U5665 ( .B1(n9672), .B2(P1_REG2_REG_17__SCAN_IN), .A(n9671), .ZN(
        n9674) );
  AOI21_X1 U5666 ( .B1(n8718), .B2(n7439), .A(n8355), .ZN(n9702) );
  NOR2_X1 U5667 ( .A1(n8536), .A2(n5363), .ZN(n5362) );
  INV_X1 U5668 ( .A(n8534), .ZN(n5363) );
  AND2_X1 U5669 ( .A1(n8266), .A2(n8265), .ZN(n9713) );
  AND2_X1 U5670 ( .A1(n8264), .A2(n8250), .ZN(n9734) );
  INV_X1 U5671 ( .A(n9927), .ZN(n5001) );
  AND2_X1 U5672 ( .A1(n8249), .A2(n8233), .ZN(n9748) );
  OR2_X1 U5673 ( .A1(n8241), .A2(n9762), .ZN(n9741) );
  NAND2_X1 U5674 ( .A1(n9829), .A2(n8641), .ZN(n9813) );
  AND2_X1 U5675 ( .A1(n8435), .A2(n8463), .ZN(n9809) );
  NAND2_X1 U5676 ( .A1(n4990), .A2(n4994), .ZN(n9821) );
  NAND2_X1 U5677 ( .A1(n9883), .A2(n4995), .ZN(n4990) );
  AND2_X1 U5678 ( .A1(n8467), .A2(n8468), .ZN(n9846) );
  AND2_X1 U5679 ( .A1(n8165), .A2(n8164), .ZN(n9861) );
  NAND2_X1 U5680 ( .A1(n9883), .A2(n8141), .ZN(n9854) );
  NAND2_X1 U5681 ( .A1(n9876), .A2(n8512), .ZN(n9858) );
  INV_X1 U5682 ( .A(n9878), .ZN(n9884) );
  AND2_X1 U5683 ( .A1(n8511), .A2(n8512), .ZN(n9878) );
  AND2_X1 U5684 ( .A1(n8280), .A2(n8507), .ZN(n9877) );
  NAND2_X1 U5685 ( .A1(n8280), .A2(n5371), .ZN(n9876) );
  AND3_X1 U5686 ( .A1(n8020), .A2(n8019), .A3(n8018), .ZN(n9880) );
  INV_X1 U5687 ( .A(n5194), .ZN(n9894) );
  NAND2_X1 U5688 ( .A1(n8044), .A2(n8043), .ZN(n9532) );
  INV_X1 U5689 ( .A(n8506), .ZN(n8374) );
  AND2_X1 U5690 ( .A1(n8052), .A2(n8051), .ZN(n9860) );
  AND2_X1 U5691 ( .A1(n8507), .A2(n8508), .ZN(n8506) );
  NAND2_X1 U5692 ( .A1(n7854), .A2(n7853), .ZN(n7946) );
  NAND2_X1 U5693 ( .A1(n7925), .A2(n8371), .ZN(n7924) );
  NAND2_X1 U5694 ( .A1(n7850), .A2(n7849), .ZN(n7923) );
  OR2_X1 U5695 ( .A1(n10616), .A2(n10003), .ZN(n7733) );
  NAND2_X1 U5696 ( .A1(n7728), .A2(n4985), .ZN(n7850) );
  INV_X1 U5697 ( .A(n8476), .ZN(n8369) );
  NAND2_X1 U5698 ( .A1(n5367), .A2(n8474), .ZN(n7748) );
  NAND2_X1 U5699 ( .A1(n5188), .A2(n5187), .ZN(n10616) );
  OR2_X1 U5700 ( .A1(n7464), .A2(n7463), .ZN(n7523) );
  INV_X1 U5701 ( .A(P1_REG3_REG_10__SCAN_IN), .ZN(n7522) );
  OR2_X1 U5702 ( .A1(n7640), .A2(n10621), .ZN(n7641) );
  NAND2_X1 U5703 ( .A1(n8402), .A2(n8410), .ZN(n7599) );
  NAND2_X1 U5704 ( .A1(n7508), .A2(n7507), .ZN(n7598) );
  AND4_X1 U5705 ( .A1(n7150), .A2(n7149), .A3(n7148), .A4(n7147), .ZN(n7519)
         );
  NAND2_X1 U5706 ( .A1(n4978), .A2(n5214), .ZN(n5480) );
  NAND2_X1 U5707 ( .A1(n4988), .A2(n7109), .ZN(n4978) );
  NAND2_X1 U5708 ( .A1(n6919), .A2(n8363), .ZN(n7110) );
  NAND2_X1 U5709 ( .A1(n6918), .A2(n6917), .ZN(n6919) );
  AND2_X1 U5710 ( .A1(n5028), .A2(n8358), .ZN(n5358) );
  NAND2_X1 U5711 ( .A1(n6990), .A2(n5357), .ZN(n5356) );
  NAND2_X1 U5712 ( .A1(n8560), .A2(n5231), .ZN(n5028) );
  OR2_X1 U5713 ( .A1(n6923), .A2(n6922), .ZN(n7208) );
  INV_X1 U5714 ( .A(n4855), .ZN(n6623) );
  OR2_X1 U5715 ( .A1(n9920), .A2(n9613), .ZN(n5225) );
  NOR2_X1 U5716 ( .A1(n9717), .A2(n5227), .ZN(n5226) );
  INV_X1 U5717 ( .A(n8258), .ZN(n5227) );
  NAND2_X1 U5718 ( .A1(n8196), .A2(n8195), .ZN(n9944) );
  OR2_X1 U5719 ( .A1(n6934), .A2(n8595), .ZN(n10597) );
  XNOR2_X1 U5720 ( .A(n8320), .B(n8319), .ZN(n8604) );
  NAND2_X1 U5721 ( .A1(n5043), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6253) );
  INV_X1 U5722 ( .A(n5047), .ZN(n5045) );
  XNOR2_X1 U5723 ( .A(n6136), .B(n6135), .ZN(n8259) );
  AOI21_X1 U5724 ( .B1(n6044), .B2(n5292), .A(n4933), .ZN(n5291) );
  INV_X1 U5725 ( .A(P1_IR_REG_24__SCAN_IN), .ZN(n6226) );
  NAND2_X1 U5726 ( .A1(n5276), .A2(n5982), .ZN(n5272) );
  INV_X1 U5727 ( .A(n5270), .ZN(n5269) );
  OAI21_X1 U5728 ( .B1(n5273), .B2(n5271), .A(n4938), .ZN(n5270) );
  INV_X1 U5729 ( .A(P1_IR_REG_21__SCAN_IN), .ZN(n6246) );
  AND2_X1 U5730 ( .A1(n5943), .A2(n5925), .ZN(n5926) );
  NAND2_X1 U5731 ( .A1(n5733), .A2(n5732), .ZN(n5759) );
  AND2_X1 U5732 ( .A1(n5696), .A2(n5673), .ZN(n5674) );
  AOI21_X1 U5733 ( .B1(n5246), .B2(n5248), .A(n5244), .ZN(n5243) );
  INV_X1 U5734 ( .A(n5669), .ZN(n5244) );
  NAND2_X1 U5735 ( .A1(n5044), .A2(n6235), .ZN(n6312) );
  NAND2_X1 U5736 ( .A1(n5563), .A2(n5564), .ZN(n5580) );
  NAND2_X1 U5737 ( .A1(n5302), .A2(n6106), .ZN(n8937) );
  NAND2_X1 U5738 ( .A1(n6103), .A2(n6102), .ZN(n5302) );
  XNOR2_X1 U5739 ( .A(n6040), .B(n6038), .ZN(n8945) );
  NAND2_X1 U5740 ( .A1(n5307), .A2(n6068), .ZN(n8990) );
  NAND2_X1 U5741 ( .A1(n6072), .A2(n6071), .ZN(n9417) );
  NAND2_X1 U5742 ( .A1(n5886), .A2(n7891), .ZN(n7896) );
  NAND2_X1 U5743 ( .A1(n7896), .A2(n5890), .ZN(n7998) );
  XNOR2_X1 U5744 ( .A(n6067), .B(n6065), .ZN(n9000) );
  AND2_X1 U5745 ( .A1(n6184), .A2(n6183), .ZN(n9009) );
  NAND2_X1 U5746 ( .A1(n5960), .A2(n8959), .ZN(n9024) );
  NAND2_X1 U5747 ( .A1(n6206), .A2(n6205), .ZN(n10284) );
  NAND2_X1 U5748 ( .A1(n5324), .A2(n6005), .ZN(n9032) );
  NAND2_X1 U5749 ( .A1(n5324), .A2(n5321), .ZN(n9034) );
  NAND2_X1 U5750 ( .A1(n7572), .A2(n5752), .ZN(n5315) );
  INV_X1 U5751 ( .A(n9015), .ZN(n10281) );
  NAND2_X1 U5752 ( .A1(n4953), .A2(n4956), .ZN(n8099) );
  OR2_X1 U5753 ( .A1(n5886), .A2(n4959), .ZN(n4953) );
  AOI21_X1 U5754 ( .B1(n5312), .B2(n7420), .A(n4911), .ZN(n5311) );
  INV_X1 U5755 ( .A(n7374), .ZN(n7330) );
  AOI21_X1 U5756 ( .B1(n7419), .B2(n5626), .A(n5313), .ZN(n5310) );
  AOI21_X1 U5757 ( .B1(n5326), .B2(n4950), .A(n4943), .ZN(n4949) );
  OR2_X1 U5758 ( .A1(n5325), .A2(n10289), .ZN(n4951) );
  INV_X1 U5759 ( .A(n5326), .ZN(n5325) );
  INV_X1 U5760 ( .A(n4950), .ZN(n5850) );
  INV_X1 U5761 ( .A(n9046), .ZN(n10293) );
  NAND2_X1 U5762 ( .A1(n6419), .A2(P2_REG0_REG_2__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U5763 ( .A1(n5589), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n5550) );
  AND2_X1 U5764 ( .A1(n5549), .A2(n5551), .ZN(n5070) );
  OR2_X1 U5765 ( .A1(n5548), .A2(n5529), .ZN(n5533) );
  NAND2_X1 U5766 ( .A1(n6640), .A2(n10413), .ZN(n9069) );
  AND2_X1 U5767 ( .A1(n5637), .A2(n5636), .ZN(n10462) );
  AND2_X1 U5768 ( .A1(n6647), .A2(n6646), .ZN(n10450) );
  INV_X1 U5769 ( .A(n9386), .ZN(n9115) );
  AOI21_X1 U5770 ( .B1(n8718), .B2(n8726), .A(n8717), .ZN(n9393) );
  NAND2_X1 U5771 ( .A1(n5440), .A2(n4864), .ZN(n9169) );
  NAND2_X1 U5772 ( .A1(n5098), .A2(n5097), .ZN(n9161) );
  AND2_X1 U5773 ( .A1(n5098), .A2(n4887), .ZN(n9160) );
  AOI21_X1 U5774 ( .B1(n5163), .B2(n9349), .A(n5160), .ZN(n9408) );
  NAND2_X1 U5775 ( .A1(n5162), .A2(n5161), .ZN(n5160) );
  XNOR2_X1 U5776 ( .A(n9184), .B(n9183), .ZN(n5163) );
  NAND2_X1 U5777 ( .A1(n9186), .A2(n9239), .ZN(n5161) );
  NAND2_X1 U5778 ( .A1(n9206), .A2(n8712), .ZN(n9199) );
  NAND2_X1 U5779 ( .A1(n9244), .A2(n5476), .ZN(n9222) );
  OR2_X1 U5780 ( .A1(n9246), .A2(n9245), .ZN(n9244) );
  NAND2_X1 U5781 ( .A1(n5468), .A2(n5465), .ZN(n9279) );
  AND2_X1 U5782 ( .A1(n5521), .A2(n5520), .ZN(n9317) );
  AND2_X1 U5783 ( .A1(n5109), .A2(n5110), .ZN(n9310) );
  NAND2_X1 U5784 ( .A1(n9327), .A2(n9336), .ZN(n5109) );
  NAND2_X1 U5785 ( .A1(n8089), .A2(n5209), .ZN(n9329) );
  NAND2_X1 U5786 ( .A1(n5461), .A2(n4861), .ZN(n9356) );
  NAND2_X1 U5787 ( .A1(n5132), .A2(n5137), .ZN(n5131) );
  NAND2_X1 U5788 ( .A1(n10678), .A2(n5483), .ZN(n7915) );
  NAND2_X1 U5789 ( .A1(n7698), .A2(n10659), .ZN(n7699) );
  AND2_X1 U5790 ( .A1(n7338), .A2(n8783), .ZN(n7480) );
  NAND2_X1 U5791 ( .A1(n7302), .A2(n8772), .ZN(n7403) );
  AND2_X1 U5792 ( .A1(n6965), .A2(n6271), .ZN(n7295) );
  NAND2_X1 U5793 ( .A1(n10521), .A2(n5212), .ZN(n10519) );
  INV_X1 U5794 ( .A(n9152), .ZN(n9380) );
  NAND2_X1 U5795 ( .A1(n9399), .A2(n5118), .ZN(n9470) );
  XNOR2_X1 U5796 ( .A(n6161), .B(P2_IR_REG_24__SCAN_IN), .ZN(n10409) );
  AND2_X1 U5797 ( .A1(n6432), .A2(P2_STATE_REG_SCAN_IN), .ZN(n10413) );
  NAND2_X1 U5798 ( .A1(n5524), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5122) );
  XNOR2_X1 U5799 ( .A(n6154), .B(P2_IR_REG_26__SCAN_IN), .ZN(n10408) );
  NAND2_X1 U5800 ( .A1(n5520), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5513) );
  INV_X1 U5801 ( .A(P1_DATAO_REG_15__SCAN_IN), .ZN(n6894) );
  NOR2_X1 U5802 ( .A1(n6597), .A2(P2_STATE_REG_SCAN_IN), .ZN(n9487) );
  AND4_X1 U5803 ( .A1(n7194), .A2(n7193), .A3(n7192), .A4(n7191), .ZN(n7562)
         );
  NAND2_X1 U5804 ( .A1(n7198), .A2(n7197), .ZN(n7520) );
  AND4_X1 U5805 ( .A1(n7662), .A2(n7661), .A3(n7660), .A4(n7659), .ZN(n7760)
         );
  OAI21_X1 U5806 ( .B1(n8299), .B2(n8298), .A(n6802), .ZN(n6840) );
  NAND2_X1 U5807 ( .A1(n9505), .A2(n9507), .ZN(n9506) );
  AND4_X1 U5808 ( .A1(n8289), .A2(n8288), .A3(n8287), .A4(n8286), .ZN(n8694)
         );
  OAI21_X1 U5809 ( .B1(n5413), .B2(n8690), .A(n5408), .ZN(n5407) );
  NAND2_X1 U5810 ( .A1(n5413), .A2(n5409), .ZN(n5408) );
  OR2_X1 U5811 ( .A1(n8690), .A2(n5417), .ZN(n5409) );
  NAND2_X1 U5812 ( .A1(n5413), .A2(n5412), .ZN(n5411) );
  INV_X1 U5813 ( .A(n8690), .ZN(n5412) );
  AND4_X1 U5814 ( .A1(n7747), .A2(n7746), .A3(n7745), .A4(n7744), .ZN(n7855)
         );
  NAND2_X1 U5815 ( .A1(n7732), .A2(n7731), .ZN(n9998) );
  NAND2_X1 U5816 ( .A1(n9553), .A2(n8659), .ZN(n9526) );
  NAND2_X1 U5817 ( .A1(n8229), .A2(n8228), .ZN(n9928) );
  INV_X1 U5818 ( .A(n9618), .ZN(n9538) );
  AND3_X1 U5819 ( .A1(n8151), .A2(n8150), .A3(n8149), .ZN(n9882) );
  OR2_X1 U5820 ( .A1(n8135), .A2(n4858), .ZN(n8140) );
  NAND2_X1 U5821 ( .A1(n6603), .A2(n10044), .ZN(n6469) );
  OR2_X1 U5822 ( .A1(n9589), .A2(n5401), .ZN(n5397) );
  OR2_X1 U5823 ( .A1(n9585), .A2(n5401), .ZN(n5400) );
  NAND2_X1 U5824 ( .A1(n8170), .A2(n8169), .ZN(n9954) );
  INV_X1 U5825 ( .A(n7946), .ZN(n8032) );
  AND4_X1 U5826 ( .A1(n7670), .A2(n7669), .A3(n7668), .A4(n7667), .ZN(n7959)
         );
  NOR2_X1 U5827 ( .A1(n5391), .A2(n4880), .ZN(n7953) );
  INV_X1 U5828 ( .A(n5394), .ZN(n5391) );
  AND2_X1 U5829 ( .A1(n8190), .A2(n8189), .ZN(n9581) );
  NAND2_X1 U5830 ( .A1(n5170), .A2(n9515), .ZN(n9575) );
  NAND2_X1 U5831 ( .A1(n5177), .A2(n5171), .ZN(n5170) );
  AND2_X1 U5832 ( .A1(n5395), .A2(n5172), .ZN(n5171) );
  AND4_X1 U5833 ( .A1(n7529), .A2(n7528), .A3(n7527), .A4(n7526), .ZN(n7767)
         );
  INV_X1 U5834 ( .A(n7763), .ZN(n5376) );
  INV_X1 U5835 ( .A(n9609), .ZN(n9590) );
  INV_X1 U5836 ( .A(n9569), .ZN(n9601) );
  INV_X1 U5837 ( .A(n7137), .ZN(n5384) );
  NAND2_X1 U5838 ( .A1(n5179), .A2(n5178), .ZN(n9599) );
  NAND2_X1 U5839 ( .A1(n4940), .A2(n4878), .ZN(n5178) );
  NAND2_X1 U5840 ( .A1(n6624), .A2(n9866), .ZN(n9607) );
  NAND2_X1 U5841 ( .A1(n6629), .A2(n6622), .ZN(n9609) );
  INV_X1 U5842 ( .A(n5239), .ZN(n5238) );
  NOR2_X1 U5843 ( .A1(n5036), .A2(n6904), .ZN(n5035) );
  OR2_X1 U5844 ( .A1(n5486), .A2(n8595), .ZN(n5236) );
  INV_X1 U5845 ( .A(n9726), .ZN(n9613) );
  INV_X1 U5846 ( .A(n9782), .ZN(n9811) );
  INV_X1 U5847 ( .A(n9848), .ZN(n9810) );
  INV_X1 U5848 ( .A(n9861), .ZN(n9824) );
  INV_X1 U5849 ( .A(n7855), .ZN(n9620) );
  INV_X1 U5850 ( .A(n7959), .ZN(n9621) );
  INV_X1 U5851 ( .A(n7519), .ZN(n9624) );
  NAND2_X1 U5852 ( .A1(n6775), .A2(P1_REG2_REG_0__SCAN_IN), .ZN(n6472) );
  OR2_X1 U5853 ( .A1(n6568), .A2(n6567), .ZN(n6565) );
  NOR2_X1 U5854 ( .A1(n7103), .A2(n7102), .ZN(n7101) );
  XNOR2_X1 U5855 ( .A(n6892), .B(n6351), .ZN(n7779) );
  AOI21_X1 U5856 ( .B1(n9655), .B2(P1_REG2_REG_16__SCAN_IN), .A(n9647), .ZN(
        n6365) );
  OR2_X1 U5857 ( .A1(n10374), .A2(n6363), .ZN(n9673) );
  NAND2_X1 U5858 ( .A1(n8393), .A2(n8392), .ZN(n9694) );
  NAND2_X1 U5859 ( .A1(n9730), .A2(n8258), .ZN(n9709) );
  OR2_X1 U5860 ( .A1(n8212), .A2(n6792), .ZN(n8215) );
  OAI21_X1 U5861 ( .B1(n9799), .B2(n5342), .A(n5340), .ZN(n9765) );
  AOI21_X1 U5862 ( .B1(n9799), .B2(n9798), .A(n8283), .ZN(n9780) );
  NAND2_X1 U5863 ( .A1(n9805), .A2(n8192), .ZN(n9793) );
  OR2_X1 U5864 ( .A1(n8179), .A2(n4858), .ZN(n8182) );
  NAND2_X1 U5865 ( .A1(n8155), .A2(n8154), .ZN(n9961) );
  OR2_X1 U5866 ( .A1(n8142), .A2(n6792), .ZN(n8144) );
  NAND2_X1 U5867 ( .A1(n5230), .A2(n8005), .ZN(n8010) );
  NAND2_X1 U5868 ( .A1(n8009), .A2(n8008), .ZN(n9986) );
  NAND2_X1 U5869 ( .A1(n7114), .A2(n8570), .ZN(n7170) );
  INV_X1 U5870 ( .A(n7111), .ZN(n7231) );
  NAND2_X1 U5871 ( .A1(n6986), .A2(n6898), .ZN(n7051) );
  INV_X1 U5872 ( .A(n9898), .ZN(n10640) );
  INV_X1 U5873 ( .A(n4947), .ZN(n4946) );
  OAI21_X1 U5874 ( .B1(n9914), .B2(n10001), .A(n9912), .ZN(n4947) );
  NAND2_X1 U5875 ( .A1(n9926), .A2(n4997), .ZN(n10012) );
  INV_X1 U5876 ( .A(n4998), .ZN(n4997) );
  OAI21_X1 U5877 ( .B1(n9927), .B2(n10582), .A(n9925), .ZN(n4998) );
  INV_X1 U5878 ( .A(P1_IR_REG_29__SCAN_IN), .ZN(n4986) );
  AOI21_X1 U5879 ( .B1(n6446), .B2(n6445), .A(n6318), .ZN(n6447) );
  NAND2_X1 U5880 ( .A1(n6231), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6225) );
  XNOR2_X1 U5881 ( .A(n6045), .B(n6044), .ZN(n8208) );
  NAND2_X1 U5882 ( .A1(n5290), .A2(n6026), .ZN(n6045) );
  OR2_X1 U5883 ( .A1(n6028), .A2(n6027), .ZN(n5290) );
  INV_X1 U5884 ( .A(n8595), .ZN(n6579) );
  NAND2_X1 U5885 ( .A1(n5834), .A2(n5854), .ZN(n7857) );
  NAND2_X1 U5886 ( .A1(n5260), .A2(n5259), .ZN(n5854) );
  NAND2_X1 U5887 ( .A1(n5283), .A2(n5280), .ZN(n5783) );
  NAND2_X1 U5888 ( .A1(n5283), .A2(n5284), .ZN(n5762) );
  AND2_X1 U5889 ( .A1(n6311), .A2(n6310), .ZN(n7441) );
  NAND2_X1 U5890 ( .A1(n5650), .A2(n5649), .ZN(n5655) );
  NAND2_X1 U5891 ( .A1(n5650), .A2(n5634), .ZN(n7025) );
  OR2_X1 U5892 ( .A1(n5607), .A2(n5606), .ZN(n5608) );
  AND2_X1 U5893 ( .A1(n6334), .A2(n6333), .ZN(n9643) );
  OR2_X1 U5894 ( .A1(n4982), .A2(n4981), .ZN(n5554) );
  NOR2_X1 U5895 ( .A1(n10350), .A2(n10349), .ZN(n10352) );
  NOR2_X1 U5896 ( .A1(n10348), .A2(n10347), .ZN(n10349) );
  NAND2_X1 U5897 ( .A1(n4879), .A2(n5435), .ZN(n5434) );
  NAND2_X1 U5898 ( .A1(n5072), .A2(n6639), .ZN(n5436) );
  INV_X1 U5899 ( .A(n8934), .ZN(n5435) );
  AOI21_X1 U5900 ( .B1(n9366), .B2(n5425), .A(n7318), .ZN(n7327) );
  NAND2_X1 U5901 ( .A1(n5117), .A2(n5115), .ZN(P2_U3549) );
  OR2_X1 U5902 ( .A1(n10701), .A2(n5116), .ZN(n5115) );
  NAND2_X1 U5903 ( .A1(n9470), .A2(n10701), .ZN(n5117) );
  INV_X1 U5904 ( .A(P2_REG1_REG_29__SCAN_IN), .ZN(n5116) );
  AND3_X1 U5905 ( .A1(n4885), .A2(n5355), .A3(n5352), .ZN(n5487) );
  NAND2_X1 U5906 ( .A1(n8294), .A2(n10632), .ZN(n5350) );
  INV_X1 U5907 ( .A(n5349), .ZN(n5348) );
  NAND2_X1 U5908 ( .A1(n5347), .A2(n10637), .ZN(n5346) );
  OAI21_X1 U5909 ( .B1(n9917), .B2(n5351), .A(n5354), .ZN(n5349) );
  AND2_X1 U5910 ( .A1(n5446), .A2(n5460), .ZN(n4861) );
  NOR2_X1 U5911 ( .A1(n5827), .A2(n5833), .ZN(n5259) );
  XNOR2_X1 U5912 ( .A(n5298), .B(n8925), .ZN(n4862) );
  INV_X2 U5913 ( .A(n8824), .ZN(n8890) );
  INV_X1 U5914 ( .A(n5621), .ZN(n5542) );
  INV_X1 U5915 ( .A(n8788), .ZN(n5053) );
  OR2_X1 U5916 ( .A1(n5758), .A2(n5757), .ZN(n4863) );
  AND2_X1 U5917 ( .A1(n9170), .A2(n8872), .ZN(n4864) );
  AND2_X1 U5918 ( .A1(n5380), .A2(n8619), .ZN(n4865) );
  NAND2_X1 U5919 ( .A1(n9266), .A2(n5442), .ZN(n9228) );
  INV_X1 U5920 ( .A(n8363), .ZN(n4988) );
  NAND2_X1 U5921 ( .A1(n6030), .A2(n6029), .ZN(n8709) );
  NOR2_X1 U5922 ( .A1(n5826), .A2(SI_13_), .ZN(n5827) );
  INV_X1 U5923 ( .A(n8805), .ZN(n5204) );
  INV_X1 U5924 ( .A(n8294), .ZN(n9917) );
  AND2_X1 U5925 ( .A1(n8318), .A2(n8279), .ZN(n8294) );
  AND2_X1 U5926 ( .A1(n5173), .A2(n9576), .ZN(n4866) );
  AND2_X1 U5927 ( .A1(n5088), .A2(n9140), .ZN(n4867) );
  NAND2_X1 U5928 ( .A1(n8823), .A2(n8822), .ZN(n5067) );
  INV_X1 U5930 ( .A(n9183), .ZN(n9178) );
  AND2_X1 U5931 ( .A1(n8872), .A2(n8870), .ZN(n9183) );
  INV_X1 U5932 ( .A(n8915), .ZN(n7843) );
  AND2_X1 U5933 ( .A1(n8818), .A2(n8819), .ZN(n8915) );
  AND2_X1 U5934 ( .A1(n5432), .A2(n9317), .ZN(n4868) );
  INV_X1 U5935 ( .A(n9328), .ZN(n9336) );
  AND2_X1 U5936 ( .A1(n8708), .A2(n8707), .ZN(n9328) );
  NOR2_X1 U5937 ( .A1(n5479), .A2(n4921), .ZN(n4869) );
  INV_X1 U5938 ( .A(n9130), .ZN(n9303) );
  AND2_X1 U5939 ( .A1(n8840), .A2(n8841), .ZN(n9130) );
  NAND2_X1 U5940 ( .A1(n9837), .A2(n8166), .ZN(n4870) );
  INV_X1 U5941 ( .A(n5259), .ZN(n5258) );
  NAND2_X1 U5942 ( .A1(n8798), .A2(n8796), .ZN(n7492) );
  INV_X1 U5943 ( .A(n7492), .ZN(n8909) );
  INV_X1 U5944 ( .A(P2_IR_REG_25__SCAN_IN), .ZN(n5451) );
  NAND2_X1 U5945 ( .A1(n5260), .A2(n5261), .ZN(n4871) );
  INV_X1 U5946 ( .A(n10521), .ZN(n6257) );
  AND2_X1 U5947 ( .A1(n5806), .A2(n5805), .ZN(n4872) );
  NAND2_X1 U5948 ( .A1(n5814), .A2(n5813), .ZN(n10294) );
  INV_X1 U5949 ( .A(n10294), .ZN(n5203) );
  NAND2_X1 U5950 ( .A1(n8889), .A2(n9317), .ZN(n4873) );
  AND2_X1 U5951 ( .A1(n5183), .A2(n5182), .ZN(n4874) );
  AND2_X1 U5952 ( .A1(n8777), .A2(n5123), .ZN(n4875) );
  AND2_X1 U5953 ( .A1(n5315), .A2(n7539), .ZN(n4876) );
  AND2_X1 U5954 ( .A1(n5317), .A2(n8966), .ZN(n4877) );
  INV_X1 U5955 ( .A(n5234), .ZN(n5233) );
  NAND2_X1 U5956 ( .A1(n7856), .A2(n7849), .ZN(n5234) );
  AND4_X1 U5957 ( .A1(n5725), .A2(n5724), .A3(n5723), .A4(n5722), .ZN(n7582)
         );
  INV_X1 U5958 ( .A(n7582), .ZN(n5120) );
  XNOR2_X1 U5959 ( .A(n8350), .B(n8349), .ZN(n9490) );
  NAND2_X1 U5960 ( .A1(n8665), .A2(n8664), .ZN(n4878) );
  INV_X1 U5961 ( .A(n9317), .ZN(n5298) );
  NAND2_X1 U5962 ( .A1(n7647), .A2(n7646), .ZN(n10641) );
  INV_X1 U5963 ( .A(n10641), .ZN(n5187) );
  NAND2_X1 U5964 ( .A1(n7558), .A2(n5403), .ZN(n7559) );
  INV_X1 U5965 ( .A(n9772), .ZN(n6904) );
  OR4_X1 U5966 ( .A1(n10050), .A2(n9371), .A3(n6646), .A4(n8932), .ZN(n4879)
         );
  NAND2_X1 U5967 ( .A1(n6603), .A2(n8387), .ZN(n6792) );
  NAND2_X1 U5968 ( .A1(n5447), .A2(n8751), .ZN(n8758) );
  AND2_X1 U5969 ( .A1(n8603), .A2(n5530), .ZN(n5590) );
  AND2_X1 U5970 ( .A1(n8526), .A2(n8527), .ZN(n9764) );
  AND2_X1 U5971 ( .A1(n7940), .A2(n7939), .ZN(n4880) );
  NOR2_X1 U5972 ( .A1(n7521), .A2(n5018), .ZN(n4881) );
  AND2_X1 U5973 ( .A1(n5053), .A2(n8783), .ZN(n4882) );
  NAND2_X1 U5974 ( .A1(n6055), .A2(n6054), .ZN(n9420) );
  INV_X1 U5975 ( .A(n9420), .ZN(n9226) );
  INV_X1 U5976 ( .A(n5466), .ZN(n5465) );
  NAND2_X1 U5977 ( .A1(n9280), .A2(n5467), .ZN(n5466) );
  XNOR2_X1 U5978 ( .A(n6325), .B(n6324), .ZN(n6602) );
  NOR2_X1 U5979 ( .A1(n6218), .A2(n6217), .ZN(n6237) );
  INV_X1 U5980 ( .A(n5281), .ZN(n5280) );
  NAND2_X1 U5981 ( .A1(n5284), .A2(n5282), .ZN(n5281) );
  NAND2_X1 U5982 ( .A1(n6303), .A2(n6236), .ZN(n6288) );
  AND2_X1 U5983 ( .A1(n10659), .A2(n5204), .ZN(n4883) );
  AND3_X1 U5984 ( .A1(n8515), .A2(n9822), .A3(n9809), .ZN(n4884) );
  NAND2_X1 U5985 ( .A1(n9220), .A2(n9139), .ZN(n9205) );
  NAND2_X1 U5986 ( .A1(n5177), .A2(n5395), .ZN(n9514) );
  OR2_X1 U5987 ( .A1(n8285), .A2(n10626), .ZN(n4885) );
  AND2_X1 U5988 ( .A1(n8848), .A2(n9230), .ZN(n9245) );
  OAI21_X1 U5989 ( .B1(n7857), .B2(n5609), .A(n5841), .ZN(n7985) );
  INV_X1 U5990 ( .A(n9743), .ZN(n9753) );
  INV_X1 U5991 ( .A(P1_IR_REG_30__SCAN_IN), .ZN(n6443) );
  NAND2_X1 U5992 ( .A1(n8882), .A2(n8868), .ZN(n9144) );
  INV_X1 U5993 ( .A(n9144), .ZN(n5078) );
  INV_X1 U5994 ( .A(n8874), .ZN(n5438) );
  INV_X1 U5995 ( .A(n8356), .ZN(n5002) );
  AND2_X1 U5996 ( .A1(n8422), .A2(n8419), .ZN(n8371) );
  INV_X1 U5997 ( .A(n5417), .ZN(n5415) );
  NOR2_X1 U5998 ( .A1(n8699), .A2(n5418), .ZN(n5417) );
  NAND2_X1 U5999 ( .A1(n9244), .A2(n5462), .ZN(n9220) );
  AND2_X1 U6000 ( .A1(n5495), .A2(n5496), .ZN(n4886) );
  NAND2_X1 U6001 ( .A1(n9405), .A2(n9143), .ZN(n4887) );
  OR2_X1 U6002 ( .A1(n7693), .A2(n7694), .ZN(n8806) );
  NAND2_X1 U6003 ( .A1(n5566), .A2(n5422), .ZN(n5610) );
  NAND2_X1 U6004 ( .A1(n8311), .A2(n5852), .ZN(n4888) );
  AND4_X1 U6005 ( .A1(n5785), .A2(n5764), .A3(n5677), .A4(n5838), .ZN(n4889)
         );
  AND2_X1 U6006 ( .A1(n5639), .A2(n5638), .ZN(n10546) );
  NAND2_X1 U6007 ( .A1(n8211), .A2(n8210), .ZN(n9939) );
  NAND2_X1 U6008 ( .A1(n5878), .A2(n5877), .ZN(n9124) );
  AND2_X1 U6009 ( .A1(n8845), .A2(n8844), .ZN(n9133) );
  NAND2_X1 U6010 ( .A1(n5947), .A2(n5946), .ZN(n9448) );
  AND2_X1 U6011 ( .A1(n6068), .A2(n5306), .ZN(n4890) );
  AND2_X1 U6012 ( .A1(n9133), .A2(n8842), .ZN(n4891) );
  AND2_X1 U6013 ( .A1(n8833), .A2(n8834), .ZN(n9347) );
  INV_X1 U6014 ( .A(n9347), .ZN(n5446) );
  AND2_X1 U6015 ( .A1(n8070), .A2(n8065), .ZN(n4892) );
  NAND2_X1 U6016 ( .A1(n8262), .A2(n8261), .ZN(n9920) );
  NAND2_X1 U6017 ( .A1(n8182), .A2(n8181), .ZN(n9950) );
  NAND2_X1 U6018 ( .A1(n9829), .A2(n5185), .ZN(n5186) );
  NAND2_X1 U6019 ( .A1(n9954), .A2(n9810), .ZN(n4893) );
  NAND2_X1 U6020 ( .A1(n5755), .A2(n5756), .ZN(n4894) );
  INV_X1 U6021 ( .A(n5286), .ZN(n5285) );
  NAND2_X1 U6022 ( .A1(n4863), .A2(n5732), .ZN(n5286) );
  AND2_X1 U6023 ( .A1(n6276), .A2(n6275), .ZN(n4895) );
  INV_X1 U6024 ( .A(n5067), .ZN(n8821) );
  NAND3_X1 U6025 ( .A1(n5552), .A2(n5550), .A3(n5070), .ZN(n9067) );
  INV_X1 U6026 ( .A(n9067), .ZN(n5071) );
  AND2_X1 U6027 ( .A1(n8514), .A2(n9846), .ZN(n4896) );
  AND2_X1 U6028 ( .A1(n9944), .A2(n9811), .ZN(n4897) );
  INV_X1 U6029 ( .A(n5137), .ZN(n5136) );
  AND2_X1 U6030 ( .A1(n4885), .A2(n5353), .ZN(n4898) );
  AND2_X1 U6031 ( .A1(n5419), .A2(n5417), .ZN(n4899) );
  NAND2_X1 U6032 ( .A1(n8447), .A2(n8401), .ZN(n8536) );
  INV_X2 U6033 ( .A(n6603), .ZN(n5192) );
  AND2_X1 U6034 ( .A1(n8929), .A2(n8928), .ZN(n4900) );
  AND2_X1 U6035 ( .A1(n9287), .A2(n9293), .ZN(n4901) );
  NAND3_X1 U6036 ( .A1(n6317), .A2(n6319), .A3(n6219), .ZN(n6314) );
  INV_X1 U6037 ( .A(n6314), .ZN(n5044) );
  AND2_X1 U6038 ( .A1(n8755), .A2(n8751), .ZN(n4902) );
  INV_X1 U6039 ( .A(n5443), .ZN(n5442) );
  NAND2_X1 U6040 ( .A1(n9245), .A2(n8852), .ZN(n5443) );
  INV_X1 U6041 ( .A(n5322), .ZN(n5321) );
  NAND2_X1 U6042 ( .A1(n5323), .A2(n6005), .ZN(n5322) );
  NOR2_X1 U6043 ( .A1(n7946), .A2(n9620), .ZN(n4903) );
  INV_X1 U6044 ( .A(P2_IR_REG_18__SCAN_IN), .ZN(n5330) );
  AND2_X1 U6045 ( .A1(n5871), .A2(n10192), .ZN(n4904) );
  AND2_X1 U6046 ( .A1(n8889), .A2(n5542), .ZN(n4905) );
  INV_X1 U6047 ( .A(n5268), .ZN(n5988) );
  OAI21_X1 U6048 ( .B1(n5927), .B2(n5272), .A(n5269), .ZN(n5268) );
  NAND2_X1 U6049 ( .A1(n4859), .A2(n5327), .ZN(n4906) );
  AND2_X1 U6050 ( .A1(n10683), .A2(n9060), .ZN(n4907) );
  NOR2_X1 U6051 ( .A1(n9400), .A2(n9185), .ZN(n4908) );
  NOR2_X1 U6052 ( .A1(n9110), .A2(n9339), .ZN(n4909) );
  NAND2_X1 U6053 ( .A1(n9883), .A2(n5235), .ZN(n9836) );
  NAND2_X1 U6054 ( .A1(n5553), .A2(n5503), .ZN(n4910) );
  AND2_X1 U6055 ( .A1(n7243), .A2(n5648), .ZN(n4911) );
  AND2_X1 U6056 ( .A1(n9217), .A2(n9233), .ZN(n4912) );
  OR2_X1 U6057 ( .A1(n6232), .A2(P1_IR_REG_23__SCAN_IN), .ZN(n4913) );
  INV_X1 U6058 ( .A(n5276), .ZN(n5275) );
  NOR2_X1 U6059 ( .A1(n5963), .A2(n5277), .ZN(n5276) );
  AND2_X1 U6060 ( .A1(n5588), .A2(n5587), .ZN(n6974) );
  AND2_X1 U6061 ( .A1(n5281), .A2(n4970), .ZN(n4914) );
  INV_X1 U6062 ( .A(n7420), .ZN(n5313) );
  AND2_X1 U6063 ( .A1(n4987), .A2(n8557), .ZN(n4915) );
  AND2_X1 U6064 ( .A1(n8784), .A2(n8785), .ZN(n4916) );
  AND2_X1 U6065 ( .A1(n5512), .A2(n5330), .ZN(n4917) );
  INV_X1 U6066 ( .A(n5097), .ZN(n5096) );
  AND2_X1 U6067 ( .A1(n9162), .A2(n4887), .ZN(n5097) );
  INV_X1 U6068 ( .A(n9170), .ZN(n9162) );
  AND2_X1 U6069 ( .A1(n8877), .A2(n8874), .ZN(n9170) );
  INV_X1 U6070 ( .A(n4969), .ZN(n4968) );
  NAND2_X1 U6071 ( .A1(n5278), .A2(n4970), .ZN(n4969) );
  AND4_X1 U6072 ( .A1(n6157), .A2(n5515), .A3(n5330), .A4(n5512), .ZN(n4918)
         );
  AND2_X1 U6073 ( .A1(n5095), .A2(n5078), .ZN(n4919) );
  OR2_X1 U6074 ( .A1(n9961), .A2(n9824), .ZN(n4920) );
  NOR2_X1 U6075 ( .A1(n9928), .A2(n9614), .ZN(n4921) );
  AND2_X1 U6076 ( .A1(n8711), .A2(n5441), .ZN(n4922) );
  NOR2_X1 U6077 ( .A1(n5445), .A2(n5444), .ZN(n4923) );
  INV_X1 U6078 ( .A(n8531), .ZN(n9727) );
  AND2_X1 U6079 ( .A1(n10290), .A2(n5849), .ZN(n4924) );
  AND2_X1 U6080 ( .A1(n7109), .A2(n6917), .ZN(n4925) );
  NOR2_X1 U6081 ( .A1(n5252), .A2(n5872), .ZN(n5251) );
  NOR2_X1 U6082 ( .A1(n5446), .A2(n5130), .ZN(n5129) );
  OR2_X1 U6083 ( .A1(n10650), .A2(n9014), .ZN(n4926) );
  AND2_X1 U6084 ( .A1(n9266), .A2(n8852), .ZN(n4927) );
  NOR2_X1 U6085 ( .A1(n8809), .A2(n5153), .ZN(n5152) );
  AND2_X1 U6086 ( .A1(n5372), .A2(n5221), .ZN(n4928) );
  AND2_X1 U6087 ( .A1(n9906), .A2(n9695), .ZN(n8591) );
  NOR2_X1 U6088 ( .A1(P2_IR_REG_28__SCAN_IN), .A2(P2_IR_REG_29__SCAN_IN), .ZN(
        n4929) );
  INV_X1 U6089 ( .A(n5827), .ZN(n5261) );
  INV_X1 U6090 ( .A(n7578), .ZN(n5454) );
  INV_X1 U6091 ( .A(n5591), .ZN(n5682) );
  INV_X2 U6092 ( .A(n5621), .ZN(n5747) );
  NAND2_X1 U6093 ( .A1(n7698), .A2(n5202), .ZN(n4930) );
  NAND2_X1 U6094 ( .A1(n7897), .A2(n5850), .ZN(n7903) );
  XOR2_X1 U6095 ( .A(n8623), .B(n8683), .Z(n4931) );
  NAND2_X1 U6096 ( .A1(n8215), .A2(n8214), .ZN(n9935) );
  INV_X1 U6097 ( .A(n9935), .ZN(n5182) );
  AND2_X1 U6098 ( .A1(n9524), .A2(n9523), .ZN(n4932) );
  AND2_X1 U6099 ( .A1(n8742), .A2(n8743), .ZN(n8830) );
  INV_X1 U6100 ( .A(n8830), .ZN(n5060) );
  NAND2_X1 U6101 ( .A1(n5790), .A2(n5789), .ZN(n8805) );
  NOR2_X1 U6102 ( .A1(n6043), .A2(SI_23_), .ZN(n4933) );
  NAND2_X1 U6103 ( .A1(n9533), .A2(n8614), .ZN(n9543) );
  NAND2_X1 U6104 ( .A1(n5103), .A2(n5102), .ZN(n9254) );
  NAND2_X1 U6105 ( .A1(n5131), .A2(n5133), .ZN(n9346) );
  INV_X1 U6106 ( .A(n9515), .ZN(n5173) );
  INV_X1 U6107 ( .A(P2_IR_REG_20__SCAN_IN), .ZN(n5493) );
  NAND2_X1 U6108 ( .A1(n5109), .A2(n5108), .ZN(n9308) );
  INV_X1 U6109 ( .A(P2_IR_REG_10__SCAN_IN), .ZN(n5764) );
  AND2_X1 U6110 ( .A1(n10678), .A2(n5471), .ZN(n4934) );
  NAND2_X1 U6111 ( .A1(n8610), .A2(n9535), .ZN(n9533) );
  INV_X1 U6112 ( .A(P2_IR_REG_6__SCAN_IN), .ZN(n5677) );
  NAND2_X1 U6113 ( .A1(n5377), .A2(n7756), .ZN(n7762) );
  INV_X1 U6114 ( .A(n5196), .ZN(n8024) );
  NOR2_X1 U6115 ( .A1(n7930), .A2(n9993), .ZN(n5196) );
  NAND2_X1 U6116 ( .A1(n8089), .A2(n5207), .ZN(n5210) );
  INV_X1 U6117 ( .A(n9223), .ZN(n9247) );
  NOR2_X1 U6118 ( .A1(n9256), .A2(n8709), .ZN(n9223) );
  INV_X1 U6119 ( .A(n5468), .ZN(n9302) );
  NAND2_X1 U6120 ( .A1(n9304), .A2(n9303), .ZN(n5468) );
  AND2_X1 U6121 ( .A1(n7850), .A2(n5233), .ZN(n4935) );
  AND2_X1 U6122 ( .A1(n6122), .A2(n6121), .ZN(n4936) );
  AND2_X1 U6123 ( .A1(n9128), .A2(n9338), .ZN(n4937) );
  OR2_X1 U6124 ( .A1(n5981), .A2(SI_20_), .ZN(n4938) );
  AND2_X1 U6125 ( .A1(n5962), .A2(n10061), .ZN(n4939) );
  OR2_X1 U6126 ( .A1(n4932), .A2(n5181), .ZN(n4940) );
  AND2_X1 U6127 ( .A1(n7728), .A2(n7727), .ZN(n4941) );
  INV_X1 U6128 ( .A(n5482), .ZN(n5110) );
  OR2_X1 U6129 ( .A1(n6744), .A2(n6743), .ZN(n10635) );
  NOR2_X1 U6130 ( .A1(n6934), .A2(n6579), .ZN(n4942) );
  INV_X1 U6131 ( .A(n7891), .ZN(n4958) );
  NAND2_X1 U6132 ( .A1(n7479), .A2(n4895), .ZN(n7491) );
  INV_X1 U6133 ( .A(P2_IR_REG_14__SCAN_IN), .ZN(n5838) );
  INV_X1 U6134 ( .A(n8570), .ZN(n5023) );
  XOR2_X1 U6135 ( .A(n7892), .B(n5868), .Z(n4943) );
  NAND2_X1 U6136 ( .A1(n5154), .A2(n8799), .ZN(n7691) );
  NAND2_X1 U6137 ( .A1(n7579), .A2(n7578), .ZN(n7619) );
  INV_X1 U6138 ( .A(n8065), .ZN(n5390) );
  NAND2_X1 U6139 ( .A1(n8140), .A2(n8139), .ZN(n9973) );
  INV_X1 U6140 ( .A(n9973), .ZN(n5193) );
  NAND2_X1 U6141 ( .A1(n7338), .A2(n4882), .ZN(n7479) );
  NAND2_X1 U6142 ( .A1(n5165), .A2(n7457), .ZN(n7558) );
  NAND2_X1 U6143 ( .A1(n6797), .A2(n8301), .ZN(n8560) );
  INV_X1 U6144 ( .A(n8560), .ZN(n5359) );
  NAND2_X1 U6145 ( .A1(n7518), .A2(n8558), .ZN(n8402) );
  INV_X1 U6146 ( .A(n8402), .ZN(n5006) );
  NAND2_X1 U6147 ( .A1(n7024), .A2(n5421), .ZN(n7125) );
  INV_X1 U6148 ( .A(n5375), .ZN(n6232) );
  NAND2_X1 U6149 ( .A1(n4859), .A2(n5478), .ZN(n6155) );
  NAND2_X1 U6150 ( .A1(n7604), .A2(n10596), .ZN(n10615) );
  INV_X1 U6151 ( .A(n10615), .ZN(n5188) );
  NAND2_X1 U6152 ( .A1(n5455), .A2(n7492), .ZN(n7579) );
  INV_X1 U6153 ( .A(n5310), .ZN(n7245) );
  AND2_X1 U6154 ( .A1(n7479), .A2(n6275), .ZN(n4944) );
  NAND4_X1 U6155 ( .A1(n5535), .A2(n5534), .A3(n5533), .A4(n5532), .ZN(n9068)
         );
  INV_X1 U6156 ( .A(n9068), .ZN(n5424) );
  NAND2_X1 U6157 ( .A1(n6607), .A2(n9772), .ZN(n8547) );
  INV_X1 U6158 ( .A(n9379), .ZN(n5212) );
  NAND2_X1 U6159 ( .A1(n7294), .A2(n6272), .ZN(n7405) );
  INV_X1 U6160 ( .A(P1_IR_REG_23__SCAN_IN), .ZN(n5374) );
  NAND2_X1 U6161 ( .A1(n5718), .A2(n5717), .ZN(n10605) );
  INV_X1 U6162 ( .A(n10605), .ZN(n5121) );
  AND2_X1 U6163 ( .A1(n7107), .A2(n6901), .ZN(n10629) );
  NAND2_X1 U6164 ( .A1(n6446), .A2(n6442), .ZN(n10029) );
  INV_X1 U6165 ( .A(P2_DATAO_REG_3__SCAN_IN), .ZN(n4963) );
  INV_X1 U6166 ( .A(P1_ADDR_REG_19__SCAN_IN), .ZN(n5085) );
  AOI21_X1 U6167 ( .B1(n4945), .B2(n10401), .A(n9691), .ZN(n9692) );
  XNOR2_X1 U6168 ( .A(n9688), .B(n9687), .ZN(n4945) );
  NAND2_X1 U6169 ( .A1(n9913), .A2(n4946), .ZN(n5215) );
  NAND2_X1 U6170 ( .A1(n10620), .A2(n7663), .ZN(n5367) );
  NAND2_X2 U6171 ( .A1(n9807), .A2(n8463), .ZN(n9799) );
  INV_X1 U6172 ( .A(n5247), .ZN(n5246) );
  NAND2_X1 U6173 ( .A1(n7925), .A2(n5336), .ZN(n5335) );
  NAND2_X1 U6174 ( .A1(n5017), .A2(n5016), .ZN(n5011) );
  NAND2_X1 U6175 ( .A1(n5245), .A2(n5243), .ZN(n5675) );
  NAND2_X1 U6176 ( .A1(n7907), .A2(n4924), .ZN(n4948) );
  NAND2_X1 U6177 ( .A1(n4952), .A2(n4954), .ZN(n5942) );
  NAND2_X1 U6178 ( .A1(n5886), .A2(n4956), .ZN(n4952) );
  NAND2_X1 U6179 ( .A1(n5480), .A2(n8362), .ZN(n7166) );
  INV_X1 U6180 ( .A(n5502), .ZN(n5500) );
  NAND2_X1 U6181 ( .A1(n5553), .A2(n4982), .ZN(n5564) );
  OAI21_X1 U6182 ( .B1(n5234), .B2(n7728), .A(n4983), .ZN(n8004) );
  NAND2_X2 U6183 ( .A1(n6470), .A2(n10041), .ZN(n8268) );
  OR2_X1 U6184 ( .A1(n5023), .A2(n4988), .ZN(n4987) );
  XNOR2_X2 U6185 ( .A(n10528), .B(n4989), .ZN(n8363) );
  INV_X1 U6186 ( .A(n5012), .ZN(n5016) );
  NAND2_X1 U6187 ( .A1(n5019), .A2(n5003), .ZN(n8477) );
  NAND3_X1 U6188 ( .A1(n5008), .A2(n5007), .A3(n5005), .ZN(n5019) );
  NAND2_X1 U6189 ( .A1(n5011), .A2(n8407), .ZN(n10620) );
  INV_X1 U6190 ( .A(n8407), .ZN(n5013) );
  NAND2_X1 U6191 ( .A1(n5017), .A2(n8416), .ZN(n8471) );
  INV_X1 U6192 ( .A(n8472), .ZN(n5014) );
  NAND3_X1 U6193 ( .A1(n5027), .A2(n9859), .A3(n8513), .ZN(n5026) );
  NAND3_X1 U6194 ( .A1(n8510), .A2(n9878), .A3(n8509), .ZN(n5027) );
  NAND2_X2 U6195 ( .A1(n6772), .A2(n6771), .ZN(n6925) );
  NAND2_X1 U6196 ( .A1(n5029), .A2(n5262), .ZN(n8550) );
  NAND3_X1 U6197 ( .A1(n5032), .A2(n5030), .A3(n5264), .ZN(n5029) );
  NAND2_X1 U6198 ( .A1(n5238), .A2(n5034), .ZN(n5037) );
  OAI21_X1 U6199 ( .B1(n8555), .B2(n8452), .A(n5035), .ZN(n5034) );
  NAND2_X1 U6200 ( .A1(n5037), .A2(n5236), .ZN(n8602) );
  NAND4_X1 U6201 ( .A1(n5045), .A2(n5372), .A3(n6237), .A4(n5044), .ZN(n5043)
         );
  NAND4_X1 U6202 ( .A1(n6221), .A2(n6222), .A3(n6223), .A4(n6220), .ZN(n5047)
         );
  OAI211_X1 U6203 ( .C1(n5048), .C2(n5053), .A(n8908), .B(n8792), .ZN(n5052)
         );
  NAND3_X1 U6204 ( .A1(n5073), .A2(n8930), .A3(n5427), .ZN(n5072) );
  AND3_X1 U6205 ( .A1(n5478), .A2(n4859), .A3(n5451), .ZN(n6152) );
  NAND3_X1 U6206 ( .A1(n5478), .A2(n4859), .A3(n5080), .ZN(n5524) );
  NAND4_X1 U6207 ( .A1(n5478), .A2(n4859), .A3(n5080), .A4(n4929), .ZN(n9485)
         );
  NAND2_X1 U6208 ( .A1(n5602), .A2(n5601), .ZN(n5607) );
  NAND2_X1 U6209 ( .A1(n5583), .A2(n5582), .ZN(n5081) );
  NAND3_X1 U6210 ( .A1(n5453), .A2(n4926), .A3(n5082), .ZN(n7621) );
  NAND3_X1 U6211 ( .A1(n5297), .A2(n5085), .A3(n5084), .ZN(n5296) );
  NAND2_X1 U6212 ( .A1(n9244), .A2(n4867), .ZN(n5086) );
  NAND2_X1 U6213 ( .A1(n5086), .A2(n5087), .ZN(n9190) );
  NAND2_X1 U6214 ( .A1(n9177), .A2(n4919), .ZN(n5090) );
  NAND2_X1 U6215 ( .A1(n9177), .A2(n9178), .ZN(n5098) );
  NAND2_X1 U6216 ( .A1(n9327), .A2(n5104), .ZN(n5103) );
  OR2_X1 U6217 ( .A1(n8310), .A2(n9059), .ZN(n5114) );
  MUX2_X1 U6218 ( .A(P2_DATAO_REG_5__SCAN_IN), .B(P1_DATAO_REG_5__SCAN_IN), 
        .S(n6597), .Z(n5629) );
  MUX2_X1 U6219 ( .A(P2_DATAO_REG_6__SCAN_IN), .B(P1_DATAO_REG_6__SCAN_IN), 
        .S(n6597), .Z(n5651) );
  MUX2_X1 U6220 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(P1_DATAO_REG_4__SCAN_IN), 
        .S(n6597), .Z(n5603) );
  MUX2_X1 U6221 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(P1_DATAO_REG_10__SCAN_IN), 
        .S(n6597), .Z(n5753) );
  MUX2_X1 U6222 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(P1_DATAO_REG_9__SCAN_IN), 
        .S(n6597), .Z(n5734) );
  MUX2_X1 U6223 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(P1_DATAO_REG_8__SCAN_IN), 
        .S(n6597), .Z(n5713) );
  MUX2_X1 U6224 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(P1_DATAO_REG_11__SCAN_IN), 
        .S(n6597), .Z(n5760) );
  OAI21_X1 U6225 ( .B1(n7302), .B2(n5125), .A(n4875), .ZN(n7328) );
  OAI21_X2 U6226 ( .B1(n4916), .B2(n7328), .A(n6260), .ZN(n7476) );
  NAND2_X1 U6227 ( .A1(n8084), .A2(n5129), .ZN(n5126) );
  OAI21_X1 U6228 ( .B1(n8084), .B2(n8083), .A(n8745), .ZN(n8706) );
  AOI21_X1 U6229 ( .B1(n8083), .B2(n8745), .A(n5138), .ZN(n5137) );
  NAND2_X1 U6230 ( .A1(n5142), .A2(n9272), .ZN(n5141) );
  OAI21_X1 U6231 ( .B1(n9272), .B2(n5144), .A(n5142), .ZN(n9227) );
  INV_X1 U6232 ( .A(n7581), .ZN(n5147) );
  NAND2_X1 U6233 ( .A1(n5152), .A2(n5147), .ZN(n5150) );
  NAND3_X1 U6234 ( .A1(n5150), .A2(n8806), .A3(n5148), .ZN(n7833) );
  NAND3_X1 U6235 ( .A1(n5150), .A2(n5149), .A3(n5148), .ZN(n7834) );
  NAND2_X1 U6236 ( .A1(n7581), .A2(n5155), .ZN(n5154) );
  INV_X1 U6237 ( .A(n5155), .ZN(n5151) );
  NAND2_X1 U6238 ( .A1(n7581), .A2(n8796), .ZN(n7615) );
  NAND2_X1 U6239 ( .A1(n6259), .A2(n6974), .ZN(n5158) );
  NAND2_X2 U6240 ( .A1(n8765), .A2(n5158), .ZN(n8900) );
  NAND2_X1 U6241 ( .A1(n7348), .A2(n5157), .ZN(n8765) );
  AND2_X1 U6242 ( .A1(n5593), .A2(n5592), .ZN(n5159) );
  NAND3_X1 U6243 ( .A1(n5403), .A2(n5402), .A3(n7558), .ZN(n7710) );
  NAND2_X1 U6244 ( .A1(n7461), .A2(n7458), .ZN(n5165) );
  NAND2_X1 U6245 ( .A1(n7461), .A2(n7460), .ZN(n7557) );
  NAND2_X2 U6246 ( .A1(n7794), .A2(n7793), .ZN(n7942) );
  NAND3_X1 U6247 ( .A1(n5377), .A2(n7756), .A3(n5376), .ZN(n7794) );
  NAND2_X1 U6248 ( .A1(n5166), .A2(n5167), .ZN(n9574) );
  NAND3_X1 U6249 ( .A1(n9585), .A2(n9589), .A3(n5168), .ZN(n5166) );
  NAND3_X1 U6250 ( .A1(n9585), .A2(n9589), .A3(n5398), .ZN(n5177) );
  NAND2_X1 U6251 ( .A1(n9554), .A2(n5180), .ZN(n5179) );
  NAND3_X1 U6252 ( .A1(n5384), .A2(n7127), .A3(n7126), .ZN(n7452) );
  NAND3_X1 U6253 ( .A1(n8111), .A2(n8112), .A3(n8116), .ZN(n8122) );
  AND2_X2 U6254 ( .A1(n9829), .A2(n4874), .ZN(n9769) );
  INV_X1 U6255 ( .A(n5186), .ZN(n9794) );
  NOR2_X2 U6256 ( .A1(n7605), .A2(n10577), .ZN(n7604) );
  INV_X2 U6257 ( .A(n10491), .ZN(n6995) );
  INV_X1 U6258 ( .A(n7054), .ZN(n5190) );
  NAND2_X1 U6259 ( .A1(n10491), .A2(n6989), .ZN(n7054) );
  AND3_X2 U6260 ( .A1(n6601), .A2(n6600), .A3(n5191), .ZN(n10491) );
  NAND2_X1 U6261 ( .A1(n9733), .A2(n5199), .ZN(n8330) );
  NAND2_X1 U6262 ( .A1(n9733), .A2(n8292), .ZN(n9710) );
  NAND2_X1 U6263 ( .A1(n5200), .A2(n7698), .ZN(n7986) );
  INV_X1 U6264 ( .A(n5210), .ZN(n9311) );
  NOR2_X2 U6265 ( .A1(n10519), .A2(n7348), .ZN(n7298) );
  NOR2_X2 U6266 ( .A1(n9191), .A2(n9405), .ZN(n9164) );
  NAND2_X2 U6267 ( .A1(n6643), .A2(n6597), .ZN(n5609) );
  NAND2_X2 U6268 ( .A1(n6188), .A2(n6646), .ZN(n6643) );
  NAND2_X1 U6269 ( .A1(n6918), .A2(n4925), .ZN(n5214) );
  MUX2_X1 U6270 ( .A(P1_REG1_REG_29__SCAN_IN), .B(n5215), .S(n10634), .Z(
        P1_U3552) );
  MUX2_X1 U6271 ( .A(P1_REG0_REG_29__SCAN_IN), .B(n5215), .S(n10637), .Z(
        P1_U3520) );
  NAND2_X1 U6272 ( .A1(n9806), .A2(n5218), .ZN(n5217) );
  NAND2_X1 U6273 ( .A1(n9730), .A2(n5226), .ZN(n5224) );
  NAND2_X1 U6274 ( .A1(n5224), .A2(n5222), .ZN(n8318) );
  NAND2_X1 U6275 ( .A1(n5224), .A2(n5225), .ZN(n8278) );
  NAND2_X1 U6276 ( .A1(n8004), .A2(n8491), .ZN(n5230) );
  NAND3_X1 U6277 ( .A1(n6986), .A2(n6898), .A3(n5231), .ZN(n7053) );
  NAND2_X1 U6278 ( .A1(n9630), .A2(n10512), .ZN(n8564) );
  NAND2_X1 U6279 ( .A1(n6988), .A2(n6987), .ZN(n6986) );
  NAND2_X2 U6280 ( .A1(n9885), .A2(n9884), .ZN(n9883) );
  NAND2_X1 U6281 ( .A1(n8257), .A2(n8531), .ZN(n9730) );
  OAI21_X1 U6282 ( .B1(n7643), .B2(n7642), .A(n7641), .ZN(n10614) );
  NAND2_X1 U6283 ( .A1(n7168), .A2(n8364), .ZN(n7203) );
  AND2_X2 U6284 ( .A1(n6932), .A2(n8569), .ZN(n7112) );
  XNOR2_X1 U6285 ( .A(n8328), .B(n8380), .ZN(n9914) );
  OAI21_X1 U6286 ( .B1(n8555), .B2(n5241), .A(n5240), .ZN(n5239) );
  AOI21_X1 U6287 ( .B1(n8554), .B2(n6904), .A(n6579), .ZN(n5240) );
  OAI21_X1 U6288 ( .B1(n5633), .B2(n5248), .A(n5246), .ZN(n5670) );
  NAND2_X1 U6289 ( .A1(n5633), .A2(n5246), .ZN(n5245) );
  NAND2_X1 U6290 ( .A1(n5829), .A2(n5251), .ZN(n5249) );
  NAND2_X1 U6291 ( .A1(n6007), .A2(n5288), .ZN(n5287) );
  NAND2_X1 U6292 ( .A1(n6007), .A2(n6006), .ZN(n6028) );
  NAND2_X1 U6293 ( .A1(n5287), .A2(n5291), .ZN(n6052) );
  NAND3_X1 U6294 ( .A1(n5498), .A2(P2_ADDR_REG_19__SCAN_IN), .A3(
        P1_ADDR_REG_19__SCAN_IN), .ZN(n5295) );
  NAND2_X2 U6295 ( .A1(n5299), .A2(n5298), .ZN(n5621) );
  NAND2_X4 U6296 ( .A1(n5523), .A2(n8926), .ZN(n10693) );
  NAND2_X1 U6298 ( .A1(n6103), .A2(n5303), .ZN(n5300) );
  NAND2_X1 U6299 ( .A1(n5300), .A2(n5301), .ZN(n6182) );
  NAND2_X1 U6300 ( .A1(n5308), .A2(n5311), .ZN(n5664) );
  NAND2_X1 U6301 ( .A1(n7224), .A2(n5309), .ZN(n5308) );
  NAND2_X1 U6302 ( .A1(n7571), .A2(n5752), .ZN(n5314) );
  NAND2_X1 U6303 ( .A1(n5314), .A2(n4876), .ZN(n7542) );
  NAND2_X1 U6304 ( .A1(n7159), .A2(n5695), .ZN(n5316) );
  NAND2_X1 U6305 ( .A1(n5316), .A2(n4877), .ZN(n8971) );
  NAND2_X1 U6306 ( .A1(n4859), .A2(n5328), .ZN(n5517) );
  OAI21_X1 U6307 ( .B1(n7925), .B2(n5332), .A(n5331), .ZN(n8013) );
  AOI21_X1 U6308 ( .B1(n5474), .B2(n7856), .A(n5337), .ZN(n5331) );
  INV_X1 U6309 ( .A(n5474), .ZN(n5332) );
  NAND2_X1 U6310 ( .A1(n5335), .A2(n5333), .ZN(n8046) );
  INV_X1 U6311 ( .A(n5334), .ZN(n5333) );
  OAI21_X1 U6312 ( .B1(n5474), .B2(n5337), .A(n8500), .ZN(n5334) );
  NOR2_X1 U6313 ( .A1(n7856), .A2(n5337), .ZN(n5336) );
  NAND2_X1 U6314 ( .A1(n7924), .A2(n5474), .ZN(n8012) );
  NAND3_X1 U6315 ( .A1(n5339), .A2(n8527), .A3(n5338), .ZN(n9752) );
  NAND3_X1 U6316 ( .A1(n5340), .A2(n9764), .A3(n5342), .ZN(n5338) );
  NAND3_X1 U6317 ( .A1(n9799), .A2(n5340), .A3(n9764), .ZN(n5339) );
  INV_X1 U6318 ( .A(n5345), .ZN(n9778) );
  INV_X1 U6319 ( .A(n5352), .ZN(n5347) );
  OAI211_X1 U6320 ( .C1(n4898), .C2(n10635), .A(n5348), .B(n5346), .ZN(
        P1_U3519) );
  NAND3_X1 U6321 ( .A1(n4898), .A2(n5350), .A3(n5352), .ZN(n10010) );
  NAND2_X1 U6322 ( .A1(n8561), .A2(n8359), .ZN(n7059) );
  NAND2_X1 U6323 ( .A1(n9718), .A2(n9717), .ZN(n9716) );
  NAND2_X1 U6324 ( .A1(n5367), .A2(n5364), .ZN(n7871) );
  OAI21_X1 U6325 ( .B1(n5371), .B2(n5370), .A(n9859), .ZN(n5369) );
  NAND2_X1 U6326 ( .A1(n8610), .A2(n4865), .ZN(n5379) );
  OAI21_X2 U6327 ( .B1(n8610), .B2(n5382), .A(n4865), .ZN(n8625) );
  NAND2_X1 U6328 ( .A1(n7127), .A2(n7126), .ZN(n7136) );
  NAND2_X1 U6329 ( .A1(n7942), .A2(n5386), .ZN(n5385) );
  NAND3_X1 U6330 ( .A1(n5400), .A2(n8632), .A3(n5397), .ZN(n9565) );
  NAND2_X1 U6331 ( .A1(n9585), .A2(n9589), .ZN(n9505) );
  NOR2_X1 U6332 ( .A1(n6314), .A2(n5404), .ZN(n6303) );
  NAND2_X1 U6333 ( .A1(n9599), .A2(n5410), .ZN(n5406) );
  OAI211_X1 U6334 ( .C1(n9599), .C2(n5411), .A(n5406), .B(n5407), .ZN(n8697)
         );
  OR2_X2 U6335 ( .A1(n9599), .A2(n9600), .ZN(n5419) );
  NAND2_X2 U6336 ( .A1(n6608), .A2(n6581), .ZN(n8686) );
  OR2_X2 U6337 ( .A1(n6578), .A2(n8595), .ZN(n6608) );
  NAND2_X1 U6338 ( .A1(n6848), .A2(n6847), .ZN(n7024) );
  NAND2_X1 U6339 ( .A1(n7024), .A2(n7023), .ZN(n7032) );
  NAND2_X1 U6340 ( .A1(n8112), .A2(n8111), .ZN(n8117) );
  NAND3_X1 U6341 ( .A1(n5566), .A2(n5422), .A3(n5491), .ZN(n5612) );
  AND3_X2 U6342 ( .A1(n5509), .A2(n5507), .A3(n5508), .ZN(n10505) );
  NAND2_X1 U6343 ( .A1(n8732), .A2(n5429), .ZN(n5426) );
  OAI211_X1 U6344 ( .C1(n8732), .C2(n5430), .A(n5426), .B(n5428), .ZN(n5427)
         );
  NAND2_X1 U6345 ( .A1(n5436), .A2(n5434), .ZN(P2_U3244) );
  NAND2_X1 U6346 ( .A1(n9184), .A2(n4864), .ZN(n5439) );
  NAND2_X1 U6347 ( .A1(n7495), .A2(n4923), .ZN(n7581) );
  NAND2_X1 U6348 ( .A1(n6262), .A2(n8908), .ZN(n7495) );
  INV_X1 U6349 ( .A(n8798), .ZN(n5445) );
  NAND2_X1 U6350 ( .A1(n4902), .A2(n5447), .ZN(n6258) );
  NAND2_X1 U6351 ( .A1(n5449), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5497) );
  NAND3_X1 U6352 ( .A1(n4859), .A2(n5450), .A3(n5478), .ZN(n5449) );
  NAND2_X1 U6353 ( .A1(n7494), .A2(n5452), .ZN(n5453) );
  NOR2_X1 U6354 ( .A1(n7618), .A2(n5454), .ZN(n5452) );
  NAND2_X1 U6355 ( .A1(n6965), .A2(n5456), .ZN(n7294) );
  OAI21_X1 U6356 ( .B1(n7405), .B2(n8775), .A(n6273), .ZN(n6274) );
  NAND2_X1 U6357 ( .A1(n8088), .A2(n4861), .ZN(n5457) );
  NAND2_X1 U6358 ( .A1(n5457), .A2(n5458), .ZN(n9327) );
  NOR2_X1 U6359 ( .A1(n9126), .A2(n9125), .ZN(n9357) );
  NOR2_X1 U6360 ( .A1(n9302), .A2(n9132), .ZN(n9281) );
  NAND2_X1 U6361 ( .A1(n6152), .A2(n5473), .ZN(n5527) );
  INV_X1 U6362 ( .A(n7924), .ZN(n7873) );
  INV_X1 U6363 ( .A(n6988), .ZN(n8360) );
  INV_X1 U6364 ( .A(n8926), .ZN(n8896) );
  XNOR2_X1 U6365 ( .A(n6108), .B(n6107), .ZN(n8243) );
  CLKBUF_X1 U6366 ( .A(n8610), .Z(n9534) );
  NAND2_X1 U6367 ( .A1(n5557), .A2(P2_DATAO_REG_2__SCAN_IN), .ZN(n5555) );
  OR2_X1 U6368 ( .A1(n8685), .A2(n6989), .ZN(n6584) );
  OAI22_X1 U6369 ( .A1(n10512), .A2(n8686), .B1(n6797), .B2(n8685), .ZN(n6798)
         );
  NOR2_X2 U6370 ( .A1(n7056), .A2(n6925), .ZN(n6932) );
  NOR2_X2 U6371 ( .A1(n9998), .A2(n7733), .ZN(n7931) );
  NAND2_X1 U6372 ( .A1(n9319), .A2(n8739), .ZN(n9291) );
  NAND2_X1 U6373 ( .A1(n9295), .A2(n8840), .ZN(n9272) );
  AND2_X2 U6374 ( .A1(n5531), .A2(n9489), .ZN(n5589) );
  OAI21_X1 U6375 ( .B1(n9145), .B2(n8883), .A(n8882), .ZN(n8723) );
  NOR2_X1 U6376 ( .A1(n8491), .A2(n8495), .ZN(n5474) );
  AND2_X2 U6377 ( .A1(n10037), .A2(n10041), .ZN(n5475) );
  INV_X1 U6378 ( .A(n9448), .ZN(n9110) );
  AOI21_X1 U6379 ( .B1(n7910), .B2(n8915), .A(n7909), .ZN(n7911) );
  AND2_X1 U6380 ( .A1(n6582), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n5477) );
  AND4_X1 U6381 ( .A1(n5494), .A2(n4918), .A3(n6172), .A4(n5511), .ZN(n5478)
         );
  AND2_X1 U6382 ( .A1(n5523), .A2(n8932), .ZN(n9458) );
  NOR2_X1 U6383 ( .A1(n9753), .A2(n9741), .ZN(n5479) );
  INV_X1 U6384 ( .A(P2_REG3_REG_9__SCAN_IN), .ZN(n5719) );
  AND2_X1 U6385 ( .A1(n9334), .A2(n9129), .ZN(n5482) );
  INV_X1 U6386 ( .A(P1_DATAO_REG_2__SCAN_IN), .ZN(n5556) );
  AND3_X1 U6387 ( .A1(n5916), .A2(n5915), .A3(n5914), .ZN(n9338) );
  AND2_X1 U6388 ( .A1(n6001), .A2(n6000), .ZN(n9293) );
  INV_X1 U6389 ( .A(n8536), .ZN(n8277) );
  INV_X1 U6390 ( .A(n9809), .ZN(n8191) );
  NOR2_X1 U6391 ( .A1(n8183), .A2(n8172), .ZN(n5485) );
  XNOR2_X1 U6392 ( .A(n9772), .B(n8594), .ZN(n5486) );
  INV_X1 U6393 ( .A(n9164), .ZN(n9179) );
  INV_X1 U6394 ( .A(n8765), .ZN(n8766) );
  NAND2_X1 U6395 ( .A1(n8878), .A2(n8890), .ZN(n8879) );
  INV_X1 U6396 ( .A(n8539), .ZN(n8540) );
  NAND2_X1 U6397 ( .A1(n8927), .A2(n8926), .ZN(n8929) );
  NOR2_X1 U6398 ( .A1(n5523), .A2(n8896), .ZN(n8897) );
  XNOR2_X1 U6399 ( .A(n8927), .B(n8895), .ZN(n8898) );
  NOR2_X1 U6400 ( .A1(n5862), .A2(n5861), .ZN(n5879) );
  NAND2_X1 U6401 ( .A1(n7020), .A2(n7022), .ZN(n7023) );
  AND2_X1 U6402 ( .A1(n8230), .A2(P1_REG3_REG_26__SCAN_IN), .ZN(n8247) );
  INV_X1 U6403 ( .A(P1_REG3_REG_7__SCAN_IN), .ZN(n7141) );
  NOR2_X1 U6404 ( .A1(n5741), .A2(n6714), .ZN(n5770) );
  NAND2_X1 U6405 ( .A1(n8898), .A2(n8897), .ZN(n8930) );
  NAND2_X1 U6406 ( .A1(n6056), .A2(P2_REG3_REG_24__SCAN_IN), .ZN(n6073) );
  NOR2_X1 U6407 ( .A1(n5933), .A2(n10267), .ZN(n5948) );
  AND2_X1 U6408 ( .A1(n5948), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n5968) );
  OR2_X1 U6409 ( .A1(n5816), .A2(n5815), .ZN(n5843) );
  NAND2_X1 U6410 ( .A1(n9111), .A2(n9458), .ZN(n9397) );
  INV_X1 U6411 ( .A(n8804), .ZN(n7840) );
  NAND2_X1 U6412 ( .A1(n6963), .A2(n6964), .ZN(n6962) );
  NOR2_X1 U6413 ( .A1(n6989), .A2(n8686), .ZN(n6587) );
  AND2_X1 U6414 ( .A1(n8171), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n8183) );
  AND3_X1 U6415 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .A3(P1_REG3_REG_5__SCAN_IN), .ZN(n6849) );
  AND2_X1 U6416 ( .A1(n8247), .A2(P1_REG3_REG_27__SCAN_IN), .ZN(n7070) );
  NOR2_X1 U6417 ( .A1(n8157), .A2(n8156), .ZN(n8171) );
  NOR2_X1 U6418 ( .A1(n7862), .A2(n7861), .ZN(n7875) );
  INV_X1 U6419 ( .A(SI_15_), .ZN(n10192) );
  NOR2_X1 U6420 ( .A1(n5685), .A2(n5683), .ZN(n5702) );
  OR2_X1 U6421 ( .A1(n6073), .A2(n8993), .ZN(n6094) );
  AND2_X1 U6422 ( .A1(n9019), .A2(n5726), .ZN(n5727) );
  OR2_X1 U6423 ( .A1(n6094), .A2(n10272), .ZN(n6126) );
  INV_X1 U6424 ( .A(P2_REG3_REG_10__SCAN_IN), .ZN(n6714) );
  NAND2_X1 U6425 ( .A1(n9164), .A2(n9168), .ZN(n9150) );
  NAND2_X1 U6426 ( .A1(n5968), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n5994) );
  INV_X1 U6427 ( .A(n9197), .ZN(n9198) );
  NAND2_X1 U6428 ( .A1(n6175), .A2(n8928), .ZN(n6953) );
  INV_X1 U6429 ( .A(P1_REG3_REG_9__SCAN_IN), .ZN(n7463) );
  AND2_X1 U6430 ( .A1(P1_REG3_REG_22__SCAN_IN), .A2(n6693), .ZN(n6694) );
  AND2_X1 U6431 ( .A1(n7875), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8014) );
  OR2_X1 U6432 ( .A1(n8147), .A2(n6692), .ZN(n8157) );
  NAND2_X1 U6433 ( .A1(n7173), .A2(n8571), .ZN(n7518) );
  NAND2_X1 U6434 ( .A1(n8326), .A2(n8325), .ZN(n8327) );
  OR2_X1 U6435 ( .A1(n6349), .A2(P1_IR_REG_15__SCAN_IN), .ZN(n6290) );
  INV_X1 U6436 ( .A(P1_IR_REG_12__SCAN_IN), .ZN(n6294) );
  XNOR2_X1 U6437 ( .A(n10521), .B(n5615), .ZN(n7220) );
  INV_X1 U6438 ( .A(n10284), .ZN(n9044) );
  AND2_X1 U6439 ( .A1(n6057), .A2(n6033), .ZN(n9248) );
  NAND2_X1 U6440 ( .A1(n6419), .A2(P2_REG0_REG_0__SCAN_IN), .ZN(n5539) );
  AND2_X1 U6441 ( .A1(n6133), .A2(n6132), .ZN(n9146) );
  INV_X1 U6442 ( .A(n9133), .ZN(n9280) );
  OR2_X1 U6443 ( .A1(n6971), .A2(n8733), .ZN(n6948) );
  INV_X1 U6444 ( .A(n8828), .ZN(n8916) );
  OR2_X1 U6445 ( .A1(n10049), .A2(n6163), .ZN(n6164) );
  INV_X1 U6446 ( .A(P2_IR_REG_23__SCAN_IN), .ZN(n6172) );
  INV_X1 U6447 ( .A(P2_IR_REG_16__SCAN_IN), .ZN(n5511) );
  OR2_X1 U6448 ( .A1(n8658), .A2(n8657), .ZN(n8659) );
  OR2_X1 U6449 ( .A1(n8631), .A2(n8630), .ZN(n8632) );
  NOR2_X1 U6450 ( .A1(n7655), .A2(n7654), .ZN(n7664) );
  OR2_X1 U6451 ( .A1(n6630), .A2(n9881), .ZN(n9569) );
  INV_X1 U6452 ( .A(n9566), .ZN(n9605) );
  NAND2_X1 U6453 ( .A1(n8598), .A2(n6623), .ZN(n8553) );
  NAND2_X1 U6454 ( .A1(n6774), .A2(P1_REG1_REG_1__SCAN_IN), .ZN(n6483) );
  AND4_X1 U6455 ( .A1(n7079), .A2(n7078), .A3(n7077), .A4(n7076), .ZN(n9721)
         );
  INV_X1 U6456 ( .A(n9939), .ZN(n9789) );
  OR3_X1 U6457 ( .A1(n10582), .A2(n6623), .A3(n8597), .ZN(n9866) );
  INV_X1 U6458 ( .A(n10618), .ZN(n10578) );
  OR2_X1 U6459 ( .A1(n6625), .A2(n6497), .ZN(n6923) );
  OR2_X1 U6460 ( .A1(n10046), .A2(P1_D_REG_0__SCAN_IN), .ZN(n6402) );
  NAND2_X1 U6461 ( .A1(n6243), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6245) );
  XNOR2_X1 U6462 ( .A(n5891), .B(n5874), .ZN(n5893) );
  INV_X1 U6463 ( .A(P1_IR_REG_31__SCAN_IN), .ZN(n6318) );
  AND2_X1 U6464 ( .A1(n6176), .A2(n9316), .ZN(n9046) );
  INV_X1 U6465 ( .A(n8939), .ZN(n10282) );
  INV_X1 U6466 ( .A(n8994), .ZN(n9049) );
  INV_X1 U6467 ( .A(n6175), .ZN(n8933) );
  AOI21_X1 U6468 ( .B1(n9180), .B2(n5591), .A(n6119), .ZN(n9053) );
  INV_X1 U6469 ( .A(n10415), .ZN(n10480) );
  OR2_X1 U6470 ( .A1(n7815), .A2(n7814), .ZN(n7969) );
  INV_X1 U6471 ( .A(n9137), .ZN(n9229) );
  INV_X1 U6472 ( .A(n9376), .ZN(n9349) );
  INV_X1 U6473 ( .A(n9359), .ZN(n9289) );
  NAND2_X1 U6474 ( .A1(n6167), .A2(n6166), .ZN(n6956) );
  INV_X1 U6475 ( .A(n10697), .ZN(n10673) );
  OR2_X1 U6476 ( .A1(n6951), .A2(n6950), .ZN(n6958) );
  NAND2_X1 U6477 ( .A1(n10408), .A2(n6164), .ZN(n10051) );
  AND2_X1 U6478 ( .A1(n5857), .A2(n5840), .ZN(n7680) );
  AND2_X1 U6479 ( .A1(n6762), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6393) );
  AOI21_X1 U6480 ( .B1(n6840), .B2(n6839), .A(n6838), .ZN(n6848) );
  AND2_X1 U6481 ( .A1(n6635), .A2(n10622), .ZN(n9566) );
  INV_X1 U6482 ( .A(n6607), .ZN(n8598) );
  AND4_X1 U6483 ( .A1(n8274), .A2(n8273), .A3(n8272), .A4(n8271), .ZN(n9726)
         );
  AND4_X1 U6484 ( .A1(n7869), .A2(n7868), .A3(n7867), .A4(n7866), .ZN(n8126)
         );
  INV_X1 U6485 ( .A(n10393), .ZN(n9678) );
  NAND2_X1 U6486 ( .A1(n8539), .A2(n8587), .ZN(n8380) );
  INV_X1 U6487 ( .A(n9764), .ZN(n9762) );
  AND2_X1 U6488 ( .A1(n9836), .A2(n9855), .ZN(n9856) );
  AND2_X1 U6489 ( .A1(n8041), .A2(n8011), .ZN(n9985) );
  INV_X1 U6490 ( .A(n10626), .ZN(n9891) );
  OR2_X1 U6491 ( .A1(n6934), .A2(n6628), .ZN(n10618) );
  OR2_X1 U6492 ( .A1(n6923), .A2(n6499), .ZN(n6744) );
  AND2_X1 U6493 ( .A1(n6299), .A2(n6298), .ZN(n7730) );
  NOR2_X1 U6494 ( .A1(n10318), .A2(n10317), .ZN(n10319) );
  NOR2_X1 U6495 ( .A1(n10344), .A2(n10343), .ZN(n10345) );
  NAND2_X1 U6496 ( .A1(n6437), .A2(n6436), .ZN(n10486) );
  INV_X1 U6497 ( .A(n6209), .ZN(n6210) );
  AND4_X1 U6498 ( .A1(n5777), .A2(n5776), .A3(n5775), .A4(n5774), .ZN(n7694)
         );
  OR2_X1 U6499 ( .A1(n10288), .A2(n5542), .ZN(n9017) );
  INV_X2 U6500 ( .A(n9009), .ZN(n10288) );
  INV_X1 U6501 ( .A(n8991), .ZN(n9186) );
  INV_X1 U6502 ( .A(n10450), .ZN(n10481) );
  NAND2_X1 U6503 ( .A1(n9378), .A2(n6282), .ZN(n9333) );
  NAND2_X1 U6504 ( .A1(n9378), .A2(n6280), .ZN(n9359) );
  OR2_X1 U6505 ( .A1(n6958), .A2(n6956), .ZN(n10699) );
  OR2_X1 U6506 ( .A1(n6958), .A2(n6957), .ZN(n10702) );
  NAND2_X1 U6507 ( .A1(n10052), .A2(n10051), .ZN(n10410) );
  INV_X1 U6508 ( .A(n7680), .ZN(n7685) );
  INV_X1 U6509 ( .A(n9607), .ZN(n9598) );
  INV_X1 U6510 ( .A(n9783), .ZN(n9754) );
  OR2_X1 U6511 ( .A1(n7880), .A2(n7879), .ZN(n9618) );
  OR2_X1 U6512 ( .A1(n10374), .A2(n10376), .ZN(n10393) );
  OR2_X1 U6513 ( .A1(P1_U3083), .A2(n6366), .ZN(n10391) );
  INV_X2 U6514 ( .A(n10633), .ZN(n10634) );
  OR2_X1 U6515 ( .A1(n6744), .A2(n6921), .ZN(n10633) );
  INV_X2 U6516 ( .A(n10635), .ZN(n10637) );
  INV_X1 U6517 ( .A(n8597), .ZN(n10047) );
  INV_X1 U6518 ( .A(P2_DATAO_REG_15__SCAN_IN), .ZN(n6893) );
  NOR2_X1 U6519 ( .A1(n10346), .A2(n10345), .ZN(n10348) );
  NOR2_X1 U6520 ( .A1(P2_IR_REG_7__SCAN_IN), .A2(P2_IR_REG_5__SCAN_IN), .ZN(
        n5489) );
  NOR2_X1 U6521 ( .A1(P2_IR_REG_11__SCAN_IN), .A2(P2_IR_REG_15__SCAN_IN), .ZN(
        n5488) );
  NAND4_X1 U6522 ( .A1(n5490), .A2(n4889), .A3(n5489), .A4(n5488), .ZN(n5492)
         );
  NAND2_X1 U6523 ( .A1(n5518), .A2(n5493), .ZN(n5514) );
  NOR2_X1 U6524 ( .A1(n5514), .A2(P2_IR_REG_24__SCAN_IN), .ZN(n5494) );
  INV_X1 U6525 ( .A(P2_IR_REG_26__SCAN_IN), .ZN(n5495) );
  INV_X1 U6526 ( .A(P2_RD_REG_SCAN_IN), .ZN(n5498) );
  NAND2_X2 U6527 ( .A1(n6643), .A2(n8387), .ZN(n5965) );
  INV_X1 U6528 ( .A(P1_DATAO_REG_1__SCAN_IN), .ZN(n6391) );
  OR2_X1 U6529 ( .A1(n5965), .A2(n6391), .ZN(n5509) );
  NAND2_X1 U6530 ( .A1(P2_IR_REG_31__SCAN_IN), .A2(P2_IR_REG_0__SCAN_IN), .ZN(
        n5499) );
  XNOR2_X1 U6531 ( .A(n5499), .B(P2_IR_REG_1__SCAN_IN), .ZN(n10421) );
  INV_X1 U6532 ( .A(n10421), .ZN(n6390) );
  OR2_X1 U6533 ( .A1(n6643), .A2(n6390), .ZN(n5508) );
  INV_X1 U6534 ( .A(P2_DATAO_REG_0__SCAN_IN), .ZN(n6467) );
  INV_X1 U6535 ( .A(SI_0_), .ZN(n5540) );
  NAND2_X1 U6536 ( .A1(n5500), .A2(SI_1_), .ZN(n5553) );
  INV_X1 U6537 ( .A(SI_1_), .ZN(n5501) );
  NAND2_X1 U6538 ( .A1(n5502), .A2(n5501), .ZN(n5503) );
  MUX2_X1 U6539 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(P2_DATAO_REG_1__SCAN_IN), 
        .S(n4854), .Z(n5504) );
  INV_X1 U6540 ( .A(n5504), .ZN(n5505) );
  NAND2_X1 U6541 ( .A1(n4910), .A2(n5505), .ZN(n5506) );
  NAND2_X1 U6542 ( .A1(n5554), .A2(n5506), .ZN(n6599) );
  OR2_X1 U6543 ( .A1(n5609), .A2(n6599), .ZN(n5507) );
  NAND2_X1 U6544 ( .A1(n4906), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5519) );
  NAND2_X1 U6545 ( .A1(n5519), .A2(n5518), .ZN(n5520) );
  NAND2_X1 U6546 ( .A1(n5517), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5516) );
  NAND2_X1 U6547 ( .A1(n8926), .A2(n8733), .ZN(n6279) );
  XNOR2_X1 U6548 ( .A(n6158), .B(n6157), .ZN(n6175) );
  OR2_X1 U6549 ( .A1(n5519), .A2(n5518), .ZN(n5521) );
  OR2_X1 U6550 ( .A1(n6175), .A2(n9317), .ZN(n5522) );
  XNOR2_X1 U6551 ( .A(n10505), .B(n6115), .ZN(n5544) );
  INV_X1 U6552 ( .A(n5531), .ZN(n8603) );
  NAND2_X1 U6553 ( .A1(n5590), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n5535) );
  INV_X1 U6554 ( .A(n5530), .ZN(n9489) );
  INV_X1 U6555 ( .A(P2_REG0_REG_1__SCAN_IN), .ZN(n5529) );
  AND2_X2 U6556 ( .A1(n5531), .A2(n5530), .ZN(n5591) );
  NAND2_X1 U6557 ( .A1(n5591), .A2(P2_REG3_REG_1__SCAN_IN), .ZN(n5532) );
  NAND2_X1 U6558 ( .A1(n5621), .A2(n9068), .ZN(n5546) );
  XNOR2_X1 U6559 ( .A(n5544), .B(n5546), .ZN(n7358) );
  NAND2_X1 U6560 ( .A1(n5589), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n5538) );
  NAND2_X1 U6561 ( .A1(n5591), .A2(P2_REG3_REG_0__SCAN_IN), .ZN(n5537) );
  NAND2_X1 U6562 ( .A1(n5590), .A2(P2_REG1_REG_0__SCAN_IN), .ZN(n5536) );
  NAND4_X1 U6563 ( .A1(n5539), .A2(n5538), .A3(n5537), .A4(n5536), .ZN(n6952)
         );
  INV_X1 U6564 ( .A(P2_IR_REG_0__SCAN_IN), .ZN(n10427) );
  NOR2_X1 U6565 ( .A1(n8387), .A2(n5540), .ZN(n5541) );
  XNOR2_X1 U6566 ( .A(n5541), .B(P1_DATAO_REG_0__SCAN_IN), .ZN(n9493) );
  MUX2_X1 U6567 ( .A(n10427), .B(n9493), .S(n6643), .Z(n7317) );
  INV_X1 U6568 ( .A(n7317), .ZN(n7313) );
  AND2_X1 U6569 ( .A1(n7317), .A2(n6115), .ZN(n7356) );
  AOI21_X1 U6570 ( .B1(n7352), .B2(n5621), .A(n7356), .ZN(n5543) );
  NAND2_X1 U6571 ( .A1(n7358), .A2(n5543), .ZN(n7357) );
  INV_X1 U6572 ( .A(n5544), .ZN(n5545) );
  NAND2_X1 U6573 ( .A1(n5546), .A2(n5545), .ZN(n5547) );
  INV_X1 U6574 ( .A(n7089), .ZN(n5575) );
  NAND2_X1 U6575 ( .A1(n5590), .A2(P2_REG1_REG_2__SCAN_IN), .ZN(n5551) );
  NAND2_X1 U6576 ( .A1(n5591), .A2(P2_REG3_REG_2__SCAN_IN), .ZN(n5549) );
  NAND2_X1 U6577 ( .A1(n5621), .A2(n9067), .ZN(n5572) );
  INV_X1 U6578 ( .A(n5564), .ZN(n5561) );
  INV_X1 U6579 ( .A(n5559), .ZN(n5558) );
  INV_X1 U6580 ( .A(SI_2_), .ZN(n10217) );
  NAND2_X1 U6581 ( .A1(n5558), .A2(n10217), .ZN(n5560) );
  NAND2_X1 U6582 ( .A1(n5559), .A2(SI_2_), .ZN(n5579) );
  NAND2_X1 U6583 ( .A1(n5560), .A2(n5579), .ZN(n5562) );
  NAND2_X1 U6584 ( .A1(n5561), .A2(n5562), .ZN(n5565) );
  INV_X1 U6585 ( .A(n5562), .ZN(n5563) );
  NAND2_X1 U6586 ( .A1(n5565), .A2(n5580), .ZN(n6791) );
  OR2_X1 U6587 ( .A1(n5609), .A2(n6791), .ZN(n5571) );
  OR2_X1 U6588 ( .A1(n5965), .A2(n5556), .ZN(n5570) );
  INV_X1 U6589 ( .A(P2_IR_REG_31__SCAN_IN), .ZN(n9484) );
  OR2_X1 U6590 ( .A1(n5566), .A2(n9484), .ZN(n5568) );
  INV_X1 U6591 ( .A(P2_IR_REG_2__SCAN_IN), .ZN(n5567) );
  NAND2_X1 U6592 ( .A1(n5568), .A2(n5567), .ZN(n5577) );
  OAI21_X1 U6593 ( .B1(n5568), .B2(n5567), .A(n5577), .ZN(n10435) );
  OR2_X1 U6594 ( .A1(n6643), .A2(n10435), .ZN(n5569) );
  NAND2_X1 U6595 ( .A1(n5572), .A2(n7220), .ZN(n5573) );
  NAND2_X1 U6596 ( .A1(n5576), .A2(n5573), .ZN(n7088) );
  INV_X1 U6597 ( .A(n7088), .ZN(n5574) );
  NAND2_X1 U6598 ( .A1(n5575), .A2(n5574), .ZN(n7223) );
  NAND2_X1 U6599 ( .A1(n7223), .A2(n5576), .ZN(n5600) );
  NAND2_X1 U6600 ( .A1(n5577), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5578) );
  XNOR2_X1 U6601 ( .A(n5578), .B(P2_IR_REG_3__SCAN_IN), .ZN(n10448) );
  AOI22_X1 U6602 ( .A1(n5945), .A2(P1_DATAO_REG_3__SCAN_IN), .B1(n6433), .B2(
        n10448), .ZN(n5588) );
  NAND2_X1 U6603 ( .A1(n5580), .A2(n5579), .ZN(n5585) );
  NAND2_X1 U6604 ( .A1(n5581), .A2(SI_3_), .ZN(n5601) );
  INV_X1 U6605 ( .A(SI_3_), .ZN(n5582) );
  OR2_X1 U6606 ( .A1(n5585), .A2(n5584), .ZN(n5586) );
  AND2_X1 U6607 ( .A1(n5602), .A2(n5586), .ZN(n6770) );
  NAND2_X1 U6608 ( .A1(n6770), .A2(n8726), .ZN(n5587) );
  XNOR2_X1 U6609 ( .A(n6974), .B(n6115), .ZN(n5596) );
  NAND2_X1 U6610 ( .A1(n5589), .A2(P2_REG2_REG_3__SCAN_IN), .ZN(n5595) );
  NAND2_X1 U6611 ( .A1(n5590), .A2(P2_REG1_REG_3__SCAN_IN), .ZN(n5594) );
  NAND2_X1 U6612 ( .A1(n6419), .A2(P2_REG0_REG_3__SCAN_IN), .ZN(n5593) );
  NAND2_X1 U6613 ( .A1(n5591), .A2(n7216), .ZN(n5592) );
  AND2_X1 U6614 ( .A1(n5621), .A2(n6259), .ZN(n5597) );
  NAND2_X1 U6615 ( .A1(n5596), .A2(n5597), .ZN(n5622) );
  INV_X1 U6616 ( .A(n5596), .ZN(n7369) );
  INV_X1 U6617 ( .A(n5597), .ZN(n5598) );
  NAND2_X1 U6618 ( .A1(n7369), .A2(n5598), .ZN(n5599) );
  AND2_X1 U6619 ( .A1(n5622), .A2(n5599), .ZN(n7221) );
  NAND2_X1 U6620 ( .A1(n5600), .A2(n7221), .ZN(n7224) );
  NAND2_X1 U6621 ( .A1(n5603), .A2(SI_4_), .ZN(n5627) );
  INV_X1 U6622 ( .A(n5603), .ZN(n5604) );
  NAND2_X1 U6623 ( .A1(n5604), .A2(n10215), .ZN(n5605) );
  NAND2_X1 U6624 ( .A1(n5607), .A2(n5606), .ZN(n5628) );
  NAND2_X1 U6625 ( .A1(n5628), .A2(n5608), .ZN(n6841) );
  NAND2_X1 U6626 ( .A1(n5610), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5611) );
  MUX2_X1 U6627 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5611), .S(
        P2_IR_REG_4__SCAN_IN), .Z(n5613) );
  AND2_X1 U6628 ( .A1(n5613), .A2(n5612), .ZN(n6659) );
  AOI22_X1 U6629 ( .A1(n5945), .A2(P1_DATAO_REG_4__SCAN_IN), .B1(n6433), .B2(
        n6659), .ZN(n5614) );
  XNOR2_X1 U6630 ( .A(n7301), .B(n5615), .ZN(n7418) );
  NAND2_X1 U6631 ( .A1(n6419), .A2(P2_REG0_REG_4__SCAN_IN), .ZN(n5620) );
  NAND2_X1 U6632 ( .A1(n5589), .A2(P2_REG2_REG_4__SCAN_IN), .ZN(n5619) );
  INV_X1 U6633 ( .A(n5640), .ZN(n5641) );
  OAI21_X1 U6634 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(P2_REG3_REG_4__SCAN_IN), 
        .A(n5641), .ZN(n7372) );
  INV_X1 U6635 ( .A(n7372), .ZN(n5616) );
  NAND2_X1 U6636 ( .A1(n5591), .A2(n5616), .ZN(n5618) );
  NAND2_X1 U6637 ( .A1(n5590), .A2(P2_REG1_REG_4__SCAN_IN), .ZN(n5617) );
  OR2_X1 U6638 ( .A1(n7217), .A2(n5747), .ZN(n5624) );
  XNOR2_X1 U6639 ( .A(n7418), .B(n5624), .ZN(n7368) );
  AND2_X1 U6640 ( .A1(n7368), .A2(n5622), .ZN(n5623) );
  INV_X1 U6641 ( .A(n7418), .ZN(n5625) );
  NAND2_X1 U6642 ( .A1(n5625), .A2(n5624), .ZN(n5626) );
  NAND2_X1 U6643 ( .A1(n5628), .A2(n5627), .ZN(n5633) );
  INV_X1 U6644 ( .A(n5629), .ZN(n5630) );
  INV_X1 U6645 ( .A(SI_5_), .ZN(n10216) );
  NAND2_X1 U6646 ( .A1(n5630), .A2(n10216), .ZN(n5631) );
  OR2_X1 U6647 ( .A1(n5633), .A2(n5632), .ZN(n5634) );
  NAND2_X1 U6648 ( .A1(n5612), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5635) );
  MUX2_X1 U6649 ( .A(P2_IR_REG_31__SCAN_IN), .B(n5635), .S(
        P2_IR_REG_5__SCAN_IN), .Z(n5637) );
  INV_X1 U6650 ( .A(n5678), .ZN(n5636) );
  AOI22_X1 U6651 ( .A1(n5945), .A2(P1_DATAO_REG_5__SCAN_IN), .B1(n6433), .B2(
        n10462), .ZN(n5638) );
  XNOR2_X1 U6652 ( .A(n10546), .B(n6115), .ZN(n5647) );
  NAND2_X1 U6653 ( .A1(n5589), .A2(P2_REG2_REG_5__SCAN_IN), .ZN(n5646) );
  NAND2_X1 U6654 ( .A1(n6419), .A2(P2_REG0_REG_5__SCAN_IN), .ZN(n5645) );
  INV_X1 U6655 ( .A(P2_REG3_REG_5__SCAN_IN), .ZN(n10251) );
  NAND2_X1 U6656 ( .A1(n5641), .A2(n10251), .ZN(n5642) );
  AND2_X1 U6657 ( .A1(n5685), .A2(n5642), .ZN(n7415) );
  NAND2_X1 U6658 ( .A1(n5591), .A2(n7415), .ZN(n5644) );
  NAND2_X1 U6659 ( .A1(n5590), .A2(P2_REG1_REG_5__SCAN_IN), .ZN(n5643) );
  NAND4_X1 U6660 ( .A1(n5646), .A2(n5645), .A3(n5644), .A4(n5643), .ZN(n7374)
         );
  NAND2_X1 U6661 ( .A1(n5621), .A2(n7374), .ZN(n5648) );
  XNOR2_X1 U6662 ( .A(n5647), .B(n5648), .ZN(n7420) );
  INV_X1 U6663 ( .A(n5647), .ZN(n7243) );
  NAND2_X1 U6664 ( .A1(n5651), .A2(SI_6_), .ZN(n5669) );
  INV_X1 U6665 ( .A(n5651), .ZN(n5652) );
  NAND2_X1 U6666 ( .A1(n5652), .A2(n10213), .ZN(n5653) );
  OR2_X1 U6667 ( .A1(n5655), .A2(n5654), .ZN(n5656) );
  NAND2_X1 U6668 ( .A1(n5670), .A2(n5656), .ZN(n7128) );
  OR2_X1 U6669 ( .A1(n7128), .A2(n5609), .ZN(n5659) );
  OR2_X1 U6670 ( .A1(n5678), .A2(n9484), .ZN(n5657) );
  XNOR2_X1 U6671 ( .A(n5657), .B(P2_IR_REG_6__SCAN_IN), .ZN(n10477) );
  AOI22_X1 U6672 ( .A1(n5945), .A2(P1_DATAO_REG_6__SCAN_IN), .B1(n6433), .B2(
        n10477), .ZN(n5658) );
  NAND2_X1 U6673 ( .A1(n5659), .A2(n5658), .ZN(n8784) );
  XNOR2_X1 U6674 ( .A(n8784), .B(n5615), .ZN(n5665) );
  NAND2_X1 U6675 ( .A1(n6419), .A2(P2_REG0_REG_6__SCAN_IN), .ZN(n5663) );
  NAND2_X1 U6676 ( .A1(n5589), .A2(P2_REG2_REG_6__SCAN_IN), .ZN(n5662) );
  XNOR2_X1 U6677 ( .A(n5685), .B(P2_REG3_REG_6__SCAN_IN), .ZN(n7240) );
  NAND2_X1 U6678 ( .A1(n5591), .A2(n7240), .ZN(n5661) );
  NAND2_X1 U6679 ( .A1(n6418), .A2(P2_REG1_REG_6__SCAN_IN), .ZN(n5660) );
  NAND4_X1 U6680 ( .A1(n5663), .A2(n5662), .A3(n5661), .A4(n5660), .ZN(n8781)
         );
  NAND2_X1 U6681 ( .A1(n5621), .A2(n8781), .ZN(n5666) );
  XNOR2_X1 U6682 ( .A(n5665), .B(n5666), .ZN(n7244) );
  NAND2_X1 U6683 ( .A1(n5664), .A2(n7244), .ZN(n7250) );
  INV_X1 U6684 ( .A(n5665), .ZN(n5667) );
  NAND2_X1 U6685 ( .A1(n5667), .A2(n5666), .ZN(n5668) );
  NAND2_X1 U6686 ( .A1(n7250), .A2(n5668), .ZN(n7159) );
  MUX2_X1 U6687 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(P2_DATAO_REG_7__SCAN_IN), 
        .S(n8387), .Z(n5671) );
  NAND2_X1 U6688 ( .A1(n5671), .A2(SI_7_), .ZN(n5696) );
  INV_X1 U6689 ( .A(n5671), .ZN(n5672) );
  NAND2_X1 U6690 ( .A1(n5672), .A2(n10210), .ZN(n5673) );
  OR2_X1 U6691 ( .A1(n5675), .A2(n5674), .ZN(n5676) );
  NAND2_X1 U6692 ( .A1(n5675), .A2(n5674), .ZN(n5697) );
  NAND2_X1 U6693 ( .A1(n5676), .A2(n5697), .ZN(n7195) );
  OR2_X1 U6694 ( .A1(n7195), .A2(n5609), .ZN(n5681) );
  NAND2_X1 U6695 ( .A1(n5678), .A2(n5677), .ZN(n5698) );
  NAND2_X1 U6696 ( .A1(n5698), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5679) );
  XNOR2_X1 U6697 ( .A(n5679), .B(P2_IR_REG_7__SCAN_IN), .ZN(n6670) );
  AOI22_X1 U6698 ( .A1(n5945), .A2(P1_DATAO_REG_7__SCAN_IN), .B1(n6433), .B2(
        n6670), .ZN(n5680) );
  NAND2_X1 U6699 ( .A1(n5681), .A2(n5680), .ZN(n8789) );
  XNOR2_X1 U6700 ( .A(n8789), .B(n5615), .ZN(n5691) );
  NAND2_X1 U6701 ( .A1(n6419), .A2(P2_REG0_REG_7__SCAN_IN), .ZN(n5690) );
  NAND2_X1 U6702 ( .A1(n5589), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n5689) );
  NAND2_X1 U6703 ( .A1(P2_REG3_REG_7__SCAN_IN), .A2(P2_REG3_REG_6__SCAN_IN), 
        .ZN(n5683) );
  INV_X1 U6704 ( .A(n5702), .ZN(n5703) );
  INV_X1 U6705 ( .A(P2_REG3_REG_6__SCAN_IN), .ZN(n5684) );
  OAI21_X1 U6706 ( .B1(n5685), .B2(n5684), .A(n10114), .ZN(n5686) );
  AND2_X1 U6707 ( .A1(n5703), .A2(n5686), .ZN(n7484) );
  NAND2_X1 U6708 ( .A1(n5591), .A2(n7484), .ZN(n5688) );
  NAND2_X1 U6709 ( .A1(n6418), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n5687) );
  NAND4_X1 U6710 ( .A1(n5690), .A2(n5689), .A3(n5688), .A4(n5687), .ZN(n9065)
         );
  AND2_X1 U6711 ( .A1(n5621), .A2(n9065), .ZN(n5692) );
  NAND2_X1 U6712 ( .A1(n5691), .A2(n5692), .ZN(n5695) );
  INV_X1 U6713 ( .A(n5691), .ZN(n8969) );
  INV_X1 U6714 ( .A(n5692), .ZN(n5693) );
  NAND2_X1 U6715 ( .A1(n8969), .A2(n5693), .ZN(n5694) );
  NAND2_X1 U6716 ( .A1(n5695), .A2(n5694), .ZN(n7160) );
  NAND2_X1 U6717 ( .A1(n5697), .A2(n5696), .ZN(n5715) );
  XNOR2_X1 U6718 ( .A(n5715), .B(n5714), .ZN(n7440) );
  NAND2_X1 U6719 ( .A1(n7440), .A2(n8726), .ZN(n5701) );
  NAND2_X1 U6720 ( .A1(n5716), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5699) );
  XNOR2_X1 U6721 ( .A(n5699), .B(P2_IR_REG_8__SCAN_IN), .ZN(n6707) );
  AOI22_X1 U6722 ( .A1(n5945), .A2(P1_DATAO_REG_8__SCAN_IN), .B1(n6433), .B2(
        n6707), .ZN(n5700) );
  NAND2_X1 U6723 ( .A1(n5701), .A2(n5700), .ZN(n8975) );
  XNOR2_X1 U6724 ( .A(n8975), .B(n5615), .ZN(n5709) );
  NAND2_X1 U6725 ( .A1(n5589), .A2(P2_REG2_REG_8__SCAN_IN), .ZN(n5708) );
  NAND2_X1 U6726 ( .A1(n6418), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n5707) );
  NAND2_X1 U6727 ( .A1(n5702), .A2(P2_REG3_REG_8__SCAN_IN), .ZN(n5720) );
  INV_X1 U6728 ( .A(P2_REG3_REG_8__SCAN_IN), .ZN(n10127) );
  NAND2_X1 U6729 ( .A1(n5703), .A2(n10127), .ZN(n5704) );
  AND2_X1 U6730 ( .A1(n5720), .A2(n5704), .ZN(n8974) );
  NAND2_X1 U6731 ( .A1(n5591), .A2(n8974), .ZN(n5706) );
  NAND2_X1 U6732 ( .A1(n6419), .A2(P2_REG0_REG_8__SCAN_IN), .ZN(n5705) );
  NOR2_X1 U6733 ( .A1(n7478), .A2(n5747), .ZN(n5710) );
  NAND2_X1 U6734 ( .A1(n5709), .A2(n5710), .ZN(n5726) );
  INV_X1 U6735 ( .A(n5709), .ZN(n9018) );
  INV_X1 U6736 ( .A(n5710), .ZN(n5711) );
  NAND2_X1 U6737 ( .A1(n9018), .A2(n5711), .ZN(n5712) );
  AND2_X1 U6738 ( .A1(n5726), .A2(n5712), .ZN(n8966) );
  XNOR2_X1 U6739 ( .A(n5733), .B(n5732), .ZN(n7511) );
  NAND2_X1 U6740 ( .A1(n7511), .A2(n8726), .ZN(n5718) );
  NAND2_X1 U6741 ( .A1(n5787), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5737) );
  XNOR2_X1 U6742 ( .A(n5737), .B(P2_IR_REG_9__SCAN_IN), .ZN(n6728) );
  AOI22_X1 U6743 ( .A1(n5945), .A2(P1_DATAO_REG_9__SCAN_IN), .B1(n6433), .B2(
        n6728), .ZN(n5717) );
  XNOR2_X1 U6744 ( .A(n10605), .B(n6115), .ZN(n5730) );
  NAND2_X1 U6745 ( .A1(n5589), .A2(P2_REG2_REG_9__SCAN_IN), .ZN(n5725) );
  NAND2_X1 U6746 ( .A1(n6418), .A2(P2_REG1_REG_9__SCAN_IN), .ZN(n5724) );
  NAND2_X1 U6747 ( .A1(n5720), .A2(n5719), .ZN(n5721) );
  AND2_X1 U6748 ( .A1(n5741), .A2(n5721), .ZN(n9011) );
  NAND2_X1 U6749 ( .A1(n5591), .A2(n9011), .ZN(n5723) );
  NAND2_X1 U6750 ( .A1(n6419), .A2(P2_REG0_REG_9__SCAN_IN), .ZN(n5722) );
  NOR2_X1 U6751 ( .A1(n7582), .A2(n5747), .ZN(n5728) );
  XNOR2_X1 U6752 ( .A(n5730), .B(n5728), .ZN(n9019) );
  NAND2_X1 U6753 ( .A1(n8971), .A2(n5727), .ZN(n9008) );
  INV_X1 U6754 ( .A(n5728), .ZN(n5729) );
  NAND2_X1 U6755 ( .A1(n5730), .A2(n5729), .ZN(n5731) );
  NAND2_X1 U6756 ( .A1(n9008), .A2(n5731), .ZN(n7571) );
  INV_X1 U6757 ( .A(n5734), .ZN(n5735) );
  NAND2_X1 U6758 ( .A1(n5735), .A2(n10203), .ZN(n5755) );
  NAND2_X1 U6759 ( .A1(n5759), .A2(n5755), .ZN(n5736) );
  XNOR2_X1 U6760 ( .A(n5753), .B(n10191), .ZN(n5757) );
  XNOR2_X1 U6761 ( .A(n5736), .B(n5757), .ZN(n7644) );
  NAND2_X1 U6762 ( .A1(n7644), .A2(n8726), .ZN(n5740) );
  NAND2_X1 U6763 ( .A1(n5737), .A2(n5785), .ZN(n5738) );
  NAND2_X1 U6764 ( .A1(n5738), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5765) );
  XNOR2_X1 U6765 ( .A(n5765), .B(P2_IR_REG_10__SCAN_IN), .ZN(n6863) );
  AOI22_X1 U6766 ( .A1(n5945), .A2(P1_DATAO_REG_10__SCAN_IN), .B1(n6433), .B2(
        n6863), .ZN(n5739) );
  NAND2_X1 U6767 ( .A1(n5740), .A2(n5739), .ZN(n7590) );
  XNOR2_X1 U6768 ( .A(n7590), .B(n5615), .ZN(n5748) );
  NAND2_X1 U6769 ( .A1(n6419), .A2(P2_REG0_REG_10__SCAN_IN), .ZN(n5746) );
  NAND2_X1 U6770 ( .A1(n5589), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n5745) );
  INV_X1 U6771 ( .A(n5770), .ZN(n5772) );
  NAND2_X1 U6772 ( .A1(n5741), .A2(n6714), .ZN(n5742) );
  AND2_X1 U6773 ( .A1(n5772), .A2(n5742), .ZN(n7589) );
  NAND2_X1 U6774 ( .A1(n5591), .A2(n7589), .ZN(n5744) );
  NAND2_X1 U6775 ( .A1(n6418), .A2(P2_REG1_REG_10__SCAN_IN), .ZN(n5743) );
  NOR2_X1 U6776 ( .A1(n9014), .A2(n5747), .ZN(n5749) );
  NAND2_X1 U6777 ( .A1(n5748), .A2(n5749), .ZN(n5752) );
  INV_X1 U6778 ( .A(n5748), .ZN(n7541) );
  INV_X1 U6779 ( .A(n5749), .ZN(n5750) );
  NAND2_X1 U6780 ( .A1(n7541), .A2(n5750), .ZN(n5751) );
  NAND2_X1 U6781 ( .A1(n5752), .A2(n5751), .ZN(n7572) );
  INV_X1 U6782 ( .A(n5753), .ZN(n5754) );
  NAND2_X1 U6783 ( .A1(n5754), .A2(n10191), .ZN(n5756) );
  INV_X1 U6784 ( .A(n5756), .ZN(n5758) );
  NAND2_X1 U6785 ( .A1(n5762), .A2(n5761), .ZN(n5763) );
  NAND2_X1 U6786 ( .A1(n5783), .A2(n5763), .ZN(n7650) );
  OR2_X1 U6787 ( .A1(n7650), .A2(n5609), .ZN(n5769) );
  NAND2_X1 U6788 ( .A1(n5765), .A2(n5764), .ZN(n5766) );
  NAND2_X1 U6789 ( .A1(n5766), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5767) );
  XNOR2_X1 U6790 ( .A(n5767), .B(P2_IR_REG_11__SCAN_IN), .ZN(n6868) );
  AOI22_X1 U6791 ( .A1(n5945), .A2(P1_DATAO_REG_11__SCAN_IN), .B1(n6433), .B2(
        n6868), .ZN(n5768) );
  XNOR2_X1 U6792 ( .A(n7693), .B(n5615), .ZN(n5778) );
  NAND2_X1 U6793 ( .A1(n6419), .A2(P2_REG0_REG_11__SCAN_IN), .ZN(n5777) );
  NAND2_X1 U6794 ( .A1(n5589), .A2(P2_REG2_REG_11__SCAN_IN), .ZN(n5776) );
  INV_X1 U6795 ( .A(n5791), .ZN(n5792) );
  INV_X1 U6796 ( .A(P2_REG3_REG_11__SCAN_IN), .ZN(n5771) );
  NAND2_X1 U6797 ( .A1(n5772), .A2(n5771), .ZN(n5773) );
  AND2_X1 U6798 ( .A1(n5792), .A2(n5773), .ZN(n7545) );
  NAND2_X1 U6799 ( .A1(n5591), .A2(n7545), .ZN(n5775) );
  NAND2_X1 U6800 ( .A1(n6418), .A2(P2_REG1_REG_11__SCAN_IN), .ZN(n5774) );
  NOR2_X1 U6801 ( .A1(n7694), .A2(n5747), .ZN(n5779) );
  NAND2_X1 U6802 ( .A1(n5778), .A2(n5779), .ZN(n5798) );
  INV_X1 U6803 ( .A(n5778), .ZN(n7629) );
  INV_X1 U6804 ( .A(n5779), .ZN(n5780) );
  NAND2_X1 U6805 ( .A1(n7629), .A2(n5780), .ZN(n5781) );
  AND2_X1 U6806 ( .A1(n5798), .A2(n5781), .ZN(n7539) );
  MUX2_X1 U6807 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(P2_DATAO_REG_12__SCAN_IN), 
        .S(n8387), .Z(n5804) );
  XNOR2_X1 U6808 ( .A(n5808), .B(n5807), .ZN(n7729) );
  NAND2_X1 U6809 ( .A1(n7729), .A2(n8726), .ZN(n5790) );
  INV_X1 U6810 ( .A(P2_IR_REG_11__SCAN_IN), .ZN(n5784) );
  NAND3_X1 U6811 ( .A1(n5785), .A2(n5764), .A3(n5784), .ZN(n5786) );
  NOR2_X1 U6812 ( .A1(n5787), .A2(n5786), .ZN(n5811) );
  OR2_X1 U6813 ( .A1(n5811), .A2(n9484), .ZN(n5788) );
  XNOR2_X1 U6814 ( .A(n5788), .B(P2_IR_REG_12__SCAN_IN), .ZN(n7253) );
  AOI22_X1 U6815 ( .A1(n5945), .A2(P1_DATAO_REG_12__SCAN_IN), .B1(n6433), .B2(
        n7253), .ZN(n5789) );
  XNOR2_X1 U6816 ( .A(n8805), .B(n6115), .ZN(n5802) );
  INV_X1 U6817 ( .A(P2_REG3_REG_12__SCAN_IN), .ZN(n10238) );
  NAND2_X1 U6818 ( .A1(n5792), .A2(n10238), .ZN(n5793) );
  AND2_X1 U6819 ( .A1(n5816), .A2(n5793), .ZN(n7701) );
  NAND2_X1 U6820 ( .A1(n5591), .A2(n7701), .ZN(n5797) );
  NAND2_X1 U6821 ( .A1(n5589), .A2(P2_REG2_REG_12__SCAN_IN), .ZN(n5796) );
  NAND2_X1 U6822 ( .A1(n6418), .A2(P2_REG1_REG_12__SCAN_IN), .ZN(n5795) );
  NAND2_X1 U6823 ( .A1(n6419), .A2(P2_REG0_REG_12__SCAN_IN), .ZN(n5794) );
  NOR2_X1 U6824 ( .A1(n8804), .A2(n5747), .ZN(n5800) );
  XNOR2_X1 U6825 ( .A(n5802), .B(n5800), .ZN(n7632) );
  AND2_X1 U6826 ( .A1(n7632), .A2(n5798), .ZN(n5799) );
  NAND2_X1 U6827 ( .A1(n7542), .A2(n5799), .ZN(n7631) );
  INV_X1 U6828 ( .A(n5800), .ZN(n5801) );
  NAND2_X1 U6829 ( .A1(n5802), .A2(n5801), .ZN(n5803) );
  NAND2_X1 U6830 ( .A1(n7631), .A2(n5803), .ZN(n10289) );
  INV_X1 U6831 ( .A(n5804), .ZN(n5806) );
  INV_X1 U6832 ( .A(SI_12_), .ZN(n5805) );
  MUX2_X1 U6833 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(P2_DATAO_REG_13__SCAN_IN), 
        .S(n8387), .Z(n5826) );
  XNOR2_X1 U6834 ( .A(n5829), .B(n5828), .ZN(n7851) );
  NAND2_X1 U6835 ( .A1(n7851), .A2(n8726), .ZN(n5814) );
  INV_X1 U6836 ( .A(P2_IR_REG_12__SCAN_IN), .ZN(n5810) );
  NAND2_X1 U6837 ( .A1(n5811), .A2(n5810), .ZN(n5812) );
  NAND2_X1 U6838 ( .A1(n5812), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5836) );
  XNOR2_X1 U6839 ( .A(n5836), .B(P2_IR_REG_13__SCAN_IN), .ZN(n7395) );
  AOI22_X1 U6840 ( .A1(n5945), .A2(P1_DATAO_REG_13__SCAN_IN), .B1(n6433), .B2(
        n7395), .ZN(n5813) );
  XNOR2_X1 U6841 ( .A(n10294), .B(n5615), .ZN(n5822) );
  NAND2_X1 U6842 ( .A1(n6419), .A2(P2_REG0_REG_13__SCAN_IN), .ZN(n5821) );
  NAND2_X1 U6843 ( .A1(n5589), .A2(P2_REG2_REG_13__SCAN_IN), .ZN(n5820) );
  INV_X1 U6844 ( .A(P2_REG3_REG_13__SCAN_IN), .ZN(n5815) );
  NAND2_X1 U6845 ( .A1(n5816), .A2(n5815), .ZN(n5817) );
  AND2_X1 U6846 ( .A1(n5843), .A2(n5817), .ZN(n10283) );
  NAND2_X1 U6847 ( .A1(n5591), .A2(n10283), .ZN(n5819) );
  NAND2_X1 U6848 ( .A1(n5590), .A2(P2_REG1_REG_13__SCAN_IN), .ZN(n5818) );
  NOR2_X1 U6849 ( .A1(n7914), .A2(n5747), .ZN(n5823) );
  NAND2_X1 U6850 ( .A1(n5822), .A2(n5823), .ZN(n5849) );
  INV_X1 U6851 ( .A(n5822), .ZN(n7898) );
  INV_X1 U6852 ( .A(n5823), .ZN(n5824) );
  NAND2_X1 U6853 ( .A1(n7898), .A2(n5824), .ZN(n5825) );
  NAND2_X1 U6854 ( .A1(n5849), .A2(n5825), .ZN(n10290) );
  MUX2_X1 U6855 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(P2_DATAO_REG_14__SCAN_IN), 
        .S(n8387), .Z(n5830) );
  INV_X1 U6856 ( .A(n5830), .ZN(n5831) );
  INV_X1 U6857 ( .A(SI_14_), .ZN(n10085) );
  NAND2_X1 U6858 ( .A1(n5831), .A2(n10085), .ZN(n5832) );
  NAND2_X1 U6859 ( .A1(n5853), .A2(n5832), .ZN(n5833) );
  NAND2_X1 U6860 ( .A1(n4871), .A2(n5833), .ZN(n5834) );
  INV_X1 U6861 ( .A(P2_IR_REG_13__SCAN_IN), .ZN(n5835) );
  NAND2_X1 U6862 ( .A1(n5836), .A2(n5835), .ZN(n5837) );
  NAND2_X1 U6863 ( .A1(n5837), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5839) );
  NAND2_X1 U6864 ( .A1(n5839), .A2(n5838), .ZN(n5857) );
  OR2_X1 U6865 ( .A1(n5839), .A2(n5838), .ZN(n5840) );
  AOI22_X1 U6866 ( .A1(n6433), .A2(n7680), .B1(n5945), .B2(
        P1_DATAO_REG_14__SCAN_IN), .ZN(n5841) );
  NAND2_X1 U6867 ( .A1(n5589), .A2(P2_REG2_REG_14__SCAN_IN), .ZN(n5848) );
  NAND2_X1 U6868 ( .A1(n6419), .A2(P2_REG0_REG_14__SCAN_IN), .ZN(n5847) );
  INV_X1 U6869 ( .A(P2_REG3_REG_14__SCAN_IN), .ZN(n5842) );
  NAND2_X1 U6870 ( .A1(n5843), .A2(n5842), .ZN(n5844) );
  AND2_X1 U6871 ( .A1(n5862), .A2(n5844), .ZN(n7917) );
  NAND2_X1 U6872 ( .A1(n5591), .A2(n7917), .ZN(n5846) );
  NAND2_X1 U6873 ( .A1(n5590), .A2(P2_REG1_REG_14__SCAN_IN), .ZN(n5845) );
  NOR2_X1 U6874 ( .A1(n9060), .A2(n5747), .ZN(n5851) );
  XNOR2_X1 U6875 ( .A(n8311), .B(n5851), .ZN(n7907) );
  INV_X1 U6876 ( .A(n5851), .ZN(n5852) );
  MUX2_X1 U6877 ( .A(n6894), .B(n6893), .S(n8387), .Z(n5871) );
  INV_X1 U6878 ( .A(n5871), .ZN(n5855) );
  XNOR2_X1 U6879 ( .A(n5855), .B(SI_15_), .ZN(n5856) );
  XNOR2_X1 U6880 ( .A(n5873), .B(n5856), .ZN(n8006) );
  NAND2_X1 U6881 ( .A1(n8006), .A2(n8726), .ZN(n5860) );
  NAND2_X1 U6882 ( .A1(n5857), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5858) );
  XNOR2_X1 U6883 ( .A(n5858), .B(P2_IR_REG_15__SCAN_IN), .ZN(n7810) );
  AOI22_X1 U6884 ( .A1(n7810), .A2(n6433), .B1(n5945), .B2(
        P1_DATAO_REG_15__SCAN_IN), .ZN(n5859) );
  XNOR2_X1 U6885 ( .A(n8310), .B(n6115), .ZN(n7892) );
  NAND2_X1 U6886 ( .A1(n6419), .A2(P2_REG0_REG_15__SCAN_IN), .ZN(n5867) );
  NAND2_X1 U6887 ( .A1(n5589), .A2(P2_REG2_REG_15__SCAN_IN), .ZN(n5866) );
  INV_X1 U6888 ( .A(P2_REG3_REG_15__SCAN_IN), .ZN(n5861) );
  INV_X1 U6889 ( .A(n5879), .ZN(n5880) );
  NAND2_X1 U6890 ( .A1(n5862), .A2(n5861), .ZN(n5863) );
  AND2_X1 U6891 ( .A1(n5880), .A2(n5863), .ZN(n8306) );
  NAND2_X1 U6892 ( .A1(n5591), .A2(n8306), .ZN(n5865) );
  NAND2_X1 U6893 ( .A1(n6418), .A2(P2_REG1_REG_15__SCAN_IN), .ZN(n5864) );
  NOR2_X1 U6894 ( .A1(n7982), .A2(n5747), .ZN(n5868) );
  INV_X1 U6895 ( .A(n5868), .ZN(n5869) );
  NAND2_X1 U6896 ( .A1(n7892), .A2(n5869), .ZN(n5870) );
  NAND2_X1 U6897 ( .A1(n8315), .A2(n5870), .ZN(n5886) );
  NOR2_X1 U6898 ( .A1(n5871), .A2(n10192), .ZN(n5872) );
  MUX2_X1 U6899 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(P2_DATAO_REG_16__SCAN_IN), 
        .S(n8387), .Z(n5891) );
  INV_X1 U6900 ( .A(SI_16_), .ZN(n5874) );
  XNOR2_X1 U6901 ( .A(n5894), .B(n5893), .ZN(n8042) );
  NAND2_X1 U6902 ( .A1(n8042), .A2(n8726), .ZN(n5878) );
  NOR2_X1 U6903 ( .A1(n4859), .A2(n9484), .ZN(n5875) );
  MUX2_X1 U6904 ( .A(n9484), .B(n5875), .S(P2_IR_REG_16__SCAN_IN), .Z(n5876)
         );
  OR2_X1 U6905 ( .A1(n5876), .A2(n5903), .ZN(n7827) );
  INV_X1 U6906 ( .A(n7827), .ZN(n7973) );
  AOI22_X1 U6907 ( .A1(n5945), .A2(P1_DATAO_REG_16__SCAN_IN), .B1(n6433), .B2(
        n7973), .ZN(n5877) );
  XNOR2_X1 U6908 ( .A(n9124), .B(n6115), .ZN(n5889) );
  NAND2_X1 U6909 ( .A1(n5589), .A2(P2_REG2_REG_16__SCAN_IN), .ZN(n5885) );
  NAND2_X1 U6910 ( .A1(n5879), .A2(P2_REG3_REG_16__SCAN_IN), .ZN(n5912) );
  INV_X1 U6911 ( .A(P2_REG3_REG_16__SCAN_IN), .ZN(n10248) );
  NAND2_X1 U6912 ( .A1(n5880), .A2(n10248), .ZN(n5881) );
  AND2_X1 U6913 ( .A1(n5912), .A2(n5881), .ZN(n7888) );
  NAND2_X1 U6914 ( .A1(n5591), .A2(n7888), .ZN(n5884) );
  NAND2_X1 U6915 ( .A1(n6419), .A2(P2_REG0_REG_16__SCAN_IN), .ZN(n5883) );
  NAND2_X1 U6916 ( .A1(n6418), .A2(P2_REG1_REG_16__SCAN_IN), .ZN(n5882) );
  NOR2_X1 U6917 ( .A1(n9058), .A2(n5542), .ZN(n5887) );
  XNOR2_X1 U6918 ( .A(n5889), .B(n5887), .ZN(n7891) );
  INV_X1 U6919 ( .A(n5887), .ZN(n5888) );
  NAND2_X1 U6920 ( .A1(n5889), .A2(n5888), .ZN(n5890) );
  NOR2_X1 U6921 ( .A1(n5891), .A2(SI_16_), .ZN(n5892) );
  AOI21_X1 U6922 ( .B1(n5894), .B2(n5893), .A(n5892), .ZN(n5899) );
  MUX2_X1 U6923 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(P2_DATAO_REG_17__SCAN_IN), 
        .S(n8387), .Z(n5895) );
  NAND2_X1 U6924 ( .A1(n5895), .A2(SI_17_), .ZN(n5921) );
  INV_X1 U6925 ( .A(n5895), .ZN(n5896) );
  INV_X1 U6926 ( .A(SI_17_), .ZN(n10188) );
  NAND2_X1 U6927 ( .A1(n5896), .A2(n10188), .ZN(n5897) );
  NAND2_X1 U6928 ( .A1(n5921), .A2(n5897), .ZN(n5900) );
  INV_X1 U6929 ( .A(n5900), .ZN(n5898) );
  NAND2_X1 U6930 ( .A1(n5899), .A2(n5898), .ZN(n5922) );
  INV_X1 U6931 ( .A(n5899), .ZN(n5901) );
  NAND2_X1 U6932 ( .A1(n5901), .A2(n5900), .ZN(n5902) );
  NAND2_X1 U6933 ( .A1(n5922), .A2(n5902), .ZN(n8135) );
  NOR2_X1 U6934 ( .A1(n5903), .A2(n9484), .ZN(n5904) );
  MUX2_X1 U6935 ( .A(n9484), .B(n5904), .S(P2_IR_REG_17__SCAN_IN), .Z(n5906)
         );
  INV_X1 U6936 ( .A(n5929), .ZN(n5905) );
  OR2_X1 U6937 ( .A1(n5906), .A2(n5905), .ZN(n9081) );
  INV_X1 U6938 ( .A(n9081), .ZN(n9073) );
  AOI22_X1 U6939 ( .A1(n5945), .A2(P1_DATAO_REG_17__SCAN_IN), .B1(n6433), .B2(
        n9073), .ZN(n5907) );
  XNOR2_X1 U6940 ( .A(n9457), .B(n6115), .ZN(n5917) );
  NAND2_X1 U6941 ( .A1(n5589), .A2(P2_REG2_REG_17__SCAN_IN), .ZN(n5910) );
  NAND2_X1 U6942 ( .A1(n6419), .A2(P2_REG0_REG_17__SCAN_IN), .ZN(n5909) );
  AND2_X1 U6943 ( .A1(n5910), .A2(n5909), .ZN(n5916) );
  INV_X1 U6944 ( .A(P2_REG3_REG_17__SCAN_IN), .ZN(n5911) );
  NAND2_X1 U6945 ( .A1(n5912), .A2(n5911), .ZN(n5913) );
  AND2_X1 U6946 ( .A1(n5933), .A2(n5913), .ZN(n9353) );
  NAND2_X1 U6947 ( .A1(n9353), .A2(n5591), .ZN(n5915) );
  NAND2_X1 U6948 ( .A1(n6418), .A2(P2_REG1_REG_17__SCAN_IN), .ZN(n5914) );
  OR2_X1 U6949 ( .A1(n9338), .A2(n5747), .ZN(n5918) );
  AND2_X1 U6950 ( .A1(n5917), .A2(n5918), .ZN(n7994) );
  INV_X1 U6951 ( .A(n5917), .ZN(n5920) );
  INV_X1 U6952 ( .A(n5918), .ZN(n5919) );
  NAND2_X1 U6953 ( .A1(n5920), .A2(n5919), .ZN(n7995) );
  NAND2_X1 U6954 ( .A1(n5922), .A2(n5921), .ZN(n5927) );
  MUX2_X1 U6955 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(P2_DATAO_REG_18__SCAN_IN), 
        .S(n8387), .Z(n5923) );
  NAND2_X1 U6956 ( .A1(n5923), .A2(SI_18_), .ZN(n5943) );
  INV_X1 U6957 ( .A(n5923), .ZN(n5924) );
  INV_X1 U6958 ( .A(SI_18_), .ZN(n10184) );
  NAND2_X1 U6959 ( .A1(n5924), .A2(n10184), .ZN(n5925) );
  OR2_X1 U6960 ( .A1(n5927), .A2(n5926), .ZN(n5928) );
  NAND2_X1 U6961 ( .A1(n5944), .A2(n5928), .ZN(n8142) );
  NAND2_X1 U6962 ( .A1(n5929), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n5930) );
  XNOR2_X1 U6963 ( .A(n5930), .B(P2_IR_REG_18__SCAN_IN), .ZN(n9090) );
  AOI22_X1 U6964 ( .A1(n5945), .A2(P1_DATAO_REG_18__SCAN_IN), .B1(n6433), .B2(
        n9090), .ZN(n5931) );
  XNOR2_X1 U6965 ( .A(n9451), .B(n6115), .ZN(n5938) );
  INV_X1 U6966 ( .A(P2_REG0_REG_18__SCAN_IN), .ZN(n5937) );
  INV_X1 U6967 ( .A(P2_REG3_REG_18__SCAN_IN), .ZN(n10267) );
  INV_X1 U6968 ( .A(n5948), .ZN(n5950) );
  NAND2_X1 U6969 ( .A1(n5933), .A2(n10267), .ZN(n5934) );
  NAND2_X1 U6970 ( .A1(n5950), .A2(n5934), .ZN(n9330) );
  OR2_X1 U6971 ( .A1(n9330), .A2(n5682), .ZN(n5936) );
  AOI22_X1 U6972 ( .A1(n5589), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n6418), .B2(
        P2_REG1_REG_18__SCAN_IN), .ZN(n5935) );
  OAI211_X1 U6973 ( .C1(n5548), .C2(n5937), .A(n5936), .B(n5935), .ZN(n9057)
         );
  NAND2_X1 U6974 ( .A1(n9057), .A2(n5621), .ZN(n5939) );
  NAND2_X1 U6975 ( .A1(n5938), .A2(n5939), .ZN(n8097) );
  INV_X1 U6976 ( .A(n5938), .ZN(n5941) );
  INV_X1 U6977 ( .A(n5939), .ZN(n5940) );
  NAND2_X1 U6978 ( .A1(n5941), .A2(n5940), .ZN(n8098) );
  NAND2_X1 U6979 ( .A1(n5942), .A2(n8098), .ZN(n8960) );
  INV_X1 U6980 ( .A(n8960), .ZN(n5956) );
  MUX2_X1 U6981 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(P2_DATAO_REG_19__SCAN_IN), 
        .S(n8387), .Z(n5961) );
  XNOR2_X1 U6982 ( .A(n5961), .B(SI_19_), .ZN(n5963) );
  XNOR2_X1 U6983 ( .A(n5964), .B(n5963), .ZN(n8152) );
  NAND2_X1 U6984 ( .A1(n8152), .A2(n8726), .ZN(n5947) );
  AOI22_X1 U6985 ( .A1(n5945), .A2(P1_DATAO_REG_19__SCAN_IN), .B1(n9317), .B2(
        n6433), .ZN(n5946) );
  XNOR2_X1 U6986 ( .A(n9448), .B(n5615), .ZN(n8957) );
  INV_X1 U6987 ( .A(n5968), .ZN(n5969) );
  INV_X1 U6988 ( .A(P2_REG3_REG_19__SCAN_IN), .ZN(n5949) );
  NAND2_X1 U6989 ( .A1(n5950), .A2(n5949), .ZN(n5951) );
  AND2_X1 U6990 ( .A1(n5969), .A2(n5951), .ZN(n9314) );
  NAND2_X1 U6991 ( .A1(n9314), .A2(n5591), .ZN(n5954) );
  AOI22_X1 U6992 ( .A1(n6419), .A2(P2_REG0_REG_19__SCAN_IN), .B1(n5589), .B2(
        P2_REG2_REG_19__SCAN_IN), .ZN(n5953) );
  NAND2_X1 U6993 ( .A1(n6418), .A2(P2_REG1_REG_19__SCAN_IN), .ZN(n5952) );
  NOR2_X1 U6994 ( .A1(n9339), .A2(n5542), .ZN(n5957) );
  AND2_X1 U6995 ( .A1(n8957), .A2(n5957), .ZN(n8954) );
  INV_X1 U6996 ( .A(n8954), .ZN(n5955) );
  INV_X1 U6997 ( .A(n8957), .ZN(n5959) );
  INV_X1 U6998 ( .A(n5957), .ZN(n5958) );
  NAND2_X1 U6999 ( .A1(n5959), .A2(n5958), .ZN(n8959) );
  INV_X1 U7000 ( .A(n5961), .ZN(n5962) );
  INV_X1 U7001 ( .A(SI_19_), .ZN(n10061) );
  MUX2_X1 U7002 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(P2_DATAO_REG_20__SCAN_IN), 
        .S(n8387), .Z(n5981) );
  INV_X1 U7003 ( .A(SI_20_), .ZN(n10062) );
  XNOR2_X1 U7004 ( .A(n5983), .B(n5982), .ZN(n8167) );
  NAND2_X1 U7005 ( .A1(n8167), .A2(n8726), .ZN(n5967) );
  INV_X1 U7006 ( .A(P1_DATAO_REG_20__SCAN_IN), .ZN(n7612) );
  OR2_X1 U7007 ( .A1(n5965), .A2(n7612), .ZN(n5966) );
  XNOR2_X1 U7008 ( .A(n9441), .B(n5615), .ZN(n5977) );
  INV_X1 U7009 ( .A(P2_REG3_REG_20__SCAN_IN), .ZN(n10057) );
  NAND2_X1 U7010 ( .A1(n5969), .A2(n10057), .ZN(n5970) );
  NAND2_X1 U7011 ( .A1(n5994), .A2(n5970), .ZN(n9301) );
  OR2_X1 U7012 ( .A1(n9301), .A2(n5682), .ZN(n5976) );
  INV_X1 U7013 ( .A(P2_REG0_REG_20__SCAN_IN), .ZN(n5973) );
  NAND2_X1 U7014 ( .A1(n6418), .A2(P2_REG1_REG_20__SCAN_IN), .ZN(n5972) );
  NAND2_X1 U7015 ( .A1(n5589), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n5971) );
  OAI211_X1 U7016 ( .C1(n5548), .C2(n5973), .A(n5972), .B(n5971), .ZN(n5974)
         );
  INV_X1 U7017 ( .A(n5974), .ZN(n5975) );
  NOR2_X1 U7018 ( .A1(n9274), .A2(n5542), .ZN(n5978) );
  XNOR2_X1 U7019 ( .A(n5977), .B(n5978), .ZN(n9025) );
  INV_X1 U7020 ( .A(n5977), .ZN(n5980) );
  INV_X1 U7021 ( .A(n5978), .ZN(n5979) );
  MUX2_X1 U7022 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(P2_DATAO_REG_21__SCAN_IN), 
        .S(n8387), .Z(n5984) );
  NAND2_X1 U7023 ( .A1(n5984), .A2(SI_21_), .ZN(n6006) );
  INV_X1 U7024 ( .A(n5984), .ZN(n5985) );
  INV_X1 U7025 ( .A(SI_21_), .ZN(n10182) );
  NAND2_X1 U7026 ( .A1(n5985), .A2(n10182), .ZN(n5986) );
  NAND2_X1 U7027 ( .A1(n6006), .A2(n5986), .ZN(n5989) );
  INV_X1 U7028 ( .A(n5989), .ZN(n5987) );
  NAND2_X1 U7029 ( .A1(n5988), .A2(n5987), .ZN(n6007) );
  NAND2_X1 U7030 ( .A1(n5268), .A2(n5989), .ZN(n5990) );
  NAND2_X1 U7031 ( .A1(n6007), .A2(n5990), .ZN(n8179) );
  INV_X1 U7032 ( .A(P1_DATAO_REG_21__SCAN_IN), .ZN(n7577) );
  OR2_X1 U7033 ( .A1(n5965), .A2(n7577), .ZN(n5991) );
  XNOR2_X1 U7034 ( .A(n9436), .B(n6115), .ZN(n6002) );
  INV_X1 U7035 ( .A(P2_REG3_REG_21__SCAN_IN), .ZN(n5993) );
  NAND2_X1 U7036 ( .A1(n5994), .A2(n5993), .ZN(n5995) );
  AND2_X1 U7037 ( .A1(n6010), .A2(n5995), .ZN(n9284) );
  NAND2_X1 U7038 ( .A1(n9284), .A2(n5591), .ZN(n6001) );
  INV_X1 U7039 ( .A(P2_REG0_REG_21__SCAN_IN), .ZN(n5998) );
  NAND2_X1 U7040 ( .A1(n6418), .A2(P2_REG1_REG_21__SCAN_IN), .ZN(n5997) );
  NAND2_X1 U7041 ( .A1(n5589), .A2(P2_REG2_REG_21__SCAN_IN), .ZN(n5996) );
  OAI211_X1 U7042 ( .C1(n5548), .C2(n5998), .A(n5997), .B(n5996), .ZN(n5999)
         );
  INV_X1 U7043 ( .A(n5999), .ZN(n6000) );
  NOR2_X1 U7044 ( .A1(n9293), .A2(n5747), .ZN(n6003) );
  XNOR2_X1 U7045 ( .A(n6002), .B(n6003), .ZN(n8980) );
  INV_X1 U7046 ( .A(n6002), .ZN(n6004) );
  NAND2_X1 U7047 ( .A1(n6004), .A2(n6003), .ZN(n6005) );
  MUX2_X1 U7048 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(P2_DATAO_REG_22__SCAN_IN), 
        .S(n8387), .Z(n6024) );
  XNOR2_X1 U7049 ( .A(n6024), .B(SI_22_), .ZN(n6027) );
  XNOR2_X1 U7050 ( .A(n6028), .B(n6027), .ZN(n8193) );
  NAND2_X1 U7051 ( .A1(n8193), .A2(n8726), .ZN(n6009) );
  INV_X1 U7052 ( .A(P1_DATAO_REG_22__SCAN_IN), .ZN(n8316) );
  OR2_X1 U7053 ( .A1(n5965), .A2(n8316), .ZN(n6008) );
  XNOR2_X1 U7054 ( .A(n9430), .B(n6115), .ZN(n6018) );
  INV_X1 U7055 ( .A(P2_REG3_REG_22__SCAN_IN), .ZN(n10264) );
  INV_X1 U7056 ( .A(n6031), .ZN(n6032) );
  NAND2_X1 U7057 ( .A1(n6010), .A2(n10264), .ZN(n6011) );
  NAND2_X1 U7058 ( .A1(n6032), .A2(n6011), .ZN(n9035) );
  OR2_X1 U7059 ( .A1(n9035), .A2(n5682), .ZN(n6017) );
  INV_X1 U7060 ( .A(P2_REG0_REG_22__SCAN_IN), .ZN(n6014) );
  NAND2_X1 U7061 ( .A1(n5589), .A2(P2_REG2_REG_22__SCAN_IN), .ZN(n6013) );
  NAND2_X1 U7062 ( .A1(n6418), .A2(P2_REG1_REG_22__SCAN_IN), .ZN(n6012) );
  OAI211_X1 U7063 ( .C1(n5548), .C2(n6014), .A(n6013), .B(n6012), .ZN(n6015)
         );
  INV_X1 U7064 ( .A(n6015), .ZN(n6016) );
  INV_X1 U7065 ( .A(n9275), .ZN(n9240) );
  NAND2_X1 U7066 ( .A1(n9240), .A2(n5621), .ZN(n6019) );
  NAND2_X1 U7067 ( .A1(n6018), .A2(n6019), .ZN(n6023) );
  INV_X1 U7068 ( .A(n6018), .ZN(n6021) );
  INV_X1 U7069 ( .A(n6019), .ZN(n6020) );
  NAND2_X1 U7070 ( .A1(n6021), .A2(n6020), .ZN(n6022) );
  NAND2_X1 U7071 ( .A1(n6023), .A2(n6022), .ZN(n9031) );
  INV_X1 U7072 ( .A(n6024), .ZN(n6025) );
  INV_X1 U7073 ( .A(SI_22_), .ZN(n10157) );
  NAND2_X1 U7074 ( .A1(n6025), .A2(n10157), .ZN(n6026) );
  MUX2_X1 U7075 ( .A(P1_DATAO_REG_23__SCAN_IN), .B(P2_DATAO_REG_23__SCAN_IN), 
        .S(n8387), .Z(n6043) );
  INV_X1 U7076 ( .A(SI_23_), .ZN(n10158) );
  XNOR2_X1 U7077 ( .A(n6043), .B(n10158), .ZN(n6044) );
  NAND2_X1 U7078 ( .A1(n8208), .A2(n8726), .ZN(n6030) );
  INV_X1 U7079 ( .A(P1_DATAO_REG_23__SCAN_IN), .ZN(n7788) );
  OR2_X1 U7080 ( .A1(n5965), .A2(n7788), .ZN(n6029) );
  XNOR2_X1 U7081 ( .A(n8709), .B(n5615), .ZN(n6038) );
  INV_X1 U7082 ( .A(n6056), .ZN(n6057) );
  INV_X1 U7083 ( .A(P2_REG3_REG_23__SCAN_IN), .ZN(n10115) );
  NAND2_X1 U7084 ( .A1(n6032), .A2(n10115), .ZN(n6033) );
  INV_X1 U7085 ( .A(P2_REG0_REG_23__SCAN_IN), .ZN(n6036) );
  NAND2_X1 U7086 ( .A1(n5589), .A2(P2_REG2_REG_23__SCAN_IN), .ZN(n6035) );
  NAND2_X1 U7087 ( .A1(n6418), .A2(P2_REG1_REG_23__SCAN_IN), .ZN(n6034) );
  OAI211_X1 U7088 ( .C1(n6036), .C2(n5548), .A(n6035), .B(n6034), .ZN(n6037)
         );
  AOI21_X1 U7089 ( .B1(n9248), .B2(n5591), .A(n6037), .ZN(n9264) );
  NOR2_X1 U7090 ( .A1(n9264), .A2(n5542), .ZN(n8944) );
  NAND2_X1 U7091 ( .A1(n8945), .A2(n8944), .ZN(n6042) );
  INV_X1 U7092 ( .A(n6038), .ZN(n6039) );
  OR2_X1 U7093 ( .A1(n6040), .A2(n6039), .ZN(n6041) );
  NAND2_X1 U7094 ( .A1(n6042), .A2(n6041), .ZN(n6067) );
  MUX2_X1 U7095 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(P2_DATAO_REG_24__SCAN_IN), 
        .S(n8387), .Z(n6046) );
  NAND2_X1 U7096 ( .A1(n6046), .A2(SI_24_), .ZN(n6069) );
  INV_X1 U7097 ( .A(n6046), .ZN(n6047) );
  INV_X1 U7098 ( .A(SI_24_), .ZN(n10179) );
  NAND2_X1 U7099 ( .A1(n6047), .A2(n10179), .ZN(n6048) );
  NAND2_X1 U7100 ( .A1(n6069), .A2(n6048), .ZN(n6051) );
  INV_X1 U7101 ( .A(n6051), .ZN(n6049) );
  NAND2_X1 U7102 ( .A1(n6050), .A2(n6049), .ZN(n6070) );
  NAND2_X1 U7103 ( .A1(n6052), .A2(n6051), .ZN(n6053) );
  NAND2_X1 U7104 ( .A1(n6070), .A2(n6053), .ZN(n8212) );
  INV_X1 U7105 ( .A(P1_DATAO_REG_24__SCAN_IN), .ZN(n7831) );
  OR2_X1 U7106 ( .A1(n5965), .A2(n7831), .ZN(n6054) );
  XNOR2_X1 U7107 ( .A(n9420), .B(n6115), .ZN(n6065) );
  INV_X1 U7108 ( .A(P2_REG3_REG_24__SCAN_IN), .ZN(n10059) );
  NAND2_X1 U7109 ( .A1(n6057), .A2(n10059), .ZN(n6058) );
  NAND2_X1 U7110 ( .A1(n6073), .A2(n6058), .ZN(n9003) );
  OR2_X1 U7111 ( .A1(n9003), .A2(n5682), .ZN(n6064) );
  INV_X1 U7112 ( .A(P2_REG0_REG_24__SCAN_IN), .ZN(n6061) );
  NAND2_X1 U7113 ( .A1(n6418), .A2(P2_REG1_REG_24__SCAN_IN), .ZN(n6060) );
  NAND2_X1 U7114 ( .A1(n5589), .A2(P2_REG2_REG_24__SCAN_IN), .ZN(n6059) );
  OAI211_X1 U7115 ( .C1(n5548), .C2(n6061), .A(n6060), .B(n6059), .ZN(n6062)
         );
  INV_X1 U7116 ( .A(n6062), .ZN(n6063) );
  NOR2_X1 U7117 ( .A1(n9138), .A2(n5747), .ZN(n8999) );
  INV_X1 U7118 ( .A(n6065), .ZN(n6066) );
  NAND2_X1 U7119 ( .A1(n6067), .A2(n6066), .ZN(n6068) );
  NAND2_X1 U7120 ( .A1(n6070), .A2(n6069), .ZN(n6091) );
  MUX2_X1 U7121 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(P2_DATAO_REG_25__SCAN_IN), 
        .S(n8387), .Z(n6087) );
  XNOR2_X1 U7122 ( .A(n6087), .B(SI_25_), .ZN(n6090) );
  XNOR2_X1 U7123 ( .A(n6091), .B(n6090), .ZN(n8226) );
  NAND2_X1 U7124 ( .A1(n8226), .A2(n8726), .ZN(n6072) );
  INV_X1 U7125 ( .A(P1_DATAO_REG_25__SCAN_IN), .ZN(n7965) );
  OR2_X1 U7126 ( .A1(n5965), .A2(n7965), .ZN(n6071) );
  XNOR2_X1 U7127 ( .A(n9417), .B(n6115), .ZN(n6081) );
  INV_X1 U7128 ( .A(P2_REG3_REG_25__SCAN_IN), .ZN(n8993) );
  NAND2_X1 U7129 ( .A1(n6073), .A2(n8993), .ZN(n6074) );
  NAND2_X1 U7130 ( .A1(n6094), .A2(n6074), .ZN(n9213) );
  OR2_X1 U7131 ( .A1(n9213), .A2(n5682), .ZN(n6080) );
  INV_X1 U7132 ( .A(P2_REG0_REG_25__SCAN_IN), .ZN(n6077) );
  NAND2_X1 U7133 ( .A1(n6418), .A2(P2_REG1_REG_25__SCAN_IN), .ZN(n6076) );
  NAND2_X1 U7134 ( .A1(n5589), .A2(P2_REG2_REG_25__SCAN_IN), .ZN(n6075) );
  OAI211_X1 U7135 ( .C1(n5548), .C2(n6077), .A(n6076), .B(n6075), .ZN(n6078)
         );
  INV_X1 U7136 ( .A(n6078), .ZN(n6079) );
  INV_X1 U7137 ( .A(n9233), .ZN(n9054) );
  NAND2_X1 U7138 ( .A1(n9054), .A2(n5621), .ZN(n6082) );
  NAND2_X1 U7139 ( .A1(n6081), .A2(n6082), .ZN(n6086) );
  INV_X1 U7140 ( .A(n6081), .ZN(n6084) );
  INV_X1 U7141 ( .A(n6082), .ZN(n6083) );
  NAND2_X1 U7142 ( .A1(n6084), .A2(n6083), .ZN(n6085) );
  NAND2_X1 U7143 ( .A1(n6086), .A2(n6085), .ZN(n8989) );
  NAND2_X1 U7144 ( .A1(n8987), .A2(n6086), .ZN(n9040) );
  INV_X1 U7145 ( .A(n9040), .ZN(n6103) );
  INV_X1 U7146 ( .A(n6087), .ZN(n6088) );
  INV_X1 U7147 ( .A(SI_25_), .ZN(n10174) );
  NAND2_X1 U7148 ( .A1(n6088), .A2(n10174), .ZN(n6089) );
  MUX2_X1 U7149 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(P2_DATAO_REG_26__SCAN_IN), 
        .S(n8387), .Z(n6109) );
  INV_X1 U7150 ( .A(SI_26_), .ZN(n10171) );
  XNOR2_X1 U7151 ( .A(n6109), .B(n10171), .ZN(n6107) );
  NAND2_X1 U7152 ( .A1(n8243), .A2(n8726), .ZN(n6093) );
  INV_X1 U7153 ( .A(P1_DATAO_REG_26__SCAN_IN), .ZN(n8080) );
  OR2_X1 U7154 ( .A1(n5965), .A2(n8080), .ZN(n6092) );
  XNOR2_X1 U7155 ( .A(n9411), .B(n5615), .ZN(n6105) );
  INV_X1 U7156 ( .A(P2_REG3_REG_26__SCAN_IN), .ZN(n10272) );
  NAND2_X1 U7157 ( .A1(n6094), .A2(n10272), .ZN(n6095) );
  NAND2_X1 U7158 ( .A1(n9194), .A2(n5591), .ZN(n6101) );
  INV_X1 U7159 ( .A(P2_REG0_REG_26__SCAN_IN), .ZN(n6098) );
  NAND2_X1 U7160 ( .A1(n6418), .A2(P2_REG1_REG_26__SCAN_IN), .ZN(n6097) );
  NAND2_X1 U7161 ( .A1(n5589), .A2(P2_REG2_REG_26__SCAN_IN), .ZN(n6096) );
  OAI211_X1 U7162 ( .C1(n5548), .C2(n6098), .A(n6097), .B(n6096), .ZN(n6099)
         );
  INV_X1 U7163 ( .A(n6099), .ZN(n6100) );
  NOR2_X1 U7164 ( .A1(n8991), .A2(n5747), .ZN(n6104) );
  XNOR2_X1 U7165 ( .A(n6105), .B(n6104), .ZN(n9041) );
  INV_X1 U7166 ( .A(n9041), .ZN(n6102) );
  NAND2_X1 U7167 ( .A1(n6105), .A2(n6104), .ZN(n6106) );
  NAND2_X1 U7168 ( .A1(n6108), .A2(n6107), .ZN(n6112) );
  INV_X1 U7169 ( .A(n6109), .ZN(n6110) );
  NAND2_X1 U7170 ( .A1(n6110), .A2(n10171), .ZN(n6111) );
  MUX2_X1 U7171 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(P2_DATAO_REG_27__SCAN_IN), 
        .S(n8387), .Z(n6137) );
  INV_X1 U7172 ( .A(SI_27_), .ZN(n10169) );
  XNOR2_X1 U7173 ( .A(n6137), .B(n10169), .ZN(n6135) );
  NAND2_X1 U7174 ( .A1(n8259), .A2(n8726), .ZN(n6114) );
  INV_X1 U7175 ( .A(P1_DATAO_REG_27__SCAN_IN), .ZN(n8105) );
  OR2_X1 U7176 ( .A1(n5965), .A2(n8105), .ZN(n6113) );
  XNOR2_X1 U7177 ( .A(n9405), .B(n6115), .ZN(n6120) );
  XNOR2_X1 U7178 ( .A(n6126), .B(P2_REG3_REG_27__SCAN_IN), .ZN(n9180) );
  INV_X1 U7179 ( .A(P2_REG0_REG_27__SCAN_IN), .ZN(n6118) );
  NAND2_X1 U7180 ( .A1(n6418), .A2(P2_REG1_REG_27__SCAN_IN), .ZN(n6117) );
  NAND2_X1 U7181 ( .A1(n5589), .A2(P2_REG2_REG_27__SCAN_IN), .ZN(n6116) );
  OAI211_X1 U7182 ( .C1(n5548), .C2(n6118), .A(n6117), .B(n6116), .ZN(n6119)
         );
  NOR2_X1 U7183 ( .A1(n9053), .A2(n5542), .ZN(n6121) );
  XNOR2_X1 U7184 ( .A(n6120), .B(n6121), .ZN(n8936) );
  INV_X1 U7185 ( .A(n6120), .ZN(n6122) );
  INV_X1 U7186 ( .A(n6126), .ZN(n6124) );
  AND2_X1 U7187 ( .A1(P2_REG3_REG_27__SCAN_IN), .A2(P2_REG3_REG_28__SCAN_IN), 
        .ZN(n6123) );
  NAND2_X1 U7188 ( .A1(n6124), .A2(n6123), .ZN(n6189) );
  INV_X1 U7189 ( .A(P2_REG3_REG_27__SCAN_IN), .ZN(n10112) );
  INV_X1 U7190 ( .A(P2_REG3_REG_28__SCAN_IN), .ZN(n6125) );
  OAI21_X1 U7191 ( .B1(n6126), .B2(n10112), .A(n6125), .ZN(n6127) );
  NAND2_X1 U7192 ( .A1(n6189), .A2(n6127), .ZN(n6198) );
  OR2_X1 U7193 ( .A1(n6198), .A2(n5682), .ZN(n6133) );
  INV_X1 U7194 ( .A(P2_REG0_REG_28__SCAN_IN), .ZN(n6130) );
  NAND2_X1 U7195 ( .A1(n6418), .A2(P2_REG1_REG_28__SCAN_IN), .ZN(n6129) );
  NAND2_X1 U7196 ( .A1(n5589), .A2(P2_REG2_REG_28__SCAN_IN), .ZN(n6128) );
  OAI211_X1 U7197 ( .C1(n5548), .C2(n6130), .A(n6129), .B(n6128), .ZN(n6131)
         );
  INV_X1 U7198 ( .A(n6131), .ZN(n6132) );
  NOR2_X1 U7199 ( .A1(n9146), .A2(n5542), .ZN(n6134) );
  MUX2_X1 U7200 ( .A(n6134), .B(n9146), .S(n5615), .Z(n6180) );
  INV_X1 U7201 ( .A(n6137), .ZN(n6138) );
  NAND2_X1 U7202 ( .A1(n6138), .A2(n10169), .ZN(n6139) );
  MUX2_X1 U7203 ( .A(P1_DATAO_REG_28__SCAN_IN), .B(P2_DATAO_REG_28__SCAN_IN), 
        .S(n8387), .Z(n8321) );
  INV_X1 U7204 ( .A(SI_28_), .ZN(n10165) );
  XNOR2_X1 U7205 ( .A(n8321), .B(n10165), .ZN(n8319) );
  NAND2_X1 U7206 ( .A1(n8604), .A2(n8726), .ZN(n6142) );
  INV_X1 U7207 ( .A(P1_DATAO_REG_28__SCAN_IN), .ZN(n8605) );
  OR2_X1 U7208 ( .A1(n5965), .A2(n8605), .ZN(n6141) );
  INV_X1 U7209 ( .A(n9400), .ZN(n9168) );
  NOR4_X1 U7210 ( .A1(P2_D_REG_27__SCAN_IN), .A2(P2_D_REG_26__SCAN_IN), .A3(
        P2_D_REG_25__SCAN_IN), .A4(P2_D_REG_24__SCAN_IN), .ZN(n6151) );
  NOR4_X1 U7211 ( .A1(P2_D_REG_23__SCAN_IN), .A2(P2_D_REG_22__SCAN_IN), .A3(
        P2_D_REG_21__SCAN_IN), .A4(P2_D_REG_20__SCAN_IN), .ZN(n6150) );
  OR4_X1 U7212 ( .A1(P2_D_REG_31__SCAN_IN), .A2(P2_D_REG_30__SCAN_IN), .A3(
        P2_D_REG_29__SCAN_IN), .A4(P2_D_REG_28__SCAN_IN), .ZN(n6148) );
  NOR4_X1 U7213 ( .A1(P2_D_REG_15__SCAN_IN), .A2(P2_D_REG_14__SCAN_IN), .A3(
        P2_D_REG_13__SCAN_IN), .A4(P2_D_REG_12__SCAN_IN), .ZN(n6146) );
  NOR4_X1 U7214 ( .A1(P2_D_REG_17__SCAN_IN), .A2(P2_D_REG_19__SCAN_IN), .A3(
        P2_D_REG_18__SCAN_IN), .A4(P2_D_REG_16__SCAN_IN), .ZN(n6145) );
  NOR4_X1 U7215 ( .A1(P2_D_REG_7__SCAN_IN), .A2(P2_D_REG_6__SCAN_IN), .A3(
        P2_D_REG_5__SCAN_IN), .A4(P2_D_REG_2__SCAN_IN), .ZN(n6144) );
  NOR4_X1 U7216 ( .A1(P2_D_REG_11__SCAN_IN), .A2(P2_D_REG_10__SCAN_IN), .A3(
        P2_D_REG_9__SCAN_IN), .A4(P2_D_REG_8__SCAN_IN), .ZN(n6143) );
  NAND4_X1 U7217 ( .A1(n6146), .A2(n6145), .A3(n6144), .A4(n6143), .ZN(n6147)
         );
  NOR4_X1 U7218 ( .A1(P2_D_REG_4__SCAN_IN), .A2(P2_D_REG_3__SCAN_IN), .A3(
        n6148), .A4(n6147), .ZN(n6149) );
  AND3_X1 U7219 ( .A1(n6151), .A2(n6150), .A3(n6149), .ZN(n6165) );
  INV_X1 U7220 ( .A(n6152), .ZN(n6153) );
  NAND2_X1 U7221 ( .A1(n6153), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6154) );
  NAND2_X1 U7222 ( .A1(n6155), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6156) );
  XNOR2_X1 U7223 ( .A(n6156), .B(P2_IR_REG_25__SCAN_IN), .ZN(n10049) );
  NAND2_X1 U7224 ( .A1(n6158), .A2(n6157), .ZN(n6159) );
  NAND2_X1 U7225 ( .A1(n6173), .A2(n6172), .ZN(n6160) );
  NAND2_X1 U7226 ( .A1(n6160), .A2(P2_IR_REG_31__SCAN_IN), .ZN(n6161) );
  INV_X1 U7227 ( .A(n10409), .ZN(n7832) );
  INV_X1 U7228 ( .A(P2_B_REG_SCAN_IN), .ZN(n6162) );
  AOI22_X1 U7229 ( .A1(P2_B_REG_SCAN_IN), .A2(n7832), .B1(n10409), .B2(n6162), 
        .ZN(n6163) );
  OR2_X1 U7230 ( .A1(n10409), .A2(n10408), .ZN(n6167) );
  OR2_X1 U7231 ( .A1(n10051), .A2(P2_D_REG_0__SCAN_IN), .ZN(n6166) );
  OR2_X1 U7232 ( .A1(n10051), .A2(P2_D_REG_1__SCAN_IN), .ZN(n6169) );
  OR2_X1 U7233 ( .A1(n10408), .A2(n10049), .ZN(n6168) );
  NAND2_X1 U7234 ( .A1(n6169), .A2(n6168), .ZN(n6947) );
  OR2_X1 U7235 ( .A1(n6956), .A2(n6947), .ZN(n6170) );
  AND2_X1 U7236 ( .A1(n10408), .A2(n10049), .ZN(n6171) );
  XNOR2_X1 U7237 ( .A(n6173), .B(n6172), .ZN(n6432) );
  INV_X1 U7238 ( .A(n10413), .ZN(n6174) );
  NOR2_X1 U7239 ( .A1(n6201), .A2(n10050), .ZN(n6184) );
  AND2_X1 U7240 ( .A1(n5523), .A2(n8896), .ZN(n6282) );
  NAND2_X1 U7241 ( .A1(n6184), .A2(n6282), .ZN(n6176) );
  NAND3_X1 U7242 ( .A1(n8926), .A2(n6175), .A3(n9317), .ZN(n6971) );
  NOR3_X1 U7243 ( .A1(n9168), .A2(n6180), .A3(n10293), .ZN(n6177) );
  AOI21_X1 U7244 ( .B1(n6180), .B2(n9168), .A(n6177), .ZN(n6178) );
  NAND3_X1 U7245 ( .A1(n9400), .A2(n6180), .A3(n9046), .ZN(n6179) );
  OAI21_X1 U7246 ( .B1(n9400), .B2(n6180), .A(n6179), .ZN(n6181) );
  NAND2_X1 U7247 ( .A1(n6182), .A2(n6181), .ZN(n6186) );
  NAND2_X1 U7248 ( .A1(n8926), .A2(n5298), .ZN(n8932) );
  NAND2_X1 U7249 ( .A1(n8933), .A2(n8733), .ZN(n6435) );
  INV_X1 U7250 ( .A(n6435), .ZN(n6642) );
  NOR2_X1 U7251 ( .A1(n9458), .A2(n6642), .ZN(n6183) );
  OAI21_X1 U7252 ( .B1(n9168), .B2(n9046), .A(n10288), .ZN(n6185) );
  NAND3_X1 U7253 ( .A1(n6187), .A2(n6186), .A3(n6185), .ZN(n6211) );
  OR2_X1 U7254 ( .A1(n9053), .A2(n9371), .ZN(n6195) );
  INV_X1 U7255 ( .A(n6189), .ZN(n9153) );
  INV_X1 U7256 ( .A(P2_REG0_REG_29__SCAN_IN), .ZN(n6192) );
  NAND2_X1 U7257 ( .A1(n6418), .A2(P2_REG1_REG_29__SCAN_IN), .ZN(n6191) );
  NAND2_X1 U7258 ( .A1(n5589), .A2(P2_REG2_REG_29__SCAN_IN), .ZN(n6190) );
  OAI211_X1 U7259 ( .C1(n5548), .C2(n6192), .A(n6191), .B(n6190), .ZN(n6193)
         );
  AOI21_X1 U7260 ( .B1(n9153), .B2(n5591), .A(n6193), .ZN(n8715) );
  INV_X1 U7261 ( .A(n6188), .ZN(n6673) );
  OR2_X1 U7262 ( .A1(n8715), .A2(n9370), .ZN(n6194) );
  NAND2_X1 U7263 ( .A1(n6195), .A2(n6194), .ZN(n9172) );
  INV_X1 U7264 ( .A(n9172), .ZN(n6208) );
  INV_X1 U7265 ( .A(n6201), .ZN(n6197) );
  NOR2_X1 U7266 ( .A1(n10050), .A2(n8932), .ZN(n6196) );
  NAND2_X1 U7267 ( .A1(n6197), .A2(n6196), .ZN(n8994) );
  INV_X1 U7268 ( .A(n6198), .ZN(n9166) );
  INV_X1 U7269 ( .A(n6282), .ZN(n6199) );
  OAI22_X1 U7270 ( .A1(n10050), .A2(n6199), .B1(n9458), .B2(P2_U3152), .ZN(
        n6200) );
  NAND2_X1 U7271 ( .A1(n6201), .A2(n6200), .ZN(n6206) );
  INV_X1 U7272 ( .A(n6432), .ZN(n6204) );
  INV_X1 U7273 ( .A(n8932), .ZN(n6202) );
  NOR2_X1 U7274 ( .A1(n6202), .A2(n6435), .ZN(n6203) );
  NAND2_X1 U7275 ( .A1(n6265), .A2(P2_STATE_REG_SCAN_IN), .ZN(n6205) );
  AOI22_X1 U7276 ( .A1(n9166), .A2(n10284), .B1(P2_REG3_REG_28__SCAN_IN), .B2(
        P2_U3152), .ZN(n6207) );
  OAI21_X1 U7277 ( .B1(n6208), .B2(n8994), .A(n6207), .ZN(n6209) );
  NAND2_X1 U7278 ( .A1(n6211), .A2(n6210), .ZN(P2_U3222) );
  NAND4_X1 U7279 ( .A1(n6214), .A2(n6213), .A3(n6212), .A4(n6294), .ZN(n6218)
         );
  NAND4_X1 U7280 ( .A1(n6357), .A2(n6354), .A3(n6216), .A4(n6215), .ZN(n6217)
         );
  NOR2_X1 U7281 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_7__SCAN_IN), .ZN(
        n6223) );
  NOR2_X1 U7282 ( .A1(P1_IR_REG_21__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n6222) );
  NOR2_X1 U7283 ( .A1(P1_IR_REG_20__SCAN_IN), .A2(P1_IR_REG_19__SCAN_IN), .ZN(
        n6221) );
  NOR2_X1 U7284 ( .A1(P1_IR_REG_6__SCAN_IN), .A2(P1_IR_REG_22__SCAN_IN), .ZN(
        n6220) );
  NAND2_X1 U7285 ( .A1(n6249), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6229) );
  INV_X1 U7286 ( .A(P1_IR_REG_25__SCAN_IN), .ZN(n6228) );
  NAND2_X1 U7287 ( .A1(n6229), .A2(n6228), .ZN(n6231) );
  INV_X1 U7288 ( .A(P1_IR_REG_26__SCAN_IN), .ZN(n6224) );
  NAND2_X1 U7289 ( .A1(n4913), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6227) );
  XNOR2_X1 U7290 ( .A(n6227), .B(n6226), .ZN(n7808) );
  OR2_X1 U7291 ( .A1(n6229), .A2(n6228), .ZN(n6230) );
  NAND2_X1 U7292 ( .A1(n6231), .A2(n6230), .ZN(n7964) );
  NAND2_X1 U7293 ( .A1(n6232), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6233) );
  XNOR2_X1 U7294 ( .A(n6233), .B(n5374), .ZN(n6762) );
  INV_X1 U7295 ( .A(n6393), .ZN(n6234) );
  NOR2_X2 U7296 ( .A1(n6581), .A2(n6234), .ZN(P1_U4006) );
  NOR2_X1 U7297 ( .A1(P1_IR_REG_8__SCAN_IN), .A2(P1_IR_REG_9__SCAN_IN), .ZN(
        n6236) );
  INV_X1 U7298 ( .A(n6237), .ZN(n6238) );
  NOR2_X2 U7299 ( .A1(n6288), .A2(n6238), .ZN(n6478) );
  NAND2_X1 U7300 ( .A1(n6478), .A2(n6239), .ZN(n6240) );
  INV_X1 U7301 ( .A(P1_IR_REG_20__SCAN_IN), .ZN(n6241) );
  NAND2_X1 U7302 ( .A1(n6477), .A2(n6241), .ZN(n6242) );
  NAND2_X1 U7303 ( .A1(n6247), .A2(n6246), .ZN(n6243) );
  INV_X1 U7304 ( .A(P1_IR_REG_22__SCAN_IN), .ZN(n6244) );
  XNOR2_X1 U7305 ( .A(n6245), .B(n6244), .ZN(n6607) );
  NAND2_X1 U7306 ( .A1(n8553), .A2(n6581), .ZN(n6248) );
  NAND2_X1 U7307 ( .A1(n6248), .A2(n6762), .ZN(n6361) );
  NAND2_X1 U7308 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_27__SCAN_IN), 
        .ZN(n6251) );
  NAND2_X1 U7309 ( .A1(n6253), .A2(n6251), .ZN(n6252) );
  XNOR2_X2 U7310 ( .A(n6252), .B(P1_IR_REG_28__SCAN_IN), .ZN(n6363) );
  XNOR2_X1 U7311 ( .A(n6253), .B(n6445), .ZN(n6362) );
  NAND2_X1 U7312 ( .A1(n6361), .A2(n6603), .ZN(n6254) );
  NAND2_X1 U7313 ( .A1(n6254), .A2(P1_STATE_REG_SCAN_IN), .ZN(P1_U3083) );
  INV_X2 U7314 ( .A(n9069), .ZN(P2_U3966) );
  INV_X2 U7315 ( .A(P1_STATE_REG_SCAN_IN), .ZN(P1_U3084) );
  NAND2_X1 U7316 ( .A1(n8933), .A2(n9317), .ZN(n8895) );
  NAND2_X1 U7317 ( .A1(n8896), .A2(n8733), .ZN(n6256) );
  OR2_X1 U7318 ( .A1(n8975), .A2(n7478), .ZN(n8793) );
  NAND2_X1 U7319 ( .A1(n8975), .A2(n7478), .ZN(n8794) );
  OR2_X1 U7320 ( .A1(n6952), .A2(n7317), .ZN(n7319) );
  NAND2_X1 U7321 ( .A1(n9068), .A2(n10505), .ZN(n8751) );
  NAND2_X1 U7322 ( .A1(n6258), .A2(n8760), .ZN(n6963) );
  INV_X1 U7323 ( .A(n8900), .ZN(n6964) );
  NAND2_X1 U7324 ( .A1(n6962), .A2(n8765), .ZN(n7303) );
  INV_X1 U7325 ( .A(n7301), .ZN(n10537) );
  NAND2_X1 U7326 ( .A1(n10537), .A2(n9066), .ZN(n8773) );
  NAND2_X1 U7327 ( .A1(n7217), .A2(n7301), .ZN(n8772) );
  NAND2_X1 U7328 ( .A1(n7303), .A2(n8903), .ZN(n7302) );
  NAND2_X1 U7329 ( .A1(n10546), .A2(n7374), .ZN(n8778) );
  INV_X1 U7330 ( .A(n10546), .ZN(n7425) );
  NAND2_X1 U7331 ( .A1(n7425), .A2(n7330), .ZN(n8777) );
  INV_X1 U7332 ( .A(n8781), .ZN(n8785) );
  OR2_X1 U7333 ( .A1(n8784), .A2(n8785), .ZN(n6260) );
  XNOR2_X1 U7334 ( .A(n8789), .B(n9065), .ZN(n8788) );
  INV_X1 U7335 ( .A(n9065), .ZN(n8970) );
  NOR2_X1 U7336 ( .A1(n8789), .A2(n8970), .ZN(n6261) );
  AOI21_X1 U7337 ( .B1(n7476), .B2(n8788), .A(n6261), .ZN(n6262) );
  OAI21_X1 U7338 ( .B1(n8908), .B2(n6262), .A(n7495), .ZN(n6263) );
  AOI222_X1 U7339 ( .A1(n9349), .A2(n6263), .B1(n5120), .B2(n9241), .C1(n9065), 
        .C2(n9239), .ZN(n6264) );
  INV_X1 U7340 ( .A(n6264), .ZN(n10589) );
  NOR2_X1 U7341 ( .A1(n6265), .A2(P2_U3152), .ZN(n6949) );
  INV_X1 U7342 ( .A(n6947), .ZN(n6266) );
  NAND3_X1 U7343 ( .A1(n6949), .A2(n6266), .A3(n6956), .ZN(n6267) );
  MUX2_X1 U7344 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n10589), .S(n9378), .Z(n6287)
         );
  NAND2_X1 U7345 ( .A1(n9365), .A2(n8754), .ZN(n9364) );
  NAND2_X1 U7346 ( .A1(n5071), .A2(n10521), .ZN(n6270) );
  NAND2_X1 U7347 ( .A1(n9364), .A2(n6270), .ZN(n6966) );
  NAND2_X1 U7348 ( .A1(n6966), .A2(n8900), .ZN(n6965) );
  NAND2_X1 U7349 ( .A1(n5157), .A2(n6974), .ZN(n6271) );
  NAND2_X1 U7350 ( .A1(n9066), .A2(n7301), .ZN(n6272) );
  AND2_X1 U7351 ( .A1(n8778), .A2(n8777), .ZN(n8775) );
  INV_X1 U7352 ( .A(n8775), .ZN(n8905) );
  NAND2_X1 U7353 ( .A1(n10546), .A2(n7330), .ZN(n6273) );
  INV_X1 U7354 ( .A(n6274), .ZN(n7337) );
  XNOR2_X1 U7355 ( .A(n8784), .B(n8785), .ZN(n8906) );
  NAND2_X1 U7356 ( .A1(n7337), .A2(n8906), .ZN(n7338) );
  NAND2_X1 U7357 ( .A1(n8784), .A2(n8781), .ZN(n8783) );
  OR2_X1 U7358 ( .A1(n8789), .A2(n9065), .ZN(n6275) );
  INV_X1 U7359 ( .A(n8908), .ZN(n6276) );
  NOR2_X1 U7360 ( .A1(n4944), .A2(n6276), .ZN(n10586) );
  INV_X1 U7361 ( .A(n7491), .ZN(n6281) );
  AND2_X1 U7362 ( .A1(n6435), .A2(n5298), .ZN(n6278) );
  NAND2_X1 U7363 ( .A1(n6279), .A2(n6175), .ZN(n6277) );
  NAND2_X1 U7364 ( .A1(n6278), .A2(n6277), .ZN(n9369) );
  OR2_X1 U7365 ( .A1(n6279), .A2(n5298), .ZN(n7347) );
  NAND2_X1 U7366 ( .A1(n9369), .A2(n7347), .ZN(n6280) );
  NOR3_X1 U7367 ( .A1(n10586), .A2(n6281), .A3(n9359), .ZN(n6286) );
  AND2_X1 U7368 ( .A1(n9378), .A2(n5298), .ZN(n9362) );
  INV_X1 U7369 ( .A(n9362), .ZN(n8093) );
  INV_X1 U7370 ( .A(n8975), .ZN(n10588) );
  NAND2_X1 U7371 ( .A1(n10505), .A2(n7317), .ZN(n9379) );
  INV_X1 U7372 ( .A(n6974), .ZN(n7348) );
  NOR2_X2 U7373 ( .A1(n7332), .A2(n8784), .ZN(n7481) );
  INV_X1 U7374 ( .A(n8789), .ZN(n10570) );
  AND2_X1 U7375 ( .A1(n7481), .A2(n10570), .ZN(n7483) );
  NAND2_X1 U7376 ( .A1(n10588), .A2(n7483), .ZN(n7500) );
  OAI211_X1 U7377 ( .C1(n10588), .C2(n7483), .A(n5299), .B(n7500), .ZN(n10587)
         );
  NOR2_X1 U7378 ( .A1(n8093), .A2(n10587), .ZN(n6285) );
  INV_X1 U7379 ( .A(n8974), .ZN(n6283) );
  OAI22_X1 U7380 ( .A1(n9333), .A2(n10588), .B1(n9316), .B2(n6283), .ZN(n6284)
         );
  OR4_X1 U7381 ( .A1(n6287), .A2(n6286), .A3(n6285), .A4(n6284), .ZN(P2_U3288)
         );
  OR2_X1 U7382 ( .A1(n6288), .A2(P1_IR_REG_10__SCAN_IN), .ZN(n6342) );
  NOR2_X1 U7383 ( .A1(n6342), .A2(P1_IR_REG_11__SCAN_IN), .ZN(n6293) );
  NOR2_X1 U7384 ( .A1(P1_IR_REG_12__SCAN_IN), .A2(P1_IR_REG_13__SCAN_IN), .ZN(
        n6289) );
  NAND2_X1 U7385 ( .A1(n6293), .A2(n6289), .ZN(n6291) );
  NAND2_X1 U7386 ( .A1(n6290), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6355) );
  XNOR2_X1 U7387 ( .A(n6355), .B(P1_IR_REG_16__SCAN_IN), .ZN(n9655) );
  NAND2_X1 U7388 ( .A1(n6291), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6292) );
  XNOR2_X1 U7389 ( .A(n6292), .B(P1_IR_REG_14__SCAN_IN), .ZN(n7858) );
  OR2_X1 U7390 ( .A1(n6293), .A2(n6318), .ZN(n6296) );
  NAND2_X1 U7391 ( .A1(n6296), .A2(n6294), .ZN(n6298) );
  NAND2_X1 U7392 ( .A1(n6298), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6295) );
  XNOR2_X1 U7393 ( .A(n6295), .B(P1_IR_REG_13__SCAN_IN), .ZN(n7852) );
  INV_X1 U7394 ( .A(n6296), .ZN(n6297) );
  NAND2_X1 U7395 ( .A1(n6297), .A2(P1_IR_REG_12__SCAN_IN), .ZN(n6299) );
  NAND2_X1 U7396 ( .A1(n6288), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6300) );
  XNOR2_X1 U7397 ( .A(n6300), .B(P1_IR_REG_10__SCAN_IN), .ZN(n7645) );
  NAND2_X1 U7398 ( .A1(P1_REG2_REG_10__SCAN_IN), .A2(n7645), .ZN(n6341) );
  INV_X1 U7399 ( .A(P1_REG2_REG_10__SCAN_IN), .ZN(n6301) );
  MUX2_X1 U7400 ( .A(n6301), .B(P1_REG2_REG_10__SCAN_IN), .S(n7645), .Z(n6302)
         );
  INV_X1 U7401 ( .A(n6302), .ZN(n6816) );
  OR2_X1 U7402 ( .A1(n6303), .A2(n6318), .ZN(n6308) );
  INV_X1 U7403 ( .A(P1_IR_REG_8__SCAN_IN), .ZN(n6304) );
  NAND2_X1 U7404 ( .A1(n6308), .A2(n6304), .ZN(n6310) );
  NAND2_X1 U7405 ( .A1(n6310), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6305) );
  XNOR2_X1 U7406 ( .A(n6305), .B(P1_IR_REG_9__SCAN_IN), .ZN(n7512) );
  NAND2_X1 U7407 ( .A1(n7512), .A2(P1_REG2_REG_9__SCAN_IN), .ZN(n6340) );
  INV_X1 U7408 ( .A(P1_REG2_REG_9__SCAN_IN), .ZN(n6306) );
  MUX2_X1 U7409 ( .A(n6306), .B(P1_REG2_REG_9__SCAN_IN), .S(n7512), .Z(n6307)
         );
  INV_X1 U7410 ( .A(n6307), .ZN(n10402) );
  INV_X1 U7411 ( .A(n6308), .ZN(n6309) );
  NAND2_X1 U7412 ( .A1(n6309), .A2(P1_IR_REG_8__SCAN_IN), .ZN(n6311) );
  INV_X1 U7413 ( .A(n7441), .ZN(n6523) );
  INV_X1 U7414 ( .A(P1_REG2_REG_8__SCAN_IN), .ZN(n6339) );
  NAND2_X1 U7415 ( .A1(n6312), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6313) );
  XNOR2_X1 U7416 ( .A(n6313), .B(P1_IR_REG_7__SCAN_IN), .ZN(n7196) );
  NOR2_X1 U7417 ( .A1(n7196), .A2(P1_REG2_REG_7__SCAN_IN), .ZN(n6338) );
  NAND2_X1 U7418 ( .A1(n6314), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6315) );
  MUX2_X1 U7419 ( .A(P1_IR_REG_31__SCAN_IN), .B(n6315), .S(
        P1_IR_REG_6__SCAN_IN), .Z(n6316) );
  AND2_X1 U7420 ( .A1(n6312), .A2(n6316), .ZN(n7129) );
  INV_X1 U7421 ( .A(n7129), .ZN(n6409) );
  INV_X1 U7422 ( .A(P1_REG2_REG_6__SCAN_IN), .ZN(n7178) );
  OR2_X1 U7423 ( .A1(n6317), .A2(n6318), .ZN(n6328) );
  OR2_X1 U7424 ( .A1(n6319), .A2(n6318), .ZN(n6320) );
  AND2_X1 U7425 ( .A1(n6328), .A2(n6320), .ZN(n6331) );
  INV_X1 U7426 ( .A(P1_IR_REG_4__SCAN_IN), .ZN(n6321) );
  NAND2_X1 U7427 ( .A1(n6331), .A2(n6321), .ZN(n6334) );
  NAND2_X1 U7428 ( .A1(n6334), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6322) );
  XNOR2_X1 U7429 ( .A(n6322), .B(P1_IR_REG_5__SCAN_IN), .ZN(n7026) );
  INV_X1 U7430 ( .A(P1_IR_REG_2__SCAN_IN), .ZN(n6327) );
  NAND2_X1 U7431 ( .A1(n6328), .A2(n6327), .ZN(n6326) );
  NAND2_X1 U7432 ( .A1(n6326), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6323) );
  XNOR2_X1 U7433 ( .A(n6323), .B(P1_IR_REG_3__SCAN_IN), .ZN(n6769) );
  INV_X1 U7434 ( .A(P1_IR_REG_1__SCAN_IN), .ZN(n6325) );
  NAND2_X1 U7435 ( .A1(P1_IR_REG_31__SCAN_IN), .A2(P1_IR_REG_0__SCAN_IN), .ZN(
        n6324) );
  INV_X1 U7436 ( .A(n6602), .ZN(n6370) );
  XNOR2_X1 U7437 ( .A(n6602), .B(P1_REG2_REG_1__SCAN_IN), .ZN(n6552) );
  AND3_X1 U7438 ( .A1(n6552), .A2(P1_IR_REG_0__SCAN_IN), .A3(
        P1_REG2_REG_0__SCAN_IN), .ZN(n6549) );
  AOI21_X1 U7439 ( .B1(n6370), .B2(P1_REG2_REG_1__SCAN_IN), .A(n6549), .ZN(
        n6568) );
  INV_X1 U7440 ( .A(P1_REG2_REG_2__SCAN_IN), .ZN(n6329) );
  OAI21_X1 U7441 ( .B1(n6328), .B2(n6327), .A(n6326), .ZN(n6793) );
  MUX2_X1 U7442 ( .A(P1_REG2_REG_2__SCAN_IN), .B(n6329), .S(n6793), .Z(n6567)
         );
  INV_X1 U7443 ( .A(n6793), .ZN(n6577) );
  NAND2_X1 U7444 ( .A1(n6577), .A2(P1_REG2_REG_2__SCAN_IN), .ZN(n6534) );
  INV_X1 U7445 ( .A(P1_REG2_REG_3__SCAN_IN), .ZN(n6330) );
  MUX2_X1 U7446 ( .A(n6330), .B(P1_REG2_REG_3__SCAN_IN), .S(n6769), .Z(n6533)
         );
  AOI21_X1 U7447 ( .B1(n6565), .B2(n6534), .A(n6533), .ZN(n6532) );
  AOI21_X1 U7448 ( .B1(P1_REG2_REG_3__SCAN_IN), .B2(n6769), .A(n6532), .ZN(
        n9640) );
  INV_X1 U7449 ( .A(P1_REG2_REG_4__SCAN_IN), .ZN(n6335) );
  INV_X1 U7450 ( .A(n6331), .ZN(n6332) );
  NAND2_X1 U7451 ( .A1(n6332), .A2(P1_IR_REG_4__SCAN_IN), .ZN(n6333) );
  MUX2_X1 U7452 ( .A(P1_REG2_REG_4__SCAN_IN), .B(n6335), .S(n9643), .Z(n9641)
         );
  INV_X1 U7453 ( .A(n9639), .ZN(n6336) );
  NOR2_X1 U7454 ( .A1(n9643), .A2(P1_REG2_REG_4__SCAN_IN), .ZN(n6506) );
  INV_X1 U7455 ( .A(P1_REG2_REG_5__SCAN_IN), .ZN(n7120) );
  MUX2_X1 U7456 ( .A(P1_REG2_REG_5__SCAN_IN), .B(n7120), .S(n7026), .Z(n6505)
         );
  OAI21_X1 U7457 ( .B1(n6336), .B2(n6506), .A(n6505), .ZN(n6510) );
  OAI21_X1 U7458 ( .B1(P1_REG2_REG_5__SCAN_IN), .B2(n7026), .A(n6510), .ZN(
        n6561) );
  MUX2_X1 U7459 ( .A(n7178), .B(P1_REG2_REG_6__SCAN_IN), .S(n7129), .Z(n6560)
         );
  INV_X1 U7460 ( .A(n6559), .ZN(n6337) );
  OAI21_X1 U7461 ( .B1(n6409), .B2(n7178), .A(n6337), .ZN(n6456) );
  INV_X1 U7462 ( .A(P1_REG2_REG_7__SCAN_IN), .ZN(n7145) );
  MUX2_X1 U7463 ( .A(n7145), .B(P1_REG2_REG_7__SCAN_IN), .S(n7196), .Z(n6457)
         );
  NOR2_X1 U7464 ( .A1(n6456), .A2(n6457), .ZN(n6455) );
  NOR2_X1 U7465 ( .A1(n6338), .A2(n6455), .ZN(n6517) );
  MUX2_X1 U7466 ( .A(n6339), .B(P1_REG2_REG_8__SCAN_IN), .S(n7441), .Z(n6516)
         );
  NOR2_X1 U7467 ( .A1(n6517), .A2(n6516), .ZN(n6515) );
  AOI21_X1 U7468 ( .B1(n6523), .B2(n6339), .A(n6515), .ZN(n10403) );
  NAND2_X1 U7469 ( .A1(n10402), .A2(n10403), .ZN(n10400) );
  NAND2_X1 U7470 ( .A1(n6340), .A2(n10400), .ZN(n6817) );
  NAND2_X1 U7471 ( .A1(n6816), .A2(n6817), .ZN(n6815) );
  NAND2_X1 U7472 ( .A1(P1_REG2_REG_11__SCAN_IN), .A2(n6881), .ZN(n6885) );
  INV_X1 U7473 ( .A(n6885), .ZN(n6344) );
  NAND2_X1 U7474 ( .A1(n6342), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6343) );
  XNOR2_X1 U7475 ( .A(n6343), .B(P1_IR_REG_11__SCAN_IN), .ZN(n7651) );
  OAI22_X1 U7476 ( .A1(n6344), .A2(n7651), .B1(P1_REG2_REG_11__SCAN_IN), .B2(
        n6881), .ZN(n7103) );
  INV_X1 U7477 ( .A(P1_REG2_REG_12__SCAN_IN), .ZN(n6345) );
  MUX2_X1 U7478 ( .A(P1_REG2_REG_12__SCAN_IN), .B(n6345), .S(n7730), .Z(n6346)
         );
  INV_X1 U7479 ( .A(n6346), .ZN(n7102) );
  AOI21_X1 U7480 ( .B1(n7730), .B2(P1_REG2_REG_12__SCAN_IN), .A(n7101), .ZN(
        n7270) );
  NAND2_X1 U7481 ( .A1(P1_REG2_REG_13__SCAN_IN), .A2(n7852), .ZN(n6347) );
  OAI21_X1 U7482 ( .B1(n7852), .B2(P1_REG2_REG_13__SCAN_IN), .A(n6347), .ZN(
        n7269) );
  AOI21_X1 U7483 ( .B1(n7852), .B2(P1_REG2_REG_13__SCAN_IN), .A(n7268), .ZN(
        n7429) );
  NAND2_X1 U7484 ( .A1(n7858), .A2(P1_REG2_REG_14__SCAN_IN), .ZN(n6348) );
  OAI21_X1 U7485 ( .B1(n7858), .B2(P1_REG2_REG_14__SCAN_IN), .A(n6348), .ZN(
        n7428) );
  AOI21_X1 U7486 ( .B1(P1_REG2_REG_14__SCAN_IN), .B2(n7858), .A(n7427), .ZN(
        n6351) );
  NAND2_X1 U7487 ( .A1(n6349), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6350) );
  XNOR2_X1 U7488 ( .A(n6350), .B(P1_IR_REG_15__SCAN_IN), .ZN(n8007) );
  INV_X1 U7489 ( .A(n8007), .ZN(n6892) );
  NOR2_X1 U7490 ( .A1(n6351), .A2(n6892), .ZN(n6352) );
  INV_X1 U7491 ( .A(P1_REG2_REG_15__SCAN_IN), .ZN(n7778) );
  NOR2_X1 U7492 ( .A1(n7778), .A2(n7779), .ZN(n7777) );
  NAND2_X1 U7493 ( .A1(P1_REG2_REG_16__SCAN_IN), .A2(n9655), .ZN(n6353) );
  OAI21_X1 U7494 ( .B1(n9655), .B2(P1_REG2_REG_16__SCAN_IN), .A(n6353), .ZN(
        n9648) );
  NOR2_X1 U7495 ( .A1(n9649), .A2(n9648), .ZN(n9647) );
  INV_X1 U7496 ( .A(P1_REG2_REG_17__SCAN_IN), .ZN(n6359) );
  NAND2_X1 U7497 ( .A1(n6355), .A2(n6354), .ZN(n6356) );
  NAND2_X1 U7498 ( .A1(n6356), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6358) );
  NAND2_X1 U7499 ( .A1(n6358), .A2(n6357), .ZN(n7185) );
  OAI21_X1 U7500 ( .B1(n6358), .B2(n6357), .A(n7185), .ZN(n9670) );
  MUX2_X1 U7501 ( .A(n6359), .B(P1_REG2_REG_17__SCAN_IN), .S(n9670), .Z(n6360)
         );
  INV_X1 U7502 ( .A(n6360), .ZN(n6364) );
  NOR2_X1 U7503 ( .A1(n6365), .A2(n6364), .ZN(n9671) );
  NAND2_X1 U7504 ( .A1(n6361), .A2(P1_STATE_REG_SCAN_IN), .ZN(n10375) );
  OR2_X1 U7505 ( .A1(n10375), .A2(n4860), .ZN(n10374) );
  AOI211_X1 U7506 ( .C1(n6365), .C2(n6364), .A(n9671), .B(n9673), .ZN(n6389)
         );
  INV_X1 U7507 ( .A(P1_REG3_REG_17__SCAN_IN), .ZN(n8146) );
  NOR2_X1 U7508 ( .A1(n8146), .A2(P1_STATE_REG_SCAN_IN), .ZN(n9547) );
  INV_X1 U7509 ( .A(n6363), .ZN(n10376) );
  INV_X1 U7510 ( .A(n6762), .ZN(n7784) );
  NOR2_X1 U7511 ( .A1(n6581), .A2(n7784), .ZN(n6366) );
  INV_X1 U7512 ( .A(P1_ADDR_REG_17__SCAN_IN), .ZN(n6367) );
  OAI22_X1 U7513 ( .A1(n10393), .A2(n9670), .B1(n10391), .B2(n6367), .ZN(n6388) );
  XNOR2_X1 U7514 ( .A(n9670), .B(P1_REG1_REG_17__SCAN_IN), .ZN(n6385) );
  INV_X1 U7515 ( .A(n9655), .ZN(n6383) );
  INV_X1 U7516 ( .A(P1_REG1_REG_16__SCAN_IN), .ZN(n6382) );
  XOR2_X1 U7517 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n9655), .Z(n9657) );
  INV_X1 U7518 ( .A(n7858), .ZN(n6706) );
  INV_X1 U7519 ( .A(P1_REG1_REG_14__SCAN_IN), .ZN(n6379) );
  INV_X1 U7520 ( .A(n7852), .ZN(n6378) );
  INV_X1 U7521 ( .A(P1_REG1_REG_13__SCAN_IN), .ZN(n6377) );
  INV_X1 U7522 ( .A(n7730), .ZN(n6376) );
  INV_X1 U7523 ( .A(P1_REG1_REG_12__SCAN_IN), .ZN(n6375) );
  INV_X1 U7524 ( .A(P1_REG1_REG_10__SCAN_IN), .ZN(n6368) );
  MUX2_X1 U7525 ( .A(P1_REG1_REG_10__SCAN_IN), .B(n6368), .S(n7645), .Z(n6822)
         );
  INV_X1 U7526 ( .A(P1_REG1_REG_9__SCAN_IN), .ZN(n10602) );
  INV_X1 U7527 ( .A(n7512), .ZN(n10392) );
  AOI22_X1 U7528 ( .A1(n7512), .A2(P1_REG1_REG_9__SCAN_IN), .B1(n10602), .B2(
        n10392), .ZN(n10396) );
  INV_X1 U7529 ( .A(P1_REG1_REG_8__SCAN_IN), .ZN(n6369) );
  MUX2_X1 U7530 ( .A(P1_REG1_REG_8__SCAN_IN), .B(n6369), .S(n7441), .Z(n6519)
         );
  XOR2_X1 U7531 ( .A(P1_REG1_REG_1__SCAN_IN), .B(n6602), .Z(n6545) );
  INV_X1 U7532 ( .A(P1_IR_REG_0__SCAN_IN), .ZN(n10383) );
  INV_X1 U7533 ( .A(P1_REG1_REG_0__SCAN_IN), .ZN(n10382) );
  NOR3_X1 U7534 ( .A1(n6545), .A2(n10383), .A3(n10382), .ZN(n6544) );
  AOI21_X1 U7535 ( .B1(n6370), .B2(P1_REG1_REG_1__SCAN_IN), .A(n6544), .ZN(
        n6571) );
  INV_X1 U7536 ( .A(P1_REG1_REG_2__SCAN_IN), .ZN(n6371) );
  MUX2_X1 U7537 ( .A(P1_REG1_REG_2__SCAN_IN), .B(n6371), .S(n6793), .Z(n6570)
         );
  NOR2_X1 U7538 ( .A1(n6571), .A2(n6570), .ZN(n6569) );
  AOI21_X1 U7539 ( .B1(P1_REG1_REG_2__SCAN_IN), .B2(n6577), .A(n6569), .ZN(
        n6530) );
  XNOR2_X1 U7540 ( .A(n6769), .B(P1_REG1_REG_3__SCAN_IN), .ZN(n6529) );
  NOR2_X1 U7541 ( .A1(n6530), .A2(n6529), .ZN(n6528) );
  AOI21_X1 U7542 ( .B1(P1_REG1_REG_3__SCAN_IN), .B2(n6769), .A(n6528), .ZN(
        n9634) );
  INV_X1 U7543 ( .A(P1_REG1_REG_4__SCAN_IN), .ZN(n6372) );
  MUX2_X1 U7544 ( .A(P1_REG1_REG_4__SCAN_IN), .B(n6372), .S(n9643), .Z(n9633)
         );
  NAND2_X1 U7545 ( .A1(n9634), .A2(n9633), .ZN(n9632) );
  OAI21_X1 U7546 ( .B1(P1_REG1_REG_4__SCAN_IN), .B2(n9643), .A(n9632), .ZN(
        n6502) );
  XNOR2_X1 U7547 ( .A(n7026), .B(P1_REG1_REG_5__SCAN_IN), .ZN(n6503) );
  NOR2_X1 U7548 ( .A1(n6502), .A2(n6503), .ZN(n6501) );
  AOI21_X1 U7549 ( .B1(n7026), .B2(P1_REG1_REG_5__SCAN_IN), .A(n6501), .ZN(
        n6557) );
  XNOR2_X1 U7550 ( .A(n7129), .B(P1_REG1_REG_6__SCAN_IN), .ZN(n6556) );
  NOR2_X1 U7551 ( .A1(n6557), .A2(n6556), .ZN(n6555) );
  AOI21_X1 U7552 ( .B1(n7129), .B2(P1_REG1_REG_6__SCAN_IN), .A(n6555), .ZN(
        n6460) );
  NOR2_X1 U7553 ( .A1(n7196), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n6373) );
  AOI21_X1 U7554 ( .B1(n7196), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6373), .ZN(
        n6459) );
  NAND2_X1 U7555 ( .A1(n6460), .A2(n6459), .ZN(n6458) );
  OAI21_X1 U7556 ( .B1(n7196), .B2(P1_REG1_REG_7__SCAN_IN), .A(n6458), .ZN(
        n6520) );
  NAND2_X1 U7557 ( .A1(n6519), .A2(n6520), .ZN(n6518) );
  OAI21_X1 U7558 ( .B1(P1_REG1_REG_8__SCAN_IN), .B2(n7441), .A(n6518), .ZN(
        n10397) );
  NAND2_X1 U7559 ( .A1(n10396), .A2(n10397), .ZN(n10395) );
  OAI21_X1 U7560 ( .B1(P1_REG1_REG_9__SCAN_IN), .B2(n7512), .A(n10395), .ZN(
        n6823) );
  NAND2_X1 U7561 ( .A1(n6822), .A2(n6823), .ZN(n6821) );
  OAI21_X1 U7562 ( .B1(P1_REG1_REG_10__SCAN_IN), .B2(n7645), .A(n6821), .ZN(
        n6879) );
  NOR2_X1 U7563 ( .A1(P1_REG1_REG_11__SCAN_IN), .A2(n7651), .ZN(n6878) );
  NAND2_X1 U7564 ( .A1(n7651), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n6374) );
  OAI21_X1 U7565 ( .B1(n6879), .B2(n6878), .A(n6374), .ZN(n7095) );
  XNOR2_X1 U7566 ( .A(n7730), .B(P1_REG1_REG_12__SCAN_IN), .ZN(n7096) );
  NOR2_X1 U7567 ( .A1(n7095), .A2(n7096), .ZN(n7094) );
  AOI21_X1 U7568 ( .B1(n6376), .B2(n6375), .A(n7094), .ZN(n7273) );
  XNOR2_X1 U7569 ( .A(n7852), .B(P1_REG1_REG_13__SCAN_IN), .ZN(n7274) );
  NOR2_X1 U7570 ( .A1(n7273), .A2(n7274), .ZN(n7272) );
  AOI21_X1 U7571 ( .B1(n6378), .B2(n6377), .A(n7272), .ZN(n7433) );
  XNOR2_X1 U7572 ( .A(n7858), .B(P1_REG1_REG_14__SCAN_IN), .ZN(n7432) );
  NOR2_X1 U7573 ( .A1(n7433), .A2(n7432), .ZN(n7431) );
  AOI21_X1 U7574 ( .B1(n6706), .B2(n6379), .A(n7431), .ZN(n6380) );
  NAND2_X1 U7575 ( .A1(n8007), .A2(n6380), .ZN(n6381) );
  XNOR2_X1 U7576 ( .A(n6892), .B(n6380), .ZN(n7774) );
  NAND2_X1 U7577 ( .A1(P1_REG1_REG_15__SCAN_IN), .A2(n7774), .ZN(n7773) );
  NAND2_X1 U7578 ( .A1(n6381), .A2(n7773), .ZN(n9658) );
  NAND2_X1 U7579 ( .A1(n9657), .A2(n9658), .ZN(n9656) );
  OAI21_X1 U7580 ( .B1(n6383), .B2(n6382), .A(n9656), .ZN(n6384) );
  INV_X1 U7581 ( .A(n4860), .ZN(n6592) );
  OR3_X1 U7582 ( .A1(n10375), .A2(n6363), .A3(n6592), .ZN(n10380) );
  INV_X1 U7583 ( .A(n10380), .ZN(n10398) );
  NAND2_X1 U7584 ( .A1(n6385), .A2(n6384), .ZN(n9662) );
  OAI211_X1 U7585 ( .C1(n6385), .C2(n6384), .A(n10398), .B(n9662), .ZN(n6386)
         );
  INV_X1 U7586 ( .A(n6386), .ZN(n6387) );
  OR4_X1 U7587 ( .A1(n6389), .A2(n9547), .A3(n6388), .A4(n6387), .ZN(P1_U3258)
         );
  INV_X1 U7588 ( .A(n9487), .ZN(n9491) );
  AND2_X1 U7589 ( .A1(n6597), .A2(P2_U3152), .ZN(n7786) );
  OAI222_X1 U7590 ( .A1(n9491), .A2(n6391), .B1(n4857), .B2(n6599), .C1(
        P2_U3152), .C2(n6390), .ZN(P2_U3357) );
  OAI222_X1 U7591 ( .A1(n9491), .A2(n5556), .B1(n4857), .B2(n6791), .C1(
        P2_U3152), .C2(n10435), .ZN(P2_U3356) );
  INV_X1 U7592 ( .A(n6770), .ZN(n6406) );
  AOI22_X1 U7593 ( .A1(n10448), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_3__SCAN_IN), .B2(n9487), .ZN(n6392) );
  OAI21_X1 U7594 ( .B1(n6406), .B2(n4857), .A(n6392), .ZN(P2_U3355) );
  NAND2_X1 U7595 ( .A1(n6581), .A2(n6393), .ZN(n8597) );
  INV_X1 U7596 ( .A(P1_D_REG_1__SCAN_IN), .ZN(n6400) );
  NAND3_X1 U7597 ( .A1(n7964), .A2(P1_B_REG_SCAN_IN), .A3(n7808), .ZN(n6395)
         );
  OAI21_X1 U7598 ( .B1(P1_B_REG_SCAN_IN), .B2(n7808), .A(n6395), .ZN(n6396) );
  OR2_X1 U7599 ( .A1(n10046), .A2(P1_D_REG_1__SCAN_IN), .ZN(n6398) );
  NAND2_X1 U7600 ( .A1(n6394), .A2(n7964), .ZN(n6397) );
  NAND2_X1 U7601 ( .A1(n6920), .A2(n10047), .ZN(n6399) );
  OAI21_X1 U7602 ( .B1(n10047), .B2(n6400), .A(n6399), .ZN(P1_U3441) );
  INV_X1 U7603 ( .A(P1_D_REG_0__SCAN_IN), .ZN(n6404) );
  NAND2_X1 U7604 ( .A1(n6394), .A2(n7808), .ZN(n6401) );
  NAND2_X1 U7605 ( .A1(n6743), .A2(n10047), .ZN(n6403) );
  OAI21_X1 U7606 ( .B1(n10047), .B2(n6404), .A(n6403), .ZN(P1_U3440) );
  INV_X1 U7607 ( .A(P1_DATAO_REG_4__SCAN_IN), .ZN(n6405) );
  INV_X1 U7608 ( .A(n6659), .ZN(n6761) );
  OAI222_X1 U7609 ( .A1(n9491), .A2(n6405), .B1(n4857), .B2(n6841), .C1(
        P2_U3152), .C2(n6761), .ZN(P2_U3354) );
  INV_X1 U7610 ( .A(P2_DATAO_REG_1__SCAN_IN), .ZN(n6598) );
  NAND2_X1 U7611 ( .A1(n8387), .A2(P1_U3084), .ZN(n10033) );
  OAI222_X1 U7612 ( .A1(n10039), .A2(n6598), .B1(n6602), .B2(P1_U3084), .C1(
        n10033), .C2(n6599), .ZN(P1_U3352) );
  INV_X1 U7613 ( .A(n6769), .ZN(n6539) );
  OAI222_X1 U7614 ( .A1(n10033), .A2(n6406), .B1(n10039), .B2(n4963), .C1(
        P1_U3084), .C2(n6539), .ZN(P1_U3350) );
  INV_X1 U7615 ( .A(P1_DATAO_REG_5__SCAN_IN), .ZN(n6407) );
  INV_X1 U7616 ( .A(n10462), .ZN(n6666) );
  OAI222_X1 U7617 ( .A1(n9491), .A2(n6407), .B1(n4857), .B2(n7025), .C1(
        P2_U3152), .C2(n6666), .ZN(P2_U3353) );
  INV_X1 U7618 ( .A(n10033), .ZN(n7783) );
  INV_X1 U7619 ( .A(n7783), .ZN(n10043) );
  INV_X1 U7620 ( .A(P2_DATAO_REG_5__SCAN_IN), .ZN(n6429) );
  INV_X1 U7621 ( .A(n7026), .ZN(n6408) );
  OAI222_X1 U7622 ( .A1(n10043), .A2(n7025), .B1(n10039), .B2(n6429), .C1(
        P1_U3084), .C2(n6408), .ZN(P1_U3348) );
  INV_X1 U7623 ( .A(P2_DATAO_REG_6__SCAN_IN), .ZN(n6431) );
  OAI222_X1 U7624 ( .A1(n10043), .A2(n7128), .B1(n10039), .B2(n6431), .C1(
        P1_U3084), .C2(n6409), .ZN(P1_U3347) );
  INV_X1 U7625 ( .A(P2_DATAO_REG_2__SCAN_IN), .ZN(n6790) );
  OAI222_X1 U7626 ( .A1(n10039), .A2(n6790), .B1(n6793), .B2(P1_U3084), .C1(
        n10043), .C2(n6791), .ZN(P1_U3351) );
  INV_X1 U7627 ( .A(P1_DATAO_REG_6__SCAN_IN), .ZN(n6410) );
  INV_X1 U7628 ( .A(n10477), .ZN(n6668) );
  OAI222_X1 U7629 ( .A1(n9491), .A2(n6410), .B1(n4857), .B2(n7128), .C1(
        P2_U3152), .C2(n6668), .ZN(P2_U3352) );
  INV_X1 U7630 ( .A(n10039), .ZN(n7017) );
  AOI22_X1 U7631 ( .A1(P2_DATAO_REG_4__SCAN_IN), .A2(n7017), .B1(n9643), .B2(
        P1_STATE_REG_SCAN_IN), .ZN(n6411) );
  OAI21_X1 U7632 ( .B1(n6841), .B2(n10033), .A(n6411), .ZN(P1_U3349) );
  AOI22_X1 U7633 ( .A1(n7196), .A2(P1_STATE_REG_SCAN_IN), .B1(n7017), .B2(
        P2_DATAO_REG_7__SCAN_IN), .ZN(n6412) );
  OAI21_X1 U7634 ( .B1(n7195), .B2(n10033), .A(n6412), .ZN(P1_U3346) );
  INV_X1 U7635 ( .A(n6670), .ZN(n6691) );
  INV_X1 U7636 ( .A(P1_DATAO_REG_7__SCAN_IN), .ZN(n6413) );
  OAI222_X1 U7637 ( .A1(P2_U3152), .A2(n6691), .B1(n4857), .B2(n7195), .C1(
        n6413), .C2(n9491), .ZN(P2_U3351) );
  INV_X1 U7638 ( .A(n7440), .ZN(n6415) );
  AOI22_X1 U7639 ( .A1(n7441), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_8__SCAN_IN), .B2(n7017), .ZN(n6414) );
  OAI21_X1 U7640 ( .B1(n6415), .B2(n10033), .A(n6414), .ZN(P1_U3345) );
  INV_X1 U7641 ( .A(P1_DATAO_REG_8__SCAN_IN), .ZN(n6416) );
  INV_X1 U7642 ( .A(n6707), .ZN(n6719) );
  OAI222_X1 U7643 ( .A1(n9491), .A2(n6416), .B1(n4857), .B2(n6415), .C1(n6719), 
        .C2(P2_U3152), .ZN(P2_U3350) );
  INV_X1 U7644 ( .A(n7511), .ZN(n6427) );
  AOI22_X1 U7645 ( .A1(n6728), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_9__SCAN_IN), .B2(n9487), .ZN(n6417) );
  OAI21_X1 U7646 ( .B1(n6427), .B2(n4857), .A(n6417), .ZN(P2_U3349) );
  INV_X1 U7647 ( .A(P2_DATAO_REG_31__SCAN_IN), .ZN(n6424) );
  NAND2_X1 U7648 ( .A1(n6418), .A2(P2_REG1_REG_31__SCAN_IN), .ZN(n6422) );
  NAND2_X1 U7649 ( .A1(n5589), .A2(P2_REG2_REG_31__SCAN_IN), .ZN(n6421) );
  NAND2_X1 U7650 ( .A1(n6419), .A2(P2_REG0_REG_31__SCAN_IN), .ZN(n6420) );
  AND3_X1 U7651 ( .A1(n6422), .A2(n6421), .A3(n6420), .ZN(n9114) );
  INV_X1 U7652 ( .A(n9114), .ZN(n8722) );
  NAND2_X1 U7653 ( .A1(n8722), .A2(P2_U3966), .ZN(n6423) );
  OAI21_X1 U7654 ( .B1(n6424), .B2(P2_U3966), .A(n6423), .ZN(P2_U3583) );
  NAND2_X1 U7655 ( .A1(n6259), .A2(P2_U3966), .ZN(n6425) );
  OAI21_X1 U7656 ( .B1(n4963), .B2(P2_U3966), .A(n6425), .ZN(P2_U3555) );
  INV_X1 U7657 ( .A(P2_DATAO_REG_9__SCAN_IN), .ZN(n6426) );
  OAI222_X1 U7658 ( .A1(n10043), .A2(n6427), .B1(n10392), .B2(P1_U3084), .C1(
        n6426), .C2(n10039), .ZN(P1_U3344) );
  NAND2_X1 U7659 ( .A1(n7374), .A2(P2_U3966), .ZN(n6428) );
  OAI21_X1 U7660 ( .B1(n6429), .B2(P2_U3966), .A(n6428), .ZN(P2_U3557) );
  NAND2_X1 U7661 ( .A1(n8781), .A2(P2_U3966), .ZN(n6430) );
  OAI21_X1 U7662 ( .B1(n6431), .B2(P2_U3966), .A(n6430), .ZN(P2_U3558) );
  OR2_X1 U7663 ( .A1(n6432), .A2(P2_U3152), .ZN(n8935) );
  NAND2_X1 U7664 ( .A1(n10050), .A2(n8935), .ZN(n6434) );
  NAND2_X1 U7665 ( .A1(n6434), .A2(n6433), .ZN(n6437) );
  OR2_X1 U7666 ( .A1(n10050), .A2(n6435), .ZN(n6436) );
  NOR2_X1 U7667 ( .A1(n10486), .A2(P2_U3966), .ZN(P2_U3151) );
  INV_X1 U7668 ( .A(n7644), .ZN(n6440) );
  AOI22_X1 U7669 ( .A1(n6863), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_10__SCAN_IN), .B2(n9487), .ZN(n6438) );
  OAI21_X1 U7670 ( .B1(n6440), .B2(n4857), .A(n6438), .ZN(P2_U3348) );
  AOI22_X1 U7671 ( .A1(n7645), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_10__SCAN_IN), .B2(n7017), .ZN(n6439) );
  OAI21_X1 U7672 ( .B1(n6440), .B2(n10033), .A(n6439), .ZN(P1_U3343) );
  AOI22_X1 U7673 ( .A1(n6868), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_11__SCAN_IN), .B2(n9487), .ZN(n6441) );
  OAI21_X1 U7674 ( .B1(n7650), .B2(n4857), .A(n6441), .ZN(P2_U3347) );
  CLKBUF_X1 U7675 ( .A(P1_U4006), .Z(n9627) );
  INV_X1 U7676 ( .A(P1_DATAO_REG_31__SCAN_IN), .ZN(n6453) );
  NOR2_X1 U7677 ( .A1(P1_IR_REG_27__SCAN_IN), .A2(P1_IR_REG_29__SCAN_IN), .ZN(
        n6442) );
  INV_X1 U7678 ( .A(P1_IR_REG_27__SCAN_IN), .ZN(n6445) );
  INV_X1 U7679 ( .A(n6774), .ZN(n8341) );
  INV_X1 U7680 ( .A(P1_REG1_REG_31__SCAN_IN), .ZN(n6451) );
  NAND2_X1 U7681 ( .A1(n6775), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n6450) );
  NAND2_X1 U7682 ( .A1(n5475), .A2(P1_REG0_REG_31__SCAN_IN), .ZN(n6449) );
  OAI211_X1 U7683 ( .C1(n8341), .C2(n6451), .A(n6450), .B(n6449), .ZN(n9695)
         );
  NAND2_X1 U7684 ( .A1(n9695), .A2(n9627), .ZN(n6452) );
  OAI21_X1 U7685 ( .B1(n9627), .B2(n6453), .A(n6452), .ZN(P1_U3586) );
  INV_X1 U7686 ( .A(n7651), .ZN(n6882) );
  INV_X1 U7687 ( .A(P2_DATAO_REG_11__SCAN_IN), .ZN(n6454) );
  OAI222_X1 U7688 ( .A1(n10043), .A2(n7650), .B1(n6882), .B2(P1_U3084), .C1(
        n6454), .C2(n10039), .ZN(P1_U3342) );
  AOI21_X1 U7689 ( .B1(n6457), .B2(n6456), .A(n6455), .ZN(n6466) );
  OAI21_X1 U7690 ( .B1(n6460), .B2(n6459), .A(n6458), .ZN(n6461) );
  NAND2_X1 U7691 ( .A1(n6461), .A2(n10398), .ZN(n6465) );
  INV_X1 U7692 ( .A(n10391), .ZN(n10386) );
  AND2_X1 U7693 ( .A1(P1_U3084), .A2(P1_REG3_REG_7__SCAN_IN), .ZN(n7287) );
  INV_X1 U7694 ( .A(n7196), .ZN(n6462) );
  NOR2_X1 U7695 ( .A1(n10393), .A2(n6462), .ZN(n6463) );
  AOI211_X1 U7696 ( .C1(n10386), .C2(P1_ADDR_REG_7__SCAN_IN), .A(n7287), .B(
        n6463), .ZN(n6464) );
  OAI211_X1 U7697 ( .C1(n6466), .C2(n9673), .A(n6465), .B(n6464), .ZN(P1_U3248) );
  NAND2_X1 U7698 ( .A1(n8387), .A2(SI_0_), .ZN(n6468) );
  XNOR2_X1 U7699 ( .A(n6468), .B(n6467), .ZN(n10044) );
  INV_X1 U7700 ( .A(n6989), .ZN(n6983) );
  NAND2_X1 U7701 ( .A1(n6607), .A2(n4855), .ZN(n6934) );
  INV_X1 U7702 ( .A(n6934), .ZN(n6486) );
  NAND2_X1 U7703 ( .A1(n5475), .A2(P1_REG0_REG_0__SCAN_IN), .ZN(n6475) );
  NAND2_X1 U7704 ( .A1(n4856), .A2(P1_REG3_REG_0__SCAN_IN), .ZN(n6474) );
  NAND2_X1 U7705 ( .A1(n6774), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6473) );
  NOR2_X1 U7706 ( .A1(n9631), .A2(n6989), .ZN(n6991) );
  INV_X1 U7707 ( .A(n9631), .ZN(n6476) );
  NOR2_X1 U7708 ( .A1(n6476), .A2(n6983), .ZN(n8559) );
  NOR2_X1 U7709 ( .A1(n6991), .A2(n8559), .ZN(n8357) );
  INV_X1 U7710 ( .A(n6478), .ZN(n6479) );
  NAND2_X1 U7711 ( .A1(n6479), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n6480) );
  NAND2_X1 U7712 ( .A1(n6579), .A2(n6904), .ZN(n8596) );
  OR2_X1 U7713 ( .A1(n8553), .A2(n8596), .ZN(n7107) );
  NAND2_X1 U7714 ( .A1(n7107), .A2(n6934), .ZN(n6485) );
  NAND2_X1 U7715 ( .A1(n4856), .A2(P1_REG3_REG_1__SCAN_IN), .ZN(n6484) );
  NAND4_X2 U7716 ( .A1(n6484), .A2(n6483), .A3(n6482), .A4(n6481), .ZN(n6896)
         );
  OAI22_X1 U7717 ( .A1(n8357), .A2(n6485), .B1(n6897), .B2(n9881), .ZN(n6982)
         );
  AOI21_X1 U7718 ( .B1(n6983), .B2(n6486), .A(n6982), .ZN(n6747) );
  INV_X1 U7719 ( .A(n8596), .ZN(n6628) );
  OR2_X1 U7720 ( .A1(n8553), .A2(n6628), .ZN(n6763) );
  NAND2_X1 U7721 ( .A1(n6763), .A2(n10047), .ZN(n6625) );
  NOR4_X1 U7722 ( .A1(P1_D_REG_23__SCAN_IN), .A2(P1_D_REG_22__SCAN_IN), .A3(
        P1_D_REG_21__SCAN_IN), .A4(P1_D_REG_20__SCAN_IN), .ZN(n6495) );
  NOR4_X1 U7723 ( .A1(P1_D_REG_27__SCAN_IN), .A2(P1_D_REG_26__SCAN_IN), .A3(
        P1_D_REG_25__SCAN_IN), .A4(P1_D_REG_24__SCAN_IN), .ZN(n6494) );
  OR4_X1 U7724 ( .A1(P1_D_REG_31__SCAN_IN), .A2(P1_D_REG_30__SCAN_IN), .A3(
        P1_D_REG_29__SCAN_IN), .A4(P1_D_REG_28__SCAN_IN), .ZN(n6492) );
  NOR4_X1 U7725 ( .A1(P1_D_REG_15__SCAN_IN), .A2(P1_D_REG_14__SCAN_IN), .A3(
        P1_D_REG_13__SCAN_IN), .A4(P1_D_REG_12__SCAN_IN), .ZN(n6490) );
  NOR4_X1 U7726 ( .A1(P1_D_REG_17__SCAN_IN), .A2(P1_D_REG_19__SCAN_IN), .A3(
        P1_D_REG_18__SCAN_IN), .A4(P1_D_REG_16__SCAN_IN), .ZN(n6489) );
  NOR4_X1 U7727 ( .A1(P1_D_REG_7__SCAN_IN), .A2(P1_D_REG_6__SCAN_IN), .A3(
        P1_D_REG_5__SCAN_IN), .A4(P1_D_REG_2__SCAN_IN), .ZN(n6488) );
  NOR4_X1 U7728 ( .A1(P1_D_REG_11__SCAN_IN), .A2(P1_D_REG_10__SCAN_IN), .A3(
        P1_D_REG_9__SCAN_IN), .A4(P1_D_REG_8__SCAN_IN), .ZN(n6487) );
  NAND4_X1 U7729 ( .A1(n6490), .A2(n6489), .A3(n6488), .A4(n6487), .ZN(n6491)
         );
  NOR4_X1 U7730 ( .A1(P1_D_REG_4__SCAN_IN), .A2(P1_D_REG_3__SCAN_IN), .A3(
        n6492), .A4(n6491), .ZN(n6493) );
  AND3_X1 U7731 ( .A1(n6495), .A2(n6494), .A3(n6493), .ZN(n6496) );
  OR2_X1 U7732 ( .A1(n10046), .A2(n6496), .ZN(n6621) );
  INV_X1 U7733 ( .A(n6621), .ZN(n6497) );
  OR2_X1 U7734 ( .A1(n8547), .A2(n8595), .ZN(n10582) );
  INV_X1 U7735 ( .A(n6920), .ZN(n6498) );
  OAI21_X1 U7736 ( .B1(n10582), .B2(n6623), .A(n6498), .ZN(n6499) );
  INV_X1 U7737 ( .A(n6743), .ZN(n6921) );
  NAND2_X1 U7738 ( .A1(n10633), .A2(P1_REG1_REG_0__SCAN_IN), .ZN(n6500) );
  OAI21_X1 U7739 ( .B1(n6747), .B2(n10633), .A(n6500), .ZN(P1_U3523) );
  INV_X1 U7740 ( .A(P1_ADDR_REG_5__SCAN_IN), .ZN(n6514) );
  AOI211_X1 U7741 ( .C1(n6503), .C2(n6502), .A(n10380), .B(n6501), .ZN(n6504)
         );
  AND2_X1 U7742 ( .A1(P1_U3084), .A2(P1_REG3_REG_5__SCAN_IN), .ZN(n7035) );
  NOR2_X1 U7743 ( .A1(n6504), .A2(n7035), .ZN(n6513) );
  INV_X1 U7744 ( .A(n6505), .ZN(n6508) );
  INV_X1 U7745 ( .A(n6506), .ZN(n6507) );
  NAND3_X1 U7746 ( .A1(n9639), .A2(n6508), .A3(n6507), .ZN(n6509) );
  AOI21_X1 U7747 ( .B1(n6510), .B2(n6509), .A(n9673), .ZN(n6511) );
  AOI21_X1 U7748 ( .B1(n9678), .B2(n7026), .A(n6511), .ZN(n6512) );
  OAI211_X1 U7749 ( .C1(n6514), .C2(n10391), .A(n6513), .B(n6512), .ZN(
        P1_U3246) );
  AOI21_X1 U7750 ( .B1(n6517), .B2(n6516), .A(n6515), .ZN(n6527) );
  OAI21_X1 U7751 ( .B1(n6520), .B2(n6519), .A(n6518), .ZN(n6525) );
  INV_X1 U7752 ( .A(P1_REG3_REG_8__SCAN_IN), .ZN(n6521) );
  NOR2_X1 U7753 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6521), .ZN(n7470) );
  AOI21_X1 U7754 ( .B1(n10386), .B2(P1_ADDR_REG_8__SCAN_IN), .A(n7470), .ZN(
        n6522) );
  OAI21_X1 U7755 ( .B1(n6523), .B2(n10393), .A(n6522), .ZN(n6524) );
  AOI21_X1 U7756 ( .B1(n6525), .B2(n10398), .A(n6524), .ZN(n6526) );
  OAI21_X1 U7757 ( .B1(n6527), .B2(n9673), .A(n6526), .ZN(P1_U3249) );
  INV_X1 U7758 ( .A(P1_REG3_REG_3__SCAN_IN), .ZN(n6941) );
  NOR2_X1 U7759 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n6941), .ZN(n6810) );
  AOI211_X1 U7760 ( .C1(n6530), .C2(n6529), .A(n6528), .B(n10380), .ZN(n6531)
         );
  AOI211_X1 U7761 ( .C1(n10386), .C2(P1_ADDR_REG_3__SCAN_IN), .A(n6810), .B(
        n6531), .ZN(n6538) );
  INV_X1 U7762 ( .A(n9673), .ZN(n10401) );
  INV_X1 U7763 ( .A(n6532), .ZN(n6536) );
  NAND3_X1 U7764 ( .A1(n6565), .A2(n6534), .A3(n6533), .ZN(n6535) );
  NAND3_X1 U7765 ( .A1(n10401), .A2(n6536), .A3(n6535), .ZN(n6537) );
  OAI211_X1 U7766 ( .C1(n10393), .C2(n6539), .A(n6538), .B(n6537), .ZN(
        P1_U3244) );
  INV_X1 U7767 ( .A(n7729), .ZN(n6542) );
  AOI22_X1 U7768 ( .A1(n7253), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_12__SCAN_IN), .B2(n9487), .ZN(n6540) );
  OAI21_X1 U7769 ( .B1(n6542), .B2(n4857), .A(n6540), .ZN(P2_U3346) );
  AOI22_X1 U7770 ( .A1(n7730), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_12__SCAN_IN), .B2(n7017), .ZN(n6541) );
  OAI21_X1 U7771 ( .B1(n6542), .B2(n10033), .A(n6541), .ZN(P1_U3341) );
  INV_X1 U7772 ( .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n6543) );
  NOR2_X1 U7773 ( .A1(n10391), .A2(n6543), .ZN(n6548) );
  NAND2_X1 U7774 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG1_REG_0__SCAN_IN), 
        .ZN(n6546) );
  AOI211_X1 U7775 ( .C1(n6546), .C2(n6545), .A(n6544), .B(n10380), .ZN(n6547)
         );
  AOI211_X1 U7776 ( .C1(P1_REG3_REG_1__SCAN_IN), .C2(P1_U3084), .A(n6548), .B(
        n6547), .ZN(n6554) );
  NAND2_X1 U7777 ( .A1(P1_IR_REG_0__SCAN_IN), .A2(P1_REG2_REG_0__SCAN_IN), 
        .ZN(n6591) );
  INV_X1 U7778 ( .A(n6591), .ZN(n6551) );
  INV_X1 U7779 ( .A(n6549), .ZN(n6550) );
  OAI211_X1 U7780 ( .C1(n6552), .C2(n6551), .A(n10401), .B(n6550), .ZN(n6553)
         );
  OAI211_X1 U7781 ( .C1(n10393), .C2(n6602), .A(n6554), .B(n6553), .ZN(
        P1_U3242) );
  INV_X1 U7782 ( .A(P1_REG3_REG_6__SCAN_IN), .ZN(n7036) );
  NOR2_X1 U7783 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7036), .ZN(n7139) );
  AOI211_X1 U7784 ( .C1(n6557), .C2(n6556), .A(n10380), .B(n6555), .ZN(n6558)
         );
  AOI211_X1 U7785 ( .C1(n10386), .C2(P1_ADDR_REG_6__SCAN_IN), .A(n7139), .B(
        n6558), .ZN(n6564) );
  AOI211_X1 U7786 ( .C1(n6561), .C2(n6560), .A(n9673), .B(n6559), .ZN(n6562)
         );
  AOI21_X1 U7787 ( .B1(n9678), .B2(n7129), .A(n6562), .ZN(n6563) );
  NAND2_X1 U7788 ( .A1(n6564), .A2(n6563), .ZN(P1_U3247) );
  INV_X1 U7789 ( .A(n6565), .ZN(n6566) );
  AOI211_X1 U7790 ( .C1(n6568), .C2(n6567), .A(n6566), .B(n9673), .ZN(n6576)
         );
  INV_X1 U7791 ( .A(P1_ADDR_REG_2__SCAN_IN), .ZN(n6574) );
  AOI211_X1 U7792 ( .C1(n6571), .C2(n6570), .A(n6569), .B(n10380), .ZN(n6572)
         );
  AOI21_X1 U7793 ( .B1(P1_REG3_REG_2__SCAN_IN), .B2(P1_U3084), .A(n6572), .ZN(
        n6573) );
  OAI21_X1 U7794 ( .B1(n6574), .B2(n10391), .A(n6573), .ZN(n6575) );
  AOI211_X1 U7795 ( .C1(n9678), .C2(n6577), .A(n6576), .B(n6575), .ZN(n6596)
         );
  NAND2_X1 U7796 ( .A1(n6607), .A2(n6628), .ZN(n6580) );
  INV_X1 U7797 ( .A(n6581), .ZN(n6582) );
  OR2_X1 U7798 ( .A1(n6581), .A2(n10383), .ZN(n6583) );
  NOR2_X1 U7799 ( .A1(n6587), .A2(n5477), .ZN(n6588) );
  NAND2_X1 U7800 ( .A1(n6589), .A2(n6588), .ZN(n6606) );
  NAND2_X1 U7801 ( .A1(n6590), .A2(n6606), .ZN(n6612) );
  OAI21_X1 U7802 ( .B1(n6590), .B2(n6606), .A(n6612), .ZN(n6827) );
  MUX2_X1 U7803 ( .A(n6591), .B(n6827), .S(n4860), .Z(n6595) );
  INV_X1 U7804 ( .A(P1_REG2_REG_0__SCAN_IN), .ZN(n10379) );
  AOI21_X1 U7805 ( .B1(n6592), .B2(n10379), .A(n6363), .ZN(n6593) );
  NOR2_X1 U7806 ( .A1(n6593), .A2(P1_IR_REG_0__SCAN_IN), .ZN(n10389) );
  INV_X1 U7807 ( .A(n10389), .ZN(n6594) );
  OAI211_X1 U7808 ( .C1(n6595), .C2(n6363), .A(P1_U4006), .B(n6594), .ZN(n9646) );
  NAND2_X1 U7809 ( .A1(n6596), .A2(n9646), .ZN(P1_U3243) );
  NAND2_X1 U7810 ( .A1(n6896), .A2(n6799), .ZN(n6605) );
  NAND2_X2 U7811 ( .A1(n6603), .A2(n6597), .ZN(n8136) );
  OR2_X1 U7812 ( .A1(n4858), .A2(n6599), .ZN(n6600) );
  NAND2_X1 U7813 ( .A1(n6995), .A2(n8678), .ZN(n6604) );
  NAND2_X1 U7814 ( .A1(n6605), .A2(n6604), .ZN(n6786) );
  INV_X1 U7815 ( .A(n6606), .ZN(n6610) );
  OR2_X1 U7816 ( .A1(n6607), .A2(n9772), .ZN(n6609) );
  NAND2_X4 U7817 ( .A1(n6609), .A2(n6608), .ZN(n8683) );
  NAND2_X1 U7818 ( .A1(n6610), .A2(n8683), .ZN(n6611) );
  NAND2_X1 U7819 ( .A1(n6612), .A2(n6611), .ZN(n6619) );
  INV_X1 U7820 ( .A(n6619), .ZN(n6617) );
  NAND2_X1 U7821 ( .A1(n6995), .A2(n6773), .ZN(n6614) );
  NAND2_X1 U7822 ( .A1(n6896), .A2(n6780), .ZN(n6613) );
  NAND2_X1 U7823 ( .A1(n6614), .A2(n6613), .ZN(n6615) );
  INV_X1 U7824 ( .A(n6618), .ZN(n6616) );
  NAND2_X1 U7825 ( .A1(n6617), .A2(n6616), .ZN(n6788) );
  NAND2_X1 U7826 ( .A1(n6619), .A2(n6618), .ZN(n6787) );
  NAND2_X1 U7827 ( .A1(n6788), .A2(n6787), .ZN(n6620) );
  XOR2_X1 U7828 ( .A(n6786), .B(n6620), .Z(n6638) );
  NAND3_X1 U7829 ( .A1(n6920), .A2(n6743), .A3(n6621), .ZN(n6626) );
  NOR2_X1 U7830 ( .A1(n6626), .A2(n8597), .ZN(n6629) );
  AND2_X1 U7831 ( .A1(n10618), .A2(n8553), .ZN(n6622) );
  NAND2_X1 U7832 ( .A1(n6629), .A2(n4942), .ZN(n6624) );
  NAND3_X1 U7833 ( .A1(n4942), .A2(n10047), .A3(n6626), .ZN(n6767) );
  INV_X1 U7834 ( .A(n6625), .ZN(n6627) );
  NAND2_X1 U7835 ( .A1(n6626), .A2(n10618), .ZN(n6764) );
  NAND3_X1 U7836 ( .A1(n6767), .A2(n6627), .A3(n6764), .ZN(n8300) );
  AOI22_X1 U7837 ( .A1(n6995), .A2(n9607), .B1(n8300), .B2(
        P1_REG3_REG_1__SCAN_IN), .ZN(n6637) );
  AND2_X1 U7838 ( .A1(n6629), .A2(n6628), .ZN(n6635) );
  INV_X1 U7839 ( .A(n6635), .ZN(n6630) );
  NAND2_X1 U7840 ( .A1(n4856), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n6633) );
  NAND2_X1 U7841 ( .A1(n6774), .A2(P1_REG1_REG_2__SCAN_IN), .ZN(n6631) );
  INV_X1 U7842 ( .A(n6797), .ZN(n9630) );
  AOI22_X1 U7843 ( .A1(n9601), .A2(n9630), .B1(n9566), .B2(n9631), .ZN(n6636)
         );
  OAI211_X1 U7844 ( .C1(n6638), .C2(n9609), .A(n6637), .B(n6636), .ZN(P1_U3220) );
  INV_X1 U7845 ( .A(n8935), .ZN(n6639) );
  AOI21_X1 U7846 ( .B1(n6640), .B2(P2_STATE_REG_SCAN_IN), .A(n6639), .ZN(n6641) );
  OAI21_X1 U7847 ( .B1(n10050), .B2(n6642), .A(n6641), .ZN(n6644) );
  NAND2_X1 U7848 ( .A1(n6644), .A2(n6643), .ZN(n6645) );
  NAND2_X1 U7849 ( .A1(n6645), .A2(n9069), .ZN(n6674) );
  NAND2_X1 U7850 ( .A1(n6674), .A2(n6188), .ZN(n10414) );
  NOR2_X1 U7851 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10127), .ZN(n6657) );
  INV_X1 U7852 ( .A(n6645), .ZN(n6647) );
  INV_X1 U7853 ( .A(P2_REG1_REG_4__SCAN_IN), .ZN(n10542) );
  MUX2_X1 U7854 ( .A(n10542), .B(P2_REG1_REG_4__SCAN_IN), .S(n6659), .Z(n6751)
         );
  INV_X1 U7855 ( .A(P2_REG1_REG_3__SCAN_IN), .ZN(n6648) );
  MUX2_X1 U7856 ( .A(P2_REG1_REG_3__SCAN_IN), .B(n6648), .S(n10448), .Z(n10451) );
  INV_X1 U7857 ( .A(P2_REG1_REG_2__SCAN_IN), .ZN(n10525) );
  MUX2_X1 U7858 ( .A(n10525), .B(P2_REG1_REG_2__SCAN_IN), .S(n10435), .Z(
        n10438) );
  NAND2_X1 U7859 ( .A1(n10421), .A2(P2_REG1_REG_1__SCAN_IN), .ZN(n6650) );
  INV_X1 U7860 ( .A(P2_REG1_REG_1__SCAN_IN), .ZN(n6649) );
  MUX2_X1 U7861 ( .A(P2_REG1_REG_1__SCAN_IN), .B(n6649), .S(n10421), .Z(n10429) );
  NAND3_X1 U7862 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG1_REG_0__SCAN_IN), 
        .A3(n10429), .ZN(n10428) );
  NAND2_X1 U7863 ( .A1(n6650), .A2(n10428), .ZN(n10439) );
  NAND2_X1 U7864 ( .A1(n10438), .A2(n10439), .ZN(n10437) );
  OAI21_X1 U7865 ( .B1(n10435), .B2(n10525), .A(n10437), .ZN(n10452) );
  NAND2_X1 U7866 ( .A1(n10451), .A2(n10452), .ZN(n10449) );
  INV_X1 U7867 ( .A(n10449), .ZN(n6651) );
  AOI21_X1 U7868 ( .B1(n10448), .B2(P2_REG1_REG_3__SCAN_IN), .A(n6651), .ZN(
        n6752) );
  NOR2_X1 U7869 ( .A1(n6751), .A2(n6752), .ZN(n6750) );
  AOI21_X1 U7870 ( .B1(n6659), .B2(P2_REG1_REG_4__SCAN_IN), .A(n6750), .ZN(
        n10465) );
  INV_X1 U7871 ( .A(P2_REG1_REG_5__SCAN_IN), .ZN(n10550) );
  MUX2_X1 U7872 ( .A(n10550), .B(P2_REG1_REG_5__SCAN_IN), .S(n10462), .Z(
        n10464) );
  NOR2_X1 U7873 ( .A1(n10465), .A2(n10464), .ZN(n10463) );
  AOI21_X1 U7874 ( .B1(n10462), .B2(P2_REG1_REG_5__SCAN_IN), .A(n10463), .ZN(
        n10484) );
  INV_X1 U7875 ( .A(P2_REG1_REG_6__SCAN_IN), .ZN(n10567) );
  MUX2_X1 U7876 ( .A(n10567), .B(P2_REG1_REG_6__SCAN_IN), .S(n10477), .Z(
        n10483) );
  NOR2_X1 U7877 ( .A1(n10484), .A2(n10483), .ZN(n10482) );
  NOR2_X1 U7878 ( .A1(n6668), .A2(n10567), .ZN(n6681) );
  INV_X1 U7879 ( .A(P2_REG1_REG_7__SCAN_IN), .ZN(n6652) );
  MUX2_X1 U7880 ( .A(P2_REG1_REG_7__SCAN_IN), .B(n6652), .S(n6670), .Z(n6680)
         );
  OAI21_X1 U7881 ( .B1(n10482), .B2(n6681), .A(n6680), .ZN(n6679) );
  NAND2_X1 U7882 ( .A1(n6670), .A2(P2_REG1_REG_7__SCAN_IN), .ZN(n6654) );
  INV_X1 U7883 ( .A(P2_REG1_REG_8__SCAN_IN), .ZN(n10592) );
  MUX2_X1 U7884 ( .A(n10592), .B(P2_REG1_REG_8__SCAN_IN), .S(n6707), .Z(n6653)
         );
  AOI21_X1 U7885 ( .B1(n6679), .B2(n6654), .A(n6653), .ZN(n6731) );
  AND3_X1 U7886 ( .A1(n6679), .A2(n6654), .A3(n6653), .ZN(n6655) );
  NOR3_X1 U7887 ( .A1(n10481), .A2(n6731), .A3(n6655), .ZN(n6656) );
  AOI211_X1 U7888 ( .C1(P2_ADDR_REG_8__SCAN_IN), .C2(n10486), .A(n6657), .B(
        n6656), .ZN(n6678) );
  INV_X1 U7889 ( .A(P2_REG2_REG_8__SCAN_IN), .ZN(n6658) );
  MUX2_X1 U7890 ( .A(P2_REG2_REG_8__SCAN_IN), .B(n6658), .S(n6707), .Z(n6676)
         );
  INV_X1 U7891 ( .A(P2_REG2_REG_7__SCAN_IN), .ZN(n6672) );
  INV_X1 U7892 ( .A(P2_REG2_REG_6__SCAN_IN), .ZN(n10474) );
  INV_X1 U7893 ( .A(P2_REG2_REG_5__SCAN_IN), .ZN(n7409) );
  MUX2_X1 U7894 ( .A(P2_REG2_REG_5__SCAN_IN), .B(n7409), .S(n10462), .Z(n10468) );
  INV_X1 U7895 ( .A(P2_REG2_REG_4__SCAN_IN), .ZN(n7307) );
  MUX2_X1 U7896 ( .A(n7307), .B(P2_REG2_REG_4__SCAN_IN), .S(n6659), .Z(n6756)
         );
  INV_X1 U7897 ( .A(P2_REG2_REG_3__SCAN_IN), .ZN(n6660) );
  MUX2_X1 U7898 ( .A(P2_REG2_REG_3__SCAN_IN), .B(n6660), .S(n10448), .Z(n10454) );
  INV_X1 U7899 ( .A(P2_REG2_REG_2__SCAN_IN), .ZN(n6664) );
  MUX2_X1 U7900 ( .A(n6664), .B(P2_REG2_REG_2__SCAN_IN), .S(n10435), .Z(n10441) );
  NAND2_X1 U7901 ( .A1(n10421), .A2(P2_REG2_REG_1__SCAN_IN), .ZN(n6663) );
  INV_X1 U7902 ( .A(P2_REG2_REG_1__SCAN_IN), .ZN(n6661) );
  MUX2_X1 U7903 ( .A(n6661), .B(P2_REG2_REG_1__SCAN_IN), .S(n10421), .Z(n6662)
         );
  INV_X1 U7904 ( .A(n6662), .ZN(n10424) );
  NAND3_X1 U7905 ( .A1(P2_IR_REG_0__SCAN_IN), .A2(P2_REG2_REG_0__SCAN_IN), 
        .A3(n10424), .ZN(n10423) );
  NAND2_X1 U7906 ( .A1(n6663), .A2(n10423), .ZN(n10442) );
  NAND2_X1 U7907 ( .A1(n10441), .A2(n10442), .ZN(n10440) );
  OAI21_X1 U7908 ( .B1(n10435), .B2(n6664), .A(n10440), .ZN(n10455) );
  NAND2_X1 U7909 ( .A1(n10454), .A2(n10455), .ZN(n10453) );
  INV_X1 U7910 ( .A(n10453), .ZN(n6665) );
  AOI21_X1 U7911 ( .B1(n10448), .B2(P2_REG2_REG_3__SCAN_IN), .A(n6665), .ZN(
        n6755) );
  OR2_X1 U7912 ( .A1(n6756), .A2(n6755), .ZN(n6758) );
  OAI21_X1 U7913 ( .B1(n7307), .B2(n6761), .A(n6758), .ZN(n10469) );
  NAND2_X1 U7914 ( .A1(n10468), .A2(n10469), .ZN(n10467) );
  OAI21_X1 U7915 ( .B1(n7409), .B2(n6666), .A(n10467), .ZN(n10476) );
  AOI21_X1 U7916 ( .B1(n10477), .B2(P2_REG2_REG_6__SCAN_IN), .A(n10476), .ZN(
        n6667) );
  AOI21_X1 U7917 ( .B1(n10474), .B2(n6668), .A(n6667), .ZN(n6687) );
  NAND2_X1 U7918 ( .A1(n6670), .A2(P2_REG2_REG_7__SCAN_IN), .ZN(n6669) );
  OAI21_X1 U7919 ( .B1(n6670), .B2(P2_REG2_REG_7__SCAN_IN), .A(n6669), .ZN(
        n6671) );
  INV_X1 U7920 ( .A(n6671), .ZN(n6688) );
  NAND2_X1 U7921 ( .A1(n6687), .A2(n6688), .ZN(n6686) );
  OAI21_X1 U7922 ( .B1(n6672), .B2(n6691), .A(n6686), .ZN(n6675) );
  INV_X1 U7923 ( .A(n6646), .ZN(n9112) );
  NAND3_X1 U7924 ( .A1(n6674), .A2(n9112), .A3(n6673), .ZN(n10415) );
  NAND2_X1 U7925 ( .A1(n6675), .A2(n6676), .ZN(n6718) );
  OAI211_X1 U7926 ( .C1(n6676), .C2(n6675), .A(n10480), .B(n6718), .ZN(n6677)
         );
  OAI211_X1 U7927 ( .C1(n10414), .C2(n6719), .A(n6678), .B(n6677), .ZN(
        P2_U3253) );
  INV_X1 U7928 ( .A(P2_REG3_REG_7__SCAN_IN), .ZN(n10114) );
  NOR2_X1 U7929 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10114), .ZN(n6685) );
  INV_X1 U7930 ( .A(n6679), .ZN(n6683) );
  NOR3_X1 U7931 ( .A1(n10482), .A2(n6681), .A3(n6680), .ZN(n6682) );
  NOR3_X1 U7932 ( .A1(n10481), .A2(n6683), .A3(n6682), .ZN(n6684) );
  AOI211_X1 U7933 ( .C1(P2_ADDR_REG_7__SCAN_IN), .C2(n10486), .A(n6685), .B(
        n6684), .ZN(n6690) );
  OAI211_X1 U7934 ( .C1(n6688), .C2(n6687), .A(n10480), .B(n6686), .ZN(n6689)
         );
  OAI211_X1 U7935 ( .C1(n10414), .C2(n6691), .A(n6690), .B(n6689), .ZN(
        P2_U3252) );
  NAND2_X1 U7936 ( .A1(n6849), .A2(P1_REG3_REG_6__SCAN_IN), .ZN(n7142) );
  NAND2_X1 U7937 ( .A1(n7188), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7464) );
  INV_X1 U7938 ( .A(P1_REG3_REG_11__SCAN_IN), .ZN(n7654) );
  NAND2_X1 U7939 ( .A1(n7664), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7740) );
  INV_X1 U7940 ( .A(P1_REG3_REG_13__SCAN_IN), .ZN(n7739) );
  INV_X1 U7941 ( .A(P1_REG3_REG_14__SCAN_IN), .ZN(n7861) );
  NAND2_X1 U7942 ( .A1(P1_REG3_REG_18__SCAN_IN), .A2(P1_REG3_REG_17__SCAN_IN), 
        .ZN(n6692) );
  INV_X1 U7943 ( .A(P1_REG3_REG_19__SCAN_IN), .ZN(n8156) );
  NAND2_X1 U7944 ( .A1(n8183), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8197) );
  INV_X1 U7945 ( .A(n8197), .ZN(n6693) );
  INV_X1 U7946 ( .A(n7069), .ZN(n8218) );
  INV_X1 U7947 ( .A(n6694), .ZN(n8199) );
  INV_X1 U7948 ( .A(P1_REG3_REG_23__SCAN_IN), .ZN(n6695) );
  NAND2_X1 U7949 ( .A1(n8199), .A2(n6695), .ZN(n6696) );
  AND2_X1 U7950 ( .A1(n8218), .A2(n6696), .ZN(n9786) );
  NAND2_X1 U7951 ( .A1(n4856), .A2(n9786), .ZN(n6702) );
  NAND2_X1 U7952 ( .A1(n6774), .A2(P1_REG1_REG_23__SCAN_IN), .ZN(n6701) );
  INV_X1 U7953 ( .A(P1_REG2_REG_23__SCAN_IN), .ZN(n6697) );
  OR2_X1 U7954 ( .A1(n8268), .A2(n6697), .ZN(n6700) );
  INV_X1 U7955 ( .A(P1_REG0_REG_23__SCAN_IN), .ZN(n6698) );
  OR2_X1 U7956 ( .A1(n8270), .A2(n6698), .ZN(n6699) );
  INV_X1 U7957 ( .A(n9766), .ZN(n9801) );
  NAND2_X1 U7958 ( .A1(n9801), .A2(P1_U4006), .ZN(n6703) );
  OAI21_X1 U7959 ( .B1(n9627), .B2(n7788), .A(n6703), .ZN(P1_U3578) );
  INV_X1 U7960 ( .A(n7851), .ZN(n6749) );
  AOI22_X1 U7961 ( .A1(n7852), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_13__SCAN_IN), .B2(n7017), .ZN(n6704) );
  OAI21_X1 U7962 ( .B1(n6749), .B2(n10033), .A(n6704), .ZN(P1_U3340) );
  INV_X1 U7963 ( .A(P2_DATAO_REG_14__SCAN_IN), .ZN(n6705) );
  OAI222_X1 U7964 ( .A1(n10043), .A2(n7857), .B1(n6706), .B2(P1_U3084), .C1(
        n6705), .C2(n10039), .ZN(P1_U3339) );
  INV_X1 U7965 ( .A(n6863), .ZN(n6867) );
  INV_X1 U7966 ( .A(P2_REG1_REG_9__SCAN_IN), .ZN(n10610) );
  INV_X1 U7967 ( .A(n6728), .ZN(n6741) );
  INV_X1 U7968 ( .A(n6731), .ZN(n6709) );
  NAND2_X1 U7969 ( .A1(n6707), .A2(P2_REG1_REG_8__SCAN_IN), .ZN(n6727) );
  MUX2_X1 U7970 ( .A(n10610), .B(P2_REG1_REG_9__SCAN_IN), .S(n6728), .Z(n6708)
         );
  AOI21_X1 U7971 ( .B1(n6709), .B2(n6727), .A(n6708), .ZN(n6733) );
  INV_X1 U7972 ( .A(n6733), .ZN(n6710) );
  OAI21_X1 U7973 ( .B1(n10610), .B2(n6741), .A(n6710), .ZN(n6713) );
  INV_X1 U7974 ( .A(P2_REG1_REG_10__SCAN_IN), .ZN(n6711) );
  MUX2_X1 U7975 ( .A(P2_REG1_REG_10__SCAN_IN), .B(n6711), .S(n6863), .Z(n6712)
         );
  NAND2_X1 U7976 ( .A1(n6712), .A2(n6713), .ZN(n6866) );
  OAI211_X1 U7977 ( .C1(n6713), .C2(n6712), .A(n6866), .B(n10450), .ZN(n6717)
         );
  NOR2_X1 U7978 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n6714), .ZN(n6715) );
  AOI21_X1 U7979 ( .B1(n10486), .B2(P2_ADDR_REG_10__SCAN_IN), .A(n6715), .ZN(
        n6716) );
  OAI211_X1 U7980 ( .C1(n10414), .C2(n6867), .A(n6717), .B(n6716), .ZN(n6726)
         );
  OAI21_X1 U7981 ( .B1(n6658), .B2(n6719), .A(n6718), .ZN(n6737) );
  INV_X1 U7982 ( .A(P2_REG2_REG_9__SCAN_IN), .ZN(n6720) );
  MUX2_X1 U7983 ( .A(P2_REG2_REG_9__SCAN_IN), .B(n6720), .S(n6728), .Z(n6738)
         );
  NAND2_X1 U7984 ( .A1(n6737), .A2(n6738), .ZN(n6736) );
  INV_X1 U7985 ( .A(n6736), .ZN(n6721) );
  AOI21_X1 U7986 ( .B1(n6728), .B2(P2_REG2_REG_9__SCAN_IN), .A(n6721), .ZN(
        n6724) );
  NAND2_X1 U7987 ( .A1(n6863), .A2(P2_REG2_REG_10__SCAN_IN), .ZN(n6722) );
  OAI21_X1 U7988 ( .B1(n6863), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6722), .ZN(
        n6723) );
  NOR2_X1 U7989 ( .A1(n6724), .A2(n6723), .ZN(n6862) );
  AOI211_X1 U7990 ( .C1(n6724), .C2(n6723), .A(n6862), .B(n10415), .ZN(n6725)
         );
  OR2_X1 U7991 ( .A1(n6726), .A2(n6725), .ZN(P2_U3255) );
  NAND2_X1 U7992 ( .A1(P2_REG3_REG_9__SCAN_IN), .A2(P2_U3152), .ZN(n9013) );
  INV_X1 U7993 ( .A(n9013), .ZN(n6735) );
  INV_X1 U7994 ( .A(n6727), .ZN(n6730) );
  MUX2_X1 U7995 ( .A(P2_REG1_REG_9__SCAN_IN), .B(n10610), .S(n6728), .Z(n6729)
         );
  NOR3_X1 U7996 ( .A1(n6731), .A2(n6730), .A3(n6729), .ZN(n6732) );
  NOR3_X1 U7997 ( .A1(n6733), .A2(n6732), .A3(n10481), .ZN(n6734) );
  AOI211_X1 U7998 ( .C1(P2_ADDR_REG_9__SCAN_IN), .C2(n10486), .A(n6735), .B(
        n6734), .ZN(n6740) );
  OAI211_X1 U7999 ( .C1(n6738), .C2(n6737), .A(n10480), .B(n6736), .ZN(n6739)
         );
  OAI211_X1 U8000 ( .C1(n10414), .C2(n6741), .A(n6740), .B(n6739), .ZN(
        P2_U3254) );
  INV_X1 U8001 ( .A(P1_DATAO_REG_14__SCAN_IN), .ZN(n6742) );
  OAI222_X1 U8002 ( .A1(P2_U3152), .A2(n7685), .B1(n4857), .B2(n7857), .C1(
        n6742), .C2(n9491), .ZN(P2_U3344) );
  INV_X1 U8003 ( .A(P1_REG0_REG_0__SCAN_IN), .ZN(n6745) );
  OR2_X1 U8004 ( .A1(n10637), .A2(n6745), .ZN(n6746) );
  OAI21_X1 U8005 ( .B1(n6747), .B2(n10635), .A(n6746), .ZN(P1_U3454) );
  INV_X1 U8006 ( .A(n7395), .ZN(n7390) );
  INV_X1 U8007 ( .A(P1_DATAO_REG_13__SCAN_IN), .ZN(n6748) );
  OAI222_X1 U8008 ( .A1(P2_U3152), .A2(n7390), .B1(n4857), .B2(n6749), .C1(
        n6748), .C2(n9491), .ZN(P2_U3345) );
  NAND2_X1 U8009 ( .A1(P2_REG3_REG_4__SCAN_IN), .A2(P2_U3152), .ZN(n7371) );
  INV_X1 U8010 ( .A(n7371), .ZN(n6754) );
  AOI211_X1 U8011 ( .C1(n6752), .C2(n6751), .A(n6750), .B(n10481), .ZN(n6753)
         );
  AOI211_X1 U8012 ( .C1(P2_ADDR_REG_4__SCAN_IN), .C2(n10486), .A(n6754), .B(
        n6753), .ZN(n6760) );
  NAND2_X1 U8013 ( .A1(n6756), .A2(n6755), .ZN(n6757) );
  NAND3_X1 U8014 ( .A1(n10480), .A2(n6758), .A3(n6757), .ZN(n6759) );
  OAI211_X1 U8015 ( .C1(n10414), .C2(n6761), .A(n6760), .B(n6759), .ZN(
        P2_U3249) );
  AND3_X1 U8016 ( .A1(n6763), .A2(n6581), .A3(n6762), .ZN(n6765) );
  NAND2_X1 U8017 ( .A1(n6765), .A2(n6764), .ZN(n6766) );
  NAND2_X1 U8018 ( .A1(n6766), .A2(P1_STATE_REG_SCAN_IN), .ZN(n6768) );
  NAND2_X1 U8019 ( .A1(n6768), .A2(n6767), .ZN(n9602) );
  INV_X1 U8020 ( .A(n9602), .ZN(n9593) );
  AOI22_X1 U8021 ( .A1(n8153), .A2(P2_DATAO_REG_3__SCAN_IN), .B1(n5192), .B2(
        n6769), .ZN(n6772) );
  NAND2_X1 U8022 ( .A1(n6770), .A2(n7439), .ZN(n6771) );
  NAND2_X1 U8023 ( .A1(n6925), .A2(n6773), .ZN(n6782) );
  NAND2_X1 U8024 ( .A1(n4856), .A2(n6941), .ZN(n6779) );
  NAND2_X1 U8025 ( .A1(n6774), .A2(P1_REG1_REG_3__SCAN_IN), .ZN(n6778) );
  NAND2_X1 U8026 ( .A1(n6775), .A2(P1_REG2_REG_3__SCAN_IN), .ZN(n6777) );
  NAND2_X1 U8027 ( .A1(n5475), .A2(P1_REG0_REG_3__SCAN_IN), .ZN(n6776) );
  NAND4_X1 U8028 ( .A1(n6779), .A2(n6778), .A3(n6777), .A4(n6776), .ZN(n9629)
         );
  NAND2_X1 U8029 ( .A1(n9629), .A2(n6780), .ZN(n6781) );
  NAND2_X1 U8030 ( .A1(n6782), .A2(n6781), .ZN(n6783) );
  XNOR2_X1 U8031 ( .A(n6783), .B(n8675), .ZN(n6837) );
  NAND2_X1 U8032 ( .A1(n9629), .A2(n6799), .ZN(n6785) );
  NAND2_X1 U8033 ( .A1(n6925), .A2(n8678), .ZN(n6784) );
  NAND2_X1 U8034 ( .A1(n6785), .A2(n6784), .ZN(n6835) );
  XNOR2_X1 U8035 ( .A(n6837), .B(n6835), .ZN(n6839) );
  NAND2_X1 U8036 ( .A1(n6787), .A2(n6786), .ZN(n6789) );
  NAND2_X1 U8037 ( .A1(n6789), .A2(n6788), .ZN(n8299) );
  OR2_X1 U8038 ( .A1(n8136), .A2(n6790), .ZN(n6796) );
  OR2_X1 U8039 ( .A1(n6792), .A2(n6791), .ZN(n6795) );
  NAND2_X1 U8040 ( .A1(n5192), .A2(n6577), .ZN(n6794) );
  XNOR2_X1 U8041 ( .A(n6798), .B(n8683), .ZN(n6801) );
  INV_X1 U8042 ( .A(n8301), .ZN(n10512) );
  OAI22_X1 U8043 ( .A1(n6797), .A2(n7033), .B1(n10512), .B2(n8685), .ZN(n6800)
         );
  XNOR2_X1 U8044 ( .A(n6801), .B(n6800), .ZN(n8298) );
  OR2_X1 U8045 ( .A1(n6801), .A2(n6800), .ZN(n6802) );
  XNOR2_X1 U8046 ( .A(n6839), .B(n6840), .ZN(n6803) );
  NAND2_X1 U8047 ( .A1(n6803), .A2(n9590), .ZN(n6812) );
  INV_X1 U8048 ( .A(P1_REG3_REG_4__SCAN_IN), .ZN(n6804) );
  XNOR2_X1 U8049 ( .A(n6804), .B(P1_REG3_REG_3__SCAN_IN), .ZN(n6834) );
  NAND2_X1 U8050 ( .A1(n4856), .A2(n6834), .ZN(n6808) );
  NAND2_X1 U8051 ( .A1(n6774), .A2(P1_REG1_REG_4__SCAN_IN), .ZN(n6807) );
  OR2_X1 U8052 ( .A1(n8268), .A2(n6335), .ZN(n6806) );
  NAND2_X1 U8053 ( .A1(n5475), .A2(P1_REG0_REG_4__SCAN_IN), .ZN(n6805) );
  OAI22_X1 U8054 ( .A1(n9605), .A2(n6797), .B1(n4989), .B2(n9569), .ZN(n6809)
         );
  AOI211_X1 U8055 ( .C1(n6925), .C2(n9607), .A(n6810), .B(n6809), .ZN(n6811)
         );
  OAI211_X1 U8056 ( .C1(P1_REG3_REG_3__SCAN_IN), .C2(n9593), .A(n6812), .B(
        n6811), .ZN(P1_U3216) );
  INV_X1 U8057 ( .A(P1_ADDR_REG_10__SCAN_IN), .ZN(n6814) );
  NOR2_X1 U8058 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7522), .ZN(n7720) );
  INV_X1 U8059 ( .A(n7720), .ZN(n6813) );
  OAI21_X1 U8060 ( .B1(n10391), .B2(n6814), .A(n6813), .ZN(n6820) );
  OAI211_X1 U8061 ( .C1(n6817), .C2(n6816), .A(n10401), .B(n6815), .ZN(n6818)
         );
  INV_X1 U8062 ( .A(n6818), .ZN(n6819) );
  AOI211_X1 U8063 ( .C1(n9678), .C2(n7645), .A(n6820), .B(n6819), .ZN(n6826)
         );
  OAI21_X1 U8064 ( .B1(n6823), .B2(n6822), .A(n6821), .ZN(n6824) );
  NAND2_X1 U8065 ( .A1(n6824), .A2(n10398), .ZN(n6825) );
  NAND2_X1 U8066 ( .A1(n6826), .A2(n6825), .ZN(P1_U3251) );
  INV_X1 U8067 ( .A(n6827), .ZN(n6832) );
  INV_X1 U8068 ( .A(n8300), .ZN(n6829) );
  INV_X1 U8069 ( .A(P1_REG3_REG_0__SCAN_IN), .ZN(n6828) );
  OAI22_X1 U8070 ( .A1(n9598), .A2(n6989), .B1(n6829), .B2(n6828), .ZN(n6830)
         );
  AOI21_X1 U8071 ( .B1(n9601), .B2(n6896), .A(n6830), .ZN(n6831) );
  OAI21_X1 U8072 ( .B1(n6832), .B2(n9609), .A(n6831), .ZN(P1_U3230) );
  NAND2_X1 U8073 ( .A1(P2_DATAO_REG_29__SCAN_IN), .A2(n9069), .ZN(n6833) );
  OAI21_X1 U8074 ( .B1(n8715), .B2(n9069), .A(n6833), .ZN(P2_U3581) );
  INV_X1 U8075 ( .A(n6834), .ZN(n6936) );
  INV_X1 U8076 ( .A(n6835), .ZN(n6836) );
  AND2_X1 U8077 ( .A1(n6837), .A2(n6836), .ZN(n6838) );
  OR2_X1 U8078 ( .A1(n6841), .A2(n6792), .ZN(n6843) );
  AOI22_X1 U8079 ( .A1(n8153), .A2(P2_DATAO_REG_4__SCAN_IN), .B1(n5192), .B2(
        n9643), .ZN(n6842) );
  NAND2_X1 U8080 ( .A1(n6843), .A2(n6842), .ZN(n10528) );
  NAND2_X1 U8081 ( .A1(n10528), .A2(n6773), .ZN(n6845) );
  NAND2_X1 U8082 ( .A1(n9628), .A2(n8678), .ZN(n6844) );
  NAND2_X1 U8083 ( .A1(n6845), .A2(n6844), .ZN(n6846) );
  XNOR2_X1 U8084 ( .A(n6846), .B(n8683), .ZN(n7020) );
  AOI22_X1 U8085 ( .A1(n10528), .A2(n8678), .B1(n6799), .B2(n9628), .ZN(n7021)
         );
  XNOR2_X1 U8086 ( .A(n7020), .B(n7021), .ZN(n6847) );
  OAI211_X1 U8087 ( .C1(n6848), .C2(n6847), .A(n7024), .B(n9590), .ZN(n6859)
         );
  AND2_X1 U8088 ( .A1(P1_U3084), .A2(P1_REG3_REG_4__SCAN_IN), .ZN(n9636) );
  INV_X1 U8089 ( .A(n9629), .ZN(n6926) );
  INV_X1 U8090 ( .A(n6849), .ZN(n7037) );
  INV_X1 U8091 ( .A(P1_REG3_REG_5__SCAN_IN), .ZN(n6851) );
  NAND2_X1 U8092 ( .A1(P1_REG3_REG_3__SCAN_IN), .A2(P1_REG3_REG_4__SCAN_IN), 
        .ZN(n6850) );
  NAND2_X1 U8093 ( .A1(n6851), .A2(n6850), .ZN(n6852) );
  AND2_X1 U8094 ( .A1(n7037), .A2(n6852), .ZN(n7118) );
  NAND2_X1 U8095 ( .A1(n4856), .A2(n7118), .ZN(n6856) );
  NAND2_X1 U8096 ( .A1(n6774), .A2(P1_REG1_REG_5__SCAN_IN), .ZN(n6855) );
  NAND2_X1 U8097 ( .A1(n5475), .A2(P1_REG0_REG_5__SCAN_IN), .ZN(n6854) );
  OR2_X1 U8098 ( .A1(n8268), .A2(n7120), .ZN(n6853) );
  NAND4_X1 U8099 ( .A1(n6856), .A2(n6855), .A3(n6854), .A4(n6853), .ZN(n9626)
         );
  INV_X1 U8100 ( .A(n9626), .ZN(n7169) );
  OAI22_X1 U8101 ( .A1(n9605), .A2(n6926), .B1(n7169), .B2(n9569), .ZN(n6857)
         );
  AOI211_X1 U8102 ( .C1(n10528), .C2(n9607), .A(n9636), .B(n6857), .ZN(n6858)
         );
  OAI211_X1 U8103 ( .C1(n9593), .C2(n6936), .A(n6859), .B(n6858), .ZN(P1_U3228) );
  INV_X1 U8104 ( .A(P2_REG2_REG_11__SCAN_IN), .ZN(n6860) );
  MUX2_X1 U8105 ( .A(n6860), .B(P2_REG2_REG_11__SCAN_IN), .S(n6868), .Z(n6861)
         );
  INV_X1 U8106 ( .A(n6861), .ZN(n6865) );
  AOI21_X1 U8107 ( .B1(n6863), .B2(P2_REG2_REG_10__SCAN_IN), .A(n6862), .ZN(
        n6864) );
  NAND2_X1 U8108 ( .A1(n6864), .A2(n6865), .ZN(n7008) );
  OAI21_X1 U8109 ( .B1(n6865), .B2(n6864), .A(n7008), .ZN(n6876) );
  INV_X1 U8110 ( .A(n6868), .ZN(n7010) );
  OAI21_X1 U8111 ( .B1(n6867), .B2(n6711), .A(n6866), .ZN(n6871) );
  INV_X1 U8112 ( .A(P2_REG1_REG_11__SCAN_IN), .ZN(n6869) );
  MUX2_X1 U8113 ( .A(P2_REG1_REG_11__SCAN_IN), .B(n6869), .S(n6868), .Z(n6870)
         );
  NAND2_X1 U8114 ( .A1(n6870), .A2(n6871), .ZN(n6999) );
  OAI211_X1 U8115 ( .C1(n6871), .C2(n6870), .A(n10450), .B(n6999), .ZN(n6874)
         );
  AND2_X1 U8116 ( .A1(P2_U3152), .A2(P2_REG3_REG_11__SCAN_IN), .ZN(n6872) );
  AOI21_X1 U8117 ( .B1(n10486), .B2(P2_ADDR_REG_11__SCAN_IN), .A(n6872), .ZN(
        n6873) );
  OAI211_X1 U8118 ( .C1(n10414), .C2(n7010), .A(n6874), .B(n6873), .ZN(n6875)
         );
  AOI21_X1 U8119 ( .B1(n10480), .B2(n6876), .A(n6875), .ZN(n6877) );
  INV_X1 U8120 ( .A(n6877), .ZN(P2_U3256) );
  AOI21_X1 U8121 ( .B1(n7651), .B2(P1_REG1_REG_11__SCAN_IN), .A(n6878), .ZN(
        n6880) );
  XOR2_X1 U8122 ( .A(n6880), .B(n6879), .Z(n6891) );
  INV_X1 U8123 ( .A(n6881), .ZN(n6883) );
  INV_X1 U8124 ( .A(P1_REG2_REG_11__SCAN_IN), .ZN(n7657) );
  NAND3_X1 U8125 ( .A1(n6883), .A2(n6882), .A3(n7657), .ZN(n6884) );
  NAND3_X1 U8126 ( .A1(n7103), .A2(n10401), .A3(n6884), .ZN(n6890) );
  OAI21_X1 U8127 ( .B1(n6885), .B2(n10374), .A(n10393), .ZN(n6888) );
  AND2_X1 U8128 ( .A1(P1_U3084), .A2(P1_REG3_REG_11__SCAN_IN), .ZN(n7765) );
  INV_X1 U8129 ( .A(P1_ADDR_REG_11__SCAN_IN), .ZN(n6886) );
  NOR2_X1 U8130 ( .A1(n10391), .A2(n6886), .ZN(n6887) );
  AOI211_X1 U8131 ( .C1(n7651), .C2(n6888), .A(n7765), .B(n6887), .ZN(n6889)
         );
  OAI211_X1 U8132 ( .C1(n6891), .C2(n10380), .A(n6890), .B(n6889), .ZN(
        P1_U3252) );
  INV_X1 U8133 ( .A(n8006), .ZN(n6895) );
  OAI222_X1 U8134 ( .A1(n10039), .A2(n6893), .B1(n10033), .B2(n6895), .C1(
        P1_U3084), .C2(n6892), .ZN(P1_U3338) );
  INV_X1 U8135 ( .A(n7810), .ZN(n7820) );
  OAI222_X1 U8136 ( .A1(n7820), .A2(P2_U3152), .B1(n4857), .B2(n6895), .C1(
        n6894), .C2(n9491), .ZN(P2_U3343) );
  INV_X1 U8137 ( .A(P1_REG0_REG_3__SCAN_IN), .ZN(n6913) );
  XNOR2_X1 U8138 ( .A(n6995), .B(n6897), .ZN(n6988) );
  NAND2_X1 U8139 ( .A1(n6896), .A2(n6995), .ZN(n6898) );
  NAND2_X1 U8140 ( .A1(n6797), .A2(n10512), .ZN(n6899) );
  NAND2_X1 U8141 ( .A1(n7053), .A2(n6899), .ZN(n6900) );
  INV_X1 U8142 ( .A(n8358), .ZN(n6903) );
  NAND2_X1 U8143 ( .A1(n6900), .A2(n6903), .ZN(n6918) );
  OAI21_X1 U8144 ( .B1(n6900), .B2(n6903), .A(n6918), .ZN(n6910) );
  INV_X1 U8145 ( .A(n6910), .ZN(n6946) );
  AOI21_X1 U8146 ( .B1(n6607), .B2(n6608), .A(n9772), .ZN(n6901) );
  OAI22_X1 U8147 ( .A1(n4989), .A2(n9881), .B1(n6797), .B2(n9879), .ZN(n6909)
         );
  NAND2_X1 U8148 ( .A1(n6897), .A2(n6995), .ZN(n6902) );
  NAND3_X1 U8149 ( .A1(n7059), .A2(n6903), .A3(n8560), .ZN(n6907) );
  OR2_X1 U8150 ( .A1(n6607), .A2(n6904), .ZN(n6906) );
  OR2_X1 U8151 ( .A1(n4855), .A2(n6579), .ZN(n6905) );
  AOI21_X1 U8152 ( .B1(n6927), .B2(n6907), .A(n10626), .ZN(n6908) );
  AOI211_X1 U8153 ( .C1(n10629), .C2(n6910), .A(n6909), .B(n6908), .ZN(n6940)
         );
  AOI21_X1 U8154 ( .B1(n6925), .B2(n7056), .A(n6932), .ZN(n6943) );
  AOI22_X1 U8155 ( .A1(n6943), .A2(n10617), .B1(n10578), .B2(n6925), .ZN(n6911) );
  OAI211_X1 U8156 ( .C1(n6946), .C2(n10582), .A(n6940), .B(n6911), .ZN(n6914)
         );
  NAND2_X1 U8157 ( .A1(n6914), .A2(n10637), .ZN(n6912) );
  OAI21_X1 U8158 ( .B1(n10637), .B2(n6913), .A(n6912), .ZN(P1_U3463) );
  INV_X1 U8159 ( .A(P1_REG1_REG_3__SCAN_IN), .ZN(n6916) );
  NAND2_X1 U8160 ( .A1(n6914), .A2(n10634), .ZN(n6915) );
  OAI21_X1 U8161 ( .B1(n10634), .B2(n6916), .A(n6915), .ZN(P1_U3526) );
  INV_X1 U8162 ( .A(n6925), .ZN(n8568) );
  NAND2_X1 U8163 ( .A1(n6926), .A2(n8568), .ZN(n6917) );
  OAI21_X1 U8164 ( .B1(n6919), .B2(n8363), .A(n7110), .ZN(n6931) );
  INV_X1 U8165 ( .A(n6931), .ZN(n10532) );
  NAND2_X1 U8166 ( .A1(n6921), .A2(n6920), .ZN(n6922) );
  AND2_X2 U8167 ( .A1(n7208), .A2(n9866), .ZN(n9896) );
  INV_X2 U8168 ( .A(n9896), .ZN(n9841) );
  NOR2_X1 U8169 ( .A1(n6608), .A2(n6904), .ZN(n6924) );
  NAND2_X1 U8170 ( .A1(n9841), .A2(n6924), .ZN(n9899) );
  OAI22_X1 U8171 ( .A1(n6926), .A2(n9879), .B1(n7169), .B2(n9881), .ZN(n6930)
         );
  NAND2_X1 U8172 ( .A1(n6926), .A2(n6925), .ZN(n8565) );
  NAND3_X1 U8173 ( .A1(n6927), .A2(n8363), .A3(n8565), .ZN(n6928) );
  AOI21_X1 U8174 ( .B1(n7114), .B2(n6928), .A(n10626), .ZN(n6929) );
  AOI211_X1 U8175 ( .C1(n6931), .C2(n10629), .A(n6930), .B(n6929), .ZN(n10531)
         );
  MUX2_X1 U8176 ( .A(n6335), .B(n10531), .S(n9841), .Z(n6939) );
  INV_X1 U8177 ( .A(n6932), .ZN(n6933) );
  INV_X1 U8178 ( .A(n10528), .ZN(n8569) );
  AOI21_X1 U8179 ( .B1(n10528), .B2(n6933), .A(n7112), .ZN(n10529) );
  OR2_X1 U8180 ( .A1(n6934), .A2(n8596), .ZN(n6935) );
  NOR2_X2 U8181 ( .A1(n9896), .A2(n6935), .ZN(n9902) );
  OAI22_X1 U8182 ( .A1(n9898), .A2(n8569), .B1(n6936), .B2(n9866), .ZN(n6937)
         );
  AOI21_X1 U8183 ( .B1(n10529), .B2(n9902), .A(n6937), .ZN(n6938) );
  OAI211_X1 U8184 ( .C1(n10532), .C2(n9899), .A(n6939), .B(n6938), .ZN(
        P1_U3287) );
  MUX2_X1 U8185 ( .A(n6330), .B(n6940), .S(n9841), .Z(n6945) );
  OAI22_X1 U8186 ( .A1(n9898), .A2(n8568), .B1(P1_REG3_REG_3__SCAN_IN), .B2(
        n9866), .ZN(n6942) );
  AOI21_X1 U8187 ( .B1(n9902), .B2(n6943), .A(n6942), .ZN(n6944) );
  OAI211_X1 U8188 ( .C1(n6946), .C2(n9899), .A(n6945), .B(n6944), .ZN(P1_U3288) );
  NAND3_X1 U8189 ( .A1(n6949), .A2(n6948), .A3(n6947), .ZN(n6950) );
  INV_X1 U8190 ( .A(P2_REG1_REG_0__SCAN_IN), .ZN(n10426) );
  INV_X1 U8191 ( .A(n7319), .ZN(n7321) );
  NAND2_X1 U8192 ( .A1(n6952), .A2(n7317), .ZN(n8752) );
  INV_X1 U8193 ( .A(n8752), .ZN(n8899) );
  NOR2_X1 U8194 ( .A1(n7321), .A2(n8899), .ZN(n7316) );
  OAI22_X1 U8195 ( .A1(n7316), .A2(n9376), .B1(n5424), .B2(n9370), .ZN(n7311)
         );
  NAND2_X1 U8196 ( .A1(n9369), .A2(n6971), .ZN(n10697) );
  OAI22_X1 U8197 ( .A1(n7316), .A2(n10673), .B1(n7317), .B2(n6953), .ZN(n6954)
         );
  OR2_X1 U8198 ( .A1(n7311), .A2(n6954), .ZN(n6959) );
  NAND2_X1 U8199 ( .A1(n10701), .A2(n6959), .ZN(n6955) );
  OAI21_X1 U8200 ( .B1(n10701), .B2(n10426), .A(n6955), .ZN(P2_U3520) );
  INV_X1 U8201 ( .A(n6956), .ZN(n6957) );
  INV_X2 U8202 ( .A(n10702), .ZN(n10613) );
  INV_X1 U8203 ( .A(P2_REG0_REG_0__SCAN_IN), .ZN(n6961) );
  NAND2_X1 U8204 ( .A1(n10613), .A2(n6959), .ZN(n6960) );
  OAI21_X1 U8205 ( .B1(n10613), .B2(n6961), .A(n6960), .ZN(P2_U3451) );
  OAI21_X1 U8206 ( .B1(n6964), .B2(n6963), .A(n6962), .ZN(n6970) );
  OAI22_X1 U8207 ( .A1(n5071), .A2(n9371), .B1(n7217), .B2(n9370), .ZN(n6969)
         );
  OAI21_X1 U8208 ( .B1(n6966), .B2(n8900), .A(n6965), .ZN(n7349) );
  INV_X1 U8209 ( .A(n7349), .ZN(n6967) );
  NOR2_X1 U8210 ( .A1(n6967), .A2(n9369), .ZN(n6968) );
  AOI211_X1 U8211 ( .C1(n9349), .C2(n6970), .A(n6969), .B(n6968), .ZN(n7343)
         );
  INV_X1 U8212 ( .A(n6971), .ZN(n10655) );
  INV_X1 U8213 ( .A(n7298), .ZN(n6973) );
  NAND2_X1 U8214 ( .A1(n10519), .A2(n7348), .ZN(n6972) );
  NAND2_X1 U8215 ( .A1(n6973), .A2(n6972), .ZN(n7344) );
  OAI22_X1 U8216 ( .A1(n7344), .A2(n10693), .B1(n6974), .B2(n10691), .ZN(n6975) );
  AOI21_X1 U8217 ( .B1(n7349), .B2(n10655), .A(n6975), .ZN(n6976) );
  NAND2_X1 U8218 ( .A1(n7343), .A2(n6976), .ZN(n6978) );
  NAND2_X1 U8219 ( .A1(n6978), .A2(n10701), .ZN(n6977) );
  OAI21_X1 U8220 ( .B1(n10701), .B2(n6648), .A(n6977), .ZN(P2_U3523) );
  INV_X1 U8221 ( .A(P2_REG0_REG_3__SCAN_IN), .ZN(n6980) );
  NAND2_X1 U8222 ( .A1(n6978), .A2(n10613), .ZN(n6979) );
  OAI21_X1 U8223 ( .B1(n10613), .B2(n6980), .A(n6979), .ZN(P2_U3460) );
  NOR2_X1 U8224 ( .A1(n9866), .A2(n6828), .ZN(n6981) );
  OAI21_X1 U8225 ( .B1(n6982), .B2(n6981), .A(n9841), .ZN(n6985) );
  OAI21_X1 U8226 ( .B1(n10640), .B2(n9902), .A(n6983), .ZN(n6984) );
  OAI211_X1 U8227 ( .C1(n10379), .C2(n9841), .A(n6985), .B(n6984), .ZN(
        P1_U3291) );
  OAI21_X1 U8228 ( .B1(n6988), .B2(n6987), .A(n6986), .ZN(n6998) );
  OAI211_X1 U8229 ( .C1(n10491), .C2(n6989), .A(n10617), .B(n7054), .ZN(n10495) );
  OAI21_X1 U8230 ( .B1(n6991), .B2(n8360), .A(n6990), .ZN(n6992) );
  INV_X1 U8231 ( .A(n6998), .ZN(n10494) );
  AOI222_X1 U8232 ( .A1(n6992), .A2(n9891), .B1(n10629), .B2(n10494), .C1(
        n9631), .C2(n10622), .ZN(n10498) );
  INV_X1 U8233 ( .A(n9866), .ZN(n10638) );
  NOR2_X1 U8234 ( .A1(n6797), .A2(n9881), .ZN(n10493) );
  AOI21_X1 U8235 ( .B1(n10638), .B2(P1_REG3_REG_1__SCAN_IN), .A(n10493), .ZN(
        n6993) );
  OAI211_X1 U8236 ( .C1(n9772), .C2(n10495), .A(n10498), .B(n6993), .ZN(n6994)
         );
  NAND2_X1 U8237 ( .A1(n6994), .A2(n9841), .ZN(n6997) );
  AOI22_X1 U8238 ( .A1(n10640), .A2(n6995), .B1(P1_REG2_REG_1__SCAN_IN), .B2(
        n9896), .ZN(n6996) );
  OAI211_X1 U8239 ( .C1(n6998), .C2(n9899), .A(n6997), .B(n6996), .ZN(P1_U3290) );
  INV_X1 U8240 ( .A(n7253), .ZN(n7259) );
  NAND2_X1 U8241 ( .A1(P2_REG3_REG_12__SCAN_IN), .A2(P2_U3152), .ZN(n7635) );
  INV_X1 U8242 ( .A(n7635), .ZN(n7006) );
  OAI21_X1 U8243 ( .B1(n7010), .B2(n6869), .A(n6999), .ZN(n7003) );
  INV_X1 U8244 ( .A(n7003), .ZN(n7001) );
  INV_X1 U8245 ( .A(P2_REG1_REG_12__SCAN_IN), .ZN(n10670) );
  MUX2_X1 U8246 ( .A(P2_REG1_REG_12__SCAN_IN), .B(n10670), .S(n7253), .Z(n7000) );
  NAND2_X1 U8247 ( .A1(n7001), .A2(n7000), .ZN(n7257) );
  MUX2_X1 U8248 ( .A(n10670), .B(P2_REG1_REG_12__SCAN_IN), .S(n7253), .Z(n7002) );
  NAND2_X1 U8249 ( .A1(n7003), .A2(n7002), .ZN(n7004) );
  AOI21_X1 U8250 ( .B1(n7257), .B2(n7004), .A(n10481), .ZN(n7005) );
  AOI211_X1 U8251 ( .C1(P2_ADDR_REG_12__SCAN_IN), .C2(n10486), .A(n7006), .B(
        n7005), .ZN(n7014) );
  INV_X1 U8252 ( .A(P2_REG2_REG_12__SCAN_IN), .ZN(n7007) );
  MUX2_X1 U8253 ( .A(P2_REG2_REG_12__SCAN_IN), .B(n7007), .S(n7253), .Z(n7012)
         );
  INV_X1 U8254 ( .A(n7008), .ZN(n7009) );
  AOI21_X1 U8255 ( .B1(n7010), .B2(n6860), .A(n7009), .ZN(n7011) );
  NAND2_X1 U8256 ( .A1(n7011), .A2(n7012), .ZN(n7251) );
  OAI211_X1 U8257 ( .C1(n7012), .C2(n7011), .A(n10480), .B(n7251), .ZN(n7013)
         );
  OAI211_X1 U8258 ( .C1(n10414), .C2(n7259), .A(n7014), .B(n7013), .ZN(
        P2_U3257) );
  INV_X1 U8259 ( .A(P2_DATAO_REG_28__SCAN_IN), .ZN(n7016) );
  INV_X1 U8260 ( .A(n9146), .ZN(n9185) );
  NAND2_X1 U8261 ( .A1(n9185), .A2(P2_U3966), .ZN(n7015) );
  OAI21_X1 U8262 ( .B1(n7016), .B2(P2_U3966), .A(n7015), .ZN(P2_U3580) );
  INV_X1 U8263 ( .A(n8042), .ZN(n7081) );
  AOI22_X1 U8264 ( .A1(n9655), .A2(P1_STATE_REG_SCAN_IN), .B1(
        P2_DATAO_REG_16__SCAN_IN), .B2(n7017), .ZN(n7018) );
  OAI21_X1 U8265 ( .B1(n7081), .B2(n10033), .A(n7018), .ZN(P1_U3337) );
  INV_X1 U8266 ( .A(P2_DATAO_REG_17__SCAN_IN), .ZN(n8137) );
  OAI222_X1 U8267 ( .A1(n10043), .A2(n8135), .B1(n9670), .B2(P1_U3084), .C1(
        n8137), .C2(n10039), .ZN(P1_U3336) );
  INV_X1 U8268 ( .A(P1_DATAO_REG_17__SCAN_IN), .ZN(n7019) );
  OAI222_X1 U8269 ( .A1(P2_U3152), .A2(n9081), .B1(n4857), .B2(n8135), .C1(
        n7019), .C2(n9491), .ZN(P2_U3341) );
  OR2_X1 U8270 ( .A1(n7025), .A2(n6792), .ZN(n7028) );
  AOI22_X1 U8271 ( .A1(n8153), .A2(P2_DATAO_REG_5__SCAN_IN), .B1(n5192), .B2(
        n7026), .ZN(n7027) );
  OAI22_X1 U8272 ( .A1(n7111), .A2(n8686), .B1(n7169), .B2(n8685), .ZN(n7029)
         );
  XNOR2_X1 U8273 ( .A(n7029), .B(n8683), .ZN(n7031) );
  INV_X1 U8274 ( .A(n7031), .ZN(n7030) );
  NAND2_X1 U8275 ( .A1(n7125), .A2(n7126), .ZN(n7034) );
  OAI22_X1 U8276 ( .A1(n7111), .A2(n8685), .B1(n7169), .B2(n8682), .ZN(n7124)
         );
  XNOR2_X1 U8277 ( .A(n7034), .B(n7124), .ZN(n7049) );
  AOI21_X1 U8278 ( .B1(n9566), .B2(n9628), .A(n7035), .ZN(n7047) );
  NAND2_X1 U8279 ( .A1(n7231), .A2(n9607), .ZN(n7046) );
  NAND2_X1 U8280 ( .A1(n9602), .A2(n7118), .ZN(n7045) );
  NAND2_X1 U8281 ( .A1(n6774), .A2(P1_REG1_REG_6__SCAN_IN), .ZN(n7043) );
  NAND2_X1 U8282 ( .A1(n7037), .A2(n7036), .ZN(n7038) );
  AND2_X1 U8283 ( .A1(n7142), .A2(n7038), .ZN(n7180) );
  NAND2_X1 U8284 ( .A1(n4856), .A2(n7180), .ZN(n7042) );
  INV_X1 U8285 ( .A(P1_REG0_REG_6__SCAN_IN), .ZN(n7039) );
  OR2_X1 U8286 ( .A1(n8270), .A2(n7039), .ZN(n7041) );
  OR2_X1 U8287 ( .A1(n8268), .A2(n7178), .ZN(n7040) );
  NAND2_X1 U8288 ( .A1(n9601), .A2(n9625), .ZN(n7044) );
  NAND4_X1 U8289 ( .A1(n7047), .A2(n7046), .A3(n7045), .A4(n7044), .ZN(n7048)
         );
  AOI21_X1 U8290 ( .B1(n7049), .B2(n9590), .A(n7048), .ZN(n7050) );
  INV_X1 U8291 ( .A(n7050), .ZN(P1_U3225) );
  INV_X1 U8292 ( .A(n9899), .ZN(n10645) );
  NAND2_X1 U8293 ( .A1(n7051), .A2(n8359), .ZN(n7052) );
  NAND2_X1 U8294 ( .A1(n7053), .A2(n7052), .ZN(n10515) );
  NAND2_X1 U8295 ( .A1(n7054), .A2(n8301), .ZN(n7055) );
  AND2_X1 U8296 ( .A1(n7056), .A2(n7055), .ZN(n10510) );
  NAND2_X1 U8297 ( .A1(n9902), .A2(n10510), .ZN(n7058) );
  NAND2_X1 U8298 ( .A1(n10638), .A2(P1_REG3_REG_2__SCAN_IN), .ZN(n7057) );
  OAI211_X1 U8299 ( .C1(n9898), .C2(n10512), .A(n7058), .B(n7057), .ZN(n7067)
         );
  NAND2_X1 U8300 ( .A1(n10515), .A2(n10629), .ZN(n7065) );
  OAI21_X1 U8301 ( .B1(n8359), .B2(n8561), .A(n7059), .ZN(n7063) );
  NAND2_X1 U8302 ( .A1(n6896), .A2(n10622), .ZN(n7061) );
  NAND2_X1 U8303 ( .A1(n9629), .A2(n10623), .ZN(n7060) );
  NAND2_X1 U8304 ( .A1(n7061), .A2(n7060), .ZN(n7062) );
  AOI21_X1 U8305 ( .B1(n7063), .B2(n9891), .A(n7062), .ZN(n7064) );
  NAND2_X1 U8306 ( .A1(n7065), .A2(n7064), .ZN(n10513) );
  MUX2_X1 U8307 ( .A(n10513), .B(P1_REG2_REG_2__SCAN_IN), .S(n9896), .Z(n7066)
         );
  AOI211_X1 U8308 ( .C1(n10645), .C2(n10515), .A(n7067), .B(n7066), .ZN(n7068)
         );
  INV_X1 U8309 ( .A(n7068), .ZN(P1_U3289) );
  INV_X1 U8310 ( .A(n8331), .ZN(n7073) );
  INV_X1 U8311 ( .A(n7070), .ZN(n8266) );
  INV_X1 U8312 ( .A(P1_REG3_REG_28__SCAN_IN), .ZN(n7071) );
  NAND2_X1 U8313 ( .A1(n8266), .A2(n7071), .ZN(n7072) );
  NAND2_X1 U8314 ( .A1(n4856), .A2(n8691), .ZN(n7079) );
  NAND2_X1 U8315 ( .A1(n6774), .A2(P1_REG1_REG_28__SCAN_IN), .ZN(n7078) );
  INV_X1 U8316 ( .A(P1_REG2_REG_28__SCAN_IN), .ZN(n7074) );
  OR2_X1 U8317 ( .A1(n8268), .A2(n7074), .ZN(n7077) );
  INV_X1 U8318 ( .A(P1_REG0_REG_28__SCAN_IN), .ZN(n7075) );
  OR2_X1 U8319 ( .A1(n8270), .A2(n7075), .ZN(n7076) );
  INV_X1 U8320 ( .A(n9721), .ZN(n8342) );
  NAND2_X1 U8321 ( .A1(n8342), .A2(n9627), .ZN(n7080) );
  OAI21_X1 U8322 ( .B1(P1_U4006), .B2(n8605), .A(n7080), .ZN(P1_U3583) );
  INV_X1 U8323 ( .A(P1_DATAO_REG_16__SCAN_IN), .ZN(n7082) );
  OAI222_X1 U8324 ( .A1(n9491), .A2(n7082), .B1(n4857), .B2(n7081), .C1(
        P2_U3152), .C2(n7827), .ZN(P2_U3342) );
  NAND2_X1 U8325 ( .A1(n9049), .A2(n9241), .ZN(n9015) );
  NOR2_X1 U8326 ( .A1(n10284), .A2(P2_U3152), .ZN(n7364) );
  INV_X1 U8327 ( .A(n7364), .ZN(n7083) );
  AOI22_X1 U8328 ( .A1(n10281), .A2(n9068), .B1(n7083), .B2(
        P2_REG3_REG_0__SCAN_IN), .ZN(n7086) );
  AOI21_X1 U8329 ( .B1(n6952), .B2(n5621), .A(n10288), .ZN(n7084) );
  OAI21_X1 U8330 ( .B1(n7084), .B2(n10293), .A(n7313), .ZN(n7085) );
  OAI211_X1 U8331 ( .C1(n9017), .C2(n8752), .A(n7086), .B(n7085), .ZN(P2_U3234) );
  INV_X1 U8332 ( .A(P2_REG3_REG_2__SCAN_IN), .ZN(n10148) );
  INV_X1 U8333 ( .A(n7223), .ZN(n7087) );
  AOI211_X1 U8334 ( .C1(n7089), .C2(n7088), .A(n7087), .B(n10288), .ZN(n7090)
         );
  AOI21_X1 U8335 ( .B1(n6257), .B2(n10293), .A(n7090), .ZN(n7092) );
  NAND2_X1 U8336 ( .A1(n9049), .A2(n9239), .ZN(n8939) );
  AOI22_X1 U8337 ( .A1(n10281), .A2(n6259), .B1(n10282), .B2(n9068), .ZN(n7091) );
  OAI211_X1 U8338 ( .C1(n7364), .C2(n10148), .A(n7092), .B(n7091), .ZN(
        P2_U3239) );
  INV_X1 U8339 ( .A(P1_ADDR_REG_12__SCAN_IN), .ZN(n7100) );
  INV_X1 U8340 ( .A(P1_REG3_REG_12__SCAN_IN), .ZN(n7093) );
  NOR2_X1 U8341 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n7093), .ZN(n7801) );
  INV_X1 U8342 ( .A(n7801), .ZN(n7099) );
  AOI21_X1 U8343 ( .B1(n7096), .B2(n7095), .A(n7094), .ZN(n7097) );
  OR2_X1 U8344 ( .A1(n10380), .A2(n7097), .ZN(n7098) );
  OAI211_X1 U8345 ( .C1(n10391), .C2(n7100), .A(n7099), .B(n7098), .ZN(n7105)
         );
  AOI211_X1 U8346 ( .C1(n7103), .C2(n7102), .A(n7101), .B(n9673), .ZN(n7104)
         );
  AOI211_X1 U8347 ( .C1(n9678), .C2(n7730), .A(n7105), .B(n7104), .ZN(n7106)
         );
  INV_X1 U8348 ( .A(n7106), .ZN(P1_U3253) );
  AND2_X1 U8349 ( .A1(n7107), .A2(n8683), .ZN(n7108) );
  NAND2_X1 U8350 ( .A1(n9841), .A2(n7108), .ZN(n9853) );
  NAND2_X1 U8351 ( .A1(n8569), .A2(n4989), .ZN(n7109) );
  NAND2_X1 U8352 ( .A1(n7111), .A2(n9626), .ZN(n8557) );
  NAND2_X1 U8353 ( .A1(n7231), .A2(n7169), .ZN(n7172) );
  NAND2_X1 U8354 ( .A1(n8557), .A2(n7172), .ZN(n8362) );
  INV_X1 U8355 ( .A(n8362), .ZN(n7115) );
  OAI21_X1 U8356 ( .B1(n5480), .B2(n8362), .A(n7166), .ZN(n7234) );
  AND2_X2 U8357 ( .A1(n7112), .A2(n7111), .ZN(n7179) );
  OAI21_X1 U8358 ( .B1(n7112), .B2(n7111), .A(n10617), .ZN(n7113) );
  OR2_X1 U8359 ( .A1(n7179), .A2(n7113), .ZN(n7229) );
  NAND2_X1 U8360 ( .A1(n10528), .A2(n4989), .ZN(n8570) );
  XNOR2_X1 U8361 ( .A(n7170), .B(n7115), .ZN(n7116) );
  AOI222_X1 U8362 ( .A1(n9628), .A2(n10622), .B1(n9625), .B2(n10623), .C1(
        n9891), .C2(n7116), .ZN(n7233) );
  OAI21_X1 U8363 ( .B1(n9772), .B2(n7229), .A(n7233), .ZN(n7117) );
  NAND2_X1 U8364 ( .A1(n7117), .A2(n9841), .ZN(n7123) );
  INV_X1 U8365 ( .A(n7118), .ZN(n7119) );
  OAI22_X1 U8366 ( .A1(n9841), .A2(n7120), .B1(n7119), .B2(n9866), .ZN(n7121)
         );
  AOI21_X1 U8367 ( .B1(n10640), .B2(n7231), .A(n7121), .ZN(n7122) );
  OAI211_X1 U8368 ( .C1(n9853), .C2(n7234), .A(n7123), .B(n7122), .ZN(P1_U3286) );
  NAND2_X1 U8369 ( .A1(n7125), .A2(n7124), .ZN(n7127) );
  OR2_X1 U8370 ( .A1(n7128), .A2(n6792), .ZN(n7131) );
  AOI22_X1 U8371 ( .A1(n8153), .A2(P2_DATAO_REG_6__SCAN_IN), .B1(n5192), .B2(
        n7129), .ZN(n7130) );
  NAND2_X1 U8372 ( .A1(n7131), .A2(n7130), .ZN(n7201) );
  NAND2_X1 U8373 ( .A1(n7201), .A2(n8672), .ZN(n7133) );
  NAND2_X1 U8374 ( .A1(n9625), .A2(n8678), .ZN(n7132) );
  NAND2_X1 U8375 ( .A1(n7133), .A2(n7132), .ZN(n7134) );
  XNOR2_X1 U8376 ( .A(n7134), .B(n8675), .ZN(n7285) );
  NOR2_X1 U8377 ( .A1(n7167), .A2(n8682), .ZN(n7135) );
  AOI21_X1 U8378 ( .B1(n7201), .B2(n8678), .A(n7135), .ZN(n7284) );
  XNOR2_X1 U8379 ( .A(n7285), .B(n7284), .ZN(n7137) );
  NAND2_X1 U8380 ( .A1(n7136), .A2(n7137), .ZN(n7138) );
  AOI21_X1 U8381 ( .B1(n7452), .B2(n7138), .A(n9609), .ZN(n7156) );
  NAND2_X1 U8382 ( .A1(n7201), .A2(n9607), .ZN(n7154) );
  AOI21_X1 U8383 ( .B1(n9566), .B2(n9626), .A(n7139), .ZN(n7153) );
  NAND2_X1 U8384 ( .A1(n9602), .A2(n7180), .ZN(n7152) );
  INV_X1 U8385 ( .A(n7188), .ZN(n7144) );
  NAND2_X1 U8386 ( .A1(n7142), .A2(n7141), .ZN(n7143) );
  AND2_X1 U8387 ( .A1(n7144), .A2(n7143), .ZN(n7288) );
  NAND2_X1 U8388 ( .A1(n4856), .A2(n7288), .ZN(n7150) );
  NAND2_X1 U8389 ( .A1(n6774), .A2(P1_REG1_REG_7__SCAN_IN), .ZN(n7149) );
  OR2_X1 U8390 ( .A1(n8268), .A2(n7145), .ZN(n7148) );
  INV_X1 U8391 ( .A(P1_REG0_REG_7__SCAN_IN), .ZN(n7146) );
  OR2_X1 U8392 ( .A1(n8270), .A2(n7146), .ZN(n7147) );
  NAND2_X1 U8393 ( .A1(n9601), .A2(n9624), .ZN(n7151) );
  NAND4_X1 U8394 ( .A1(n7154), .A2(n7153), .A3(n7152), .A4(n7151), .ZN(n7155)
         );
  OR2_X1 U8395 ( .A1(n7156), .A2(n7155), .ZN(P1_U3237) );
  AOI22_X1 U8396 ( .A1(n9090), .A2(P2_STATE_REG_SCAN_IN), .B1(
        P1_DATAO_REG_18__SCAN_IN), .B2(n9487), .ZN(n7157) );
  OAI21_X1 U8397 ( .B1(n8142), .B2(n4857), .A(n7157), .ZN(P2_U3340) );
  INV_X1 U8398 ( .A(n8968), .ZN(n7158) );
  AOI211_X1 U8399 ( .C1(n7160), .C2(n7159), .A(n10288), .B(n7158), .ZN(n7164)
         );
  INV_X1 U8400 ( .A(n7478), .ZN(n9064) );
  AOI22_X1 U8401 ( .A1(n10282), .A2(n8781), .B1(n10281), .B2(n9064), .ZN(n7162) );
  AOI22_X1 U8402 ( .A1(n10284), .A2(n7484), .B1(P2_U3152), .B2(
        P2_REG3_REG_7__SCAN_IN), .ZN(n7161) );
  OAI211_X1 U8403 ( .C1(n10570), .C2(n9046), .A(n7162), .B(n7161), .ZN(n7163)
         );
  OR2_X1 U8404 ( .A1(n7164), .A2(n7163), .ZN(P2_U3215) );
  NAND2_X1 U8405 ( .A1(n7231), .A2(n9626), .ZN(n7165) );
  OR2_X1 U8406 ( .A1(n7201), .A2(n7167), .ZN(n7516) );
  NAND2_X1 U8407 ( .A1(n7201), .A2(n7167), .ZN(n8577) );
  NAND2_X1 U8408 ( .A1(n7516), .A2(n8577), .ZN(n8364) );
  OAI21_X1 U8409 ( .B1(n7168), .B2(n8364), .A(n7203), .ZN(n10558) );
  OAI22_X1 U8410 ( .A1(n7169), .A2(n9879), .B1(n7519), .B2(n9881), .ZN(n7177)
         );
  AND2_X1 U8411 ( .A1(n8577), .A2(n7172), .ZN(n8571) );
  INV_X1 U8412 ( .A(n7518), .ZN(n7175) );
  INV_X1 U8413 ( .A(n8364), .ZN(n7171) );
  AOI21_X1 U8414 ( .B1(n7173), .B2(n7172), .A(n7171), .ZN(n7174) );
  AOI211_X1 U8415 ( .C1(n7175), .C2(n7516), .A(n10626), .B(n7174), .ZN(n7176)
         );
  AOI211_X1 U8416 ( .C1(n10629), .C2(n10558), .A(n7177), .B(n7176), .ZN(n10555) );
  MUX2_X1 U8417 ( .A(n7178), .B(n10555), .S(n9841), .Z(n7184) );
  INV_X1 U8418 ( .A(n7201), .ZN(n10553) );
  NAND2_X1 U8419 ( .A1(n7179), .A2(n10553), .ZN(n7206) );
  OAI21_X1 U8420 ( .B1(n7179), .B2(n10553), .A(n7206), .ZN(n10554) );
  INV_X1 U8421 ( .A(n9902), .ZN(n9870) );
  AOI22_X1 U8422 ( .A1(n10640), .A2(n7201), .B1(n7180), .B2(n10638), .ZN(n7181) );
  OAI21_X1 U8423 ( .B1(n10554), .B2(n9870), .A(n7181), .ZN(n7182) );
  AOI21_X1 U8424 ( .B1(n10558), .B2(n10645), .A(n7182), .ZN(n7183) );
  NAND2_X1 U8425 ( .A1(n7184), .A2(n7183), .ZN(P1_U3285) );
  NAND2_X1 U8426 ( .A1(n7185), .A2(P1_IR_REG_31__SCAN_IN), .ZN(n7186) );
  XNOR2_X1 U8427 ( .A(n7186), .B(P1_IR_REG_18__SCAN_IN), .ZN(n9686) );
  INV_X1 U8428 ( .A(n9686), .ZN(n9682) );
  INV_X1 U8429 ( .A(P2_DATAO_REG_18__SCAN_IN), .ZN(n7187) );
  OAI222_X1 U8430 ( .A1(n10043), .A2(n8142), .B1(n9682), .B2(P1_U3084), .C1(
        n7187), .C2(n10039), .ZN(P1_U3335) );
  OR2_X1 U8431 ( .A1(n7188), .A2(P1_REG3_REG_8__SCAN_IN), .ZN(n7189) );
  AND2_X1 U8432 ( .A1(n7464), .A2(n7189), .ZN(n7606) );
  NAND2_X1 U8433 ( .A1(n4856), .A2(n7606), .ZN(n7194) );
  NAND2_X1 U8434 ( .A1(n6774), .A2(P1_REG1_REG_8__SCAN_IN), .ZN(n7193) );
  OR2_X1 U8435 ( .A1(n8268), .A2(n6339), .ZN(n7192) );
  INV_X1 U8436 ( .A(P1_REG0_REG_8__SCAN_IN), .ZN(n7190) );
  OR2_X1 U8437 ( .A1(n8270), .A2(n7190), .ZN(n7191) );
  INV_X1 U8438 ( .A(n7562), .ZN(n9623) );
  NAND2_X1 U8439 ( .A1(n7518), .A2(n7516), .ZN(n7199) );
  OR2_X1 U8440 ( .A1(n7195), .A2(n6792), .ZN(n7198) );
  AOI22_X1 U8441 ( .A1(n8153), .A2(P2_DATAO_REG_7__SCAN_IN), .B1(n5192), .B2(
        n7196), .ZN(n7197) );
  XNOR2_X1 U8442 ( .A(n7520), .B(n9624), .ZN(n8365) );
  INV_X1 U8443 ( .A(n8365), .ZN(n7204) );
  XNOR2_X1 U8444 ( .A(n7199), .B(n7204), .ZN(n7200) );
  AOI222_X1 U8445 ( .A1(n9625), .A2(n10622), .B1(n9623), .B2(n10623), .C1(
        n9891), .C2(n7200), .ZN(n7383) );
  OR2_X1 U8446 ( .A1(n7201), .A2(n9625), .ZN(n7202) );
  NAND2_X1 U8447 ( .A1(n7203), .A2(n7202), .ZN(n7205) );
  OAI21_X1 U8448 ( .B1(n7205), .B2(n7204), .A(n7508), .ZN(n7380) );
  INV_X1 U8449 ( .A(n9853), .ZN(n7214) );
  INV_X1 U8450 ( .A(n7520), .ZN(n7212) );
  AOI21_X1 U8451 ( .B1(n7206), .B2(n7520), .A(n10597), .ZN(n7207) );
  OR2_X2 U8452 ( .A1(n7206), .A2(n7520), .ZN(n7605) );
  AND2_X1 U8453 ( .A1(n7207), .A2(n7605), .ZN(n7381) );
  INV_X1 U8454 ( .A(n7208), .ZN(n7209) );
  NAND2_X1 U8455 ( .A1(n7209), .A2(n6904), .ZN(n8060) );
  INV_X1 U8456 ( .A(n8060), .ZN(n10644) );
  NAND2_X1 U8457 ( .A1(n7381), .A2(n10644), .ZN(n7211) );
  AOI22_X1 U8458 ( .A1(n9896), .A2(P1_REG2_REG_7__SCAN_IN), .B1(n7288), .B2(
        n10638), .ZN(n7210) );
  OAI211_X1 U8459 ( .C1(n7212), .C2(n9898), .A(n7211), .B(n7210), .ZN(n7213)
         );
  AOI21_X1 U8460 ( .B1(n7380), .B2(n7214), .A(n7213), .ZN(n7215) );
  OAI21_X1 U8461 ( .B1(n7383), .B2(n9896), .A(n7215), .ZN(P1_U3284) );
  INV_X1 U8462 ( .A(P2_REG3_REG_3__SCAN_IN), .ZN(n7216) );
  OAI22_X1 U8463 ( .A1(n9044), .A2(P2_REG3_REG_3__SCAN_IN), .B1(
        P2_STATE_REG_SCAN_IN), .B2(n7216), .ZN(n7219) );
  OAI22_X1 U8464 ( .A1(n5071), .A2(n8939), .B1(n9015), .B2(n7217), .ZN(n7218)
         );
  AOI211_X1 U8465 ( .C1(n7348), .C2(n10293), .A(n7219), .B(n7218), .ZN(n7228)
         );
  NOR3_X1 U8466 ( .A1(n9017), .A2(n5071), .A3(n7220), .ZN(n7226) );
  INV_X1 U8467 ( .A(n7221), .ZN(n7222) );
  AOI21_X1 U8468 ( .B1(n7223), .B2(n7222), .A(n10288), .ZN(n7225) );
  OAI21_X1 U8469 ( .B1(n7226), .B2(n7225), .A(n7224), .ZN(n7227) );
  NAND2_X1 U8470 ( .A1(n7228), .A2(n7227), .ZN(P2_U3220) );
  INV_X1 U8471 ( .A(P1_REG0_REG_5__SCAN_IN), .ZN(n7236) );
  INV_X1 U8472 ( .A(n10582), .ZN(n10632) );
  NOR2_X2 U8473 ( .A1(n10629), .A2(n10632), .ZN(n10001) );
  INV_X1 U8474 ( .A(n7229), .ZN(n7230) );
  AOI21_X1 U8475 ( .B1(n10578), .B2(n7231), .A(n7230), .ZN(n7232) );
  OAI211_X1 U8476 ( .C1(n10001), .C2(n7234), .A(n7233), .B(n7232), .ZN(n7237)
         );
  NAND2_X1 U8477 ( .A1(n7237), .A2(n10637), .ZN(n7235) );
  OAI21_X1 U8478 ( .B1(n10637), .B2(n7236), .A(n7235), .ZN(P1_U3469) );
  INV_X1 U8479 ( .A(P1_REG1_REG_5__SCAN_IN), .ZN(n7239) );
  NAND2_X1 U8480 ( .A1(n7237), .A2(n10634), .ZN(n7238) );
  OAI21_X1 U8481 ( .B1(n10634), .B2(n7239), .A(n7238), .ZN(P1_U3528) );
  INV_X1 U8482 ( .A(n7240), .ZN(n7331) );
  NAND2_X1 U8483 ( .A1(P2_REG3_REG_6__SCAN_IN), .A2(P2_U3152), .ZN(n10489) );
  OAI21_X1 U8484 ( .B1(n9044), .B2(n7331), .A(n10489), .ZN(n7242) );
  OAI22_X1 U8485 ( .A1(n7330), .A2(n8939), .B1(n9015), .B2(n8970), .ZN(n7241)
         );
  AOI211_X1 U8486 ( .C1(n8784), .C2(n10293), .A(n7242), .B(n7241), .ZN(n7249)
         );
  OAI22_X1 U8487 ( .A1(n9017), .A2(n7330), .B1(n7243), .B2(n10288), .ZN(n7247)
         );
  INV_X1 U8488 ( .A(n7244), .ZN(n7246) );
  NAND3_X1 U8489 ( .A1(n7247), .A2(n7246), .A3(n7245), .ZN(n7248) );
  OAI211_X1 U8490 ( .C1(n10288), .C2(n7250), .A(n7249), .B(n7248), .ZN(
        P2_U3241) );
  INV_X1 U8491 ( .A(n7251), .ZN(n7252) );
  AOI21_X1 U8492 ( .B1(P2_REG2_REG_12__SCAN_IN), .B2(n7253), .A(n7252), .ZN(
        n7256) );
  INV_X1 U8493 ( .A(P2_REG2_REG_13__SCAN_IN), .ZN(n7254) );
  AOI22_X1 U8494 ( .A1(n7395), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n7254), .B2(
        n7390), .ZN(n7255) );
  NAND2_X1 U8495 ( .A1(n7256), .A2(n7255), .ZN(n7394) );
  OAI21_X1 U8496 ( .B1(n7256), .B2(n7255), .A(n7394), .ZN(n7266) );
  INV_X1 U8497 ( .A(n7257), .ZN(n7258) );
  AOI21_X1 U8498 ( .B1(n10670), .B2(n7259), .A(n7258), .ZN(n7261) );
  INV_X1 U8499 ( .A(P2_REG1_REG_13__SCAN_IN), .ZN(n10680) );
  AOI22_X1 U8500 ( .A1(n7395), .A2(n10680), .B1(P2_REG1_REG_13__SCAN_IN), .B2(
        n7390), .ZN(n7260) );
  NOR2_X1 U8501 ( .A1(n7261), .A2(n7260), .ZN(n7389) );
  AOI21_X1 U8502 ( .B1(n7261), .B2(n7260), .A(n7389), .ZN(n7264) );
  INV_X1 U8503 ( .A(n10414), .ZN(n10478) );
  NAND2_X1 U8504 ( .A1(n10478), .A2(n7395), .ZN(n7263) );
  AOI22_X1 U8505 ( .A1(n10486), .A2(P2_ADDR_REG_13__SCAN_IN), .B1(
        P2_REG3_REG_13__SCAN_IN), .B2(P2_U3152), .ZN(n7262) );
  OAI211_X1 U8506 ( .C1(n10481), .C2(n7264), .A(n7263), .B(n7262), .ZN(n7265)
         );
  AOI21_X1 U8507 ( .B1(n10480), .B2(n7266), .A(n7265), .ZN(n7267) );
  INV_X1 U8508 ( .A(n7267), .ZN(P2_U3258) );
  INV_X1 U8509 ( .A(P1_ADDR_REG_13__SCAN_IN), .ZN(n7279) );
  AOI211_X1 U8510 ( .C1(n7270), .C2(n7269), .A(n7268), .B(n9673), .ZN(n7271)
         );
  AOI21_X1 U8511 ( .B1(n9678), .B2(n7852), .A(n7271), .ZN(n7278) );
  AOI21_X1 U8512 ( .B1(n7274), .B2(n7273), .A(n7272), .ZN(n7275) );
  NOR2_X1 U8513 ( .A1(n10380), .A2(n7275), .ZN(n7276) );
  AND2_X1 U8514 ( .A1(P1_U3084), .A2(P1_REG3_REG_13__SCAN_IN), .ZN(n7957) );
  NOR2_X1 U8515 ( .A1(n7276), .A2(n7957), .ZN(n7277) );
  OAI211_X1 U8516 ( .C1(n7279), .C2(n10391), .A(n7278), .B(n7277), .ZN(
        P1_U3254) );
  NAND2_X1 U8517 ( .A1(n7520), .A2(n8672), .ZN(n7281) );
  NAND2_X1 U8518 ( .A1(n9624), .A2(n8678), .ZN(n7280) );
  NAND2_X1 U8519 ( .A1(n7281), .A2(n7280), .ZN(n7282) );
  XNOR2_X1 U8520 ( .A(n7282), .B(n8683), .ZN(n7447) );
  NOR2_X1 U8521 ( .A1(n7519), .A2(n8682), .ZN(n7283) );
  AOI21_X1 U8522 ( .B1(n7520), .B2(n8678), .A(n7283), .ZN(n7448) );
  XNOR2_X1 U8523 ( .A(n7447), .B(n7448), .ZN(n7454) );
  NAND2_X1 U8524 ( .A1(n7285), .A2(n7284), .ZN(n7450) );
  NAND2_X1 U8525 ( .A1(n7452), .A2(n7450), .ZN(n7286) );
  XOR2_X1 U8526 ( .A(n7454), .B(n7286), .Z(n7293) );
  AOI21_X1 U8527 ( .B1(n9566), .B2(n9625), .A(n7287), .ZN(n7290) );
  NAND2_X1 U8528 ( .A1(n9602), .A2(n7288), .ZN(n7289) );
  OAI211_X1 U8529 ( .C1(n7562), .C2(n9569), .A(n7290), .B(n7289), .ZN(n7291)
         );
  AOI21_X1 U8530 ( .B1(n7520), .B2(n9607), .A(n7291), .ZN(n7292) );
  OAI21_X1 U8531 ( .B1(n7293), .B2(n9609), .A(n7292), .ZN(P1_U3211) );
  OAI21_X1 U8532 ( .B1(n7295), .B2(n8768), .A(n7294), .ZN(n10536) );
  INV_X1 U8533 ( .A(n7296), .ZN(n7297) );
  NAND2_X1 U8534 ( .A1(n7297), .A2(n5542), .ZN(n9152) );
  OR2_X1 U8535 ( .A1(n7298), .A2(n10537), .ZN(n7299) );
  NAND2_X1 U8536 ( .A1(n7406), .A2(n7299), .ZN(n10538) );
  OAI22_X1 U8537 ( .A1(n9152), .A2(n10538), .B1(n7372), .B2(n9316), .ZN(n7300)
         );
  AOI21_X1 U8538 ( .B1(n9366), .B2(n7301), .A(n7300), .ZN(n7310) );
  OAI21_X1 U8539 ( .B1(n8903), .B2(n7303), .A(n7302), .ZN(n7304) );
  NAND2_X1 U8540 ( .A1(n7304), .A2(n9349), .ZN(n7306) );
  AOI22_X1 U8541 ( .A1(n9239), .A2(n6259), .B1(n7374), .B2(n9241), .ZN(n7305)
         );
  NAND2_X1 U8542 ( .A1(n7306), .A2(n7305), .ZN(n10539) );
  NOR2_X1 U8543 ( .A1(n9378), .A2(n7307), .ZN(n7308) );
  AOI21_X1 U8544 ( .B1(n9378), .B2(n10539), .A(n7308), .ZN(n7309) );
  OAI211_X1 U8545 ( .C1(n9359), .C2(n10536), .A(n7310), .B(n7309), .ZN(
        P2_U3292) );
  INV_X1 U8546 ( .A(P2_REG2_REG_0__SCAN_IN), .ZN(n10422) );
  AOI21_X1 U8547 ( .B1(P2_REG3_REG_0__SCAN_IN), .B2(n9377), .A(n7311), .ZN(
        n7312) );
  MUX2_X1 U8548 ( .A(n10422), .B(n7312), .S(n9378), .Z(n7315) );
  OAI21_X1 U8549 ( .B1(n9366), .B2(n9380), .A(n7313), .ZN(n7314) );
  OAI211_X1 U8550 ( .C1(n7316), .C2(n9359), .A(n7315), .B(n7314), .ZN(P2_U3296) );
  NAND2_X1 U8551 ( .A1(n8753), .A2(n8751), .ZN(n7322) );
  XNOR2_X1 U8552 ( .A(n7322), .B(n7352), .ZN(n10502) );
  NOR2_X1 U8553 ( .A1(n10505), .A2(n7317), .ZN(n10503) );
  NOR3_X1 U8554 ( .A1(n9152), .A2(n5212), .A3(n10503), .ZN(n7318) );
  INV_X1 U8555 ( .A(n7322), .ZN(n7320) );
  OAI21_X1 U8556 ( .B1(n7320), .B2(n7319), .A(n9349), .ZN(n7324) );
  NOR2_X1 U8557 ( .A1(n7322), .A2(n7321), .ZN(n8901) );
  AOI22_X1 U8558 ( .A1(n9239), .A2(n6952), .B1(n9067), .B2(n9241), .ZN(n7323)
         );
  OAI21_X1 U8559 ( .B1(n7324), .B2(n8901), .A(n7323), .ZN(n10506) );
  AOI21_X1 U8560 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(n9377), .A(n10506), .ZN(
        n7325) );
  MUX2_X1 U8561 ( .A(n6661), .B(n7325), .S(n9378), .Z(n7326) );
  OAI211_X1 U8562 ( .C1(n10502), .C2(n9359), .A(n7327), .B(n7326), .ZN(
        P2_U3295) );
  XNOR2_X1 U8563 ( .A(n7328), .B(n8906), .ZN(n7329) );
  OAI222_X1 U8564 ( .A1(n9370), .A2(n8970), .B1(n9371), .B2(n7330), .C1(n9376), 
        .C2(n7329), .ZN(n10564) );
  INV_X1 U8565 ( .A(n10564), .ZN(n7342) );
  OAI22_X1 U8566 ( .A1(n9378), .A2(n10474), .B1(n7331), .B2(n9316), .ZN(n7336)
         );
  INV_X1 U8567 ( .A(n7481), .ZN(n7334) );
  NAND2_X1 U8568 ( .A1(n7332), .A2(n8784), .ZN(n7333) );
  NAND2_X1 U8569 ( .A1(n7334), .A2(n7333), .ZN(n10563) );
  NOR2_X1 U8570 ( .A1(n9152), .A2(n10563), .ZN(n7335) );
  AOI211_X1 U8571 ( .C1(n9366), .C2(n8784), .A(n7336), .B(n7335), .ZN(n7341)
         );
  NOR2_X1 U8572 ( .A1(n7337), .A2(n8906), .ZN(n10561) );
  INV_X1 U8573 ( .A(n10561), .ZN(n7339) );
  NAND3_X1 U8574 ( .A1(n7339), .A2(n9289), .A3(n7338), .ZN(n7340) );
  OAI211_X1 U8575 ( .C1(n7342), .C2(n9268), .A(n7341), .B(n7340), .ZN(P2_U3290) );
  OAI22_X1 U8576 ( .A1(n7343), .A2(n9268), .B1(P2_REG3_REG_3__SCAN_IN), .B2(
        n9316), .ZN(n7346) );
  OAI22_X1 U8577 ( .A1(n9152), .A2(n7344), .B1(n9378), .B2(n6660), .ZN(n7345)
         );
  NOR2_X1 U8578 ( .A1(n7346), .A2(n7345), .ZN(n7351) );
  NOR2_X1 U8579 ( .A1(n9268), .A2(n7347), .ZN(n9367) );
  AOI22_X1 U8580 ( .A1(n9367), .A2(n7349), .B1(n9366), .B2(n7348), .ZN(n7350)
         );
  NAND2_X1 U8581 ( .A1(n7351), .A2(n7350), .ZN(P2_U3293) );
  INV_X1 U8582 ( .A(P2_REG3_REG_1__SCAN_IN), .ZN(n7363) );
  NOR2_X1 U8583 ( .A1(n9046), .A2(n10505), .ZN(n7355) );
  INV_X1 U8584 ( .A(n7352), .ZN(n7353) );
  NOR3_X1 U8585 ( .A1(n9017), .A2(n7358), .A3(n7353), .ZN(n7354) );
  AOI211_X1 U8586 ( .C1(n10282), .C2(n6952), .A(n7355), .B(n7354), .ZN(n7362)
         );
  INV_X1 U8587 ( .A(n7356), .ZN(n7359) );
  OAI21_X1 U8588 ( .B1(n7359), .B2(n7358), .A(n7357), .ZN(n7360) );
  AOI22_X1 U8589 ( .A1(n10281), .A2(n9067), .B1(n9009), .B2(n7360), .ZN(n7361)
         );
  OAI211_X1 U8590 ( .C1(n7364), .C2(n7363), .A(n7362), .B(n7361), .ZN(P2_U3224) );
  INV_X1 U8591 ( .A(n8152), .ZN(n7366) );
  INV_X1 U8592 ( .A(P1_DATAO_REG_19__SCAN_IN), .ZN(n7365) );
  OAI222_X1 U8593 ( .A1(n5298), .A2(P2_U3152), .B1(n4857), .B2(n7366), .C1(
        n7365), .C2(n9491), .ZN(P2_U3339) );
  INV_X1 U8594 ( .A(P2_DATAO_REG_19__SCAN_IN), .ZN(n7367) );
  OAI222_X1 U8595 ( .A1(n10039), .A2(n7367), .B1(n10033), .B2(n7366), .C1(
        P1_U3084), .C2(n6904), .ZN(P1_U3334) );
  OAI21_X1 U8596 ( .B1(n7368), .B2(n7224), .A(n7419), .ZN(n7378) );
  NOR3_X1 U8597 ( .A1(n9017), .A2(n7369), .A3(n7368), .ZN(n7370) );
  OAI21_X1 U8598 ( .B1(n7370), .B2(n10282), .A(n6259), .ZN(n7376) );
  OAI21_X1 U8599 ( .B1(n9044), .B2(n7372), .A(n7371), .ZN(n7373) );
  AOI21_X1 U8600 ( .B1(n10281), .B2(n7374), .A(n7373), .ZN(n7375) );
  OAI211_X1 U8601 ( .C1(n10537), .C2(n9046), .A(n7376), .B(n7375), .ZN(n7377)
         );
  AOI21_X1 U8602 ( .B1(n9009), .B2(n7378), .A(n7377), .ZN(n7379) );
  INV_X1 U8603 ( .A(n7379), .ZN(P2_U3232) );
  INV_X1 U8604 ( .A(n7380), .ZN(n7384) );
  AOI21_X1 U8605 ( .B1(n10578), .B2(n7520), .A(n7381), .ZN(n7382) );
  OAI211_X1 U8606 ( .C1(n10001), .C2(n7384), .A(n7383), .B(n7382), .ZN(n7386)
         );
  NAND2_X1 U8607 ( .A1(n7386), .A2(n10637), .ZN(n7385) );
  OAI21_X1 U8608 ( .B1(n10637), .B2(n7146), .A(n7385), .ZN(P1_U3475) );
  INV_X1 U8609 ( .A(P1_REG1_REG_7__SCAN_IN), .ZN(n7388) );
  NAND2_X1 U8610 ( .A1(n7386), .A2(n10634), .ZN(n7387) );
  OAI21_X1 U8611 ( .B1(n10634), .B2(n7388), .A(n7387), .ZN(P1_U3530) );
  AOI21_X1 U8612 ( .B1(n7390), .B2(n10680), .A(n7389), .ZN(n7392) );
  INV_X1 U8613 ( .A(P2_REG1_REG_14__SCAN_IN), .ZN(n10688) );
  AOI22_X1 U8614 ( .A1(n7680), .A2(n10688), .B1(P2_REG1_REG_14__SCAN_IN), .B2(
        n7685), .ZN(n7391) );
  NOR2_X1 U8615 ( .A1(n7392), .A2(n7391), .ZN(n7684) );
  AOI21_X1 U8616 ( .B1(n7392), .B2(n7391), .A(n7684), .ZN(n7402) );
  INV_X1 U8617 ( .A(P2_REG2_REG_14__SCAN_IN), .ZN(n7393) );
  AOI22_X1 U8618 ( .A1(n7680), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7393), .B2(
        n7685), .ZN(n7397) );
  OAI21_X1 U8619 ( .B1(n7395), .B2(P2_REG2_REG_13__SCAN_IN), .A(n7394), .ZN(
        n7396) );
  NAND2_X1 U8620 ( .A1(n7397), .A2(n7396), .ZN(n7679) );
  OAI21_X1 U8621 ( .B1(n7397), .B2(n7396), .A(n7679), .ZN(n7400) );
  NAND2_X1 U8622 ( .A1(P2_U3152), .A2(P2_REG3_REG_14__SCAN_IN), .ZN(n7900) );
  NAND2_X1 U8623 ( .A1(n10486), .A2(P2_ADDR_REG_14__SCAN_IN), .ZN(n7398) );
  OAI211_X1 U8624 ( .C1(n10414), .C2(n7685), .A(n7900), .B(n7398), .ZN(n7399)
         );
  AOI21_X1 U8625 ( .B1(n7400), .B2(n10480), .A(n7399), .ZN(n7401) );
  OAI21_X1 U8626 ( .B1(n7402), .B2(n10481), .A(n7401), .ZN(P2_U3259) );
  XNOR2_X1 U8627 ( .A(n7403), .B(n8905), .ZN(n7404) );
  AOI22_X1 U8628 ( .A1(n9066), .A2(n9239), .B1(n9241), .B2(n8781), .ZN(n7417)
         );
  OAI21_X1 U8629 ( .B1(n7404), .B2(n9376), .A(n7417), .ZN(n10547) );
  INV_X1 U8630 ( .A(n10547), .ZN(n7414) );
  XNOR2_X1 U8631 ( .A(n8775), .B(n7405), .ZN(n10549) );
  XNOR2_X1 U8632 ( .A(n7406), .B(n10546), .ZN(n7407) );
  NAND2_X1 U8633 ( .A1(n7407), .A2(n5299), .ZN(n10545) );
  INV_X1 U8634 ( .A(n7415), .ZN(n7408) );
  OAI22_X1 U8635 ( .A1(n9378), .A2(n7409), .B1(n7408), .B2(n9316), .ZN(n7410)
         );
  AOI21_X1 U8636 ( .B1(n9366), .B2(n7425), .A(n7410), .ZN(n7411) );
  OAI21_X1 U8637 ( .B1(n8093), .B2(n10545), .A(n7411), .ZN(n7412) );
  AOI21_X1 U8638 ( .B1(n9289), .B2(n10549), .A(n7412), .ZN(n7413) );
  OAI21_X1 U8639 ( .B1(n9268), .B2(n7414), .A(n7413), .ZN(P2_U3291) );
  NAND2_X1 U8640 ( .A1(P2_U3152), .A2(P2_REG3_REG_5__SCAN_IN), .ZN(n10460) );
  NAND2_X1 U8641 ( .A1(n10284), .A2(n7415), .ZN(n7416) );
  OAI211_X1 U8642 ( .C1(n8994), .C2(n7417), .A(n10460), .B(n7416), .ZN(n7424)
         );
  INV_X1 U8643 ( .A(n9017), .ZN(n8956) );
  AOI22_X1 U8644 ( .A1(n8956), .A2(n9066), .B1(n9009), .B2(n7418), .ZN(n7422)
         );
  INV_X1 U8645 ( .A(n7419), .ZN(n7421) );
  NOR3_X1 U8646 ( .A1(n7422), .A2(n7421), .A3(n7420), .ZN(n7423) );
  AOI211_X1 U8647 ( .C1(n7425), .C2(n10293), .A(n7424), .B(n7423), .ZN(n7426)
         );
  OAI21_X1 U8648 ( .B1(n7245), .B2(n10288), .A(n7426), .ZN(P2_U3229) );
  INV_X1 U8649 ( .A(P1_ADDR_REG_14__SCAN_IN), .ZN(n7438) );
  AOI211_X1 U8650 ( .C1(n7429), .C2(n7428), .A(n7427), .B(n9673), .ZN(n7430)
         );
  AOI21_X1 U8651 ( .B1(n9678), .B2(n7858), .A(n7430), .ZN(n7437) );
  AOI21_X1 U8652 ( .B1(n7433), .B2(n7432), .A(n7431), .ZN(n7434) );
  NOR2_X1 U8653 ( .A1(n10380), .A2(n7434), .ZN(n7435) );
  NOR2_X1 U8654 ( .A1(n7861), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8073) );
  NOR2_X1 U8655 ( .A1(n7435), .A2(n8073), .ZN(n7436) );
  OAI211_X1 U8656 ( .C1(n7438), .C2(n10391), .A(n7437), .B(n7436), .ZN(
        P1_U3255) );
  NAND2_X1 U8657 ( .A1(n7440), .A2(n7439), .ZN(n7443) );
  AOI22_X1 U8658 ( .A1(n8153), .A2(P2_DATAO_REG_8__SCAN_IN), .B1(n5192), .B2(
        n7441), .ZN(n7442) );
  NAND2_X1 U8659 ( .A1(n7443), .A2(n7442), .ZN(n10577) );
  NAND2_X1 U8660 ( .A1(n10577), .A2(n6773), .ZN(n7445) );
  NAND2_X1 U8661 ( .A1(n9623), .A2(n8678), .ZN(n7444) );
  NAND2_X1 U8662 ( .A1(n7445), .A2(n7444), .ZN(n7446) );
  XNOR2_X1 U8663 ( .A(n7446), .B(n8683), .ZN(n7556) );
  INV_X1 U8664 ( .A(n7447), .ZN(n7449) );
  NAND2_X1 U8665 ( .A1(n7449), .A2(n7448), .ZN(n7453) );
  AND2_X1 U8666 ( .A1(n7450), .A2(n7453), .ZN(n7451) );
  INV_X1 U8667 ( .A(n7453), .ZN(n7455) );
  NOR2_X1 U8668 ( .A1(n7562), .A2(n8682), .ZN(n7456) );
  AOI21_X1 U8669 ( .B1(n10577), .B2(n8678), .A(n7456), .ZN(n7459) );
  INV_X1 U8670 ( .A(n7459), .ZN(n7457) );
  AND2_X1 U8671 ( .A1(n7459), .A2(n7458), .ZN(n7460) );
  NAND2_X1 U8672 ( .A1(n7558), .A2(n7557), .ZN(n7462) );
  XOR2_X1 U8673 ( .A(n7556), .B(n7462), .Z(n7475) );
  NAND2_X1 U8674 ( .A1(n6774), .A2(P1_REG1_REG_9__SCAN_IN), .ZN(n7469) );
  NAND2_X1 U8675 ( .A1(n7464), .A2(n7463), .ZN(n7465) );
  AND2_X1 U8676 ( .A1(n7523), .A2(n7465), .ZN(n7565) );
  NAND2_X1 U8677 ( .A1(n4856), .A2(n7565), .ZN(n7468) );
  NAND2_X1 U8678 ( .A1(n5475), .A2(P1_REG0_REG_9__SCAN_IN), .ZN(n7467) );
  OR2_X1 U8679 ( .A1(n8268), .A2(n6306), .ZN(n7466) );
  NAND4_X1 U8680 ( .A1(n7469), .A2(n7468), .A3(n7467), .A4(n7466), .ZN(n10621)
         );
  INV_X1 U8681 ( .A(n10621), .ZN(n7515) );
  AOI21_X1 U8682 ( .B1(n9566), .B2(n9624), .A(n7470), .ZN(n7472) );
  NAND2_X1 U8683 ( .A1(n9602), .A2(n7606), .ZN(n7471) );
  OAI211_X1 U8684 ( .C1(n7515), .C2(n9569), .A(n7472), .B(n7471), .ZN(n7473)
         );
  AOI21_X1 U8685 ( .B1(n10577), .B2(n9607), .A(n7473), .ZN(n7474) );
  OAI21_X1 U8686 ( .B1(n7475), .B2(n9609), .A(n7474), .ZN(P1_U3219) );
  XNOR2_X1 U8687 ( .A(n7476), .B(n8788), .ZN(n7477) );
  OAI222_X1 U8688 ( .A1(n9370), .A2(n7478), .B1(n7477), .B2(n9376), .C1(n9371), 
        .C2(n8785), .ZN(n10572) );
  INV_X1 U8689 ( .A(n10572), .ZN(n7489) );
  OAI21_X1 U8690 ( .B1(n7480), .B2(n5053), .A(n7479), .ZN(n10574) );
  NOR2_X1 U8691 ( .A1(n7481), .A2(n10570), .ZN(n7482) );
  OR2_X1 U8692 ( .A1(n7483), .A2(n7482), .ZN(n10571) );
  AOI22_X1 U8693 ( .A1(n9268), .A2(P2_REG2_REG_7__SCAN_IN), .B1(n7484), .B2(
        n9377), .ZN(n7486) );
  NAND2_X1 U8694 ( .A1(n9366), .A2(n8789), .ZN(n7485) );
  OAI211_X1 U8695 ( .C1(n9152), .C2(n10571), .A(n7486), .B(n7485), .ZN(n7487)
         );
  AOI21_X1 U8696 ( .B1(n10574), .B2(n9289), .A(n7487), .ZN(n7488) );
  OAI21_X1 U8697 ( .B1(n7489), .B2(n9268), .A(n7488), .ZN(P2_U3289) );
  NAND2_X1 U8698 ( .A1(n10605), .A2(n7582), .ZN(n8798) );
  NAND2_X1 U8699 ( .A1(n8975), .A2(n9064), .ZN(n7490) );
  NAND2_X1 U8700 ( .A1(n7491), .A2(n7490), .ZN(n7494) );
  INV_X1 U8701 ( .A(n7579), .ZN(n7493) );
  AOI21_X1 U8702 ( .B1(n8909), .B2(n7494), .A(n7493), .ZN(n7499) );
  INV_X1 U8703 ( .A(n9014), .ZN(n9063) );
  AOI22_X1 U8704 ( .A1(n9239), .A2(n9064), .B1(n9063), .B2(n9241), .ZN(n7498)
         );
  XNOR2_X1 U8705 ( .A(n7580), .B(n8909), .ZN(n7496) );
  NAND2_X1 U8706 ( .A1(n7496), .A2(n9349), .ZN(n7497) );
  OAI211_X1 U8707 ( .C1(n7499), .C2(n9369), .A(n7498), .B(n7497), .ZN(n10607)
         );
  INV_X1 U8708 ( .A(n10607), .ZN(n7506) );
  INV_X1 U8709 ( .A(n7499), .ZN(n10609) );
  OR2_X2 U8710 ( .A1(n7500), .A2(n10605), .ZN(n7587) );
  NAND2_X1 U8711 ( .A1(n7500), .A2(n10605), .ZN(n7501) );
  NAND2_X1 U8712 ( .A1(n7587), .A2(n7501), .ZN(n10606) );
  AOI22_X1 U8713 ( .A1(n9268), .A2(P2_REG2_REG_9__SCAN_IN), .B1(n9011), .B2(
        n9377), .ZN(n7503) );
  NAND2_X1 U8714 ( .A1(n9366), .A2(n10605), .ZN(n7502) );
  OAI211_X1 U8715 ( .C1(n10606), .C2(n9152), .A(n7503), .B(n7502), .ZN(n7504)
         );
  AOI21_X1 U8716 ( .B1(n10609), .B2(n9367), .A(n7504), .ZN(n7505) );
  OAI21_X1 U8717 ( .B1(n7506), .B2(n9268), .A(n7505), .ZN(P2_U3287) );
  OR2_X1 U8718 ( .A1(n7520), .A2(n9624), .ZN(n7507) );
  OR2_X1 U8719 ( .A1(n10577), .A2(n7562), .ZN(n8416) );
  AND2_X1 U8720 ( .A1(n10577), .A2(n7562), .ZN(n7521) );
  INV_X1 U8721 ( .A(n7521), .ZN(n8411) );
  INV_X1 U8722 ( .A(n8367), .ZN(n7509) );
  NAND2_X1 U8723 ( .A1(n10577), .A2(n9623), .ZN(n7510) );
  NAND2_X1 U8724 ( .A1(n7596), .A2(n7510), .ZN(n7643) );
  NAND2_X1 U8725 ( .A1(n7511), .A2(n7439), .ZN(n7514) );
  AOI22_X1 U8726 ( .A1(n8153), .A2(P2_DATAO_REG_9__SCAN_IN), .B1(n5192), .B2(
        n7512), .ZN(n7513) );
  OR2_X1 U8727 ( .A1(n7640), .A2(n7515), .ZN(n8472) );
  NAND2_X1 U8728 ( .A1(n7640), .A2(n7515), .ZN(n8407) );
  NAND2_X1 U8729 ( .A1(n8472), .A2(n8407), .ZN(n8356) );
  XNOR2_X1 U8730 ( .A(n7643), .B(n8356), .ZN(n10595) );
  INV_X1 U8731 ( .A(n10629), .ZN(n9887) );
  OR2_X1 U8732 ( .A1(n7520), .A2(n7519), .ZN(n7517) );
  AND2_X1 U8733 ( .A1(n7517), .A2(n7516), .ZN(n8558) );
  NAND2_X1 U8734 ( .A1(n7520), .A2(n7519), .ZN(n8410) );
  XNOR2_X1 U8735 ( .A(n8471), .B(n8356), .ZN(n7531) );
  NAND2_X1 U8736 ( .A1(n7523), .A2(n7522), .ZN(n7524) );
  AND2_X1 U8737 ( .A1(n7655), .A2(n7524), .ZN(n10639) );
  NAND2_X1 U8738 ( .A1(n4856), .A2(n10639), .ZN(n7529) );
  NAND2_X1 U8739 ( .A1(n6774), .A2(P1_REG1_REG_10__SCAN_IN), .ZN(n7528) );
  OR2_X1 U8740 ( .A1(n8268), .A2(n6301), .ZN(n7527) );
  INV_X1 U8741 ( .A(P1_REG0_REG_10__SCAN_IN), .ZN(n7525) );
  OR2_X1 U8742 ( .A1(n8270), .A2(n7525), .ZN(n7526) );
  OAI22_X1 U8743 ( .A1(n7767), .A2(n9881), .B1(n7562), .B2(n9879), .ZN(n7530)
         );
  AOI21_X1 U8744 ( .B1(n7531), .B2(n9891), .A(n7530), .ZN(n7532) );
  OAI21_X1 U8745 ( .B1(n10595), .B2(n9887), .A(n7532), .ZN(n10599) );
  NAND2_X1 U8746 ( .A1(n10599), .A2(n9841), .ZN(n7538) );
  INV_X1 U8747 ( .A(n7565), .ZN(n7533) );
  OAI22_X1 U8748 ( .A1(n9841), .A2(n6306), .B1(n7533), .B2(n9866), .ZN(n7536)
         );
  INV_X1 U8749 ( .A(n7640), .ZN(n10596) );
  OR2_X1 U8750 ( .A1(n10596), .A2(n7604), .ZN(n7534) );
  NAND2_X1 U8751 ( .A1(n10615), .A2(n7534), .ZN(n10598) );
  NOR2_X1 U8752 ( .A1(n10598), .A2(n9870), .ZN(n7535) );
  AOI211_X1 U8753 ( .C1(n10640), .C2(n7640), .A(n7536), .B(n7535), .ZN(n7537)
         );
  OAI211_X1 U8754 ( .C1(n10595), .C2(n9899), .A(n7538), .B(n7537), .ZN(
        P1_U3282) );
  INV_X1 U8755 ( .A(n7539), .ZN(n7540) );
  AOI21_X1 U8756 ( .B1(n7569), .B2(n7540), .A(n10288), .ZN(n7544) );
  NOR3_X1 U8757 ( .A1(n7541), .A2(n9014), .A3(n9017), .ZN(n7543) );
  OAI21_X1 U8758 ( .B1(n7544), .B2(n7543), .A(n7542), .ZN(n7551) );
  INV_X1 U8759 ( .A(n7545), .ZN(n7624) );
  OR2_X1 U8760 ( .A1(n9014), .A2(n9371), .ZN(n7547) );
  OR2_X1 U8761 ( .A1(n8804), .A2(n9370), .ZN(n7546) );
  NAND2_X1 U8762 ( .A1(n7547), .A2(n7546), .ZN(n7616) );
  AOI22_X1 U8763 ( .A1(n9049), .A2(n7616), .B1(P2_REG3_REG_11__SCAN_IN), .B2(
        P2_U3152), .ZN(n7548) );
  OAI21_X1 U8764 ( .B1(n9044), .B2(n7624), .A(n7548), .ZN(n7549) );
  AOI21_X1 U8765 ( .B1(n7693), .B2(n10293), .A(n7549), .ZN(n7550) );
  NAND2_X1 U8766 ( .A1(n7551), .A2(n7550), .ZN(P2_U3238) );
  NAND2_X1 U8767 ( .A1(n7640), .A2(n8672), .ZN(n7553) );
  NAND2_X1 U8768 ( .A1(n10621), .A2(n8678), .ZN(n7552) );
  NAND2_X1 U8769 ( .A1(n7553), .A2(n7552), .ZN(n7554) );
  XNOR2_X1 U8770 ( .A(n7554), .B(n8675), .ZN(n7708) );
  AND2_X1 U8771 ( .A1(n10621), .A2(n6799), .ZN(n7555) );
  AOI21_X1 U8772 ( .B1(n7640), .B2(n8678), .A(n7555), .ZN(n7707) );
  XNOR2_X1 U8773 ( .A(n7708), .B(n7707), .ZN(n7561) );
  INV_X1 U8774 ( .A(n7710), .ZN(n7560) );
  AOI21_X1 U8775 ( .B1(n7561), .B2(n7559), .A(n7560), .ZN(n7568) );
  NOR2_X1 U8776 ( .A1(n9569), .A2(n7767), .ZN(n7564) );
  OAI22_X1 U8777 ( .A1(n9605), .A2(n7562), .B1(P1_STATE_REG_SCAN_IN), .B2(
        n7463), .ZN(n7563) );
  AOI211_X1 U8778 ( .C1(n7565), .C2(n9602), .A(n7564), .B(n7563), .ZN(n7567)
         );
  NAND2_X1 U8779 ( .A1(n7640), .A2(n9607), .ZN(n7566) );
  OAI211_X1 U8780 ( .C1(n7568), .C2(n9609), .A(n7567), .B(n7566), .ZN(P1_U3229) );
  INV_X1 U8781 ( .A(n7569), .ZN(n7570) );
  AOI211_X1 U8782 ( .C1(n7572), .C2(n7571), .A(n10288), .B(n7570), .ZN(n7576)
         );
  INV_X1 U8783 ( .A(n7590), .ZN(n10650) );
  INV_X1 U8784 ( .A(n7694), .ZN(n9062) );
  AOI22_X1 U8785 ( .A1(n10282), .A2(n5120), .B1(n10281), .B2(n9062), .ZN(n7574) );
  AOI22_X1 U8786 ( .A1(n10284), .A2(n7589), .B1(P2_REG3_REG_10__SCAN_IN), .B2(
        P2_U3152), .ZN(n7573) );
  OAI211_X1 U8787 ( .C1(n10650), .C2(n9046), .A(n7574), .B(n7573), .ZN(n7575)
         );
  OR2_X1 U8788 ( .A1(n7576), .A2(n7575), .ZN(P2_U3219) );
  INV_X1 U8789 ( .A(n8167), .ZN(n7613) );
  INV_X1 U8790 ( .A(P2_DATAO_REG_20__SCAN_IN), .ZN(n8168) );
  OAI222_X1 U8791 ( .A1(n10043), .A2(n7613), .B1(n6579), .B2(P1_U3084), .C1(
        n8168), .C2(n10039), .ZN(P1_U3333) );
  OAI222_X1 U8792 ( .A1(P2_U3152), .A2(n8928), .B1(n4857), .B2(n8179), .C1(
        n7577), .C2(n9491), .ZN(P2_U3337) );
  OR2_X1 U8793 ( .A1(n10605), .A2(n5120), .ZN(n7578) );
  OR2_X1 U8794 ( .A1(n7590), .A2(n9014), .ZN(n8750) );
  NAND2_X1 U8795 ( .A1(n7590), .A2(n9014), .ZN(n8799) );
  NAND2_X1 U8796 ( .A1(n8750), .A2(n8799), .ZN(n8912) );
  INV_X1 U8797 ( .A(n8912), .ZN(n7618) );
  XNOR2_X1 U8798 ( .A(n7619), .B(n7618), .ZN(n7586) );
  XNOR2_X1 U8799 ( .A(n7615), .B(n8912), .ZN(n7584) );
  OAI22_X1 U8800 ( .A1(n7694), .A2(n9370), .B1(n7582), .B2(n9371), .ZN(n7583)
         );
  AOI21_X1 U8801 ( .B1(n7584), .B2(n9349), .A(n7583), .ZN(n7585) );
  OAI21_X1 U8802 ( .B1(n7586), .B2(n9369), .A(n7585), .ZN(n10652) );
  INV_X1 U8803 ( .A(n10652), .ZN(n7595) );
  INV_X1 U8804 ( .A(n7586), .ZN(n10654) );
  AND2_X1 U8805 ( .A1(n7590), .A2(n7587), .ZN(n7588) );
  OR2_X1 U8806 ( .A1(n7698), .A2(n7588), .ZN(n10651) );
  AOI22_X1 U8807 ( .A1(n9268), .A2(P2_REG2_REG_10__SCAN_IN), .B1(n7589), .B2(
        n9377), .ZN(n7592) );
  NAND2_X1 U8808 ( .A1(n7590), .A2(n9366), .ZN(n7591) );
  OAI211_X1 U8809 ( .C1(n10651), .C2(n9152), .A(n7592), .B(n7591), .ZN(n7593)
         );
  AOI21_X1 U8810 ( .B1(n10654), .B2(n9367), .A(n7593), .ZN(n7594) );
  OAI21_X1 U8811 ( .B1(n7595), .B2(n9268), .A(n7594), .ZN(P2_U3286) );
  INV_X1 U8812 ( .A(n7596), .ZN(n7597) );
  AOI21_X1 U8813 ( .B1(n8367), .B2(n7598), .A(n7597), .ZN(n7603) );
  INV_X1 U8814 ( .A(n7603), .ZN(n10583) );
  XOR2_X1 U8815 ( .A(n8367), .B(n7599), .Z(n7601) );
  AOI22_X1 U8816 ( .A1(n9624), .A2(n10622), .B1(n10623), .B2(n10621), .ZN(
        n7600) );
  OAI21_X1 U8817 ( .B1(n7601), .B2(n10626), .A(n7600), .ZN(n7602) );
  AOI21_X1 U8818 ( .B1(n7603), .B2(n10629), .A(n7602), .ZN(n10581) );
  MUX2_X1 U8819 ( .A(n6339), .B(n10581), .S(n9841), .Z(n7611) );
  AOI21_X1 U8820 ( .B1(n10577), .B2(n7605), .A(n7604), .ZN(n10579) );
  INV_X1 U8821 ( .A(n10577), .ZN(n7608) );
  INV_X1 U8822 ( .A(n7606), .ZN(n7607) );
  OAI22_X1 U8823 ( .A1(n7608), .A2(n9898), .B1(n7607), .B2(n9866), .ZN(n7609)
         );
  AOI21_X1 U8824 ( .B1(n10579), .B2(n9902), .A(n7609), .ZN(n7610) );
  OAI211_X1 U8825 ( .C1(n10583), .C2(n9899), .A(n7611), .B(n7610), .ZN(
        P1_U3283) );
  OAI222_X1 U8826 ( .A1(P2_U3152), .A2(n8926), .B1(n4857), .B2(n7613), .C1(
        n7612), .C2(n9491), .ZN(P2_U3338) );
  INV_X1 U8827 ( .A(n8750), .ZN(n7614) );
  INV_X1 U8828 ( .A(n8809), .ZN(n8747) );
  XNOR2_X1 U8829 ( .A(n7691), .B(n8910), .ZN(n7617) );
  AOI21_X1 U8830 ( .B1(n7617), .B2(n9349), .A(n7616), .ZN(n10662) );
  INV_X1 U8831 ( .A(n8910), .ZN(n7620) );
  NAND2_X1 U8832 ( .A1(n7621), .A2(n7620), .ZN(n7695) );
  OR2_X1 U8833 ( .A1(n7621), .A2(n7620), .ZN(n7622) );
  AND2_X1 U8834 ( .A1(n7695), .A2(n7622), .ZN(n10661) );
  XNOR2_X1 U8835 ( .A(n7698), .B(n7693), .ZN(n7623) );
  NAND2_X1 U8836 ( .A1(n7623), .A2(n5299), .ZN(n10658) );
  OAI22_X1 U8837 ( .A1(n9378), .A2(n6860), .B1(n7624), .B2(n9316), .ZN(n7625)
         );
  AOI21_X1 U8838 ( .B1(n7693), .B2(n9366), .A(n7625), .ZN(n7626) );
  OAI21_X1 U8839 ( .B1(n10658), .B2(n8093), .A(n7626), .ZN(n7627) );
  AOI21_X1 U8840 ( .B1(n10661), .B2(n9289), .A(n7627), .ZN(n7628) );
  OAI21_X1 U8841 ( .B1(n9268), .B2(n10662), .A(n7628), .ZN(P2_U3285) );
  INV_X1 U8842 ( .A(P2_DATAO_REG_21__SCAN_IN), .ZN(n8180) );
  OAI222_X1 U8843 ( .A1(n10043), .A2(n8179), .B1(P1_U3084), .B2(n4855), .C1(
        n8180), .C2(n10039), .ZN(P1_U3332) );
  NOR3_X1 U8844 ( .A1(n7632), .A2(n7629), .A3(n9017), .ZN(n7630) );
  NOR2_X1 U8845 ( .A1(n7630), .A2(n10282), .ZN(n7639) );
  OAI21_X1 U8846 ( .B1(n7542), .B2(n7632), .A(n7631), .ZN(n7633) );
  NAND2_X1 U8847 ( .A1(n7633), .A2(n9009), .ZN(n7638) );
  NAND2_X1 U8848 ( .A1(n10284), .A2(n7701), .ZN(n7634) );
  OAI211_X1 U8849 ( .C1(n9015), .C2(n7914), .A(n7635), .B(n7634), .ZN(n7636)
         );
  AOI21_X1 U8850 ( .B1(n8805), .B2(n10293), .A(n7636), .ZN(n7637) );
  OAI211_X1 U8851 ( .C1(n7639), .C2(n7694), .A(n7638), .B(n7637), .ZN(P2_U3226) );
  AND2_X1 U8852 ( .A1(n7640), .A2(n10621), .ZN(n7642) );
  NAND2_X1 U8853 ( .A1(n7644), .A2(n7439), .ZN(n7647) );
  AOI22_X1 U8854 ( .A1(n8153), .A2(P2_DATAO_REG_10__SCAN_IN), .B1(n5192), .B2(
        n7645), .ZN(n7646) );
  OR2_X1 U8855 ( .A1(n10641), .A2(n7767), .ZN(n8473) );
  NAND2_X1 U8856 ( .A1(n10641), .A2(n7767), .ZN(n8474) );
  NAND2_X1 U8857 ( .A1(n8473), .A2(n8474), .ZN(n10619) );
  NAND2_X1 U8858 ( .A1(n10614), .A2(n10619), .ZN(n7649) );
  INV_X1 U8859 ( .A(n7767), .ZN(n9622) );
  OR2_X1 U8860 ( .A1(n10641), .A2(n9622), .ZN(n7648) );
  NAND2_X1 U8861 ( .A1(n7649), .A2(n7648), .ZN(n7726) );
  AOI22_X1 U8862 ( .A1(n8153), .A2(P2_DATAO_REG_11__SCAN_IN), .B1(n5192), .B2(
        n7651), .ZN(n7652) );
  AND2_X1 U8863 ( .A1(n7655), .A2(n7654), .ZN(n7656) );
  NOR2_X1 U8864 ( .A1(n7664), .A2(n7656), .ZN(n7769) );
  NAND2_X1 U8865 ( .A1(n4856), .A2(n7769), .ZN(n7662) );
  NAND2_X1 U8866 ( .A1(n6774), .A2(P1_REG1_REG_11__SCAN_IN), .ZN(n7661) );
  OR2_X1 U8867 ( .A1(n8268), .A2(n7657), .ZN(n7660) );
  INV_X1 U8868 ( .A(P1_REG0_REG_11__SCAN_IN), .ZN(n7658) );
  OR2_X1 U8869 ( .A1(n8270), .A2(n7658), .ZN(n7659) );
  OR2_X1 U8870 ( .A1(n10003), .A2(n7760), .ZN(n8478) );
  NAND2_X1 U8871 ( .A1(n10003), .A2(n7760), .ZN(n8479) );
  XNOR2_X1 U8872 ( .A(n7726), .B(n8369), .ZN(n10002) );
  INV_X1 U8873 ( .A(n10619), .ZN(n7663) );
  XNOR2_X1 U8874 ( .A(n7748), .B(n8369), .ZN(n7672) );
  OR2_X1 U8875 ( .A1(n7664), .A2(P1_REG3_REG_12__SCAN_IN), .ZN(n7665) );
  AND2_X1 U8876 ( .A1(n7665), .A2(n7740), .ZN(n7802) );
  NAND2_X1 U8877 ( .A1(n4856), .A2(n7802), .ZN(n7670) );
  NAND2_X1 U8878 ( .A1(n6774), .A2(P1_REG1_REG_12__SCAN_IN), .ZN(n7669) );
  OR2_X1 U8879 ( .A1(n8268), .A2(n6345), .ZN(n7668) );
  INV_X1 U8880 ( .A(P1_REG0_REG_12__SCAN_IN), .ZN(n7666) );
  OR2_X1 U8881 ( .A1(n8270), .A2(n7666), .ZN(n7667) );
  AOI22_X1 U8882 ( .A1(n10622), .A2(n9622), .B1(n9621), .B2(n10623), .ZN(n7671) );
  OAI21_X1 U8883 ( .B1(n7672), .B2(n10626), .A(n7671), .ZN(n7673) );
  AOI21_X1 U8884 ( .B1(n10002), .B2(n10629), .A(n7673), .ZN(n10006) );
  INV_X1 U8885 ( .A(n10003), .ZN(n7772) );
  INV_X1 U8886 ( .A(n7733), .ZN(n7674) );
  AOI21_X1 U8887 ( .B1(n10003), .B2(n10616), .A(n7674), .ZN(n10004) );
  NAND2_X1 U8888 ( .A1(n10004), .A2(n9902), .ZN(n7676) );
  AOI22_X1 U8889 ( .A1(n9896), .A2(P1_REG2_REG_11__SCAN_IN), .B1(n7769), .B2(
        n10638), .ZN(n7675) );
  OAI211_X1 U8890 ( .C1(n7772), .C2(n9898), .A(n7676), .B(n7675), .ZN(n7677)
         );
  AOI21_X1 U8891 ( .B1(n10002), .B2(n10645), .A(n7677), .ZN(n7678) );
  OAI21_X1 U8892 ( .B1(n10006), .B2(n9896), .A(n7678), .ZN(P1_U3280) );
  OAI21_X1 U8893 ( .B1(n7680), .B2(P2_REG2_REG_14__SCAN_IN), .A(n7679), .ZN(
        n7819) );
  XNOR2_X1 U8894 ( .A(n7819), .B(n7810), .ZN(n7682) );
  INV_X1 U8895 ( .A(P2_REG2_REG_15__SCAN_IN), .ZN(n7681) );
  NAND2_X1 U8896 ( .A1(n7682), .A2(n7681), .ZN(n7821) );
  OAI21_X1 U8897 ( .B1(n7682), .B2(n7681), .A(n7821), .ZN(n7683) );
  INV_X1 U8898 ( .A(n7683), .ZN(n7690) );
  AOI21_X1 U8899 ( .B1(n7685), .B2(n10688), .A(n7684), .ZN(n7809) );
  XNOR2_X1 U8900 ( .A(n7809), .B(n7820), .ZN(n7686) );
  NAND2_X1 U8901 ( .A1(P2_REG1_REG_15__SCAN_IN), .A2(n7686), .ZN(n7811) );
  OAI211_X1 U8902 ( .C1(n7686), .C2(P2_REG1_REG_15__SCAN_IN), .A(n10450), .B(
        n7811), .ZN(n7689) );
  AND2_X1 U8903 ( .A1(P2_REG3_REG_15__SCAN_IN), .A2(P2_U3152), .ZN(n8305) );
  NOR2_X1 U8904 ( .A1(n10414), .A2(n7820), .ZN(n7687) );
  AOI211_X1 U8905 ( .C1(P2_ADDR_REG_15__SCAN_IN), .C2(n10486), .A(n8305), .B(
        n7687), .ZN(n7688) );
  OAI211_X1 U8906 ( .C1(n7690), .C2(n10415), .A(n7689), .B(n7688), .ZN(
        P2_U3260) );
  OR2_X1 U8907 ( .A1(n8805), .A2(n8804), .ZN(n8810) );
  NAND2_X1 U8908 ( .A1(n8805), .A2(n8804), .ZN(n8811) );
  XNOR2_X1 U8909 ( .A(n7833), .B(n8801), .ZN(n7692) );
  OAI222_X1 U8910 ( .A1(n9370), .A2(n7914), .B1(n9371), .B2(n7694), .C1(n9376), 
        .C2(n7692), .ZN(n10668) );
  INV_X1 U8911 ( .A(n10668), .ZN(n7706) );
  INV_X1 U8912 ( .A(n7693), .ZN(n10659) );
  NAND2_X1 U8913 ( .A1(n7695), .A2(n5484), .ZN(n7696) );
  NOR2_X1 U8914 ( .A1(n7696), .A2(n8801), .ZN(n7842) );
  AOI21_X1 U8915 ( .B1(n8801), .B2(n7696), .A(n7842), .ZN(n7697) );
  INV_X1 U8916 ( .A(n7697), .ZN(n10669) );
  NAND2_X1 U8917 ( .A1(n8805), .A2(n7699), .ZN(n7700) );
  NAND2_X1 U8918 ( .A1(n7836), .A2(n7700), .ZN(n10666) );
  AOI22_X1 U8919 ( .A1(n9268), .A2(P2_REG2_REG_12__SCAN_IN), .B1(n7701), .B2(
        n9377), .ZN(n7703) );
  NAND2_X1 U8920 ( .A1(n8805), .A2(n9366), .ZN(n7702) );
  OAI211_X1 U8921 ( .C1(n10666), .C2(n9152), .A(n7703), .B(n7702), .ZN(n7704)
         );
  AOI21_X1 U8922 ( .B1(n10669), .B2(n9289), .A(n7704), .ZN(n7705) );
  OAI21_X1 U8923 ( .B1(n9268), .B2(n7706), .A(n7705), .ZN(P2_U3284) );
  NAND2_X1 U8924 ( .A1(n7708), .A2(n7707), .ZN(n7709) );
  NAND2_X1 U8925 ( .A1(n10641), .A2(n8672), .ZN(n7712) );
  NAND2_X1 U8926 ( .A1(n9622), .A2(n8678), .ZN(n7711) );
  NAND2_X1 U8927 ( .A1(n7712), .A2(n7711), .ZN(n7713) );
  XNOR2_X1 U8928 ( .A(n7713), .B(n8683), .ZN(n7715) );
  NAND2_X1 U8929 ( .A1(n7714), .A2(n7715), .ZN(n7755) );
  INV_X1 U8930 ( .A(n7714), .ZN(n7717) );
  INV_X1 U8931 ( .A(n7715), .ZN(n7716) );
  NAND2_X1 U8932 ( .A1(n7755), .A2(n7756), .ZN(n7719) );
  NOR2_X1 U8933 ( .A1(n7767), .A2(n8682), .ZN(n7718) );
  AOI21_X1 U8934 ( .B1(n10641), .B2(n8678), .A(n7718), .ZN(n7754) );
  XNOR2_X1 U8935 ( .A(n7719), .B(n7754), .ZN(n7725) );
  AOI21_X1 U8936 ( .B1(n9566), .B2(n10621), .A(n7720), .ZN(n7722) );
  NAND2_X1 U8937 ( .A1(n9602), .A2(n10639), .ZN(n7721) );
  OAI211_X1 U8938 ( .C1(n7760), .C2(n9569), .A(n7722), .B(n7721), .ZN(n7723)
         );
  AOI21_X1 U8939 ( .B1(n10641), .B2(n9607), .A(n7723), .ZN(n7724) );
  OAI21_X1 U8940 ( .B1(n7725), .B2(n9609), .A(n7724), .ZN(P1_U3215) );
  NAND2_X1 U8941 ( .A1(n7726), .A2(n8369), .ZN(n7728) );
  INV_X1 U8942 ( .A(n7760), .ZN(n10624) );
  OR2_X1 U8943 ( .A1(n10003), .A2(n10624), .ZN(n7727) );
  NAND2_X1 U8944 ( .A1(n7729), .A2(n7439), .ZN(n7732) );
  AOI22_X1 U8945 ( .A1(n8153), .A2(P2_DATAO_REG_12__SCAN_IN), .B1(n5192), .B2(
        n7730), .ZN(n7731) );
  OR2_X1 U8946 ( .A1(n9998), .A2(n7959), .ZN(n8485) );
  NAND2_X1 U8947 ( .A1(n9998), .A2(n7959), .ZN(n8486) );
  NAND2_X1 U8948 ( .A1(n8485), .A2(n8486), .ZN(n8482) );
  INV_X1 U8949 ( .A(n8482), .ZN(n7749) );
  OAI21_X1 U8950 ( .B1(n4941), .B2(n8482), .A(n7850), .ZN(n10000) );
  NAND2_X1 U8951 ( .A1(n9998), .A2(n7733), .ZN(n7734) );
  NAND2_X1 U8952 ( .A1(n7734), .A2(n10617), .ZN(n7735) );
  NOR2_X1 U8953 ( .A1(n7931), .A2(n7735), .ZN(n9997) );
  NAND2_X1 U8954 ( .A1(n9998), .A2(n10640), .ZN(n7737) );
  AOI22_X1 U8955 ( .A1(n9896), .A2(P1_REG2_REG_12__SCAN_IN), .B1(n7802), .B2(
        n10638), .ZN(n7736) );
  NAND2_X1 U8956 ( .A1(n7737), .A2(n7736), .ZN(n7738) );
  AOI21_X1 U8957 ( .B1(n9997), .B2(n10644), .A(n7738), .ZN(n7753) );
  NAND2_X1 U8958 ( .A1(n7740), .A2(n7739), .ZN(n7741) );
  AND2_X1 U8959 ( .A1(n7862), .A2(n7741), .ZN(n7961) );
  NAND2_X1 U8960 ( .A1(n4856), .A2(n7961), .ZN(n7747) );
  NAND2_X1 U8961 ( .A1(n6774), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n7746) );
  INV_X1 U8962 ( .A(P1_REG0_REG_13__SCAN_IN), .ZN(n7742) );
  OR2_X1 U8963 ( .A1(n8270), .A2(n7742), .ZN(n7745) );
  INV_X1 U8964 ( .A(P1_REG2_REG_13__SCAN_IN), .ZN(n7743) );
  OR2_X1 U8965 ( .A1(n8268), .A2(n7743), .ZN(n7744) );
  NAND2_X1 U8966 ( .A1(n7871), .A2(n8478), .ZN(n7750) );
  XNOR2_X1 U8967 ( .A(n7750), .B(n7749), .ZN(n7751) );
  OAI222_X1 U8968 ( .A1(n9881), .A2(n7855), .B1(n9879), .B2(n7760), .C1(n10626), .C2(n7751), .ZN(n9996) );
  NAND2_X1 U8969 ( .A1(n9996), .A2(n9841), .ZN(n7752) );
  OAI211_X1 U8970 ( .C1(n10000), .C2(n9853), .A(n7753), .B(n7752), .ZN(
        P1_U3279) );
  NAND2_X1 U8971 ( .A1(n10003), .A2(n6773), .ZN(n7758) );
  NAND2_X1 U8972 ( .A1(n10624), .A2(n8678), .ZN(n7757) );
  NAND2_X1 U8973 ( .A1(n7758), .A2(n7757), .ZN(n7759) );
  XNOR2_X1 U8974 ( .A(n7759), .B(n8675), .ZN(n7789) );
  NOR2_X1 U8975 ( .A1(n7760), .A2(n8682), .ZN(n7761) );
  AOI21_X1 U8976 ( .B1(n10003), .B2(n8678), .A(n7761), .ZN(n7790) );
  XNOR2_X1 U8977 ( .A(n7789), .B(n7790), .ZN(n7763) );
  AOI21_X1 U8978 ( .B1(n7762), .B2(n7763), .A(n9609), .ZN(n7764) );
  NAND2_X1 U8979 ( .A1(n7764), .A2(n7794), .ZN(n7771) );
  AOI21_X1 U8980 ( .B1(n9601), .B2(n9621), .A(n7765), .ZN(n7766) );
  OAI21_X1 U8981 ( .B1(n9605), .B2(n7767), .A(n7766), .ZN(n7768) );
  AOI21_X1 U8982 ( .B1(n7769), .B2(n9602), .A(n7768), .ZN(n7770) );
  OAI211_X1 U8983 ( .C1(n7772), .C2(n9598), .A(n7771), .B(n7770), .ZN(P1_U3234) );
  INV_X1 U8984 ( .A(P1_ADDR_REG_15__SCAN_IN), .ZN(n7776) );
  OAI211_X1 U8985 ( .C1(P1_REG1_REG_15__SCAN_IN), .C2(n7774), .A(n10398), .B(
        n7773), .ZN(n7775) );
  NAND2_X1 U8986 ( .A1(P1_U3084), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n8125) );
  OAI211_X1 U8987 ( .C1(n7776), .C2(n10391), .A(n7775), .B(n8125), .ZN(n7781)
         );
  AOI211_X1 U8988 ( .C1(n7779), .C2(n7778), .A(n7777), .B(n9673), .ZN(n7780)
         );
  AOI211_X1 U8989 ( .C1(n9678), .C2(n8007), .A(n7781), .B(n7780), .ZN(n7782)
         );
  INV_X1 U8990 ( .A(n7782), .ZN(P1_U3256) );
  INV_X1 U8991 ( .A(P2_DATAO_REG_23__SCAN_IN), .ZN(n8209) );
  NAND2_X1 U8992 ( .A1(n8208), .A2(n7783), .ZN(n7785) );
  NAND2_X1 U8993 ( .A1(n7784), .A2(P1_STATE_REG_SCAN_IN), .ZN(n8601) );
  OAI211_X1 U8994 ( .C1(n8209), .C2(n10039), .A(n7785), .B(n8601), .ZN(
        P1_U3330) );
  NAND2_X1 U8995 ( .A1(n8208), .A2(n7786), .ZN(n7787) );
  OAI211_X1 U8996 ( .C1(n7788), .C2(n9491), .A(n7787), .B(n8935), .ZN(P2_U3335) );
  INV_X1 U8997 ( .A(n7789), .ZN(n7792) );
  INV_X1 U8998 ( .A(n7790), .ZN(n7791) );
  NAND2_X1 U8999 ( .A1(n7792), .A2(n7791), .ZN(n7793) );
  NAND2_X1 U9000 ( .A1(n9998), .A2(n8672), .ZN(n7796) );
  NAND2_X1 U9001 ( .A1(n9621), .A2(n8678), .ZN(n7795) );
  NAND2_X1 U9002 ( .A1(n7796), .A2(n7795), .ZN(n7797) );
  XNOR2_X1 U9003 ( .A(n7797), .B(n8683), .ZN(n7940) );
  NAND2_X1 U9004 ( .A1(n9998), .A2(n8678), .ZN(n7799) );
  NAND2_X1 U9005 ( .A1(n9621), .A2(n6799), .ZN(n7798) );
  NAND2_X1 U9006 ( .A1(n7799), .A2(n7798), .ZN(n7939) );
  INV_X1 U9007 ( .A(n7939), .ZN(n7937) );
  XNOR2_X1 U9008 ( .A(n7940), .B(n7937), .ZN(n7800) );
  XNOR2_X1 U9009 ( .A(n7942), .B(n7800), .ZN(n7807) );
  AOI21_X1 U9010 ( .B1(n9566), .B2(n10624), .A(n7801), .ZN(n7804) );
  NAND2_X1 U9011 ( .A1(n9602), .A2(n7802), .ZN(n7803) );
  OAI211_X1 U9012 ( .C1(n7855), .C2(n9569), .A(n7804), .B(n7803), .ZN(n7805)
         );
  AOI21_X1 U9013 ( .B1(n9998), .B2(n9607), .A(n7805), .ZN(n7806) );
  OAI21_X1 U9014 ( .B1(n7807), .B2(n9609), .A(n7806), .ZN(P1_U3222) );
  INV_X1 U9015 ( .A(P2_DATAO_REG_24__SCAN_IN), .ZN(n8213) );
  OAI222_X1 U9016 ( .A1(n10043), .A2(n8212), .B1(P1_U3084), .B2(n7808), .C1(
        n8213), .C2(n10039), .ZN(P1_U3329) );
  NAND2_X1 U9017 ( .A1(n7810), .A2(n7809), .ZN(n7812) );
  NAND2_X1 U9018 ( .A1(n7812), .A2(n7811), .ZN(n7815) );
  INV_X1 U9019 ( .A(P2_REG1_REG_16__SCAN_IN), .ZN(n7813) );
  NAND2_X1 U9020 ( .A1(n7827), .A2(n7813), .ZN(n7968) );
  OAI21_X1 U9021 ( .B1(n7827), .B2(n7813), .A(n7968), .ZN(n7814) );
  NAND2_X1 U9022 ( .A1(n7815), .A2(n7814), .ZN(n7816) );
  AOI21_X1 U9023 ( .B1(n7969), .B2(n7816), .A(n10481), .ZN(n7830) );
  INV_X1 U9024 ( .A(P2_REG2_REG_16__SCAN_IN), .ZN(n7818) );
  NOR2_X1 U9025 ( .A1(n7973), .A2(n7818), .ZN(n7817) );
  AOI21_X1 U9026 ( .B1(n7973), .B2(n7818), .A(n7817), .ZN(n7824) );
  NAND2_X1 U9027 ( .A1(n7820), .A2(n7819), .ZN(n7822) );
  NAND2_X1 U9028 ( .A1(n7822), .A2(n7821), .ZN(n7823) );
  NOR2_X1 U9029 ( .A1(n7823), .A2(n7824), .ZN(n7972) );
  AOI211_X1 U9030 ( .C1(n7824), .C2(n7823), .A(n10415), .B(n7972), .ZN(n7829)
         );
  NOR2_X1 U9031 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n10248), .ZN(n7825) );
  AOI21_X1 U9032 ( .B1(n10486), .B2(P2_ADDR_REG_16__SCAN_IN), .A(n7825), .ZN(
        n7826) );
  OAI21_X1 U9033 ( .B1(n10414), .B2(n7827), .A(n7826), .ZN(n7828) );
  OR3_X1 U9034 ( .A1(n7830), .A2(n7829), .A3(n7828), .ZN(P2_U3261) );
  OAI222_X1 U9035 ( .A1(n7832), .A2(P2_U3152), .B1(n4857), .B2(n8212), .C1(
        n7831), .C2(n9491), .ZN(P2_U3334) );
  INV_X1 U9036 ( .A(n8801), .ZN(n8913) );
  NAND2_X1 U9037 ( .A1(n7834), .A2(n8811), .ZN(n7910) );
  OR2_X1 U9038 ( .A1(n10294), .A2(n7914), .ZN(n8818) );
  NAND2_X1 U9039 ( .A1(n10294), .A2(n7914), .ZN(n8819) );
  XNOR2_X1 U9040 ( .A(n7910), .B(n7843), .ZN(n7835) );
  OAI222_X1 U9041 ( .A1(n9370), .A2(n9060), .B1(n7835), .B2(n9376), .C1(n9371), 
        .C2(n8804), .ZN(n10677) );
  INV_X1 U9042 ( .A(n7836), .ZN(n7837) );
  OAI21_X1 U9043 ( .B1(n5203), .B2(n7837), .A(n4930), .ZN(n10675) );
  AOI22_X1 U9044 ( .A1(n9268), .A2(P2_REG2_REG_13__SCAN_IN), .B1(n10283), .B2(
        n9377), .ZN(n7839) );
  NAND2_X1 U9045 ( .A1(n10294), .A2(n9366), .ZN(n7838) );
  OAI211_X1 U9046 ( .C1(n10675), .C2(n9152), .A(n7839), .B(n7838), .ZN(n7847)
         );
  NOR2_X1 U9047 ( .A1(n7844), .A2(n7843), .ZN(n10674) );
  INV_X1 U9048 ( .A(n10678), .ZN(n7845) );
  NOR3_X1 U9049 ( .A1(n10674), .A2(n7845), .A3(n9359), .ZN(n7846) );
  AOI211_X1 U9050 ( .C1(n9378), .C2(n10677), .A(n7847), .B(n7846), .ZN(n7848)
         );
  INV_X1 U9051 ( .A(n7848), .ZN(P2_U3283) );
  NAND2_X1 U9052 ( .A1(n9998), .A2(n9621), .ZN(n7849) );
  NAND2_X1 U9053 ( .A1(n7851), .A2(n7439), .ZN(n7854) );
  AOI22_X1 U9054 ( .A1(n8153), .A2(P2_DATAO_REG_13__SCAN_IN), .B1(n7852), .B2(
        n5192), .ZN(n7853) );
  INV_X1 U9055 ( .A(n8493), .ZN(n8422) );
  INV_X1 U9056 ( .A(n8495), .ZN(n8419) );
  INV_X1 U9057 ( .A(n8371), .ZN(n7856) );
  AOI22_X1 U9058 ( .A1(n8153), .A2(P2_DATAO_REG_14__SCAN_IN), .B1(n5192), .B2(
        n7858), .ZN(n7859) );
  AND2_X1 U9059 ( .A1(n7862), .A2(n7861), .ZN(n7863) );
  NOR2_X1 U9060 ( .A1(n7875), .A2(n7863), .ZN(n8074) );
  NAND2_X1 U9061 ( .A1(n4856), .A2(n8074), .ZN(n7869) );
  NAND2_X1 U9062 ( .A1(n6774), .A2(P1_REG1_REG_14__SCAN_IN), .ZN(n7868) );
  INV_X1 U9063 ( .A(P1_REG2_REG_14__SCAN_IN), .ZN(n7864) );
  OR2_X1 U9064 ( .A1(n8268), .A2(n7864), .ZN(n7867) );
  INV_X1 U9065 ( .A(P1_REG0_REG_14__SCAN_IN), .ZN(n7865) );
  OR2_X1 U9066 ( .A1(n8270), .A2(n7865), .ZN(n7866) );
  NAND2_X1 U9067 ( .A1(n9993), .A2(n8126), .ZN(n8494) );
  NAND2_X1 U9068 ( .A1(n8496), .A2(n8494), .ZN(n8491) );
  INV_X1 U9069 ( .A(n8491), .ZN(n8372) );
  XNOR2_X1 U9070 ( .A(n8004), .B(n8372), .ZN(n9995) );
  NAND2_X1 U9071 ( .A1(n8485), .A2(n8478), .ZN(n8421) );
  INV_X1 U9072 ( .A(n8421), .ZN(n7870) );
  NAND2_X1 U9073 ( .A1(n7871), .A2(n7870), .ZN(n7872) );
  NAND2_X1 U9074 ( .A1(n7872), .A2(n8486), .ZN(n7925) );
  OAI21_X1 U9075 ( .B1(n7873), .B2(n8495), .A(n8491), .ZN(n7874) );
  NAND3_X1 U9076 ( .A1(n7874), .A2(n8012), .A3(n9891), .ZN(n7882) );
  NOR2_X1 U9077 ( .A1(n7875), .A2(P1_REG3_REG_15__SCAN_IN), .ZN(n7876) );
  OR2_X1 U9078 ( .A1(n8014), .A2(n7876), .ZN(n8129) );
  INV_X1 U9079 ( .A(n4856), .ZN(n8160) );
  OAI22_X1 U9080 ( .A1(n8129), .A2(n8160), .B1(n8268), .B2(n7778), .ZN(n7880)
         );
  INV_X1 U9081 ( .A(P1_REG1_REG_15__SCAN_IN), .ZN(n7878) );
  NAND2_X1 U9082 ( .A1(n5475), .A2(P1_REG0_REG_15__SCAN_IN), .ZN(n7877) );
  OAI21_X1 U9083 ( .B1(n8341), .B2(n7878), .A(n7877), .ZN(n7879) );
  AOI22_X1 U9084 ( .A1(n9620), .A2(n10622), .B1(n10623), .B2(n9618), .ZN(n7881) );
  NAND2_X1 U9085 ( .A1(n7882), .A2(n7881), .ZN(n9992) );
  INV_X1 U9086 ( .A(n9993), .ZN(n7885) );
  NAND2_X1 U9087 ( .A1(n8032), .A2(n7931), .ZN(n7930) );
  AOI211_X1 U9088 ( .C1(n9993), .C2(n7930), .A(n10597), .B(n5196), .ZN(n9991)
         );
  NAND2_X1 U9089 ( .A1(n9991), .A2(n10644), .ZN(n7884) );
  AOI22_X1 U9090 ( .A1(n9896), .A2(P1_REG2_REG_14__SCAN_IN), .B1(n8074), .B2(
        n10638), .ZN(n7883) );
  OAI211_X1 U9091 ( .C1(n7885), .C2(n9898), .A(n7884), .B(n7883), .ZN(n7886)
         );
  AOI21_X1 U9092 ( .B1(n9841), .B2(n9992), .A(n7886), .ZN(n7887) );
  OAI21_X1 U9093 ( .B1(n9995), .B2(n9853), .A(n7887), .ZN(P1_U3277) );
  INV_X1 U9094 ( .A(n7888), .ZN(n8090) );
  NOR2_X1 U9095 ( .A1(n9044), .A2(n8090), .ZN(n7890) );
  INV_X1 U9096 ( .A(n9338), .ZN(n9127) );
  INV_X1 U9097 ( .A(n7982), .ZN(n9059) );
  AOI22_X1 U9098 ( .A1(n9127), .A2(n9241), .B1(n9059), .B2(n9239), .ZN(n8085)
         );
  OAI22_X1 U9099 ( .A1(n8994), .A2(n8085), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10248), .ZN(n7889) );
  AOI211_X1 U9100 ( .C1(n9124), .C2(n10293), .A(n7890), .B(n7889), .ZN(n7895)
         );
  OAI22_X1 U9101 ( .A1(n7892), .A2(n10288), .B1(n7982), .B2(n9017), .ZN(n7893)
         );
  NAND3_X1 U9102 ( .A1(n4958), .A2(n8315), .A3(n7893), .ZN(n7894) );
  OAI211_X1 U9103 ( .C1(n7896), .C2(n10288), .A(n7895), .B(n7894), .ZN(
        P2_U3228) );
  INV_X1 U9104 ( .A(n7897), .ZN(n10287) );
  NOR3_X1 U9105 ( .A1(n7898), .A2(n7914), .A3(n9017), .ZN(n7899) );
  AOI21_X1 U9106 ( .B1(n10287), .B2(n9009), .A(n7899), .ZN(n7908) );
  INV_X1 U9107 ( .A(n7917), .ZN(n7902) );
  INV_X1 U9108 ( .A(n7914), .ZN(n9061) );
  AOI22_X1 U9109 ( .A1(n10282), .A2(n9061), .B1(n10281), .B2(n9059), .ZN(n7901) );
  OAI211_X1 U9110 ( .C1(n9044), .C2(n7902), .A(n7901), .B(n7900), .ZN(n7905)
         );
  NOR2_X1 U9111 ( .A1(n7903), .A2(n10288), .ZN(n7904) );
  AOI211_X1 U9112 ( .C1(n7985), .C2(n10293), .A(n7905), .B(n7904), .ZN(n7906)
         );
  OAI21_X1 U9113 ( .B1(n7908), .B2(n7907), .A(n7906), .ZN(P2_U3217) );
  INV_X1 U9114 ( .A(n8819), .ZN(n7909) );
  NAND2_X1 U9115 ( .A1(n7985), .A2(n9060), .ZN(n8822) );
  NAND2_X1 U9116 ( .A1(n7911), .A2(n8821), .ZN(n7983) );
  OAI211_X1 U9117 ( .C1(n7911), .C2(n8821), .A(n9349), .B(n7983), .ZN(n7913)
         );
  NAND2_X1 U9118 ( .A1(n9059), .A2(n9241), .ZN(n7912) );
  OAI211_X1 U9119 ( .C1(n7914), .C2(n9371), .A(n7913), .B(n7912), .ZN(n10686)
         );
  INV_X1 U9120 ( .A(n10686), .ZN(n7922) );
  AOI21_X1 U9121 ( .B1(n8821), .B2(n7915), .A(n4934), .ZN(n7916) );
  INV_X1 U9122 ( .A(n7916), .ZN(n10687) );
  XNOR2_X1 U9123 ( .A(n7985), .B(n4930), .ZN(n10684) );
  AOI22_X1 U9124 ( .A1(n9268), .A2(P2_REG2_REG_14__SCAN_IN), .B1(n7917), .B2(
        n9377), .ZN(n7919) );
  NAND2_X1 U9125 ( .A1(n7985), .A2(n9366), .ZN(n7918) );
  OAI211_X1 U9126 ( .C1(n10684), .C2(n9152), .A(n7919), .B(n7918), .ZN(n7920)
         );
  AOI21_X1 U9127 ( .B1(n10687), .B2(n9289), .A(n7920), .ZN(n7921) );
  OAI21_X1 U9128 ( .B1(n9268), .B2(n7922), .A(n7921), .ZN(P2_U3282) );
  AOI21_X1 U9129 ( .B1(n8371), .B2(n7923), .A(n4935), .ZN(n7929) );
  OAI21_X1 U9130 ( .B1(n8371), .B2(n7925), .A(n7924), .ZN(n7927) );
  OAI22_X1 U9131 ( .A1(n8126), .A2(n9881), .B1(n7959), .B2(n9879), .ZN(n7926)
         );
  AOI21_X1 U9132 ( .B1(n7927), .B2(n9891), .A(n7926), .ZN(n7928) );
  OAI21_X1 U9133 ( .B1(n7929), .B2(n9887), .A(n7928), .ZN(n8034) );
  INV_X1 U9134 ( .A(n8034), .ZN(n7936) );
  INV_X1 U9135 ( .A(n7929), .ZN(n8036) );
  OAI21_X1 U9136 ( .B1(n8032), .B2(n7931), .A(n7930), .ZN(n8033) );
  AOI22_X1 U9137 ( .A1(n9896), .A2(P1_REG2_REG_13__SCAN_IN), .B1(n7961), .B2(
        n10638), .ZN(n7933) );
  NAND2_X1 U9138 ( .A1(n7946), .A2(n10640), .ZN(n7932) );
  OAI211_X1 U9139 ( .C1(n8033), .C2(n9870), .A(n7933), .B(n7932), .ZN(n7934)
         );
  AOI21_X1 U9140 ( .B1(n8036), .B2(n10645), .A(n7934), .ZN(n7935) );
  OAI21_X1 U9141 ( .B1(n7936), .B2(n9896), .A(n7935), .ZN(P1_U3278) );
  INV_X1 U9142 ( .A(n7940), .ZN(n7938) );
  NAND2_X1 U9143 ( .A1(n7938), .A2(n7937), .ZN(n7941) );
  NAND2_X1 U9144 ( .A1(n7946), .A2(n6773), .ZN(n7944) );
  NAND2_X1 U9145 ( .A1(n9620), .A2(n8678), .ZN(n7943) );
  NAND2_X1 U9146 ( .A1(n7944), .A2(n7943), .ZN(n7945) );
  XNOR2_X1 U9147 ( .A(n7945), .B(n8683), .ZN(n7949) );
  NAND2_X1 U9148 ( .A1(n7946), .A2(n8678), .ZN(n7948) );
  NAND2_X1 U9149 ( .A1(n9620), .A2(n6799), .ZN(n7947) );
  NAND2_X1 U9150 ( .A1(n7948), .A2(n7947), .ZN(n7950) );
  NAND2_X1 U9151 ( .A1(n7949), .A2(n7950), .ZN(n7954) );
  INV_X1 U9152 ( .A(n7949), .ZN(n7952) );
  INV_X1 U9153 ( .A(n7950), .ZN(n7951) );
  NAND2_X1 U9154 ( .A1(n7952), .A2(n7951), .ZN(n8065) );
  NOR2_X1 U9155 ( .A1(n8066), .A2(n5390), .ZN(n7956) );
  AOI21_X1 U9156 ( .B1(n8065), .B2(n7954), .A(n7953), .ZN(n7955) );
  OAI21_X1 U9157 ( .B1(n7956), .B2(n7955), .A(n9590), .ZN(n7963) );
  INV_X1 U9158 ( .A(n8126), .ZN(n9619) );
  AOI21_X1 U9159 ( .B1(n9601), .B2(n9619), .A(n7957), .ZN(n7958) );
  OAI21_X1 U9160 ( .B1(n9605), .B2(n7959), .A(n7958), .ZN(n7960) );
  AOI21_X1 U9161 ( .B1(n7961), .B2(n9602), .A(n7960), .ZN(n7962) );
  OAI211_X1 U9162 ( .C1(n8032), .C2(n9598), .A(n7963), .B(n7962), .ZN(P1_U3232) );
  INV_X1 U9163 ( .A(P2_DATAO_REG_25__SCAN_IN), .ZN(n8227) );
  INV_X1 U9164 ( .A(n8226), .ZN(n7966) );
  OAI222_X1 U9165 ( .A1(n10039), .A2(n8227), .B1(n10033), .B2(n7966), .C1(
        n7964), .C2(P1_U3084), .ZN(P1_U3328) );
  INV_X1 U9166 ( .A(n10049), .ZN(n7967) );
  OAI222_X1 U9167 ( .A1(P2_U3152), .A2(n7967), .B1(n4857), .B2(n7966), .C1(
        n7965), .C2(n9491), .ZN(P2_U3333) );
  NAND2_X1 U9168 ( .A1(n7969), .A2(n7968), .ZN(n9077) );
  XNOR2_X1 U9169 ( .A(n9081), .B(P2_REG1_REG_17__SCAN_IN), .ZN(n9078) );
  XNOR2_X1 U9170 ( .A(n9077), .B(n9078), .ZN(n7980) );
  NOR2_X1 U9171 ( .A1(P2_STATE_REG_SCAN_IN), .A2(n5911), .ZN(n7970) );
  AOI21_X1 U9172 ( .B1(n10486), .B2(P2_ADDR_REG_17__SCAN_IN), .A(n7970), .ZN(
        n7971) );
  OAI21_X1 U9173 ( .B1(n10414), .B2(n9081), .A(n7971), .ZN(n7979) );
  AOI21_X1 U9174 ( .B1(n7973), .B2(P2_REG2_REG_16__SCAN_IN), .A(n7972), .ZN(
        n7977) );
  INV_X1 U9175 ( .A(P2_REG2_REG_17__SCAN_IN), .ZN(n7975) );
  NOR2_X1 U9176 ( .A1(n9073), .A2(n7975), .ZN(n7974) );
  AOI21_X1 U9177 ( .B1(n9073), .B2(n7975), .A(n7974), .ZN(n7976) );
  NOR2_X1 U9178 ( .A1(n7977), .A2(n7976), .ZN(n9072) );
  AOI211_X1 U9179 ( .C1(n7977), .C2(n7976), .A(n10415), .B(n9072), .ZN(n7978)
         );
  AOI211_X1 U9180 ( .C1(n10450), .C2(n7980), .A(n7979), .B(n7978), .ZN(n7981)
         );
  INV_X1 U9181 ( .A(n7981), .ZN(P2_U3262) );
  INV_X1 U9182 ( .A(n7985), .ZN(n10683) );
  NAND2_X1 U9183 ( .A1(n8310), .A2(n7982), .ZN(n8745) );
  NAND2_X1 U9184 ( .A1(n8744), .A2(n8745), .ZN(n8828) );
  XNOR2_X1 U9185 ( .A(n8087), .B(n8916), .ZN(n10698) );
  INV_X1 U9186 ( .A(n10698), .ZN(n7993) );
  NAND2_X1 U9187 ( .A1(n7983), .A2(n8823), .ZN(n8084) );
  XNOR2_X1 U9188 ( .A(n8084), .B(n8916), .ZN(n7984) );
  OAI222_X1 U9189 ( .A1(n9370), .A2(n9058), .B1(n9371), .B2(n9060), .C1(n9376), 
        .C2(n7984), .ZN(n10696) );
  INV_X1 U9190 ( .A(n8310), .ZN(n10692) );
  INV_X1 U9191 ( .A(n7986), .ZN(n7988) );
  NOR2_X2 U9192 ( .A1(n8310), .A2(n7986), .ZN(n8089) );
  INV_X1 U9193 ( .A(n8089), .ZN(n7987) );
  OAI21_X1 U9194 ( .B1(n10692), .B2(n7988), .A(n7987), .ZN(n10694) );
  AOI22_X1 U9195 ( .A1(n9268), .A2(P2_REG2_REG_15__SCAN_IN), .B1(n8306), .B2(
        n9377), .ZN(n7990) );
  NAND2_X1 U9196 ( .A1(n8310), .A2(n9366), .ZN(n7989) );
  OAI211_X1 U9197 ( .C1(n10694), .C2(n9152), .A(n7990), .B(n7989), .ZN(n7991)
         );
  AOI21_X1 U9198 ( .B1(n10696), .B2(n9378), .A(n7991), .ZN(n7992) );
  OAI21_X1 U9199 ( .B1(n7993), .B2(n9359), .A(n7992), .ZN(P2_U3281) );
  INV_X1 U9200 ( .A(n7994), .ZN(n7996) );
  NAND2_X1 U9201 ( .A1(n7996), .A2(n7995), .ZN(n7997) );
  XNOR2_X1 U9202 ( .A(n7998), .B(n7997), .ZN(n8003) );
  INV_X1 U9203 ( .A(n9353), .ZN(n8000) );
  INV_X1 U9204 ( .A(n9057), .ZN(n9129) );
  OAI22_X1 U9205 ( .A1(n9129), .A2(n9370), .B1(n9058), .B2(n9371), .ZN(n9348)
         );
  AOI22_X1 U9206 ( .A1(n9049), .A2(n9348), .B1(P2_REG3_REG_17__SCAN_IN), .B2(
        P2_U3152), .ZN(n7999) );
  OAI21_X1 U9207 ( .B1(n9044), .B2(n8000), .A(n7999), .ZN(n8001) );
  AOI21_X1 U9208 ( .B1(n9457), .B2(n10293), .A(n8001), .ZN(n8002) );
  OAI21_X1 U9209 ( .B1(n8003), .B2(n10288), .A(n8002), .ZN(P2_U3230) );
  OR2_X1 U9210 ( .A1(n9993), .A2(n9619), .ZN(n8005) );
  NAND2_X1 U9211 ( .A1(n8006), .A2(n7439), .ZN(n8009) );
  AOI22_X1 U9212 ( .A1(n8153), .A2(P2_DATAO_REG_15__SCAN_IN), .B1(n8007), .B2(
        n5192), .ZN(n8008) );
  NAND2_X1 U9213 ( .A1(n9986), .A2(n9538), .ZN(n8503) );
  NAND2_X1 U9214 ( .A1(n8010), .A2(n8500), .ZN(n8011) );
  OAI211_X1 U9215 ( .C1(n8500), .C2(n8013), .A(n8046), .B(n9891), .ZN(n8022)
         );
  OR2_X1 U9216 ( .A1(n8014), .A2(P1_REG3_REG_16__SCAN_IN), .ZN(n8015) );
  AND2_X1 U9217 ( .A1(n8147), .A2(n8015), .ZN(n9540) );
  NAND2_X1 U9218 ( .A1(n9540), .A2(n4856), .ZN(n8020) );
  NAND2_X1 U9219 ( .A1(n5475), .A2(P1_REG0_REG_16__SCAN_IN), .ZN(n8017) );
  NAND2_X1 U9220 ( .A1(n6775), .A2(P1_REG2_REG_16__SCAN_IN), .ZN(n8016) );
  AND2_X1 U9221 ( .A1(n8017), .A2(n8016), .ZN(n8019) );
  NAND2_X1 U9222 ( .A1(n6774), .A2(P1_REG1_REG_16__SCAN_IN), .ZN(n8018) );
  INV_X1 U9223 ( .A(n9880), .ZN(n9617) );
  NAND2_X1 U9224 ( .A1(n9617), .A2(n10623), .ZN(n8021) );
  OAI211_X1 U9225 ( .C1(n8126), .C2(n9879), .A(n8022), .B(n8021), .ZN(n8023)
         );
  AOI21_X1 U9226 ( .B1(n9985), .B2(n10629), .A(n8023), .ZN(n9989) );
  NAND2_X1 U9227 ( .A1(n9986), .A2(n8024), .ZN(n8025) );
  AND2_X1 U9228 ( .A1(n8056), .A2(n8025), .ZN(n9987) );
  NAND2_X1 U9229 ( .A1(n9987), .A2(n9902), .ZN(n8029) );
  NAND2_X1 U9230 ( .A1(n9896), .A2(P1_REG2_REG_15__SCAN_IN), .ZN(n8026) );
  OAI21_X1 U9231 ( .B1(n9866), .B2(n8129), .A(n8026), .ZN(n8027) );
  AOI21_X1 U9232 ( .B1(n9986), .B2(n10640), .A(n8027), .ZN(n8028) );
  NAND2_X1 U9233 ( .A1(n8029), .A2(n8028), .ZN(n8030) );
  AOI21_X1 U9234 ( .B1(n9985), .B2(n10645), .A(n8030), .ZN(n8031) );
  OAI21_X1 U9235 ( .B1(n9989), .B2(n9896), .A(n8031), .ZN(P1_U3276) );
  OAI22_X1 U9236 ( .A1(n8033), .A2(n10597), .B1(n8032), .B2(n10618), .ZN(n8035) );
  AOI211_X1 U9237 ( .C1(n10632), .C2(n8036), .A(n8035), .B(n8034), .ZN(n8039)
         );
  NAND2_X1 U9238 ( .A1(n10633), .A2(P1_REG1_REG_13__SCAN_IN), .ZN(n8037) );
  OAI21_X1 U9239 ( .B1(n8039), .B2(n10633), .A(n8037), .ZN(P1_U3536) );
  NAND2_X1 U9240 ( .A1(n10635), .A2(P1_REG0_REG_13__SCAN_IN), .ZN(n8038) );
  OAI21_X1 U9241 ( .B1(n8039), .B2(n10635), .A(n8038), .ZN(P1_U3493) );
  NAND2_X1 U9242 ( .A1(n9986), .A2(n9618), .ZN(n8040) );
  NAND2_X1 U9243 ( .A1(n8041), .A2(n8040), .ZN(n8045) );
  NAND2_X1 U9244 ( .A1(n8042), .A2(n7439), .ZN(n8044) );
  AOI22_X1 U9245 ( .A1(n9655), .A2(n5192), .B1(n8153), .B2(
        P2_DATAO_REG_16__SCAN_IN), .ZN(n8043) );
  NAND2_X1 U9246 ( .A1(n9532), .A2(n9880), .ZN(n8508) );
  NAND2_X1 U9247 ( .A1(n8045), .A2(n8374), .ZN(n8134) );
  OAI21_X1 U9248 ( .B1(n8045), .B2(n8374), .A(n8134), .ZN(n9978) );
  NAND2_X1 U9249 ( .A1(n8046), .A2(n8502), .ZN(n8047) );
  OAI211_X1 U9250 ( .C1(n8047), .C2(n8506), .A(n8280), .B(n9891), .ZN(n8055)
         );
  XNOR2_X1 U9251 ( .A(n8147), .B(P1_REG3_REG_17__SCAN_IN), .ZN(n9895) );
  NAND2_X1 U9252 ( .A1(n9895), .A2(n4856), .ZN(n8052) );
  INV_X1 U9253 ( .A(P1_REG1_REG_17__SCAN_IN), .ZN(n9663) );
  NAND2_X1 U9254 ( .A1(n6775), .A2(P1_REG2_REG_17__SCAN_IN), .ZN(n8049) );
  NAND2_X1 U9255 ( .A1(n5475), .A2(P1_REG0_REG_17__SCAN_IN), .ZN(n8048) );
  OAI211_X1 U9256 ( .C1(n9663), .C2(n8341), .A(n8049), .B(n8048), .ZN(n8050)
         );
  INV_X1 U9257 ( .A(n8050), .ZN(n8051) );
  OAI22_X1 U9258 ( .A1(n9860), .A2(n9881), .B1(n9538), .B2(n9879), .ZN(n8053)
         );
  INV_X1 U9259 ( .A(n8053), .ZN(n8054) );
  NAND2_X1 U9260 ( .A1(n8055), .A2(n8054), .ZN(n9982) );
  AOI21_X1 U9261 ( .B1(n9532), .B2(n8056), .A(n10597), .ZN(n8057) );
  NAND2_X1 U9262 ( .A1(n8057), .A2(n9894), .ZN(n9979) );
  AOI22_X1 U9263 ( .A1(n9896), .A2(P1_REG2_REG_16__SCAN_IN), .B1(n9540), .B2(
        n10638), .ZN(n8059) );
  NAND2_X1 U9264 ( .A1(n9532), .A2(n10640), .ZN(n8058) );
  OAI211_X1 U9265 ( .C1(n9979), .C2(n8060), .A(n8059), .B(n8058), .ZN(n8061)
         );
  AOI21_X1 U9266 ( .B1(n9982), .B2(n9841), .A(n8061), .ZN(n8062) );
  OAI21_X1 U9267 ( .B1(n9978), .B2(n9853), .A(n8062), .ZN(P1_U3275) );
  INV_X1 U9268 ( .A(n8243), .ZN(n8081) );
  INV_X1 U9269 ( .A(P2_DATAO_REG_26__SCAN_IN), .ZN(n8244) );
  OAI222_X1 U9270 ( .A1(n10043), .A2(n8081), .B1(P1_U3084), .B2(n6394), .C1(
        n8244), .C2(n10039), .ZN(P1_U3327) );
  NAND2_X1 U9271 ( .A1(n9993), .A2(n8678), .ZN(n8064) );
  NAND2_X1 U9272 ( .A1(n9619), .A2(n6799), .ZN(n8063) );
  NAND2_X1 U9273 ( .A1(n8064), .A2(n8063), .ZN(n8109) );
  NAND2_X1 U9274 ( .A1(n9993), .A2(n8672), .ZN(n8068) );
  NAND2_X1 U9275 ( .A1(n9619), .A2(n8678), .ZN(n8067) );
  NAND2_X1 U9276 ( .A1(n8068), .A2(n8067), .ZN(n8069) );
  XNOR2_X1 U9277 ( .A(n8069), .B(n8675), .ZN(n8071) );
  INV_X1 U9278 ( .A(n8071), .ZN(n8070) );
  NAND2_X1 U9279 ( .A1(n8111), .A2(n8110), .ZN(n8072) );
  XOR2_X1 U9280 ( .A(n8109), .B(n8072), .Z(n8079) );
  AOI21_X1 U9281 ( .B1(n9566), .B2(n9620), .A(n8073), .ZN(n8076) );
  NAND2_X1 U9282 ( .A1(n9602), .A2(n8074), .ZN(n8075) );
  OAI211_X1 U9283 ( .C1(n9538), .C2(n9569), .A(n8076), .B(n8075), .ZN(n8077)
         );
  AOI21_X1 U9284 ( .B1(n9993), .B2(n9607), .A(n8077), .ZN(n8078) );
  OAI21_X1 U9285 ( .B1(n8079), .B2(n9609), .A(n8078), .ZN(P1_U3213) );
  INV_X1 U9286 ( .A(n10408), .ZN(n8082) );
  OAI222_X1 U9287 ( .A1(n8082), .A2(P2_U3152), .B1(n4857), .B2(n8081), .C1(
        n8080), .C2(n9491), .ZN(P2_U3332) );
  INV_X1 U9288 ( .A(n8744), .ZN(n8083) );
  NAND2_X1 U9289 ( .A1(n9124), .A2(n9058), .ZN(n8743) );
  XNOR2_X1 U9290 ( .A(n8706), .B(n5060), .ZN(n8086) );
  OAI21_X1 U9291 ( .B1(n8086), .B2(n9376), .A(n8085), .ZN(n9465) );
  INV_X1 U9292 ( .A(n9465), .ZN(n8096) );
  AOI21_X1 U9293 ( .B1(n8830), .B2(n8088), .A(n9126), .ZN(n9466) );
  INV_X1 U9294 ( .A(n9124), .ZN(n9463) );
  OAI211_X1 U9295 ( .C1(n9463), .C2(n8089), .A(n5299), .B(n9351), .ZN(n9462)
         );
  OAI22_X1 U9296 ( .A1(n9378), .A2(n7818), .B1(n8090), .B2(n9316), .ZN(n8091)
         );
  AOI21_X1 U9297 ( .B1(n9124), .B2(n9366), .A(n8091), .ZN(n8092) );
  OAI21_X1 U9298 ( .B1(n9462), .B2(n8093), .A(n8092), .ZN(n8094) );
  AOI21_X1 U9299 ( .B1(n9466), .B2(n9289), .A(n8094), .ZN(n8095) );
  OAI21_X1 U9300 ( .B1(n9268), .B2(n8096), .A(n8095), .ZN(P2_U3280) );
  INV_X1 U9301 ( .A(n8259), .ZN(n8106) );
  INV_X1 U9302 ( .A(P2_DATAO_REG_27__SCAN_IN), .ZN(n8260) );
  OAI222_X1 U9303 ( .A1(n10043), .A2(n8106), .B1(n4860), .B2(P1_U3084), .C1(
        n8260), .C2(n10039), .ZN(P1_U3326) );
  NAND2_X1 U9304 ( .A1(n8098), .A2(n8097), .ZN(n8100) );
  XOR2_X1 U9305 ( .A(n8100), .B(n8099), .Z(n8104) );
  INV_X1 U9306 ( .A(n9339), .ZN(n9056) );
  AOI22_X1 U9307 ( .A1(n10282), .A2(n9127), .B1(n10281), .B2(n9056), .ZN(n8101) );
  NAND2_X1 U9308 ( .A1(P2_U3152), .A2(P2_REG3_REG_18__SCAN_IN), .ZN(n9087) );
  OAI211_X1 U9309 ( .C1(n9044), .C2(n9330), .A(n8101), .B(n9087), .ZN(n8102)
         );
  AOI21_X1 U9310 ( .B1(n9451), .B2(n10293), .A(n8102), .ZN(n8103) );
  OAI21_X1 U9311 ( .B1(n8104), .B2(n10288), .A(n8103), .ZN(P2_U3240) );
  OAI222_X1 U9312 ( .A1(P2_U3152), .A2(n6646), .B1(n4857), .B2(n8106), .C1(
        n8105), .C2(n9491), .ZN(P2_U3331) );
  NAND2_X1 U9313 ( .A1(n9986), .A2(n8678), .ZN(n8108) );
  NAND2_X1 U9314 ( .A1(n9618), .A2(n6799), .ZN(n8107) );
  NAND2_X1 U9315 ( .A1(n8108), .A2(n8107), .ZN(n8124) );
  NAND2_X1 U9316 ( .A1(n8110), .A2(n8109), .ZN(n8112) );
  NAND2_X1 U9317 ( .A1(n9986), .A2(n6773), .ZN(n8114) );
  NAND2_X1 U9318 ( .A1(n9618), .A2(n8678), .ZN(n8113) );
  NAND2_X1 U9319 ( .A1(n8114), .A2(n8113), .ZN(n8115) );
  XNOR2_X1 U9320 ( .A(n8115), .B(n8683), .ZN(n8118) );
  INV_X1 U9321 ( .A(n8118), .ZN(n8116) );
  INV_X1 U9322 ( .A(n8121), .ZN(n8119) );
  NAND2_X1 U9323 ( .A1(n8117), .A2(n8118), .ZN(n8120) );
  NAND2_X1 U9324 ( .A1(n8119), .A2(n8120), .ZN(n8123) );
  AND2_X2 U9325 ( .A1(n8121), .A2(n8120), .ZN(n8610) );
  AOI22_X1 U9326 ( .A1(n8124), .A2(n8123), .B1(n8122), .B2(n9534), .ZN(n8132)
         );
  OAI21_X1 U9327 ( .B1(n9605), .B2(n8126), .A(n8125), .ZN(n8127) );
  AOI21_X1 U9328 ( .B1(n9601), .B2(n9617), .A(n8127), .ZN(n8128) );
  OAI21_X1 U9329 ( .B1(n9593), .B2(n8129), .A(n8128), .ZN(n8130) );
  AOI21_X1 U9330 ( .B1(n9986), .B2(n9607), .A(n8130), .ZN(n8131) );
  OAI21_X1 U9331 ( .B1(n8132), .B2(n9609), .A(n8131), .ZN(P1_U3239) );
  INV_X1 U9332 ( .A(P2_DATAO_REG_22__SCAN_IN), .ZN(n8194) );
  INV_X1 U9333 ( .A(n8193), .ZN(n8317) );
  OAI222_X1 U9334 ( .A1(n10039), .A2(n8194), .B1(n10033), .B2(n8317), .C1(
        n6607), .C2(P1_U3084), .ZN(P1_U3331) );
  NAND2_X1 U9335 ( .A1(n9532), .A2(n9617), .ZN(n8133) );
  OAI22_X1 U9336 ( .A1(n9670), .A2(n6603), .B1(n8136), .B2(n8137), .ZN(n8138)
         );
  INV_X1 U9337 ( .A(n8138), .ZN(n8139) );
  OR2_X1 U9338 ( .A1(n9973), .A2(n9860), .ZN(n8511) );
  NAND2_X1 U9339 ( .A1(n9973), .A2(n9860), .ZN(n8512) );
  INV_X1 U9340 ( .A(n9860), .ZN(n9616) );
  OR2_X1 U9341 ( .A1(n9973), .A2(n9616), .ZN(n8141) );
  AOI22_X1 U9342 ( .A1(n9686), .A2(n5192), .B1(n8153), .B2(
        P2_DATAO_REG_18__SCAN_IN), .ZN(n8143) );
  INV_X1 U9343 ( .A(P1_REG3_REG_18__SCAN_IN), .ZN(n8145) );
  OAI21_X1 U9344 ( .B1(n8147), .B2(n8146), .A(n8145), .ZN(n8148) );
  NAND2_X1 U9345 ( .A1(n8148), .A2(n8157), .ZN(n9867) );
  OR2_X1 U9346 ( .A1(n9867), .A2(n8160), .ZN(n8151) );
  AOI22_X1 U9347 ( .A1(n6775), .A2(P1_REG2_REG_18__SCAN_IN), .B1(n5475), .B2(
        P1_REG0_REG_18__SCAN_IN), .ZN(n8150) );
  NAND2_X1 U9348 ( .A1(n6774), .A2(P1_REG1_REG_18__SCAN_IN), .ZN(n8149) );
  OR2_X1 U9349 ( .A1(n9873), .A2(n9882), .ZN(n8469) );
  NAND2_X1 U9350 ( .A1(n9873), .A2(n9882), .ZN(n8470) );
  INV_X1 U9351 ( .A(n9882), .ZN(n9615) );
  NAND2_X1 U9352 ( .A1(n9873), .A2(n9615), .ZN(n9837) );
  NAND2_X1 U9353 ( .A1(n8152), .A2(n7439), .ZN(n8155) );
  AOI22_X1 U9354 ( .A1(n8153), .A2(P2_DATAO_REG_19__SCAN_IN), .B1(n9772), .B2(
        n5192), .ZN(n8154) );
  INV_X1 U9355 ( .A(n8171), .ZN(n8159) );
  NAND2_X1 U9356 ( .A1(n8157), .A2(n8156), .ZN(n8158) );
  NAND2_X1 U9357 ( .A1(n8159), .A2(n8158), .ZN(n9839) );
  OR2_X1 U9358 ( .A1(n9839), .A2(n8160), .ZN(n8165) );
  INV_X1 U9359 ( .A(P1_REG2_REG_19__SCAN_IN), .ZN(n9840) );
  NAND2_X1 U9360 ( .A1(n6774), .A2(P1_REG1_REG_19__SCAN_IN), .ZN(n8162) );
  NAND2_X1 U9361 ( .A1(n5475), .A2(P1_REG0_REG_19__SCAN_IN), .ZN(n8161) );
  OAI211_X1 U9362 ( .C1(n8268), .C2(n9840), .A(n8162), .B(n8161), .ZN(n8163)
         );
  INV_X1 U9363 ( .A(n8163), .ZN(n8164) );
  NAND2_X1 U9364 ( .A1(n9961), .A2(n9824), .ZN(n8166) );
  NAND2_X1 U9365 ( .A1(n8167), .A2(n7439), .ZN(n8170) );
  OR2_X1 U9366 ( .A1(n8136), .A2(n8168), .ZN(n8169) );
  NOR2_X1 U9367 ( .A1(n8171), .A2(P1_REG3_REG_20__SCAN_IN), .ZN(n8172) );
  NAND2_X1 U9368 ( .A1(n5485), .A2(n4856), .ZN(n8178) );
  INV_X1 U9369 ( .A(P1_REG1_REG_20__SCAN_IN), .ZN(n8175) );
  NAND2_X1 U9370 ( .A1(n5475), .A2(P1_REG0_REG_20__SCAN_IN), .ZN(n8174) );
  NAND2_X1 U9371 ( .A1(n6775), .A2(P1_REG2_REG_20__SCAN_IN), .ZN(n8173) );
  OAI211_X1 U9372 ( .C1(n8175), .C2(n8341), .A(n8174), .B(n8173), .ZN(n8176)
         );
  INV_X1 U9373 ( .A(n8176), .ZN(n8177) );
  OR2_X1 U9374 ( .A1(n8136), .A2(n8180), .ZN(n8181) );
  OR2_X1 U9375 ( .A1(n8183), .A2(P1_REG3_REG_21__SCAN_IN), .ZN(n8184) );
  AND2_X1 U9376 ( .A1(n8184), .A2(n8197), .ZN(n9816) );
  NAND2_X1 U9377 ( .A1(n9816), .A2(n4856), .ZN(n8190) );
  INV_X1 U9378 ( .A(P1_REG1_REG_21__SCAN_IN), .ZN(n8187) );
  NAND2_X1 U9379 ( .A1(n6775), .A2(P1_REG2_REG_21__SCAN_IN), .ZN(n8186) );
  NAND2_X1 U9380 ( .A1(n5475), .A2(P1_REG0_REG_21__SCAN_IN), .ZN(n8185) );
  OAI211_X1 U9381 ( .C1(n8187), .C2(n8341), .A(n8186), .B(n8185), .ZN(n8188)
         );
  INV_X1 U9382 ( .A(n8188), .ZN(n8189) );
  OR2_X1 U9383 ( .A1(n9950), .A2(n9581), .ZN(n8435) );
  NAND2_X1 U9384 ( .A1(n9950), .A2(n9581), .ZN(n8463) );
  INV_X1 U9385 ( .A(n9581), .ZN(n9825) );
  NAND2_X1 U9386 ( .A1(n9950), .A2(n9825), .ZN(n8192) );
  NAND2_X1 U9387 ( .A1(n8193), .A2(n7439), .ZN(n8196) );
  OR2_X1 U9388 ( .A1(n8136), .A2(n8194), .ZN(n8195) );
  NAND2_X1 U9389 ( .A1(n6774), .A2(P1_REG1_REG_22__SCAN_IN), .ZN(n8206) );
  INV_X1 U9390 ( .A(P1_REG3_REG_22__SCAN_IN), .ZN(n8198) );
  NAND2_X1 U9391 ( .A1(n8198), .A2(n8197), .ZN(n8200) );
  AND2_X1 U9392 ( .A1(n8200), .A2(n8199), .ZN(n9795) );
  NAND2_X1 U9393 ( .A1(n4856), .A2(n9795), .ZN(n8205) );
  INV_X1 U9394 ( .A(P1_REG0_REG_22__SCAN_IN), .ZN(n8201) );
  OR2_X1 U9395 ( .A1(n8270), .A2(n8201), .ZN(n8204) );
  INV_X1 U9396 ( .A(P1_REG2_REG_22__SCAN_IN), .ZN(n8202) );
  OR2_X1 U9397 ( .A1(n8268), .A2(n8202), .ZN(n8203) );
  OR2_X1 U9398 ( .A1(n9944), .A2(n9811), .ZN(n8207) );
  NAND2_X1 U9399 ( .A1(n8208), .A2(n7439), .ZN(n8211) );
  OR2_X1 U9400 ( .A1(n8136), .A2(n8209), .ZN(n8210) );
  OR2_X1 U9401 ( .A1(n9939), .A2(n9766), .ZN(n8521) );
  NAND2_X1 U9402 ( .A1(n9939), .A2(n9766), .ZN(n8522) );
  NAND2_X1 U9403 ( .A1(n9939), .A2(n9801), .ZN(n9760) );
  OR2_X1 U9404 ( .A1(n8136), .A2(n8213), .ZN(n8214) );
  INV_X1 U9405 ( .A(n8216), .ZN(n8232) );
  INV_X1 U9406 ( .A(P1_REG3_REG_24__SCAN_IN), .ZN(n8217) );
  NAND2_X1 U9407 ( .A1(n8218), .A2(n8217), .ZN(n8219) );
  AND2_X1 U9408 ( .A1(n8232), .A2(n8219), .ZN(n9770) );
  NAND2_X1 U9409 ( .A1(n4856), .A2(n9770), .ZN(n8225) );
  NAND2_X1 U9410 ( .A1(n6774), .A2(P1_REG1_REG_24__SCAN_IN), .ZN(n8224) );
  INV_X1 U9411 ( .A(P1_REG2_REG_24__SCAN_IN), .ZN(n8220) );
  OR2_X1 U9412 ( .A1(n8268), .A2(n8220), .ZN(n8223) );
  INV_X1 U9413 ( .A(P1_REG0_REG_24__SCAN_IN), .ZN(n8221) );
  OR2_X1 U9414 ( .A1(n8270), .A2(n8221), .ZN(n8222) );
  NAND2_X1 U9415 ( .A1(n9935), .A2(n9754), .ZN(n8240) );
  AND2_X1 U9416 ( .A1(n9760), .A2(n8240), .ZN(n9740) );
  NAND2_X1 U9417 ( .A1(n8226), .A2(n7439), .ZN(n8229) );
  OR2_X1 U9418 ( .A1(n8136), .A2(n8227), .ZN(n8228) );
  INV_X1 U9419 ( .A(n8230), .ZN(n8249) );
  INV_X1 U9420 ( .A(P1_REG3_REG_25__SCAN_IN), .ZN(n8231) );
  NAND2_X1 U9421 ( .A1(n8232), .A2(n8231), .ZN(n8233) );
  NAND2_X1 U9422 ( .A1(n4856), .A2(n9748), .ZN(n8239) );
  NAND2_X1 U9423 ( .A1(n6774), .A2(P1_REG1_REG_25__SCAN_IN), .ZN(n8238) );
  INV_X1 U9424 ( .A(P1_REG2_REG_25__SCAN_IN), .ZN(n8234) );
  OR2_X1 U9425 ( .A1(n8268), .A2(n8234), .ZN(n8237) );
  INV_X1 U9426 ( .A(P1_REG0_REG_25__SCAN_IN), .ZN(n8235) );
  OR2_X1 U9427 ( .A1(n8270), .A2(n8235), .ZN(n8236) );
  NAND2_X1 U9428 ( .A1(n9928), .A2(n9768), .ZN(n8457) );
  NAND2_X1 U9429 ( .A1(n8458), .A2(n8457), .ZN(n9743) );
  AND2_X1 U9430 ( .A1(n9740), .A2(n9743), .ZN(n8242) );
  INV_X1 U9431 ( .A(n8240), .ZN(n8241) );
  OR2_X1 U9432 ( .A1(n9935), .A2(n9783), .ZN(n8526) );
  NAND2_X1 U9433 ( .A1(n9935), .A2(n9783), .ZN(n8527) );
  INV_X1 U9434 ( .A(n9768), .ZN(n9614) );
  INV_X1 U9435 ( .A(n9728), .ZN(n8257) );
  NAND2_X1 U9436 ( .A1(n8243), .A2(n7439), .ZN(n8246) );
  OR2_X1 U9437 ( .A1(n8136), .A2(n8244), .ZN(n8245) );
  INV_X1 U9438 ( .A(n8247), .ZN(n8264) );
  INV_X1 U9439 ( .A(P1_REG3_REG_26__SCAN_IN), .ZN(n8248) );
  NAND2_X1 U9440 ( .A1(n8249), .A2(n8248), .ZN(n8250) );
  NAND2_X1 U9441 ( .A1(n4856), .A2(n9734), .ZN(n8256) );
  NAND2_X1 U9442 ( .A1(n6774), .A2(P1_REG1_REG_26__SCAN_IN), .ZN(n8255) );
  INV_X1 U9443 ( .A(P1_REG2_REG_26__SCAN_IN), .ZN(n8251) );
  OR2_X1 U9444 ( .A1(n8268), .A2(n8251), .ZN(n8254) );
  INV_X1 U9445 ( .A(P1_REG0_REG_26__SCAN_IN), .ZN(n8252) );
  OR2_X1 U9446 ( .A1(n8270), .A2(n8252), .ZN(n8253) );
  NAND2_X1 U9447 ( .A1(n9923), .A2(n8667), .ZN(n8284) );
  NAND2_X1 U9448 ( .A1(n8454), .A2(n8284), .ZN(n8531) );
  NAND2_X1 U9449 ( .A1(n9923), .A2(n9755), .ZN(n8258) );
  NAND2_X1 U9450 ( .A1(n8259), .A2(n7439), .ZN(n8262) );
  OR2_X1 U9451 ( .A1(n8136), .A2(n8260), .ZN(n8261) );
  INV_X1 U9452 ( .A(P1_REG3_REG_27__SCAN_IN), .ZN(n8263) );
  NAND2_X1 U9453 ( .A1(n8264), .A2(n8263), .ZN(n8265) );
  NAND2_X1 U9454 ( .A1(n4856), .A2(n9713), .ZN(n8274) );
  NAND2_X1 U9455 ( .A1(n6774), .A2(P1_REG1_REG_27__SCAN_IN), .ZN(n8273) );
  INV_X1 U9456 ( .A(P1_REG2_REG_27__SCAN_IN), .ZN(n8267) );
  OR2_X1 U9457 ( .A1(n8268), .A2(n8267), .ZN(n8272) );
  INV_X1 U9458 ( .A(P1_REG0_REG_27__SCAN_IN), .ZN(n8269) );
  OR2_X1 U9459 ( .A1(n8270), .A2(n8269), .ZN(n8271) );
  NAND2_X1 U9460 ( .A1(n9920), .A2(n9726), .ZN(n8535) );
  NAND2_X1 U9461 ( .A1(n8604), .A2(n7439), .ZN(n8276) );
  OR2_X1 U9462 ( .A1(n8136), .A2(n7016), .ZN(n8275) );
  NAND2_X1 U9463 ( .A1(n8278), .A2(n8277), .ZN(n8279) );
  NAND2_X1 U9464 ( .A1(n9857), .A2(n8470), .ZN(n9845) );
  OR2_X1 U9465 ( .A1(n9961), .A2(n9861), .ZN(n8467) );
  NAND2_X1 U9466 ( .A1(n9961), .A2(n9861), .ZN(n8468) );
  INV_X1 U9467 ( .A(n8468), .ZN(n8405) );
  AOI21_X2 U9468 ( .B1(n9845), .B2(n9846), .A(n8405), .ZN(n9823) );
  XNOR2_X1 U9469 ( .A(n9954), .B(n9810), .ZN(n9822) );
  INV_X1 U9470 ( .A(n9822), .ZN(n8282) );
  AND2_X1 U9471 ( .A1(n9954), .A2(n9848), .ZN(n8403) );
  INV_X1 U9472 ( .A(n8403), .ZN(n8281) );
  NAND2_X1 U9473 ( .A1(n9808), .A2(n9809), .ZN(n9807) );
  OR2_X1 U9474 ( .A1(n9944), .A2(n9782), .ZN(n8461) );
  NAND2_X1 U9475 ( .A1(n9944), .A2(n9782), .ZN(n8462) );
  INV_X1 U9476 ( .A(n8462), .ZN(n8283) );
  INV_X1 U9477 ( .A(n8522), .ZN(n8415) );
  NAND2_X1 U9478 ( .A1(n9752), .A2(n9753), .ZN(n9751) );
  NAND2_X1 U9479 ( .A1(n9751), .A2(n8457), .ZN(n9725) );
  INV_X1 U9480 ( .A(n8284), .ZN(n8456) );
  AOI21_X1 U9481 ( .B1(n9725), .B2(n9727), .A(n8456), .ZN(n9718) );
  NAND2_X1 U9482 ( .A1(n4856), .A2(n8331), .ZN(n8289) );
  NAND2_X1 U9483 ( .A1(n6774), .A2(P1_REG1_REG_29__SCAN_IN), .ZN(n8288) );
  NAND2_X1 U9484 ( .A1(n6775), .A2(P1_REG2_REG_29__SCAN_IN), .ZN(n8287) );
  NAND2_X1 U9485 ( .A1(n5475), .A2(P1_REG0_REG_29__SCAN_IN), .ZN(n8286) );
  OAI22_X1 U9486 ( .A1(n8694), .A2(n9881), .B1(n9726), .B2(n9879), .ZN(n8290)
         );
  INV_X1 U9487 ( .A(n9920), .ZN(n8292) );
  INV_X1 U9488 ( .A(n9928), .ZN(n9750) );
  INV_X1 U9489 ( .A(n9950), .ZN(n8641) );
  INV_X1 U9490 ( .A(n9961), .ZN(n9513) );
  NAND2_X1 U9491 ( .A1(n9868), .A2(n9513), .ZN(n9842) );
  NOR2_X2 U9492 ( .A1(n9842), .A2(n9954), .ZN(n9829) );
  NAND2_X1 U9493 ( .A1(n9750), .A2(n9769), .ZN(n9745) );
  NOR2_X2 U9494 ( .A1(n9745), .A2(n9923), .ZN(n9733) );
  AOI21_X1 U9495 ( .B1(n8291), .B2(n9710), .A(n8329), .ZN(n9915) );
  INV_X1 U9496 ( .A(n8291), .ZN(n8687) );
  AOI22_X1 U9497 ( .A1(n9896), .A2(P1_REG2_REG_28__SCAN_IN), .B1(n8691), .B2(
        n10638), .ZN(n8293) );
  OAI21_X1 U9498 ( .B1(n8687), .B2(n9898), .A(n8293), .ZN(n8296) );
  NOR2_X1 U9499 ( .A1(n9917), .A2(n9899), .ZN(n8295) );
  AOI211_X1 U9500 ( .C1(n9902), .C2(n9915), .A(n8296), .B(n8295), .ZN(n8297)
         );
  OAI21_X1 U9501 ( .B1(n5487), .B2(n9896), .A(n8297), .ZN(P1_U3263) );
  XOR2_X1 U9502 ( .A(n8299), .B(n8298), .Z(n8304) );
  AOI22_X1 U9503 ( .A1(n8301), .A2(n9607), .B1(n8300), .B2(
        P1_REG3_REG_2__SCAN_IN), .ZN(n8303) );
  AOI22_X1 U9504 ( .A1(n9601), .A2(n9629), .B1(n9566), .B2(n6896), .ZN(n8302)
         );
  OAI211_X1 U9505 ( .C1(n8304), .C2(n9609), .A(n8303), .B(n8302), .ZN(P1_U3235) );
  OR2_X1 U9506 ( .A1(n8939), .A2(n9060), .ZN(n8308) );
  AOI21_X1 U9507 ( .B1(n10284), .B2(n8306), .A(n8305), .ZN(n8307) );
  OAI211_X1 U9508 ( .C1(n9058), .C2(n9015), .A(n8308), .B(n8307), .ZN(n8309)
         );
  AOI21_X1 U9509 ( .B1(n8310), .B2(n10293), .A(n8309), .ZN(n8314) );
  OAI22_X1 U9510 ( .A1(n8311), .A2(n10288), .B1(n9060), .B2(n9017), .ZN(n8312)
         );
  NAND3_X1 U9511 ( .A1(n4943), .A2(n7903), .A3(n8312), .ZN(n8313) );
  OAI211_X1 U9512 ( .C1(n8315), .C2(n10288), .A(n8314), .B(n8313), .ZN(
        P2_U3243) );
  OAI222_X1 U9513 ( .A1(n6175), .A2(P2_U3152), .B1(n4857), .B2(n8317), .C1(
        n8316), .C2(n9491), .ZN(P2_U3336) );
  OAI21_X1 U9514 ( .B1(n8687), .B2(n9721), .A(n8318), .ZN(n8328) );
  NAND2_X1 U9515 ( .A1(n8320), .A2(n8319), .ZN(n8324) );
  INV_X1 U9516 ( .A(n8321), .ZN(n8322) );
  NAND2_X1 U9517 ( .A1(n8322), .A2(n10165), .ZN(n8323) );
  MUX2_X1 U9518 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(P2_DATAO_REG_29__SCAN_IN), 
        .S(n8387), .Z(n8351) );
  INV_X1 U9519 ( .A(SI_29_), .ZN(n10164) );
  XNOR2_X1 U9520 ( .A(n8351), .B(n10164), .ZN(n8349) );
  NAND2_X1 U9521 ( .A1(n9490), .A2(n7439), .ZN(n8326) );
  INV_X1 U9522 ( .A(P2_DATAO_REG_29__SCAN_IN), .ZN(n10040) );
  OR2_X1 U9523 ( .A1(n8136), .A2(n10040), .ZN(n8325) );
  INV_X1 U9524 ( .A(n8327), .ZN(n8333) );
  INV_X1 U9525 ( .A(n8694), .ZN(n9612) );
  AOI21_X1 U9526 ( .B1(n8327), .B2(n8330), .A(n9703), .ZN(n9911) );
  AOI22_X1 U9527 ( .A1(n9896), .A2(P1_REG2_REG_29__SCAN_IN), .B1(n8331), .B2(
        n10638), .ZN(n8332) );
  OAI21_X1 U9528 ( .B1(n8333), .B2(n9898), .A(n8332), .ZN(n8347) );
  NOR2_X1 U9529 ( .A1(n8334), .A2(n8453), .ZN(n8335) );
  XNOR2_X1 U9530 ( .A(n8335), .B(n8380), .ZN(n8345) );
  INV_X1 U9531 ( .A(P1_B_REG_SCAN_IN), .ZN(n8336) );
  NOR2_X1 U9532 ( .A1(n4860), .A2(n8336), .ZN(n8337) );
  NOR2_X1 U9533 ( .A1(n9881), .A2(n8337), .ZN(n9696) );
  INV_X1 U9534 ( .A(P1_REG1_REG_30__SCAN_IN), .ZN(n8340) );
  NAND2_X1 U9535 ( .A1(n6775), .A2(P1_REG2_REG_30__SCAN_IN), .ZN(n8339) );
  NAND2_X1 U9536 ( .A1(n5475), .A2(P1_REG0_REG_30__SCAN_IN), .ZN(n8338) );
  OAI211_X1 U9537 ( .C1(n8341), .C2(n8340), .A(n8339), .B(n8338), .ZN(n9611)
         );
  NOR2_X1 U9538 ( .A1(n9913), .A2(n9896), .ZN(n8346) );
  OAI21_X1 U9539 ( .B1(n9853), .B2(n9914), .A(n8348), .ZN(P1_U3355) );
  INV_X1 U9540 ( .A(n8351), .ZN(n8352) );
  NAND2_X1 U9541 ( .A1(n8352), .A2(n10164), .ZN(n8353) );
  MUX2_X1 U9542 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(P2_DATAO_REG_30__SCAN_IN), 
        .S(n8387), .Z(n8383) );
  INV_X1 U9543 ( .A(SI_30_), .ZN(n10161) );
  XNOR2_X1 U9544 ( .A(n8383), .B(n10161), .ZN(n8381) );
  INV_X1 U9545 ( .A(P2_DATAO_REG_30__SCAN_IN), .ZN(n10035) );
  NOR2_X1 U9546 ( .A1(n8136), .A2(n10035), .ZN(n8355) );
  NOR2_X1 U9547 ( .A1(n9702), .A2(n9611), .ZN(n8586) );
  INV_X1 U9548 ( .A(n9798), .ZN(n9792) );
  INV_X1 U9549 ( .A(n9859), .ZN(n8375) );
  NAND4_X1 U9550 ( .A1(n8360), .A2(n8359), .A3(n8358), .A4(n8357), .ZN(n8361)
         );
  NOR4_X1 U9551 ( .A1(n8364), .A2(n8363), .A3(n8362), .A4(n8361), .ZN(n8366)
         );
  NAND4_X1 U9552 ( .A1(n5002), .A2(n8367), .A3(n8366), .A4(n8365), .ZN(n8368)
         );
  NOR4_X1 U9553 ( .A1(n8369), .A2(n10619), .A3(n8482), .A4(n8368), .ZN(n8370)
         );
  NAND4_X1 U9554 ( .A1(n8372), .A2(n8500), .A3(n8371), .A4(n8370), .ZN(n8373)
         );
  NOR4_X1 U9555 ( .A1(n8375), .A2(n8374), .A3(n9884), .A4(n8373), .ZN(n8376)
         );
  NAND4_X1 U9556 ( .A1(n9809), .A2(n9846), .A3(n8376), .A4(n9822), .ZN(n8377)
         );
  NOR4_X1 U9557 ( .A1(n9762), .A2(n9779), .A3(n9792), .A4(n8377), .ZN(n8378)
         );
  NAND4_X1 U9558 ( .A1(n9717), .A2(n9727), .A3(n9753), .A4(n8378), .ZN(n8379)
         );
  NOR4_X1 U9559 ( .A1(n8586), .A2(n8536), .A3(n8380), .A4(n8379), .ZN(n8395)
         );
  NAND2_X1 U9560 ( .A1(n8382), .A2(n8381), .ZN(n8386) );
  INV_X1 U9561 ( .A(n8383), .ZN(n8384) );
  NAND2_X1 U9562 ( .A1(n8384), .A2(n10161), .ZN(n8385) );
  MUX2_X1 U9563 ( .A(P1_DATAO_REG_31__SCAN_IN), .B(P2_DATAO_REG_31__SCAN_IN), 
        .S(n8387), .Z(n8389) );
  INV_X1 U9564 ( .A(SI_31_), .ZN(n8388) );
  XNOR2_X1 U9565 ( .A(n8389), .B(n8388), .ZN(n8390) );
  NAND2_X1 U9566 ( .A1(n8727), .A2(n7439), .ZN(n8393) );
  OR2_X1 U9567 ( .A1(n8136), .A2(n6424), .ZN(n8392) );
  INV_X1 U9568 ( .A(n8591), .ZN(n8394) );
  NAND2_X1 U9569 ( .A1(n8395), .A2(n8394), .ZN(n8398) );
  INV_X1 U9570 ( .A(n9695), .ZN(n8396) );
  AND2_X1 U9571 ( .A1(n9694), .A2(n8396), .ZN(n8399) );
  INV_X1 U9572 ( .A(n8399), .ZN(n8551) );
  AND2_X1 U9573 ( .A1(n9702), .A2(n9611), .ZN(n8545) );
  INV_X1 U9574 ( .A(n8545), .ZN(n8397) );
  NAND2_X1 U9575 ( .A1(n8551), .A2(n8397), .ZN(n8556) );
  OAI21_X1 U9576 ( .B1(n8398), .B2(n8556), .A(n4855), .ZN(n8552) );
  INV_X1 U9577 ( .A(n8552), .ZN(n8452) );
  AOI21_X1 U9578 ( .B1(n8545), .B2(n9695), .A(n8399), .ZN(n8548) );
  NAND2_X1 U9579 ( .A1(n8534), .A2(n8456), .ZN(n8400) );
  NAND3_X1 U9580 ( .A1(n8401), .A2(n8535), .A3(n8400), .ZN(n8584) );
  NAND2_X1 U9581 ( .A1(n8457), .A2(n8527), .ZN(n8443) );
  NAND2_X1 U9582 ( .A1(n8435), .A2(n8403), .ZN(n8404) );
  AND2_X1 U9583 ( .A1(n8404), .A2(n8463), .ZN(n8465) );
  NAND2_X1 U9584 ( .A1(n8465), .A2(n8462), .ZN(n8438) );
  OR2_X1 U9585 ( .A1(n8438), .A2(n8405), .ZN(n8433) );
  AND2_X1 U9586 ( .A1(n8512), .A2(n8508), .ZN(n8406) );
  NAND2_X1 U9587 ( .A1(n8470), .A2(n8406), .ZN(n8430) );
  NAND2_X1 U9588 ( .A1(n8503), .A2(n8494), .ZN(n8424) );
  NAND2_X1 U9589 ( .A1(n8474), .A2(n8407), .ZN(n8408) );
  NAND2_X1 U9590 ( .A1(n8408), .A2(n8473), .ZN(n8409) );
  NAND2_X1 U9591 ( .A1(n8479), .A2(n8409), .ZN(n8418) );
  INV_X1 U9592 ( .A(n8418), .ZN(n8412) );
  NAND4_X1 U9593 ( .A1(n8486), .A2(n8412), .A3(n8411), .A4(n8410), .ZN(n8413)
         );
  OR4_X1 U9594 ( .A1(n8430), .A2(n8495), .A3(n8424), .A4(n8413), .ZN(n8414) );
  OR4_X1 U9595 ( .A1(n8443), .A2(n8415), .A3(n8433), .A4(n8414), .ZN(n8580) );
  AND3_X1 U9596 ( .A1(n8473), .A2(n8416), .A3(n8472), .ZN(n8417) );
  NOR2_X1 U9597 ( .A1(n8418), .A2(n8417), .ZN(n8420) );
  OAI211_X1 U9598 ( .C1(n8421), .C2(n8420), .A(n8419), .B(n8486), .ZN(n8423)
         );
  AND3_X1 U9599 ( .A1(n8496), .A2(n8423), .A3(n8422), .ZN(n8425) );
  OAI211_X1 U9600 ( .C1(n8425), .C2(n8424), .A(n8507), .B(n8502), .ZN(n8426)
         );
  INV_X1 U9601 ( .A(n8426), .ZN(n8429) );
  INV_X1 U9602 ( .A(n8511), .ZN(n8427) );
  NAND2_X1 U9603 ( .A1(n8470), .A2(n8427), .ZN(n8428) );
  OAI211_X1 U9604 ( .C1(n8430), .C2(n8429), .A(n8469), .B(n8428), .ZN(n8431)
         );
  INV_X1 U9605 ( .A(n8431), .ZN(n8432) );
  NOR2_X1 U9606 ( .A1(n8433), .A2(n8432), .ZN(n8440) );
  OR2_X1 U9607 ( .A1(n9954), .A2(n9848), .ZN(n8434) );
  NAND2_X1 U9608 ( .A1(n8435), .A2(n8434), .ZN(n8464) );
  INV_X1 U9609 ( .A(n8467), .ZN(n8436) );
  NOR2_X1 U9610 ( .A1(n8464), .A2(n8436), .ZN(n8437) );
  OAI211_X1 U9611 ( .C1(n8438), .C2(n8437), .A(n8521), .B(n8461), .ZN(n8439)
         );
  OAI21_X1 U9612 ( .B1(n8440), .B2(n8439), .A(n8522), .ZN(n8441) );
  AND2_X1 U9613 ( .A1(n8441), .A2(n8526), .ZN(n8442) );
  OR2_X1 U9614 ( .A1(n8443), .A2(n8442), .ZN(n8444) );
  AND3_X1 U9615 ( .A1(n8454), .A2(n8444), .A3(n8458), .ZN(n8581) );
  OAI211_X1 U9616 ( .C1(n5006), .C2(n8580), .A(n8581), .B(n8534), .ZN(n8445)
         );
  INV_X1 U9617 ( .A(n8445), .ZN(n8446) );
  NOR2_X1 U9618 ( .A1(n8584), .A2(n8446), .ZN(n8449) );
  AND2_X1 U9619 ( .A1(n8539), .A2(n8447), .ZN(n8544) );
  INV_X1 U9620 ( .A(n8544), .ZN(n8589) );
  INV_X1 U9621 ( .A(n9702), .ZN(n9907) );
  NAND2_X1 U9622 ( .A1(n9695), .A2(n9611), .ZN(n8448) );
  NAND2_X1 U9623 ( .A1(n9907), .A2(n8448), .ZN(n8546) );
  OAI211_X1 U9624 ( .C1(n8449), .C2(n8589), .A(n8546), .B(n8587), .ZN(n8450)
         );
  AOI211_X1 U9625 ( .C1(n8548), .C2(n8450), .A(n8591), .B(n4855), .ZN(n8451)
         );
  NOR2_X1 U9626 ( .A1(n8452), .A2(n8451), .ZN(n8554) );
  NOR2_X1 U9627 ( .A1(n8542), .A2(n8453), .ZN(n8541) );
  INV_X1 U9628 ( .A(n8454), .ZN(n8455) );
  MUX2_X1 U9629 ( .A(n8456), .B(n8455), .S(n8547), .Z(n8532) );
  INV_X1 U9630 ( .A(n8457), .ZN(n8460) );
  INV_X1 U9631 ( .A(n8458), .ZN(n8459) );
  INV_X1 U9632 ( .A(n8547), .ZN(n8533) );
  MUX2_X1 U9633 ( .A(n8460), .B(n8459), .S(n8533), .Z(n8530) );
  MUX2_X1 U9634 ( .A(n8462), .B(n8461), .S(n8547), .Z(n8519) );
  NAND2_X1 U9635 ( .A1(n8464), .A2(n8463), .ZN(n8466) );
  MUX2_X1 U9636 ( .A(n8466), .B(n8465), .S(n8547), .Z(n8517) );
  MUX2_X1 U9637 ( .A(n8468), .B(n8467), .S(n8547), .Z(n8515) );
  MUX2_X1 U9638 ( .A(n8470), .B(n8469), .S(n8533), .Z(n8514) );
  MUX2_X1 U9639 ( .A(n8474), .B(n8473), .S(n8533), .Z(n8475) );
  OAI211_X1 U9640 ( .C1(n8477), .C2(n10619), .A(n8476), .B(n8475), .ZN(n8484)
         );
  MUX2_X1 U9641 ( .A(n8479), .B(n8478), .S(n8547), .Z(n8480) );
  INV_X1 U9642 ( .A(n8480), .ZN(n8481) );
  NOR2_X1 U9643 ( .A1(n8482), .A2(n8481), .ZN(n8483) );
  NAND2_X1 U9644 ( .A1(n8484), .A2(n8483), .ZN(n8487) );
  AOI21_X1 U9645 ( .B1(n8487), .B2(n8485), .A(n8495), .ZN(n8489) );
  AOI21_X1 U9646 ( .B1(n8487), .B2(n8486), .A(n8493), .ZN(n8488) );
  MUX2_X1 U9647 ( .A(n8489), .B(n8488), .S(n8547), .Z(n8492) );
  MUX2_X1 U9648 ( .A(n8494), .B(n8496), .S(n8547), .Z(n8490) );
  OAI21_X1 U9649 ( .B1(n8492), .B2(n8491), .A(n8490), .ZN(n8501) );
  NAND2_X1 U9650 ( .A1(n8494), .A2(n8493), .ZN(n8498) );
  NAND2_X1 U9651 ( .A1(n8496), .A2(n8495), .ZN(n8497) );
  MUX2_X1 U9652 ( .A(n8498), .B(n8497), .S(n8547), .Z(n8499) );
  NAND3_X1 U9653 ( .A1(n8501), .A2(n8500), .A3(n8499), .ZN(n8505) );
  MUX2_X1 U9654 ( .A(n8503), .B(n8502), .S(n8547), .Z(n8504) );
  NAND3_X1 U9655 ( .A1(n8506), .A2(n8505), .A3(n8504), .ZN(n8510) );
  MUX2_X1 U9656 ( .A(n8508), .B(n8507), .S(n8533), .Z(n8509) );
  MUX2_X1 U9657 ( .A(n8512), .B(n8511), .S(n8547), .Z(n8513) );
  NAND3_X1 U9658 ( .A1(n9798), .A2(n8517), .A3(n8516), .ZN(n8518) );
  NAND3_X1 U9659 ( .A1(n8520), .A2(n8519), .A3(n8518), .ZN(n8524) );
  MUX2_X1 U9660 ( .A(n8522), .B(n8521), .S(n8533), .Z(n8523) );
  NAND2_X1 U9661 ( .A1(n8524), .A2(n8523), .ZN(n8525) );
  NAND2_X1 U9662 ( .A1(n9764), .A2(n8525), .ZN(n8529) );
  MUX2_X1 U9663 ( .A(n8527), .B(n8526), .S(n8533), .Z(n8528) );
  MUX2_X1 U9664 ( .A(n8535), .B(n8534), .S(n8533), .Z(n8537) );
  NAND3_X1 U9665 ( .A1(n8538), .A2(n8537), .A3(n8277), .ZN(n8543) );
  NOR2_X1 U9666 ( .A1(n8548), .A2(n8547), .ZN(n8549) );
  AOI211_X1 U9667 ( .C1(n8551), .C2(n8550), .A(n8591), .B(n8549), .ZN(n8555)
         );
  INV_X1 U9668 ( .A(n8556), .ZN(n8593) );
  INV_X1 U9669 ( .A(n8557), .ZN(n8578) );
  INV_X1 U9670 ( .A(n8558), .ZN(n8576) );
  AOI21_X1 U9671 ( .B1(n6896), .B2(n10491), .A(n4855), .ZN(n8563) );
  INV_X1 U9672 ( .A(n8559), .ZN(n8562) );
  AOI211_X1 U9673 ( .C1(n8563), .C2(n8562), .A(n5359), .B(n8561), .ZN(n8567)
         );
  INV_X1 U9674 ( .A(n8564), .ZN(n8566) );
  OAI21_X1 U9675 ( .B1(n8567), .B2(n8566), .A(n8565), .ZN(n8574) );
  AOI22_X1 U9676 ( .A1(n8569), .A2(n9628), .B1(n8568), .B2(n9629), .ZN(n8573)
         );
  INV_X1 U9677 ( .A(n8571), .ZN(n8572) );
  AOI211_X1 U9678 ( .C1(n8574), .C2(n8573), .A(n5023), .B(n8572), .ZN(n8575)
         );
  AOI211_X1 U9679 ( .C1(n8578), .C2(n8577), .A(n8576), .B(n8575), .ZN(n8579)
         );
  NOR2_X1 U9680 ( .A1(n8580), .A2(n8579), .ZN(n8583) );
  INV_X1 U9681 ( .A(n8581), .ZN(n8582) );
  NOR3_X1 U9682 ( .A1(n9708), .A2(n8583), .A3(n8582), .ZN(n8585) );
  NOR2_X1 U9683 ( .A1(n8585), .A2(n8584), .ZN(n8590) );
  INV_X1 U9684 ( .A(n8586), .ZN(n8588) );
  OAI211_X1 U9685 ( .C1(n8590), .C2(n8589), .A(n8588), .B(n8587), .ZN(n8592)
         );
  AOI21_X1 U9686 ( .B1(n8593), .B2(n8592), .A(n8591), .ZN(n8594) );
  NOR4_X1 U9687 ( .A1(n9879), .A2(n8597), .A3(n8596), .A4(n4860), .ZN(n8600)
         );
  OAI21_X1 U9688 ( .B1(n8598), .B2(n8601), .A(P1_B_REG_SCAN_IN), .ZN(n8599) );
  OAI22_X1 U9689 ( .A1(n8602), .A2(n8601), .B1(n8600), .B2(n8599), .ZN(
        P1_U3240) );
  INV_X1 U9690 ( .A(n8718), .ZN(n10038) );
  INV_X1 U9691 ( .A(P1_DATAO_REG_30__SCAN_IN), .ZN(n8716) );
  OAI222_X1 U9692 ( .A1(P2_U3152), .A2(n8603), .B1(n4857), .B2(n10038), .C1(
        n8716), .C2(n9491), .ZN(P2_U3328) );
  INV_X1 U9693 ( .A(n8604), .ZN(n8698) );
  OAI222_X1 U9694 ( .A1(P2_U3152), .A2(n6188), .B1(n4857), .B2(n8698), .C1(
        n8605), .C2(n9491), .ZN(P2_U3330) );
  NAND2_X1 U9695 ( .A1(n9532), .A2(n8672), .ZN(n8607) );
  NAND2_X1 U9696 ( .A1(n9617), .A2(n8678), .ZN(n8606) );
  NAND2_X1 U9697 ( .A1(n8607), .A2(n8606), .ZN(n8608) );
  XNOR2_X1 U9698 ( .A(n8608), .B(n8683), .ZN(n8611) );
  NOR2_X1 U9699 ( .A1(n9880), .A2(n8682), .ZN(n8609) );
  AOI21_X1 U9700 ( .B1(n9532), .B2(n8678), .A(n8609), .ZN(n8612) );
  XNOR2_X1 U9701 ( .A(n8611), .B(n8612), .ZN(n9535) );
  INV_X1 U9702 ( .A(n8611), .ZN(n8613) );
  NAND2_X1 U9703 ( .A1(n8613), .A2(n8612), .ZN(n8614) );
  NAND2_X1 U9704 ( .A1(n9973), .A2(n6773), .ZN(n8616) );
  OR2_X1 U9705 ( .A1(n9860), .A2(n8685), .ZN(n8615) );
  NAND2_X1 U9706 ( .A1(n8616), .A2(n8615), .ZN(n8617) );
  XNOR2_X1 U9707 ( .A(n8617), .B(n8675), .ZN(n9545) );
  NOR2_X1 U9708 ( .A1(n9860), .A2(n8682), .ZN(n8618) );
  AOI21_X1 U9709 ( .B1(n9973), .B2(n8678), .A(n8618), .ZN(n9544) );
  AND2_X1 U9710 ( .A1(n9545), .A2(n9544), .ZN(n8620) );
  NAND2_X1 U9711 ( .A1(n9873), .A2(n6773), .ZN(n8622) );
  NAND2_X1 U9712 ( .A1(n9615), .A2(n8678), .ZN(n8621) );
  NAND2_X1 U9713 ( .A1(n8622), .A2(n8621), .ZN(n8623) );
  NOR2_X1 U9714 ( .A1(n9882), .A2(n8682), .ZN(n8624) );
  AOI21_X1 U9715 ( .B1(n9873), .B2(n8678), .A(n8624), .ZN(n9587) );
  NAND2_X1 U9716 ( .A1(n9588), .A2(n9587), .ZN(n9585) );
  INV_X1 U9717 ( .A(n8625), .ZN(n8626) );
  NAND2_X2 U9718 ( .A1(n8626), .A2(n4931), .ZN(n9589) );
  OAI22_X1 U9719 ( .A1(n9513), .A2(n8685), .B1(n9861), .B2(n8682), .ZN(n8630)
         );
  NAND2_X1 U9720 ( .A1(n9961), .A2(n8672), .ZN(n8628) );
  NAND2_X1 U9721 ( .A1(n9824), .A2(n8678), .ZN(n8627) );
  NAND2_X1 U9722 ( .A1(n8628), .A2(n8627), .ZN(n8629) );
  XNOR2_X1 U9723 ( .A(n8629), .B(n8683), .ZN(n8631) );
  XOR2_X1 U9724 ( .A(n8630), .B(n8631), .Z(n9507) );
  NAND2_X1 U9725 ( .A1(n9954), .A2(n8672), .ZN(n8634) );
  OR2_X1 U9726 ( .A1(n9848), .A2(n8685), .ZN(n8633) );
  NAND2_X1 U9727 ( .A1(n8634), .A2(n8633), .ZN(n8635) );
  XNOR2_X1 U9728 ( .A(n8635), .B(n8675), .ZN(n8637) );
  NOR2_X1 U9729 ( .A1(n9848), .A2(n8682), .ZN(n8636) );
  AOI21_X1 U9730 ( .B1(n9954), .B2(n8678), .A(n8636), .ZN(n8638) );
  AND2_X1 U9731 ( .A1(n8637), .A2(n8638), .ZN(n9561) );
  INV_X1 U9732 ( .A(n8637), .ZN(n8640) );
  INV_X1 U9733 ( .A(n8638), .ZN(n8639) );
  NAND2_X1 U9734 ( .A1(n8640), .A2(n8639), .ZN(n9562) );
  OAI22_X1 U9735 ( .A1(n8641), .A2(n8686), .B1(n9581), .B2(n8685), .ZN(n8642)
         );
  XOR2_X1 U9736 ( .A(n8683), .B(n8642), .Z(n8644) );
  AOI22_X1 U9737 ( .A1(n9950), .A2(n8678), .B1(n6799), .B2(n9825), .ZN(n8643)
         );
  NOR2_X1 U9738 ( .A1(n8644), .A2(n8643), .ZN(n9516) );
  NAND2_X1 U9739 ( .A1(n8644), .A2(n8643), .ZN(n9515) );
  NAND2_X1 U9740 ( .A1(n9944), .A2(n6773), .ZN(n8646) );
  NAND2_X1 U9741 ( .A1(n9811), .A2(n8678), .ZN(n8645) );
  NAND2_X1 U9742 ( .A1(n8646), .A2(n8645), .ZN(n8647) );
  XNOR2_X1 U9743 ( .A(n8647), .B(n8675), .ZN(n8650) );
  NOR2_X1 U9744 ( .A1(n9782), .A2(n8682), .ZN(n8648) );
  AOI21_X1 U9745 ( .B1(n9944), .B2(n8678), .A(n8648), .ZN(n8649) );
  OR2_X1 U9746 ( .A1(n8650), .A2(n8649), .ZN(n9576) );
  NAND2_X1 U9747 ( .A1(n8650), .A2(n8649), .ZN(n9577) );
  NAND2_X1 U9748 ( .A1(n9574), .A2(n9577), .ZN(n8653) );
  OAI22_X1 U9749 ( .A1(n9789), .A2(n8686), .B1(n9766), .B2(n8685), .ZN(n8651)
         );
  XOR2_X1 U9750 ( .A(n8683), .B(n8651), .Z(n8652) );
  NAND2_X1 U9751 ( .A1(n8653), .A2(n8652), .ZN(n9495) );
  OAI22_X1 U9752 ( .A1(n9789), .A2(n8685), .B1(n9766), .B2(n8682), .ZN(n9498)
         );
  NOR2_X2 U9753 ( .A1(n8653), .A2(n8652), .ZN(n9497) );
  OAI22_X1 U9754 ( .A1(n5182), .A2(n8685), .B1(n9783), .B2(n8682), .ZN(n8657)
         );
  NAND2_X1 U9755 ( .A1(n9935), .A2(n8672), .ZN(n8655) );
  NAND2_X1 U9756 ( .A1(n9754), .A2(n8678), .ZN(n8654) );
  NAND2_X1 U9757 ( .A1(n8655), .A2(n8654), .ZN(n8656) );
  XNOR2_X1 U9758 ( .A(n8656), .B(n8683), .ZN(n8658) );
  XOR2_X1 U9759 ( .A(n8657), .B(n8658), .Z(n9555) );
  NAND2_X1 U9760 ( .A1(n9928), .A2(n6773), .ZN(n8661) );
  NAND2_X1 U9761 ( .A1(n9614), .A2(n8678), .ZN(n8660) );
  NAND2_X1 U9762 ( .A1(n8661), .A2(n8660), .ZN(n8662) );
  XNOR2_X1 U9763 ( .A(n8662), .B(n8675), .ZN(n9524) );
  NOR2_X1 U9764 ( .A1(n9768), .A2(n8682), .ZN(n8663) );
  AOI21_X1 U9765 ( .B1(n9928), .B2(n8678), .A(n8663), .ZN(n9523) );
  INV_X1 U9766 ( .A(n9524), .ZN(n8665) );
  INV_X1 U9767 ( .A(n9523), .ZN(n8664) );
  NOR2_X1 U9768 ( .A1(n8667), .A2(n8682), .ZN(n8666) );
  AOI21_X1 U9769 ( .B1(n9923), .B2(n8678), .A(n8666), .ZN(n8671) );
  INV_X1 U9770 ( .A(n9923), .ZN(n9736) );
  OAI22_X1 U9771 ( .A1(n9736), .A2(n8686), .B1(n8667), .B2(n8685), .ZN(n8668)
         );
  XNOR2_X1 U9772 ( .A(n8668), .B(n8683), .ZN(n8669) );
  XOR2_X1 U9773 ( .A(n8671), .B(n8669), .Z(n9600) );
  INV_X1 U9774 ( .A(n8669), .ZN(n8670) );
  NAND2_X1 U9775 ( .A1(n9920), .A2(n8672), .ZN(n8674) );
  NAND2_X1 U9776 ( .A1(n9613), .A2(n8678), .ZN(n8673) );
  NAND2_X1 U9777 ( .A1(n8674), .A2(n8673), .ZN(n8676) );
  XNOR2_X1 U9778 ( .A(n8676), .B(n8675), .ZN(n8680) );
  NOR2_X1 U9779 ( .A1(n9726), .A2(n8682), .ZN(n8677) );
  AOI21_X1 U9780 ( .B1(n9920), .B2(n8678), .A(n8677), .ZN(n8679) );
  NAND2_X1 U9781 ( .A1(n8680), .A2(n8679), .ZN(n8681) );
  OAI21_X1 U9782 ( .B1(n8680), .B2(n8679), .A(n8681), .ZN(n8699) );
  OAI22_X1 U9783 ( .A1(n8687), .A2(n8685), .B1(n9721), .B2(n8682), .ZN(n8684)
         );
  XNOR2_X1 U9784 ( .A(n8684), .B(n8683), .ZN(n8689) );
  OAI22_X1 U9785 ( .A1(n8687), .A2(n8686), .B1(n9721), .B2(n8685), .ZN(n8688)
         );
  XNOR2_X1 U9786 ( .A(n8689), .B(n8688), .ZN(n8690) );
  AOI22_X1 U9787 ( .A1(n9566), .A2(n9613), .B1(P1_REG3_REG_28__SCAN_IN), .B2(
        P1_U3084), .ZN(n8693) );
  NAND2_X1 U9788 ( .A1(n9602), .A2(n8691), .ZN(n8692) );
  OAI211_X1 U9789 ( .C1(n8694), .C2(n9569), .A(n8693), .B(n8692), .ZN(n8695)
         );
  AOI21_X1 U9790 ( .B1(n8291), .B2(n9607), .A(n8695), .ZN(n8696) );
  OAI21_X1 U9791 ( .B1(n8697), .B2(n9609), .A(n8696), .ZN(P1_U3218) );
  OAI222_X1 U9792 ( .A1(n10039), .A2(n7016), .B1(P1_U3084), .B2(n6363), .C1(
        n10033), .C2(n8698), .ZN(P1_U3325) );
  AOI21_X1 U9793 ( .B1(n8700), .B2(n8699), .A(n4899), .ZN(n8705) );
  AOI22_X1 U9794 ( .A1(n9566), .A2(n9755), .B1(P1_REG3_REG_27__SCAN_IN), .B2(
        P1_U3084), .ZN(n8702) );
  NAND2_X1 U9795 ( .A1(n9602), .A2(n9713), .ZN(n8701) );
  OAI211_X1 U9796 ( .C1(n9721), .C2(n9569), .A(n8702), .B(n8701), .ZN(n8703)
         );
  AOI21_X1 U9797 ( .B1(n9920), .B2(n9607), .A(n8703), .ZN(n8704) );
  OAI21_X1 U9798 ( .B1(n8705), .B2(n9609), .A(n8704), .ZN(P1_U3212) );
  NAND2_X1 U9799 ( .A1(n9457), .A2(n9338), .ZN(n8834) );
  NAND2_X1 U9800 ( .A1(n9451), .A2(n9129), .ZN(n8707) );
  NAND2_X1 U9801 ( .A1(n9335), .A2(n9328), .ZN(n9341) );
  NAND2_X1 U9802 ( .A1(n9341), .A2(n8708), .ZN(n9321) );
  NAND2_X1 U9803 ( .A1(n9448), .A2(n9339), .ZN(n8738) );
  NAND2_X1 U9804 ( .A1(n8739), .A2(n8738), .ZN(n9309) );
  INV_X1 U9805 ( .A(n9309), .ZN(n9320) );
  NAND2_X1 U9806 ( .A1(n9321), .A2(n9320), .ZN(n9319) );
  NAND2_X1 U9807 ( .A1(n9441), .A2(n9274), .ZN(n8841) );
  NAND2_X1 U9808 ( .A1(n9291), .A2(n9130), .ZN(n9295) );
  NAND2_X1 U9809 ( .A1(n9436), .A2(n9293), .ZN(n8844) );
  NAND2_X1 U9810 ( .A1(n9430), .A2(n9275), .ZN(n8847) );
  NAND2_X1 U9811 ( .A1(n8852), .A2(n8847), .ZN(n9262) );
  INV_X1 U9812 ( .A(n9262), .ZN(n9255) );
  NAND2_X1 U9813 ( .A1(n8709), .A2(n9264), .ZN(n9230) );
  INV_X1 U9814 ( .A(n9245), .ZN(n8920) );
  AND2_X1 U9815 ( .A1(n9420), .A2(n9138), .ZN(n8855) );
  INV_X1 U9816 ( .A(n8855), .ZN(n8850) );
  NAND2_X1 U9817 ( .A1(n8856), .A2(n8850), .ZN(n9137) );
  INV_X1 U9818 ( .A(n9230), .ZN(n8710) );
  NOR2_X1 U9819 ( .A1(n9137), .A2(n8710), .ZN(n8711) );
  NOR2_X1 U9820 ( .A1(n9417), .A2(n9233), .ZN(n8860) );
  INV_X1 U9821 ( .A(n8860), .ZN(n8712) );
  NAND2_X1 U9822 ( .A1(n9417), .A2(n9233), .ZN(n8862) );
  INV_X1 U9823 ( .A(n8861), .ZN(n8866) );
  NAND2_X1 U9824 ( .A1(n9411), .A2(n8991), .ZN(n8869) );
  NAND2_X1 U9825 ( .A1(n9405), .A2(n9053), .ZN(n8870) );
  NAND2_X1 U9826 ( .A1(n9400), .A2(n9146), .ZN(n8874) );
  NAND2_X1 U9827 ( .A1(n9490), .A2(n8726), .ZN(n8714) );
  INV_X1 U9828 ( .A(P1_DATAO_REG_29__SCAN_IN), .ZN(n9492) );
  OR2_X1 U9829 ( .A1(n5965), .A2(n9492), .ZN(n8713) );
  NAND2_X1 U9830 ( .A1(n9111), .A2(n8715), .ZN(n8868) );
  INV_X1 U9831 ( .A(n8868), .ZN(n8883) );
  NOR2_X1 U9832 ( .A1(n5965), .A2(n8716), .ZN(n8717) );
  INV_X1 U9833 ( .A(P2_REG0_REG_30__SCAN_IN), .ZN(n8721) );
  NAND2_X1 U9834 ( .A1(n5589), .A2(P2_REG2_REG_30__SCAN_IN), .ZN(n8720) );
  NAND2_X1 U9835 ( .A1(n6418), .A2(P2_REG1_REG_30__SCAN_IN), .ZN(n8719) );
  OAI211_X1 U9836 ( .C1(n5548), .C2(n8721), .A(n8720), .B(n8719), .ZN(n9052)
         );
  AND2_X1 U9837 ( .A1(n9393), .A2(n9052), .ZN(n8887) );
  OAI22_X1 U9838 ( .A1(n8723), .A2(n8887), .B1(n8928), .B2(n8722), .ZN(n8725)
         );
  NAND2_X1 U9839 ( .A1(n8723), .A2(n9393), .ZN(n8724) );
  NAND2_X1 U9840 ( .A1(n8725), .A2(n8724), .ZN(n8732) );
  NAND2_X1 U9841 ( .A1(n8727), .A2(n8726), .ZN(n8729) );
  OR2_X1 U9842 ( .A1(n5965), .A2(n6453), .ZN(n8728) );
  OR2_X1 U9843 ( .A1(n9386), .A2(n9114), .ZN(n8731) );
  INV_X1 U9844 ( .A(n9393), .ZN(n9119) );
  INV_X1 U9845 ( .A(n9052), .ZN(n9148) );
  AND2_X1 U9846 ( .A1(n9119), .A2(n9148), .ZN(n8886) );
  INV_X1 U9847 ( .A(n8886), .ZN(n8730) );
  NAND2_X1 U9848 ( .A1(n8731), .A2(n8730), .ZN(n8923) );
  NAND2_X1 U9849 ( .A1(n9386), .A2(n9114), .ZN(n8889) );
  AND2_X1 U9850 ( .A1(n8896), .A2(n8733), .ZN(n8931) );
  INV_X1 U9851 ( .A(n8870), .ZN(n8735) );
  AND2_X1 U9852 ( .A1(n8733), .A2(n9317), .ZN(n8734) );
  AND2_X1 U9853 ( .A1(n6175), .A2(n8734), .ZN(n8824) );
  NOR3_X1 U9854 ( .A1(n5438), .A2(n8735), .A3(n8824), .ZN(n8881) );
  NAND2_X1 U9855 ( .A1(n9451), .A2(n9057), .ZN(n8737) );
  MUX2_X1 U9856 ( .A(n9057), .B(n9451), .S(n8890), .Z(n8736) );
  AOI21_X1 U9857 ( .B1(n8737), .B2(n8736), .A(n9309), .ZN(n8839) );
  INV_X1 U9858 ( .A(n8738), .ZN(n8741) );
  INV_X1 U9859 ( .A(n8739), .ZN(n8740) );
  MUX2_X1 U9860 ( .A(n8741), .B(n8740), .S(n8890), .Z(n8838) );
  MUX2_X1 U9861 ( .A(n8743), .B(n8742), .S(n8824), .Z(n8832) );
  MUX2_X1 U9862 ( .A(n8745), .B(n8744), .S(n8890), .Z(n8829) );
  NAND2_X1 U9863 ( .A1(n8750), .A2(n5445), .ZN(n8746) );
  NAND3_X1 U9864 ( .A1(n8747), .A2(n8799), .A3(n8746), .ZN(n8749) );
  NAND2_X1 U9865 ( .A1(n8806), .A2(n8750), .ZN(n8748) );
  MUX2_X1 U9866 ( .A(n8749), .B(n8748), .S(n8890), .Z(n8817) );
  AOI21_X1 U9867 ( .B1(n8750), .B2(n8796), .A(n8890), .ZN(n8803) );
  NAND2_X1 U9868 ( .A1(n8752), .A2(n8751), .ZN(n8759) );
  AND2_X1 U9869 ( .A1(n8759), .A2(n8753), .ZN(n8757) );
  INV_X1 U9870 ( .A(n8754), .ZN(n9368) );
  INV_X1 U9871 ( .A(n8755), .ZN(n8756) );
  AOI21_X1 U9872 ( .B1(n8757), .B2(n9368), .A(n8756), .ZN(n8764) );
  OAI21_X1 U9873 ( .B1(n8759), .B2(n8928), .A(n8758), .ZN(n8762) );
  INV_X1 U9874 ( .A(n8760), .ZN(n8761) );
  AOI21_X1 U9875 ( .B1(n8762), .B2(n9368), .A(n8761), .ZN(n8763) );
  MUX2_X1 U9876 ( .A(n8764), .B(n8763), .S(n8890), .Z(n8771) );
  MUX2_X1 U9877 ( .A(n8767), .B(n8766), .S(n8890), .Z(n8769) );
  NOR2_X1 U9878 ( .A1(n8769), .A2(n8768), .ZN(n8770) );
  OAI21_X1 U9879 ( .B1(n8771), .B2(n8900), .A(n8770), .ZN(n8776) );
  MUX2_X1 U9880 ( .A(n8773), .B(n8772), .S(n8824), .Z(n8774) );
  NAND3_X1 U9881 ( .A1(n8776), .A2(n8775), .A3(n8774), .ZN(n8780) );
  MUX2_X1 U9882 ( .A(n8778), .B(n8777), .S(n8890), .Z(n8779) );
  NAND2_X1 U9883 ( .A1(n8780), .A2(n8779), .ZN(n8786) );
  MUX2_X1 U9884 ( .A(n8781), .B(n8784), .S(n8890), .Z(n8782) );
  INV_X1 U9885 ( .A(n8784), .ZN(n10562) );
  NAND3_X1 U9886 ( .A1(n8786), .A2(n8785), .A3(n10562), .ZN(n8787) );
  OR2_X1 U9887 ( .A1(n8789), .A2(n8890), .ZN(n8791) );
  NAND2_X1 U9888 ( .A1(n8789), .A2(n8890), .ZN(n8790) );
  MUX2_X1 U9889 ( .A(n8791), .B(n8790), .S(n8970), .Z(n8792) );
  MUX2_X1 U9890 ( .A(n8794), .B(n8793), .S(n8890), .Z(n8795) );
  NAND3_X1 U9891 ( .A1(n8797), .A2(n8796), .A3(n8795), .ZN(n8800) );
  NAND3_X1 U9892 ( .A1(n8800), .A2(n8799), .A3(n8798), .ZN(n8802) );
  OAI21_X1 U9893 ( .B1(n8803), .B2(n8802), .A(n8801), .ZN(n8816) );
  NAND2_X1 U9894 ( .A1(n8805), .A2(n8806), .ZN(n8808) );
  INV_X1 U9895 ( .A(n8806), .ZN(n8807) );
  AOI22_X1 U9896 ( .A1(n7840), .A2(n8808), .B1(n5204), .B2(n8807), .ZN(n8814)
         );
  NAND2_X1 U9897 ( .A1(n8810), .A2(n8809), .ZN(n8812) );
  AND2_X1 U9898 ( .A1(n8812), .A2(n8811), .ZN(n8813) );
  MUX2_X1 U9899 ( .A(n8814), .B(n8813), .S(n8890), .Z(n8815) );
  MUX2_X1 U9900 ( .A(n8819), .B(n8818), .S(n8890), .Z(n8820) );
  INV_X1 U9901 ( .A(n8822), .ZN(n8826) );
  INV_X1 U9902 ( .A(n8823), .ZN(n8825) );
  MUX2_X1 U9903 ( .A(n8826), .B(n8825), .S(n8824), .Z(n8827) );
  NAND3_X1 U9904 ( .A1(n9347), .A2(n8832), .A3(n8831), .ZN(n8836) );
  MUX2_X1 U9905 ( .A(n8834), .B(n8833), .S(n8890), .Z(n8835) );
  NAND4_X1 U9906 ( .A1(n9328), .A2(n9320), .A3(n8836), .A4(n8835), .ZN(n8837)
         );
  OAI211_X1 U9907 ( .C1(n8839), .C2(n8838), .A(n9130), .B(n8837), .ZN(n8843)
         );
  MUX2_X1 U9908 ( .A(n8841), .B(n8840), .S(n8890), .Z(n8842) );
  MUX2_X1 U9909 ( .A(n8845), .B(n8844), .S(n8890), .Z(n8846) );
  INV_X1 U9910 ( .A(n8847), .ZN(n8849) );
  OAI211_X1 U9911 ( .C1(n8854), .C2(n8849), .A(n8848), .B(n8856), .ZN(n8851)
         );
  NAND2_X1 U9912 ( .A1(n8851), .A2(n8850), .ZN(n8859) );
  INV_X1 U9913 ( .A(n8852), .ZN(n8853) );
  AOI21_X1 U9914 ( .B1(n8857), .B2(n8856), .A(n8855), .ZN(n8858) );
  NOR2_X1 U9915 ( .A1(n8861), .A2(n8860), .ZN(n8863) );
  MUX2_X1 U9916 ( .A(n8863), .B(n8862), .S(n8890), .Z(n8864) );
  INV_X1 U9917 ( .A(n8869), .ZN(n8867) );
  OAI211_X1 U9918 ( .C1(n8871), .C2(n8867), .A(n8872), .B(n8866), .ZN(n8880)
         );
  NAND3_X1 U9919 ( .A1(n8871), .A2(n8870), .A3(n8869), .ZN(n8873) );
  NAND3_X1 U9920 ( .A1(n8873), .A2(n8877), .A3(n8872), .ZN(n8875) );
  NAND2_X1 U9921 ( .A1(n8875), .A2(n8874), .ZN(n8876) );
  INV_X1 U9922 ( .A(n8877), .ZN(n8878) );
  INV_X1 U9923 ( .A(n8882), .ZN(n8884) );
  INV_X1 U9924 ( .A(n8887), .ZN(n8888) );
  NAND2_X1 U9925 ( .A1(n8889), .A2(n8888), .ZN(n8924) );
  MUX2_X1 U9926 ( .A(n8923), .B(n8924), .S(n8890), .Z(n8893) );
  MUX2_X1 U9927 ( .A(n9115), .B(n9114), .S(n8890), .Z(n8892) );
  NOR2_X1 U9928 ( .A1(n9115), .A2(n9114), .ZN(n8891) );
  NOR4_X1 U9929 ( .A1(n8900), .A2(n8899), .A3(n8754), .A4(n8926), .ZN(n8902)
         );
  NAND3_X1 U9930 ( .A1(n8903), .A2(n8902), .A3(n8901), .ZN(n8904) );
  NOR4_X1 U9931 ( .A1(n5053), .A2(n8906), .A3(n8905), .A4(n8904), .ZN(n8907)
         );
  NAND4_X1 U9932 ( .A1(n8910), .A2(n8909), .A3(n8908), .A4(n8907), .ZN(n8911)
         );
  NOR4_X1 U9933 ( .A1(n5067), .A2(n8913), .A3(n8912), .A4(n8911), .ZN(n8914)
         );
  NAND4_X1 U9934 ( .A1(n9347), .A2(n8916), .A3(n8915), .A4(n8914), .ZN(n8917)
         );
  NOR4_X1 U9935 ( .A1(n9336), .A2(n9309), .A3(n5060), .A4(n8917), .ZN(n8918)
         );
  NAND4_X1 U9936 ( .A1(n9133), .A2(n9255), .A3(n9130), .A4(n8918), .ZN(n8919)
         );
  NOR4_X1 U9937 ( .A1(n9140), .A2(n8920), .A3(n9137), .A4(n8919), .ZN(n8921)
         );
  NAND4_X1 U9938 ( .A1(n9170), .A2(n9183), .A3(n9197), .A4(n8921), .ZN(n8922)
         );
  OAI21_X1 U9939 ( .B1(n8935), .B2(n8933), .A(P2_B_REG_SCAN_IN), .ZN(n8934) );
  XNOR2_X1 U9940 ( .A(n8937), .B(n8936), .ZN(n8943) );
  INV_X1 U9941 ( .A(n9180), .ZN(n8938) );
  OAI22_X1 U9942 ( .A1(n8938), .A2(n9044), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10112), .ZN(n8941) );
  OAI22_X1 U9943 ( .A1(n9146), .A2(n9015), .B1(n8991), .B2(n8939), .ZN(n8940)
         );
  AOI211_X1 U9944 ( .C1(n9405), .C2(n10293), .A(n8941), .B(n8940), .ZN(n8942)
         );
  OAI21_X1 U9945 ( .B1(n8943), .B2(n10288), .A(n8942), .ZN(P2_U3216) );
  NOR2_X1 U9946 ( .A1(n9017), .A2(n9264), .ZN(n8947) );
  NOR2_X1 U9947 ( .A1(n10288), .A2(n8944), .ZN(n8946) );
  MUX2_X1 U9948 ( .A(n8947), .B(n8946), .S(n8945), .Z(n8951) );
  INV_X1 U9949 ( .A(n8709), .ZN(n9250) );
  AOI22_X1 U9950 ( .A1(n10284), .A2(n9248), .B1(P2_REG3_REG_23__SCAN_IN), .B2(
        P2_U3152), .ZN(n8949) );
  INV_X1 U9951 ( .A(n9138), .ZN(n9242) );
  AOI22_X1 U9952 ( .A1(n10282), .A2(n9240), .B1(n10281), .B2(n9242), .ZN(n8948) );
  OAI211_X1 U9953 ( .C1(n9250), .C2(n9046), .A(n8949), .B(n8948), .ZN(n8950)
         );
  OR2_X1 U9954 ( .A1(n8951), .A2(n8950), .ZN(P2_U3218) );
  OAI22_X1 U9955 ( .A1(n9274), .A2(n9370), .B1(n9129), .B2(n9371), .ZN(n8952)
         );
  INV_X1 U9956 ( .A(n8952), .ZN(n9322) );
  NAND2_X1 U9957 ( .A1(P2_U3152), .A2(P2_REG3_REG_19__SCAN_IN), .ZN(n9105) );
  NAND2_X1 U9958 ( .A1(n10284), .A2(n9314), .ZN(n8953) );
  OAI211_X1 U9959 ( .C1(n8994), .C2(n9322), .A(n9105), .B(n8953), .ZN(n8964)
         );
  INV_X1 U9960 ( .A(n8959), .ZN(n8955) );
  NOR3_X1 U9961 ( .A1(n8955), .A2(n8954), .A3(n10288), .ZN(n8962) );
  NAND3_X1 U9962 ( .A1(n8957), .A2(n8956), .A3(n9056), .ZN(n8958) );
  OAI21_X1 U9963 ( .B1(n8959), .B2(n10288), .A(n8958), .ZN(n8961) );
  MUX2_X1 U9964 ( .A(n8962), .B(n8961), .S(n8960), .Z(n8963) );
  AOI211_X1 U9965 ( .C1(n9448), .C2(n10293), .A(n8964), .B(n8963), .ZN(n8965)
         );
  INV_X1 U9966 ( .A(n8965), .ZN(P2_U3221) );
  INV_X1 U9967 ( .A(n8966), .ZN(n8967) );
  AOI21_X1 U9968 ( .B1(n8968), .B2(n8967), .A(n10288), .ZN(n8973) );
  NOR3_X1 U9969 ( .A1(n9017), .A2(n8970), .A3(n8969), .ZN(n8972) );
  OAI21_X1 U9970 ( .B1(n8973), .B2(n8972), .A(n8971), .ZN(n8979) );
  AOI22_X1 U9971 ( .A1(n10284), .A2(n8974), .B1(P2_REG3_REG_8__SCAN_IN), .B2(
        P2_U3152), .ZN(n8978) );
  AOI22_X1 U9972 ( .A1(n10282), .A2(n9065), .B1(n10281), .B2(n5120), .ZN(n8977) );
  NAND2_X1 U9973 ( .A1(n10293), .A2(n8975), .ZN(n8976) );
  NAND4_X1 U9974 ( .A1(n8979), .A2(n8978), .A3(n8977), .A4(n8976), .ZN(
        P2_U3223) );
  XNOR2_X1 U9975 ( .A(n8981), .B(n8980), .ZN(n8986) );
  INV_X1 U9976 ( .A(n9436), .ZN(n9287) );
  AOI22_X1 U9977 ( .A1(n10284), .A2(n9284), .B1(P2_REG3_REG_21__SCAN_IN), .B2(
        P2_U3152), .ZN(n8983) );
  INV_X1 U9978 ( .A(n9274), .ZN(n9131) );
  AOI22_X1 U9979 ( .A1(n10282), .A2(n9131), .B1(n10281), .B2(n9240), .ZN(n8982) );
  OAI211_X1 U9980 ( .C1(n9287), .C2(n9046), .A(n8983), .B(n8982), .ZN(n8984)
         );
  INV_X1 U9981 ( .A(n8984), .ZN(n8985) );
  OAI21_X1 U9982 ( .B1(n8986), .B2(n10288), .A(n8985), .ZN(P2_U3225) );
  INV_X1 U9983 ( .A(n8987), .ZN(n8988) );
  AOI21_X1 U9984 ( .B1(n8990), .B2(n8989), .A(n8988), .ZN(n8998) );
  NOR2_X1 U9985 ( .A1(n9044), .A2(n9213), .ZN(n8996) );
  NOR2_X1 U9986 ( .A1(n9138), .A2(n9371), .ZN(n8992) );
  AOI21_X1 U9987 ( .B1(n9186), .B2(n9241), .A(n8992), .ZN(n9209) );
  OAI22_X1 U9988 ( .A1(n9209), .A2(n8994), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n8993), .ZN(n8995) );
  AOI211_X1 U9989 ( .C1(n9417), .C2(n10293), .A(n8996), .B(n8995), .ZN(n8997)
         );
  OAI21_X1 U9990 ( .B1(n8998), .B2(n10288), .A(n8997), .ZN(P2_U3227) );
  NOR2_X1 U9991 ( .A1(n9017), .A2(n9138), .ZN(n9002) );
  NOR2_X1 U9992 ( .A1(n8999), .A2(n10288), .ZN(n9001) );
  MUX2_X1 U9993 ( .A(n9002), .B(n9001), .S(n9000), .Z(n9007) );
  INV_X1 U9994 ( .A(n9003), .ZN(n9224) );
  AOI22_X1 U9995 ( .A1(n10284), .A2(n9224), .B1(P2_REG3_REG_24__SCAN_IN), .B2(
        P2_U3152), .ZN(n9005) );
  INV_X1 U9996 ( .A(n9264), .ZN(n9055) );
  AOI22_X1 U9997 ( .A1(n10282), .A2(n9055), .B1(n10281), .B2(n9054), .ZN(n9004) );
  OAI211_X1 U9998 ( .C1(n9226), .C2(n9046), .A(n9005), .B(n9004), .ZN(n9006)
         );
  OR2_X1 U9999 ( .A1(n9007), .A2(n9006), .ZN(P2_U3231) );
  OAI21_X1 U10000 ( .B1(n8971), .B2(n9019), .A(n9008), .ZN(n9010) );
  NAND2_X1 U10001 ( .A1(n9010), .A2(n9009), .ZN(n9023) );
  NAND2_X1 U10002 ( .A1(n10284), .A2(n9011), .ZN(n9012) );
  OAI211_X1 U10003 ( .C1(n9015), .C2(n9014), .A(n9013), .B(n9012), .ZN(n9016)
         );
  AOI21_X1 U10004 ( .B1(n10605), .B2(n10293), .A(n9016), .ZN(n9022) );
  NOR3_X1 U10005 ( .A1(n9019), .A2(n9018), .A3(n9017), .ZN(n9020) );
  OAI21_X1 U10006 ( .B1(n9020), .B2(n10282), .A(n9064), .ZN(n9021) );
  NAND3_X1 U10007 ( .A1(n9023), .A2(n9022), .A3(n9021), .ZN(P2_U3233) );
  XNOR2_X1 U10008 ( .A(n9025), .B(n9024), .ZN(n9030) );
  INV_X1 U10009 ( .A(n9293), .ZN(n9134) );
  AOI22_X1 U10010 ( .A1(n10282), .A2(n9056), .B1(n10281), .B2(n9134), .ZN(
        n9027) );
  NAND2_X1 U10011 ( .A1(P2_U3152), .A2(P2_REG3_REG_20__SCAN_IN), .ZN(n9026) );
  OAI211_X1 U10012 ( .C1(n9044), .C2(n9301), .A(n9027), .B(n9026), .ZN(n9028)
         );
  AOI21_X1 U10013 ( .B1(n9441), .B2(n10293), .A(n9028), .ZN(n9029) );
  OAI21_X1 U10014 ( .B1(n9030), .B2(n10288), .A(n9029), .ZN(P2_U3235) );
  NAND2_X1 U10015 ( .A1(n9032), .A2(n9031), .ZN(n9033) );
  AOI21_X1 U10016 ( .B1(n9034), .B2(n9033), .A(n10288), .ZN(n9039) );
  INV_X1 U10017 ( .A(n9430), .ZN(n9260) );
  INV_X1 U10018 ( .A(n9035), .ZN(n9258) );
  AOI22_X1 U10019 ( .A1(n10284), .A2(n9258), .B1(P2_REG3_REG_22__SCAN_IN), 
        .B2(P2_U3152), .ZN(n9037) );
  AOI22_X1 U10020 ( .A1(n10282), .A2(n9134), .B1(n10281), .B2(n9055), .ZN(
        n9036) );
  OAI211_X1 U10021 ( .C1(n9260), .C2(n9046), .A(n9037), .B(n9036), .ZN(n9038)
         );
  OR2_X1 U10022 ( .A1(n9039), .A2(n9038), .ZN(P2_U3237) );
  XNOR2_X1 U10023 ( .A(n9040), .B(n9041), .ZN(n9051) );
  OR2_X1 U10024 ( .A1(n9053), .A2(n9370), .ZN(n9043) );
  NAND2_X1 U10025 ( .A1(n9054), .A2(n9239), .ZN(n9042) );
  NAND2_X1 U10026 ( .A1(n9043), .A2(n9042), .ZN(n9200) );
  INV_X1 U10027 ( .A(n9194), .ZN(n9045) );
  OAI22_X1 U10028 ( .A1(n9045), .A2(n9044), .B1(P2_STATE_REG_SCAN_IN), .B2(
        n10272), .ZN(n9048) );
  INV_X1 U10029 ( .A(n9411), .ZN(n9196) );
  NOR2_X1 U10030 ( .A1(n9196), .A2(n9046), .ZN(n9047) );
  AOI211_X1 U10031 ( .C1(n9049), .C2(n9200), .A(n9048), .B(n9047), .ZN(n9050)
         );
  OAI21_X1 U10032 ( .B1(n9051), .B2(n10288), .A(n9050), .ZN(P2_U3242) );
  MUX2_X1 U10033 ( .A(n9052), .B(P2_DATAO_REG_30__SCAN_IN), .S(n9069), .Z(
        P2_U3582) );
  INV_X1 U10034 ( .A(n9053), .ZN(n9143) );
  MUX2_X1 U10035 ( .A(P2_DATAO_REG_27__SCAN_IN), .B(n9143), .S(P2_U3966), .Z(
        P2_U3579) );
  MUX2_X1 U10036 ( .A(n9186), .B(P2_DATAO_REG_26__SCAN_IN), .S(n9069), .Z(
        P2_U3578) );
  MUX2_X1 U10037 ( .A(n9054), .B(P2_DATAO_REG_25__SCAN_IN), .S(n9069), .Z(
        P2_U3577) );
  MUX2_X1 U10038 ( .A(n9242), .B(P2_DATAO_REG_24__SCAN_IN), .S(n9069), .Z(
        P2_U3576) );
  MUX2_X1 U10039 ( .A(P2_DATAO_REG_23__SCAN_IN), .B(n9055), .S(P2_U3966), .Z(
        P2_U3575) );
  MUX2_X1 U10040 ( .A(P2_DATAO_REG_22__SCAN_IN), .B(n9240), .S(P2_U3966), .Z(
        P2_U3574) );
  MUX2_X1 U10041 ( .A(P2_DATAO_REG_21__SCAN_IN), .B(n9134), .S(P2_U3966), .Z(
        P2_U3573) );
  MUX2_X1 U10042 ( .A(n9131), .B(P2_DATAO_REG_20__SCAN_IN), .S(n9069), .Z(
        P2_U3572) );
  MUX2_X1 U10043 ( .A(P2_DATAO_REG_19__SCAN_IN), .B(n9056), .S(P2_U3966), .Z(
        P2_U3571) );
  MUX2_X1 U10044 ( .A(n9057), .B(P2_DATAO_REG_18__SCAN_IN), .S(n9069), .Z(
        P2_U3570) );
  MUX2_X1 U10045 ( .A(P2_DATAO_REG_17__SCAN_IN), .B(n9127), .S(P2_U3966), .Z(
        P2_U3569) );
  INV_X1 U10046 ( .A(n9058), .ZN(n9123) );
  MUX2_X1 U10047 ( .A(P2_DATAO_REG_16__SCAN_IN), .B(n9123), .S(P2_U3966), .Z(
        P2_U3568) );
  MUX2_X1 U10048 ( .A(P2_DATAO_REG_15__SCAN_IN), .B(n9059), .S(P2_U3966), .Z(
        P2_U3567) );
  INV_X1 U10049 ( .A(n9060), .ZN(n10280) );
  MUX2_X1 U10050 ( .A(P2_DATAO_REG_14__SCAN_IN), .B(n10280), .S(P2_U3966), .Z(
        P2_U3566) );
  MUX2_X1 U10051 ( .A(P2_DATAO_REG_13__SCAN_IN), .B(n9061), .S(P2_U3966), .Z(
        P2_U3565) );
  MUX2_X1 U10052 ( .A(P2_DATAO_REG_12__SCAN_IN), .B(n7840), .S(P2_U3966), .Z(
        P2_U3564) );
  MUX2_X1 U10053 ( .A(P2_DATAO_REG_11__SCAN_IN), .B(n9062), .S(P2_U3966), .Z(
        P2_U3563) );
  MUX2_X1 U10054 ( .A(P2_DATAO_REG_10__SCAN_IN), .B(n9063), .S(P2_U3966), .Z(
        P2_U3562) );
  MUX2_X1 U10055 ( .A(P2_DATAO_REG_9__SCAN_IN), .B(n5120), .S(P2_U3966), .Z(
        P2_U3561) );
  MUX2_X1 U10056 ( .A(P2_DATAO_REG_8__SCAN_IN), .B(n9064), .S(P2_U3966), .Z(
        P2_U3560) );
  MUX2_X1 U10057 ( .A(n9065), .B(P2_DATAO_REG_7__SCAN_IN), .S(n9069), .Z(
        P2_U3559) );
  MUX2_X1 U10058 ( .A(P2_DATAO_REG_4__SCAN_IN), .B(n9066), .S(P2_U3966), .Z(
        P2_U3556) );
  MUX2_X1 U10059 ( .A(n9067), .B(P2_DATAO_REG_2__SCAN_IN), .S(n9069), .Z(
        P2_U3554) );
  MUX2_X1 U10060 ( .A(n9068), .B(P2_DATAO_REG_1__SCAN_IN), .S(n9069), .Z(
        P2_U3553) );
  MUX2_X1 U10061 ( .A(n6952), .B(P2_DATAO_REG_0__SCAN_IN), .S(n9069), .Z(
        P2_U3552) );
  OR2_X1 U10062 ( .A1(n9090), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9071) );
  NAND2_X1 U10063 ( .A1(n9090), .A2(P2_REG2_REG_18__SCAN_IN), .ZN(n9070) );
  NAND2_X1 U10064 ( .A1(n9071), .A2(n9070), .ZN(n9076) );
  AOI21_X1 U10065 ( .B1(P2_REG2_REG_17__SCAN_IN), .B2(n9073), .A(n9072), .ZN(
        n9074) );
  INV_X1 U10066 ( .A(n9074), .ZN(n9075) );
  NOR2_X1 U10067 ( .A1(n9076), .A2(n9075), .ZN(n9093) );
  AOI21_X1 U10068 ( .B1(n9076), .B2(n9075), .A(n9093), .ZN(n9092) );
  INV_X1 U10069 ( .A(P2_REG1_REG_17__SCAN_IN), .ZN(n9082) );
  INV_X1 U10070 ( .A(n9077), .ZN(n9079) );
  NAND2_X1 U10071 ( .A1(n9079), .A2(n9078), .ZN(n9080) );
  OAI21_X1 U10072 ( .B1(n9082), .B2(n9081), .A(n9080), .ZN(n9085) );
  INV_X1 U10073 ( .A(n9090), .ZN(n9095) );
  INV_X1 U10074 ( .A(P2_REG1_REG_18__SCAN_IN), .ZN(n9083) );
  NAND2_X1 U10075 ( .A1(n9095), .A2(n9083), .ZN(n9099) );
  OAI21_X1 U10076 ( .B1(n9095), .B2(n9083), .A(n9099), .ZN(n9084) );
  NOR2_X1 U10077 ( .A1(n9084), .A2(n9085), .ZN(n9101) );
  AOI21_X1 U10078 ( .B1(n9085), .B2(n9084), .A(n9101), .ZN(n9088) );
  NAND2_X1 U10079 ( .A1(n10486), .A2(P2_ADDR_REG_18__SCAN_IN), .ZN(n9086) );
  OAI211_X1 U10080 ( .C1(n10481), .C2(n9088), .A(n9087), .B(n9086), .ZN(n9089)
         );
  AOI21_X1 U10081 ( .B1(n9090), .B2(n10478), .A(n9089), .ZN(n9091) );
  OAI21_X1 U10082 ( .B1(n9092), .B2(n10415), .A(n9091), .ZN(P2_U3263) );
  INV_X1 U10083 ( .A(P2_REG2_REG_18__SCAN_IN), .ZN(n9094) );
  AOI21_X1 U10084 ( .B1(n9095), .B2(n9094), .A(n9093), .ZN(n9098) );
  INV_X1 U10085 ( .A(P2_REG2_REG_19__SCAN_IN), .ZN(n9096) );
  MUX2_X1 U10086 ( .A(P2_REG2_REG_19__SCAN_IN), .B(n9096), .S(n9317), .Z(n9097) );
  XNOR2_X1 U10087 ( .A(n9098), .B(n9097), .ZN(n9109) );
  INV_X1 U10088 ( .A(n9099), .ZN(n9100) );
  NOR2_X1 U10089 ( .A1(n9101), .A2(n9100), .ZN(n9103) );
  XNOR2_X1 U10090 ( .A(n5298), .B(P2_REG1_REG_19__SCAN_IN), .ZN(n9102) );
  XNOR2_X1 U10091 ( .A(n9103), .B(n9102), .ZN(n9106) );
  NAND2_X1 U10092 ( .A1(n10486), .A2(P2_ADDR_REG_19__SCAN_IN), .ZN(n9104) );
  OAI211_X1 U10093 ( .C1(n10481), .C2(n9106), .A(n9105), .B(n9104), .ZN(n9107)
         );
  AOI21_X1 U10094 ( .B1(n9317), .B2(n10478), .A(n9107), .ZN(n9108) );
  OAI21_X1 U10095 ( .B1(n10415), .B2(n9109), .A(n9108), .ZN(P2_U3264) );
  NOR2_X2 U10096 ( .A1(n9441), .A2(n9312), .ZN(n9298) );
  NAND2_X1 U10097 ( .A1(n9287), .A2(n9298), .ZN(n9283) );
  OR2_X2 U10098 ( .A1(n9430), .A2(n9283), .ZN(n9256) );
  OR2_X2 U10099 ( .A1(n9150), .A2(n9111), .ZN(n9151) );
  XNOR2_X1 U10100 ( .A(n9118), .B(n9115), .ZN(n9388) );
  NAND2_X1 U10101 ( .A1(n9112), .A2(P2_B_REG_SCAN_IN), .ZN(n9113) );
  NAND2_X1 U10102 ( .A1(n9241), .A2(n9113), .ZN(n9149) );
  NOR2_X1 U10103 ( .A1(n9114), .A2(n9149), .ZN(n9385) );
  INV_X1 U10104 ( .A(n9385), .ZN(n9391) );
  NOR2_X1 U10105 ( .A1(n9268), .A2(n9391), .ZN(n9120) );
  NOR2_X1 U10106 ( .A1(n9115), .A2(n9333), .ZN(n9116) );
  AOI211_X1 U10107 ( .C1(n9268), .C2(P2_REG2_REG_31__SCAN_IN), .A(n9120), .B(
        n9116), .ZN(n9117) );
  OAI21_X1 U10108 ( .B1(n9388), .B2(n9152), .A(n9117), .ZN(P2_U3265) );
  INV_X1 U10109 ( .A(n9118), .ZN(n9390) );
  NAND2_X1 U10110 ( .A1(n9151), .A2(n9119), .ZN(n9389) );
  NAND3_X1 U10111 ( .A1(n9390), .A2(n9380), .A3(n9389), .ZN(n9122) );
  AOI21_X1 U10112 ( .B1(n9268), .B2(P2_REG2_REG_30__SCAN_IN), .A(n9120), .ZN(
        n9121) );
  OAI211_X1 U10113 ( .C1(n9393), .C2(n9333), .A(n9122), .B(n9121), .ZN(
        P2_U3266) );
  INV_X1 U10114 ( .A(n9457), .ZN(n9128) );
  INV_X1 U10115 ( .A(n9451), .ZN(n9334) );
  NAND2_X1 U10116 ( .A1(n9254), .A2(n9262), .ZN(n9136) );
  NAND2_X1 U10117 ( .A1(n9260), .A2(n9275), .ZN(n9135) );
  NAND2_X1 U10118 ( .A1(n9136), .A2(n9135), .ZN(n9246) );
  NAND2_X1 U10119 ( .A1(n9226), .A2(n9138), .ZN(n9139) );
  INV_X1 U10120 ( .A(n9417), .ZN(n9217) );
  NOR2_X1 U10121 ( .A1(n9411), .A2(n9186), .ZN(n9142) );
  NAND2_X1 U10122 ( .A1(n9411), .A2(n9186), .ZN(n9141) );
  INV_X1 U10123 ( .A(n9394), .ZN(n9159) );
  XNOR2_X1 U10124 ( .A(n9145), .B(n9144), .ZN(n9147) );
  OAI222_X1 U10125 ( .A1(n9149), .A2(n9148), .B1(n9147), .B2(n9376), .C1(n9371), .C2(n9146), .ZN(n9395) );
  INV_X1 U10126 ( .A(n9111), .ZN(n9155) );
  INV_X1 U10127 ( .A(n9150), .ZN(n9165) );
  OAI21_X1 U10128 ( .B1(n9155), .B2(n9165), .A(n9151), .ZN(n9396) );
  NOR2_X1 U10129 ( .A1(n9396), .A2(n9152), .ZN(n9157) );
  AOI22_X1 U10130 ( .A1(n9153), .A2(n9377), .B1(P2_REG2_REG_29__SCAN_IN), .B2(
        n9268), .ZN(n9154) );
  OAI21_X1 U10131 ( .B1(n9155), .B2(n9333), .A(n9154), .ZN(n9156) );
  AOI211_X1 U10132 ( .C1(n9395), .C2(n9378), .A(n9157), .B(n9156), .ZN(n9158)
         );
  OAI21_X1 U10133 ( .B1(n9159), .B2(n9359), .A(n9158), .ZN(P2_U3267) );
  OAI21_X1 U10134 ( .B1(n9160), .B2(n9162), .A(n9161), .ZN(n9163) );
  INV_X1 U10135 ( .A(n9163), .ZN(n9404) );
  AOI21_X1 U10136 ( .B1(n9400), .B2(n9179), .A(n9165), .ZN(n9401) );
  AOI22_X1 U10137 ( .A1(n9166), .A2(n9377), .B1(P2_REG2_REG_28__SCAN_IN), .B2(
        n9268), .ZN(n9167) );
  OAI21_X1 U10138 ( .B1(n9168), .B2(n9333), .A(n9167), .ZN(n9175) );
  OAI21_X1 U10139 ( .B1(n9171), .B2(n9170), .A(n9169), .ZN(n9173) );
  AOI21_X1 U10140 ( .B1(n9173), .B2(n9349), .A(n9172), .ZN(n9403) );
  NOR2_X1 U10141 ( .A1(n9403), .A2(n9268), .ZN(n9174) );
  AOI211_X1 U10142 ( .C1(n9401), .C2(n9380), .A(n9175), .B(n9174), .ZN(n9176)
         );
  OAI21_X1 U10143 ( .B1(n9404), .B2(n9359), .A(n9176), .ZN(P2_U3268) );
  XNOR2_X1 U10144 ( .A(n9177), .B(n9178), .ZN(n9409) );
  AOI21_X1 U10145 ( .B1(n9405), .B2(n9191), .A(n9164), .ZN(n9406) );
  INV_X1 U10146 ( .A(n9405), .ZN(n9182) );
  AOI22_X1 U10147 ( .A1(n9180), .A2(n9377), .B1(P2_REG2_REG_27__SCAN_IN), .B2(
        n9268), .ZN(n9181) );
  OAI21_X1 U10148 ( .B1(n9182), .B2(n9333), .A(n9181), .ZN(n9188) );
  NOR2_X1 U10149 ( .A1(n9408), .A2(n9268), .ZN(n9187) );
  AOI211_X1 U10150 ( .C1(n9380), .C2(n9406), .A(n9188), .B(n9187), .ZN(n9189)
         );
  OAI21_X1 U10151 ( .B1(n9409), .B2(n9359), .A(n9189), .ZN(P2_U3269) );
  XNOR2_X1 U10152 ( .A(n9190), .B(n9197), .ZN(n9414) );
  INV_X1 U10153 ( .A(n9211), .ZN(n9193) );
  INV_X1 U10154 ( .A(n9191), .ZN(n9192) );
  AOI211_X1 U10155 ( .C1(n9411), .C2(n9193), .A(n10693), .B(n9192), .ZN(n9410)
         );
  AOI22_X1 U10156 ( .A1(n9194), .A2(n9377), .B1(n9268), .B2(
        P2_REG2_REG_26__SCAN_IN), .ZN(n9195) );
  OAI21_X1 U10157 ( .B1(n9196), .B2(n9333), .A(n9195), .ZN(n9203) );
  XNOR2_X1 U10158 ( .A(n9199), .B(n9198), .ZN(n9201) );
  AOI21_X1 U10159 ( .B1(n9201), .B2(n9349), .A(n9200), .ZN(n9413) );
  NOR2_X1 U10160 ( .A1(n9413), .A2(n9268), .ZN(n9202) );
  AOI211_X1 U10161 ( .C1(n9410), .C2(n9362), .A(n9203), .B(n9202), .ZN(n9204)
         );
  OAI21_X1 U10162 ( .B1(n9414), .B2(n9359), .A(n9204), .ZN(P2_U3270) );
  XNOR2_X1 U10163 ( .A(n9205), .B(n9207), .ZN(n9419) );
  OAI211_X1 U10164 ( .C1(n9208), .C2(n9207), .A(n9206), .B(n9349), .ZN(n9210)
         );
  NAND2_X1 U10165 ( .A1(n9210), .A2(n9209), .ZN(n9416) );
  AOI211_X1 U10166 ( .C1(n9417), .C2(n9212), .A(n10693), .B(n9211), .ZN(n9415)
         );
  NAND2_X1 U10167 ( .A1(n9415), .A2(n9362), .ZN(n9216) );
  INV_X1 U10168 ( .A(n9213), .ZN(n9214) );
  AOI22_X1 U10169 ( .A1(n9268), .A2(P2_REG2_REG_25__SCAN_IN), .B1(n9214), .B2(
        n9377), .ZN(n9215) );
  OAI211_X1 U10170 ( .C1(n9217), .C2(n9333), .A(n9216), .B(n9215), .ZN(n9218)
         );
  AOI21_X1 U10171 ( .B1(n9378), .B2(n9416), .A(n9218), .ZN(n9219) );
  OAI21_X1 U10172 ( .B1(n9419), .B2(n9359), .A(n9219), .ZN(P2_U3271) );
  INV_X1 U10173 ( .A(n9220), .ZN(n9221) );
  AOI21_X1 U10174 ( .B1(n9229), .B2(n9222), .A(n9221), .ZN(n9424) );
  XNOR2_X1 U10175 ( .A(n9226), .B(n9247), .ZN(n9421) );
  AOI22_X1 U10176 ( .A1(n9268), .A2(P2_REG2_REG_24__SCAN_IN), .B1(n9224), .B2(
        n9377), .ZN(n9225) );
  OAI21_X1 U10177 ( .B1(n9226), .B2(n9333), .A(n9225), .ZN(n9237) );
  INV_X1 U10178 ( .A(n9227), .ZN(n9232) );
  AOI21_X1 U10179 ( .B1(n9228), .B2(n9230), .A(n9229), .ZN(n9231) );
  NOR3_X1 U10180 ( .A1(n9232), .A2(n9231), .A3(n9376), .ZN(n9235) );
  OAI22_X1 U10181 ( .A1(n9233), .A2(n9370), .B1(n9264), .B2(n9371), .ZN(n9234)
         );
  NOR2_X1 U10182 ( .A1(n9235), .A2(n9234), .ZN(n9423) );
  NOR2_X1 U10183 ( .A1(n9423), .A2(n9268), .ZN(n9236) );
  AOI211_X1 U10184 ( .C1(n9421), .C2(n9380), .A(n9237), .B(n9236), .ZN(n9238)
         );
  OAI21_X1 U10185 ( .B1(n9424), .B2(n9359), .A(n9238), .ZN(P2_U3272) );
  OAI21_X1 U10186 ( .B1(n4927), .B2(n9245), .A(n9228), .ZN(n9243) );
  AOI222_X1 U10187 ( .A1(n9349), .A2(n9243), .B1(n9242), .B2(n9241), .C1(n9240), .C2(n9239), .ZN(n9428) );
  NAND2_X1 U10188 ( .A1(n9246), .A2(n9245), .ZN(n9425) );
  NAND3_X1 U10189 ( .A1(n9244), .A2(n9425), .A3(n9289), .ZN(n9253) );
  AOI21_X1 U10190 ( .B1(n8709), .B2(n9256), .A(n9223), .ZN(n9426) );
  AOI22_X1 U10191 ( .A1(n9268), .A2(P2_REG2_REG_23__SCAN_IN), .B1(n9248), .B2(
        n9377), .ZN(n9249) );
  OAI21_X1 U10192 ( .B1(n9250), .B2(n9333), .A(n9249), .ZN(n9251) );
  AOI21_X1 U10193 ( .B1(n9426), .B2(n9380), .A(n9251), .ZN(n9252) );
  OAI211_X1 U10194 ( .C1(n9268), .C2(n9428), .A(n9253), .B(n9252), .ZN(
        P2_U3273) );
  XNOR2_X1 U10195 ( .A(n9254), .B(n9255), .ZN(n9434) );
  INV_X1 U10196 ( .A(n9256), .ZN(n9257) );
  AOI21_X1 U10197 ( .B1(n9430), .B2(n9283), .A(n9257), .ZN(n9431) );
  AOI22_X1 U10198 ( .A1(n9268), .A2(P2_REG2_REG_22__SCAN_IN), .B1(n9258), .B2(
        n9377), .ZN(n9259) );
  OAI21_X1 U10199 ( .B1(n9260), .B2(n9333), .A(n9259), .ZN(n9270) );
  INV_X1 U10200 ( .A(n9261), .ZN(n9263) );
  AOI21_X1 U10201 ( .B1(n9263), .B2(n9262), .A(n9376), .ZN(n9267) );
  OAI22_X1 U10202 ( .A1(n9264), .A2(n9370), .B1(n9293), .B2(n9371), .ZN(n9265)
         );
  AOI21_X1 U10203 ( .B1(n9267), .B2(n9266), .A(n9265), .ZN(n9433) );
  NOR2_X1 U10204 ( .A1(n9433), .A2(n9268), .ZN(n9269) );
  AOI211_X1 U10205 ( .C1(n9431), .C2(n9380), .A(n9270), .B(n9269), .ZN(n9271)
         );
  OAI21_X1 U10206 ( .B1(n9434), .B2(n9359), .A(n9271), .ZN(P2_U3274) );
  INV_X1 U10207 ( .A(n9272), .ZN(n9273) );
  AOI21_X1 U10208 ( .B1(n9273), .B2(n9280), .A(n9376), .ZN(n9278) );
  OAI22_X1 U10209 ( .A1(n9275), .A2(n9370), .B1(n9274), .B2(n9371), .ZN(n9276)
         );
  AOI21_X1 U10210 ( .B1(n9278), .B2(n9277), .A(n9276), .ZN(n9439) );
  OAI21_X1 U10211 ( .B1(n9281), .B2(n9280), .A(n9279), .ZN(n9435) );
  OR2_X1 U10212 ( .A1(n9287), .A2(n9298), .ZN(n9282) );
  AND2_X1 U10213 ( .A1(n9283), .A2(n9282), .ZN(n9437) );
  NAND2_X1 U10214 ( .A1(n9437), .A2(n9380), .ZN(n9286) );
  AOI22_X1 U10215 ( .A1(n9268), .A2(P2_REG2_REG_21__SCAN_IN), .B1(n9284), .B2(
        n9377), .ZN(n9285) );
  OAI211_X1 U10216 ( .C1(n9287), .C2(n9333), .A(n9286), .B(n9285), .ZN(n9288)
         );
  AOI21_X1 U10217 ( .B1(n9435), .B2(n9289), .A(n9288), .ZN(n9290) );
  OAI21_X1 U10218 ( .B1(n9268), .B2(n9439), .A(n9290), .ZN(P2_U3275) );
  INV_X1 U10219 ( .A(n9291), .ZN(n9292) );
  AOI21_X1 U10220 ( .B1(n9292), .B2(n9303), .A(n9376), .ZN(n9296) );
  OAI22_X1 U10221 ( .A1(n9293), .A2(n9370), .B1(n9339), .B2(n9371), .ZN(n9294)
         );
  AOI21_X1 U10222 ( .B1(n9296), .B2(n9295), .A(n9294), .ZN(n9444) );
  AND2_X1 U10223 ( .A1(n9441), .A2(n9312), .ZN(n9297) );
  NOR2_X1 U10224 ( .A1(n9298), .A2(n9297), .ZN(n9442) );
  NAND2_X1 U10225 ( .A1(n9441), .A2(n9366), .ZN(n9300) );
  NAND2_X1 U10226 ( .A1(n9268), .A2(P2_REG2_REG_20__SCAN_IN), .ZN(n9299) );
  OAI211_X1 U10227 ( .C1(n9316), .C2(n9301), .A(n9300), .B(n9299), .ZN(n9306)
         );
  OAI21_X1 U10228 ( .B1(n9304), .B2(n9303), .A(n5468), .ZN(n9445) );
  NOR2_X1 U10229 ( .A1(n9445), .A2(n9359), .ZN(n9305) );
  AOI211_X1 U10230 ( .C1(n9442), .C2(n9380), .A(n9306), .B(n9305), .ZN(n9307)
         );
  OAI21_X1 U10231 ( .B1(n9268), .B2(n9444), .A(n9307), .ZN(P2_U3276) );
  OAI21_X1 U10232 ( .B1(n9310), .B2(n9309), .A(n9308), .ZN(n9450) );
  AOI22_X1 U10233 ( .A1(n9448), .A2(n9366), .B1(P2_REG2_REG_19__SCAN_IN), .B2(
        n9268), .ZN(n9326) );
  INV_X1 U10234 ( .A(n9312), .ZN(n9313) );
  AOI211_X1 U10235 ( .C1(n9448), .C2(n5210), .A(n10693), .B(n9313), .ZN(n9447)
         );
  INV_X1 U10236 ( .A(n9447), .ZN(n9318) );
  INV_X1 U10237 ( .A(n9314), .ZN(n9315) );
  OAI22_X1 U10238 ( .A1(n9318), .A2(n9317), .B1(n9316), .B2(n9315), .ZN(n9324)
         );
  OAI211_X1 U10239 ( .C1(n9321), .C2(n9320), .A(n9319), .B(n9349), .ZN(n9323)
         );
  NAND2_X1 U10240 ( .A1(n9323), .A2(n9322), .ZN(n9446) );
  OAI21_X1 U10241 ( .B1(n9324), .B2(n9446), .A(n9378), .ZN(n9325) );
  OAI211_X1 U10242 ( .C1(n9450), .C2(n9359), .A(n9326), .B(n9325), .ZN(
        P2_U3277) );
  XNOR2_X1 U10243 ( .A(n9327), .B(n9328), .ZN(n9455) );
  AOI21_X1 U10244 ( .B1(n9451), .B2(n9329), .A(n9311), .ZN(n9452) );
  INV_X1 U10245 ( .A(n9330), .ZN(n9331) );
  AOI22_X1 U10246 ( .A1(n9268), .A2(P2_REG2_REG_18__SCAN_IN), .B1(n9331), .B2(
        n9377), .ZN(n9332) );
  OAI21_X1 U10247 ( .B1(n9334), .B2(n9333), .A(n9332), .ZN(n9344) );
  INV_X1 U10248 ( .A(n9335), .ZN(n9337) );
  AOI21_X1 U10249 ( .B1(n9337), .B2(n9336), .A(n9376), .ZN(n9342) );
  OAI22_X1 U10250 ( .A1(n9339), .A2(n9370), .B1(n9338), .B2(n9371), .ZN(n9340)
         );
  AOI21_X1 U10251 ( .B1(n9342), .B2(n9341), .A(n9340), .ZN(n9454) );
  NOR2_X1 U10252 ( .A1(n9454), .A2(n9268), .ZN(n9343) );
  AOI211_X1 U10253 ( .C1(n9452), .C2(n9380), .A(n9344), .B(n9343), .ZN(n9345)
         );
  OAI21_X1 U10254 ( .B1(n9455), .B2(n9359), .A(n9345), .ZN(P2_U3278) );
  XNOR2_X1 U10255 ( .A(n9346), .B(n9347), .ZN(n9350) );
  AOI21_X1 U10256 ( .B1(n9350), .B2(n9349), .A(n9348), .ZN(n9460) );
  XNOR2_X1 U10257 ( .A(n9351), .B(n9457), .ZN(n9352) );
  NOR2_X1 U10258 ( .A1(n9352), .A2(n10693), .ZN(n9456) );
  NAND2_X1 U10259 ( .A1(n9457), .A2(n9366), .ZN(n9355) );
  NAND2_X1 U10260 ( .A1(n9377), .A2(n9353), .ZN(n9354) );
  OAI211_X1 U10261 ( .C1(n9378), .C2(n7975), .A(n9355), .B(n9354), .ZN(n9361)
         );
  OAI21_X1 U10262 ( .B1(n9357), .B2(n5446), .A(n9356), .ZN(n9358) );
  INV_X1 U10263 ( .A(n9358), .ZN(n9461) );
  NOR2_X1 U10264 ( .A1(n9461), .A2(n9359), .ZN(n9360) );
  AOI211_X1 U10265 ( .C1(n9456), .C2(n9362), .A(n9361), .B(n9360), .ZN(n9363)
         );
  OAI21_X1 U10266 ( .B1(n9268), .B2(n9460), .A(n9363), .ZN(P2_U3279) );
  OAI21_X1 U10267 ( .B1(n9365), .B2(n8754), .A(n9364), .ZN(n10524) );
  AOI22_X1 U10268 ( .A1(n9367), .A2(n10524), .B1(n9366), .B2(n6257), .ZN(n9384) );
  XNOR2_X1 U10269 ( .A(n8758), .B(n9368), .ZN(n9375) );
  INV_X1 U10270 ( .A(n9369), .ZN(n9373) );
  OAI22_X1 U10271 ( .A1(n5424), .A2(n9371), .B1(n5157), .B2(n9370), .ZN(n9372)
         );
  AOI21_X1 U10272 ( .B1(n10524), .B2(n9373), .A(n9372), .ZN(n9374) );
  OAI21_X1 U10273 ( .B1(n9376), .B2(n9375), .A(n9374), .ZN(n10522) );
  AOI22_X1 U10274 ( .A1(n9378), .A2(n10522), .B1(P2_REG3_REG_2__SCAN_IN), .B2(
        n9377), .ZN(n9383) );
  NAND2_X1 U10275 ( .A1(n9379), .A2(n6257), .ZN(n10518) );
  NAND3_X1 U10276 ( .A1(n9380), .A2(n10519), .A3(n10518), .ZN(n9382) );
  NAND2_X1 U10277 ( .A1(n9268), .A2(P2_REG2_REG_2__SCAN_IN), .ZN(n9381) );
  NAND4_X1 U10278 ( .A1(n9384), .A2(n9383), .A3(n9382), .A4(n9381), .ZN(
        P2_U3294) );
  AOI21_X1 U10279 ( .B1(n9386), .B2(n9458), .A(n9385), .ZN(n9387) );
  OAI21_X1 U10280 ( .B1(n9388), .B2(n10693), .A(n9387), .ZN(n9468) );
  MUX2_X1 U10281 ( .A(P2_REG1_REG_31__SCAN_IN), .B(n9468), .S(n10701), .Z(
        P2_U3551) );
  NAND3_X1 U10282 ( .A1(n9390), .A2(n5299), .A3(n9389), .ZN(n9392) );
  OAI211_X1 U10283 ( .C1(n9393), .C2(n10691), .A(n9392), .B(n9391), .ZN(n9469)
         );
  INV_X2 U10284 ( .A(n10699), .ZN(n10701) );
  MUX2_X1 U10285 ( .A(P2_REG1_REG_30__SCAN_IN), .B(n9469), .S(n10701), .Z(
        P2_U3550) );
  NAND2_X1 U10286 ( .A1(n9394), .A2(n10697), .ZN(n9399) );
  INV_X1 U10287 ( .A(n9395), .ZN(n9398) );
  AOI22_X1 U10288 ( .A1(n9401), .A2(n5299), .B1(n9458), .B2(n9400), .ZN(n9402)
         );
  OAI211_X1 U10289 ( .C1(n9404), .C2(n10673), .A(n9403), .B(n9402), .ZN(n9471)
         );
  MUX2_X1 U10290 ( .A(P2_REG1_REG_28__SCAN_IN), .B(n9471), .S(n10701), .Z(
        P2_U3548) );
  AOI22_X1 U10291 ( .A1(n9406), .A2(n5299), .B1(n9458), .B2(n9405), .ZN(n9407)
         );
  OAI211_X1 U10292 ( .C1(n9409), .C2(n10673), .A(n9408), .B(n9407), .ZN(n9472)
         );
  MUX2_X1 U10293 ( .A(P2_REG1_REG_27__SCAN_IN), .B(n9472), .S(n10701), .Z(
        P2_U3547) );
  AOI21_X1 U10294 ( .B1(n9458), .B2(n9411), .A(n9410), .ZN(n9412) );
  OAI211_X1 U10295 ( .C1(n9414), .C2(n10673), .A(n9413), .B(n9412), .ZN(n9473)
         );
  MUX2_X1 U10296 ( .A(P2_REG1_REG_26__SCAN_IN), .B(n9473), .S(n10701), .Z(
        P2_U3546) );
  AOI211_X1 U10297 ( .C1(n9458), .C2(n9417), .A(n9416), .B(n9415), .ZN(n9418)
         );
  OAI21_X1 U10298 ( .B1(n9419), .B2(n10673), .A(n9418), .ZN(n9474) );
  MUX2_X1 U10299 ( .A(P2_REG1_REG_25__SCAN_IN), .B(n9474), .S(n10701), .Z(
        P2_U3545) );
  AOI22_X1 U10300 ( .A1(n9421), .A2(n5299), .B1(n9458), .B2(n9420), .ZN(n9422)
         );
  OAI211_X1 U10301 ( .C1(n9424), .C2(n10673), .A(n9423), .B(n9422), .ZN(n9475)
         );
  MUX2_X1 U10302 ( .A(P2_REG1_REG_24__SCAN_IN), .B(n9475), .S(n10701), .Z(
        P2_U3544) );
  NAND3_X1 U10303 ( .A1(n9244), .A2(n9425), .A3(n10697), .ZN(n9429) );
  AOI22_X1 U10304 ( .A1(n9426), .A2(n5299), .B1(n9458), .B2(n8709), .ZN(n9427)
         );
  NAND3_X1 U10305 ( .A1(n9429), .A2(n9428), .A3(n9427), .ZN(n9476) );
  MUX2_X1 U10306 ( .A(P2_REG1_REG_23__SCAN_IN), .B(n9476), .S(n10701), .Z(
        P2_U3543) );
  AOI22_X1 U10307 ( .A1(n9431), .A2(n5299), .B1(n9458), .B2(n9430), .ZN(n9432)
         );
  OAI211_X1 U10308 ( .C1(n9434), .C2(n10673), .A(n9433), .B(n9432), .ZN(n9477)
         );
  MUX2_X1 U10309 ( .A(P2_REG1_REG_22__SCAN_IN), .B(n9477), .S(n10701), .Z(
        P2_U3542) );
  INV_X1 U10310 ( .A(n9435), .ZN(n9440) );
  AOI22_X1 U10311 ( .A1(n9437), .A2(n5299), .B1(n9458), .B2(n9436), .ZN(n9438)
         );
  OAI211_X1 U10312 ( .C1(n9440), .C2(n10673), .A(n9439), .B(n9438), .ZN(n9478)
         );
  MUX2_X1 U10313 ( .A(P2_REG1_REG_21__SCAN_IN), .B(n9478), .S(n10701), .Z(
        P2_U3541) );
  AOI22_X1 U10314 ( .A1(n9442), .A2(n5299), .B1(n9458), .B2(n9441), .ZN(n9443)
         );
  OAI211_X1 U10315 ( .C1(n9445), .C2(n10673), .A(n9444), .B(n9443), .ZN(n9479)
         );
  MUX2_X1 U10316 ( .A(P2_REG1_REG_20__SCAN_IN), .B(n9479), .S(n10701), .Z(
        P2_U3540) );
  AOI211_X1 U10317 ( .C1(n9458), .C2(n9448), .A(n9447), .B(n9446), .ZN(n9449)
         );
  OAI21_X1 U10318 ( .B1(n9450), .B2(n10673), .A(n9449), .ZN(n9480) );
  MUX2_X1 U10319 ( .A(P2_REG1_REG_19__SCAN_IN), .B(n9480), .S(n10701), .Z(
        P2_U3539) );
  AOI22_X1 U10320 ( .A1(n9452), .A2(n5299), .B1(n9458), .B2(n9451), .ZN(n9453)
         );
  OAI211_X1 U10321 ( .C1(n9455), .C2(n10673), .A(n9454), .B(n9453), .ZN(n9481)
         );
  MUX2_X1 U10322 ( .A(P2_REG1_REG_18__SCAN_IN), .B(n9481), .S(n10701), .Z(
        P2_U3538) );
  AOI21_X1 U10323 ( .B1(n9458), .B2(n9457), .A(n9456), .ZN(n9459) );
  OAI211_X1 U10324 ( .C1(n9461), .C2(n10673), .A(n9460), .B(n9459), .ZN(n9482)
         );
  MUX2_X1 U10325 ( .A(P2_REG1_REG_17__SCAN_IN), .B(n9482), .S(n10701), .Z(
        P2_U3537) );
  OAI21_X1 U10326 ( .B1(n9463), .B2(n10691), .A(n9462), .ZN(n9464) );
  AOI211_X1 U10327 ( .C1(n9466), .C2(n10697), .A(n9465), .B(n9464), .ZN(n9467)
         );
  INV_X1 U10328 ( .A(n9467), .ZN(n9483) );
  MUX2_X1 U10329 ( .A(P2_REG1_REG_16__SCAN_IN), .B(n9483), .S(n10701), .Z(
        P2_U3536) );
  MUX2_X1 U10330 ( .A(P2_REG0_REG_31__SCAN_IN), .B(n9468), .S(n10613), .Z(
        P2_U3519) );
  MUX2_X1 U10331 ( .A(P2_REG0_REG_30__SCAN_IN), .B(n9469), .S(n10613), .Z(
        P2_U3518) );
  MUX2_X1 U10332 ( .A(P2_REG0_REG_29__SCAN_IN), .B(n9470), .S(n10613), .Z(
        P2_U3517) );
  MUX2_X1 U10333 ( .A(P2_REG0_REG_28__SCAN_IN), .B(n9471), .S(n10613), .Z(
        P2_U3516) );
  MUX2_X1 U10334 ( .A(P2_REG0_REG_27__SCAN_IN), .B(n9472), .S(n10613), .Z(
        P2_U3515) );
  MUX2_X1 U10335 ( .A(P2_REG0_REG_26__SCAN_IN), .B(n9473), .S(n10613), .Z(
        P2_U3514) );
  MUX2_X1 U10336 ( .A(P2_REG0_REG_25__SCAN_IN), .B(n9474), .S(n10613), .Z(
        P2_U3513) );
  MUX2_X1 U10337 ( .A(P2_REG0_REG_24__SCAN_IN), .B(n9475), .S(n10613), .Z(
        P2_U3512) );
  MUX2_X1 U10338 ( .A(P2_REG0_REG_23__SCAN_IN), .B(n9476), .S(n10613), .Z(
        P2_U3511) );
  MUX2_X1 U10339 ( .A(P2_REG0_REG_22__SCAN_IN), .B(n9477), .S(n10613), .Z(
        P2_U3510) );
  MUX2_X1 U10340 ( .A(P2_REG0_REG_21__SCAN_IN), .B(n9478), .S(n10613), .Z(
        P2_U3509) );
  MUX2_X1 U10341 ( .A(P2_REG0_REG_20__SCAN_IN), .B(n9479), .S(n10613), .Z(
        P2_U3508) );
  MUX2_X1 U10342 ( .A(P2_REG0_REG_19__SCAN_IN), .B(n9480), .S(n10613), .Z(
        P2_U3507) );
  MUX2_X1 U10343 ( .A(P2_REG0_REG_18__SCAN_IN), .B(n9481), .S(n10613), .Z(
        P2_U3505) );
  MUX2_X1 U10344 ( .A(P2_REG0_REG_17__SCAN_IN), .B(n9482), .S(n10613), .Z(
        P2_U3502) );
  MUX2_X1 U10345 ( .A(P2_REG0_REG_16__SCAN_IN), .B(n9483), .S(n10613), .Z(
        P2_U3499) );
  INV_X1 U10346 ( .A(n8727), .ZN(n10034) );
  NOR4_X1 U10347 ( .A1(n9485), .A2(P2_IR_REG_30__SCAN_IN), .A3(P2_U3152), .A4(
        n9484), .ZN(n9486) );
  AOI21_X1 U10348 ( .B1(n9487), .B2(P1_DATAO_REG_31__SCAN_IN), .A(n9486), .ZN(
        n9488) );
  OAI21_X1 U10349 ( .B1(n10034), .B2(n4857), .A(n9488), .ZN(P2_U3327) );
  INV_X1 U10350 ( .A(n9490), .ZN(n10042) );
  OAI222_X1 U10351 ( .A1(P2_U3152), .A2(n9489), .B1(n4857), .B2(n10042), .C1(
        n9492), .C2(n9491), .ZN(P2_U3329) );
  INV_X1 U10352 ( .A(n9493), .ZN(n9494) );
  MUX2_X1 U10353 ( .A(P2_IR_REG_0__SCAN_IN), .B(n9494), .S(P2_U3152), .Z(
        P2_U3358) );
  INV_X1 U10354 ( .A(n9495), .ZN(n9496) );
  NOR2_X1 U10355 ( .A1(n9497), .A2(n9496), .ZN(n9499) );
  XNOR2_X1 U10356 ( .A(n9499), .B(n9498), .ZN(n9504) );
  AOI22_X1 U10357 ( .A1(n9601), .A2(n9754), .B1(P1_REG3_REG_23__SCAN_IN), .B2(
        P1_U3084), .ZN(n9501) );
  NAND2_X1 U10358 ( .A1(n9602), .A2(n9786), .ZN(n9500) );
  OAI211_X1 U10359 ( .C1(n9782), .C2(n9605), .A(n9501), .B(n9500), .ZN(n9502)
         );
  AOI21_X1 U10360 ( .B1(n9939), .B2(n9607), .A(n9502), .ZN(n9503) );
  OAI21_X1 U10361 ( .B1(n9504), .B2(n9609), .A(n9503), .ZN(P1_U3214) );
  OAI21_X1 U10362 ( .B1(n9507), .B2(n9505), .A(n9506), .ZN(n9508) );
  NAND2_X1 U10363 ( .A1(n9508), .A2(n9590), .ZN(n9512) );
  NOR2_X1 U10364 ( .A1(n9593), .A2(n9839), .ZN(n9510) );
  NAND2_X1 U10365 ( .A1(P1_U3084), .A2(P1_REG3_REG_19__SCAN_IN), .ZN(n9690) );
  OAI21_X1 U10366 ( .B1(n9605), .B2(n9882), .A(n9690), .ZN(n9509) );
  AOI211_X1 U10367 ( .C1(n9601), .C2(n9810), .A(n9510), .B(n9509), .ZN(n9511)
         );
  OAI211_X1 U10368 ( .C1(n9513), .C2(n9598), .A(n9512), .B(n9511), .ZN(
        P1_U3217) );
  NOR2_X1 U10369 ( .A1(n9516), .A2(n5173), .ZN(n9517) );
  XNOR2_X1 U10370 ( .A(n9514), .B(n9517), .ZN(n9522) );
  AOI22_X1 U10371 ( .A1(n9810), .A2(n9566), .B1(P1_REG3_REG_21__SCAN_IN), .B2(
        P1_U3084), .ZN(n9519) );
  NAND2_X1 U10372 ( .A1(n9816), .A2(n9602), .ZN(n9518) );
  OAI211_X1 U10373 ( .C1(n9782), .C2(n9569), .A(n9519), .B(n9518), .ZN(n9520)
         );
  AOI21_X1 U10374 ( .B1(n9950), .B2(n9607), .A(n9520), .ZN(n9521) );
  OAI21_X1 U10375 ( .B1(n9522), .B2(n9609), .A(n9521), .ZN(P1_U3221) );
  XNOR2_X1 U10376 ( .A(n9524), .B(n9523), .ZN(n9525) );
  XNOR2_X1 U10377 ( .A(n9526), .B(n9525), .ZN(n9531) );
  AOI22_X1 U10378 ( .A1(n9601), .A2(n9755), .B1(P1_REG3_REG_25__SCAN_IN), .B2(
        P1_U3084), .ZN(n9528) );
  NAND2_X1 U10379 ( .A1(n9602), .A2(n9748), .ZN(n9527) );
  OAI211_X1 U10380 ( .C1(n9783), .C2(n9605), .A(n9528), .B(n9527), .ZN(n9529)
         );
  AOI21_X1 U10381 ( .B1(n9928), .B2(n9607), .A(n9529), .ZN(n9530) );
  OAI21_X1 U10382 ( .B1(n9531), .B2(n9609), .A(n9530), .ZN(P1_U3223) );
  INV_X1 U10383 ( .A(n9532), .ZN(n9980) );
  OAI21_X1 U10384 ( .B1(n9535), .B2(n9534), .A(n9533), .ZN(n9536) );
  NAND2_X1 U10385 ( .A1(n9536), .A2(n9590), .ZN(n9542) );
  AOI22_X1 U10386 ( .A1(n9601), .A2(n9616), .B1(P1_REG3_REG_16__SCAN_IN), .B2(
        P1_U3084), .ZN(n9537) );
  OAI21_X1 U10387 ( .B1(n9538), .B2(n9605), .A(n9537), .ZN(n9539) );
  AOI21_X1 U10388 ( .B1(n9540), .B2(n9602), .A(n9539), .ZN(n9541) );
  OAI211_X1 U10389 ( .C1(n9980), .C2(n9598), .A(n9542), .B(n9541), .ZN(
        P1_U3224) );
  XNOR2_X1 U10390 ( .A(n9545), .B(n9544), .ZN(n9546) );
  XNOR2_X1 U10391 ( .A(n9543), .B(n9546), .ZN(n9552) );
  AOI21_X1 U10392 ( .B1(n9566), .B2(n9617), .A(n9547), .ZN(n9549) );
  NAND2_X1 U10393 ( .A1(n9602), .A2(n9895), .ZN(n9548) );
  OAI211_X1 U10394 ( .C1(n9882), .C2(n9569), .A(n9549), .B(n9548), .ZN(n9550)
         );
  AOI21_X1 U10395 ( .B1(n9973), .B2(n9607), .A(n9550), .ZN(n9551) );
  OAI21_X1 U10396 ( .B1(n9552), .B2(n9609), .A(n9551), .ZN(P1_U3226) );
  OAI21_X1 U10397 ( .B1(n9555), .B2(n9554), .A(n9553), .ZN(n9556) );
  NAND2_X1 U10398 ( .A1(n9556), .A2(n9590), .ZN(n9560) );
  AOI22_X1 U10399 ( .A1(n9601), .A2(n9614), .B1(P1_REG3_REG_24__SCAN_IN), .B2(
        P1_U3084), .ZN(n9557) );
  OAI21_X1 U10400 ( .B1(n9766), .B2(n9605), .A(n9557), .ZN(n9558) );
  AOI21_X1 U10401 ( .B1(n9770), .B2(n9602), .A(n9558), .ZN(n9559) );
  OAI211_X1 U10402 ( .C1(n5182), .C2(n9598), .A(n9560), .B(n9559), .ZN(
        P1_U3227) );
  INV_X1 U10403 ( .A(n9561), .ZN(n9563) );
  NAND2_X1 U10404 ( .A1(n9563), .A2(n9562), .ZN(n9564) );
  XNOR2_X1 U10405 ( .A(n9565), .B(n9564), .ZN(n9572) );
  AOI22_X1 U10406 ( .A1(n9824), .A2(n9566), .B1(P1_REG3_REG_20__SCAN_IN), .B2(
        P1_U3084), .ZN(n9568) );
  NAND2_X1 U10407 ( .A1(n5485), .A2(n9602), .ZN(n9567) );
  OAI211_X1 U10408 ( .C1(n9581), .C2(n9569), .A(n9568), .B(n9567), .ZN(n9570)
         );
  AOI21_X1 U10409 ( .B1(n9954), .B2(n9607), .A(n9570), .ZN(n9571) );
  OAI21_X1 U10410 ( .B1(n9572), .B2(n9609), .A(n9571), .ZN(P1_U3231) );
  INV_X1 U10411 ( .A(n9944), .ZN(n9797) );
  INV_X1 U10412 ( .A(n9577), .ZN(n9573) );
  NOR2_X1 U10413 ( .A1(n9574), .A2(n9573), .ZN(n9579) );
  AOI21_X1 U10414 ( .B1(n9577), .B2(n9576), .A(n9575), .ZN(n9578) );
  OAI21_X1 U10415 ( .B1(n9579), .B2(n9578), .A(n9590), .ZN(n9584) );
  AOI22_X1 U10416 ( .A1(n9601), .A2(n9801), .B1(P1_REG3_REG_22__SCAN_IN), .B2(
        P1_U3084), .ZN(n9580) );
  OAI21_X1 U10417 ( .B1(n9581), .B2(n9605), .A(n9580), .ZN(n9582) );
  AOI21_X1 U10418 ( .B1(n9795), .B2(n9602), .A(n9582), .ZN(n9583) );
  OAI211_X1 U10419 ( .C1(n9797), .C2(n9598), .A(n9584), .B(n9583), .ZN(
        P1_U3233) );
  INV_X1 U10420 ( .A(n9873), .ZN(n9964) );
  INV_X1 U10421 ( .A(n9589), .ZN(n9586) );
  NOR2_X1 U10422 ( .A1(n9586), .A2(n9585), .ZN(n9592) );
  AOI21_X1 U10423 ( .B1(n9589), .B2(n9588), .A(n9587), .ZN(n9591) );
  OAI21_X1 U10424 ( .B1(n9592), .B2(n9591), .A(n9590), .ZN(n9597) );
  NOR2_X1 U10425 ( .A1(n9593), .A2(n9867), .ZN(n9595) );
  NAND2_X1 U10426 ( .A1(P1_U3084), .A2(P1_REG3_REG_18__SCAN_IN), .ZN(n9666) );
  OAI21_X1 U10427 ( .B1(n9605), .B2(n9860), .A(n9666), .ZN(n9594) );
  AOI211_X1 U10428 ( .C1(n9601), .C2(n9824), .A(n9595), .B(n9594), .ZN(n9596)
         );
  OAI211_X1 U10429 ( .C1(n9964), .C2(n9598), .A(n9597), .B(n9596), .ZN(
        P1_U3236) );
  XNOR2_X1 U10430 ( .A(n9599), .B(n9600), .ZN(n9610) );
  AOI22_X1 U10431 ( .A1(n9601), .A2(n9613), .B1(P1_REG3_REG_26__SCAN_IN), .B2(
        P1_U3084), .ZN(n9604) );
  NAND2_X1 U10432 ( .A1(n9602), .A2(n9734), .ZN(n9603) );
  OAI211_X1 U10433 ( .C1(n9768), .C2(n9605), .A(n9604), .B(n9603), .ZN(n9606)
         );
  AOI21_X1 U10434 ( .B1(n9923), .B2(n9607), .A(n9606), .ZN(n9608) );
  OAI21_X1 U10435 ( .B1(n9610), .B2(n9609), .A(n9608), .ZN(P1_U3238) );
  MUX2_X1 U10436 ( .A(P1_DATAO_REG_30__SCAN_IN), .B(n9611), .S(n9627), .Z(
        P1_U3585) );
  MUX2_X1 U10437 ( .A(P1_DATAO_REG_29__SCAN_IN), .B(n9612), .S(n9627), .Z(
        P1_U3584) );
  MUX2_X1 U10438 ( .A(P1_DATAO_REG_27__SCAN_IN), .B(n9613), .S(P1_U4006), .Z(
        P1_U3582) );
  MUX2_X1 U10439 ( .A(P1_DATAO_REG_26__SCAN_IN), .B(n9755), .S(P1_U4006), .Z(
        P1_U3581) );
  MUX2_X1 U10440 ( .A(P1_DATAO_REG_25__SCAN_IN), .B(n9614), .S(P1_U4006), .Z(
        P1_U3580) );
  MUX2_X1 U10441 ( .A(P1_DATAO_REG_24__SCAN_IN), .B(n9754), .S(P1_U4006), .Z(
        P1_U3579) );
  MUX2_X1 U10442 ( .A(P1_DATAO_REG_22__SCAN_IN), .B(n9811), .S(P1_U4006), .Z(
        P1_U3577) );
  MUX2_X1 U10443 ( .A(P1_DATAO_REG_21__SCAN_IN), .B(n9825), .S(P1_U4006), .Z(
        P1_U3576) );
  MUX2_X1 U10444 ( .A(P1_DATAO_REG_20__SCAN_IN), .B(n9810), .S(P1_U4006), .Z(
        P1_U3575) );
  MUX2_X1 U10445 ( .A(P1_DATAO_REG_19__SCAN_IN), .B(n9824), .S(P1_U4006), .Z(
        P1_U3574) );
  MUX2_X1 U10446 ( .A(P1_DATAO_REG_18__SCAN_IN), .B(n9615), .S(P1_U4006), .Z(
        P1_U3573) );
  MUX2_X1 U10447 ( .A(P1_DATAO_REG_17__SCAN_IN), .B(n9616), .S(P1_U4006), .Z(
        P1_U3572) );
  MUX2_X1 U10448 ( .A(P1_DATAO_REG_16__SCAN_IN), .B(n9617), .S(n9627), .Z(
        P1_U3571) );
  MUX2_X1 U10449 ( .A(P1_DATAO_REG_15__SCAN_IN), .B(n9618), .S(n9627), .Z(
        P1_U3570) );
  MUX2_X1 U10450 ( .A(P1_DATAO_REG_14__SCAN_IN), .B(n9619), .S(n9627), .Z(
        P1_U3569) );
  MUX2_X1 U10451 ( .A(P1_DATAO_REG_13__SCAN_IN), .B(n9620), .S(n9627), .Z(
        P1_U3568) );
  MUX2_X1 U10452 ( .A(P1_DATAO_REG_12__SCAN_IN), .B(n9621), .S(n9627), .Z(
        P1_U3567) );
  MUX2_X1 U10453 ( .A(P1_DATAO_REG_11__SCAN_IN), .B(n10624), .S(n9627), .Z(
        P1_U3566) );
  MUX2_X1 U10454 ( .A(P1_DATAO_REG_10__SCAN_IN), .B(n9622), .S(n9627), .Z(
        P1_U3565) );
  MUX2_X1 U10455 ( .A(P1_DATAO_REG_9__SCAN_IN), .B(n10621), .S(n9627), .Z(
        P1_U3564) );
  MUX2_X1 U10456 ( .A(P1_DATAO_REG_8__SCAN_IN), .B(n9623), .S(n9627), .Z(
        P1_U3563) );
  MUX2_X1 U10457 ( .A(P1_DATAO_REG_7__SCAN_IN), .B(n9624), .S(n9627), .Z(
        P1_U3562) );
  MUX2_X1 U10458 ( .A(P1_DATAO_REG_6__SCAN_IN), .B(n9625), .S(n9627), .Z(
        P1_U3561) );
  MUX2_X1 U10459 ( .A(P1_DATAO_REG_5__SCAN_IN), .B(n9626), .S(n9627), .Z(
        P1_U3560) );
  MUX2_X1 U10460 ( .A(P1_DATAO_REG_4__SCAN_IN), .B(n9628), .S(n9627), .Z(
        P1_U3559) );
  MUX2_X1 U10461 ( .A(P1_DATAO_REG_3__SCAN_IN), .B(n9629), .S(P1_U4006), .Z(
        P1_U3558) );
  MUX2_X1 U10462 ( .A(P1_DATAO_REG_2__SCAN_IN), .B(n9630), .S(P1_U4006), .Z(
        P1_U3557) );
  MUX2_X1 U10463 ( .A(P1_DATAO_REG_1__SCAN_IN), .B(n6896), .S(P1_U4006), .Z(
        P1_U3556) );
  MUX2_X1 U10464 ( .A(P1_DATAO_REG_0__SCAN_IN), .B(n9631), .S(P1_U4006), .Z(
        P1_U3555) );
  OAI21_X1 U10465 ( .B1(n9634), .B2(n9633), .A(n9632), .ZN(n9638) );
  INV_X1 U10466 ( .A(P1_ADDR_REG_4__SCAN_IN), .ZN(n9635) );
  NOR2_X1 U10467 ( .A1(n10391), .A2(n9635), .ZN(n9637) );
  AOI211_X1 U10468 ( .C1(n9638), .C2(n10398), .A(n9637), .B(n9636), .ZN(n9645)
         );
  OAI21_X1 U10469 ( .B1(n9641), .B2(n9640), .A(n9639), .ZN(n9642) );
  AOI22_X1 U10470 ( .A1(n9643), .A2(n9678), .B1(n10401), .B2(n9642), .ZN(n9644) );
  NAND3_X1 U10471 ( .A1(n9646), .A2(n9645), .A3(n9644), .ZN(P1_U3245) );
  AOI211_X1 U10472 ( .C1(n9649), .C2(n9648), .A(n9647), .B(n9673), .ZN(n9650)
         );
  INV_X1 U10473 ( .A(n9650), .ZN(n9661) );
  INV_X1 U10474 ( .A(P1_REG3_REG_16__SCAN_IN), .ZN(n9651) );
  NOR2_X1 U10475 ( .A1(P1_STATE_REG_SCAN_IN), .A2(n9651), .ZN(n9654) );
  INV_X1 U10476 ( .A(P1_ADDR_REG_16__SCAN_IN), .ZN(n9652) );
  NOR2_X1 U10477 ( .A1(n10391), .A2(n9652), .ZN(n9653) );
  AOI211_X1 U10478 ( .C1(n9678), .C2(n9655), .A(n9654), .B(n9653), .ZN(n9660)
         );
  OAI211_X1 U10479 ( .C1(n9658), .C2(n9657), .A(n10398), .B(n9656), .ZN(n9659)
         );
  NAND3_X1 U10480 ( .A1(n9661), .A2(n9660), .A3(n9659), .ZN(P1_U3257) );
  OAI21_X1 U10481 ( .B1(n9663), .B2(n9670), .A(n9662), .ZN(n9665) );
  INV_X1 U10482 ( .A(P1_REG1_REG_18__SCAN_IN), .ZN(n9971) );
  AOI22_X1 U10483 ( .A1(n9686), .A2(n9971), .B1(P1_REG1_REG_18__SCAN_IN), .B2(
        n9682), .ZN(n9664) );
  NOR2_X1 U10484 ( .A1(n9665), .A2(n9664), .ZN(n9681) );
  AOI21_X1 U10485 ( .B1(n9665), .B2(n9664), .A(n9681), .ZN(n9680) );
  INV_X1 U10486 ( .A(P1_ADDR_REG_18__SCAN_IN), .ZN(n9667) );
  OAI21_X1 U10487 ( .B1(n10391), .B2(n9667), .A(n9666), .ZN(n9677) );
  INV_X1 U10488 ( .A(P1_REG2_REG_18__SCAN_IN), .ZN(n9668) );
  MUX2_X1 U10489 ( .A(P1_REG2_REG_18__SCAN_IN), .B(n9668), .S(n9686), .Z(n9669) );
  INV_X1 U10490 ( .A(n9669), .ZN(n9675) );
  INV_X1 U10491 ( .A(n9670), .ZN(n9672) );
  NOR2_X1 U10492 ( .A1(n9674), .A2(n9675), .ZN(n9685) );
  AOI211_X1 U10493 ( .C1(n9675), .C2(n9674), .A(n9685), .B(n9673), .ZN(n9676)
         );
  AOI211_X1 U10494 ( .C1(n9678), .C2(n9686), .A(n9677), .B(n9676), .ZN(n9679)
         );
  OAI21_X1 U10495 ( .B1(n9680), .B2(n10380), .A(n9679), .ZN(P1_U3259) );
  AOI21_X1 U10496 ( .B1(n9971), .B2(n9682), .A(n9681), .ZN(n9684) );
  XNOR2_X1 U10497 ( .A(n6904), .B(P1_REG1_REG_19__SCAN_IN), .ZN(n9683) );
  XNOR2_X1 U10498 ( .A(n9684), .B(n9683), .ZN(n9693) );
  AOI21_X1 U10499 ( .B1(n9686), .B2(P1_REG2_REG_18__SCAN_IN), .A(n9685), .ZN(
        n9688) );
  MUX2_X1 U10500 ( .A(P1_REG2_REG_19__SCAN_IN), .B(n9840), .S(n9772), .Z(n9687) );
  OR2_X1 U10501 ( .A1(n10391), .A2(n5085), .ZN(n9689) );
  OAI211_X1 U10502 ( .C1(n10393), .C2(n6904), .A(n9690), .B(n9689), .ZN(n9691)
         );
  OAI21_X1 U10503 ( .B1(n9693), .B2(n10380), .A(n9692), .ZN(P1_U3260) );
  NAND2_X1 U10504 ( .A1(n9703), .A2(n9702), .ZN(n9701) );
  XNOR2_X1 U10505 ( .A(n9701), .B(n9906), .ZN(n9904) );
  NAND2_X1 U10506 ( .A1(n9904), .A2(n9902), .ZN(n9700) );
  NAND2_X1 U10507 ( .A1(n9694), .A2(n10640), .ZN(n9699) );
  NAND2_X1 U10508 ( .A1(n9696), .A2(n9695), .ZN(n9909) );
  INV_X1 U10509 ( .A(n9909), .ZN(n9697) );
  NAND2_X1 U10510 ( .A1(n9841), .A2(n9697), .ZN(n9704) );
  NAND2_X1 U10511 ( .A1(n9896), .A2(P1_REG2_REG_31__SCAN_IN), .ZN(n9698) );
  NAND4_X1 U10512 ( .A1(n9700), .A2(n9699), .A3(n9704), .A4(n9698), .ZN(
        P1_U3261) );
  OAI21_X1 U10513 ( .B1(n9703), .B2(n9702), .A(n9701), .ZN(n9910) );
  INV_X1 U10514 ( .A(P1_REG2_REG_30__SCAN_IN), .ZN(n9705) );
  OAI21_X1 U10515 ( .B1(n9841), .B2(n9705), .A(n9704), .ZN(n9706) );
  AOI21_X1 U10516 ( .B1(n9907), .B2(n10640), .A(n9706), .ZN(n9707) );
  OAI21_X1 U10517 ( .B1(n9910), .B2(n9870), .A(n9707), .ZN(P1_U3262) );
  XNOR2_X1 U10518 ( .A(n9709), .B(n9708), .ZN(n9922) );
  INV_X1 U10519 ( .A(n9733), .ZN(n9712) );
  INV_X1 U10520 ( .A(n9710), .ZN(n9711) );
  AOI211_X1 U10521 ( .C1(n9920), .C2(n9712), .A(n10597), .B(n9711), .ZN(n9919)
         );
  INV_X1 U10522 ( .A(n9919), .ZN(n9715) );
  INV_X1 U10523 ( .A(n9713), .ZN(n9714) );
  OAI22_X1 U10524 ( .A1(n9715), .A2(n9772), .B1(n9866), .B2(n9714), .ZN(n9722)
         );
  OAI211_X1 U10525 ( .C1(n9718), .C2(n9717), .A(n9716), .B(n9891), .ZN(n9720)
         );
  NAND2_X1 U10526 ( .A1(n9755), .A2(n10622), .ZN(n9719) );
  OAI211_X1 U10527 ( .C1(n9721), .C2(n9881), .A(n9720), .B(n9719), .ZN(n9918)
         );
  OAI21_X1 U10528 ( .B1(n9722), .B2(n9918), .A(n9841), .ZN(n9724) );
  AOI22_X1 U10529 ( .A1(n9920), .A2(n10640), .B1(P1_REG2_REG_27__SCAN_IN), 
        .B2(n9896), .ZN(n9723) );
  OAI211_X1 U10530 ( .C1(n9853), .C2(n9922), .A(n9724), .B(n9723), .ZN(
        P1_U3264) );
  XNOR2_X1 U10531 ( .A(n9725), .B(n9727), .ZN(n9732) );
  OAI22_X1 U10532 ( .A1(n9726), .A2(n9881), .B1(n9768), .B2(n9879), .ZN(n9731)
         );
  NAND2_X1 U10533 ( .A1(n9728), .A2(n9727), .ZN(n9729) );
  AOI21_X1 U10534 ( .B1(n9923), .B2(n9745), .A(n9733), .ZN(n9924) );
  AOI22_X1 U10535 ( .A1(n9896), .A2(P1_REG2_REG_26__SCAN_IN), .B1(n9734), .B2(
        n10638), .ZN(n9735) );
  OAI21_X1 U10536 ( .B1(n9736), .B2(n9898), .A(n9735), .ZN(n9738) );
  NOR2_X1 U10537 ( .A1(n9927), .A2(n9899), .ZN(n9737) );
  AOI211_X1 U10538 ( .C1(n9924), .C2(n9902), .A(n9738), .B(n9737), .ZN(n9739)
         );
  OAI21_X1 U10539 ( .B1(n9926), .B2(n9896), .A(n9739), .ZN(P1_U3265) );
  NAND2_X1 U10540 ( .A1(n9761), .A2(n9740), .ZN(n9742) );
  AND2_X1 U10541 ( .A1(n9742), .A2(n9741), .ZN(n9744) );
  XNOR2_X1 U10542 ( .A(n9744), .B(n9743), .ZN(n9932) );
  INV_X1 U10543 ( .A(n9769), .ZN(n9747) );
  INV_X1 U10544 ( .A(n9745), .ZN(n9746) );
  AOI21_X1 U10545 ( .B1(n9928), .B2(n9747), .A(n9746), .ZN(n9929) );
  AOI22_X1 U10546 ( .A1(n9896), .A2(P1_REG2_REG_25__SCAN_IN), .B1(n9748), .B2(
        n10638), .ZN(n9749) );
  OAI21_X1 U10547 ( .B1(n9750), .B2(n9898), .A(n9749), .ZN(n9758) );
  OAI21_X1 U10548 ( .B1(n9753), .B2(n9752), .A(n9751), .ZN(n9756) );
  AOI222_X1 U10549 ( .A1(n9891), .A2(n9756), .B1(n9755), .B2(n10623), .C1(
        n9754), .C2(n10622), .ZN(n9931) );
  NOR2_X1 U10550 ( .A1(n9931), .A2(n9896), .ZN(n9757) );
  AOI211_X1 U10551 ( .C1(n9929), .C2(n9902), .A(n9758), .B(n9757), .ZN(n9759)
         );
  OAI21_X1 U10552 ( .B1(n9853), .B2(n9932), .A(n9759), .ZN(P1_U3266) );
  NAND2_X1 U10553 ( .A1(n9761), .A2(n9760), .ZN(n9763) );
  XNOR2_X1 U10554 ( .A(n9763), .B(n9762), .ZN(n9937) );
  XNOR2_X1 U10555 ( .A(n9765), .B(n9764), .ZN(n9767) );
  OAI222_X1 U10556 ( .A1(n9881), .A2(n9768), .B1(n9767), .B2(n10626), .C1(
        n9879), .C2(n9766), .ZN(n9933) );
  AOI211_X1 U10557 ( .C1(n9935), .C2(n9784), .A(n10597), .B(n9769), .ZN(n9934)
         );
  INV_X1 U10558 ( .A(n9934), .ZN(n9773) );
  INV_X1 U10559 ( .A(n9770), .ZN(n9771) );
  OAI22_X1 U10560 ( .A1(n9773), .A2(n9772), .B1(n9866), .B2(n9771), .ZN(n9774)
         );
  OAI21_X1 U10561 ( .B1(n9933), .B2(n9774), .A(n9841), .ZN(n9776) );
  AOI22_X1 U10562 ( .A1(n9935), .A2(n10640), .B1(n9896), .B2(
        P1_REG2_REG_24__SCAN_IN), .ZN(n9775) );
  OAI211_X1 U10563 ( .C1(n9937), .C2(n9853), .A(n9776), .B(n9775), .ZN(
        P1_U3267) );
  XNOR2_X1 U10564 ( .A(n9777), .B(n9779), .ZN(n9943) );
  AOI21_X1 U10565 ( .B1(n9780), .B2(n9779), .A(n9778), .ZN(n9781) );
  OAI222_X1 U10566 ( .A1(n9881), .A2(n9783), .B1(n9879), .B2(n9782), .C1(
        n10626), .C2(n9781), .ZN(n9938) );
  INV_X1 U10567 ( .A(n9784), .ZN(n9785) );
  AOI21_X1 U10568 ( .B1(n9939), .B2(n5186), .A(n9785), .ZN(n9940) );
  NAND2_X1 U10569 ( .A1(n9940), .A2(n9902), .ZN(n9788) );
  AOI22_X1 U10570 ( .A1(n9896), .A2(P1_REG2_REG_23__SCAN_IN), .B1(n9786), .B2(
        n10638), .ZN(n9787) );
  OAI211_X1 U10571 ( .C1(n9789), .C2(n9898), .A(n9788), .B(n9787), .ZN(n9790)
         );
  AOI21_X1 U10572 ( .B1(n9938), .B2(n9841), .A(n9790), .ZN(n9791) );
  OAI21_X1 U10573 ( .B1(n9853), .B2(n9943), .A(n9791), .ZN(P1_U3268) );
  XNOR2_X1 U10574 ( .A(n9793), .B(n9792), .ZN(n9948) );
  AOI21_X1 U10575 ( .B1(n9944), .B2(n9813), .A(n9794), .ZN(n9945) );
  AOI22_X1 U10576 ( .A1(n9896), .A2(P1_REG2_REG_22__SCAN_IN), .B1(n9795), .B2(
        n10638), .ZN(n9796) );
  OAI21_X1 U10577 ( .B1(n9797), .B2(n9898), .A(n9796), .ZN(n9803) );
  XNOR2_X1 U10578 ( .A(n9799), .B(n9798), .ZN(n9800) );
  AOI222_X1 U10579 ( .A1(n9825), .A2(n10622), .B1(n9801), .B2(n10623), .C1(
        n9891), .C2(n9800), .ZN(n9947) );
  NOR2_X1 U10580 ( .A1(n9947), .A2(n9896), .ZN(n9802) );
  AOI211_X1 U10581 ( .C1(n9945), .C2(n9902), .A(n9803), .B(n9802), .ZN(n9804)
         );
  OAI21_X1 U10582 ( .B1(n9853), .B2(n9948), .A(n9804), .ZN(P1_U3269) );
  OAI21_X1 U10583 ( .B1(n9806), .B2(n8191), .A(n9805), .ZN(n9953) );
  AOI22_X1 U10584 ( .A1(n9950), .A2(n10640), .B1(P1_REG2_REG_21__SCAN_IN), 
        .B2(n9896), .ZN(n9820) );
  OAI21_X1 U10585 ( .B1(n9809), .B2(n9808), .A(n9807), .ZN(n9812) );
  AOI222_X1 U10586 ( .A1(n9891), .A2(n9812), .B1(n9811), .B2(n10623), .C1(
        n9810), .C2(n10622), .ZN(n9952) );
  INV_X1 U10587 ( .A(n9829), .ZN(n9815) );
  INV_X1 U10588 ( .A(n9813), .ZN(n9814) );
  AOI211_X1 U10589 ( .C1(n9950), .C2(n9815), .A(n10597), .B(n9814), .ZN(n9949)
         );
  AOI22_X1 U10590 ( .A1(n9949), .A2(n6904), .B1(n10638), .B2(n9816), .ZN(n9817) );
  AOI21_X1 U10591 ( .B1(n9952), .B2(n9817), .A(n9896), .ZN(n9818) );
  INV_X1 U10592 ( .A(n9818), .ZN(n9819) );
  OAI211_X1 U10593 ( .C1(n9953), .C2(n9853), .A(n9820), .B(n9819), .ZN(
        P1_U3270) );
  XNOR2_X1 U10594 ( .A(n9821), .B(n9822), .ZN(n9832) );
  XNOR2_X1 U10595 ( .A(n9823), .B(n9822), .ZN(n9827) );
  AOI22_X1 U10596 ( .A1(n9825), .A2(n10623), .B1(n10622), .B2(n9824), .ZN(
        n9826) );
  OAI21_X1 U10597 ( .B1(n9827), .B2(n10626), .A(n9826), .ZN(n9828) );
  AOI21_X1 U10598 ( .B1(n9832), .B2(n10629), .A(n9828), .ZN(n9957) );
  AOI21_X1 U10599 ( .B1(n9954), .B2(n9842), .A(n9829), .ZN(n9955) );
  INV_X1 U10600 ( .A(n9954), .ZN(n9831) );
  AOI22_X1 U10601 ( .A1(n5485), .A2(n10638), .B1(n9896), .B2(
        P1_REG2_REG_20__SCAN_IN), .ZN(n9830) );
  OAI21_X1 U10602 ( .B1(n9831), .B2(n9898), .A(n9830), .ZN(n9834) );
  INV_X1 U10603 ( .A(n9832), .ZN(n9958) );
  NOR2_X1 U10604 ( .A1(n9958), .A2(n9899), .ZN(n9833) );
  AOI211_X1 U10605 ( .C1(n9955), .C2(n9902), .A(n9834), .B(n9833), .ZN(n9835)
         );
  OAI21_X1 U10606 ( .B1(n9896), .B2(n9957), .A(n9835), .ZN(P1_U3271) );
  NAND2_X1 U10607 ( .A1(n9836), .A2(n9837), .ZN(n9838) );
  XOR2_X1 U10608 ( .A(n9838), .B(n9846), .Z(n9963) );
  OAI22_X1 U10609 ( .A1(n9841), .A2(n9840), .B1(n9839), .B2(n9866), .ZN(n9851)
         );
  INV_X1 U10610 ( .A(n9868), .ZN(n9844) );
  INV_X1 U10611 ( .A(n9842), .ZN(n9843) );
  AOI211_X1 U10612 ( .C1(n9961), .C2(n9844), .A(n10597), .B(n9843), .ZN(n9960)
         );
  XOR2_X1 U10613 ( .A(n9845), .B(n9846), .Z(n9847) );
  OAI222_X1 U10614 ( .A1(n9881), .A2(n9848), .B1(n9847), .B2(n10626), .C1(
        n9879), .C2(n9882), .ZN(n9959) );
  AOI21_X1 U10615 ( .B1(n9960), .B2(n6904), .A(n9959), .ZN(n9849) );
  NOR2_X1 U10616 ( .A1(n9849), .A2(n9896), .ZN(n9850) );
  AOI211_X1 U10617 ( .C1(n10640), .C2(n9961), .A(n9851), .B(n9850), .ZN(n9852)
         );
  OAI21_X1 U10618 ( .B1(n9853), .B2(n9963), .A(n9852), .ZN(P1_U3272) );
  NAND2_X1 U10619 ( .A1(n9854), .A2(n9859), .ZN(n9855) );
  INV_X1 U10620 ( .A(n9856), .ZN(n9968) );
  NAND2_X1 U10621 ( .A1(n9856), .A2(n10629), .ZN(n9865) );
  OAI21_X1 U10622 ( .B1(n9859), .B2(n9858), .A(n9857), .ZN(n9863) );
  OAI22_X1 U10623 ( .A1(n9861), .A2(n9881), .B1(n9860), .B2(n9879), .ZN(n9862)
         );
  AOI21_X1 U10624 ( .B1(n9863), .B2(n9891), .A(n9862), .ZN(n9864) );
  NAND2_X1 U10625 ( .A1(n9865), .A2(n9864), .ZN(n9970) );
  NAND2_X1 U10626 ( .A1(n9970), .A2(n9841), .ZN(n9875) );
  OAI22_X1 U10627 ( .A1(n9841), .A2(n9668), .B1(n9867), .B2(n9866), .ZN(n9872)
         );
  AND2_X1 U10628 ( .A1(n9873), .A2(n9892), .ZN(n9869) );
  OR2_X1 U10629 ( .A1(n9869), .A2(n9868), .ZN(n9965) );
  NOR2_X1 U10630 ( .A1(n9965), .A2(n9870), .ZN(n9871) );
  AOI211_X1 U10631 ( .C1(n10640), .C2(n9873), .A(n9872), .B(n9871), .ZN(n9874)
         );
  OAI211_X1 U10632 ( .C1(n9968), .C2(n9899), .A(n9875), .B(n9874), .ZN(
        P1_U3273) );
  OAI21_X1 U10633 ( .B1(n9878), .B2(n9877), .A(n9876), .ZN(n9890) );
  OAI22_X1 U10634 ( .A1(n9882), .A2(n9881), .B1(n9880), .B2(n9879), .ZN(n9889)
         );
  OAI21_X1 U10635 ( .B1(n9885), .B2(n9884), .A(n9883), .ZN(n9886) );
  INV_X1 U10636 ( .A(n9886), .ZN(n9977) );
  NOR2_X1 U10637 ( .A1(n9977), .A2(n9887), .ZN(n9888) );
  AOI211_X1 U10638 ( .C1(n9891), .C2(n9890), .A(n9889), .B(n9888), .ZN(n9976)
         );
  INV_X1 U10639 ( .A(n9892), .ZN(n9893) );
  AOI21_X1 U10640 ( .B1(n9973), .B2(n9894), .A(n9893), .ZN(n9974) );
  AOI22_X1 U10641 ( .A1(n9896), .A2(P1_REG2_REG_17__SCAN_IN), .B1(n9895), .B2(
        n10638), .ZN(n9897) );
  OAI21_X1 U10642 ( .B1(n5193), .B2(n9898), .A(n9897), .ZN(n9901) );
  NOR2_X1 U10643 ( .A1(n9977), .A2(n9899), .ZN(n9900) );
  AOI211_X1 U10644 ( .C1(n9974), .C2(n9902), .A(n9901), .B(n9900), .ZN(n9903)
         );
  OAI21_X1 U10645 ( .B1(n9976), .B2(n9896), .A(n9903), .ZN(P1_U3274) );
  NAND2_X1 U10646 ( .A1(n9904), .A2(n10617), .ZN(n9905) );
  OAI211_X1 U10647 ( .C1(n9906), .C2(n10618), .A(n9905), .B(n9909), .ZN(n10008) );
  MUX2_X1 U10648 ( .A(P1_REG1_REG_31__SCAN_IN), .B(n10008), .S(n10634), .Z(
        P1_U3554) );
  NAND2_X1 U10649 ( .A1(n9907), .A2(n10578), .ZN(n9908) );
  OAI211_X1 U10650 ( .C1(n9910), .C2(n10597), .A(n9909), .B(n9908), .ZN(n10009) );
  MUX2_X1 U10651 ( .A(P1_REG1_REG_30__SCAN_IN), .B(n10009), .S(n10634), .Z(
        P1_U3553) );
  AOI22_X1 U10652 ( .A1(n9911), .A2(n10617), .B1(n10578), .B2(n8327), .ZN(
        n9912) );
  AOI22_X1 U10653 ( .A1(n9915), .A2(n10617), .B1(n10578), .B2(n8291), .ZN(
        n9916) );
  MUX2_X1 U10654 ( .A(P1_REG1_REG_28__SCAN_IN), .B(n10010), .S(n10634), .Z(
        P1_U3551) );
  OAI21_X1 U10655 ( .B1(n10001), .B2(n9922), .A(n9921), .ZN(n10011) );
  MUX2_X1 U10656 ( .A(P1_REG1_REG_27__SCAN_IN), .B(n10011), .S(n10634), .Z(
        P1_U3550) );
  AOI22_X1 U10657 ( .A1(n9924), .A2(n10617), .B1(n10578), .B2(n9923), .ZN(
        n9925) );
  MUX2_X1 U10658 ( .A(P1_REG1_REG_26__SCAN_IN), .B(n10012), .S(n10634), .Z(
        P1_U3549) );
  AOI22_X1 U10659 ( .A1(n9929), .A2(n10617), .B1(n10578), .B2(n9928), .ZN(
        n9930) );
  OAI211_X1 U10660 ( .C1(n10001), .C2(n9932), .A(n9931), .B(n9930), .ZN(n10013) );
  MUX2_X1 U10661 ( .A(P1_REG1_REG_25__SCAN_IN), .B(n10013), .S(n10634), .Z(
        P1_U3548) );
  AOI211_X1 U10662 ( .C1(n10578), .C2(n9935), .A(n9934), .B(n9933), .ZN(n9936)
         );
  OAI21_X1 U10663 ( .B1(n10001), .B2(n9937), .A(n9936), .ZN(n10014) );
  MUX2_X1 U10664 ( .A(P1_REG1_REG_24__SCAN_IN), .B(n10014), .S(n10634), .Z(
        P1_U3547) );
  INV_X1 U10665 ( .A(n9938), .ZN(n9942) );
  AOI22_X1 U10666 ( .A1(n9940), .A2(n10617), .B1(n10578), .B2(n9939), .ZN(
        n9941) );
  OAI211_X1 U10667 ( .C1(n10001), .C2(n9943), .A(n9942), .B(n9941), .ZN(n10015) );
  MUX2_X1 U10668 ( .A(P1_REG1_REG_23__SCAN_IN), .B(n10015), .S(n10634), .Z(
        P1_U3546) );
  AOI22_X1 U10669 ( .A1(n9945), .A2(n10617), .B1(n10578), .B2(n9944), .ZN(
        n9946) );
  OAI211_X1 U10670 ( .C1(n9948), .C2(n10001), .A(n9947), .B(n9946), .ZN(n10016) );
  MUX2_X1 U10671 ( .A(P1_REG1_REG_22__SCAN_IN), .B(n10016), .S(n10634), .Z(
        P1_U3545) );
  AOI21_X1 U10672 ( .B1(n10578), .B2(n9950), .A(n9949), .ZN(n9951) );
  OAI211_X1 U10673 ( .C1(n9953), .C2(n10001), .A(n9952), .B(n9951), .ZN(n10017) );
  MUX2_X1 U10674 ( .A(P1_REG1_REG_21__SCAN_IN), .B(n10017), .S(n10634), .Z(
        P1_U3544) );
  AOI22_X1 U10675 ( .A1(n9955), .A2(n10617), .B1(n10578), .B2(n9954), .ZN(
        n9956) );
  OAI211_X1 U10676 ( .C1(n9958), .C2(n10582), .A(n9957), .B(n9956), .ZN(n10018) );
  MUX2_X1 U10677 ( .A(P1_REG1_REG_20__SCAN_IN), .B(n10018), .S(n10634), .Z(
        P1_U3543) );
  AOI211_X1 U10678 ( .C1(n10578), .C2(n9961), .A(n9960), .B(n9959), .ZN(n9962)
         );
  OAI21_X1 U10679 ( .B1(n9963), .B2(n10001), .A(n9962), .ZN(n10019) );
  MUX2_X1 U10680 ( .A(P1_REG1_REG_19__SCAN_IN), .B(n10019), .S(n10634), .Z(
        P1_U3542) );
  OAI22_X1 U10681 ( .A1(n9965), .A2(n10597), .B1(n9964), .B2(n10618), .ZN(
        n9966) );
  INV_X1 U10682 ( .A(n9966), .ZN(n9967) );
  OAI21_X1 U10683 ( .B1(n9968), .B2(n10582), .A(n9967), .ZN(n9969) );
  NOR2_X1 U10684 ( .A1(n9970), .A2(n9969), .ZN(n10020) );
  MUX2_X1 U10685 ( .A(n9971), .B(n10020), .S(n10634), .Z(n9972) );
  INV_X1 U10686 ( .A(n9972), .ZN(P1_U3541) );
  AOI22_X1 U10687 ( .A1(n9974), .A2(n10617), .B1(n10578), .B2(n9973), .ZN(
        n9975) );
  OAI211_X1 U10688 ( .C1(n9977), .C2(n10582), .A(n9976), .B(n9975), .ZN(n10023) );
  MUX2_X1 U10689 ( .A(P1_REG1_REG_17__SCAN_IN), .B(n10023), .S(n10634), .Z(
        P1_U3540) );
  OR2_X1 U10690 ( .A1(n9978), .A2(n10001), .ZN(n9984) );
  OAI21_X1 U10691 ( .B1(n9980), .B2(n10618), .A(n9979), .ZN(n9981) );
  NOR2_X1 U10692 ( .A1(n9982), .A2(n9981), .ZN(n9983) );
  NAND2_X1 U10693 ( .A1(n9984), .A2(n9983), .ZN(n10024) );
  MUX2_X1 U10694 ( .A(P1_REG1_REG_16__SCAN_IN), .B(n10024), .S(n10634), .Z(
        P1_U3539) );
  INV_X1 U10695 ( .A(n9985), .ZN(n9990) );
  AOI22_X1 U10696 ( .A1(n9987), .A2(n10617), .B1(n10578), .B2(n9986), .ZN(
        n9988) );
  OAI211_X1 U10697 ( .C1(n10582), .C2(n9990), .A(n9989), .B(n9988), .ZN(n10025) );
  MUX2_X1 U10698 ( .A(n10025), .B(P1_REG1_REG_15__SCAN_IN), .S(n10633), .Z(
        P1_U3538) );
  AOI211_X1 U10699 ( .C1(n10578), .C2(n9993), .A(n9992), .B(n9991), .ZN(n9994)
         );
  OAI21_X1 U10700 ( .B1(n9995), .B2(n10001), .A(n9994), .ZN(n10026) );
  MUX2_X1 U10701 ( .A(n10026), .B(P1_REG1_REG_14__SCAN_IN), .S(n10633), .Z(
        P1_U3537) );
  AOI211_X1 U10702 ( .C1(n10578), .C2(n9998), .A(n9997), .B(n9996), .ZN(n9999)
         );
  OAI21_X1 U10703 ( .B1(n10001), .B2(n10000), .A(n9999), .ZN(n10027) );
  MUX2_X1 U10704 ( .A(P1_REG1_REG_12__SCAN_IN), .B(n10027), .S(n10634), .Z(
        P1_U3535) );
  INV_X1 U10705 ( .A(n10002), .ZN(n10007) );
  AOI22_X1 U10706 ( .A1(n10004), .A2(n10617), .B1(n10578), .B2(n10003), .ZN(
        n10005) );
  OAI211_X1 U10707 ( .C1(n10007), .C2(n10582), .A(n10006), .B(n10005), .ZN(
        n10028) );
  MUX2_X1 U10708 ( .A(P1_REG1_REG_11__SCAN_IN), .B(n10028), .S(n10634), .Z(
        P1_U3534) );
  MUX2_X1 U10709 ( .A(P1_REG0_REG_31__SCAN_IN), .B(n10008), .S(n10637), .Z(
        P1_U3522) );
  MUX2_X1 U10710 ( .A(P1_REG0_REG_30__SCAN_IN), .B(n10009), .S(n10637), .Z(
        P1_U3521) );
  MUX2_X1 U10711 ( .A(P1_REG0_REG_27__SCAN_IN), .B(n10011), .S(n10637), .Z(
        P1_U3518) );
  MUX2_X1 U10712 ( .A(P1_REG0_REG_26__SCAN_IN), .B(n10012), .S(n10637), .Z(
        P1_U3517) );
  MUX2_X1 U10713 ( .A(P1_REG0_REG_25__SCAN_IN), .B(n10013), .S(n10637), .Z(
        P1_U3516) );
  MUX2_X1 U10714 ( .A(P1_REG0_REG_24__SCAN_IN), .B(n10014), .S(n10637), .Z(
        P1_U3515) );
  MUX2_X1 U10715 ( .A(P1_REG0_REG_23__SCAN_IN), .B(n10015), .S(n10637), .Z(
        P1_U3514) );
  MUX2_X1 U10716 ( .A(P1_REG0_REG_22__SCAN_IN), .B(n10016), .S(n10637), .Z(
        P1_U3513) );
  MUX2_X1 U10717 ( .A(P1_REG0_REG_21__SCAN_IN), .B(n10017), .S(n10637), .Z(
        P1_U3512) );
  MUX2_X1 U10718 ( .A(P1_REG0_REG_20__SCAN_IN), .B(n10018), .S(n10637), .Z(
        P1_U3511) );
  MUX2_X1 U10719 ( .A(P1_REG0_REG_19__SCAN_IN), .B(n10019), .S(n10637), .Z(
        P1_U3510) );
  INV_X1 U10720 ( .A(P1_REG0_REG_18__SCAN_IN), .ZN(n10021) );
  MUX2_X1 U10721 ( .A(n10021), .B(n10020), .S(n10637), .Z(n10022) );
  INV_X1 U10722 ( .A(n10022), .ZN(P1_U3508) );
  MUX2_X1 U10723 ( .A(P1_REG0_REG_17__SCAN_IN), .B(n10023), .S(n10637), .Z(
        P1_U3505) );
  MUX2_X1 U10724 ( .A(P1_REG0_REG_16__SCAN_IN), .B(n10024), .S(n10637), .Z(
        P1_U3502) );
  MUX2_X1 U10725 ( .A(n10025), .B(P1_REG0_REG_15__SCAN_IN), .S(n10635), .Z(
        P1_U3499) );
  MUX2_X1 U10726 ( .A(P1_REG0_REG_14__SCAN_IN), .B(n10026), .S(n10637), .Z(
        P1_U3496) );
  MUX2_X1 U10727 ( .A(P1_REG0_REG_12__SCAN_IN), .B(n10027), .S(n10637), .Z(
        P1_U3490) );
  MUX2_X1 U10728 ( .A(P1_REG0_REG_11__SCAN_IN), .B(n10028), .S(n10637), .Z(
        P1_U3487) );
  NAND3_X1 U10729 ( .A1(n6443), .A2(P1_STATE_REG_SCAN_IN), .A3(
        P1_IR_REG_31__SCAN_IN), .ZN(n10030) );
  OAI22_X1 U10730 ( .A1(n10029), .A2(n10030), .B1(n6424), .B2(n10039), .ZN(
        n10031) );
  INV_X1 U10731 ( .A(n10031), .ZN(n10032) );
  OAI21_X1 U10732 ( .B1(n10034), .B2(n10033), .A(n10032), .ZN(P1_U3322) );
  OAI222_X1 U10733 ( .A1(n10043), .A2(n10038), .B1(n10037), .B2(P1_U3084), 
        .C1(n10035), .C2(n10039), .ZN(P1_U3323) );
  OAI222_X1 U10734 ( .A1(n10043), .A2(n10042), .B1(P1_U3084), .B2(n10041), 
        .C1(n10040), .C2(n10039), .ZN(P1_U3324) );
  INV_X1 U10735 ( .A(n10044), .ZN(n10045) );
  MUX2_X1 U10736 ( .A(n10045), .B(P1_IR_REG_0__SCAN_IN), .S(
        P1_STATE_REG_SCAN_IN), .Z(P1_U3353) );
  NAND2_X1 U10737 ( .A1(n10047), .A2(n10046), .ZN(n10048) );
  AND2_X1 U10738 ( .A1(P1_D_REG_2__SCAN_IN), .A2(n10048), .ZN(P1_U3321) );
  AND2_X1 U10739 ( .A1(P1_D_REG_3__SCAN_IN), .A2(n10048), .ZN(P1_U3320) );
  AND2_X1 U10740 ( .A1(P1_D_REG_4__SCAN_IN), .A2(n10048), .ZN(P1_U3319) );
  AND2_X1 U10741 ( .A1(P1_D_REG_5__SCAN_IN), .A2(n10048), .ZN(P1_U3318) );
  AND2_X1 U10742 ( .A1(P1_D_REG_6__SCAN_IN), .A2(n10048), .ZN(P1_U3317) );
  AND2_X1 U10743 ( .A1(P1_D_REG_7__SCAN_IN), .A2(n10048), .ZN(P1_U3316) );
  AND2_X1 U10744 ( .A1(P1_D_REG_8__SCAN_IN), .A2(n10048), .ZN(P1_U3315) );
  AND2_X1 U10745 ( .A1(P1_D_REG_9__SCAN_IN), .A2(n10048), .ZN(P1_U3314) );
  AND2_X1 U10746 ( .A1(P1_D_REG_10__SCAN_IN), .A2(n10048), .ZN(P1_U3313) );
  AND2_X1 U10747 ( .A1(P1_D_REG_11__SCAN_IN), .A2(n10048), .ZN(P1_U3312) );
  AND2_X1 U10748 ( .A1(P1_D_REG_12__SCAN_IN), .A2(n10048), .ZN(P1_U3311) );
  AND2_X1 U10749 ( .A1(P1_D_REG_13__SCAN_IN), .A2(n10048), .ZN(P1_U3310) );
  AND2_X1 U10750 ( .A1(P1_D_REG_14__SCAN_IN), .A2(n10048), .ZN(P1_U3309) );
  AND2_X1 U10751 ( .A1(P1_D_REG_15__SCAN_IN), .A2(n10048), .ZN(P1_U3308) );
  AND2_X1 U10752 ( .A1(P1_D_REG_16__SCAN_IN), .A2(n10048), .ZN(P1_U3307) );
  AND2_X1 U10753 ( .A1(P1_D_REG_17__SCAN_IN), .A2(n10048), .ZN(P1_U3306) );
  AND2_X1 U10754 ( .A1(P1_D_REG_18__SCAN_IN), .A2(n10048), .ZN(P1_U3305) );
  AND2_X1 U10755 ( .A1(P1_D_REG_19__SCAN_IN), .A2(n10048), .ZN(P1_U3304) );
  AND2_X1 U10756 ( .A1(P1_D_REG_20__SCAN_IN), .A2(n10048), .ZN(P1_U3303) );
  AND2_X1 U10757 ( .A1(P1_D_REG_21__SCAN_IN), .A2(n10048), .ZN(P1_U3302) );
  AND2_X1 U10758 ( .A1(P1_D_REG_22__SCAN_IN), .A2(n10048), .ZN(P1_U3301) );
  AND2_X1 U10759 ( .A1(P1_D_REG_23__SCAN_IN), .A2(n10048), .ZN(P1_U3300) );
  AND2_X1 U10760 ( .A1(P1_D_REG_24__SCAN_IN), .A2(n10048), .ZN(P1_U3299) );
  AND2_X1 U10761 ( .A1(P1_D_REG_25__SCAN_IN), .A2(n10048), .ZN(P1_U3298) );
  AND2_X1 U10762 ( .A1(P1_D_REG_26__SCAN_IN), .A2(n10048), .ZN(P1_U3297) );
  AND2_X1 U10763 ( .A1(P1_D_REG_27__SCAN_IN), .A2(n10048), .ZN(P1_U3296) );
  AND2_X1 U10764 ( .A1(P1_D_REG_28__SCAN_IN), .A2(n10048), .ZN(P1_U3295) );
  AND2_X1 U10765 ( .A1(P1_D_REG_29__SCAN_IN), .A2(n10048), .ZN(P1_U3294) );
  AND2_X1 U10766 ( .A1(P1_D_REG_30__SCAN_IN), .A2(n10048), .ZN(P1_U3293) );
  AND2_X1 U10767 ( .A1(P1_D_REG_31__SCAN_IN), .A2(n10048), .ZN(P1_U3292) );
  NOR2_X1 U10768 ( .A1(n10049), .A2(n10408), .ZN(n10054) );
  INV_X1 U10769 ( .A(P2_D_REG_1__SCAN_IN), .ZN(n10053) );
  INV_X1 U10770 ( .A(n10050), .ZN(n10052) );
  AOI22_X1 U10771 ( .A1(n10413), .A2(n10054), .B1(n10053), .B2(n10410), .ZN(
        P2_U3438) );
  AND2_X1 U10772 ( .A1(P2_D_REG_2__SCAN_IN), .A2(n10410), .ZN(P2_U3326) );
  AND2_X1 U10773 ( .A1(P2_D_REG_3__SCAN_IN), .A2(n10410), .ZN(P2_U3325) );
  AND2_X1 U10774 ( .A1(P2_D_REG_4__SCAN_IN), .A2(n10410), .ZN(P2_U3324) );
  AND2_X1 U10775 ( .A1(P2_D_REG_5__SCAN_IN), .A2(n10410), .ZN(P2_U3323) );
  AND2_X1 U10776 ( .A1(P2_D_REG_6__SCAN_IN), .A2(n10410), .ZN(P2_U3322) );
  AND2_X1 U10777 ( .A1(P2_D_REG_7__SCAN_IN), .A2(n10410), .ZN(P2_U3321) );
  AND2_X1 U10778 ( .A1(P2_D_REG_8__SCAN_IN), .A2(n10410), .ZN(P2_U3320) );
  AND2_X1 U10779 ( .A1(P2_D_REG_9__SCAN_IN), .A2(n10410), .ZN(P2_U3319) );
  AND2_X1 U10780 ( .A1(P2_D_REG_10__SCAN_IN), .A2(n10410), .ZN(P2_U3318) );
  AND2_X1 U10781 ( .A1(P2_D_REG_11__SCAN_IN), .A2(n10410), .ZN(P2_U3317) );
  AND2_X1 U10782 ( .A1(P2_D_REG_12__SCAN_IN), .A2(n10410), .ZN(P2_U3316) );
  AND2_X1 U10783 ( .A1(P2_D_REG_13__SCAN_IN), .A2(n10410), .ZN(P2_U3315) );
  AND2_X1 U10784 ( .A1(P2_D_REG_14__SCAN_IN), .A2(n10410), .ZN(P2_U3314) );
  AND2_X1 U10785 ( .A1(P2_D_REG_15__SCAN_IN), .A2(n10410), .ZN(P2_U3313) );
  AND2_X1 U10786 ( .A1(P2_D_REG_16__SCAN_IN), .A2(n10410), .ZN(P2_U3312) );
  AND2_X1 U10787 ( .A1(P2_D_REG_17__SCAN_IN), .A2(n10410), .ZN(P2_U3311) );
  AND2_X1 U10788 ( .A1(P2_D_REG_18__SCAN_IN), .A2(n10410), .ZN(P2_U3310) );
  AND2_X1 U10789 ( .A1(P2_D_REG_19__SCAN_IN), .A2(n10410), .ZN(P2_U3309) );
  AND2_X1 U10790 ( .A1(P2_D_REG_20__SCAN_IN), .A2(n10410), .ZN(P2_U3308) );
  AND2_X1 U10791 ( .A1(P2_D_REG_21__SCAN_IN), .A2(n10410), .ZN(P2_U3307) );
  AND2_X1 U10792 ( .A1(P2_D_REG_22__SCAN_IN), .A2(n10410), .ZN(P2_U3306) );
  AND2_X1 U10793 ( .A1(P2_D_REG_23__SCAN_IN), .A2(n10410), .ZN(P2_U3305) );
  AND2_X1 U10794 ( .A1(P2_D_REG_24__SCAN_IN), .A2(n10410), .ZN(P2_U3304) );
  AND2_X1 U10795 ( .A1(P2_D_REG_25__SCAN_IN), .A2(n10410), .ZN(P2_U3303) );
  AND2_X1 U10796 ( .A1(P2_D_REG_26__SCAN_IN), .A2(n10410), .ZN(P2_U3302) );
  AND2_X1 U10797 ( .A1(P2_D_REG_27__SCAN_IN), .A2(n10410), .ZN(P2_U3301) );
  AND2_X1 U10798 ( .A1(P2_D_REG_28__SCAN_IN), .A2(n10410), .ZN(P2_U3300) );
  AND2_X1 U10799 ( .A1(P2_D_REG_29__SCAN_IN), .A2(n10410), .ZN(P2_U3299) );
  AND2_X1 U10800 ( .A1(P2_D_REG_30__SCAN_IN), .A2(n10410), .ZN(P2_U3298) );
  AND2_X1 U10801 ( .A1(P2_D_REG_31__SCAN_IN), .A2(n10410), .ZN(P2_U3297) );
  OAI22_X1 U10802 ( .A1(n5684), .A2(keyinput_125), .B1(n10267), .B2(
        keyinput_124), .ZN(n10055) );
  AOI221_X1 U10803 ( .B1(n5684), .B2(keyinput_125), .C1(keyinput_124), .C2(
        n10267), .A(n10055), .ZN(n10153) );
  XOR2_X1 U10804 ( .A(n10264), .B(keyinput_121), .Z(n10151) );
  INV_X1 U10805 ( .A(keyinput_120), .ZN(n10146) );
  INV_X1 U10806 ( .A(P2_REG3_REG_0__SCAN_IN), .ZN(n10259) );
  OAI22_X1 U10807 ( .A1(n5719), .A2(keyinput_117), .B1(n10057), .B2(
        keyinput_119), .ZN(n10056) );
  AOI221_X1 U10808 ( .B1(n5719), .B2(keyinput_117), .C1(keyinput_119), .C2(
        n10057), .A(n10056), .ZN(n10143) );
  AOI22_X1 U10809 ( .A1(n10059), .A2(keyinput_115), .B1(n5911), .B2(
        keyinput_114), .ZN(n10058) );
  OAI221_X1 U10810 ( .B1(n10059), .B2(keyinput_115), .C1(n5911), .C2(
        keyinput_114), .A(n10058), .ZN(n10141) );
  INV_X1 U10811 ( .A(keyinput_113), .ZN(n10138) );
  INV_X1 U10812 ( .A(keyinput_112), .ZN(n10136) );
  INV_X1 U10813 ( .A(keyinput_111), .ZN(n10134) );
  XOR2_X1 U10814 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_106), .Z(n10132)
         );
  INV_X1 U10815 ( .A(keyinput_105), .ZN(n10125) );
  XOR2_X1 U10816 ( .A(P2_RD_REG_SCAN_IN), .B(keyinput_97), .Z(n10123) );
  INV_X1 U10817 ( .A(keyinput_90), .ZN(n10101) );
  INV_X1 U10818 ( .A(keyinput_89), .ZN(n10099) );
  INV_X1 U10819 ( .A(SI_8_), .ZN(n10206) );
  INV_X1 U10820 ( .A(keyinput_88), .ZN(n10097) );
  INV_X1 U10821 ( .A(keyinput_87), .ZN(n10095) );
  OAI22_X1 U10822 ( .A1(n10062), .A2(keyinput_76), .B1(n10061), .B2(
        keyinput_77), .ZN(n10060) );
  AOI221_X1 U10823 ( .B1(n10062), .B2(keyinput_76), .C1(keyinput_77), .C2(
        n10061), .A(n10060), .ZN(n10081) );
  INV_X1 U10824 ( .A(keyinput_75), .ZN(n10079) );
  INV_X1 U10825 ( .A(keyinput_71), .ZN(n10073) );
  INV_X1 U10826 ( .A(keyinput_70), .ZN(n10071) );
  OAI22_X1 U10827 ( .A1(n10165), .A2(keyinput_68), .B1(SI_29_), .B2(
        keyinput_67), .ZN(n10063) );
  AOI221_X1 U10828 ( .B1(n10165), .B2(keyinput_68), .C1(keyinput_67), .C2(
        SI_29_), .A(n10063), .ZN(n10068) );
  INV_X1 U10829 ( .A(keyinput_66), .ZN(n10066) );
  OAI22_X1 U10830 ( .A1(SI_31_), .A2(keyinput_65), .B1(keyinput_64), .B2(
        P2_WR_REG_SCAN_IN), .ZN(n10064) );
  AOI221_X1 U10831 ( .B1(SI_31_), .B2(keyinput_65), .C1(P2_WR_REG_SCAN_IN), 
        .C2(keyinput_64), .A(n10064), .ZN(n10065) );
  OAI221_X1 U10832 ( .B1(SI_30_), .B2(n10066), .C1(n10161), .C2(keyinput_66), 
        .A(n10065), .ZN(n10067) );
  OAI211_X1 U10833 ( .C1(n10169), .C2(keyinput_69), .A(n10068), .B(n10067), 
        .ZN(n10069) );
  AOI21_X1 U10834 ( .B1(n10169), .B2(keyinput_69), .A(n10069), .ZN(n10070) );
  AOI221_X1 U10835 ( .B1(SI_26_), .B2(n10071), .C1(n10171), .C2(keyinput_70), 
        .A(n10070), .ZN(n10072) );
  AOI221_X1 U10836 ( .B1(SI_25_), .B2(keyinput_71), .C1(n10174), .C2(n10073), 
        .A(n10072), .ZN(n10076) );
  AOI22_X1 U10837 ( .A1(SI_22_), .A2(keyinput_74), .B1(n10158), .B2(
        keyinput_73), .ZN(n10074) );
  OAI221_X1 U10838 ( .B1(SI_22_), .B2(keyinput_74), .C1(n10158), .C2(
        keyinput_73), .A(n10074), .ZN(n10075) );
  AOI211_X1 U10839 ( .C1(SI_24_), .C2(keyinput_72), .A(n10076), .B(n10075), 
        .ZN(n10077) );
  OAI21_X1 U10840 ( .B1(SI_24_), .B2(keyinput_72), .A(n10077), .ZN(n10078) );
  OAI221_X1 U10841 ( .B1(SI_21_), .B2(keyinput_75), .C1(n10182), .C2(n10079), 
        .A(n10078), .ZN(n10080) );
  OAI211_X1 U10842 ( .C1(n10184), .C2(keyinput_78), .A(n10081), .B(n10080), 
        .ZN(n10082) );
  AOI21_X1 U10843 ( .B1(n10184), .B2(keyinput_78), .A(n10082), .ZN(n10093) );
  XNOR2_X1 U10844 ( .A(keyinput_79), .B(n10188), .ZN(n10092) );
  OAI22_X1 U10845 ( .A1(SI_12_), .A2(keyinput_84), .B1(SI_11_), .B2(
        keyinput_85), .ZN(n10083) );
  AOI221_X1 U10846 ( .B1(SI_12_), .B2(keyinput_84), .C1(keyinput_85), .C2(
        SI_11_), .A(n10083), .ZN(n10091) );
  OAI22_X1 U10847 ( .A1(n10085), .A2(keyinput_82), .B1(keyinput_83), .B2(
        SI_13_), .ZN(n10084) );
  AOI221_X1 U10848 ( .B1(n10085), .B2(keyinput_82), .C1(SI_13_), .C2(
        keyinput_83), .A(n10084), .ZN(n10088) );
  OAI22_X1 U10849 ( .A1(n10192), .A2(keyinput_81), .B1(keyinput_86), .B2(
        SI_10_), .ZN(n10086) );
  AOI221_X1 U10850 ( .B1(n10192), .B2(keyinput_81), .C1(SI_10_), .C2(
        keyinput_86), .A(n10086), .ZN(n10087) );
  OAI211_X1 U10851 ( .C1(SI_16_), .C2(keyinput_80), .A(n10088), .B(n10087), 
        .ZN(n10089) );
  AOI21_X1 U10852 ( .B1(SI_16_), .B2(keyinput_80), .A(n10089), .ZN(n10090) );
  OAI211_X1 U10853 ( .C1(n10093), .C2(n10092), .A(n10091), .B(n10090), .ZN(
        n10094) );
  OAI221_X1 U10854 ( .B1(SI_9_), .B2(n10095), .C1(n10203), .C2(keyinput_87), 
        .A(n10094), .ZN(n10096) );
  OAI221_X1 U10855 ( .B1(SI_8_), .B2(keyinput_88), .C1(n10206), .C2(n10097), 
        .A(n10096), .ZN(n10098) );
  OAI221_X1 U10856 ( .B1(SI_7_), .B2(keyinput_89), .C1(n10210), .C2(n10099), 
        .A(n10098), .ZN(n10100) );
  OAI221_X1 U10857 ( .B1(SI_6_), .B2(keyinput_90), .C1(n10213), .C2(n10101), 
        .A(n10100), .ZN(n10106) );
  OAI22_X1 U10858 ( .A1(n10215), .A2(keyinput_92), .B1(SI_5_), .B2(keyinput_91), .ZN(n10102) );
  AOI221_X1 U10859 ( .B1(n10215), .B2(keyinput_92), .C1(keyinput_91), .C2(
        SI_5_), .A(n10102), .ZN(n10105) );
  XNOR2_X1 U10860 ( .A(n10217), .B(keyinput_94), .ZN(n10104) );
  XNOR2_X1 U10861 ( .A(SI_3_), .B(keyinput_93), .ZN(n10103) );
  AOI211_X1 U10862 ( .C1(n10106), .C2(n10105), .A(n10104), .B(n10103), .ZN(
        n10107) );
  INV_X1 U10863 ( .A(n10107), .ZN(n10110) );
  OAI22_X1 U10864 ( .A1(SI_0_), .A2(keyinput_96), .B1(keyinput_95), .B2(SI_1_), 
        .ZN(n10108) );
  AOI221_X1 U10865 ( .B1(SI_0_), .B2(keyinput_96), .C1(SI_1_), .C2(keyinput_95), .A(n10108), .ZN(n10109) );
  NAND2_X1 U10866 ( .A1(n10110), .A2(n10109), .ZN(n10122) );
  OAI22_X1 U10867 ( .A1(n10112), .A2(keyinput_100), .B1(keyinput_104), .B2(
        P2_REG3_REG_3__SCAN_IN), .ZN(n10111) );
  AOI221_X1 U10868 ( .B1(n10112), .B2(keyinput_100), .C1(
        P2_REG3_REG_3__SCAN_IN), .C2(keyinput_104), .A(n10111), .ZN(n10121) );
  AOI22_X1 U10869 ( .A1(n10115), .A2(keyinput_102), .B1(n10114), .B2(
        keyinput_99), .ZN(n10113) );
  OAI221_X1 U10870 ( .B1(n10115), .B2(keyinput_102), .C1(n10114), .C2(
        keyinput_99), .A(n10113), .ZN(n10119) );
  OAI22_X1 U10871 ( .A1(P2_U3152), .A2(keyinput_98), .B1(keyinput_101), .B2(
        P2_REG3_REG_14__SCAN_IN), .ZN(n10116) );
  AOI221_X1 U10872 ( .B1(P2_U3152), .B2(keyinput_98), .C1(
        P2_REG3_REG_14__SCAN_IN), .C2(keyinput_101), .A(n10116), .ZN(n10117)
         );
  OAI21_X1 U10873 ( .B1(keyinput_103), .B2(P2_REG3_REG_10__SCAN_IN), .A(n10117), .ZN(n10118) );
  AOI211_X1 U10874 ( .C1(keyinput_103), .C2(P2_REG3_REG_10__SCAN_IN), .A(
        n10119), .B(n10118), .ZN(n10120) );
  OAI211_X1 U10875 ( .C1(n10123), .C2(n10122), .A(n10121), .B(n10120), .ZN(
        n10124) );
  OAI221_X1 U10876 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(n10125), .C1(n5949), 
        .C2(keyinput_105), .A(n10124), .ZN(n10131) );
  AOI22_X1 U10877 ( .A1(n10127), .A2(keyinput_107), .B1(keyinput_109), .B2(
        n5993), .ZN(n10126) );
  OAI221_X1 U10878 ( .B1(n10127), .B2(keyinput_107), .C1(n5993), .C2(
        keyinput_109), .A(n10126), .ZN(n10130) );
  AOI22_X1 U10879 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_108), .B1(
        P2_REG3_REG_12__SCAN_IN), .B2(keyinput_110), .ZN(n10128) );
  OAI221_X1 U10880 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_108), .C1(
        P2_REG3_REG_12__SCAN_IN), .C2(keyinput_110), .A(n10128), .ZN(n10129)
         );
  AOI211_X1 U10881 ( .C1(n10132), .C2(n10131), .A(n10130), .B(n10129), .ZN(
        n10133) );
  AOI221_X1 U10882 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(keyinput_111), .C1(
        n8993), .C2(n10134), .A(n10133), .ZN(n10135) );
  AOI221_X1 U10883 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(n10136), .C1(n10248), 
        .C2(keyinput_112), .A(n10135), .ZN(n10137) );
  AOI221_X1 U10884 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_113), .C1(
        n10251), .C2(n10138), .A(n10137), .ZN(n10140) );
  INV_X1 U10885 ( .A(P2_REG3_REG_4__SCAN_IN), .ZN(n10253) );
  NAND2_X1 U10886 ( .A1(n10253), .A2(keyinput_116), .ZN(n10139) );
  OAI221_X1 U10887 ( .B1(n10141), .B2(n10140), .C1(n10253), .C2(keyinput_116), 
        .A(n10139), .ZN(n10142) );
  OAI211_X1 U10888 ( .C1(n10259), .C2(keyinput_118), .A(n10143), .B(n10142), 
        .ZN(n10144) );
  AOI21_X1 U10889 ( .B1(n10259), .B2(keyinput_118), .A(n10144), .ZN(n10145) );
  AOI221_X1 U10890 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(keyinput_120), .C1(
        n5815), .C2(n10146), .A(n10145), .ZN(n10150) );
  OAI22_X1 U10891 ( .A1(n10148), .A2(keyinput_123), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput_122), .ZN(n10147) );
  AOI221_X1 U10892 ( .B1(n10148), .B2(keyinput_123), .C1(keyinput_122), .C2(
        P2_REG3_REG_11__SCAN_IN), .A(n10147), .ZN(n10149) );
  OAI21_X1 U10893 ( .B1(n10151), .B2(n10150), .A(n10149), .ZN(n10152) );
  AOI22_X1 U10894 ( .A1(P2_REG3_REG_26__SCAN_IN), .A2(keyinput_126), .B1(
        n10153), .B2(n10152), .ZN(n10279) );
  INV_X1 U10895 ( .A(keyinput_62), .ZN(n10273) );
  INV_X1 U10896 ( .A(keyinput_57), .ZN(n10263) );
  INV_X1 U10897 ( .A(keyinput_56), .ZN(n10261) );
  OAI22_X1 U10898 ( .A1(n5719), .A2(keyinput_53), .B1(P2_REG3_REG_20__SCAN_IN), 
        .B2(keyinput_55), .ZN(n10154) );
  AOI221_X1 U10899 ( .B1(n5719), .B2(keyinput_53), .C1(keyinput_55), .C2(
        P2_REG3_REG_20__SCAN_IN), .A(n10154), .ZN(n10257) );
  AOI22_X1 U10900 ( .A1(P2_REG3_REG_24__SCAN_IN), .A2(keyinput_51), .B1(n5911), 
        .B2(keyinput_50), .ZN(n10155) );
  OAI221_X1 U10901 ( .B1(P2_REG3_REG_24__SCAN_IN), .B2(keyinput_51), .C1(n5911), .C2(keyinput_50), .A(n10155), .ZN(n10255) );
  INV_X1 U10902 ( .A(keyinput_49), .ZN(n10250) );
  INV_X1 U10903 ( .A(keyinput_48), .ZN(n10247) );
  INV_X1 U10904 ( .A(keyinput_47), .ZN(n10245) );
  XNOR2_X1 U10905 ( .A(P2_REG3_REG_28__SCAN_IN), .B(keyinput_42), .ZN(n10243)
         );
  INV_X1 U10906 ( .A(keyinput_41), .ZN(n10236) );
  INV_X1 U10907 ( .A(keyinput_26), .ZN(n10212) );
  INV_X1 U10908 ( .A(keyinput_25), .ZN(n10209) );
  INV_X1 U10909 ( .A(keyinput_24), .ZN(n10207) );
  INV_X1 U10910 ( .A(keyinput_23), .ZN(n10204) );
  INV_X1 U10911 ( .A(keyinput_11), .ZN(n10181) );
  OAI22_X1 U10912 ( .A1(n10158), .A2(keyinput_9), .B1(n10157), .B2(keyinput_10), .ZN(n10156) );
  AOI221_X1 U10913 ( .B1(n10158), .B2(keyinput_9), .C1(keyinput_10), .C2(
        n10157), .A(n10156), .ZN(n10177) );
  INV_X1 U10914 ( .A(keyinput_7), .ZN(n10175) );
  INV_X1 U10915 ( .A(keyinput_6), .ZN(n10172) );
  INV_X1 U10916 ( .A(keyinput_2), .ZN(n10162) );
  AOI22_X1 U10917 ( .A1(P2_WR_REG_SCAN_IN), .A2(keyinput_0), .B1(SI_31_), .B2(
        keyinput_1), .ZN(n10159) );
  OAI221_X1 U10918 ( .B1(P2_WR_REG_SCAN_IN), .B2(keyinput_0), .C1(SI_31_), 
        .C2(keyinput_1), .A(n10159), .ZN(n10160) );
  AOI221_X1 U10919 ( .B1(SI_30_), .B2(n10162), .C1(n10161), .C2(keyinput_2), 
        .A(n10160), .ZN(n10167) );
  AOI22_X1 U10920 ( .A1(n10165), .A2(keyinput_4), .B1(n10164), .B2(keyinput_3), 
        .ZN(n10163) );
  OAI221_X1 U10921 ( .B1(n10165), .B2(keyinput_4), .C1(n10164), .C2(keyinput_3), .A(n10163), .ZN(n10166) );
  AOI211_X1 U10922 ( .C1(n10169), .C2(keyinput_5), .A(n10167), .B(n10166), 
        .ZN(n10168) );
  OAI21_X1 U10923 ( .B1(n10169), .B2(keyinput_5), .A(n10168), .ZN(n10170) );
  OAI221_X1 U10924 ( .B1(SI_26_), .B2(n10172), .C1(n10171), .C2(keyinput_6), 
        .A(n10170), .ZN(n10173) );
  OAI221_X1 U10925 ( .B1(SI_25_), .B2(n10175), .C1(n10174), .C2(keyinput_7), 
        .A(n10173), .ZN(n10176) );
  OAI211_X1 U10926 ( .C1(n10179), .C2(keyinput_8), .A(n10177), .B(n10176), 
        .ZN(n10178) );
  AOI21_X1 U10927 ( .B1(n10179), .B2(keyinput_8), .A(n10178), .ZN(n10180) );
  AOI221_X1 U10928 ( .B1(SI_21_), .B2(keyinput_11), .C1(n10182), .C2(n10181), 
        .A(n10180), .ZN(n10187) );
  OAI22_X1 U10929 ( .A1(n10184), .A2(keyinput_14), .B1(keyinput_12), .B2(
        SI_20_), .ZN(n10183) );
  AOI221_X1 U10930 ( .B1(n10184), .B2(keyinput_14), .C1(SI_20_), .C2(
        keyinput_12), .A(n10183), .ZN(n10185) );
  OAI21_X1 U10931 ( .B1(keyinput_13), .B2(SI_19_), .A(n10185), .ZN(n10186) );
  AOI211_X1 U10932 ( .C1(keyinput_13), .C2(SI_19_), .A(n10187), .B(n10186), 
        .ZN(n10201) );
  XNOR2_X1 U10933 ( .A(keyinput_15), .B(n10188), .ZN(n10200) );
  OAI22_X1 U10934 ( .A1(SI_14_), .A2(keyinput_18), .B1(keyinput_19), .B2(
        SI_13_), .ZN(n10189) );
  AOI221_X1 U10935 ( .B1(SI_14_), .B2(keyinput_18), .C1(SI_13_), .C2(
        keyinput_19), .A(n10189), .ZN(n10199) );
  AOI22_X1 U10936 ( .A1(n10192), .A2(keyinput_17), .B1(n10191), .B2(
        keyinput_22), .ZN(n10190) );
  OAI221_X1 U10937 ( .B1(n10192), .B2(keyinput_17), .C1(n10191), .C2(
        keyinput_22), .A(n10190), .ZN(n10197) );
  INV_X1 U10938 ( .A(SI_11_), .ZN(n10194) );
  OAI22_X1 U10939 ( .A1(n10194), .A2(keyinput_21), .B1(keyinput_20), .B2(
        SI_12_), .ZN(n10193) );
  AOI221_X1 U10940 ( .B1(n10194), .B2(keyinput_21), .C1(SI_12_), .C2(
        keyinput_20), .A(n10193), .ZN(n10195) );
  OAI21_X1 U10941 ( .B1(keyinput_16), .B2(SI_16_), .A(n10195), .ZN(n10196) );
  AOI211_X1 U10942 ( .C1(keyinput_16), .C2(SI_16_), .A(n10197), .B(n10196), 
        .ZN(n10198) );
  OAI211_X1 U10943 ( .C1(n10201), .C2(n10200), .A(n10199), .B(n10198), .ZN(
        n10202) );
  OAI221_X1 U10944 ( .B1(SI_9_), .B2(n10204), .C1(n10203), .C2(keyinput_23), 
        .A(n10202), .ZN(n10205) );
  OAI221_X1 U10945 ( .B1(SI_8_), .B2(n10207), .C1(n10206), .C2(keyinput_24), 
        .A(n10205), .ZN(n10208) );
  OAI221_X1 U10946 ( .B1(SI_7_), .B2(keyinput_25), .C1(n10210), .C2(n10209), 
        .A(n10208), .ZN(n10211) );
  OAI221_X1 U10947 ( .B1(SI_6_), .B2(keyinput_26), .C1(n10213), .C2(n10212), 
        .A(n10211), .ZN(n10221) );
  OAI22_X1 U10948 ( .A1(n10216), .A2(keyinput_27), .B1(n10215), .B2(
        keyinput_28), .ZN(n10214) );
  AOI221_X1 U10949 ( .B1(n10216), .B2(keyinput_27), .C1(keyinput_28), .C2(
        n10215), .A(n10214), .ZN(n10220) );
  XNOR2_X1 U10950 ( .A(n10217), .B(keyinput_30), .ZN(n10219) );
  XNOR2_X1 U10951 ( .A(SI_3_), .B(keyinput_29), .ZN(n10218) );
  AOI211_X1 U10952 ( .C1(n10221), .C2(n10220), .A(n10219), .B(n10218), .ZN(
        n10234) );
  XOR2_X1 U10953 ( .A(keyinput_33), .B(n5498), .Z(n10224) );
  XNOR2_X1 U10954 ( .A(SI_0_), .B(keyinput_32), .ZN(n10223) );
  XNOR2_X1 U10955 ( .A(SI_1_), .B(keyinput_31), .ZN(n10222) );
  NAND3_X1 U10956 ( .A1(n10224), .A2(n10223), .A3(n10222), .ZN(n10233) );
  OAI22_X1 U10957 ( .A1(P2_REG3_REG_14__SCAN_IN), .A2(keyinput_37), .B1(
        P2_STATE_REG_SCAN_IN), .B2(keyinput_34), .ZN(n10225) );
  AOI221_X1 U10958 ( .B1(P2_REG3_REG_14__SCAN_IN), .B2(keyinput_37), .C1(
        keyinput_34), .C2(P2_STATE_REG_SCAN_IN), .A(n10225), .ZN(n10228) );
  OAI22_X1 U10959 ( .A1(P2_REG3_REG_10__SCAN_IN), .A2(keyinput_39), .B1(
        keyinput_38), .B2(P2_REG3_REG_23__SCAN_IN), .ZN(n10226) );
  AOI221_X1 U10960 ( .B1(P2_REG3_REG_10__SCAN_IN), .B2(keyinput_39), .C1(
        P2_REG3_REG_23__SCAN_IN), .C2(keyinput_38), .A(n10226), .ZN(n10227) );
  OAI211_X1 U10961 ( .C1(P2_REG3_REG_7__SCAN_IN), .C2(keyinput_35), .A(n10228), 
        .B(n10227), .ZN(n10229) );
  AOI21_X1 U10962 ( .B1(P2_REG3_REG_7__SCAN_IN), .B2(keyinput_35), .A(n10229), 
        .ZN(n10232) );
  OAI22_X1 U10963 ( .A1(P2_REG3_REG_3__SCAN_IN), .A2(keyinput_40), .B1(
        keyinput_36), .B2(P2_REG3_REG_27__SCAN_IN), .ZN(n10230) );
  AOI221_X1 U10964 ( .B1(P2_REG3_REG_3__SCAN_IN), .B2(keyinput_40), .C1(
        P2_REG3_REG_27__SCAN_IN), .C2(keyinput_36), .A(n10230), .ZN(n10231) );
  OAI211_X1 U10965 ( .C1(n10234), .C2(n10233), .A(n10232), .B(n10231), .ZN(
        n10235) );
  OAI221_X1 U10966 ( .B1(P2_REG3_REG_19__SCAN_IN), .B2(n10236), .C1(n5949), 
        .C2(keyinput_41), .A(n10235), .ZN(n10242) );
  AOI22_X1 U10967 ( .A1(n5993), .A2(keyinput_45), .B1(n10238), .B2(keyinput_46), .ZN(n10237) );
  OAI221_X1 U10968 ( .B1(n5993), .B2(keyinput_45), .C1(n10238), .C2(
        keyinput_46), .A(n10237), .ZN(n10241) );
  AOI22_X1 U10969 ( .A1(P2_REG3_REG_1__SCAN_IN), .A2(keyinput_44), .B1(
        P2_REG3_REG_8__SCAN_IN), .B2(keyinput_43), .ZN(n10239) );
  OAI221_X1 U10970 ( .B1(P2_REG3_REG_1__SCAN_IN), .B2(keyinput_44), .C1(
        P2_REG3_REG_8__SCAN_IN), .C2(keyinput_43), .A(n10239), .ZN(n10240) );
  AOI211_X1 U10971 ( .C1(n10243), .C2(n10242), .A(n10241), .B(n10240), .ZN(
        n10244) );
  AOI221_X1 U10972 ( .B1(P2_REG3_REG_25__SCAN_IN), .B2(n10245), .C1(n8993), 
        .C2(keyinput_47), .A(n10244), .ZN(n10246) );
  AOI221_X1 U10973 ( .B1(P2_REG3_REG_16__SCAN_IN), .B2(keyinput_48), .C1(
        n10248), .C2(n10247), .A(n10246), .ZN(n10249) );
  AOI221_X1 U10974 ( .B1(P2_REG3_REG_5__SCAN_IN), .B2(keyinput_49), .C1(n10251), .C2(n10250), .A(n10249), .ZN(n10254) );
  NAND2_X1 U10975 ( .A1(n10253), .A2(keyinput_52), .ZN(n10252) );
  OAI221_X1 U10976 ( .B1(n10255), .B2(n10254), .C1(n10253), .C2(keyinput_52), 
        .A(n10252), .ZN(n10256) );
  OAI211_X1 U10977 ( .C1(n10259), .C2(keyinput_54), .A(n10257), .B(n10256), 
        .ZN(n10258) );
  AOI21_X1 U10978 ( .B1(n10259), .B2(keyinput_54), .A(n10258), .ZN(n10260) );
  AOI221_X1 U10979 ( .B1(P2_REG3_REG_13__SCAN_IN), .B2(n10261), .C1(n5815), 
        .C2(keyinput_56), .A(n10260), .ZN(n10262) );
  AOI221_X1 U10980 ( .B1(P2_REG3_REG_22__SCAN_IN), .B2(keyinput_57), .C1(
        n10264), .C2(n10263), .A(n10262), .ZN(n10270) );
  AOI22_X1 U10981 ( .A1(P2_REG3_REG_2__SCAN_IN), .A2(keyinput_59), .B1(
        P2_REG3_REG_11__SCAN_IN), .B2(keyinput_58), .ZN(n10265) );
  OAI221_X1 U10982 ( .B1(P2_REG3_REG_2__SCAN_IN), .B2(keyinput_59), .C1(
        P2_REG3_REG_11__SCAN_IN), .C2(keyinput_58), .A(n10265), .ZN(n10269) );
  OAI22_X1 U10983 ( .A1(n5684), .A2(keyinput_61), .B1(n10267), .B2(keyinput_60), .ZN(n10266) );
  AOI221_X1 U10984 ( .B1(n5684), .B2(keyinput_61), .C1(keyinput_60), .C2(
        n10267), .A(n10266), .ZN(n10268) );
  OAI21_X1 U10985 ( .B1(n10270), .B2(n10269), .A(n10268), .ZN(n10271) );
  OAI221_X1 U10986 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(n10273), .C1(n10272), 
        .C2(keyinput_62), .A(n10271), .ZN(n10275) );
  AOI21_X1 U10987 ( .B1(keyinput_63), .B2(n10275), .A(P2_REG3_REG_15__SCAN_IN), 
        .ZN(n10277) );
  INV_X1 U10988 ( .A(keyinput_63), .ZN(n10274) );
  AOI21_X1 U10989 ( .B1(n10275), .B2(n10274), .A(keyinput_127), .ZN(n10276) );
  AOI22_X1 U10990 ( .A1(keyinput_127), .A2(n10277), .B1(
        P2_REG3_REG_15__SCAN_IN), .B2(n10276), .ZN(n10278) );
  AOI221_X1 U10991 ( .B1(P2_REG3_REG_26__SCAN_IN), .B2(n10279), .C1(
        keyinput_126), .C2(n10279), .A(n10278), .ZN(n10296) );
  AOI22_X1 U10992 ( .A1(n10282), .A2(n7840), .B1(n10281), .B2(n10280), .ZN(
        n10286) );
  NAND2_X1 U10993 ( .A1(n10284), .A2(n10283), .ZN(n10285) );
  OAI211_X1 U10994 ( .C1(P2_STATE_REG_SCAN_IN), .C2(n5815), .A(n10286), .B(
        n10285), .ZN(n10292) );
  AOI211_X1 U10995 ( .C1(n10290), .C2(n10289), .A(n10288), .B(n10287), .ZN(
        n10291) );
  AOI211_X1 U10996 ( .C1(n10294), .C2(n10293), .A(n10292), .B(n10291), .ZN(
        n10295) );
  XNOR2_X1 U10997 ( .A(n10296), .B(n10295), .ZN(P2_U3236) );
  XOR2_X1 U10998 ( .A(P2_ADDR_REG_0__SCAN_IN), .B(P1_ADDR_REG_0__SCAN_IN), .Z(
        ADD_1071_U46) );
  NAND3_X1 U10999 ( .A1(P1_ADDR_REG_1__SCAN_IN), .A2(P2_ADDR_REG_0__SCAN_IN), 
        .A3(P1_ADDR_REG_0__SCAN_IN), .ZN(n10299) );
  AOI21_X1 U11000 ( .B1(P2_ADDR_REG_0__SCAN_IN), .B2(P1_ADDR_REG_0__SCAN_IN), 
        .A(P1_ADDR_REG_1__SCAN_IN), .ZN(n10301) );
  INV_X1 U11001 ( .A(n10301), .ZN(n10297) );
  NAND2_X1 U11002 ( .A1(n10299), .A2(n10297), .ZN(n10298) );
  XNOR2_X1 U11003 ( .A(P2_ADDR_REG_1__SCAN_IN), .B(n10298), .ZN(ADD_1071_U5)
         );
  XOR2_X1 U11004 ( .A(P1_ADDR_REG_2__SCAN_IN), .B(P2_ADDR_REG_2__SCAN_IN), .Z(
        n10303) );
  INV_X1 U11005 ( .A(P2_ADDR_REG_1__SCAN_IN), .ZN(n10300) );
  OAI21_X1 U11006 ( .B1(n10301), .B2(n10300), .A(n10299), .ZN(n10302) );
  XOR2_X1 U11007 ( .A(n10303), .B(n10302), .Z(ADD_1071_U54) );
  XOR2_X1 U11008 ( .A(P2_ADDR_REG_3__SCAN_IN), .B(P1_ADDR_REG_3__SCAN_IN), .Z(
        n10307) );
  NAND2_X1 U11009 ( .A1(P1_ADDR_REG_2__SCAN_IN), .A2(P2_ADDR_REG_2__SCAN_IN), 
        .ZN(n10305) );
  NAND2_X1 U11010 ( .A1(n10303), .A2(n10302), .ZN(n10304) );
  NAND2_X1 U11011 ( .A1(n10305), .A2(n10304), .ZN(n10306) );
  XOR2_X1 U11012 ( .A(n10307), .B(n10306), .Z(ADD_1071_U53) );
  XNOR2_X1 U11013 ( .A(P1_ADDR_REG_4__SCAN_IN), .B(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10311) );
  NAND2_X1 U11014 ( .A1(P2_ADDR_REG_3__SCAN_IN), .A2(P1_ADDR_REG_3__SCAN_IN), 
        .ZN(n10309) );
  NAND2_X1 U11015 ( .A1(n10307), .A2(n10306), .ZN(n10308) );
  NAND2_X1 U11016 ( .A1(n10309), .A2(n10308), .ZN(n10310) );
  XNOR2_X1 U11017 ( .A(n10311), .B(n10310), .ZN(ADD_1071_U52) );
  NOR2_X1 U11018 ( .A1(P1_ADDR_REG_4__SCAN_IN), .A2(P2_ADDR_REG_4__SCAN_IN), 
        .ZN(n10313) );
  NOR2_X1 U11019 ( .A1(n10311), .A2(n10310), .ZN(n10312) );
  NOR2_X1 U11020 ( .A1(n10313), .A2(n10312), .ZN(n10314) );
  NOR2_X1 U11021 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10314), .ZN(n10318) );
  AND2_X1 U11022 ( .A1(P1_ADDR_REG_5__SCAN_IN), .A2(n10314), .ZN(n10316) );
  NOR2_X1 U11023 ( .A1(n10318), .A2(n10316), .ZN(n10315) );
  XOR2_X1 U11024 ( .A(P2_ADDR_REG_5__SCAN_IN), .B(n10315), .Z(ADD_1071_U51) );
  NOR2_X1 U11025 ( .A1(P2_ADDR_REG_5__SCAN_IN), .A2(n10316), .ZN(n10317) );
  XOR2_X1 U11026 ( .A(P1_ADDR_REG_6__SCAN_IN), .B(n10319), .Z(n10320) );
  XOR2_X1 U11027 ( .A(P2_ADDR_REG_6__SCAN_IN), .B(n10320), .Z(ADD_1071_U50) );
  NAND2_X1 U11028 ( .A1(P1_ADDR_REG_6__SCAN_IN), .A2(n10319), .ZN(n10322) );
  NAND2_X1 U11029 ( .A1(P2_ADDR_REG_6__SCAN_IN), .A2(n10320), .ZN(n10321) );
  NAND2_X1 U11030 ( .A1(n10322), .A2(n10321), .ZN(n10323) );
  XOR2_X1 U11031 ( .A(P1_ADDR_REG_7__SCAN_IN), .B(n10323), .Z(n10324) );
  XOR2_X1 U11032 ( .A(P2_ADDR_REG_7__SCAN_IN), .B(n10324), .Z(ADD_1071_U49) );
  NAND2_X1 U11033 ( .A1(P1_ADDR_REG_7__SCAN_IN), .A2(n10323), .ZN(n10326) );
  NAND2_X1 U11034 ( .A1(P2_ADDR_REG_7__SCAN_IN), .A2(n10324), .ZN(n10325) );
  NAND2_X1 U11035 ( .A1(n10326), .A2(n10325), .ZN(n10327) );
  XOR2_X1 U11036 ( .A(P1_ADDR_REG_8__SCAN_IN), .B(n10327), .Z(n10328) );
  XOR2_X1 U11037 ( .A(P2_ADDR_REG_8__SCAN_IN), .B(n10328), .Z(ADD_1071_U48) );
  NAND2_X1 U11038 ( .A1(P1_ADDR_REG_8__SCAN_IN), .A2(n10327), .ZN(n10330) );
  NAND2_X1 U11039 ( .A1(P2_ADDR_REG_8__SCAN_IN), .A2(n10328), .ZN(n10329) );
  NAND2_X1 U11040 ( .A1(n10330), .A2(n10329), .ZN(n10331) );
  XOR2_X1 U11041 ( .A(P1_ADDR_REG_9__SCAN_IN), .B(n10331), .Z(n10332) );
  XOR2_X1 U11042 ( .A(P2_ADDR_REG_9__SCAN_IN), .B(n10332), .Z(ADD_1071_U47) );
  XOR2_X1 U11043 ( .A(P2_ADDR_REG_10__SCAN_IN), .B(P1_ADDR_REG_10__SCAN_IN), 
        .Z(n10336) );
  NAND2_X1 U11044 ( .A1(P1_ADDR_REG_9__SCAN_IN), .A2(n10331), .ZN(n10334) );
  NAND2_X1 U11045 ( .A1(P2_ADDR_REG_9__SCAN_IN), .A2(n10332), .ZN(n10333) );
  NAND2_X1 U11046 ( .A1(n10334), .A2(n10333), .ZN(n10335) );
  XOR2_X1 U11047 ( .A(n10336), .B(n10335), .Z(ADD_1071_U63) );
  XOR2_X1 U11048 ( .A(P2_ADDR_REG_11__SCAN_IN), .B(P1_ADDR_REG_11__SCAN_IN), 
        .Z(n10340) );
  NAND2_X1 U11049 ( .A1(P2_ADDR_REG_10__SCAN_IN), .A2(P1_ADDR_REG_10__SCAN_IN), 
        .ZN(n10338) );
  NAND2_X1 U11050 ( .A1(n10336), .A2(n10335), .ZN(n10337) );
  NAND2_X1 U11051 ( .A1(n10338), .A2(n10337), .ZN(n10339) );
  XOR2_X1 U11052 ( .A(n10340), .B(n10339), .Z(ADD_1071_U62) );
  NAND2_X1 U11053 ( .A1(P2_ADDR_REG_11__SCAN_IN), .A2(P1_ADDR_REG_11__SCAN_IN), 
        .ZN(n10342) );
  NAND2_X1 U11054 ( .A1(n10340), .A2(n10339), .ZN(n10341) );
  NAND2_X1 U11055 ( .A1(n10342), .A2(n10341), .ZN(n10344) );
  XNOR2_X1 U11056 ( .A(P2_ADDR_REG_12__SCAN_IN), .B(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10343) );
  XNOR2_X1 U11057 ( .A(n10344), .B(n10343), .ZN(ADD_1071_U61) );
  NOR2_X1 U11058 ( .A1(P2_ADDR_REG_12__SCAN_IN), .A2(P1_ADDR_REG_12__SCAN_IN), 
        .ZN(n10346) );
  XNOR2_X1 U11059 ( .A(P2_ADDR_REG_13__SCAN_IN), .B(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10347) );
  XNOR2_X1 U11060 ( .A(n10348), .B(n10347), .ZN(ADD_1071_U60) );
  NOR2_X1 U11061 ( .A1(P2_ADDR_REG_13__SCAN_IN), .A2(P1_ADDR_REG_13__SCAN_IN), 
        .ZN(n10350) );
  XNOR2_X1 U11062 ( .A(P2_ADDR_REG_14__SCAN_IN), .B(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10351) );
  XNOR2_X1 U11063 ( .A(n10352), .B(n10351), .ZN(ADD_1071_U59) );
  NOR2_X1 U11064 ( .A1(P2_ADDR_REG_14__SCAN_IN), .A2(P1_ADDR_REG_14__SCAN_IN), 
        .ZN(n10354) );
  NOR2_X1 U11065 ( .A1(n10352), .A2(n10351), .ZN(n10353) );
  NOR2_X1 U11066 ( .A1(n10354), .A2(n10353), .ZN(n10356) );
  XNOR2_X1 U11067 ( .A(P2_ADDR_REG_15__SCAN_IN), .B(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10355) );
  XNOR2_X1 U11068 ( .A(n10356), .B(n10355), .ZN(ADD_1071_U58) );
  NOR2_X1 U11069 ( .A1(P2_ADDR_REG_15__SCAN_IN), .A2(P1_ADDR_REG_15__SCAN_IN), 
        .ZN(n10358) );
  NOR2_X1 U11070 ( .A1(n10356), .A2(n10355), .ZN(n10357) );
  NOR2_X1 U11071 ( .A1(n10358), .A2(n10357), .ZN(n10360) );
  XNOR2_X1 U11072 ( .A(P2_ADDR_REG_16__SCAN_IN), .B(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10359) );
  XNOR2_X1 U11073 ( .A(n10360), .B(n10359), .ZN(ADD_1071_U57) );
  NOR2_X1 U11074 ( .A1(P2_ADDR_REG_16__SCAN_IN), .A2(P1_ADDR_REG_16__SCAN_IN), 
        .ZN(n10362) );
  NOR2_X1 U11075 ( .A1(n10360), .A2(n10359), .ZN(n10361) );
  NOR2_X1 U11076 ( .A1(n10362), .A2(n10361), .ZN(n10364) );
  XNOR2_X1 U11077 ( .A(P2_ADDR_REG_17__SCAN_IN), .B(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10363) );
  XNOR2_X1 U11078 ( .A(n10364), .B(n10363), .ZN(ADD_1071_U56) );
  NOR2_X1 U11079 ( .A1(P2_ADDR_REG_17__SCAN_IN), .A2(P1_ADDR_REG_17__SCAN_IN), 
        .ZN(n10366) );
  NOR2_X1 U11080 ( .A1(n10364), .A2(n10363), .ZN(n10365) );
  NOR2_X1 U11081 ( .A1(n10366), .A2(n10365), .ZN(n10367) );
  NOR2_X1 U11082 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10367), .ZN(n10370) );
  AND2_X1 U11083 ( .A1(P2_ADDR_REG_18__SCAN_IN), .A2(n10367), .ZN(n10369) );
  NOR2_X1 U11084 ( .A1(n10370), .A2(n10369), .ZN(n10368) );
  XOR2_X1 U11085 ( .A(P1_ADDR_REG_18__SCAN_IN), .B(n10368), .Z(ADD_1071_U55)
         );
  NOR2_X1 U11086 ( .A1(P1_ADDR_REG_18__SCAN_IN), .A2(n10369), .ZN(n10371) );
  NOR2_X1 U11087 ( .A1(n10371), .A2(n10370), .ZN(n10373) );
  XNOR2_X1 U11088 ( .A(P2_ADDR_REG_19__SCAN_IN), .B(P1_ADDR_REG_19__SCAN_IN), 
        .ZN(n10372) );
  XNOR2_X1 U11089 ( .A(n10373), .B(n10372), .ZN(ADD_1071_U4) );
  INV_X1 U11090 ( .A(n10374), .ZN(n10378) );
  AOI21_X1 U11091 ( .B1(P1_IR_REG_0__SCAN_IN), .B2(n10376), .A(n10375), .ZN(
        n10377) );
  AOI21_X1 U11092 ( .B1(n10379), .B2(n10378), .A(n10377), .ZN(n10381) );
  OAI22_X1 U11093 ( .A1(n10381), .A2(n5192), .B1(P1_REG1_REG_0__SCAN_IN), .B2(
        n10380), .ZN(n10385) );
  NAND3_X1 U11094 ( .A1(n4860), .A2(n10383), .A3(n10382), .ZN(n10384) );
  NAND2_X1 U11095 ( .A1(n10385), .A2(n10384), .ZN(n10388) );
  AOI22_X1 U11096 ( .A1(n10386), .A2(P1_ADDR_REG_0__SCAN_IN), .B1(
        P1_REG3_REG_0__SCAN_IN), .B2(P1_U3084), .ZN(n10387) );
  OAI21_X1 U11097 ( .B1(n10389), .B2(n10388), .A(n10387), .ZN(P1_U3241) );
  INV_X1 U11098 ( .A(P1_ADDR_REG_9__SCAN_IN), .ZN(n10390) );
  OAI22_X1 U11099 ( .A1(n10393), .A2(n10392), .B1(n10391), .B2(n10390), .ZN(
        n10394) );
  INV_X1 U11100 ( .A(n10394), .ZN(n10407) );
  NAND2_X1 U11101 ( .A1(P1_REG3_REG_9__SCAN_IN), .A2(P1_U3084), .ZN(n10406) );
  OAI21_X1 U11102 ( .B1(n10397), .B2(n10396), .A(n10395), .ZN(n10399) );
  NAND2_X1 U11103 ( .A1(n10399), .A2(n10398), .ZN(n10405) );
  OAI211_X1 U11104 ( .C1(n10403), .C2(n10402), .A(n10401), .B(n10400), .ZN(
        n10404) );
  NAND4_X1 U11105 ( .A1(n10407), .A2(n10406), .A3(n10405), .A4(n10404), .ZN(
        P1_U3250) );
  NOR2_X1 U11106 ( .A1(n10409), .A2(n10408), .ZN(n10412) );
  INV_X1 U11107 ( .A(P2_D_REG_0__SCAN_IN), .ZN(n10411) );
  AOI22_X1 U11108 ( .A1(n10413), .A2(n10412), .B1(n10411), .B2(n10410), .ZN(
        P2_U3437) );
  AOI22_X1 U11109 ( .A1(n10480), .A2(P2_REG2_REG_0__SCAN_IN), .B1(
        P2_REG1_REG_0__SCAN_IN), .B2(n10450), .ZN(n10420) );
  AOI22_X1 U11110 ( .A1(n10486), .A2(P2_ADDR_REG_0__SCAN_IN), .B1(
        P2_REG3_REG_0__SCAN_IN), .B2(P2_U3152), .ZN(n10419) );
  OAI21_X1 U11111 ( .B1(n10481), .B2(P2_REG1_REG_0__SCAN_IN), .A(n10414), .ZN(
        n10417) );
  NOR2_X1 U11112 ( .A1(n10415), .A2(P2_REG2_REG_0__SCAN_IN), .ZN(n10416) );
  OAI21_X1 U11113 ( .B1(n10417), .B2(n10416), .A(P2_IR_REG_0__SCAN_IN), .ZN(
        n10418) );
  OAI211_X1 U11114 ( .C1(P2_IR_REG_0__SCAN_IN), .C2(n10420), .A(n10419), .B(
        n10418), .ZN(P2_U3245) );
  AOI22_X1 U11115 ( .A1(n10486), .A2(P2_ADDR_REG_1__SCAN_IN), .B1(
        P2_REG3_REG_1__SCAN_IN), .B2(P2_U3152), .ZN(n10434) );
  NAND2_X1 U11116 ( .A1(n10478), .A2(n10421), .ZN(n10433) );
  NOR2_X1 U11117 ( .A1(n10427), .A2(n10422), .ZN(n10425) );
  OAI211_X1 U11118 ( .C1(n10425), .C2(n10424), .A(n10480), .B(n10423), .ZN(
        n10432) );
  NOR2_X1 U11119 ( .A1(n10427), .A2(n10426), .ZN(n10430) );
  OAI211_X1 U11120 ( .C1(n10430), .C2(n10429), .A(n10450), .B(n10428), .ZN(
        n10431) );
  NAND4_X1 U11121 ( .A1(n10434), .A2(n10433), .A3(n10432), .A4(n10431), .ZN(
        P2_U3246) );
  AOI22_X1 U11122 ( .A1(n10486), .A2(P2_ADDR_REG_2__SCAN_IN), .B1(
        P2_REG3_REG_2__SCAN_IN), .B2(P2_U3152), .ZN(n10446) );
  INV_X1 U11123 ( .A(n10435), .ZN(n10436) );
  NAND2_X1 U11124 ( .A1(n10478), .A2(n10436), .ZN(n10445) );
  OAI211_X1 U11125 ( .C1(n10439), .C2(n10438), .A(n10450), .B(n10437), .ZN(
        n10444) );
  OAI211_X1 U11126 ( .C1(n10442), .C2(n10441), .A(n10480), .B(n10440), .ZN(
        n10443) );
  NAND4_X1 U11127 ( .A1(n10446), .A2(n10445), .A3(n10444), .A4(n10443), .ZN(
        P2_U3247) );
  AOI22_X1 U11128 ( .A1(n10486), .A2(P2_ADDR_REG_3__SCAN_IN), .B1(
        P2_REG3_REG_3__SCAN_IN), .B2(P2_U3152), .ZN(n10459) );
  NAND2_X1 U11129 ( .A1(n10478), .A2(n10448), .ZN(n10458) );
  OAI211_X1 U11130 ( .C1(n10452), .C2(n10451), .A(n10450), .B(n10449), .ZN(
        n10457) );
  OAI211_X1 U11131 ( .C1(n10455), .C2(n10454), .A(n10480), .B(n10453), .ZN(
        n10456) );
  NAND4_X1 U11132 ( .A1(n10459), .A2(n10458), .A3(n10457), .A4(n10456), .ZN(
        P2_U3248) );
  INV_X1 U11133 ( .A(n10460), .ZN(n10461) );
  AOI21_X1 U11134 ( .B1(n10486), .B2(P2_ADDR_REG_5__SCAN_IN), .A(n10461), .ZN(
        n10473) );
  NAND2_X1 U11135 ( .A1(n10478), .A2(n10462), .ZN(n10472) );
  AOI211_X1 U11136 ( .C1(n10465), .C2(n10464), .A(n10463), .B(n10481), .ZN(
        n10466) );
  INV_X1 U11137 ( .A(n10466), .ZN(n10471) );
  OAI211_X1 U11138 ( .C1(n10469), .C2(n10468), .A(n10480), .B(n10467), .ZN(
        n10470) );
  NAND4_X1 U11139 ( .A1(n10473), .A2(n10472), .A3(n10471), .A4(n10470), .ZN(
        P2_U3250) );
  XOR2_X1 U11140 ( .A(n10474), .B(n10477), .Z(n10475) );
  XNOR2_X1 U11141 ( .A(n10476), .B(n10475), .ZN(n10479) );
  AOI22_X1 U11142 ( .A1(n10480), .A2(n10479), .B1(n10478), .B2(n10477), .ZN(
        n10490) );
  AOI211_X1 U11143 ( .C1(n10484), .C2(n10483), .A(n10482), .B(n10481), .ZN(
        n10485) );
  INV_X1 U11144 ( .A(n10485), .ZN(n10488) );
  NAND2_X1 U11145 ( .A1(n10486), .A2(P2_ADDR_REG_6__SCAN_IN), .ZN(n10487) );
  NAND4_X1 U11146 ( .A1(n10490), .A2(n10489), .A3(n10488), .A4(n10487), .ZN(
        P2_U3251) );
  XNOR2_X1 U11147 ( .A(P1_RD_REG_SCAN_IN), .B(P2_RD_REG_SCAN_IN), .ZN(U126) );
  NOR2_X1 U11148 ( .A1(n10491), .A2(n10618), .ZN(n10492) );
  NOR2_X1 U11149 ( .A1(n10493), .A2(n10492), .ZN(n10497) );
  NAND2_X1 U11150 ( .A1(n10494), .A2(n10632), .ZN(n10496) );
  AND4_X1 U11151 ( .A1(n10498), .A2(n10497), .A3(n10496), .A4(n10495), .ZN(
        n10501) );
  INV_X1 U11152 ( .A(P1_REG1_REG_1__SCAN_IN), .ZN(n10499) );
  AOI22_X1 U11153 ( .A1(n10634), .A2(n10501), .B1(n10499), .B2(n10633), .ZN(
        P1_U3524) );
  INV_X1 U11154 ( .A(P1_REG0_REG_1__SCAN_IN), .ZN(n10500) );
  AOI22_X1 U11155 ( .A1(n10637), .A2(n10501), .B1(n10500), .B2(n10635), .ZN(
        P1_U3457) );
  INV_X1 U11156 ( .A(n10502), .ZN(n10508) );
  OR3_X1 U11157 ( .A1(n10503), .A2(n5212), .A3(n10693), .ZN(n10504) );
  OAI21_X1 U11158 ( .B1(n10505), .B2(n10691), .A(n10504), .ZN(n10507) );
  AOI211_X1 U11159 ( .C1(n10697), .C2(n10508), .A(n10507), .B(n10506), .ZN(
        n10509) );
  AOI22_X1 U11160 ( .A1(n10701), .A2(n10509), .B1(n6649), .B2(n10699), .ZN(
        P2_U3521) );
  AOI22_X1 U11161 ( .A1(n10613), .A2(n10509), .B1(n5529), .B2(n10702), .ZN(
        P2_U3454) );
  NAND2_X1 U11162 ( .A1(n10510), .A2(n10617), .ZN(n10511) );
  OAI21_X1 U11163 ( .B1(n10512), .B2(n10618), .A(n10511), .ZN(n10514) );
  AOI211_X1 U11164 ( .C1(n10632), .C2(n10515), .A(n10514), .B(n10513), .ZN(
        n10517) );
  AOI22_X1 U11165 ( .A1(n10634), .A2(n10517), .B1(n6371), .B2(n10633), .ZN(
        P1_U3525) );
  INV_X1 U11166 ( .A(P1_REG0_REG_2__SCAN_IN), .ZN(n10516) );
  AOI22_X1 U11167 ( .A1(n10637), .A2(n10517), .B1(n10516), .B2(n10635), .ZN(
        P1_U3460) );
  NAND3_X1 U11168 ( .A1(n10519), .A2(n10518), .A3(n5299), .ZN(n10520) );
  OAI21_X1 U11169 ( .B1(n10521), .B2(n10691), .A(n10520), .ZN(n10523) );
  AOI211_X1 U11170 ( .C1(n10655), .C2(n10524), .A(n10523), .B(n10522), .ZN(
        n10527) );
  AOI22_X1 U11171 ( .A1(n10701), .A2(n10527), .B1(n10525), .B2(n10699), .ZN(
        P2_U3522) );
  INV_X1 U11172 ( .A(P2_REG0_REG_2__SCAN_IN), .ZN(n10526) );
  AOI22_X1 U11173 ( .A1(n10613), .A2(n10527), .B1(n10526), .B2(n10702), .ZN(
        P2_U3457) );
  AOI22_X1 U11174 ( .A1(n10529), .A2(n10617), .B1(n10578), .B2(n10528), .ZN(
        n10530) );
  OAI211_X1 U11175 ( .C1(n10532), .C2(n10582), .A(n10531), .B(n10530), .ZN(
        n10533) );
  INV_X1 U11176 ( .A(n10533), .ZN(n10535) );
  AOI22_X1 U11177 ( .A1(n10634), .A2(n10535), .B1(n6372), .B2(n10633), .ZN(
        P1_U3527) );
  INV_X1 U11178 ( .A(P1_REG0_REG_4__SCAN_IN), .ZN(n10534) );
  AOI22_X1 U11179 ( .A1(n10637), .A2(n10535), .B1(n10534), .B2(n10635), .ZN(
        P1_U3466) );
  INV_X1 U11180 ( .A(n10536), .ZN(n10541) );
  OAI22_X1 U11181 ( .A1(n10538), .A2(n10693), .B1(n10537), .B2(n10691), .ZN(
        n10540) );
  AOI211_X1 U11182 ( .C1(n10541), .C2(n10697), .A(n10540), .B(n10539), .ZN(
        n10544) );
  AOI22_X1 U11183 ( .A1(n10701), .A2(n10544), .B1(n10542), .B2(n10699), .ZN(
        P2_U3524) );
  INV_X1 U11184 ( .A(P2_REG0_REG_4__SCAN_IN), .ZN(n10543) );
  AOI22_X1 U11185 ( .A1(n10613), .A2(n10544), .B1(n10543), .B2(n10702), .ZN(
        P2_U3463) );
  OAI21_X1 U11186 ( .B1(n10546), .B2(n10691), .A(n10545), .ZN(n10548) );
  AOI211_X1 U11187 ( .C1(n10549), .C2(n10697), .A(n10548), .B(n10547), .ZN(
        n10552) );
  AOI22_X1 U11188 ( .A1(n10701), .A2(n10552), .B1(n10550), .B2(n10699), .ZN(
        P2_U3525) );
  INV_X1 U11189 ( .A(P2_REG0_REG_5__SCAN_IN), .ZN(n10551) );
  AOI22_X1 U11190 ( .A1(n10613), .A2(n10552), .B1(n10551), .B2(n10702), .ZN(
        P2_U3466) );
  OAI22_X1 U11191 ( .A1(n10554), .A2(n10597), .B1(n10553), .B2(n10618), .ZN(
        n10557) );
  INV_X1 U11192 ( .A(n10555), .ZN(n10556) );
  AOI211_X1 U11193 ( .C1(n10632), .C2(n10558), .A(n10557), .B(n10556), .ZN(
        n10560) );
  INV_X1 U11194 ( .A(P1_REG1_REG_6__SCAN_IN), .ZN(n10559) );
  AOI22_X1 U11195 ( .A1(n10634), .A2(n10560), .B1(n10559), .B2(n10633), .ZN(
        P1_U3529) );
  AOI22_X1 U11196 ( .A1(n10637), .A2(n10560), .B1(n7039), .B2(n10635), .ZN(
        P1_U3472) );
  NOR2_X1 U11197 ( .A1(n10561), .A2(n10673), .ZN(n10566) );
  OAI22_X1 U11198 ( .A1(n10563), .A2(n10693), .B1(n10562), .B2(n10691), .ZN(
        n10565) );
  AOI211_X1 U11199 ( .C1(n10566), .C2(n7338), .A(n10565), .B(n10564), .ZN(
        n10569) );
  AOI22_X1 U11200 ( .A1(n10701), .A2(n10569), .B1(n10567), .B2(n10699), .ZN(
        P2_U3526) );
  INV_X1 U11201 ( .A(P2_REG0_REG_6__SCAN_IN), .ZN(n10568) );
  AOI22_X1 U11202 ( .A1(n10613), .A2(n10569), .B1(n10568), .B2(n10702), .ZN(
        P2_U3469) );
  OAI22_X1 U11203 ( .A1(n10571), .A2(n10693), .B1(n10570), .B2(n10691), .ZN(
        n10573) );
  AOI211_X1 U11204 ( .C1(n10697), .C2(n10574), .A(n10573), .B(n10572), .ZN(
        n10576) );
  AOI22_X1 U11205 ( .A1(n10701), .A2(n10576), .B1(n6652), .B2(n10699), .ZN(
        P2_U3527) );
  INV_X1 U11206 ( .A(P2_REG0_REG_7__SCAN_IN), .ZN(n10575) );
  AOI22_X1 U11207 ( .A1(n10613), .A2(n10576), .B1(n10575), .B2(n10702), .ZN(
        P2_U3472) );
  AOI22_X1 U11208 ( .A1(n10579), .A2(n10617), .B1(n10578), .B2(n10577), .ZN(
        n10580) );
  OAI211_X1 U11209 ( .C1(n10583), .C2(n10582), .A(n10581), .B(n10580), .ZN(
        n10584) );
  INV_X1 U11210 ( .A(n10584), .ZN(n10585) );
  AOI22_X1 U11211 ( .A1(n10634), .A2(n10585), .B1(n6369), .B2(n10633), .ZN(
        P1_U3531) );
  AOI22_X1 U11212 ( .A1(n10637), .A2(n10585), .B1(n7190), .B2(n10635), .ZN(
        P1_U3478) );
  NOR2_X1 U11213 ( .A1(n10586), .A2(n10673), .ZN(n10591) );
  OAI21_X1 U11214 ( .B1(n10588), .B2(n10691), .A(n10587), .ZN(n10590) );
  AOI211_X1 U11215 ( .C1(n10591), .C2(n7491), .A(n10590), .B(n10589), .ZN(
        n10594) );
  AOI22_X1 U11216 ( .A1(n10701), .A2(n10594), .B1(n10592), .B2(n10699), .ZN(
        P2_U3528) );
  INV_X1 U11217 ( .A(P2_REG0_REG_8__SCAN_IN), .ZN(n10593) );
  AOI22_X1 U11218 ( .A1(n10613), .A2(n10594), .B1(n10593), .B2(n10702), .ZN(
        P2_U3475) );
  INV_X1 U11219 ( .A(n10595), .ZN(n10601) );
  OAI22_X1 U11220 ( .A1(n10598), .A2(n10597), .B1(n10596), .B2(n10618), .ZN(
        n10600) );
  AOI211_X1 U11221 ( .C1(n10632), .C2(n10601), .A(n10600), .B(n10599), .ZN(
        n10604) );
  AOI22_X1 U11222 ( .A1(n10634), .A2(n10604), .B1(n10602), .B2(n10633), .ZN(
        P1_U3532) );
  INV_X1 U11223 ( .A(P1_REG0_REG_9__SCAN_IN), .ZN(n10603) );
  AOI22_X1 U11224 ( .A1(n10637), .A2(n10604), .B1(n10603), .B2(n10635), .ZN(
        P1_U3481) );
  OAI22_X1 U11225 ( .A1(n10606), .A2(n10693), .B1(n5121), .B2(n10691), .ZN(
        n10608) );
  AOI211_X1 U11226 ( .C1(n10655), .C2(n10609), .A(n10608), .B(n10607), .ZN(
        n10612) );
  AOI22_X1 U11227 ( .A1(n10701), .A2(n10612), .B1(n10610), .B2(n10699), .ZN(
        P2_U3529) );
  INV_X1 U11228 ( .A(P2_REG0_REG_9__SCAN_IN), .ZN(n10611) );
  AOI22_X1 U11229 ( .A1(n10613), .A2(n10612), .B1(n10611), .B2(n10702), .ZN(
        P2_U3478) );
  XNOR2_X1 U11230 ( .A(n10614), .B(n10619), .ZN(n10646) );
  OAI211_X1 U11231 ( .C1(n5187), .C2(n5188), .A(n10617), .B(n10616), .ZN(
        n10642) );
  OAI21_X1 U11232 ( .B1(n5187), .B2(n10618), .A(n10642), .ZN(n10631) );
  XNOR2_X1 U11233 ( .A(n10620), .B(n10619), .ZN(n10627) );
  AOI22_X1 U11234 ( .A1(n10624), .A2(n10623), .B1(n10622), .B2(n10621), .ZN(
        n10625) );
  OAI21_X1 U11235 ( .B1(n10627), .B2(n10626), .A(n10625), .ZN(n10628) );
  AOI21_X1 U11236 ( .B1(n10646), .B2(n10629), .A(n10628), .ZN(n10649) );
  INV_X1 U11237 ( .A(n10649), .ZN(n10630) );
  AOI211_X1 U11238 ( .C1(n10632), .C2(n10646), .A(n10631), .B(n10630), .ZN(
        n10636) );
  AOI22_X1 U11239 ( .A1(n10634), .A2(n10636), .B1(n6368), .B2(n10633), .ZN(
        P1_U3533) );
  AOI22_X1 U11240 ( .A1(n10637), .A2(n10636), .B1(n7525), .B2(n10635), .ZN(
        P1_U3484) );
  AOI222_X1 U11241 ( .A1(n10641), .A2(n10640), .B1(n10639), .B2(n10638), .C1(
        P1_REG2_REG_10__SCAN_IN), .C2(n9896), .ZN(n10648) );
  INV_X1 U11242 ( .A(n10642), .ZN(n10643) );
  AOI22_X1 U11243 ( .A1(n10646), .A2(n10645), .B1(n10644), .B2(n10643), .ZN(
        n10647) );
  OAI211_X1 U11244 ( .C1(n9896), .C2(n10649), .A(n10648), .B(n10647), .ZN(
        P1_U3281) );
  OAI22_X1 U11245 ( .A1(n10651), .A2(n10693), .B1(n10650), .B2(n10691), .ZN(
        n10653) );
  AOI211_X1 U11246 ( .C1(n10655), .C2(n10654), .A(n10653), .B(n10652), .ZN(
        n10657) );
  AOI22_X1 U11247 ( .A1(n10701), .A2(n10657), .B1(n6711), .B2(n10699), .ZN(
        P2_U3530) );
  INV_X1 U11248 ( .A(P2_REG0_REG_10__SCAN_IN), .ZN(n10656) );
  AOI22_X1 U11249 ( .A1(n10613), .A2(n10657), .B1(n10656), .B2(n10702), .ZN(
        P2_U3481) );
  OAI21_X1 U11250 ( .B1(n10659), .B2(n10691), .A(n10658), .ZN(n10660) );
  AOI21_X1 U11251 ( .B1(n10661), .B2(n10697), .A(n10660), .ZN(n10663) );
  AND2_X1 U11252 ( .A1(n10663), .A2(n10662), .ZN(n10665) );
  AOI22_X1 U11253 ( .A1(n10701), .A2(n10665), .B1(n6869), .B2(n10699), .ZN(
        P2_U3531) );
  INV_X1 U11254 ( .A(P2_REG0_REG_11__SCAN_IN), .ZN(n10664) );
  AOI22_X1 U11255 ( .A1(n10613), .A2(n10665), .B1(n10664), .B2(n10702), .ZN(
        P2_U3484) );
  OAI22_X1 U11256 ( .A1(n10666), .A2(n10693), .B1(n5204), .B2(n10691), .ZN(
        n10667) );
  AOI211_X1 U11257 ( .C1(n10669), .C2(n10697), .A(n10668), .B(n10667), .ZN(
        n10672) );
  AOI22_X1 U11258 ( .A1(n10701), .A2(n10672), .B1(n10670), .B2(n10699), .ZN(
        P2_U3532) );
  INV_X1 U11259 ( .A(P2_REG0_REG_12__SCAN_IN), .ZN(n10671) );
  AOI22_X1 U11260 ( .A1(n10613), .A2(n10672), .B1(n10671), .B2(n10702), .ZN(
        P2_U3487) );
  NOR2_X1 U11261 ( .A1(n10674), .A2(n10673), .ZN(n10679) );
  OAI22_X1 U11262 ( .A1(n10675), .A2(n10693), .B1(n5203), .B2(n10691), .ZN(
        n10676) );
  AOI211_X1 U11263 ( .C1(n10679), .C2(n10678), .A(n10677), .B(n10676), .ZN(
        n10682) );
  AOI22_X1 U11264 ( .A1(n10701), .A2(n10682), .B1(n10680), .B2(n10699), .ZN(
        P2_U3533) );
  INV_X1 U11265 ( .A(P2_REG0_REG_13__SCAN_IN), .ZN(n10681) );
  AOI22_X1 U11266 ( .A1(n10613), .A2(n10682), .B1(n10681), .B2(n10702), .ZN(
        P2_U3490) );
  OAI22_X1 U11267 ( .A1(n10684), .A2(n10693), .B1(n10683), .B2(n10691), .ZN(
        n10685) );
  AOI211_X1 U11268 ( .C1(n10687), .C2(n10697), .A(n10686), .B(n10685), .ZN(
        n10690) );
  AOI22_X1 U11269 ( .A1(n10701), .A2(n10690), .B1(n10688), .B2(n10699), .ZN(
        P2_U3534) );
  INV_X1 U11270 ( .A(P2_REG0_REG_14__SCAN_IN), .ZN(n10689) );
  AOI22_X1 U11271 ( .A1(n10613), .A2(n10690), .B1(n10689), .B2(n10702), .ZN(
        P2_U3493) );
  OAI22_X1 U11272 ( .A1(n10694), .A2(n10693), .B1(n10692), .B2(n10691), .ZN(
        n10695) );
  AOI211_X1 U11273 ( .C1(n10698), .C2(n10697), .A(n10696), .B(n10695), .ZN(
        n10704) );
  INV_X1 U11274 ( .A(P2_REG1_REG_15__SCAN_IN), .ZN(n10700) );
  AOI22_X1 U11275 ( .A1(n10701), .A2(n10704), .B1(n10700), .B2(n10699), .ZN(
        P2_U3535) );
  INV_X1 U11276 ( .A(P2_REG0_REG_15__SCAN_IN), .ZN(n10703) );
  AOI22_X1 U11277 ( .A1(n10613), .A2(n10704), .B1(n10703), .B2(n10702), .ZN(
        P2_U3496) );
  XNOR2_X1 U11278 ( .A(P2_WR_REG_SCAN_IN), .B(P1_WR_REG_SCAN_IN), .ZN(U123) );
  INV_X2 U4922 ( .A(n5548), .ZN(n6419) );
  CLKBUF_X1 U4932 ( .A(n5590), .Z(n6418) );
  INV_X1 U4933 ( .A(n6953), .ZN(n5523) );
  INV_X4 U4942 ( .A(n10693), .ZN(n5299) );
  CLKBUF_X1 U4949 ( .A(n7033), .Z(n8682) );
  OR2_X2 U4989 ( .A1(n5531), .A2(n5530), .ZN(n5548) );
  CLKBUF_X1 U5929 ( .A(n6578), .Z(n4855) );
endmodule

