

module b14_C_lock ( keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, 
        keyinput_5, keyinput_6, keyinput_7, keyinput_8, keyinput_9, 
        keyinput_10, keyinput_11, keyinput_12, keyinput_13, keyinput_14, 
        keyinput_15, keyinput_16, keyinput_17, keyinput_18, keyinput_19, 
        keyinput_20, keyinput_21, keyinput_22, keyinput_23, keyinput_24, 
        keyinput_25, keyinput_26, keyinput_27, keyinput_28, keyinput_29, 
        keyinput_30, keyinput_31, keyinput_32, keyinput_33, keyinput_34, 
        keyinput_35, keyinput_36, keyinput_37, keyinput_38, keyinput_39, 
        keyinput_40, keyinput_41, keyinput_42, keyinput_43, keyinput_44, 
        keyinput_45, keyinput_46, keyinput_47, keyinput_48, keyinput_49, 
        keyinput_50, keyinput_51, keyinput_52, keyinput_53, keyinput_54, 
        keyinput_55, keyinput_56, keyinput_57, keyinput_58, keyinput_59, 
        keyinput_60, keyinput_61, keyinput_62, keyinput_63, keyinput_64, 
        keyinput_65, keyinput_66, keyinput_67, keyinput_68, keyinput_69, 
        keyinput_70, keyinput_71, keyinput_72, keyinput_73, keyinput_74, 
        keyinput_75, keyinput_76, keyinput_77, keyinput_78, keyinput_79, 
        keyinput_80, keyinput_81, keyinput_82, keyinput_83, keyinput_84, 
        keyinput_85, keyinput_86, keyinput_87, keyinput_88, keyinput_89, 
        keyinput_90, keyinput_91, keyinput_92, keyinput_93, keyinput_94, 
        keyinput_95, keyinput_96, keyinput_97, keyinput_98, keyinput_99, 
        keyinput_100, keyinput_101, keyinput_102, keyinput_103, keyinput_104, 
        keyinput_105, keyinput_106, keyinput_107, keyinput_108, keyinput_109, 
        keyinput_110, keyinput_111, keyinput_112, keyinput_113, keyinput_114, 
        keyinput_115, keyinput_116, keyinput_117, keyinput_118, keyinput_119, 
        keyinput_120, keyinput_121, keyinput_122, keyinput_123, keyinput_124, 
        keyinput_125, keyinput_126, keyinput_127, keyinput_128, keyinput_129, 
        keyinput_130, keyinput_131, keyinput_132, keyinput_133, keyinput_134, 
        keyinput_135, keyinput_136, keyinput_137, keyinput_138, keyinput_139, 
        keyinput_140, keyinput_141, keyinput_142, keyinput_143, keyinput_144, 
        keyinput_145, keyinput_146, keyinput_147, keyinput_148, keyinput_149, 
        keyinput_150, keyinput_151, keyinput_152, keyinput_153, keyinput_154, 
        keyinput_155, keyinput_156, keyinput_157, keyinput_158, keyinput_159, 
        keyinput_160, keyinput_161, keyinput_162, keyinput_163, keyinput_164, 
        keyinput_165, keyinput_166, keyinput_167, keyinput_168, keyinput_169, 
        keyinput_170, keyinput_171, keyinput_172, keyinput_173, keyinput_174, 
        keyinput_175, keyinput_176, keyinput_177, keyinput_178, keyinput_179, 
        keyinput_180, keyinput_181, keyinput_182, keyinput_183, keyinput_184, 
        keyinput_185, keyinput_186, keyinput_187, keyinput_188, keyinput_189, 
        keyinput_190, keyinput_191, keyinput_192, keyinput_193, keyinput_194, 
        keyinput_195, keyinput_196, keyinput_197, keyinput_198, keyinput_199, 
        keyinput_200, keyinput_201, keyinput_202, keyinput_203, keyinput_204, 
        keyinput_205, keyinput_206, keyinput_207, keyinput_208, keyinput_209, 
        keyinput_210, keyinput_211, keyinput_212, keyinput_213, keyinput_214, 
        keyinput_215, keyinput_216, keyinput_217, keyinput_218, keyinput_219, 
        keyinput_220, keyinput_221, keyinput_222, keyinput_223, keyinput_224, 
        keyinput_225, keyinput_226, keyinput_227, keyinput_228, keyinput_229, 
        keyinput_230, keyinput_231, keyinput_232, keyinput_233, keyinput_234, 
        keyinput_235, keyinput_236, keyinput_237, keyinput_238, keyinput_239, 
        keyinput_240, keyinput_241, keyinput_242, keyinput_243, keyinput_244, 
        keyinput_245, keyinput_246, keyinput_247, keyinput_248, keyinput_249, 
        keyinput_250, keyinput_251, keyinput_252, keyinput_253, keyinput_254, 
        keyinput_255, DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, 
        DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, 
        DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, 
        DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, 
        DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, 
        DATAI_1_, DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN, 
        REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN, 
        REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN, 
        REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN, 
        REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN, 
        REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN, 
        REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN, 
        REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN, 
        IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN, 
        IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN, 
        IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN, 
        IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN, 
        IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN, 
        IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN, 
        IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN, 
        IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN, 
        IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN, 
        IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN, 
        IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN, 
        D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN, D_REG_4__SCAN_IN, 
        D_REG_5__SCAN_IN, D_REG_6__SCAN_IN, D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, 
        D_REG_9__SCAN_IN, D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, 
        D_REG_12__SCAN_IN, D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, 
        D_REG_15__SCAN_IN, D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, 
        D_REG_18__SCAN_IN, D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, 
        D_REG_21__SCAN_IN, D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, 
        D_REG_24__SCAN_IN, D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, 
        D_REG_27__SCAN_IN, D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, 
        D_REG_30__SCAN_IN, D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, 
        REG0_REG_1__SCAN_IN, REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, 
        REG0_REG_4__SCAN_IN, REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, 
        REG0_REG_7__SCAN_IN, REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, 
        REG0_REG_10__SCAN_IN, REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, 
        REG0_REG_13__SCAN_IN, REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, 
        REG0_REG_16__SCAN_IN, REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, 
        REG0_REG_19__SCAN_IN, REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, 
        REG0_REG_22__SCAN_IN, REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, 
        REG0_REG_25__SCAN_IN, REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, 
        REG0_REG_28__SCAN_IN, REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, 
        REG0_REG_31__SCAN_IN, REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, 
        REG1_REG_2__SCAN_IN, REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, 
        REG1_REG_5__SCAN_IN, REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, 
        REG1_REG_8__SCAN_IN, REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, 
        REG1_REG_11__SCAN_IN, REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, 
        REG1_REG_14__SCAN_IN, REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, 
        REG1_REG_17__SCAN_IN, REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, 
        REG1_REG_20__SCAN_IN, REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, 
        REG1_REG_23__SCAN_IN, REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, 
        REG1_REG_26__SCAN_IN, REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, 
        REG1_REG_29__SCAN_IN, REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, 
        REG2_REG_0__SCAN_IN, REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, 
        REG2_REG_3__SCAN_IN, REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, 
        REG2_REG_6__SCAN_IN, REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, 
        REG2_REG_9__SCAN_IN, REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, 
        REG2_REG_12__SCAN_IN, REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, 
        REG2_REG_15__SCAN_IN, REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, 
        REG2_REG_18__SCAN_IN, REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, 
        REG2_REG_21__SCAN_IN, REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, 
        REG2_REG_24__SCAN_IN, REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, 
        REG2_REG_27__SCAN_IN, REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, 
        REG2_REG_30__SCAN_IN, REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, 
        ADDR_REG_18__SCAN_IN, ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, 
        ADDR_REG_15__SCAN_IN, ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, 
        ADDR_REG_12__SCAN_IN, ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, 
        ADDR_REG_9__SCAN_IN, ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, 
        ADDR_REG_6__SCAN_IN, ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, 
        ADDR_REG_3__SCAN_IN, ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, 
        ADDR_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        B_REG_SCAN_IN, REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, 
        REG3_REG_6__SCAN_IN, REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, 
        REG3_REG_11__SCAN_IN, REG3_REG_22__SCAN_IN, U3352, U3351, U3350, U3349, 
        U3348, U3347, U3346, U3345, U3344, U3343, U3342, U3341, U3340, U3339, 
        U3338, U3337, U3336, U3335, U3334, U3333, U3332, U3331, U3330, U3329, 
        U3328, U3327, U3326, U3325, U3324, U3323, U3322, U3321, U3458, U3459, 
        U3320, U3319, U3318, U3317, U3316, U3315, U3314, U3313, U3312, U3311, 
        U3310, U3309, U3308, U3307, U3306, U3305, U3304, U3303, U3302, U3301, 
        U3300, U3299, U3298, U3297, U3296, U3295, U3294, U3293, U3292, U3291, 
        U3467, U3469, U3471, U3473, U3475, U3477, U3479, U3481, U3483, U3485, 
        U3487, U3489, U3491, U3493, U3495, U3497, U3499, U3501, U3503, U3505, 
        U3506, U3507, U3508, U3509, U3510, U3511, U3512, U3513, U3514, U3515, 
        U3516, U3517, U3518, U3519, U3520, U3521, U3522, U3523, U3524, U3525, 
        U3526, U3527, U3528, U3529, U3530, U3531, U3532, U3533, U3534, U3535, 
        U3536, U3537, U3538, U3539, U3540, U3541, U3542, U3543, U3544, U3545, 
        U3546, U3547, U3548, U3549, U3290, U3289, U3288, U3287, U3286, U3285, 
        U3284, U3283, U3282, U3281, U3280, U3279, U3278, U3277, U3276, U3275, 
        U3274, U3273, U3272, U3271, U3270, U3269, U3268, U3267, U3266, U3265, 
        U3264, U3263, U3262, U3354, U3261, U3260, U3259, U3258, U3257, U3256, 
        U3255, U3254, U3253, U3252, U3251, U3250, U3249, U3248, U3247, U3246, 
        U3245, U3244, U3243, U3242, U3241, U3240, U3550, U3551, U3552, U3553, 
        U3554, U3555, U3556, U3557, U3558, U3559, U3560, U3561, U3562, U3563, 
        U3564, U3565, U3566, U3567, U3568, U3569, U3570, U3571, U3572, U3573, 
        U3574, U3575, U3576, U3577, U3578, U3579, U3580, U3581, U3239, U3238, 
        U3237, U3236, U3235, U3234, U3233, U3232, U3231, U3230, U3229, U3228, 
        U3227, U3226, U3225, U3224, U3223, U3222, U3221, U3220, U3219, U3218, 
        U3217, U3216, U3215, U3214, U3213, U3212, U3211, U3210, U3149, U3148, 
        U4043 );
  input keyinput_0, keyinput_1, keyinput_2, keyinput_3, keyinput_4, keyinput_5,
         keyinput_6, keyinput_7, keyinput_8, keyinput_9, keyinput_10,
         keyinput_11, keyinput_12, keyinput_13, keyinput_14, keyinput_15,
         keyinput_16, keyinput_17, keyinput_18, keyinput_19, keyinput_20,
         keyinput_21, keyinput_22, keyinput_23, keyinput_24, keyinput_25,
         keyinput_26, keyinput_27, keyinput_28, keyinput_29, keyinput_30,
         keyinput_31, keyinput_32, keyinput_33, keyinput_34, keyinput_35,
         keyinput_36, keyinput_37, keyinput_38, keyinput_39, keyinput_40,
         keyinput_41, keyinput_42, keyinput_43, keyinput_44, keyinput_45,
         keyinput_46, keyinput_47, keyinput_48, keyinput_49, keyinput_50,
         keyinput_51, keyinput_52, keyinput_53, keyinput_54, keyinput_55,
         keyinput_56, keyinput_57, keyinput_58, keyinput_59, keyinput_60,
         keyinput_61, keyinput_62, keyinput_63, keyinput_64, keyinput_65,
         keyinput_66, keyinput_67, keyinput_68, keyinput_69, keyinput_70,
         keyinput_71, keyinput_72, keyinput_73, keyinput_74, keyinput_75,
         keyinput_76, keyinput_77, keyinput_78, keyinput_79, keyinput_80,
         keyinput_81, keyinput_82, keyinput_83, keyinput_84, keyinput_85,
         keyinput_86, keyinput_87, keyinput_88, keyinput_89, keyinput_90,
         keyinput_91, keyinput_92, keyinput_93, keyinput_94, keyinput_95,
         keyinput_96, keyinput_97, keyinput_98, keyinput_99, keyinput_100,
         keyinput_101, keyinput_102, keyinput_103, keyinput_104, keyinput_105,
         keyinput_106, keyinput_107, keyinput_108, keyinput_109, keyinput_110,
         keyinput_111, keyinput_112, keyinput_113, keyinput_114, keyinput_115,
         keyinput_116, keyinput_117, keyinput_118, keyinput_119, keyinput_120,
         keyinput_121, keyinput_122, keyinput_123, keyinput_124, keyinput_125,
         keyinput_126, keyinput_127, keyinput_128, keyinput_129, keyinput_130,
         keyinput_131, keyinput_132, keyinput_133, keyinput_134, keyinput_135,
         keyinput_136, keyinput_137, keyinput_138, keyinput_139, keyinput_140,
         keyinput_141, keyinput_142, keyinput_143, keyinput_144, keyinput_145,
         keyinput_146, keyinput_147, keyinput_148, keyinput_149, keyinput_150,
         keyinput_151, keyinput_152, keyinput_153, keyinput_154, keyinput_155,
         keyinput_156, keyinput_157, keyinput_158, keyinput_159, keyinput_160,
         keyinput_161, keyinput_162, keyinput_163, keyinput_164, keyinput_165,
         keyinput_166, keyinput_167, keyinput_168, keyinput_169, keyinput_170,
         keyinput_171, keyinput_172, keyinput_173, keyinput_174, keyinput_175,
         keyinput_176, keyinput_177, keyinput_178, keyinput_179, keyinput_180,
         keyinput_181, keyinput_182, keyinput_183, keyinput_184, keyinput_185,
         keyinput_186, keyinput_187, keyinput_188, keyinput_189, keyinput_190,
         keyinput_191, keyinput_192, keyinput_193, keyinput_194, keyinput_195,
         keyinput_196, keyinput_197, keyinput_198, keyinput_199, keyinput_200,
         keyinput_201, keyinput_202, keyinput_203, keyinput_204, keyinput_205,
         keyinput_206, keyinput_207, keyinput_208, keyinput_209, keyinput_210,
         keyinput_211, keyinput_212, keyinput_213, keyinput_214, keyinput_215,
         keyinput_216, keyinput_217, keyinput_218, keyinput_219, keyinput_220,
         keyinput_221, keyinput_222, keyinput_223, keyinput_224, keyinput_225,
         keyinput_226, keyinput_227, keyinput_228, keyinput_229, keyinput_230,
         keyinput_231, keyinput_232, keyinput_233, keyinput_234, keyinput_235,
         keyinput_236, keyinput_237, keyinput_238, keyinput_239, keyinput_240,
         keyinput_241, keyinput_242, keyinput_243, keyinput_244, keyinput_245,
         keyinput_246, keyinput_247, keyinput_248, keyinput_249, keyinput_250,
         keyinput_251, keyinput_252, keyinput_253, keyinput_254, keyinput_255,
         DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, STATE_REG_SCAN_IN, REG3_REG_7__SCAN_IN,
         REG3_REG_27__SCAN_IN, REG3_REG_14__SCAN_IN, REG3_REG_23__SCAN_IN,
         REG3_REG_10__SCAN_IN, REG3_REG_3__SCAN_IN, REG3_REG_19__SCAN_IN,
         REG3_REG_28__SCAN_IN, REG3_REG_8__SCAN_IN, REG3_REG_1__SCAN_IN,
         REG3_REG_21__SCAN_IN, REG3_REG_12__SCAN_IN, REG3_REG_25__SCAN_IN,
         REG3_REG_16__SCAN_IN, REG3_REG_5__SCAN_IN, REG3_REG_17__SCAN_IN,
         REG3_REG_24__SCAN_IN, REG3_REG_4__SCAN_IN, REG3_REG_9__SCAN_IN,
         REG3_REG_0__SCAN_IN, REG3_REG_20__SCAN_IN, REG3_REG_13__SCAN_IN,
         IR_REG_0__SCAN_IN, IR_REG_1__SCAN_IN, IR_REG_2__SCAN_IN,
         IR_REG_3__SCAN_IN, IR_REG_4__SCAN_IN, IR_REG_5__SCAN_IN,
         IR_REG_6__SCAN_IN, IR_REG_7__SCAN_IN, IR_REG_8__SCAN_IN,
         IR_REG_9__SCAN_IN, IR_REG_10__SCAN_IN, IR_REG_11__SCAN_IN,
         IR_REG_12__SCAN_IN, IR_REG_13__SCAN_IN, IR_REG_14__SCAN_IN,
         IR_REG_15__SCAN_IN, IR_REG_16__SCAN_IN, IR_REG_17__SCAN_IN,
         IR_REG_18__SCAN_IN, IR_REG_19__SCAN_IN, IR_REG_20__SCAN_IN,
         IR_REG_21__SCAN_IN, IR_REG_22__SCAN_IN, IR_REG_23__SCAN_IN,
         IR_REG_24__SCAN_IN, IR_REG_25__SCAN_IN, IR_REG_26__SCAN_IN,
         IR_REG_27__SCAN_IN, IR_REG_28__SCAN_IN, IR_REG_29__SCAN_IN,
         IR_REG_30__SCAN_IN, IR_REG_31__SCAN_IN, D_REG_0__SCAN_IN,
         D_REG_1__SCAN_IN, D_REG_2__SCAN_IN, D_REG_3__SCAN_IN,
         D_REG_4__SCAN_IN, D_REG_5__SCAN_IN, D_REG_6__SCAN_IN,
         D_REG_7__SCAN_IN, D_REG_8__SCAN_IN, D_REG_9__SCAN_IN,
         D_REG_10__SCAN_IN, D_REG_11__SCAN_IN, D_REG_12__SCAN_IN,
         D_REG_13__SCAN_IN, D_REG_14__SCAN_IN, D_REG_15__SCAN_IN,
         D_REG_16__SCAN_IN, D_REG_17__SCAN_IN, D_REG_18__SCAN_IN,
         D_REG_19__SCAN_IN, D_REG_20__SCAN_IN, D_REG_21__SCAN_IN,
         D_REG_22__SCAN_IN, D_REG_23__SCAN_IN, D_REG_24__SCAN_IN,
         D_REG_25__SCAN_IN, D_REG_26__SCAN_IN, D_REG_27__SCAN_IN,
         D_REG_28__SCAN_IN, D_REG_29__SCAN_IN, D_REG_30__SCAN_IN,
         D_REG_31__SCAN_IN, REG0_REG_0__SCAN_IN, REG0_REG_1__SCAN_IN,
         REG0_REG_2__SCAN_IN, REG0_REG_3__SCAN_IN, REG0_REG_4__SCAN_IN,
         REG0_REG_5__SCAN_IN, REG0_REG_6__SCAN_IN, REG0_REG_7__SCAN_IN,
         REG0_REG_8__SCAN_IN, REG0_REG_9__SCAN_IN, REG0_REG_10__SCAN_IN,
         REG0_REG_11__SCAN_IN, REG0_REG_12__SCAN_IN, REG0_REG_13__SCAN_IN,
         REG0_REG_14__SCAN_IN, REG0_REG_15__SCAN_IN, REG0_REG_16__SCAN_IN,
         REG0_REG_17__SCAN_IN, REG0_REG_18__SCAN_IN, REG0_REG_19__SCAN_IN,
         REG0_REG_20__SCAN_IN, REG0_REG_21__SCAN_IN, REG0_REG_22__SCAN_IN,
         REG0_REG_23__SCAN_IN, REG0_REG_24__SCAN_IN, REG0_REG_25__SCAN_IN,
         REG0_REG_26__SCAN_IN, REG0_REG_27__SCAN_IN, REG0_REG_28__SCAN_IN,
         REG0_REG_29__SCAN_IN, REG0_REG_30__SCAN_IN, REG0_REG_31__SCAN_IN,
         REG1_REG_0__SCAN_IN, REG1_REG_1__SCAN_IN, REG1_REG_2__SCAN_IN,
         REG1_REG_3__SCAN_IN, REG1_REG_4__SCAN_IN, REG1_REG_5__SCAN_IN,
         REG1_REG_6__SCAN_IN, REG1_REG_7__SCAN_IN, REG1_REG_8__SCAN_IN,
         REG1_REG_9__SCAN_IN, REG1_REG_10__SCAN_IN, REG1_REG_11__SCAN_IN,
         REG1_REG_12__SCAN_IN, REG1_REG_13__SCAN_IN, REG1_REG_14__SCAN_IN,
         REG1_REG_15__SCAN_IN, REG1_REG_16__SCAN_IN, REG1_REG_17__SCAN_IN,
         REG1_REG_18__SCAN_IN, REG1_REG_19__SCAN_IN, REG1_REG_20__SCAN_IN,
         REG1_REG_21__SCAN_IN, REG1_REG_22__SCAN_IN, REG1_REG_23__SCAN_IN,
         REG1_REG_24__SCAN_IN, REG1_REG_25__SCAN_IN, REG1_REG_26__SCAN_IN,
         REG1_REG_27__SCAN_IN, REG1_REG_28__SCAN_IN, REG1_REG_29__SCAN_IN,
         REG1_REG_30__SCAN_IN, REG1_REG_31__SCAN_IN, REG2_REG_0__SCAN_IN,
         REG2_REG_1__SCAN_IN, REG2_REG_2__SCAN_IN, REG2_REG_3__SCAN_IN,
         REG2_REG_4__SCAN_IN, REG2_REG_5__SCAN_IN, REG2_REG_6__SCAN_IN,
         REG2_REG_7__SCAN_IN, REG2_REG_8__SCAN_IN, REG2_REG_9__SCAN_IN,
         REG2_REG_10__SCAN_IN, REG2_REG_11__SCAN_IN, REG2_REG_12__SCAN_IN,
         REG2_REG_13__SCAN_IN, REG2_REG_14__SCAN_IN, REG2_REG_15__SCAN_IN,
         REG2_REG_16__SCAN_IN, REG2_REG_17__SCAN_IN, REG2_REG_18__SCAN_IN,
         REG2_REG_19__SCAN_IN, REG2_REG_20__SCAN_IN, REG2_REG_21__SCAN_IN,
         REG2_REG_22__SCAN_IN, REG2_REG_23__SCAN_IN, REG2_REG_24__SCAN_IN,
         REG2_REG_25__SCAN_IN, REG2_REG_26__SCAN_IN, REG2_REG_27__SCAN_IN,
         REG2_REG_28__SCAN_IN, REG2_REG_29__SCAN_IN, REG2_REG_30__SCAN_IN,
         REG2_REG_31__SCAN_IN, ADDR_REG_19__SCAN_IN, ADDR_REG_18__SCAN_IN,
         ADDR_REG_17__SCAN_IN, ADDR_REG_16__SCAN_IN, ADDR_REG_15__SCAN_IN,
         ADDR_REG_14__SCAN_IN, ADDR_REG_13__SCAN_IN, ADDR_REG_12__SCAN_IN,
         ADDR_REG_11__SCAN_IN, ADDR_REG_10__SCAN_IN, ADDR_REG_9__SCAN_IN,
         ADDR_REG_8__SCAN_IN, ADDR_REG_7__SCAN_IN, ADDR_REG_6__SCAN_IN,
         ADDR_REG_5__SCAN_IN, ADDR_REG_4__SCAN_IN, ADDR_REG_3__SCAN_IN,
         ADDR_REG_2__SCAN_IN, ADDR_REG_1__SCAN_IN, ADDR_REG_0__SCAN_IN,
         DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, DATAO_REG_2__SCAN_IN,
         DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, DATAO_REG_5__SCAN_IN,
         DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, DATAO_REG_8__SCAN_IN,
         DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, DATAO_REG_11__SCAN_IN,
         DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, DATAO_REG_14__SCAN_IN,
         DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, DATAO_REG_17__SCAN_IN,
         DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, DATAO_REG_20__SCAN_IN,
         DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, DATAO_REG_23__SCAN_IN,
         DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, DATAO_REG_26__SCAN_IN,
         DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, DATAO_REG_29__SCAN_IN,
         DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, B_REG_SCAN_IN,
         REG3_REG_15__SCAN_IN, REG3_REG_26__SCAN_IN, REG3_REG_6__SCAN_IN,
         REG3_REG_18__SCAN_IN, REG3_REG_2__SCAN_IN, REG3_REG_11__SCAN_IN,
         REG3_REG_22__SCAN_IN;
  output U3352, U3351, U3350, U3349, U3348, U3347, U3346, U3345, U3344, U3343,
         U3342, U3341, U3340, U3339, U3338, U3337, U3336, U3335, U3334, U3333,
         U3332, U3331, U3330, U3329, U3328, U3327, U3326, U3325, U3324, U3323,
         U3322, U3321, U3458, U3459, U3320, U3319, U3318, U3317, U3316, U3315,
         U3314, U3313, U3312, U3311, U3310, U3309, U3308, U3307, U3306, U3305,
         U3304, U3303, U3302, U3301, U3300, U3299, U3298, U3297, U3296, U3295,
         U3294, U3293, U3292, U3291, U3467, U3469, U3471, U3473, U3475, U3477,
         U3479, U3481, U3483, U3485, U3487, U3489, U3491, U3493, U3495, U3497,
         U3499, U3501, U3503, U3505, U3506, U3507, U3508, U3509, U3510, U3511,
         U3512, U3513, U3514, U3515, U3516, U3517, U3518, U3519, U3520, U3521,
         U3522, U3523, U3524, U3525, U3526, U3527, U3528, U3529, U3530, U3531,
         U3532, U3533, U3534, U3535, U3536, U3537, U3538, U3539, U3540, U3541,
         U3542, U3543, U3544, U3545, U3546, U3547, U3548, U3549, U3290, U3289,
         U3288, U3287, U3286, U3285, U3284, U3283, U3282, U3281, U3280, U3279,
         U3278, U3277, U3276, U3275, U3274, U3273, U3272, U3271, U3270, U3269,
         U3268, U3267, U3266, U3265, U3264, U3263, U3262, U3354, U3261, U3260,
         U3259, U3258, U3257, U3256, U3255, U3254, U3253, U3252, U3251, U3250,
         U3249, U3248, U3247, U3246, U3245, U3244, U3243, U3242, U3241, U3240,
         U3550, U3551, U3552, U3553, U3554, U3555, U3556, U3557, U3558, U3559,
         U3560, U3561, U3562, U3563, U3564, U3565, U3566, U3567, U3568, U3569,
         U3570, U3571, U3572, U3573, U3574, U3575, U3576, U3577, U3578, U3579,
         U3580, U3581, U3239, U3238, U3237, U3236, U3235, U3234, U3233, U3232,
         U3231, U3230, U3229, U3228, U3227, U3226, U3225, U3224, U3223, U3222,
         U3221, U3220, U3219, U3218, U3217, U3216, U3215, U3214, U3213, U3212,
         U3211, U3210, U3149, U3148, U4043;
  wire   n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341;

  INV_X1 U2530 ( .A(n4591), .ZN(n3508) );
  INV_X1 U2531 ( .A(n3251), .ZN(n3237) );
  NAND2_X1 U2532 ( .A1(n2818), .A2(n3284), .ZN(n3464) );
  INV_X4 U2533 ( .A(n3254), .ZN(n2875) );
  NAND2_X1 U2534 ( .A1(n3286), .A2(n5041), .ZN(n2818) );
  INV_X1 U2535 ( .A(IR_REG_31__SCAN_IN), .ZN(n3093) );
  INV_X1 U2536 ( .A(n2978), .ZN(n2495) );
  AND2_X2 U2537 ( .A1(n4954), .A2(n4953), .ZN(n4955) );
  NAND2_X2 U2538 ( .A1(n2815), .A2(n2777), .ZN(n2798) );
  INV_X2 U2539 ( .A(n2814), .ZN(n2815) );
  XNOR2_X2 U2540 ( .A(n4743), .B(n4742), .ZN(n4981) );
  INV_X1 U2541 ( .A(n3493), .ZN(n3507) );
  NAND2_X2 U2543 ( .A1(n3285), .A2(n4710), .ZN(n2872) );
  NOR2_X1 U2544 ( .A1(IR_REG_1__SCAN_IN), .A2(IR_REG_0__SCAN_IN), .ZN(n2826)
         );
  AND2_X1 U2545 ( .A1(n4979), .A2(n2641), .ZN(n2640) );
  OR2_X1 U2546 ( .A1(n4269), .A2(n4270), .ZN(n4271) );
  OR2_X1 U2547 ( .A1(n4699), .A2(n2610), .ZN(n2607) );
  AOI21_X1 U2548 ( .B1(n4876), .B2(n4240), .A(n4544), .ZN(n4860) );
  OAI21_X1 U2549 ( .B1(n4948), .B2(n2637), .A(n2526), .ZN(n4876) );
  NAND2_X1 U2550 ( .A1(n4234), .A2(n4443), .ZN(n4948) );
  OR2_X1 U2551 ( .A1(n4194), .A2(n4202), .ZN(n4234) );
  OR2_X1 U2552 ( .A1(n4615), .A2(n2728), .ZN(n4616) );
  NOR2_X1 U2553 ( .A1(n4828), .A2(n4827), .ZN(n4830) );
  OR2_X1 U2554 ( .A1(n2500), .A2(n4273), .ZN(n4828) );
  AOI21_X1 U2555 ( .B1(n3586), .B2(n4436), .A(n4439), .ZN(n3639) );
  OAI211_X1 U2556 ( .C1(n5185), .C2(n2632), .A(n2629), .B(n4451), .ZN(n3574)
         );
  OR2_X1 U2557 ( .A1(n3452), .A2(n3453), .ZN(n4361) );
  NAND2_X2 U2558 ( .A1(n3290), .A2(n5210), .ZN(n5276) );
  AND2_X1 U2559 ( .A1(n4433), .A2(n4451), .ZN(n4537) );
  INV_X1 U2560 ( .A(n5187), .ZN(n4590) );
  NAND2_X1 U2561 ( .A1(n2724), .A2(n2723), .ZN(n3366) );
  NAND4_X2 U2562 ( .A1(n2825), .A2(n2824), .A3(n2823), .A4(n2822), .ZN(n5156)
         );
  AND4_X1 U2563 ( .A1(n2852), .A2(n2851), .A3(n2850), .A4(n2849), .ZN(n5187)
         );
  NAND4_X1 U2564 ( .A1(n2871), .A2(n2870), .A3(n2869), .A4(n2868), .ZN(n4593)
         );
  OR2_X2 U2565 ( .A1(n2830), .A2(n3477), .ZN(n3251) );
  NAND2_X1 U2566 ( .A1(n2649), .A2(n2648), .ZN(n4304) );
  NAND2_X2 U2567 ( .A1(n2878), .A2(n5169), .ZN(n3254) );
  INV_X2 U2568 ( .A(n2495), .ZN(n2496) );
  CLKBUF_X3 U2569 ( .A(n2867), .Z(n3293) );
  MUX2_X1 U2570 ( .A(n5057), .B(DATAI_2_), .S(n2872), .Z(n3493) );
  NAND2_X1 U2571 ( .A1(n4567), .A2(n3288), .ZN(n5319) );
  BUF_X2 U2572 ( .A(n2872), .Z(n4491) );
  NAND2_X1 U2573 ( .A1(n3392), .A2(n3363), .ZN(n3364) );
  NAND2_X1 U2574 ( .A1(n2819), .A2(IR_REG_31__SCAN_IN), .ZN(n2820) );
  XNOR2_X1 U2575 ( .A(n2821), .B(n4016), .ZN(n4710) );
  OR2_X1 U2576 ( .A1(n2782), .A2(n3093), .ZN(n2781) );
  NAND2_X1 U2577 ( .A1(n2688), .A2(IR_REG_31__SCAN_IN), .ZN(n2821) );
  OR2_X1 U2578 ( .A1(n2762), .A2(n2779), .ZN(n2503) );
  AND4_X1 U2579 ( .A1(n2826), .A2(n2771), .A3(n2773), .A4(n2770), .ZN(n2606)
         );
  INV_X1 U2580 ( .A(IR_REG_21__SCAN_IN), .ZN(n3808) );
  NOR2_X1 U2581 ( .A1(IR_REG_16__SCAN_IN), .A2(IR_REG_15__SCAN_IN), .ZN(n2803)
         );
  INV_X1 U2582 ( .A(IR_REG_24__SCAN_IN), .ZN(n4011) );
  INV_X1 U2583 ( .A(IR_REG_4__SCAN_IN), .ZN(n3980) );
  NOR2_X1 U2584 ( .A1(IR_REG_3__SCAN_IN), .A2(IR_REG_2__SCAN_IN), .ZN(n2769)
         );
  NOR2_X1 U2585 ( .A1(IR_REG_10__SCAN_IN), .A2(IR_REG_12__SCAN_IN), .ZN(n2770)
         );
  NOR2_X1 U2586 ( .A1(IR_REG_28__SCAN_IN), .A2(IR_REG_27__SCAN_IN), .ZN(n2780)
         );
  NOR2_X1 U2587 ( .A1(IR_REG_11__SCAN_IN), .A2(IR_REG_8__SCAN_IN), .ZN(n2773)
         );
  NOR2_X1 U2588 ( .A1(IR_REG_7__SCAN_IN), .A2(IR_REG_5__SCAN_IN), .ZN(n2771)
         );
  INV_X2 U2589 ( .A(n2495), .ZN(n2497) );
  AND2_X4 U2590 ( .A1(n5035), .A2(n5036), .ZN(n2866) );
  AND2_X1 U2591 ( .A1(n2785), .A2(n2786), .ZN(n2978) );
  AND2_X4 U2592 ( .A1(n2785), .A2(n5036), .ZN(n2865) );
  XNOR2_X2 U2593 ( .A(n2781), .B(n3827), .ZN(n2785) );
  INV_X1 U2594 ( .A(n4787), .ZN(n4745) );
  INV_X1 U2595 ( .A(n4535), .ZN(n2671) );
  NAND2_X1 U2596 ( .A1(n4936), .A2(n4227), .ZN(n4228) );
  INV_X1 U2597 ( .A(n3383), .ZN(n2713) );
  NAND2_X1 U2598 ( .A1(n2616), .A2(n2615), .ZN(n2614) );
  INV_X1 U2599 ( .A(n4698), .ZN(n2615) );
  INV_X1 U2600 ( .A(n4700), .ZN(n2616) );
  AND2_X1 U2601 ( .A1(n2741), .A2(n2568), .ZN(n2567) );
  AOI21_X1 U2602 ( .B1(n2742), .B2(n2744), .A(n2525), .ZN(n2741) );
  NAND2_X1 U2603 ( .A1(n2742), .A2(n2569), .ZN(n2568) );
  AOI21_X1 U2604 ( .B1(n2652), .B2(n2654), .A(n2523), .ZN(n2650) );
  NAND2_X1 U2605 ( .A1(n4421), .A2(n3483), .ZN(n3458) );
  AND2_X1 U2606 ( .A1(n4900), .A2(n4229), .ZN(n2655) );
  NOR2_X1 U2607 ( .A1(n2605), .A2(IR_REG_22__SCAN_IN), .ZN(n2602) );
  INV_X1 U2608 ( .A(n2751), .ZN(n2603) );
  NAND2_X1 U2609 ( .A1(n5057), .A2(REG2_REG_2__SCAN_IN), .ZN(n2689) );
  NAND2_X1 U2610 ( .A1(n5098), .A2(n3365), .ZN(n2726) );
  NAND2_X1 U2611 ( .A1(n2726), .A2(n2725), .ZN(n2724) );
  INV_X1 U2612 ( .A(n3379), .ZN(n2725) );
  NAND2_X1 U2613 ( .A1(n3537), .A2(n3538), .ZN(n3541) );
  AND2_X1 U2614 ( .A1(n5051), .A2(REG2_REG_9__SCAN_IN), .ZN(n3616) );
  OR2_X1 U2615 ( .A1(n4603), .A2(n4604), .ZN(n2566) );
  NAND2_X1 U2616 ( .A1(n2566), .A2(n2565), .ZN(n4620) );
  INV_X1 U2617 ( .A(n4608), .ZN(n2565) );
  NAND2_X1 U2618 ( .A1(n4680), .A2(n4681), .ZN(n4690) );
  NAND2_X1 U2619 ( .A1(n2561), .A2(n2560), .ZN(n2692) );
  INV_X1 U2620 ( .A(n4675), .ZN(n2560) );
  AOI21_X1 U2621 ( .B1(n4764), .B2(n2665), .A(n2532), .ZN(n2664) );
  INV_X1 U2622 ( .A(n4728), .ZN(n2665) );
  NOR2_X1 U2623 ( .A1(n4530), .A2(n4702), .ZN(n4783) );
  NAND2_X1 U2624 ( .A1(n4957), .A2(n4929), .ZN(n2683) );
  NOR2_X1 U2625 ( .A1(n4960), .A2(n2682), .ZN(n2681) );
  INV_X1 U2626 ( .A(n4225), .ZN(n2682) );
  NAND2_X1 U2627 ( .A1(n2668), .A2(n2667), .ZN(n4121) );
  NAND2_X1 U2628 ( .A1(n2670), .A2(n2679), .ZN(n2667) );
  INV_X1 U2629 ( .A(IR_REG_28__SCAN_IN), .ZN(n4021) );
  INV_X1 U2630 ( .A(IR_REG_27__SCAN_IN), .ZN(n4016) );
  NAND2_X1 U2631 ( .A1(n2810), .A2(n2812), .ZN(n2811) );
  NOR2_X1 U2632 ( .A1(n2905), .A2(IR_REG_5__SCAN_IN), .ZN(n2937) );
  AOI21_X1 U2633 ( .B1(n3627), .B2(n3628), .A(n2977), .ZN(n4281) );
  OR2_X1 U2634 ( .A1(n4673), .A2(n2693), .ZN(n2561) );
  AND2_X1 U2635 ( .A1(n5043), .A2(REG2_REG_17__SCAN_IN), .ZN(n2693) );
  OR2_X1 U2636 ( .A1(n5093), .A2(n2505), .ZN(n2711) );
  AOI21_X1 U2637 ( .B1(n3354), .B2(n2713), .A(n2514), .ZN(n2712) );
  INV_X1 U2638 ( .A(n4703), .ZN(n2617) );
  NAND2_X1 U2639 ( .A1(n2612), .A2(n2614), .ZN(n2611) );
  NAND2_X1 U2640 ( .A1(n4898), .A2(n4867), .ZN(n2596) );
  INV_X1 U2641 ( .A(n4469), .ZN(n2638) );
  NOR2_X1 U2642 ( .A1(n2636), .A2(n4960), .ZN(n2635) );
  INV_X1 U2643 ( .A(n2639), .ZN(n2636) );
  NOR2_X1 U2644 ( .A1(n4470), .A2(n4471), .ZN(n2639) );
  INV_X1 U2645 ( .A(n2626), .ZN(n2625) );
  OAI21_X1 U2646 ( .B1(n4535), .B2(n2627), .A(n4461), .ZN(n2626) );
  NAND2_X1 U2647 ( .A1(n4101), .A2(n4102), .ZN(n2679) );
  NOR2_X1 U2648 ( .A1(n2979), .A2(n3746), .ZN(n2996) );
  AND2_X1 U2649 ( .A1(n2630), .A2(n4537), .ZN(n2628) );
  INV_X1 U2650 ( .A(n4430), .ZN(n2630) );
  AND2_X1 U2651 ( .A1(n5040), .A2(n5041), .ZN(n3465) );
  NAND2_X1 U2652 ( .A1(n4223), .A2(n4222), .ZN(n4225) );
  INV_X1 U2653 ( .A(n5192), .ZN(n5180) );
  NAND2_X1 U2654 ( .A1(n2659), .A2(n3487), .ZN(n2657) );
  AND2_X1 U2655 ( .A1(n3470), .A2(n2817), .ZN(n3288) );
  NAND2_X1 U2656 ( .A1(n2780), .A2(n2793), .ZN(n2762) );
  NOR2_X1 U2657 ( .A1(n2798), .A2(n2503), .ZN(n2601) );
  AND4_X1 U2658 ( .A1(n2803), .A2(n2775), .A3(n2774), .A4(n3996), .ZN(n2776)
         );
  NOR2_X1 U2659 ( .A1(IR_REG_20__SCAN_IN), .A2(IR_REG_19__SCAN_IN), .ZN(n2775)
         );
  NOR2_X1 U2660 ( .A1(IR_REG_18__SCAN_IN), .A2(IR_REG_17__SCAN_IN), .ZN(n2774)
         );
  NAND2_X1 U2661 ( .A1(n2776), .A2(n2753), .ZN(n2751) );
  AND2_X1 U2662 ( .A1(n2754), .A2(n3808), .ZN(n2753) );
  NOR2_X1 U2663 ( .A1(n2804), .A2(IR_REG_14__SCAN_IN), .ZN(n2587) );
  AND2_X1 U2664 ( .A1(n3241), .A2(n3240), .ZN(n3282) );
  AOI21_X1 U2665 ( .B1(n2578), .B2(n2580), .A(n2577), .ZN(n2576) );
  INV_X1 U2666 ( .A(n4372), .ZN(n2577) );
  INV_X1 U2667 ( .A(n3213), .ZN(n4321) );
  NAND2_X1 U2668 ( .A1(n4330), .A2(n4331), .ZN(n2757) );
  NAND2_X1 U2669 ( .A1(n2760), .A2(n2759), .ZN(n2758) );
  INV_X1 U2670 ( .A(n4331), .ZN(n2759) );
  INV_X1 U2671 ( .A(n4330), .ZN(n2760) );
  NAND2_X1 U2672 ( .A1(n4350), .A2(n4351), .ZN(n2740) );
  INV_X1 U2673 ( .A(n3286), .ZN(n4567) );
  NAND2_X1 U2674 ( .A1(n5202), .A2(n5040), .ZN(n3284) );
  OAI211_X1 U2675 ( .C1(n2556), .C2(n2554), .A(n2553), .B(n2552), .ZN(n3339)
         );
  NOR2_X1 U2676 ( .A1(n3339), .A2(n3399), .ZN(n3349) );
  NOR2_X1 U2677 ( .A1(n3410), .A2(n2765), .ZN(n3350) );
  XNOR2_X1 U2678 ( .A(n3353), .B(n3352), .ZN(n5093) );
  NOR2_X1 U2679 ( .A1(n5093), .A2(n5092), .ZN(n5091) );
  NAND2_X1 U2680 ( .A1(n5055), .A2(REG1_REG_5__SCAN_IN), .ZN(n2723) );
  NOR2_X1 U2681 ( .A1(n3441), .A2(n2562), .ZN(n3532) );
  AND2_X1 U2682 ( .A1(n5053), .A2(REG2_REG_7__SCAN_IN), .ZN(n2562) );
  NAND2_X1 U2683 ( .A1(n3541), .A2(n3540), .ZN(n3613) );
  INV_X1 U2684 ( .A(n3656), .ZN(n2700) );
  INV_X1 U2685 ( .A(n3620), .ZN(n2703) );
  AOI21_X1 U2686 ( .B1(REG2_REG_11__SCAN_IN), .B2(n5049), .A(n4171), .ZN(n4602) );
  NAND2_X1 U2687 ( .A1(n4174), .A2(n4175), .ZN(n4594) );
  INV_X1 U2688 ( .A(REG3_REG_13__SCAN_IN), .ZN(n4164) );
  NOR2_X1 U2689 ( .A1(n4614), .A2(n5259), .ZN(n2728) );
  NAND2_X1 U2690 ( .A1(n4620), .A2(n2544), .ZN(n2716) );
  NAND2_X1 U2691 ( .A1(n2716), .A2(REG2_REG_14__SCAN_IN), .ZN(n2715) );
  OR2_X1 U2692 ( .A1(n4644), .A2(n2564), .ZN(n2563) );
  AND2_X1 U2693 ( .A1(n5045), .A2(REG2_REG_15__SCAN_IN), .ZN(n2564) );
  INV_X1 U2694 ( .A(n5043), .ZN(n4679) );
  NAND2_X1 U2695 ( .A1(n4812), .A2(n2546), .ZN(n4752) );
  NAND2_X1 U2696 ( .A1(n4491), .A2(DATAI_27_), .ZN(n4770) );
  NAND2_X1 U2697 ( .A1(n4812), .A2(n2597), .ZN(n4769) );
  INV_X1 U2698 ( .A(n4839), .ZN(n4821) );
  AOI21_X1 U2699 ( .B1(n2655), .B2(n2653), .A(n2507), .ZN(n2652) );
  INV_X1 U2700 ( .A(n2655), .ZN(n2654) );
  NAND2_X1 U2701 ( .A1(n2684), .A2(n2524), .ZN(n4932) );
  AND2_X1 U2702 ( .A1(n4235), .A2(n4506), .ZN(n4960) );
  NAND2_X1 U2703 ( .A1(n5273), .A2(n4199), .ZN(n4200) );
  NOR2_X1 U2704 ( .A1(n3020), .A2(n4164), .ZN(n3041) );
  NOR2_X1 U2705 ( .A1(n4533), .A2(n2678), .ZN(n2677) );
  INV_X1 U2706 ( .A(n3635), .ZN(n2678) );
  INV_X1 U2707 ( .A(n2675), .ZN(n2674) );
  OAI21_X1 U2708 ( .B1(n4533), .B2(n2676), .A(n2680), .ZN(n2675) );
  NAND2_X1 U2709 ( .A1(n3636), .A2(n3635), .ZN(n2676) );
  INV_X1 U2710 ( .A(IR_REG_19__SCAN_IN), .ZN(n2812) );
  OAI211_X1 U2711 ( .C1(n3482), .C2(n2620), .A(n4422), .B(n2618), .ZN(n4211)
         );
  NAND2_X1 U2712 ( .A1(n2619), .A2(n4425), .ZN(n2618) );
  NAND2_X1 U2713 ( .A1(n2621), .A2(n4425), .ZN(n2620) );
  INV_X1 U2714 ( .A(n3487), .ZN(n2660) );
  NAND2_X1 U2715 ( .A1(n3285), .A2(n3465), .ZN(n5188) );
  INV_X1 U2716 ( .A(DATAI_0_), .ZN(n2590) );
  NAND2_X1 U2717 ( .A1(n3286), .A2(n3288), .ZN(n5264) );
  AND2_X1 U2718 ( .A1(n2878), .A2(n3313), .ZN(n4571) );
  OR2_X1 U2719 ( .A1(n2791), .A2(n2792), .ZN(n2795) );
  NAND2_X1 U2720 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_26__SCAN_IN), .ZN(n2792) );
  NOR2_X1 U2721 ( .A1(n2686), .A2(IR_REG_26__SCAN_IN), .ZN(n2685) );
  NAND2_X1 U2722 ( .A1(n2687), .A2(n2777), .ZN(n2686) );
  INV_X1 U2723 ( .A(n2779), .ZN(n2687) );
  NAND2_X1 U2724 ( .A1(n2798), .A2(IR_REG_31__SCAN_IN), .ZN(n2801) );
  XNOR2_X1 U2725 ( .A(n3275), .B(n2777), .ZN(n3329) );
  INV_X1 U2726 ( .A(n2605), .ZN(n2604) );
  NAND2_X1 U2727 ( .A1(n2776), .A2(n2754), .ZN(n2752) );
  INV_X1 U2728 ( .A(IR_REG_20__SCAN_IN), .ZN(n3807) );
  NAND2_X1 U2729 ( .A1(n3047), .A2(n2586), .ZN(n3113) );
  AND2_X1 U2730 ( .A1(n2587), .A2(n3803), .ZN(n2586) );
  NAND2_X1 U2731 ( .A1(n3047), .A2(n3996), .ZN(n3062) );
  INV_X1 U2732 ( .A(IR_REG_11__SCAN_IN), .ZN(n3795) );
  NAND2_X1 U2733 ( .A1(n2904), .A2(n2826), .ZN(n2905) );
  NAND2_X1 U2734 ( .A1(n3780), .A2(n2826), .ZN(n2827) );
  INV_X1 U2735 ( .A(IR_REG_3__SCAN_IN), .ZN(n3977) );
  AND4_X1 U2736 ( .A1(n2968), .A2(n2967), .A3(n2966), .A4(n2965), .ZN(n3643)
         );
  NAND2_X1 U2737 ( .A1(n3285), .A2(n2504), .ZN(n2649) );
  NAND2_X1 U2738 ( .A1(n2872), .A2(DATAI_1_), .ZN(n2648) );
  NAND2_X1 U2739 ( .A1(n2534), .A2(n2506), .ZN(n2746) );
  NAND2_X1 U2740 ( .A1(n2740), .A2(n2585), .ZN(n2584) );
  AND2_X1 U2741 ( .A1(n4491), .A2(DATAI_25_), .ZN(n4724) );
  INV_X1 U2742 ( .A(n5271), .ZN(n4414) );
  INV_X1 U2743 ( .A(n5272), .ZN(n4410) );
  NAND4_X1 U2744 ( .A1(n3220), .A2(n3219), .A3(n3218), .A4(n3217), .ZN(n4809)
         );
  NAND4_X1 U2745 ( .A1(n2790), .A2(n2789), .A3(n2788), .A4(n2787), .ZN(n4720)
         );
  INV_X1 U2746 ( .A(n3643), .ZN(n4586) );
  INV_X1 U2747 ( .A(n5056), .ZN(n3396) );
  NAND2_X1 U2748 ( .A1(n5100), .A2(REG1_REG_4__SCAN_IN), .ZN(n5098) );
  OR2_X1 U2749 ( .A1(n3442), .A2(n3581), .ZN(n2708) );
  NOR2_X1 U2750 ( .A1(n4172), .A2(n4173), .ZN(n4603) );
  INV_X1 U2751 ( .A(n5045), .ZN(n4648) );
  INV_X1 U2752 ( .A(n2692), .ZN(n4687) );
  OR2_X1 U2753 ( .A1(n3338), .A2(n4572), .ZN(n5090) );
  XNOR2_X1 U2754 ( .A(n2549), .B(n2547), .ZN(n2548) );
  NAND2_X1 U2755 ( .A1(n4690), .A2(n2718), .ZN(n2549) );
  NAND2_X1 U2756 ( .A1(n5042), .A2(REG1_REG_18__SCAN_IN), .ZN(n2718) );
  XNOR2_X1 U2757 ( .A(n2559), .B(n2690), .ZN(n4692) );
  INV_X1 U2758 ( .A(n4689), .ZN(n2690) );
  NAND2_X1 U2759 ( .A1(n2692), .A2(n2691), .ZN(n2559) );
  INV_X1 U2760 ( .A(n4671), .ZN(n5099) );
  NAND2_X1 U2761 ( .A1(n2663), .A2(n2664), .ZN(n4743) );
  AND2_X1 U2762 ( .A1(n2645), .A2(n2643), .ZN(n4980) );
  NOR2_X1 U2763 ( .A1(n4749), .A2(n2644), .ZN(n2643) );
  AND2_X1 U2764 ( .A1(n4750), .A2(n5154), .ZN(n2644) );
  NAND2_X1 U2765 ( .A1(n2588), .A2(n2811), .ZN(n5202) );
  OR2_X1 U2766 ( .A1(n2810), .A2(n2812), .ZN(n2588) );
  AND2_X1 U2767 ( .A1(n2969), .A2(n2955), .ZN(n5052) );
  INV_X1 U2768 ( .A(n4111), .ZN(n2569) );
  INV_X1 U2769 ( .A(n3040), .ZN(n2744) );
  INV_X1 U2770 ( .A(n4445), .ZN(n2627) );
  NOR2_X1 U2771 ( .A1(n2627), .A2(n2624), .ZN(n2623) );
  INV_X1 U2772 ( .A(n4444), .ZN(n2624) );
  INV_X1 U2773 ( .A(IR_REG_6__SCAN_IN), .ZN(n3787) );
  AND2_X1 U2774 ( .A1(n2739), .A2(n2731), .ZN(n2730) );
  NAND2_X1 U2775 ( .A1(n2732), .A2(n4351), .ZN(n2731) );
  NOR2_X1 U2776 ( .A1(n2521), .A2(n4406), .ZN(n2739) );
  INV_X1 U2777 ( .A(n3202), .ZN(n2732) );
  INV_X1 U2778 ( .A(n4351), .ZN(n2733) );
  INV_X1 U2779 ( .A(n2579), .ZN(n2578) );
  OAI21_X1 U2780 ( .B1(n4292), .B2(n2580), .A(n4373), .ZN(n2579) );
  INV_X1 U2781 ( .A(n3142), .ZN(n2580) );
  OR2_X1 U2782 ( .A1(n2890), .A2(n2834), .ZN(n2892) );
  INV_X1 U2783 ( .A(n2572), .ZN(n2571) );
  OAI21_X1 U2784 ( .B1(n2912), .B2(n2573), .A(n3546), .ZN(n2572) );
  AND2_X1 U2785 ( .A1(n3212), .A2(n3211), .ZN(n3213) );
  INV_X1 U2786 ( .A(REG2_REG_1__SCAN_IN), .ZN(n2555) );
  AND2_X1 U2787 ( .A1(n4770), .A2(n4785), .ZN(n2597) );
  AND2_X1 U2788 ( .A1(n3185), .A2(REG3_REG_24__SCAN_IN), .ZN(n3204) );
  AND2_X1 U2789 ( .A1(n3156), .A2(REG3_REG_21__SCAN_IN), .ZN(n3170) );
  AND2_X1 U2790 ( .A1(n3143), .A2(REG3_REG_20__SCAN_IN), .ZN(n3156) );
  INV_X1 U2791 ( .A(REG3_REG_10__SCAN_IN), .ZN(n3746) );
  NAND2_X1 U2792 ( .A1(n4907), .A2(n4889), .ZN(n2656) );
  INV_X1 U2793 ( .A(n4304), .ZN(n3478) );
  INV_X1 U2794 ( .A(IR_REG_30__SCAN_IN), .ZN(n3827) );
  NAND2_X1 U2795 ( .A1(n2778), .A2(n4011), .ZN(n2779) );
  NAND3_X1 U2796 ( .A1(n2772), .A2(n3980), .A3(n2769), .ZN(n2605) );
  INV_X1 U2797 ( .A(IR_REG_17__SCAN_IN), .ZN(n3803) );
  INV_X1 U2798 ( .A(IR_REG_9__SCAN_IN), .ZN(n3988) );
  INV_X1 U2799 ( .A(IR_REG_2__SCAN_IN), .ZN(n3780) );
  INV_X1 U2800 ( .A(IR_REG_1__SCAN_IN), .ZN(n2558) );
  NAND2_X1 U2801 ( .A1(IR_REG_0__SCAN_IN), .A2(IR_REG_31__SCAN_IN), .ZN(n2550)
         );
  NAND2_X1 U2802 ( .A1(n2749), .A2(n2748), .ZN(n4269) );
  AOI21_X1 U2803 ( .B1(n4310), .B2(n2499), .A(n2508), .ZN(n2748) );
  OAI21_X1 U2804 ( .B1(n4349), .B2(n2735), .A(n2734), .ZN(n4264) );
  AND2_X1 U2805 ( .A1(n2737), .A2(n4407), .ZN(n2734) );
  OAI21_X1 U2806 ( .B1(n3203), .B2(n2733), .A(n2730), .ZN(n2735) );
  NAND2_X1 U2807 ( .A1(n2738), .A2(n2530), .ZN(n2737) );
  NAND2_X1 U2808 ( .A1(n3683), .A2(n3684), .ZN(n2747) );
  AND2_X1 U2809 ( .A1(n2996), .A2(REG3_REG_11__SCAN_IN), .ZN(n3009) );
  OAI22_X1 U2810 ( .A1(n5187), .A2(n3254), .B1(n2830), .B2(n5150), .ZN(n2855)
         );
  NAND2_X1 U2811 ( .A1(n3203), .A2(n3202), .ZN(n4350) );
  INV_X1 U2812 ( .A(REG3_REG_9__SCAN_IN), .ZN(n3770) );
  NAND2_X1 U2813 ( .A1(n4291), .A2(n4292), .ZN(n4290) );
  NAND2_X1 U2814 ( .A1(n4112), .A2(n4111), .ZN(n4158) );
  NAND2_X1 U2815 ( .A1(n2756), .A2(n2755), .ZN(n4396) );
  AND2_X1 U2816 ( .A1(n2763), .A2(n2757), .ZN(n2755) );
  NAND2_X1 U2817 ( .A1(n2574), .A2(n2912), .ZN(n3522) );
  NAND2_X1 U2818 ( .A1(n3069), .A2(n3070), .ZN(n5278) );
  NAND2_X1 U2819 ( .A1(n3072), .A2(n3071), .ZN(n5279) );
  INV_X1 U2820 ( .A(n3070), .ZN(n3071) );
  AND4_X1 U2821 ( .A1(n2936), .A2(n2935), .A3(n2934), .A4(n2933), .ZN(n3555)
         );
  NOR2_X1 U2822 ( .A1(n3341), .A2(n3340), .ZN(n3361) );
  NOR2_X1 U2823 ( .A1(n3349), .A2(n3348), .ZN(n3412) );
  NOR2_X1 U2824 ( .A1(n3361), .A2(n2727), .ZN(n3408) );
  AND2_X1 U2825 ( .A1(n3347), .A2(REG1_REG_1__SCAN_IN), .ZN(n2727) );
  OAI22_X1 U2826 ( .A1(n3408), .A2(n3409), .B1(n5137), .B2(n3417), .ZN(n3362)
         );
  NAND2_X1 U2827 ( .A1(n2711), .A2(n2712), .ZN(n3356) );
  NAND2_X1 U2828 ( .A1(n2694), .A2(n2502), .ZN(n2695) );
  AND2_X1 U2829 ( .A1(n3357), .A2(REG2_REG_6__SCAN_IN), .ZN(n2694) );
  OAI21_X1 U2830 ( .B1(n3419), .B2(n3367), .A(n2516), .ZN(n3371) );
  INV_X1 U2831 ( .A(n3366), .ZN(n3368) );
  NAND2_X1 U2832 ( .A1(n3371), .A2(n3370), .ZN(n3443) );
  NAND2_X1 U2833 ( .A1(n3613), .A2(n2527), .ZN(n3658) );
  NAND2_X1 U2834 ( .A1(n3663), .A2(n3662), .ZN(n4174) );
  XNOR2_X1 U2835 ( .A(n4594), .B(n4601), .ZN(n4176) );
  INV_X1 U2836 ( .A(REG3_REG_15__SCAN_IN), .ZN(n4639) );
  OAI22_X1 U2837 ( .A1(n4634), .A2(n4633), .B1(n4635), .B2(n2717), .ZN(n4638)
         );
  INV_X1 U2838 ( .A(n4616), .ZN(n4635) );
  NAND2_X1 U2839 ( .A1(n4662), .A2(n4663), .ZN(n4664) );
  INV_X1 U2840 ( .A(n2563), .ZN(n4661) );
  XNOR2_X1 U2841 ( .A(n4655), .B(n5044), .ZN(n4649) );
  NOR2_X1 U2842 ( .A1(n4649), .A2(REG1_REG_16__SCAN_IN), .ZN(n4656) );
  INV_X1 U2843 ( .A(REG3_REG_17__SCAN_IN), .ZN(n4342) );
  NAND2_X1 U2844 ( .A1(n5042), .A2(REG2_REG_18__SCAN_IN), .ZN(n2691) );
  NAND2_X1 U2845 ( .A1(n4733), .A2(n4732), .ZN(n5325) );
  INV_X1 U2846 ( .A(n4752), .ZN(n4733) );
  INV_X1 U2847 ( .A(n4748), .ZN(n2647) );
  INV_X1 U2848 ( .A(n4809), .ZN(n4761) );
  AOI21_X1 U2849 ( .B1(n2609), .B2(n4701), .A(n4702), .ZN(n2608) );
  INV_X1 U2850 ( .A(n2613), .ZN(n4803) );
  INV_X1 U2851 ( .A(n4724), .ZN(n4810) );
  OR2_X1 U2852 ( .A1(n4699), .A2(n4698), .ZN(n4820) );
  NAND2_X1 U2853 ( .A1(n4491), .A2(DATAI_23_), .ZN(n4716) );
  AOI21_X1 U2854 ( .B1(n4845), .B2(n4233), .A(n4232), .ZN(n4719) );
  NAND2_X1 U2855 ( .A1(n2595), .A2(n2594), .ZN(n2593) );
  NOR2_X1 U2856 ( .A1(n4376), .A2(n4385), .ZN(n2594) );
  INV_X1 U2857 ( .A(n2596), .ZN(n2595) );
  AND4_X1 U2858 ( .A1(n3175), .A2(n3174), .A3(n3173), .A4(n3172), .ZN(n4861)
         );
  NAND2_X1 U2859 ( .A1(n2872), .A2(DATAI_21_), .ZN(n4867) );
  NAND2_X1 U2860 ( .A1(n2638), .A2(n2639), .ZN(n2637) );
  NAND2_X1 U2861 ( .A1(n2638), .A2(n2635), .ZN(n2634) );
  NOR3_X1 U2862 ( .A1(n4917), .A2(n4376), .A3(n4294), .ZN(n4882) );
  NOR2_X1 U2863 ( .A1(n4917), .A2(n4294), .ZN(n4896) );
  NAND2_X1 U2864 ( .A1(n4947), .A2(n2639), .ZN(n4911) );
  OR2_X1 U2865 ( .A1(n4938), .A2(n4916), .ZN(n4917) );
  NAND2_X1 U2866 ( .A1(n4955), .A2(n4936), .ZN(n4938) );
  NOR2_X1 U2867 ( .A1(n3054), .A2(n4639), .ZN(n3074) );
  NAND2_X1 U2868 ( .A1(n3074), .A2(REG3_REG_16__SCAN_IN), .ZN(n3087) );
  NAND2_X1 U2869 ( .A1(n4948), .A2(n4960), .ZN(n4947) );
  NOR2_X1 U2870 ( .A1(n4203), .A2(n5277), .ZN(n4954) );
  NAND2_X1 U2871 ( .A1(n3041), .A2(REG3_REG_14__SCAN_IN), .ZN(n3054) );
  NAND2_X1 U2872 ( .A1(n4149), .A2(n4148), .ZN(n4150) );
  OR2_X1 U2873 ( .A1(n4150), .A2(n4198), .ZN(n4203) );
  AND4_X1 U2874 ( .A1(n3024), .A2(n3023), .A3(n3022), .A4(n3021), .ZN(n4128)
         );
  NAND2_X1 U2875 ( .A1(n4096), .A2(n4445), .ZN(n4126) );
  AND2_X1 U2876 ( .A1(n4461), .A2(n4134), .ZN(n4536) );
  NOR2_X1 U2877 ( .A1(n4103), .A2(n4120), .ZN(n4149) );
  NAND2_X1 U2878 ( .A1(n2589), .A2(n4101), .ZN(n4103) );
  AND4_X1 U2879 ( .A1(n2984), .A2(n2983), .A3(n2982), .A4(n2981), .ZN(n3677)
         );
  AND4_X1 U2880 ( .A1(n3014), .A2(n3013), .A3(n3012), .A4(n3011), .ZN(n4139)
         );
  NAND2_X1 U2881 ( .A1(n3675), .A2(n4444), .ZN(n3676) );
  NAND2_X1 U2882 ( .A1(n3676), .A2(n4535), .ZN(n4096) );
  INV_X1 U2883 ( .A(n4282), .ZN(n3669) );
  AND4_X1 U2884 ( .A1(n3002), .A2(n3001), .A3(n3000), .A4(n2999), .ZN(n4102)
         );
  AND3_X1 U2885 ( .A1(n5181), .A2(n2501), .A3(n2518), .ZN(n3595) );
  NAND2_X1 U2886 ( .A1(n2633), .A2(n4537), .ZN(n2632) );
  NAND2_X1 U2887 ( .A1(n2633), .A2(n2628), .ZN(n2629) );
  NAND2_X1 U2888 ( .A1(n5184), .A2(n4430), .ZN(n2633) );
  NAND2_X1 U2889 ( .A1(n2631), .A2(n4430), .ZN(n3554) );
  OR2_X1 U2890 ( .A1(n5185), .A2(n5184), .ZN(n2631) );
  NAND2_X1 U2891 ( .A1(n5181), .A2(n5180), .ZN(n5183) );
  NAND2_X1 U2892 ( .A1(n5181), .A2(n2501), .ZN(n3564) );
  AND2_X1 U2893 ( .A1(REG3_REG_4__SCAN_IN), .A2(REG3_REG_3__SCAN_IN), .ZN(
        n2898) );
  INV_X1 U2894 ( .A(n5158), .ZN(n5150) );
  AND2_X1 U2895 ( .A1(n5151), .A2(n5150), .ZN(n5181) );
  INV_X1 U2896 ( .A(n5188), .ZN(n5154) );
  OR2_X1 U2897 ( .A1(n3494), .A2(n3493), .ZN(n4217) );
  AND4_X2 U2898 ( .A1(n2861), .A2(n2860), .A3(n2859), .A4(n2858), .ZN(n5110)
         );
  NAND2_X1 U2899 ( .A1(n2866), .A2(REG3_REG_1__SCAN_IN), .ZN(n2861) );
  OAI21_X1 U2900 ( .B1(n3274), .B2(n3273), .A(n3317), .ZN(n4976) );
  AND2_X1 U2901 ( .A1(n4571), .A2(n3428), .ZN(n4977) );
  NAND2_X1 U2902 ( .A1(n2656), .A2(n2655), .ZN(n5010) );
  NAND2_X1 U2903 ( .A1(n4226), .A2(n4225), .ZN(n4961) );
  INV_X1 U2904 ( .A(n5264), .ZN(n5333) );
  INV_X1 U2905 ( .A(n2599), .ZN(n2598) );
  OAI22_X1 U2906 ( .A1(n2601), .A2(n2600), .B1(IR_REG_29__SCAN_IN), .B2(
        IR_REG_31__SCAN_IN), .ZN(n2599) );
  NAND2_X1 U2907 ( .A1(IR_REG_31__SCAN_IN), .A2(IR_REG_29__SCAN_IN), .ZN(n2600) );
  INV_X1 U2908 ( .A(IR_REG_8__SCAN_IN), .ZN(n2985) );
  AND2_X1 U2909 ( .A1(n2550), .A2(IR_REG_1__SCAN_IN), .ZN(n2556) );
  NAND2_X1 U2910 ( .A1(n2583), .A2(n2941), .ZN(n4253) );
  NAND2_X1 U2911 ( .A1(n4159), .A2(n3040), .ZN(n4183) );
  INV_X1 U2912 ( .A(n4716), .ZN(n4273) );
  NAND2_X1 U2913 ( .A1(n4281), .A2(n4280), .ZN(n4279) );
  NAND2_X1 U2914 ( .A1(n3309), .A2(n3308), .ZN(n3310) );
  AND2_X1 U2915 ( .A1(n4253), .A2(n2944), .ZN(n3603) );
  OR2_X1 U2916 ( .A1(n4309), .A2(n4310), .ZN(n4313) );
  INV_X1 U2917 ( .A(n4822), .ZN(n4827) );
  MUX2_X1 U2918 ( .A(n5096), .B(DATAI_4_), .S(n2872), .Z(n5158) );
  AOI21_X1 U2919 ( .B1(n2761), .B2(n4251), .A(n2528), .ZN(n2582) );
  INV_X1 U2920 ( .A(n5107), .ZN(n4419) );
  NAND2_X1 U2921 ( .A1(n4290), .A2(n3142), .ZN(n4375) );
  NAND2_X1 U2922 ( .A1(n4313), .A2(n4308), .ZN(n4383) );
  NAND2_X1 U2923 ( .A1(n4279), .A2(n2995), .ZN(n3686) );
  INV_X1 U2924 ( .A(n4918), .ZN(n4916) );
  NAND2_X1 U2925 ( .A1(n3522), .A2(n2915), .ZN(n3547) );
  AOI21_X1 U2926 ( .B1(n2736), .B2(n2740), .A(n2530), .ZN(n4409) );
  NOR2_X1 U2927 ( .A1(n4349), .A2(n2521), .ZN(n2736) );
  NAND2_X1 U2928 ( .A1(n3302), .A2(STATE_REG_SCAN_IN), .ZN(n5287) );
  INV_X1 U2929 ( .A(n4417), .ZN(n5282) );
  NAND4_X1 U2930 ( .A1(n3233), .A2(n3232), .A3(n3231), .A4(n3230), .ZN(n4787)
         );
  INV_X1 U2931 ( .A(n4823), .ZN(n4725) );
  NAND4_X1 U2932 ( .A1(n3189), .A2(n3188), .A3(n3187), .A4(n3186), .ZN(n4839)
         );
  INV_X1 U2933 ( .A(n4139), .ZN(n4583) );
  INV_X1 U2934 ( .A(n4102), .ZN(n4584) );
  INV_X1 U2935 ( .A(n3677), .ZN(n4585) );
  INV_X1 U2936 ( .A(n3555), .ZN(n4588) );
  NAND2_X1 U2937 ( .A1(n2865), .A2(REG1_REG_3__SCAN_IN), .ZN(n2823) );
  OR2_X1 U2938 ( .A1(n2878), .A2(n3319), .ZN(n4592) );
  XNOR2_X1 U2939 ( .A(n3364), .B(n3352), .ZN(n5100) );
  NOR2_X1 U2940 ( .A1(n5091), .A2(n3354), .ZN(n3384) );
  INV_X1 U2941 ( .A(n2726), .ZN(n3380) );
  INV_X1 U2942 ( .A(n2724), .ZN(n3378) );
  INV_X1 U2943 ( .A(n2695), .ZN(n3422) );
  XNOR2_X1 U2944 ( .A(n3366), .B(n5054), .ZN(n3419) );
  NAND2_X1 U2945 ( .A1(n2695), .A2(n3357), .ZN(n2697) );
  AND2_X1 U2946 ( .A1(n2697), .A2(n2696), .ZN(n3441) );
  INV_X1 U2947 ( .A(n3359), .ZN(n2696) );
  INV_X1 U2948 ( .A(n3534), .ZN(n2707) );
  OAI21_X1 U2949 ( .B1(n3442), .B2(n2706), .A(n2705), .ZN(n3617) );
  NAND2_X1 U2950 ( .A1(n2709), .A2(REG2_REG_8__SCAN_IN), .ZN(n2706) );
  INV_X1 U2951 ( .A(n3535), .ZN(n2709) );
  NAND2_X1 U2952 ( .A1(n2702), .A2(n2509), .ZN(n2704) );
  OAI21_X1 U2953 ( .B1(n2701), .B2(n2699), .A(n2698), .ZN(n4171) );
  INV_X1 U2954 ( .A(n2702), .ZN(n2701) );
  OR2_X1 U2955 ( .A1(n2509), .A2(n3656), .ZN(n2698) );
  XNOR2_X1 U2956 ( .A(n4602), .B(n4601), .ZN(n4172) );
  INV_X1 U2957 ( .A(n2566), .ZN(n4609) );
  AND2_X1 U2958 ( .A1(n4598), .A2(n2729), .ZN(n4615) );
  AOI21_X1 U2959 ( .B1(n4614), .B2(n5259), .A(n4597), .ZN(n2729) );
  XNOR2_X1 U2960 ( .A(n4616), .B(n5046), .ZN(n4634) );
  NOR2_X1 U2961 ( .A1(n2715), .A2(n4629), .ZN(n4628) );
  AND2_X1 U2962 ( .A1(n2715), .A2(n2714), .ZN(n4632) );
  XNOR2_X1 U2963 ( .A(n2563), .B(n4660), .ZN(n4645) );
  NAND2_X1 U2964 ( .A1(n4645), .A2(n4959), .ZN(n4662) );
  OAI21_X1 U2965 ( .B1(n4649), .B2(n2720), .A(n2719), .ZN(n4678) );
  NAND2_X1 U2966 ( .A1(n2722), .A2(n2721), .ZN(n2720) );
  NAND2_X1 U2967 ( .A1(n4657), .A2(n2722), .ZN(n2719) );
  INV_X1 U2968 ( .A(n4659), .ZN(n2722) );
  NAND2_X1 U2969 ( .A1(n2662), .A2(n2661), .ZN(n4731) );
  AOI21_X1 U2970 ( .B1(n2498), .B2(n2666), .A(n2531), .ZN(n2661) );
  AND2_X1 U2971 ( .A1(n4812), .A2(n4785), .ZN(n4771) );
  OR2_X1 U2972 ( .A1(n4851), .A2(n4850), .ZN(n5000) );
  OAI21_X1 U2973 ( .B1(n4907), .B2(n2654), .A(n2652), .ZN(n4874) );
  AND2_X1 U2974 ( .A1(n2684), .A2(n2683), .ZN(n4934) );
  NAND2_X1 U2975 ( .A1(n2672), .A2(n2674), .ZN(n3671) );
  NAND2_X1 U2976 ( .A1(n3637), .A2(n2677), .ZN(n2672) );
  NAND2_X1 U2977 ( .A1(n2673), .A2(n3635), .ZN(n3670) );
  OR2_X1 U2978 ( .A1(n3637), .A2(n3636), .ZN(n2673) );
  AND2_X1 U2979 ( .A1(n5208), .A2(n5199), .ZN(n4935) );
  INV_X1 U2980 ( .A(n4974), .ZN(n3289) );
  NAND2_X1 U2981 ( .A1(n3510), .A2(n3509), .ZN(n4210) );
  INV_X1 U2982 ( .A(n5210), .ZN(n5118) );
  OR2_X1 U2983 ( .A1(n5019), .A2(n4978), .ZN(n5335) );
  INV_X2 U2984 ( .A(n5335), .ZN(n5337) );
  NAND2_X1 U2985 ( .A1(n2642), .A2(n5304), .ZN(n2641) );
  INV_X1 U2986 ( .A(n4981), .ZN(n2642) );
  OR2_X1 U2987 ( .A1(n5019), .A2(n5018), .ZN(n5338) );
  INV_X2 U2988 ( .A(n5338), .ZN(n5341) );
  NAND2_X1 U2989 ( .A1(n4571), .A2(n3318), .ZN(n5086) );
  INV_X1 U2990 ( .A(n2782), .ZN(n5033) );
  NAND2_X1 U2991 ( .A1(n2821), .A2(n4016), .ZN(n2819) );
  NOR2_X1 U2992 ( .A1(n2797), .A2(n2796), .ZN(n5037) );
  NAND2_X1 U2993 ( .A1(n2795), .A2(n2794), .ZN(n2797) );
  NAND2_X1 U2994 ( .A1(n3093), .A2(n2793), .ZN(n2794) );
  XNOR2_X1 U2995 ( .A(n2800), .B(IR_REG_25__SCAN_IN), .ZN(n5038) );
  XNOR2_X1 U2996 ( .A(n2801), .B(IR_REG_24__SCAN_IN), .ZN(n5039) );
  AND2_X1 U2997 ( .A1(n3329), .A2(STATE_REG_SCAN_IN), .ZN(n3313) );
  NOR2_X1 U2998 ( .A1(n2816), .A2(n2815), .ZN(n5040) );
  NOR2_X1 U2999 ( .A1(n2809), .A2(n2808), .ZN(n5041) );
  NAND2_X1 U3000 ( .A1(n2811), .A2(IR_REG_31__SCAN_IN), .ZN(n2805) );
  AND2_X1 U3001 ( .A1(n3096), .A2(n3113), .ZN(n5043) );
  AND2_X1 U3002 ( .A1(n3065), .A2(n3080), .ZN(n5045) );
  AND2_X1 U3003 ( .A1(n3015), .A2(n3005), .ZN(n5049) );
  XNOR2_X1 U3004 ( .A(n2952), .B(IR_REG_7__SCAN_IN), .ZN(n5053) );
  AND2_X1 U3005 ( .A1(n2908), .A2(n2907), .ZN(n5055) );
  AND2_X1 U3006 ( .A1(n2853), .A2(n2829), .ZN(n5056) );
  OR2_X1 U3007 ( .A1(n2826), .A2(n3093), .ZN(n2840) );
  XNOR2_X1 U3008 ( .A(n2584), .B(n2522), .ZN(n4328) );
  INV_X1 U3009 ( .A(n2708), .ZN(n3533) );
  INV_X1 U3010 ( .A(n2561), .ZN(n4676) );
  AOI22_X1 U3011 ( .A1(n4692), .A2(n4691), .B1(n2548), .B2(n5099), .ZN(n4695)
         );
  AND2_X1 U3012 ( .A1(n4747), .A2(n2664), .ZN(n2498) );
  NOR2_X1 U3013 ( .A1(n4384), .A2(n2750), .ZN(n2499) );
  OR2_X1 U3014 ( .A1(n4917), .A2(n2593), .ZN(n2500) );
  AND2_X1 U3015 ( .A1(n5180), .A2(n3503), .ZN(n2501) );
  NAND3_X1 U3016 ( .A1(n2711), .A2(n2710), .A3(n2712), .ZN(n2502) );
  AND2_X1 U3017 ( .A1(n4710), .A2(n3347), .ZN(n2504) );
  INV_X1 U3018 ( .A(n4701), .ZN(n2612) );
  INV_X1 U3019 ( .A(n2688), .ZN(n2796) );
  NAND2_X1 U3020 ( .A1(n2713), .A2(REG2_REG_4__SCAN_IN), .ZN(n2505) );
  INV_X1 U3021 ( .A(n4764), .ZN(n2666) );
  OR2_X1 U3022 ( .A1(n3683), .A2(n3684), .ZN(n2506) );
  OR2_X1 U3023 ( .A1(n2802), .A2(n3093), .ZN(n3047) );
  INV_X1 U3024 ( .A(n3687), .ZN(n4101) );
  AND2_X1 U3025 ( .A1(n4580), .A2(n4294), .ZN(n2507) );
  INV_X1 U3026 ( .A(n4470), .ZN(n4235) );
  AND2_X1 U3027 ( .A1(n3182), .A2(n3181), .ZN(n2508) );
  INV_X1 U3028 ( .A(n2830), .ZN(n2956) );
  NAND2_X2 U3029 ( .A1(n2878), .A2(n2818), .ZN(n2830) );
  NOR2_X1 U3030 ( .A1(n3025), .A2(n2751), .ZN(n2808) );
  OR2_X1 U3031 ( .A1(n3619), .A2(n3618), .ZN(n2509) );
  NOR2_X1 U3032 ( .A1(n2785), .A2(n5036), .ZN(n2867) );
  INV_X1 U3033 ( .A(n5110), .ZN(n3457) );
  NOR2_X1 U3034 ( .A1(n3203), .A2(n3202), .ZN(n4349) );
  INV_X1 U3035 ( .A(n4349), .ZN(n2585) );
  NAND3_X1 U3036 ( .A1(n2603), .A2(n2606), .A3(n2602), .ZN(n2814) );
  OR2_X1 U3037 ( .A1(n5192), .A2(n5155), .ZN(n2510) );
  NOR2_X1 U3038 ( .A1(n2752), .A2(n3025), .ZN(n2806) );
  NAND2_X1 U3039 ( .A1(n4760), .A2(n4764), .ZN(n4759) );
  OR2_X1 U3040 ( .A1(n5156), .A2(n4218), .ZN(n2511) );
  AND2_X1 U3041 ( .A1(n2613), .A2(n2612), .ZN(n2512) );
  NAND2_X1 U3042 ( .A1(n2651), .A2(n2650), .ZN(n4845) );
  NOR2_X1 U3043 ( .A1(n4656), .A2(n4657), .ZN(n2513) );
  NAND2_X1 U3044 ( .A1(n2551), .A2(n2557), .ZN(n3347) );
  AND2_X1 U3045 ( .A1(n3604), .A2(n2944), .ZN(n2761) );
  NAND2_X1 U3046 ( .A1(n3356), .A2(n5054), .ZN(n3357) );
  INV_X1 U3047 ( .A(n3605), .ZN(n3585) );
  AND2_X1 U3048 ( .A1(n5055), .A2(REG2_REG_5__SCAN_IN), .ZN(n2514) );
  INV_X1 U3049 ( .A(IR_REG_14__SCAN_IN), .ZN(n3996) );
  OR2_X1 U3050 ( .A1(n2503), .A2(IR_REG_29__SCAN_IN), .ZN(n2515) );
  OR2_X1 U3051 ( .A1(n3368), .A2(n2710), .ZN(n2516) );
  INV_X1 U3052 ( .A(IR_REG_22__SCAN_IN), .ZN(n3815) );
  INV_X1 U3053 ( .A(n2670), .ZN(n2669) );
  NAND2_X1 U3054 ( .A1(n2674), .A2(n2671), .ZN(n2670) );
  AND2_X1 U3055 ( .A1(n2677), .A2(n2679), .ZN(n2517) );
  OAI21_X1 U3056 ( .B1(n3113), .B2(IR_REG_18__SCAN_IN), .A(IR_REG_31__SCAN_IN), 
        .ZN(n2810) );
  INV_X1 U3057 ( .A(n2915), .ZN(n2573) );
  AND2_X1 U3058 ( .A1(n3559), .A2(n3585), .ZN(n2518) );
  INV_X1 U3059 ( .A(n2610), .ZN(n2609) );
  NAND2_X1 U3060 ( .A1(n2617), .A2(n2611), .ZN(n2610) );
  AND2_X1 U3061 ( .A1(IR_REG_1__SCAN_IN), .A2(REG2_REG_1__SCAN_IN), .ZN(n2519)
         );
  AND2_X1 U3062 ( .A1(IR_REG_31__SCAN_IN), .A2(REG2_REG_1__SCAN_IN), .ZN(n2520) );
  INV_X1 U3063 ( .A(n5054), .ZN(n2710) );
  XNOR2_X1 U3064 ( .A(n2805), .B(n3807), .ZN(n3286) );
  AND2_X1 U3065 ( .A1(n4322), .A2(n3213), .ZN(n2521) );
  NAND2_X1 U3066 ( .A1(n2756), .A2(n2757), .ZN(n4338) );
  NAND3_X1 U3067 ( .A1(n5037), .A2(n5038), .A3(n5039), .ZN(n2878) );
  NAND2_X1 U3068 ( .A1(n4343), .A2(n4918), .ZN(n4229) );
  XOR2_X1 U3069 ( .A(n4322), .B(n4321), .Z(n2522) );
  NAND2_X1 U3070 ( .A1(n4158), .A2(n3035), .ZN(n4159) );
  AND2_X1 U3071 ( .A1(n4862), .A2(n4881), .ZN(n2523) );
  NAND2_X1 U3072 ( .A1(n2606), .A2(n2604), .ZN(n3025) );
  AND2_X1 U3073 ( .A1(n4933), .A2(n2683), .ZN(n2524) );
  AND2_X1 U3074 ( .A1(n3053), .A2(n3052), .ZN(n2525) );
  AND2_X1 U3075 ( .A1(n4476), .A2(n2634), .ZN(n2526) );
  INV_X1 U3076 ( .A(n4223), .ZN(n4950) );
  OR2_X1 U3077 ( .A1(n3614), .A2(n3539), .ZN(n2527) );
  INV_X1 U3078 ( .A(n2592), .ZN(n4866) );
  NOR3_X1 U3079 ( .A1(n4917), .A2(n2596), .A3(n4376), .ZN(n2592) );
  AND2_X1 U3080 ( .A1(n2962), .A2(n2961), .ZN(n2528) );
  NAND2_X1 U3081 ( .A1(n4396), .A2(n4395), .ZN(n2529) );
  AND2_X1 U3082 ( .A1(n4621), .A2(n5046), .ZN(n4629) );
  AND2_X1 U3083 ( .A1(n3214), .A2(n4321), .ZN(n2530) );
  INV_X1 U3084 ( .A(n4471), .ZN(n4236) );
  NOR2_X1 U3085 ( .A1(n4729), .A2(n4744), .ZN(n2531) );
  AND2_X1 U3086 ( .A1(n4745), .A2(n4770), .ZN(n2532) );
  AND2_X1 U3087 ( .A1(n4280), .A2(n2506), .ZN(n2533) );
  NAND2_X1 U3088 ( .A1(n2995), .A2(n2747), .ZN(n2534) );
  AND2_X1 U3089 ( .A1(n4947), .A2(n4235), .ZN(n2535) );
  OR2_X1 U3090 ( .A1(n4223), .A2(n4222), .ZN(n2536) );
  AND2_X1 U3091 ( .A1(n3047), .A2(n2587), .ZN(n3092) );
  AND2_X1 U3092 ( .A1(n4706), .A2(n4523), .ZN(n4742) );
  INV_X1 U3093 ( .A(n2743), .ZN(n2742) );
  OAI21_X1 U3094 ( .B1(n3035), .B2(n2744), .A(n4182), .ZN(n2743) );
  AND2_X1 U3095 ( .A1(n2656), .A2(n4229), .ZN(n2537) );
  INV_X1 U3096 ( .A(n4889), .ZN(n2653) );
  NOR2_X1 U3097 ( .A1(n3648), .A2(n4282), .ZN(n2589) );
  INV_X1 U3098 ( .A(IR_REG_13__SCAN_IN), .ZN(n2754) );
  AND3_X1 U3099 ( .A1(n5181), .A2(n2501), .A3(n3559), .ZN(n2538) );
  NOR3_X1 U3100 ( .A1(n3595), .A2(n3579), .A3(n5264), .ZN(n2539) );
  INV_X1 U3101 ( .A(n4308), .ZN(n2750) );
  OAI21_X1 U3102 ( .B1(n5178), .B2(n3514), .A(n2510), .ZN(n3561) );
  NAND2_X1 U3103 ( .A1(n3513), .A2(n3512), .ZN(n5178) );
  CLKBUF_X1 U3104 ( .A(n3458), .Z(n3482) );
  NAND2_X1 U3105 ( .A1(n4253), .A2(n2761), .ZN(n3602) );
  INV_X1 U3106 ( .A(n4898), .ZN(n4294) );
  AND2_X1 U3107 ( .A1(n2708), .A2(n2707), .ZN(n2540) );
  AND2_X1 U3108 ( .A1(n2672), .A2(n2669), .ZN(n2541) );
  AND2_X1 U3109 ( .A1(n2893), .A2(n2894), .ZN(n2542) );
  AND2_X1 U3110 ( .A1(n2704), .A2(n2509), .ZN(n2543) );
  INV_X1 U3111 ( .A(n5046), .ZN(n2717) );
  INV_X1 U3112 ( .A(IR_REG_23__SCAN_IN), .ZN(n2777) );
  INV_X1 U3113 ( .A(n4751), .ZN(n4744) );
  AND2_X1 U3114 ( .A1(n3472), .A2(n3471), .ZN(n5194) );
  INV_X1 U3115 ( .A(n5304), .ZN(n5294) );
  NAND2_X1 U3116 ( .A1(n4968), .A2(n5140), .ZN(n5304) );
  AND2_X1 U3117 ( .A1(n4619), .A2(n2717), .ZN(n2544) );
  NOR2_X1 U3118 ( .A1(n3384), .A2(n3383), .ZN(n2545) );
  AND2_X1 U3119 ( .A1(n2597), .A2(n4744), .ZN(n2546) );
  INV_X1 U3120 ( .A(IR_REG_0__SCAN_IN), .ZN(n2591) );
  XOR2_X1 U3121 ( .A(n5202), .B(REG1_REG_19__SCAN_IN), .Z(n2547) );
  INV_X1 U3122 ( .A(REG1_REG_16__SCAN_IN), .ZN(n2721) );
  INV_X1 U3123 ( .A(n3660), .ZN(n3663) );
  MUX2_X1 U3124 ( .A(n5130), .B(REG1_REG_1__SCAN_IN), .S(n3347), .Z(n3341) );
  NAND2_X1 U3125 ( .A1(n2550), .A2(n2519), .ZN(n2552) );
  XNOR2_X1 U3126 ( .A(n3658), .B(n3618), .ZN(n3659) );
  NAND3_X1 U3127 ( .A1(IR_REG_0__SCAN_IN), .A2(n2558), .A3(IR_REG_31__SCAN_IN), 
        .ZN(n2557) );
  NAND3_X1 U3128 ( .A1(IR_REG_0__SCAN_IN), .A2(n2520), .A3(n2558), .ZN(n2553)
         );
  INV_X1 U3129 ( .A(n2556), .ZN(n2551) );
  NAND2_X1 U3130 ( .A1(n2557), .A2(n2555), .ZN(n2554) );
  NOR2_X1 U3131 ( .A1(n3389), .A2(n3351), .ZN(n3353) );
  OAI21_X1 U3132 ( .B1(n4112), .B2(n2743), .A(n2567), .ZN(n3069) );
  INV_X1 U3133 ( .A(n3524), .ZN(n2574) );
  NAND2_X1 U3134 ( .A1(n2570), .A2(n2571), .ZN(n2928) );
  NAND2_X1 U3135 ( .A1(n3524), .A2(n2915), .ZN(n2570) );
  NAND2_X1 U3136 ( .A1(n4291), .A2(n2578), .ZN(n2575) );
  NAND2_X1 U3137 ( .A1(n2575), .A2(n2576), .ZN(n4309) );
  NAND2_X1 U3138 ( .A1(n4252), .A2(n2761), .ZN(n2581) );
  NAND2_X1 U3139 ( .A1(n2581), .A2(n2582), .ZN(n3627) );
  INV_X1 U3140 ( .A(n4252), .ZN(n2583) );
  MUX2_X1 U3141 ( .A(n2591), .B(n2590), .S(n2872), .Z(n5107) );
  XNOR2_X2 U3142 ( .A(n2820), .B(n4021), .ZN(n3285) );
  NOR2_X2 U3143 ( .A1(n2798), .A2(n2515), .ZN(n2782) );
  NAND2_X1 U3144 ( .A1(n2598), .A2(n5033), .ZN(n2786) );
  NAND2_X1 U3145 ( .A1(n2607), .A2(n2608), .ZN(n4763) );
  OR2_X1 U3146 ( .A1(n4699), .A2(n2614), .ZN(n2613) );
  INV_X1 U3147 ( .A(n3483), .ZN(n2619) );
  INV_X1 U31480 ( .A(n5104), .ZN(n2621) );
  AND2_X2 U31490 ( .A1(n4422), .A2(n4425), .ZN(n4534) );
  OAI21_X1 U3150 ( .B1(n3482), .B2(n5104), .A(n3483), .ZN(n3499) );
  INV_X1 U3151 ( .A(n4534), .ZN(n3486) );
  NAND2_X1 U3152 ( .A1(n2622), .A2(n2625), .ZN(n4135) );
  NAND2_X1 U3153 ( .A1(n3675), .A2(n2623), .ZN(n2622) );
  NAND2_X1 U3154 ( .A1(n4980), .A2(n2640), .ZN(n5021) );
  OAI21_X1 U3155 ( .B1(n4746), .B2(n2646), .A(n5108), .ZN(n2645) );
  NOR2_X1 U3156 ( .A1(n4742), .A2(n2647), .ZN(n2646) );
  NAND2_X1 U3157 ( .A1(n3502), .A2(n4428), .ZN(n5185) );
  NAND2_X1 U3158 ( .A1(n4193), .A2(n4507), .ZN(n4194) );
  NOR2_X1 U3159 ( .A1(n4763), .A2(n4764), .ZN(n4762) );
  OAI21_X1 U3160 ( .B1(n3574), .B2(n3573), .A(n4434), .ZN(n3586) );
  NAND2_X1 U3161 ( .A1(n3457), .A2(n3478), .ZN(n4421) );
  NAND2_X1 U3162 ( .A1(n3642), .A2(n4533), .ZN(n3675) );
  NOR2_X1 U3163 ( .A1(n4762), .A2(n4705), .ZN(n4748) );
  AOI21_X1 U3164 ( .B1(n4860), .B2(n4697), .A(n4696), .ZN(n4699) );
  INV_X2 U3165 ( .A(n2786), .ZN(n5036) );
  NAND2_X1 U3166 ( .A1(n4907), .A2(n2652), .ZN(n2651) );
  OAI211_X1 U3167 ( .C1(n3486), .C2(n2658), .A(n2657), .B(n3511), .ZN(n5148)
         );
  INV_X1 U3168 ( .A(n2659), .ZN(n2658) );
  AND2_X1 U3169 ( .A1(n2511), .A2(n3509), .ZN(n2659) );
  NAND2_X1 U3170 ( .A1(n2660), .A2(n3486), .ZN(n3510) );
  OR2_X1 U3171 ( .A1(n4778), .A2(n2666), .ZN(n2663) );
  NAND2_X1 U3172 ( .A1(n4778), .A2(n2498), .ZN(n2662) );
  NAND2_X1 U3173 ( .A1(n4778), .A2(n4728), .ZN(n4760) );
  NAND2_X1 U3174 ( .A1(n3637), .A2(n2517), .ZN(n2668) );
  OR2_X1 U3175 ( .A1(n3669), .A2(n3677), .ZN(n2680) );
  OAI21_X2 U3176 ( .B1(n3561), .B2(n3560), .A(n3563), .ZN(n3571) );
  NAND2_X1 U3177 ( .A1(n4226), .A2(n2681), .ZN(n2684) );
  INV_X1 U3178 ( .A(n2684), .ZN(n5296) );
  NAND2_X1 U3179 ( .A1(n2815), .A2(n2685), .ZN(n2688) );
  OAI21_X1 U3180 ( .B1(n5057), .B2(REG2_REG_2__SCAN_IN), .A(n2689), .ZN(n3411)
         );
  INV_X1 U3181 ( .A(n5057), .ZN(n3417) );
  NAND2_X1 U3182 ( .A1(n2502), .A2(n3357), .ZN(n3423) );
  INV_X1 U3183 ( .A(n2697), .ZN(n3360) );
  NAND2_X1 U3184 ( .A1(n2509), .A2(n2700), .ZN(n2699) );
  NAND2_X1 U3185 ( .A1(n2509), .A2(n3620), .ZN(n3621) );
  NOR2_X1 U3186 ( .A1(n2703), .A2(n3622), .ZN(n2702) );
  INV_X1 U3187 ( .A(n2704), .ZN(n3654) );
  NAND2_X1 U3188 ( .A1(n3534), .A2(n2709), .ZN(n2705) );
  XNOR2_X1 U3189 ( .A(n3532), .B(n3531), .ZN(n3442) );
  NAND2_X1 U3190 ( .A1(n4620), .A2(n4619), .ZN(n4621) );
  INV_X1 U3191 ( .A(n4629), .ZN(n2714) );
  NAND2_X1 U3192 ( .A1(n2714), .A2(n2716), .ZN(n4622) );
  INV_X1 U3193 ( .A(n4406), .ZN(n2738) );
  NAND2_X1 U3194 ( .A1(n2745), .A2(n2746), .ZN(n4112) );
  NAND2_X1 U3195 ( .A1(n4281), .A2(n2533), .ZN(n2745) );
  NAND3_X1 U3196 ( .A1(n2894), .A2(n2893), .A3(n2897), .ZN(n3524) );
  NAND2_X1 U3197 ( .A1(n4309), .A2(n2499), .ZN(n2749) );
  NOR2_X1 U3198 ( .A1(n3025), .A2(IR_REG_13__SCAN_IN), .ZN(n2802) );
  NAND2_X1 U3199 ( .A1(n4329), .A2(n2758), .ZN(n2756) );
  NOR2_X1 U3200 ( .A1(n2798), .A2(n2779), .ZN(n2791) );
  OAI22_X1 U3201 ( .A1(n5110), .A2(n3254), .B1(n2830), .B2(n3478), .ZN(n2862)
         );
  OR2_X2 U3202 ( .A1(n4777), .A2(n4783), .ZN(n4778) );
  AOI21_X2 U3203 ( .B1(n4128), .B2(n4148), .A(n4144), .ZN(n4147) );
  OAI22_X2 U3204 ( .A1(n4121), .A2(n4536), .B1(n4120), .B2(n4583), .ZN(n4144)
         );
  INV_X1 U3205 ( .A(n3069), .ZN(n3072) );
  OR2_X1 U3206 ( .A1(n4363), .A2(n4364), .ZN(n2893) );
  AOI21_X2 U3207 ( .B1(n3593), .B2(n3592), .A(n3591), .ZN(n3637) );
  AND2_X2 U3208 ( .A1(n3462), .A2(n5210), .ZN(n5330) );
  NOR2_X1 U3209 ( .A1(n4340), .A2(n3125), .ZN(n2763) );
  AND3_X1 U32100 ( .A1(n3281), .A2(n3280), .A3(n5282), .ZN(n2764) );
  INV_X1 U32110 ( .A(n4862), .ZN(n4892) );
  AND2_X1 U32120 ( .A1(n5057), .A2(REG2_REG_2__SCAN_IN), .ZN(n2765) );
  AND4_X1 U32130 ( .A1(n3046), .A2(n3045), .A3(n3044), .A4(n3043), .ZN(n5273)
         );
  INV_X1 U32140 ( .A(IR_REG_26__SCAN_IN), .ZN(n2793) );
  INV_X1 U32150 ( .A(n4222), .ZN(n5277) );
  NAND2_X1 U32160 ( .A1(n3073), .A2(n5279), .ZN(n4329) );
  INV_X1 U32170 ( .A(n4198), .ZN(n4199) );
  OR2_X1 U32180 ( .A1(n3402), .A2(n3464), .ZN(n2766) );
  NOR2_X1 U32190 ( .A1(n4847), .A2(n4231), .ZN(n2767) );
  NOR2_X1 U32200 ( .A1(n4383), .A2(n4384), .ZN(n2768) );
  AND2_X1 U32210 ( .A1(n4491), .A2(DATAI_20_), .ZN(n4376) );
  INV_X1 U32220 ( .A(n4376), .ZN(n4881) );
  INV_X1 U32230 ( .A(IR_REG_25__SCAN_IN), .ZN(n2778) );
  NAND2_X1 U32240 ( .A1(n2892), .A2(n3433), .ZN(n4359) );
  AND2_X1 U32250 ( .A1(n3204), .A2(REG3_REG_25__SCAN_IN), .ZN(n3215) );
  INV_X1 U32260 ( .A(n2818), .ZN(n5169) );
  AND2_X1 U32270 ( .A1(n3170), .A2(REG3_REG_22__SCAN_IN), .ZN(n3183) );
  INV_X1 U32280 ( .A(n3107), .ZN(n3128) );
  INV_X1 U32290 ( .A(n3525), .ZN(n2912) );
  AND2_X1 U32300 ( .A1(n3215), .A2(REG3_REG_26__SCAN_IN), .ZN(n3227) );
  INV_X1 U32310 ( .A(n5096), .ZN(n3352) );
  AND2_X1 U32320 ( .A1(n4736), .A2(n3246), .ZN(n4754) );
  INV_X1 U32330 ( .A(n4949), .ZN(n4227) );
  AND2_X1 U32340 ( .A1(n4491), .A2(DATAI_28_), .ZN(n4751) );
  OR2_X1 U32350 ( .A1(n3285), .A2(n3466), .ZN(n5186) );
  INV_X1 U32360 ( .A(n5186), .ZN(n5157) );
  INV_X1 U32370 ( .A(n4251), .ZN(n2941) );
  AND2_X1 U32380 ( .A1(n3183), .A2(REG3_REG_23__SCAN_IN), .ZN(n3185) );
  AND2_X1 U32390 ( .A1(REG3_REG_19__SCAN_IN), .A2(n3128), .ZN(n3143) );
  NAND2_X1 U32400 ( .A1(n3009), .A2(REG3_REG_12__SCAN_IN), .ZN(n3020) );
  NOR2_X1 U32410 ( .A1(n3087), .A2(n4342), .ZN(n3108) );
  OR2_X1 U32420 ( .A1(n2963), .A2(n3770), .ZN(n2979) );
  OR2_X1 U32430 ( .A1(n3291), .A2(n3337), .ZN(n5271) );
  AND2_X1 U32440 ( .A1(n4478), .A2(n4480), .ZN(n4850) );
  INV_X1 U32450 ( .A(n4943), .ZN(n4922) );
  NOR2_X1 U32460 ( .A1(n4147), .A2(n4143), .ZN(n4122) );
  AND2_X1 U32470 ( .A1(n4573), .A2(n3464), .ZN(n5199) );
  INV_X1 U32480 ( .A(n5328), .ZN(n4904) );
  AND2_X1 U32490 ( .A1(n4454), .A2(n4444), .ZN(n4533) );
  OR2_X1 U32500 ( .A1(n5264), .A2(n5202), .ZN(n4974) );
  AND2_X1 U32510 ( .A1(n3258), .A2(n5037), .ZN(n3317) );
  OR3_X1 U32520 ( .A1(n2987), .A2(IR_REG_7__SCAN_IN), .A3(n2986), .ZN(n3003)
         );
  AND2_X1 U32530 ( .A1(n3245), .A2(n3229), .ZN(n4772) );
  NOR2_X1 U32540 ( .A1(n3281), .A2(n4417), .ZN(n3278) );
  AND2_X1 U32550 ( .A1(n4491), .A2(DATAI_22_), .ZN(n4385) );
  NOR2_X1 U32560 ( .A1(n3291), .A2(n3285), .ZN(n4399) );
  AND4_X1 U32570 ( .A1(n3250), .A2(n3249), .A3(n3248), .A4(n3247), .ZN(n4729)
         );
  AND4_X1 U32580 ( .A1(n3209), .A2(n3208), .A3(n3207), .A4(n3206), .ZN(n4823)
         );
  AND4_X1 U32590 ( .A1(n3148), .A2(n3147), .A3(n3146), .A4(n3145), .ZN(n4862)
         );
  AND4_X1 U32600 ( .A1(n3061), .A2(n3060), .A3(n3059), .A4(n3058), .ZN(n4223)
         );
  INV_X1 U32610 ( .A(n5052), .ZN(n3531) );
  INV_X1 U32620 ( .A(n5042), .ZN(n4684) );
  INV_X1 U32630 ( .A(n5194), .ZN(n5108) );
  AND2_X1 U32640 ( .A1(n4460), .A2(n4445), .ZN(n4535) );
  NOR2_X1 U32650 ( .A1(n5330), .A2(n5114), .ZN(n4943) );
  AND2_X1 U32660 ( .A1(n4427), .A2(n4424), .ZN(n4538) );
  NAND2_X1 U32670 ( .A1(n3260), .A2(n3320), .ZN(n4978) );
  INV_X1 U32680 ( .A(n4978), .ZN(n5018) );
  AOI21_X1 U32690 ( .B1(n4262), .B2(n2764), .A(n3310), .ZN(n3311) );
  OR2_X1 U32700 ( .A1(n3287), .A2(n3277), .ZN(n4417) );
  INV_X1 U32710 ( .A(n4729), .ZN(n4768) );
  INV_X1 U32720 ( .A(n4861), .ZN(n4579) );
  INV_X1 U32730 ( .A(n5273), .ZN(n4581) );
  OR2_X1 U32740 ( .A1(n3338), .A2(n4093), .ZN(n4671) );
  OR2_X1 U32750 ( .A1(n3338), .A2(n3337), .ZN(n5089) );
  INV_X1 U32760 ( .A(n4935), .ZN(n4962) );
  NAND2_X1 U32770 ( .A1(n4571), .A2(n3289), .ZN(n5210) );
  INV_X2 U32780 ( .A(n5086), .ZN(n5085) );
  INV_X1 U32790 ( .A(n4592), .ZN(U4043) );
  NOR2_X1 U32800 ( .A1(IR_REG_9__SCAN_IN), .A2(IR_REG_6__SCAN_IN), .ZN(n2772)
         );
  NAND2_X1 U32810 ( .A1(n2497), .A2(REG0_REG_24__SCAN_IN), .ZN(n2790) );
  NAND2_X1 U32820 ( .A1(n2865), .A2(REG1_REG_24__SCAN_IN), .ZN(n2789) );
  INV_X1 U32830 ( .A(n2785), .ZN(n5035) );
  NAND2_X1 U32840 ( .A1(n2898), .A2(REG3_REG_5__SCAN_IN), .ZN(n2929) );
  NAND2_X1 U32850 ( .A1(REG3_REG_7__SCAN_IN), .A2(REG3_REG_6__SCAN_IN), .ZN(
        n2783) );
  NOR2_X1 U32860 ( .A1(n2929), .A2(n2783), .ZN(n2945) );
  NAND2_X1 U32870 ( .A1(n2945), .A2(REG3_REG_8__SCAN_IN), .ZN(n2963) );
  NAND2_X1 U32880 ( .A1(n3108), .A2(REG3_REG_18__SCAN_IN), .ZN(n3107) );
  NOR2_X1 U32890 ( .A1(n3185), .A2(REG3_REG_24__SCAN_IN), .ZN(n2784) );
  NOR2_X1 U32900 ( .A1(n3204), .A2(n2784), .ZN(n4832) );
  NAND2_X1 U32910 ( .A1(n2866), .A2(n4832), .ZN(n2788) );
  NAND2_X1 U32920 ( .A1(n3293), .A2(REG2_REG_24__SCAN_IN), .ZN(n2787) );
  NAND2_X1 U32930 ( .A1(n2801), .A2(n4011), .ZN(n2799) );
  NAND2_X1 U32940 ( .A1(n2799), .A2(IR_REG_31__SCAN_IN), .ZN(n2800) );
  INV_X1 U32950 ( .A(n2803), .ZN(n2804) );
  NOR2_X1 U32960 ( .A1(n2806), .A2(n3093), .ZN(n2807) );
  MUX2_X1 U32970 ( .A(n3093), .B(n2807), .S(IR_REG_21__SCAN_IN), .Z(n2809) );
  NAND2_X1 U32980 ( .A1(n3286), .A2(n5202), .ZN(n3300) );
  NOR2_X1 U32990 ( .A1(n2808), .A2(n3093), .ZN(n2813) );
  MUX2_X1 U33000 ( .A(n3093), .B(n2813), .S(IR_REG_22__SCAN_IN), .Z(n2816) );
  INV_X1 U33010 ( .A(n5040), .ZN(n3470) );
  INV_X1 U33020 ( .A(n5041), .ZN(n2817) );
  INV_X1 U33030 ( .A(n3288), .ZN(n5106) );
  NOR2_X1 U33040 ( .A1(n3300), .A2(n5106), .ZN(n3477) );
  NAND2_X1 U33050 ( .A1(n2872), .A2(DATAI_24_), .ZN(n4822) );
  AOI22_X1 U33060 ( .A1(n4720), .A2(n3237), .B1(n2875), .B2(n4827), .ZN(n4351)
         );
  NAND2_X1 U33070 ( .A1(n2497), .A2(REG0_REG_3__SCAN_IN), .ZN(n2825) );
  INV_X1 U33080 ( .A(REG3_REG_3__SCAN_IN), .ZN(n3944) );
  NAND2_X1 U33090 ( .A1(n2866), .A2(n3944), .ZN(n2824) );
  NAND2_X1 U33100 ( .A1(n2867), .A2(REG2_REG_3__SCAN_IN), .ZN(n2822) );
  NAND2_X1 U33110 ( .A1(n5156), .A2(n2875), .ZN(n2832) );
  NAND2_X1 U33120 ( .A1(n2827), .A2(IR_REG_31__SCAN_IN), .ZN(n2828) );
  NAND2_X1 U33130 ( .A1(n2828), .A2(n3977), .ZN(n2853) );
  OR2_X1 U33140 ( .A1(n2828), .A2(n3977), .ZN(n2829) );
  MUX2_X1 U33150 ( .A(n5056), .B(DATAI_3_), .S(n2872), .Z(n4218) );
  NAND2_X1 U33160 ( .A1(n4218), .A2(n2956), .ZN(n2831) );
  NAND2_X1 U33170 ( .A1(n2832), .A2(n2831), .ZN(n2833) );
  XNOR2_X1 U33180 ( .A(n2833), .B(n3464), .ZN(n2890) );
  AOI22_X1 U33190 ( .A1(n5156), .A2(n3237), .B1(n2875), .B2(n4218), .ZN(n2889)
         );
  INV_X1 U33200 ( .A(n2889), .ZN(n2834) );
  NAND2_X1 U33210 ( .A1(n2496), .A2(REG0_REG_2__SCAN_IN), .ZN(n2837) );
  NAND2_X1 U33220 ( .A1(n2866), .A2(REG3_REG_2__SCAN_IN), .ZN(n2836) );
  NAND2_X1 U33230 ( .A1(n2865), .A2(REG1_REG_2__SCAN_IN), .ZN(n2835) );
  AND3_X1 U33240 ( .A1(n2837), .A2(n2836), .A3(n2835), .ZN(n2839) );
  NAND2_X1 U33250 ( .A1(n2867), .A2(REG2_REG_2__SCAN_IN), .ZN(n2838) );
  NAND2_X2 U33260 ( .A1(n2839), .A2(n2838), .ZN(n4591) );
  XNOR2_X2 U33270 ( .A(n2840), .B(IR_REG_2__SCAN_IN), .ZN(n5057) );
  OAI22_X1 U33280 ( .A1(n3508), .A2(n3254), .B1(n2830), .B2(n3507), .ZN(n2841)
         );
  XNOR2_X1 U33290 ( .A(n2841), .B(n3464), .ZN(n2887) );
  INV_X1 U33300 ( .A(n2887), .ZN(n2845) );
  OR2_X1 U33310 ( .A1(n3508), .A2(n3251), .ZN(n2843) );
  NAND2_X1 U33320 ( .A1(n3493), .A2(n2875), .ZN(n2842) );
  NAND2_X1 U33330 ( .A1(n2843), .A2(n2842), .ZN(n2886) );
  INV_X1 U33340 ( .A(n2886), .ZN(n2844) );
  NAND2_X1 U33350 ( .A1(n2845), .A2(n2844), .ZN(n3433) );
  NAND2_X1 U33360 ( .A1(n2496), .A2(REG0_REG_4__SCAN_IN), .ZN(n2852) );
  NAND2_X1 U33370 ( .A1(n2867), .A2(REG2_REG_4__SCAN_IN), .ZN(n2851) );
  INV_X1 U33380 ( .A(n2898), .ZN(n2847) );
  INV_X1 U33390 ( .A(REG3_REG_4__SCAN_IN), .ZN(n4367) );
  NAND2_X1 U33400 ( .A1(n4367), .A2(n3944), .ZN(n2846) );
  NAND2_X1 U33410 ( .A1(n2847), .A2(n2846), .ZN(n5177) );
  INV_X1 U33420 ( .A(n5177), .ZN(n2848) );
  NAND2_X1 U33430 ( .A1(n2866), .A2(n2848), .ZN(n2850) );
  NAND2_X1 U33440 ( .A1(n2865), .A2(REG1_REG_4__SCAN_IN), .ZN(n2849) );
  NAND2_X1 U33450 ( .A1(n2853), .A2(IR_REG_31__SCAN_IN), .ZN(n2854) );
  XNOR2_X1 U33460 ( .A(n2854), .B(IR_REG_4__SCAN_IN), .ZN(n5096) );
  XNOR2_X1 U33470 ( .A(n2855), .B(n3464), .ZN(n2896) );
  OR2_X1 U33480 ( .A1(n5187), .A2(n3251), .ZN(n2857) );
  NAND2_X1 U33490 ( .A1(n5158), .A2(n2875), .ZN(n2856) );
  NAND2_X1 U33500 ( .A1(n2857), .A2(n2856), .ZN(n2895) );
  XNOR2_X1 U33510 ( .A(n2896), .B(n2895), .ZN(n4364) );
  NOR2_X1 U33520 ( .A1(n4359), .A2(n4364), .ZN(n2888) );
  NAND2_X1 U3353 ( .A1(n2867), .A2(REG2_REG_1__SCAN_IN), .ZN(n2860) );
  NAND2_X1 U33540 ( .A1(n2978), .A2(REG0_REG_1__SCAN_IN), .ZN(n2859) );
  NAND2_X1 U3355 ( .A1(n2865), .A2(REG1_REG_1__SCAN_IN), .ZN(n2858) );
  INV_X1 U3356 ( .A(n3347), .ZN(n3346) );
  XNOR2_X1 U3357 ( .A(n2862), .B(n3252), .ZN(n2882) );
  OR2_X1 U3358 ( .A1(n5110), .A2(n3251), .ZN(n2864) );
  NAND2_X1 U3359 ( .A1(n4304), .A2(n2875), .ZN(n2863) );
  NAND2_X1 U3360 ( .A1(n2864), .A2(n2863), .ZN(n2883) );
  XNOR2_X1 U3361 ( .A(n2882), .B(n2883), .ZN(n4302) );
  NAND2_X1 U3362 ( .A1(n2865), .A2(REG1_REG_0__SCAN_IN), .ZN(n2871) );
  NAND2_X1 U3363 ( .A1(n2497), .A2(REG0_REG_0__SCAN_IN), .ZN(n2870) );
  NAND2_X1 U3364 ( .A1(n2866), .A2(REG3_REG_0__SCAN_IN), .ZN(n2869) );
  NAND2_X1 U3365 ( .A1(n2867), .A2(REG2_REG_0__SCAN_IN), .ZN(n2868) );
  NAND2_X1 U3366 ( .A1(n4593), .A2(n2875), .ZN(n2874) );
  NAND2_X1 U3367 ( .A1(n4419), .A2(n2956), .ZN(n2873) );
  NAND2_X1 U3368 ( .A1(n2874), .A2(n2873), .ZN(n3402) );
  NAND2_X1 U3369 ( .A1(n4593), .A2(n3237), .ZN(n2877) );
  NAND2_X1 U3370 ( .A1(n4419), .A2(n2875), .ZN(n2876) );
  NAND2_X1 U3371 ( .A1(n2877), .A2(n2876), .ZN(n3401) );
  NAND2_X1 U3372 ( .A1(n3401), .A2(n3402), .ZN(n2880) );
  NAND2_X1 U3373 ( .A1(IR_REG_0__SCAN_IN), .A2(REG1_REG_0__SCAN_IN), .ZN(n3340) );
  OR2_X1 U3374 ( .A1(n2878), .A2(n3340), .ZN(n2879) );
  NAND2_X1 U3375 ( .A1(n2880), .A2(n2879), .ZN(n3403) );
  INV_X1 U3376 ( .A(n3403), .ZN(n2881) );
  NAND2_X1 U3377 ( .A1(n2766), .A2(n2881), .ZN(n4301) );
  NAND2_X1 U3378 ( .A1(n4302), .A2(n4301), .ZN(n4300) );
  INV_X1 U3379 ( .A(n2882), .ZN(n2884) );
  NAND2_X1 U3380 ( .A1(n2884), .A2(n2883), .ZN(n2885) );
  NAND2_X1 U3381 ( .A1(n4300), .A2(n2885), .ZN(n3452) );
  XNOR2_X1 U3382 ( .A(n2887), .B(n2886), .ZN(n3453) );
  NAND2_X1 U3383 ( .A1(n2888), .A2(n4361), .ZN(n2894) );
  XNOR2_X1 U3384 ( .A(n2890), .B(n2889), .ZN(n3435) );
  INV_X1 U3385 ( .A(n3435), .ZN(n2891) );
  NAND2_X1 U3386 ( .A1(n2892), .A2(n2891), .ZN(n4363) );
  NAND2_X1 U3387 ( .A1(n2896), .A2(n2895), .ZN(n2897) );
  NAND2_X1 U3388 ( .A1(n2865), .A2(REG1_REG_5__SCAN_IN), .ZN(n2903) );
  NAND2_X1 U3389 ( .A1(n2497), .A2(REG0_REG_5__SCAN_IN), .ZN(n2902) );
  OAI21_X1 U3390 ( .B1(n2898), .B2(REG3_REG_5__SCAN_IN), .A(n2929), .ZN(n5211)
         );
  INV_X1 U3391 ( .A(n5211), .ZN(n2899) );
  NAND2_X1 U3392 ( .A1(n2866), .A2(n2899), .ZN(n2901) );
  NAND2_X1 U3393 ( .A1(n3293), .A2(REG2_REG_5__SCAN_IN), .ZN(n2900) );
  NAND4_X1 U3394 ( .A1(n2903), .A2(n2902), .A3(n2901), .A4(n2900), .ZN(n5155)
         );
  NAND2_X1 U3395 ( .A1(n5155), .A2(n2875), .ZN(n2910) );
  AND3_X1 U3396 ( .A1(n3980), .A2(n3977), .A3(n3780), .ZN(n2904) );
  INV_X1 U3397 ( .A(n2937), .ZN(n2908) );
  NAND2_X1 U3398 ( .A1(n2905), .A2(IR_REG_31__SCAN_IN), .ZN(n2906) );
  MUX2_X1 U3399 ( .A(IR_REG_31__SCAN_IN), .B(n2906), .S(IR_REG_5__SCAN_IN), 
        .Z(n2907) );
  MUX2_X1 U3400 ( .A(n5055), .B(DATAI_5_), .S(n4491), .Z(n5192) );
  NAND2_X1 U3401 ( .A1(n5192), .A2(n2956), .ZN(n2909) );
  NAND2_X1 U3402 ( .A1(n2910), .A2(n2909), .ZN(n2911) );
  XNOR2_X1 U3403 ( .A(n2911), .B(n3252), .ZN(n2914) );
  AOI22_X1 U3404 ( .A1(n5155), .A2(n3237), .B1(n2875), .B2(n5192), .ZN(n2913)
         );
  XNOR2_X1 U3405 ( .A(n2914), .B(n2913), .ZN(n3525) );
  NAND2_X1 U3406 ( .A1(n2914), .A2(n2913), .ZN(n2915) );
  NAND2_X1 U3407 ( .A1(n2497), .A2(REG0_REG_6__SCAN_IN), .ZN(n2919) );
  NAND2_X1 U3408 ( .A1(n2865), .A2(REG1_REG_6__SCAN_IN), .ZN(n2918) );
  XNOR2_X1 U3409 ( .A(n2929), .B(REG3_REG_6__SCAN_IN), .ZN(n3550) );
  NAND2_X1 U3410 ( .A1(n2866), .A2(n3550), .ZN(n2917) );
  NAND2_X1 U3411 ( .A1(n3293), .A2(REG2_REG_6__SCAN_IN), .ZN(n2916) );
  NAND4_X1 U3412 ( .A1(n2919), .A2(n2918), .A3(n2917), .A4(n2916), .ZN(n4589)
         );
  NAND2_X1 U3413 ( .A1(n4589), .A2(n2875), .ZN(n2922) );
  OR2_X1 U3414 ( .A1(n2937), .A2(n3093), .ZN(n2920) );
  XNOR2_X1 U3415 ( .A(n2920), .B(IR_REG_6__SCAN_IN), .ZN(n5054) );
  MUX2_X1 U3416 ( .A(n5054), .B(DATAI_6_), .S(n4491), .Z(n3562) );
  NAND2_X1 U3417 ( .A1(n3562), .A2(n2956), .ZN(n2921) );
  NAND2_X1 U3418 ( .A1(n2922), .A2(n2921), .ZN(n2923) );
  XNOR2_X1 U3419 ( .A(n2923), .B(n3464), .ZN(n2924) );
  AOI22_X1 U3420 ( .A1(n4589), .A2(n3237), .B1(n2875), .B2(n3562), .ZN(n2925)
         );
  XNOR2_X1 U3421 ( .A(n2924), .B(n2925), .ZN(n3546) );
  INV_X1 U3422 ( .A(n2924), .ZN(n2926) );
  NAND2_X1 U3423 ( .A1(n2926), .A2(n2925), .ZN(n2927) );
  NAND2_X1 U3424 ( .A1(n2928), .A2(n2927), .ZN(n4252) );
  NAND2_X1 U3425 ( .A1(n2497), .A2(REG0_REG_7__SCAN_IN), .ZN(n2936) );
  NAND2_X1 U3426 ( .A1(n2865), .A2(REG1_REG_7__SCAN_IN), .ZN(n2935) );
  INV_X1 U3427 ( .A(n2929), .ZN(n2930) );
  AOI21_X1 U3428 ( .B1(n2930), .B2(REG3_REG_6__SCAN_IN), .A(
        REG3_REG_7__SCAN_IN), .ZN(n2931) );
  OR2_X1 U3429 ( .A1(n2931), .A2(n2945), .ZN(n4256) );
  INV_X1 U3430 ( .A(n4256), .ZN(n2932) );
  NAND2_X1 U3431 ( .A1(n2866), .A2(n2932), .ZN(n2934) );
  NAND2_X1 U3432 ( .A1(n3293), .A2(REG2_REG_7__SCAN_IN), .ZN(n2933) );
  NAND2_X1 U3433 ( .A1(n2937), .A2(n3787), .ZN(n2987) );
  NAND2_X1 U3434 ( .A1(n2987), .A2(IR_REG_31__SCAN_IN), .ZN(n2952) );
  MUX2_X1 U3435 ( .A(n5053), .B(DATAI_7_), .S(n4491), .Z(n4255) );
  INV_X1 U3436 ( .A(n4255), .ZN(n3559) );
  OAI22_X1 U3437 ( .A1(n3555), .A2(n3254), .B1(n2830), .B2(n3559), .ZN(n2938)
         );
  XNOR2_X1 U3438 ( .A(n2938), .B(n3464), .ZN(n2943) );
  OR2_X1 U3439 ( .A1(n3555), .A2(n3251), .ZN(n2940) );
  NAND2_X1 U3440 ( .A1(n4255), .A2(n2875), .ZN(n2939) );
  NAND2_X1 U3441 ( .A1(n2940), .A2(n2939), .ZN(n2942) );
  XNOR2_X1 U3442 ( .A(n2943), .B(n2942), .ZN(n4251) );
  NAND2_X1 U3443 ( .A1(n2943), .A2(n2942), .ZN(n2944) );
  NAND2_X1 U3444 ( .A1(n2865), .A2(REG1_REG_8__SCAN_IN), .ZN(n2950) );
  NAND2_X1 U3445 ( .A1(n2497), .A2(REG0_REG_8__SCAN_IN), .ZN(n2949) );
  OR2_X1 U3446 ( .A1(n2945), .A2(REG3_REG_8__SCAN_IN), .ZN(n2946) );
  AND2_X1 U3447 ( .A1(n2963), .A2(n2946), .ZN(n3607) );
  NAND2_X1 U3448 ( .A1(n2866), .A2(n3607), .ZN(n2948) );
  NAND2_X1 U3449 ( .A1(n3293), .A2(REG2_REG_8__SCAN_IN), .ZN(n2947) );
  NAND4_X1 U3450 ( .A1(n2950), .A2(n2949), .A3(n2948), .A4(n2947), .ZN(n4587)
         );
  NAND2_X1 U3451 ( .A1(n4587), .A2(n2875), .ZN(n2958) );
  INV_X1 U3452 ( .A(IR_REG_7__SCAN_IN), .ZN(n2951) );
  NAND2_X1 U3453 ( .A1(n2952), .A2(n2951), .ZN(n2953) );
  NAND2_X1 U3454 ( .A1(n2953), .A2(IR_REG_31__SCAN_IN), .ZN(n2954) );
  NAND2_X1 U3455 ( .A1(n2954), .A2(n2985), .ZN(n2969) );
  OR2_X1 U3456 ( .A1(n2954), .A2(n2985), .ZN(n2955) );
  MUX2_X1 U3457 ( .A(n5052), .B(DATAI_8_), .S(n2872), .Z(n3605) );
  NAND2_X1 U34580 ( .A1(n3605), .A2(n2956), .ZN(n2957) );
  NAND2_X1 U34590 ( .A1(n2958), .A2(n2957), .ZN(n2959) );
  XNOR2_X1 U3460 ( .A(n2959), .B(n3464), .ZN(n2960) );
  AOI22_X1 U3461 ( .A1(n4587), .A2(n3237), .B1(n2875), .B2(n3605), .ZN(n2961)
         );
  XNOR2_X1 U3462 ( .A(n2960), .B(n2961), .ZN(n3604) );
  INV_X1 U3463 ( .A(n2960), .ZN(n2962) );
  NAND2_X1 U3464 ( .A1(n2865), .A2(REG1_REG_9__SCAN_IN), .ZN(n2968) );
  NAND2_X1 U3465 ( .A1(n2497), .A2(REG0_REG_9__SCAN_IN), .ZN(n2967) );
  NAND2_X1 U3466 ( .A1(n2963), .A2(n3770), .ZN(n2964) );
  AND2_X1 U34670 ( .A1(n2979), .A2(n2964), .ZN(n3631) );
  NAND2_X1 U3468 ( .A1(n2866), .A2(n3631), .ZN(n2966) );
  NAND2_X1 U34690 ( .A1(n3293), .A2(REG2_REG_9__SCAN_IN), .ZN(n2965) );
  NAND2_X1 U3470 ( .A1(n2969), .A2(IR_REG_31__SCAN_IN), .ZN(n2970) );
  XNOR2_X1 U34710 ( .A(n2970), .B(IR_REG_9__SCAN_IN), .ZN(n5051) );
  INV_X1 U3472 ( .A(n5051), .ZN(n3614) );
  INV_X1 U34730 ( .A(DATAI_9_), .ZN(n3921) );
  MUX2_X1 U3474 ( .A(n3614), .B(n3921), .S(n2872), .Z(n3640) );
  OAI22_X1 U34750 ( .A1(n3643), .A2(n3254), .B1(n2830), .B2(n3640), .ZN(n2971)
         );
  XNOR2_X1 U3476 ( .A(n2971), .B(n3252), .ZN(n2976) );
  OR2_X1 U34770 ( .A1(n3643), .A2(n3251), .ZN(n2973) );
  OR2_X1 U3478 ( .A1(n3640), .A2(n3254), .ZN(n2972) );
  NAND2_X1 U34790 ( .A1(n2973), .A2(n2972), .ZN(n2974) );
  XNOR2_X1 U3480 ( .A(n2976), .B(n2974), .ZN(n3628) );
  INV_X1 U34810 ( .A(n2974), .ZN(n2975) );
  AND2_X1 U3482 ( .A1(n2976), .A2(n2975), .ZN(n2977) );
  NAND2_X1 U34830 ( .A1(n2865), .A2(REG1_REG_10__SCAN_IN), .ZN(n2984) );
  NAND2_X1 U3484 ( .A1(n2496), .A2(REG0_REG_10__SCAN_IN), .ZN(n2983) );
  AND2_X1 U34850 ( .A1(n2979), .A2(n3746), .ZN(n2980) );
  NOR2_X1 U3486 ( .A1(n2996), .A2(n2980), .ZN(n3649) );
  NAND2_X1 U34870 ( .A1(n2866), .A2(n3649), .ZN(n2982) );
  NAND2_X1 U3488 ( .A1(n3293), .A2(REG2_REG_10__SCAN_IN), .ZN(n2981) );
  NAND2_X1 U34890 ( .A1(n2985), .A2(n3988), .ZN(n2986) );
  NAND2_X1 U3490 ( .A1(n3003), .A2(IR_REG_31__SCAN_IN), .ZN(n2988) );
  XNOR2_X1 U34910 ( .A(n2988), .B(IR_REG_10__SCAN_IN), .ZN(n5050) );
  MUX2_X1 U3492 ( .A(n5050), .B(DATAI_10_), .S(n4491), .Z(n4282) );
  OAI22_X1 U34930 ( .A1(n3677), .A2(n3254), .B1(n2830), .B2(n3669), .ZN(n2989)
         );
  XNOR2_X1 U3494 ( .A(n2989), .B(n3252), .ZN(n2992) );
  OR2_X1 U34950 ( .A1(n3677), .A2(n3251), .ZN(n2991) );
  NAND2_X1 U3496 ( .A1(n4282), .A2(n2875), .ZN(n2990) );
  NAND2_X1 U34970 ( .A1(n2991), .A2(n2990), .ZN(n2993) );
  XNOR2_X1 U3498 ( .A(n2992), .B(n2993), .ZN(n4280) );
  INV_X1 U34990 ( .A(n2992), .ZN(n2994) );
  NAND2_X1 U3500 ( .A1(n2994), .A2(n2993), .ZN(n2995) );
  NAND2_X1 U35010 ( .A1(n2865), .A2(REG1_REG_11__SCAN_IN), .ZN(n3002) );
  NAND2_X1 U3502 ( .A1(n2496), .A2(REG0_REG_11__SCAN_IN), .ZN(n3001) );
  NOR2_X1 U35030 ( .A1(n2996), .A2(REG3_REG_11__SCAN_IN), .ZN(n2997) );
  OR2_X1 U3504 ( .A1(n3009), .A2(n2997), .ZN(n3689) );
  INV_X1 U35050 ( .A(n3689), .ZN(n2998) );
  NAND2_X1 U35060 ( .A1(n2866), .A2(n2998), .ZN(n3000) );
  NAND2_X1 U35070 ( .A1(n3293), .A2(REG2_REG_11__SCAN_IN), .ZN(n2999) );
  OAI21_X1 U35080 ( .B1(n3003), .B2(IR_REG_10__SCAN_IN), .A(IR_REG_31__SCAN_IN), .ZN(n3004) );
  NAND2_X1 U35090 ( .A1(n3004), .A2(n3795), .ZN(n3015) );
  OR2_X1 U35100 ( .A1(n3004), .A2(n3795), .ZN(n3005) );
  MUX2_X1 U35110 ( .A(n5049), .B(DATAI_11_), .S(n2872), .Z(n3687) );
  OAI22_X1 U35120 ( .A1(n4102), .A2(n3254), .B1(n2830), .B2(n4101), .ZN(n3006)
         );
  XNOR2_X1 U35130 ( .A(n3006), .B(n3464), .ZN(n3683) );
  OR2_X1 U35140 ( .A1(n4102), .A2(n3251), .ZN(n3008) );
  NAND2_X1 U35150 ( .A1(n3687), .A2(n2875), .ZN(n3007) );
  NAND2_X1 U35160 ( .A1(n3008), .A2(n3007), .ZN(n3684) );
  NAND2_X1 U35170 ( .A1(n2497), .A2(REG0_REG_12__SCAN_IN), .ZN(n3014) );
  NAND2_X1 U35180 ( .A1(n2865), .A2(REG1_REG_12__SCAN_IN), .ZN(n3013) );
  OR2_X1 U35190 ( .A1(n3009), .A2(REG3_REG_12__SCAN_IN), .ZN(n3010) );
  AND2_X1 U35200 ( .A1(n3010), .A2(n3020), .ZN(n4116) );
  NAND2_X1 U35210 ( .A1(n2866), .A2(n4116), .ZN(n3012) );
  NAND2_X1 U35220 ( .A1(n3293), .A2(REG2_REG_12__SCAN_IN), .ZN(n3011) );
  NAND2_X1 U35230 ( .A1(n3015), .A2(IR_REG_31__SCAN_IN), .ZN(n3016) );
  XNOR2_X1 U35240 ( .A(n3016), .B(IR_REG_12__SCAN_IN), .ZN(n5048) );
  MUX2_X1 U35250 ( .A(n5048), .B(DATAI_12_), .S(n4491), .Z(n4120) );
  INV_X1 U35260 ( .A(n4120), .ZN(n4097) );
  OAI22_X1 U35270 ( .A1(n4139), .A2(n3254), .B1(n2830), .B2(n4097), .ZN(n3017)
         );
  XNOR2_X1 U35280 ( .A(n3017), .B(n3252), .ZN(n3030) );
  OR2_X1 U35290 ( .A1(n4139), .A2(n3251), .ZN(n3019) );
  NAND2_X1 U35300 ( .A1(n4120), .A2(n2875), .ZN(n3018) );
  AND2_X1 U35310 ( .A1(n3019), .A2(n3018), .ZN(n3031) );
  NAND2_X1 U35320 ( .A1(n3030), .A2(n3031), .ZN(n4111) );
  NAND2_X1 U35330 ( .A1(n2865), .A2(REG1_REG_13__SCAN_IN), .ZN(n3024) );
  NAND2_X1 U35340 ( .A1(n2496), .A2(REG0_REG_13__SCAN_IN), .ZN(n3023) );
  AOI21_X1 U35350 ( .B1(n3020), .B2(n4164), .A(n3041), .ZN(n4151) );
  NAND2_X1 U35360 ( .A1(n2866), .A2(n4151), .ZN(n3022) );
  NAND2_X1 U35370 ( .A1(n3293), .A2(REG2_REG_13__SCAN_IN), .ZN(n3021) );
  NAND2_X1 U35380 ( .A1(n3025), .A2(IR_REG_31__SCAN_IN), .ZN(n3026) );
  XNOR2_X1 U35390 ( .A(n3026), .B(n2754), .ZN(n4614) );
  INV_X1 U35400 ( .A(DATAI_13_), .ZN(n3719) );
  MUX2_X1 U35410 ( .A(n4614), .B(n3719), .S(n4491), .Z(n4148) );
  OAI22_X1 U35420 ( .A1(n4128), .A2(n3254), .B1(n2830), .B2(n4148), .ZN(n3027)
         );
  XNOR2_X1 U35430 ( .A(n3027), .B(n3464), .ZN(n3036) );
  OR2_X1 U35440 ( .A1(n4128), .A2(n3251), .ZN(n3029) );
  OR2_X1 U35450 ( .A1(n4148), .A2(n3254), .ZN(n3028) );
  NAND2_X1 U35460 ( .A1(n3029), .A2(n3028), .ZN(n3037) );
  XNOR2_X1 U35470 ( .A(n3036), .B(n3037), .ZN(n4162) );
  INV_X1 U35480 ( .A(n4162), .ZN(n3034) );
  INV_X1 U35490 ( .A(n3030), .ZN(n3033) );
  INV_X1 U35500 ( .A(n3031), .ZN(n3032) );
  NAND2_X1 U35510 ( .A1(n3033), .A2(n3032), .ZN(n4157) );
  AND2_X1 U35520 ( .A1(n3034), .A2(n4157), .ZN(n3035) );
  INV_X1 U35530 ( .A(n3036), .ZN(n3039) );
  INV_X1 U35540 ( .A(n3037), .ZN(n3038) );
  NAND2_X1 U35550 ( .A1(n3039), .A2(n3038), .ZN(n3040) );
  NAND2_X1 U35560 ( .A1(n2497), .A2(REG0_REG_14__SCAN_IN), .ZN(n3046) );
  NAND2_X1 U35570 ( .A1(n3293), .A2(REG2_REG_14__SCAN_IN), .ZN(n3045) );
  OAI21_X1 U35580 ( .B1(n3041), .B2(REG3_REG_14__SCAN_IN), .A(n3054), .ZN(
        n4186) );
  INV_X1 U35590 ( .A(n4186), .ZN(n3042) );
  NAND2_X1 U35600 ( .A1(n2866), .A2(n3042), .ZN(n3044) );
  NAND2_X1 U35610 ( .A1(n2865), .A2(REG1_REG_14__SCAN_IN), .ZN(n3043) );
  XNOR2_X1 U35620 ( .A(n3047), .B(IR_REG_14__SCAN_IN), .ZN(n5046) );
  MUX2_X1 U35630 ( .A(n5046), .B(DATAI_14_), .S(n4491), .Z(n4198) );
  OAI22_X1 U35640 ( .A1(n5273), .A2(n3254), .B1(n2830), .B2(n4199), .ZN(n3048)
         );
  XNOR2_X1 U35650 ( .A(n3048), .B(n3252), .ZN(n3053) );
  OR2_X1 U35660 ( .A1(n5273), .A2(n3251), .ZN(n3050) );
  NAND2_X1 U35670 ( .A1(n4198), .A2(n2875), .ZN(n3049) );
  NAND2_X1 U35680 ( .A1(n3050), .A2(n3049), .ZN(n3051) );
  XNOR2_X1 U35690 ( .A(n3053), .B(n3051), .ZN(n4182) );
  INV_X1 U35700 ( .A(n3051), .ZN(n3052) );
  NAND2_X1 U35710 ( .A1(n2865), .A2(REG1_REG_15__SCAN_IN), .ZN(n3061) );
  NAND2_X1 U35720 ( .A1(n2496), .A2(REG0_REG_15__SCAN_IN), .ZN(n3060) );
  NAND2_X1 U35730 ( .A1(n3054), .A2(n4639), .ZN(n3056) );
  INV_X1 U35740 ( .A(n3074), .ZN(n3055) );
  NAND2_X1 U35750 ( .A1(n3056), .A2(n3055), .ZN(n5286) );
  INV_X1 U35760 ( .A(n5286), .ZN(n3057) );
  NAND2_X1 U35770 ( .A1(n2866), .A2(n3057), .ZN(n3059) );
  NAND2_X1 U35780 ( .A1(n3293), .A2(REG2_REG_15__SCAN_IN), .ZN(n3058) );
  NAND2_X1 U35790 ( .A1(n3062), .A2(IR_REG_31__SCAN_IN), .ZN(n3064) );
  INV_X1 U35800 ( .A(n3064), .ZN(n3063) );
  NAND2_X1 U35810 ( .A1(n3063), .A2(IR_REG_15__SCAN_IN), .ZN(n3065) );
  INV_X1 U3582 ( .A(IR_REG_15__SCAN_IN), .ZN(n3997) );
  NAND2_X1 U3583 ( .A1(n3064), .A2(n3997), .ZN(n3080) );
  INV_X1 U3584 ( .A(DATAI_15_), .ZN(n3905) );
  MUX2_X1 U3585 ( .A(n4648), .B(n3905), .S(n4491), .Z(n4222) );
  OAI22_X1 U3586 ( .A1(n4223), .A2(n3254), .B1(n2830), .B2(n4222), .ZN(n3066)
         );
  XNOR2_X1 U3587 ( .A(n3066), .B(n3252), .ZN(n3070) );
  OR2_X1 U3588 ( .A1(n4223), .A2(n3251), .ZN(n3068) );
  OR2_X1 U3589 ( .A1(n4222), .A2(n3254), .ZN(n3067) );
  NAND2_X1 U3590 ( .A1(n3068), .A2(n3067), .ZN(n5280) );
  NAND2_X1 U3591 ( .A1(n5278), .A2(n5280), .ZN(n3073) );
  NAND2_X1 U3592 ( .A1(n2865), .A2(REG1_REG_16__SCAN_IN), .ZN(n3079) );
  NAND2_X1 U3593 ( .A1(n2497), .A2(REG0_REG_16__SCAN_IN), .ZN(n3078) );
  OAI21_X1 U3594 ( .B1(REG3_REG_16__SCAN_IN), .B2(n3074), .A(n3087), .ZN(n4958) );
  INV_X1 U3595 ( .A(n4958), .ZN(n3075) );
  NAND2_X1 U3596 ( .A1(n2866), .A2(n3075), .ZN(n3077) );
  NAND2_X1 U3597 ( .A1(n3293), .A2(REG2_REG_16__SCAN_IN), .ZN(n3076) );
  NAND4_X1 U3598 ( .A1(n3079), .A2(n3078), .A3(n3077), .A4(n3076), .ZN(n4929)
         );
  NAND2_X1 U3599 ( .A1(n4929), .A2(n2875), .ZN(n3083) );
  NAND2_X1 U3600 ( .A1(n3080), .A2(IR_REG_31__SCAN_IN), .ZN(n3081) );
  XNOR2_X1 U3601 ( .A(n3081), .B(IR_REG_16__SCAN_IN), .ZN(n5044) );
  INV_X1 U3602 ( .A(n5044), .ZN(n4660) );
  INV_X1 U3603 ( .A(DATAI_16_), .ZN(n3903) );
  MUX2_X1 U3604 ( .A(n4660), .B(n3903), .S(n4491), .Z(n4953) );
  OR2_X1 U3605 ( .A1(n4953), .A2(n2830), .ZN(n3082) );
  NAND2_X1 U3606 ( .A1(n3083), .A2(n3082), .ZN(n3084) );
  XNOR2_X1 U3607 ( .A(n3084), .B(n3464), .ZN(n4330) );
  NAND2_X1 U3608 ( .A1(n4929), .A2(n3237), .ZN(n3086) );
  OR2_X1 U3609 ( .A1(n4953), .A2(n3254), .ZN(n3085) );
  NAND2_X1 U3610 ( .A1(n3086), .A2(n3085), .ZN(n4331) );
  NAND2_X1 U3611 ( .A1(n2865), .A2(REG1_REG_17__SCAN_IN), .ZN(n3091) );
  NAND2_X1 U3612 ( .A1(n2496), .A2(REG0_REG_17__SCAN_IN), .ZN(n3090) );
  AOI21_X1 U3613 ( .B1(n4342), .B2(n3087), .A(n3108), .ZN(n4939) );
  NAND2_X1 U3614 ( .A1(n2866), .A2(n4939), .ZN(n3089) );
  NAND2_X1 U3615 ( .A1(n3293), .A2(REG2_REG_17__SCAN_IN), .ZN(n3088) );
  NAND4_X1 U3616 ( .A1(n3091), .A2(n3090), .A3(n3089), .A4(n3088), .ZN(n4949)
         );
  NAND2_X1 U3617 ( .A1(n4949), .A2(n2875), .ZN(n3098) );
  NOR2_X1 U3618 ( .A1(n3092), .A2(n3093), .ZN(n3094) );
  MUX2_X1 U3619 ( .A(n3093), .B(n3094), .S(IR_REG_17__SCAN_IN), .Z(n3095) );
  INV_X1 U3620 ( .A(n3095), .ZN(n3096) );
  INV_X1 U3621 ( .A(DATAI_17_), .ZN(n3904) );
  MUX2_X1 U3622 ( .A(n4679), .B(n3904), .S(n4491), .Z(n4936) );
  OR2_X1 U3623 ( .A1(n4936), .A2(n2830), .ZN(n3097) );
  NAND2_X1 U3624 ( .A1(n3098), .A2(n3097), .ZN(n3099) );
  XNOR2_X1 U3625 ( .A(n3099), .B(n3252), .ZN(n3102) );
  NAND2_X1 U3626 ( .A1(n4949), .A2(n3237), .ZN(n3101) );
  OR2_X1 U3627 ( .A1(n4936), .A2(n3254), .ZN(n3100) );
  AND2_X1 U3628 ( .A1(n3101), .A2(n3100), .ZN(n3103) );
  NAND2_X1 U3629 ( .A1(n3102), .A2(n3103), .ZN(n4392) );
  INV_X1 U3630 ( .A(n3102), .ZN(n3105) );
  INV_X1 U3631 ( .A(n3103), .ZN(n3104) );
  NAND2_X1 U3632 ( .A1(n3105), .A2(n3104), .ZN(n3106) );
  NAND2_X1 U3633 ( .A1(n4392), .A2(n3106), .ZN(n4340) );
  NAND2_X1 U3634 ( .A1(n2865), .A2(REG1_REG_18__SCAN_IN), .ZN(n3112) );
  NAND2_X1 U3635 ( .A1(n2497), .A2(REG0_REG_18__SCAN_IN), .ZN(n3111) );
  OAI21_X1 U3636 ( .B1(REG3_REG_18__SCAN_IN), .B2(n3108), .A(n3107), .ZN(n4401) );
  INV_X1 U3637 ( .A(n4401), .ZN(n4920) );
  NAND2_X1 U3638 ( .A1(n2866), .A2(n4920), .ZN(n3110) );
  NAND2_X1 U3639 ( .A1(n3293), .A2(REG2_REG_18__SCAN_IN), .ZN(n3109) );
  NAND4_X1 U3640 ( .A1(n3112), .A2(n3111), .A3(n3110), .A4(n3109), .ZN(n4928)
         );
  NAND2_X1 U3641 ( .A1(n4928), .A2(n2875), .ZN(n3116) );
  NAND2_X1 U3642 ( .A1(n3113), .A2(IR_REG_31__SCAN_IN), .ZN(n3114) );
  XNOR2_X1 U3643 ( .A(n3114), .B(IR_REG_18__SCAN_IN), .ZN(n5042) );
  INV_X1 U3644 ( .A(DATAI_18_), .ZN(n3910) );
  MUX2_X1 U3645 ( .A(n4684), .B(n3910), .S(n4491), .Z(n4918) );
  OR2_X1 U3646 ( .A1(n4918), .A2(n2830), .ZN(n3115) );
  NAND2_X1 U3647 ( .A1(n3116), .A2(n3115), .ZN(n3117) );
  XNOR2_X1 U3648 ( .A(n3117), .B(n3252), .ZN(n3120) );
  NAND2_X1 U3649 ( .A1(n4928), .A2(n3237), .ZN(n3119) );
  OR2_X1 U3650 ( .A1(n4918), .A2(n3254), .ZN(n3118) );
  AND2_X1 U3651 ( .A1(n3119), .A2(n3118), .ZN(n3121) );
  NAND2_X1 U3652 ( .A1(n3120), .A2(n3121), .ZN(n3126) );
  INV_X1 U3653 ( .A(n3120), .ZN(n3123) );
  INV_X1 U3654 ( .A(n3121), .ZN(n3122) );
  NAND2_X1 U3655 ( .A1(n3123), .A2(n3122), .ZN(n3124) );
  AND2_X1 U3656 ( .A1(n3126), .A2(n3124), .ZN(n4394) );
  INV_X1 U3657 ( .A(n4394), .ZN(n3125) );
  OR2_X1 U3658 ( .A1(n3125), .A2(n4392), .ZN(n4395) );
  AND2_X1 U3659 ( .A1(n3126), .A2(n4395), .ZN(n3127) );
  NAND2_X1 U3660 ( .A1(n4396), .A2(n3127), .ZN(n4291) );
  NAND2_X1 U3661 ( .A1(n2865), .A2(REG1_REG_19__SCAN_IN), .ZN(n3133) );
  NAND2_X1 U3662 ( .A1(n2497), .A2(REG0_REG_19__SCAN_IN), .ZN(n3132) );
  NOR2_X1 U3663 ( .A1(REG3_REG_19__SCAN_IN), .A2(n3128), .ZN(n3129) );
  NOR2_X1 U3664 ( .A1(n3143), .A2(n3129), .ZN(n4901) );
  NAND2_X1 U3665 ( .A1(n2866), .A2(n4901), .ZN(n3131) );
  NAND2_X1 U3666 ( .A1(n3293), .A2(REG2_REG_19__SCAN_IN), .ZN(n3130) );
  NAND4_X1 U3667 ( .A1(n3133), .A2(n3132), .A3(n3131), .A4(n3130), .ZN(n4580)
         );
  NAND2_X1 U3668 ( .A1(n4580), .A2(n2875), .ZN(n3135) );
  INV_X1 U3669 ( .A(DATAI_19_), .ZN(n3707) );
  MUX2_X1 U3670 ( .A(n5202), .B(n3707), .S(n4491), .Z(n4898) );
  OR2_X1 U3671 ( .A1(n4898), .A2(n2830), .ZN(n3134) );
  NAND2_X1 U3672 ( .A1(n3135), .A2(n3134), .ZN(n3136) );
  XNOR2_X1 U3673 ( .A(n3136), .B(n3252), .ZN(n3141) );
  NAND2_X1 U3674 ( .A1(n4580), .A2(n3237), .ZN(n3138) );
  OR2_X1 U3675 ( .A1(n4898), .A2(n3254), .ZN(n3137) );
  NAND2_X1 U3676 ( .A1(n3138), .A2(n3137), .ZN(n3139) );
  XNOR2_X1 U3677 ( .A(n3141), .B(n3139), .ZN(n4292) );
  INV_X1 U3678 ( .A(n3139), .ZN(n3140) );
  NAND2_X1 U3679 ( .A1(n3141), .A2(n3140), .ZN(n3142) );
  NAND2_X1 U3680 ( .A1(n2496), .A2(REG0_REG_20__SCAN_IN), .ZN(n3148) );
  NAND2_X1 U3681 ( .A1(n2865), .A2(REG1_REG_20__SCAN_IN), .ZN(n3147) );
  NOR2_X1 U3682 ( .A1(n3143), .A2(REG3_REG_20__SCAN_IN), .ZN(n3144) );
  NOR2_X1 U3683 ( .A1(n3156), .A2(n3144), .ZN(n4884) );
  NAND2_X1 U3684 ( .A1(n2866), .A2(n4884), .ZN(n3146) );
  NAND2_X1 U3685 ( .A1(n3293), .A2(REG2_REG_20__SCAN_IN), .ZN(n3145) );
  OAI22_X1 U3686 ( .A1(n4862), .A2(n3254), .B1(n2830), .B2(n4881), .ZN(n3149)
         );
  XNOR2_X1 U3687 ( .A(n3149), .B(n3464), .ZN(n3152) );
  OR2_X1 U3688 ( .A1(n4862), .A2(n3251), .ZN(n3151) );
  NAND2_X1 U3689 ( .A1(n4376), .A2(n2875), .ZN(n3150) );
  NAND2_X1 U3690 ( .A1(n3151), .A2(n3150), .ZN(n3153) );
  NAND2_X1 U3691 ( .A1(n3152), .A2(n3153), .ZN(n4373) );
  INV_X1 U3692 ( .A(n3152), .ZN(n3155) );
  INV_X1 U3693 ( .A(n3153), .ZN(n3154) );
  NAND2_X1 U3694 ( .A1(n3155), .A2(n3154), .ZN(n4372) );
  NAND2_X1 U3695 ( .A1(n2865), .A2(REG1_REG_21__SCAN_IN), .ZN(n3161) );
  NAND2_X1 U3696 ( .A1(n2497), .A2(REG0_REG_21__SCAN_IN), .ZN(n3160) );
  NOR2_X1 U3697 ( .A1(n3156), .A2(REG3_REG_21__SCAN_IN), .ZN(n3157) );
  NOR2_X1 U3698 ( .A1(n3170), .A2(n3157), .ZN(n4868) );
  NAND2_X1 U3699 ( .A1(n2866), .A2(n4868), .ZN(n3159) );
  NAND2_X1 U3700 ( .A1(n3293), .A2(REG2_REG_21__SCAN_IN), .ZN(n3158) );
  NAND4_X1 U3701 ( .A1(n3161), .A2(n3160), .A3(n3159), .A4(n3158), .ZN(n4840)
         );
  NAND2_X1 U3702 ( .A1(n4840), .A2(n2875), .ZN(n3163) );
  OR2_X1 U3703 ( .A1(n4867), .A2(n2830), .ZN(n3162) );
  NAND2_X1 U3704 ( .A1(n3163), .A2(n3162), .ZN(n3164) );
  XNOR2_X1 U3705 ( .A(n3164), .B(n3252), .ZN(n3166) );
  NOR2_X1 U3706 ( .A1(n4867), .A2(n3254), .ZN(n3165) );
  AOI21_X1 U3707 ( .B1(n4840), .B2(n3237), .A(n3165), .ZN(n3167) );
  AND2_X1 U3708 ( .A1(n3166), .A2(n3167), .ZN(n4310) );
  INV_X1 U3709 ( .A(n3166), .ZN(n3169) );
  INV_X1 U3710 ( .A(n3167), .ZN(n3168) );
  NAND2_X1 U3711 ( .A1(n3169), .A2(n3168), .ZN(n4308) );
  NAND2_X1 U3712 ( .A1(n2865), .A2(REG1_REG_22__SCAN_IN), .ZN(n3175) );
  NAND2_X1 U3713 ( .A1(n2497), .A2(REG0_REG_22__SCAN_IN), .ZN(n3174) );
  NOR2_X1 U3714 ( .A1(n3170), .A2(REG3_REG_22__SCAN_IN), .ZN(n3171) );
  NOR2_X1 U3715 ( .A1(n3183), .A2(n3171), .ZN(n4853) );
  NAND2_X1 U3716 ( .A1(n2866), .A2(n4853), .ZN(n3173) );
  NAND2_X1 U3717 ( .A1(n3293), .A2(REG2_REG_22__SCAN_IN), .ZN(n3172) );
  INV_X1 U3718 ( .A(n4385), .ZN(n4852) );
  OAI22_X1 U3719 ( .A1(n4861), .A2(n3254), .B1(n2830), .B2(n4852), .ZN(n3176)
         );
  XNOR2_X1 U3720 ( .A(n3176), .B(n3464), .ZN(n3179) );
  OR2_X1 U3721 ( .A1(n4861), .A2(n3251), .ZN(n3178) );
  NAND2_X1 U3722 ( .A1(n4385), .A2(n2875), .ZN(n3177) );
  NAND2_X1 U3723 ( .A1(n3178), .A2(n3177), .ZN(n3180) );
  XNOR2_X1 U3724 ( .A(n3179), .B(n3180), .ZN(n4384) );
  INV_X1 U3725 ( .A(n3179), .ZN(n3182) );
  INV_X1 U3726 ( .A(n3180), .ZN(n3181) );
  NAND2_X1 U3727 ( .A1(n2865), .A2(REG1_REG_23__SCAN_IN), .ZN(n3189) );
  NAND2_X1 U3728 ( .A1(n2497), .A2(REG0_REG_23__SCAN_IN), .ZN(n3188) );
  NOR2_X1 U3729 ( .A1(n3183), .A2(REG3_REG_23__SCAN_IN), .ZN(n3184) );
  NOR2_X1 U3730 ( .A1(n3185), .A2(n3184), .ZN(n4274) );
  NAND2_X1 U3731 ( .A1(n2866), .A2(n4274), .ZN(n3187) );
  NAND2_X1 U3732 ( .A1(n3293), .A2(REG2_REG_23__SCAN_IN), .ZN(n3186) );
  NAND2_X1 U3733 ( .A1(n4839), .A2(n2875), .ZN(n3191) );
  OR2_X1 U3734 ( .A1(n4716), .A2(n2830), .ZN(n3190) );
  NAND2_X1 U3735 ( .A1(n3191), .A2(n3190), .ZN(n3192) );
  XNOR2_X1 U3736 ( .A(n3192), .B(n3252), .ZN(n3194) );
  NOR2_X1 U3737 ( .A1(n4716), .A2(n3254), .ZN(n3193) );
  AOI21_X1 U3738 ( .B1(n4839), .B2(n3237), .A(n3193), .ZN(n3195) );
  XNOR2_X1 U3739 ( .A(n3194), .B(n3195), .ZN(n4270) );
  INV_X1 U3740 ( .A(n3194), .ZN(n3197) );
  INV_X1 U3741 ( .A(n3195), .ZN(n3196) );
  NAND2_X1 U3742 ( .A1(n3197), .A2(n3196), .ZN(n3198) );
  NAND2_X1 U3743 ( .A1(n4271), .A2(n3198), .ZN(n3203) );
  NAND2_X1 U3744 ( .A1(n4720), .A2(n2875), .ZN(n3200) );
  OR2_X1 U3745 ( .A1(n4822), .A2(n2830), .ZN(n3199) );
  NAND2_X1 U3746 ( .A1(n3200), .A2(n3199), .ZN(n3201) );
  XNOR2_X1 U3747 ( .A(n3201), .B(n3464), .ZN(n3202) );
  NAND2_X1 U3748 ( .A1(n2496), .A2(REG0_REG_25__SCAN_IN), .ZN(n3209) );
  NAND2_X1 U3749 ( .A1(n2865), .A2(REG1_REG_25__SCAN_IN), .ZN(n3208) );
  NOR2_X1 U3750 ( .A1(n3204), .A2(REG3_REG_25__SCAN_IN), .ZN(n3205) );
  NOR2_X1 U3751 ( .A1(n3215), .A2(n3205), .ZN(n4813) );
  NAND2_X1 U3752 ( .A1(n2866), .A2(n4813), .ZN(n3207) );
  NAND2_X1 U3753 ( .A1(n3293), .A2(REG2_REG_25__SCAN_IN), .ZN(n3206) );
  OAI22_X1 U3754 ( .A1(n4823), .A2(n3254), .B1(n2830), .B2(n4810), .ZN(n3210)
         );
  XNOR2_X1 U3755 ( .A(n3210), .B(n3252), .ZN(n4322) );
  OR2_X1 U3756 ( .A1(n4823), .A2(n3251), .ZN(n3212) );
  NAND2_X1 U3757 ( .A1(n4724), .A2(n2875), .ZN(n3211) );
  INV_X1 U3758 ( .A(n4322), .ZN(n3214) );
  NAND2_X1 U3759 ( .A1(n2865), .A2(REG1_REG_26__SCAN_IN), .ZN(n3220) );
  NAND2_X1 U3760 ( .A1(n2497), .A2(REG0_REG_26__SCAN_IN), .ZN(n3219) );
  NOR2_X1 U3761 ( .A1(n3215), .A2(REG3_REG_26__SCAN_IN), .ZN(n3216) );
  NOR2_X1 U3762 ( .A1(n3227), .A2(n3216), .ZN(n4411) );
  NAND2_X1 U3763 ( .A1(n2866), .A2(n4411), .ZN(n3218) );
  NAND2_X1 U3764 ( .A1(n3293), .A2(REG2_REG_26__SCAN_IN), .ZN(n3217) );
  NAND2_X1 U3765 ( .A1(n4809), .A2(n2875), .ZN(n3222) );
  NAND2_X1 U3766 ( .A1(n2872), .A2(DATAI_26_), .ZN(n4785) );
  OR2_X1 U3767 ( .A1(n4785), .A2(n2830), .ZN(n3221) );
  NAND2_X1 U3768 ( .A1(n3222), .A2(n3221), .ZN(n3223) );
  XNOR2_X1 U3769 ( .A(n3223), .B(n3252), .ZN(n3226) );
  NOR2_X1 U3770 ( .A1(n4785), .A2(n3254), .ZN(n3224) );
  AOI21_X1 U3771 ( .B1(n4809), .B2(n3237), .A(n3224), .ZN(n3225) );
  AND2_X1 U3772 ( .A1(n3226), .A2(n3225), .ZN(n4406) );
  OR2_X1 U3773 ( .A1(n3226), .A2(n3225), .ZN(n4407) );
  NAND2_X1 U3774 ( .A1(n2865), .A2(REG1_REG_27__SCAN_IN), .ZN(n3233) );
  NAND2_X1 U3775 ( .A1(n2496), .A2(REG0_REG_27__SCAN_IN), .ZN(n3232) );
  NAND2_X1 U3776 ( .A1(n3227), .A2(REG3_REG_27__SCAN_IN), .ZN(n3245) );
  INV_X1 U3777 ( .A(n3227), .ZN(n3228) );
  INV_X1 U3778 ( .A(REG3_REG_27__SCAN_IN), .ZN(n3742) );
  NAND2_X1 U3779 ( .A1(n3228), .A2(n3742), .ZN(n3229) );
  NAND2_X1 U3780 ( .A1(n2866), .A2(n4772), .ZN(n3231) );
  NAND2_X1 U3781 ( .A1(n3293), .A2(REG2_REG_27__SCAN_IN), .ZN(n3230) );
  NAND2_X1 U3782 ( .A1(n4787), .A2(n2875), .ZN(n3235) );
  OR2_X1 U3783 ( .A1(n4770), .A2(n2830), .ZN(n3234) );
  NAND2_X1 U3784 ( .A1(n3235), .A2(n3234), .ZN(n3236) );
  XNOR2_X1 U3785 ( .A(n3236), .B(n3464), .ZN(n3241) );
  INV_X1 U3786 ( .A(n3241), .ZN(n3243) );
  NAND2_X1 U3787 ( .A1(n4787), .A2(n3237), .ZN(n3239) );
  OR2_X1 U3788 ( .A1(n4770), .A2(n3254), .ZN(n3238) );
  NAND2_X1 U3789 ( .A1(n3239), .A2(n3238), .ZN(n3240) );
  INV_X1 U3790 ( .A(n3240), .ZN(n3242) );
  AOI21_X1 U3791 ( .B1(n3243), .B2(n3242), .A(n3282), .ZN(n4263) );
  NAND2_X1 U3792 ( .A1(n4264), .A2(n4263), .ZN(n4262) );
  INV_X1 U3793 ( .A(n4262), .ZN(n3279) );
  NAND2_X1 U3794 ( .A1(n2497), .A2(REG0_REG_28__SCAN_IN), .ZN(n3250) );
  NAND2_X1 U3795 ( .A1(n2865), .A2(REG1_REG_28__SCAN_IN), .ZN(n3249) );
  INV_X1 U3796 ( .A(n3245), .ZN(n3244) );
  NAND2_X1 U3797 ( .A1(n3244), .A2(REG3_REG_28__SCAN_IN), .ZN(n4736) );
  INV_X1 U3798 ( .A(REG3_REG_28__SCAN_IN), .ZN(n3303) );
  NAND2_X1 U3799 ( .A1(n3245), .A2(n3303), .ZN(n3246) );
  NAND2_X1 U3800 ( .A1(n2866), .A2(n4754), .ZN(n3248) );
  NAND2_X1 U3801 ( .A1(n3293), .A2(REG2_REG_28__SCAN_IN), .ZN(n3247) );
  OAI22_X1 U3802 ( .A1(n4729), .A2(n3251), .B1(n3254), .B2(n4744), .ZN(n3253)
         );
  XNOR2_X1 U3803 ( .A(n3253), .B(n3252), .ZN(n3256) );
  OAI22_X1 U3804 ( .A1(n4729), .A2(n3254), .B1(n2830), .B2(n4744), .ZN(n3255)
         );
  XNOR2_X1 U3805 ( .A(n3256), .B(n3255), .ZN(n3281) );
  INV_X1 U3806 ( .A(n5038), .ZN(n3262) );
  NAND2_X1 U3807 ( .A1(n3262), .A2(B_REG_SCAN_IN), .ZN(n3257) );
  MUX2_X1 U3808 ( .A(n3257), .B(B_REG_SCAN_IN), .S(n5039), .Z(n3258) );
  INV_X1 U3809 ( .A(D_REG_0__SCAN_IN), .ZN(n3322) );
  NAND2_X1 U3810 ( .A1(n3317), .A2(n3322), .ZN(n3260) );
  INV_X1 U3811 ( .A(n5037), .ZN(n3263) );
  INV_X1 U3812 ( .A(n5039), .ZN(n3259) );
  NAND2_X1 U3813 ( .A1(n3263), .A2(n3259), .ZN(n3320) );
  INV_X1 U3814 ( .A(D_REG_1__SCAN_IN), .ZN(n3261) );
  NAND2_X1 U3815 ( .A1(n3317), .A2(n3261), .ZN(n3264) );
  NAND2_X1 U3816 ( .A1(n3263), .A2(n3262), .ZN(n5032) );
  NAND2_X1 U3817 ( .A1(n3264), .A2(n5032), .ZN(n4975) );
  INV_X1 U3818 ( .A(n4975), .ZN(n3461) );
  NOR2_X1 U3819 ( .A1(D_REG_10__SCAN_IN), .A2(D_REG_13__SCAN_IN), .ZN(n3268)
         );
  NOR4_X1 U3820 ( .A1(D_REG_31__SCAN_IN), .A2(D_REG_25__SCAN_IN), .A3(
        D_REG_16__SCAN_IN), .A4(D_REG_17__SCAN_IN), .ZN(n3267) );
  NOR4_X1 U3821 ( .A1(D_REG_26__SCAN_IN), .A2(D_REG_27__SCAN_IN), .A3(
        D_REG_30__SCAN_IN), .A4(D_REG_8__SCAN_IN), .ZN(n3266) );
  NOR4_X1 U3822 ( .A1(D_REG_15__SCAN_IN), .A2(D_REG_12__SCAN_IN), .A3(
        D_REG_9__SCAN_IN), .A4(D_REG_2__SCAN_IN), .ZN(n3265) );
  NAND4_X1 U3823 ( .A1(n3268), .A2(n3267), .A3(n3266), .A4(n3265), .ZN(n3274)
         );
  NOR4_X1 U3824 ( .A1(D_REG_11__SCAN_IN), .A2(D_REG_14__SCAN_IN), .A3(
        D_REG_18__SCAN_IN), .A4(D_REG_19__SCAN_IN), .ZN(n3272) );
  NOR4_X1 U3825 ( .A1(D_REG_6__SCAN_IN), .A2(D_REG_4__SCAN_IN), .A3(
        D_REG_5__SCAN_IN), .A4(D_REG_7__SCAN_IN), .ZN(n3271) );
  NOR4_X1 U3826 ( .A1(D_REG_24__SCAN_IN), .A2(D_REG_28__SCAN_IN), .A3(
        D_REG_29__SCAN_IN), .A4(D_REG_3__SCAN_IN), .ZN(n3270) );
  NOR4_X1 U3827 ( .A1(D_REG_20__SCAN_IN), .A2(D_REG_21__SCAN_IN), .A3(
        D_REG_23__SCAN_IN), .A4(D_REG_22__SCAN_IN), .ZN(n3269) );
  NAND4_X1 U3828 ( .A1(n3272), .A2(n3271), .A3(n3270), .A4(n3269), .ZN(n3273)
         );
  NAND3_X1 U3829 ( .A1(n5018), .A2(n3461), .A3(n4976), .ZN(n3298) );
  INV_X1 U3830 ( .A(n3298), .ZN(n3276) );
  NAND2_X1 U3831 ( .A1(n2814), .A2(IR_REG_31__SCAN_IN), .ZN(n3275) );
  NAND2_X1 U3832 ( .A1(n3276), .A2(n4571), .ZN(n3287) );
  NAND2_X1 U3833 ( .A1(n3300), .A2(n3288), .ZN(n3299) );
  INV_X1 U3834 ( .A(n3465), .ZN(n3466) );
  NAND2_X1 U3835 ( .A1(n3299), .A2(n3466), .ZN(n3277) );
  NAND2_X1 U3836 ( .A1(n3279), .A2(n3278), .ZN(n3312) );
  INV_X1 U3837 ( .A(n3282), .ZN(n3280) );
  INV_X1 U3838 ( .A(n3281), .ZN(n3283) );
  NAND3_X1 U3839 ( .A1(n3283), .A2(n5282), .A3(n3282), .ZN(n3309) );
  OR2_X1 U3840 ( .A1(n2818), .A2(n3284), .ZN(n4573) );
  OR2_X1 U3841 ( .A1(n3287), .A2(n4573), .ZN(n3291) );
  INV_X1 U3842 ( .A(n4399), .ZN(n5272) );
  OR2_X1 U3843 ( .A1(n3287), .A2(n5319), .ZN(n3290) );
  AOI22_X1 U3844 ( .A1(n4410), .A2(n4787), .B1(n4751), .B2(n5276), .ZN(n3307)
         );
  INV_X1 U3845 ( .A(n3285), .ZN(n3337) );
  NAND2_X1 U3846 ( .A1(n2496), .A2(REG0_REG_29__SCAN_IN), .ZN(n3297) );
  NAND2_X1 U3847 ( .A1(n2865), .A2(REG1_REG_29__SCAN_IN), .ZN(n3296) );
  INV_X1 U3848 ( .A(n4736), .ZN(n3292) );
  NAND2_X1 U3849 ( .A1(n2866), .A2(n3292), .ZN(n3295) );
  NAND2_X1 U3850 ( .A1(n3293), .A2(REG2_REG_29__SCAN_IN), .ZN(n3294) );
  NAND4_X1 U3851 ( .A1(n3297), .A2(n3296), .A3(n3295), .A4(n3294), .ZN(n4750)
         );
  OAI21_X1 U3852 ( .B1(n4567), .B2(n3299), .A(n3298), .ZN(n3429) );
  NAND2_X1 U3853 ( .A1(n3300), .A2(n3465), .ZN(n3428) );
  AND3_X1 U3854 ( .A1(n2878), .A2(n3329), .A3(n3428), .ZN(n3301) );
  NAND2_X1 U3855 ( .A1(n3429), .A2(n3301), .ZN(n3302) );
  INV_X1 U3856 ( .A(n4754), .ZN(n3304) );
  OAI22_X1 U3857 ( .A1(n5287), .A2(n3304), .B1(STATE_REG_SCAN_IN), .B2(n3303), 
        .ZN(n3305) );
  AOI21_X1 U3858 ( .B1(n4414), .B2(n4750), .A(n3305), .ZN(n3306) );
  AND2_X1 U3859 ( .A1(n3307), .A2(n3306), .ZN(n3308) );
  NAND2_X1 U3860 ( .A1(n3312), .A2(n3311), .ZN(U3217) );
  INV_X1 U3861 ( .A(n3313), .ZN(n3319) );
  INV_X2 U3862 ( .A(STATE_REG_SCAN_IN), .ZN(U3149) );
  INV_X1 U3863 ( .A(DATAI_23_), .ZN(n3314) );
  AOI21_X1 U3864 ( .B1(n3314), .B2(U3149), .A(n3313), .ZN(U3329) );
  INV_X1 U3865 ( .A(DATAI_20_), .ZN(n3315) );
  MUX2_X1 U3866 ( .A(n3315), .B(n3286), .S(STATE_REG_SCAN_IN), .Z(n3316) );
  INV_X1 U3867 ( .A(n3316), .ZN(U3332) );
  INV_X1 U3868 ( .A(n3317), .ZN(n3318) );
  NOR2_X1 U3869 ( .A1(n3320), .A2(n3319), .ZN(n3321) );
  AOI21_X1 U3870 ( .B1(n5086), .B2(n3322), .A(n3321), .ZN(U3458) );
  INV_X1 U3871 ( .A(DATAI_28_), .ZN(n3323) );
  MUX2_X1 U3872 ( .A(n3285), .B(n3323), .S(U3149), .Z(n3324) );
  INV_X1 U3873 ( .A(n3324), .ZN(U3324) );
  INV_X1 U3874 ( .A(REG1_REG_0__SCAN_IN), .ZN(n5111) );
  NOR2_X1 U3875 ( .A1(n4710), .A2(REG2_REG_0__SCAN_IN), .ZN(n3325) );
  OR2_X1 U3876 ( .A1(n3325), .A2(n3285), .ZN(n3407) );
  AOI21_X1 U3877 ( .B1(n5111), .B2(n4710), .A(n3407), .ZN(n3326) );
  MUX2_X1 U3878 ( .A(n3326), .B(n3407), .S(IR_REG_0__SCAN_IN), .Z(n3327) );
  INV_X1 U3879 ( .A(n3327), .ZN(n3336) );
  OR2_X1 U3880 ( .A1(n3329), .A2(U3149), .ZN(n4577) );
  INV_X1 U3881 ( .A(n4577), .ZN(n3328) );
  OR2_X1 U3882 ( .A1(n4571), .A2(n3328), .ZN(n3331) );
  NAND2_X1 U3883 ( .A1(n3465), .A2(n3329), .ZN(n3330) );
  AND2_X1 U3884 ( .A1(n4491), .A2(n3330), .ZN(n3332) );
  NAND2_X1 U3885 ( .A1(n3331), .A2(n3332), .ZN(n3338) );
  INV_X1 U3886 ( .A(n3331), .ZN(n3333) );
  NOR2_X2 U3887 ( .A1(n3333), .A2(n3332), .ZN(n5088) );
  AOI22_X1 U3888 ( .A1(n5088), .A2(ADDR_REG_0__SCAN_IN), .B1(
        REG3_REG_0__SCAN_IN), .B2(U3149), .ZN(n3335) );
  INV_X1 U3889 ( .A(n4710), .ZN(n4093) );
  NAND3_X1 U3890 ( .A1(n5099), .A2(IR_REG_0__SCAN_IN), .A3(n5111), .ZN(n3334)
         );
  OAI211_X1 U3891 ( .C1(n3336), .C2(n3338), .A(n3335), .B(n3334), .ZN(U3240)
         );
  NAND2_X1 U3892 ( .A1(IR_REG_0__SCAN_IN), .A2(REG2_REG_0__SCAN_IN), .ZN(n3399) );
  OR2_X1 U3893 ( .A1(n3285), .A2(n4710), .ZN(n4572) );
  AOI211_X1 U3894 ( .C1(n3399), .C2(n3339), .A(n3349), .B(n5090), .ZN(n3343)
         );
  INV_X1 U3895 ( .A(REG1_REG_1__SCAN_IN), .ZN(n5130) );
  AOI211_X1 U3896 ( .C1(n3341), .C2(n3340), .A(n3361), .B(n4671), .ZN(n3342)
         );
  NOR2_X1 U3897 ( .A1(n3343), .A2(n3342), .ZN(n3345) );
  AOI22_X1 U3898 ( .A1(n5088), .A2(ADDR_REG_1__SCAN_IN), .B1(
        REG3_REG_1__SCAN_IN), .B2(U3149), .ZN(n3344) );
  OAI211_X1 U3899 ( .C1(n3346), .C2(n5089), .A(n3345), .B(n3344), .ZN(U3241)
         );
  NOR2_X1 U3900 ( .A1(n5088), .A2(U4043), .ZN(U3148) );
  AND2_X1 U3901 ( .A1(n3347), .A2(REG2_REG_1__SCAN_IN), .ZN(n3348) );
  NOR2_X1 U3902 ( .A1(n3412), .A2(n3411), .ZN(n3410) );
  NOR2_X1 U3903 ( .A1(n3350), .A2(n3396), .ZN(n3351) );
  INV_X1 U3904 ( .A(REG2_REG_3__SCAN_IN), .ZN(n3391) );
  XNOR2_X1 U3905 ( .A(n3350), .B(n3396), .ZN(n3390) );
  NOR2_X1 U3906 ( .A1(n3391), .A2(n3390), .ZN(n3389) );
  INV_X1 U3907 ( .A(REG2_REG_4__SCAN_IN), .ZN(n5092) );
  NOR2_X1 U3908 ( .A1(n3353), .A2(n3352), .ZN(n3354) );
  INV_X1 U3909 ( .A(REG2_REG_5__SCAN_IN), .ZN(n3355) );
  MUX2_X1 U3910 ( .A(n3355), .B(REG2_REG_5__SCAN_IN), .S(n5055), .Z(n3383) );
  INV_X1 U3911 ( .A(REG2_REG_6__SCAN_IN), .ZN(n3517) );
  NAND2_X1 U3912 ( .A1(n5053), .A2(REG2_REG_7__SCAN_IN), .ZN(n3358) );
  OAI21_X1 U3913 ( .B1(n5053), .B2(REG2_REG_7__SCAN_IN), .A(n3358), .ZN(n3359)
         );
  AOI211_X1 U3914 ( .C1(n3360), .C2(n3359), .A(n3441), .B(n5090), .ZN(n3377)
         );
  INV_X1 U3915 ( .A(n5053), .ZN(n3375) );
  INV_X1 U3916 ( .A(REG1_REG_2__SCAN_IN), .ZN(n5137) );
  MUX2_X1 U3917 ( .A(n5137), .B(REG1_REG_2__SCAN_IN), .S(n5057), .Z(n3409) );
  NAND2_X1 U3918 ( .A1(n5056), .A2(n3362), .ZN(n3363) );
  XNOR2_X1 U3919 ( .A(n3396), .B(n3362), .ZN(n3393) );
  NAND2_X1 U3920 ( .A1(REG1_REG_3__SCAN_IN), .A2(n3393), .ZN(n3392) );
  NAND2_X1 U3921 ( .A1(n5096), .A2(n3364), .ZN(n3365) );
  INV_X1 U3922 ( .A(REG1_REG_5__SCAN_IN), .ZN(n5196) );
  MUX2_X1 U3923 ( .A(n5196), .B(REG1_REG_5__SCAN_IN), .S(n5055), .Z(n3379) );
  INV_X1 U3924 ( .A(REG1_REG_6__SCAN_IN), .ZN(n3367) );
  INV_X1 U3925 ( .A(REG1_REG_7__SCAN_IN), .ZN(n3369) );
  MUX2_X1 U3926 ( .A(REG1_REG_7__SCAN_IN), .B(n3369), .S(n5053), .Z(n3370) );
  OAI211_X1 U3927 ( .C1(n3371), .C2(n3370), .A(n5099), .B(n3443), .ZN(n3374)
         );
  INV_X1 U3928 ( .A(REG3_REG_7__SCAN_IN), .ZN(n3372) );
  NOR2_X1 U3929 ( .A1(STATE_REG_SCAN_IN), .A2(n3372), .ZN(n4258) );
  AOI21_X1 U3930 ( .B1(n5088), .B2(ADDR_REG_7__SCAN_IN), .A(n4258), .ZN(n3373)
         );
  OAI211_X1 U3931 ( .C1(n5089), .C2(n3375), .A(n3374), .B(n3373), .ZN(n3376)
         );
  OR2_X1 U3932 ( .A1(n3377), .A2(n3376), .ZN(U3247) );
  INV_X1 U3933 ( .A(n5055), .ZN(n3388) );
  AOI211_X1 U3934 ( .C1(n3380), .C2(n3379), .A(n4671), .B(n3378), .ZN(n3381)
         );
  INV_X1 U3935 ( .A(n3381), .ZN(n3387) );
  INV_X1 U3936 ( .A(REG3_REG_5__SCAN_IN), .ZN(n3382) );
  NOR2_X1 U3937 ( .A1(STATE_REG_SCAN_IN), .A2(n3382), .ZN(n3527) );
  AOI211_X1 U3938 ( .C1(n3384), .C2(n3383), .A(n2545), .B(n5090), .ZN(n3385)
         );
  AOI211_X1 U3939 ( .C1(n5088), .C2(ADDR_REG_5__SCAN_IN), .A(n3527), .B(n3385), 
        .ZN(n3386) );
  OAI211_X1 U3940 ( .C1(n5089), .C2(n3388), .A(n3387), .B(n3386), .ZN(U3245)
         );
  AOI211_X1 U3941 ( .C1(n3391), .C2(n3390), .A(n3389), .B(n5090), .ZN(n3398)
         );
  OAI211_X1 U3942 ( .C1(REG1_REG_3__SCAN_IN), .C2(n3393), .A(n5099), .B(n3392), 
        .ZN(n3395) );
  NOR2_X1 U3943 ( .A1(STATE_REG_SCAN_IN), .A2(n3944), .ZN(n3437) );
  AOI21_X1 U3944 ( .B1(n5088), .B2(ADDR_REG_3__SCAN_IN), .A(n3437), .ZN(n3394)
         );
  OAI211_X1 U3945 ( .C1(n5089), .C2(n3396), .A(n3395), .B(n3394), .ZN(n3397)
         );
  OR2_X1 U3946 ( .A1(n3398), .A2(n3397), .ZN(U3243) );
  OAI21_X1 U3947 ( .B1(n3399), .B2(n4572), .A(U4043), .ZN(n3406) );
  AOI21_X1 U3948 ( .B1(n2591), .B2(n5111), .A(n2878), .ZN(n3400) );
  NOR3_X1 U3949 ( .A1(n3402), .A2(n3401), .A3(n3400), .ZN(n3404) );
  NOR2_X1 U3950 ( .A1(n3404), .A2(n3403), .ZN(n3430) );
  NOR3_X1 U3951 ( .A1(n3430), .A2(n4093), .A3(n3285), .ZN(n3405) );
  AOI211_X1 U3952 ( .C1(n2591), .C2(n3407), .A(n3406), .B(n3405), .ZN(n5094)
         );
  XOR2_X1 U3953 ( .A(n3409), .B(n3408), .Z(n3414) );
  AOI211_X1 U3954 ( .C1(n3412), .C2(n3411), .A(n3410), .B(n5090), .ZN(n3413)
         );
  AOI21_X1 U3955 ( .B1(n5099), .B2(n3414), .A(n3413), .ZN(n3416) );
  AOI22_X1 U3956 ( .A1(n5088), .A2(ADDR_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(U3149), .ZN(n3415) );
  OAI211_X1 U3957 ( .C1(n3417), .C2(n5089), .A(n3416), .B(n3415), .ZN(n3418)
         );
  OR2_X1 U3958 ( .A1(n5094), .A2(n3418), .ZN(U3242) );
  XNOR2_X1 U3959 ( .A(n3419), .B(REG1_REG_6__SCAN_IN), .ZN(n3426) );
  INV_X1 U3960 ( .A(REG3_REG_6__SCAN_IN), .ZN(n3420) );
  NOR2_X1 U3961 ( .A1(n3420), .A2(STATE_REG_SCAN_IN), .ZN(n3549) );
  AOI21_X1 U3962 ( .B1(n5088), .B2(ADDR_REG_6__SCAN_IN), .A(n3549), .ZN(n3421)
         );
  OAI21_X1 U3963 ( .B1(n2710), .B2(n5089), .A(n3421), .ZN(n3425) );
  AOI211_X1 U3964 ( .C1(n3423), .C2(n3517), .A(n3422), .B(n5090), .ZN(n3424)
         );
  AOI211_X1 U3965 ( .C1(n5099), .C2(n3426), .A(n3425), .B(n3424), .ZN(n3427)
         );
  INV_X1 U3966 ( .A(n3427), .ZN(U3246) );
  NAND2_X1 U3967 ( .A1(n3429), .A2(n4977), .ZN(n4303) );
  AOI22_X1 U3968 ( .A1(n3430), .A2(n5282), .B1(REG3_REG_0__SCAN_IN), .B2(n4303), .ZN(n3432) );
  AOI22_X1 U3969 ( .A1(n4414), .A2(n3457), .B1(n4419), .B2(n5276), .ZN(n3431)
         );
  NAND2_X1 U3970 ( .A1(n3432), .A2(n3431), .ZN(U3229) );
  NAND2_X1 U3971 ( .A1(n4361), .A2(n3433), .ZN(n3434) );
  XOR2_X1 U3972 ( .A(n3435), .B(n3434), .Z(n3440) );
  AOI22_X1 U3973 ( .A1(n4410), .A2(n4591), .B1(n4218), .B2(n5276), .ZN(n3439)
         );
  NOR2_X1 U3974 ( .A1(n5287), .A2(REG3_REG_3__SCAN_IN), .ZN(n3436) );
  AOI211_X1 U3975 ( .C1(n4414), .C2(n4590), .A(n3437), .B(n3436), .ZN(n3438)
         );
  OAI211_X1 U3976 ( .C1(n3440), .C2(n4417), .A(n3439), .B(n3438), .ZN(U3215)
         );
  INV_X1 U3977 ( .A(REG2_REG_8__SCAN_IN), .ZN(n3581) );
  AOI211_X1 U3978 ( .C1(n3581), .C2(n3442), .A(n3533), .B(n5090), .ZN(n3450)
         );
  NAND2_X1 U3979 ( .A1(n5053), .A2(REG1_REG_7__SCAN_IN), .ZN(n3444) );
  NAND2_X1 U3980 ( .A1(n3444), .A2(n3443), .ZN(n3536) );
  XNOR2_X1 U3981 ( .A(n3536), .B(n3531), .ZN(n3445) );
  NAND2_X1 U3982 ( .A1(REG1_REG_8__SCAN_IN), .A2(n3445), .ZN(n3537) );
  OAI211_X1 U3983 ( .C1(n3445), .C2(REG1_REG_8__SCAN_IN), .A(n5099), .B(n3537), 
        .ZN(n3448) );
  INV_X1 U3984 ( .A(REG3_REG_8__SCAN_IN), .ZN(n3446) );
  NOR2_X1 U3985 ( .A1(STATE_REG_SCAN_IN), .A2(n3446), .ZN(n3606) );
  AOI21_X1 U3986 ( .B1(n5088), .B2(ADDR_REG_8__SCAN_IN), .A(n3606), .ZN(n3447)
         );
  OAI211_X1 U3987 ( .C1(n5089), .C2(n3531), .A(n3448), .B(n3447), .ZN(n3449)
         );
  OR2_X1 U3988 ( .A1(n3450), .A2(n3449), .ZN(U3248) );
  INV_X1 U3989 ( .A(n4361), .ZN(n3451) );
  AOI21_X1 U3990 ( .B1(n3453), .B2(n3452), .A(n3451), .ZN(n3456) );
  AOI22_X1 U3991 ( .A1(n5276), .A2(n3493), .B1(REG3_REG_2__SCAN_IN), .B2(n4303), .ZN(n3455) );
  AOI22_X1 U3992 ( .A1(n4414), .A2(n5156), .B1(n4410), .B2(n3457), .ZN(n3454)
         );
  OAI211_X1 U3993 ( .C1(n3456), .C2(n4417), .A(n3455), .B(n3454), .ZN(U3234)
         );
  NAND2_X1 U3994 ( .A1(n5110), .A2(n4304), .ZN(n3483) );
  AND2_X1 U3995 ( .A1(n4593), .A2(n4419), .ZN(n3459) );
  NAND2_X1 U3996 ( .A1(n3458), .A2(n3459), .ZN(n3485) );
  OR2_X1 U3997 ( .A1(n3482), .A2(n3459), .ZN(n3460) );
  NAND2_X1 U3998 ( .A1(n3485), .A2(n3460), .ZN(n5124) );
  NAND4_X1 U3999 ( .A1(n4977), .A2(n3461), .A3(n4978), .A4(n4976), .ZN(n3462)
         );
  INV_X2 U4000 ( .A(n5330), .ZN(n5208) );
  NOR2_X1 U4001 ( .A1(n2818), .A2(n5202), .ZN(n3463) );
  NAND2_X1 U4002 ( .A1(n5208), .A2(n3463), .ZN(n4795) );
  NAND2_X1 U4003 ( .A1(n5199), .A2(n5202), .ZN(n4968) );
  NAND2_X1 U4004 ( .A1(n4593), .A2(n5157), .ZN(n3468) );
  INV_X1 U4005 ( .A(n5319), .ZN(n5191) );
  NAND2_X1 U4006 ( .A1(n4304), .A2(n5191), .ZN(n3467) );
  OAI211_X1 U4007 ( .C1(n3508), .C2(n5188), .A(n3468), .B(n3467), .ZN(n3469)
         );
  INV_X1 U4008 ( .A(n3469), .ZN(n3475) );
  INV_X1 U4009 ( .A(n4593), .ZN(n4420) );
  NAND2_X1 U4010 ( .A1(n4420), .A2(n4419), .ZN(n5104) );
  XNOR2_X1 U4011 ( .A(n3482), .B(n5104), .ZN(n3473) );
  NAND2_X1 U4012 ( .A1(n4567), .A2(n5041), .ZN(n3472) );
  OR2_X1 U4013 ( .A1(n5202), .A2(n3470), .ZN(n3471) );
  NAND2_X1 U4014 ( .A1(n3473), .A2(n5108), .ZN(n3474) );
  OAI211_X1 U4015 ( .C1(n5124), .C2(n4968), .A(n3475), .B(n3474), .ZN(n5127)
         );
  MUX2_X1 U4016 ( .A(n5127), .B(REG2_REG_1__SCAN_IN), .S(n5330), .Z(n3476) );
  INV_X1 U4017 ( .A(n3476), .ZN(n3481) );
  AND2_X1 U4018 ( .A1(n5208), .A2(n3477), .ZN(n5328) );
  NOR2_X1 U4019 ( .A1(n3478), .A2(n5107), .ZN(n5126) );
  NAND2_X1 U4020 ( .A1(n3478), .A2(n5107), .ZN(n3494) );
  INV_X1 U4021 ( .A(n3494), .ZN(n5125) );
  NOR3_X1 U4022 ( .A1(n4904), .A2(n5126), .A3(n5125), .ZN(n3479) );
  AOI21_X1 U4023 ( .B1(n5118), .B2(REG3_REG_1__SCAN_IN), .A(n3479), .ZN(n3480)
         );
  OAI211_X1 U4024 ( .C1(n5124), .C2(n4795), .A(n3481), .B(n3480), .ZN(U3289)
         );
  NAND2_X1 U4025 ( .A1(n4591), .A2(n3507), .ZN(n4425) );
  NAND2_X1 U4026 ( .A1(n3508), .A2(n3493), .ZN(n4422) );
  XOR2_X1 U4027 ( .A(n4534), .B(n3499), .Z(n3492) );
  NAND2_X1 U4028 ( .A1(n3457), .A2(n4304), .ZN(n3484) );
  NAND2_X1 U4029 ( .A1(n3485), .A2(n3484), .ZN(n3487) );
  NAND2_X1 U4030 ( .A1(n3487), .A2(n4534), .ZN(n3488) );
  NAND2_X1 U4031 ( .A1(n3510), .A2(n3488), .ZN(n5136) );
  INV_X1 U4032 ( .A(n4968), .ZN(n5163) );
  AOI22_X1 U4033 ( .A1(n3457), .A2(n5157), .B1(n5154), .B2(n5156), .ZN(n3489)
         );
  OAI21_X1 U4034 ( .B1(n3507), .B2(n5319), .A(n3489), .ZN(n3490) );
  AOI21_X1 U4035 ( .B1(n5136), .B2(n5163), .A(n3490), .ZN(n3491) );
  OAI21_X1 U4036 ( .B1(n3492), .B2(n5194), .A(n3491), .ZN(n5134) );
  INV_X1 U4037 ( .A(n5134), .ZN(n3498) );
  INV_X1 U4038 ( .A(n4795), .ZN(n5119) );
  OAI21_X1 U4039 ( .B1(n5125), .B2(n3507), .A(n4217), .ZN(n5133) );
  AOI22_X1 U4040 ( .A1(n5330), .A2(REG2_REG_2__SCAN_IN), .B1(
        REG3_REG_2__SCAN_IN), .B2(n5118), .ZN(n3495) );
  OAI21_X1 U4041 ( .B1(n5133), .B2(n4904), .A(n3495), .ZN(n3496) );
  AOI21_X1 U4042 ( .B1(n5136), .B2(n5119), .A(n3496), .ZN(n3497) );
  OAI21_X1 U40430 ( .B1(n3498), .B2(n5330), .A(n3497), .ZN(U3288) );
  INV_X1 U4044 ( .A(n5156), .ZN(n3500) );
  NAND2_X1 U4045 ( .A1(n3500), .A2(n4218), .ZN(n4427) );
  INV_X1 U4046 ( .A(n4218), .ZN(n4213) );
  NAND2_X1 U4047 ( .A1(n5156), .A2(n4213), .ZN(n4424) );
  NAND2_X1 U4048 ( .A1(n4211), .A2(n4538), .ZN(n3501) );
  NAND2_X1 U4049 ( .A1(n3501), .A2(n4427), .ZN(n5152) );
  NAND2_X1 U4050 ( .A1(n4590), .A2(n5150), .ZN(n4432) );
  NAND2_X1 U4051 ( .A1(n5152), .A2(n4432), .ZN(n3502) );
  NAND2_X1 U4052 ( .A1(n5187), .A2(n5158), .ZN(n4428) );
  XNOR2_X1 U4053 ( .A(n5155), .B(n5180), .ZN(n5184) );
  NAND2_X1 U4054 ( .A1(n5155), .A2(n5180), .ZN(n4430) );
  INV_X1 U4055 ( .A(n4589), .ZN(n5189) );
  NAND2_X1 U4056 ( .A1(n5189), .A2(n3562), .ZN(n4433) );
  INV_X1 U4057 ( .A(n3562), .ZN(n3503) );
  NAND2_X1 U4058 ( .A1(n4589), .A2(n3503), .ZN(n4451) );
  XNOR2_X1 U4059 ( .A(n3554), .B(n4537), .ZN(n3506) );
  AOI22_X1 U4060 ( .A1(n4588), .A2(n5154), .B1(n5157), .B2(n5155), .ZN(n3505)
         );
  NAND2_X1 U4061 ( .A1(n3562), .A2(n5191), .ZN(n3504) );
  OAI211_X1 U4062 ( .C1(n3506), .C2(n5194), .A(n3505), .B(n3504), .ZN(n5212)
         );
  INV_X1 U4063 ( .A(n5212), .ZN(n3521) );
  NAND2_X1 U4064 ( .A1(n3508), .A2(n3507), .ZN(n3509) );
  NAND2_X1 U4065 ( .A1(n5156), .A2(n4218), .ZN(n3511) );
  NAND2_X1 U4066 ( .A1(n4428), .A2(n4432), .ZN(n5153) );
  NAND2_X1 U4067 ( .A1(n5148), .A2(n5153), .ZN(n3513) );
  NAND2_X1 U4068 ( .A1(n4590), .A2(n5158), .ZN(n3512) );
  AND2_X1 U4069 ( .A1(n5155), .A2(n5192), .ZN(n3514) );
  XOR2_X1 U4070 ( .A(n3561), .B(n4537), .Z(n5214) );
  NAND2_X1 U4071 ( .A1(n5214), .A2(n4935), .ZN(n3520) );
  NOR2_X1 U4072 ( .A1(n4217), .A2(n4218), .ZN(n5151) );
  INV_X1 U4073 ( .A(n3564), .ZN(n3515) );
  AOI211_X1 U4074 ( .C1(n3562), .C2(n5183), .A(n5264), .B(n3515), .ZN(n5213)
         );
  INV_X1 U4075 ( .A(n5202), .ZN(n5114) );
  INV_X1 U4076 ( .A(n3550), .ZN(n3516) );
  OAI22_X1 U4077 ( .A1(n5208), .A2(n3517), .B1(n3516), .B2(n5210), .ZN(n3518)
         );
  AOI21_X1 U4078 ( .B1(n5213), .B2(n4943), .A(n3518), .ZN(n3519) );
  OAI211_X1 U4079 ( .C1(n3521), .C2(n5330), .A(n3520), .B(n3519), .ZN(U3284)
         );
  INV_X1 U4080 ( .A(n3522), .ZN(n3523) );
  AOI21_X1 U4081 ( .B1(n3525), .B2(n3524), .A(n3523), .ZN(n3530) );
  AOI22_X1 U4082 ( .A1(n4399), .A2(n4590), .B1(n5192), .B2(n5276), .ZN(n3529)
         );
  NOR2_X1 U4083 ( .A1(n5287), .A2(n5211), .ZN(n3526) );
  AOI211_X1 U4084 ( .C1(n4414), .C2(n4589), .A(n3527), .B(n3526), .ZN(n3528)
         );
  OAI211_X1 U4085 ( .C1(n3530), .C2(n4417), .A(n3529), .B(n3528), .ZN(U3224)
         );
  NOR2_X1 U4086 ( .A1(n3532), .A2(n3531), .ZN(n3534) );
  INV_X1 U4087 ( .A(REG2_REG_9__SCAN_IN), .ZN(n3597) );
  AOI22_X1 U4088 ( .A1(n5051), .A2(n3597), .B1(REG2_REG_9__SCAN_IN), .B2(n3614), .ZN(n3535) );
  AOI211_X1 U4089 ( .C1(n2540), .C2(n3535), .A(n3617), .B(n5090), .ZN(n3545)
         );
  NAND2_X1 U4090 ( .A1(n5052), .A2(n3536), .ZN(n3538) );
  INV_X1 U4091 ( .A(REG1_REG_9__SCAN_IN), .ZN(n3539) );
  MUX2_X1 U4092 ( .A(REG1_REG_9__SCAN_IN), .B(n3539), .S(n5051), .Z(n3540) );
  OAI211_X1 U4093 ( .C1(n3541), .C2(n3540), .A(n3613), .B(n5099), .ZN(n3543)
         );
  AND2_X1 U4094 ( .A1(U3149), .A2(REG3_REG_9__SCAN_IN), .ZN(n3630) );
  AOI21_X1 U4095 ( .B1(n5088), .B2(ADDR_REG_9__SCAN_IN), .A(n3630), .ZN(n3542)
         );
  OAI211_X1 U4096 ( .C1(n5089), .C2(n3614), .A(n3543), .B(n3542), .ZN(n3544)
         );
  OR2_X1 U4097 ( .A1(n3545), .A2(n3544), .ZN(U3249) );
  XOR2_X1 U4098 ( .A(n3547), .B(n3546), .Z(n3553) );
  AOI22_X1 U4099 ( .A1(n4399), .A2(n5155), .B1(n3562), .B2(n5276), .ZN(n3552)
         );
  INV_X1 U4100 ( .A(n5287), .ZN(n4345) );
  NOR2_X1 U4101 ( .A1(n5271), .A2(n3555), .ZN(n3548) );
  AOI211_X1 U4102 ( .C1(n4345), .C2(n3550), .A(n3549), .B(n3548), .ZN(n3551)
         );
  OAI211_X1 U4103 ( .C1(n3553), .C2(n4417), .A(n3552), .B(n3551), .ZN(U3236)
         );
  NAND2_X1 U4104 ( .A1(n3555), .A2(n4255), .ZN(n4434) );
  NAND2_X1 U4105 ( .A1(n4588), .A2(n3559), .ZN(n4437) );
  NAND2_X1 U4106 ( .A1(n4434), .A2(n4437), .ZN(n4548) );
  XNOR2_X1 U4107 ( .A(n3574), .B(n4548), .ZN(n3556) );
  NAND2_X1 U4108 ( .A1(n3556), .A2(n5108), .ZN(n3558) );
  AOI22_X1 U4109 ( .A1(n5157), .A2(n4589), .B1(n4587), .B2(n5154), .ZN(n3557)
         );
  OAI211_X1 U4110 ( .C1(n5319), .C2(n3559), .A(n3558), .B(n3557), .ZN(n5217)
         );
  INV_X1 U4111 ( .A(n5217), .ZN(n3569) );
  NOR2_X1 U4112 ( .A1(n4589), .A2(n3562), .ZN(n3560) );
  NAND2_X1 U4113 ( .A1(n4589), .A2(n3562), .ZN(n3563) );
  XOR2_X1 U4114 ( .A(n4548), .B(n3571), .Z(n5219) );
  NAND2_X1 U4115 ( .A1(n5219), .A2(n4935), .ZN(n3568) );
  AOI211_X1 U4116 ( .C1(n4255), .C2(n3564), .A(n5264), .B(n2538), .ZN(n5218)
         );
  INV_X1 U4117 ( .A(REG2_REG_7__SCAN_IN), .ZN(n3565) );
  OAI22_X1 U4118 ( .A1(n5208), .A2(n3565), .B1(n4256), .B2(n5210), .ZN(n3566)
         );
  AOI21_X1 U4119 ( .B1(n5218), .B2(n4943), .A(n3566), .ZN(n3567) );
  OAI211_X1 U4120 ( .C1(n5330), .C2(n3569), .A(n3568), .B(n3567), .ZN(U3283)
         );
  AND2_X1 U4121 ( .A1(n4588), .A2(n4255), .ZN(n3570) );
  AOI21_X2 U4122 ( .B1(n3571), .B2(n4548), .A(n3570), .ZN(n3593) );
  NAND2_X1 U4123 ( .A1(n4587), .A2(n3605), .ZN(n3592) );
  INV_X1 U4124 ( .A(n3592), .ZN(n3572) );
  NOR2_X1 U4125 ( .A1(n4587), .A2(n3605), .ZN(n3591) );
  OR2_X1 U4126 ( .A1(n3572), .A2(n3591), .ZN(n4547) );
  XNOR2_X1 U4127 ( .A(n3593), .B(n4547), .ZN(n5222) );
  INV_X1 U4128 ( .A(n4437), .ZN(n3573) );
  XNOR2_X1 U4129 ( .A(n3586), .B(n4547), .ZN(n3577) );
  AOI22_X1 U4130 ( .A1(n5154), .A2(n4586), .B1(n4588), .B2(n5157), .ZN(n3575)
         );
  OAI21_X1 U4131 ( .B1(n3585), .B2(n5319), .A(n3575), .ZN(n3576) );
  AOI21_X1 U4132 ( .B1(n3577), .B2(n5108), .A(n3576), .ZN(n3578) );
  OAI21_X1 U4133 ( .B1(n5222), .B2(n4968), .A(n3578), .ZN(n5223) );
  NAND2_X1 U4134 ( .A1(n5223), .A2(n5208), .ZN(n3584) );
  NOR2_X1 U4135 ( .A1(n2538), .A2(n3585), .ZN(n3579) );
  INV_X1 U4136 ( .A(n3607), .ZN(n3580) );
  OAI22_X1 U4137 ( .A1(n5208), .A2(n3581), .B1(n3580), .B2(n5210), .ZN(n3582)
         );
  AOI21_X1 U4138 ( .B1(n2539), .B2(n4943), .A(n3582), .ZN(n3583) );
  OAI211_X1 U4139 ( .C1(n5222), .C2(n4795), .A(n3584), .B(n3583), .ZN(U3282)
         );
  NAND2_X1 U4140 ( .A1(n4587), .A2(n3585), .ZN(n4436) );
  NOR2_X1 U4141 ( .A1(n4587), .A2(n3585), .ZN(n4439) );
  INV_X1 U4142 ( .A(n3640), .ZN(n3638) );
  AND2_X1 U4143 ( .A1(n4586), .A2(n3638), .ZN(n3636) );
  INV_X1 U4144 ( .A(n3636), .ZN(n3587) );
  NAND2_X1 U4145 ( .A1(n3643), .A2(n3640), .ZN(n3635) );
  NAND2_X1 U4146 ( .A1(n3587), .A2(n3635), .ZN(n3594) );
  INV_X1 U4147 ( .A(n3594), .ZN(n4550) );
  XNOR2_X1 U4148 ( .A(n3639), .B(n4550), .ZN(n3588) );
  NAND2_X1 U4149 ( .A1(n3588), .A2(n5108), .ZN(n3590) );
  AOI22_X1 U4150 ( .A1(n4585), .A2(n5154), .B1(n5157), .B2(n4587), .ZN(n3589)
         );
  OAI211_X1 U4151 ( .C1(n5319), .C2(n3640), .A(n3590), .B(n3589), .ZN(n5230)
         );
  INV_X1 U4152 ( .A(n5230), .ZN(n3601) );
  XNOR2_X1 U4153 ( .A(n3637), .B(n3594), .ZN(n5232) );
  NAND2_X1 U4154 ( .A1(n3595), .A2(n3640), .ZN(n3648) );
  OAI21_X1 U4155 ( .B1(n3595), .B2(n3640), .A(n3648), .ZN(n5229) );
  NOR2_X1 U4156 ( .A1(n5229), .A2(n4904), .ZN(n3599) );
  INV_X1 U4157 ( .A(n3631), .ZN(n3596) );
  OAI22_X1 U4158 ( .A1(n5208), .A2(n3597), .B1(n3596), .B2(n5210), .ZN(n3598)
         );
  AOI211_X1 U4159 ( .C1(n5232), .C2(n4935), .A(n3599), .B(n3598), .ZN(n3600)
         );
  OAI21_X1 U4160 ( .B1(n5330), .B2(n3601), .A(n3600), .ZN(U3281) );
  OAI21_X1 U4161 ( .B1(n3604), .B2(n3603), .A(n3602), .ZN(n3611) );
  AOI22_X1 U4162 ( .A1(n4410), .A2(n4588), .B1(n3605), .B2(n5276), .ZN(n3609)
         );
  AOI21_X1 U4163 ( .B1(n4345), .B2(n3607), .A(n3606), .ZN(n3608) );
  OAI211_X1 U4164 ( .C1(n5271), .C2(n3643), .A(n3609), .B(n3608), .ZN(n3610)
         );
  AOI21_X1 U4165 ( .B1(n3611), .B2(n5282), .A(n3610), .ZN(n3612) );
  INV_X1 U4166 ( .A(n3612), .ZN(U3218) );
  XOR2_X1 U4167 ( .A(REG1_REG_10__SCAN_IN), .B(n3659), .Z(n3625) );
  INV_X1 U4168 ( .A(n5050), .ZN(n3618) );
  NOR2_X1 U4169 ( .A1(n3746), .A2(STATE_REG_SCAN_IN), .ZN(n4283) );
  AOI21_X1 U4170 ( .B1(n5088), .B2(ADDR_REG_10__SCAN_IN), .A(n4283), .ZN(n3615) );
  OAI21_X1 U4171 ( .B1(n3618), .B2(n5089), .A(n3615), .ZN(n3624) );
  INV_X1 U4172 ( .A(REG2_REG_10__SCAN_IN), .ZN(n3622) );
  NOR2_X1 U4173 ( .A1(n3617), .A2(n3616), .ZN(n3619) );
  NAND2_X1 U4174 ( .A1(n3619), .A2(n3618), .ZN(n3620) );
  AOI211_X1 U4175 ( .C1(n3622), .C2(n3621), .A(n3654), .B(n5090), .ZN(n3623)
         );
  AOI211_X1 U4176 ( .C1(n5099), .C2(n3625), .A(n3624), .B(n3623), .ZN(n3626)
         );
  INV_X1 U4177 ( .A(n3626), .ZN(U3250) );
  XOR2_X1 U4178 ( .A(n3628), .B(n3627), .Z(n3634) );
  AOI22_X1 U4179 ( .A1(n4399), .A2(n4587), .B1(n3638), .B2(n5276), .ZN(n3633)
         );
  NOR2_X1 U4180 ( .A1(n5271), .A2(n3677), .ZN(n3629) );
  AOI211_X1 U4181 ( .C1(n4345), .C2(n3631), .A(n3630), .B(n3629), .ZN(n3632)
         );
  OAI211_X1 U4182 ( .C1(n3634), .C2(n4417), .A(n3633), .B(n3632), .ZN(U3228)
         );
  NAND2_X1 U4183 ( .A1(n3677), .A2(n4282), .ZN(n4454) );
  NAND2_X1 U4184 ( .A1(n4585), .A2(n3669), .ZN(n4444) );
  XOR2_X1 U4185 ( .A(n3670), .B(n4533), .Z(n5238) );
  INV_X1 U4186 ( .A(n5238), .ZN(n3653) );
  NAND2_X1 U4187 ( .A1(n3643), .A2(n3638), .ZN(n4438) );
  NAND2_X1 U4188 ( .A1(n3639), .A2(n4438), .ZN(n3641) );
  NAND2_X1 U4189 ( .A1(n4586), .A2(n3640), .ZN(n4452) );
  NAND2_X1 U4190 ( .A1(n3641), .A2(n4452), .ZN(n3642) );
  OAI211_X1 U4191 ( .C1(n3642), .C2(n4533), .A(n3675), .B(n5108), .ZN(n3646)
         );
  OAI22_X1 U4192 ( .A1(n3643), .A2(n5186), .B1(n4102), .B2(n5188), .ZN(n3644)
         );
  INV_X1 U4193 ( .A(n3644), .ZN(n3645) );
  OAI211_X1 U4194 ( .C1(n5319), .C2(n3669), .A(n3646), .B(n3645), .ZN(n5236)
         );
  INV_X1 U4195 ( .A(n3648), .ZN(n3647) );
  NOR2_X1 U4196 ( .A1(n3647), .A2(n3669), .ZN(n5235) );
  NOR3_X1 U4197 ( .A1(n5235), .A2(n2589), .A3(n4904), .ZN(n3651) );
  INV_X1 U4198 ( .A(n3649), .ZN(n4285) );
  OAI22_X1 U4199 ( .A1(n5208), .A2(n3622), .B1(n4285), .B2(n5210), .ZN(n3650)
         );
  AOI211_X1 U4200 ( .C1(n5236), .C2(n5208), .A(n3651), .B(n3650), .ZN(n3652)
         );
  OAI21_X1 U4201 ( .B1(n3653), .B2(n4962), .A(n3652), .ZN(U3280) );
  NAND2_X1 U4202 ( .A1(n5049), .A2(REG2_REG_11__SCAN_IN), .ZN(n3655) );
  OAI21_X1 U4203 ( .B1(n5049), .B2(REG2_REG_11__SCAN_IN), .A(n3655), .ZN(n3656) );
  AOI211_X1 U4204 ( .C1(n2543), .C2(n3656), .A(n4171), .B(n5090), .ZN(n3668)
         );
  INV_X1 U4205 ( .A(n5049), .ZN(n3666) );
  NAND2_X1 U4206 ( .A1(U3149), .A2(REG3_REG_11__SCAN_IN), .ZN(n3688) );
  INV_X1 U4207 ( .A(n3688), .ZN(n3657) );
  AOI21_X1 U4208 ( .B1(n5088), .B2(ADDR_REG_11__SCAN_IN), .A(n3657), .ZN(n3665) );
  AOI22_X1 U4209 ( .A1(n3659), .A2(REG1_REG_10__SCAN_IN), .B1(n5050), .B2(
        n3658), .ZN(n3660) );
  INV_X1 U4210 ( .A(REG1_REG_11__SCAN_IN), .ZN(n3661) );
  MUX2_X1 U4211 ( .A(REG1_REG_11__SCAN_IN), .B(n3661), .S(n5049), .Z(n3662) );
  OAI211_X1 U4212 ( .C1(n3663), .C2(n3662), .A(n5099), .B(n4174), .ZN(n3664)
         );
  OAI211_X1 U4213 ( .C1(n5089), .C2(n3666), .A(n3665), .B(n3664), .ZN(n3667)
         );
  OR2_X1 U4214 ( .A1(n3668), .A2(n3667), .ZN(U3251) );
  NAND2_X1 U4215 ( .A1(n4102), .A2(n3687), .ZN(n4460) );
  NAND2_X1 U4216 ( .A1(n4584), .A2(n4101), .ZN(n4445) );
  AOI21_X1 U4217 ( .B1(n4535), .B2(n3671), .A(n2541), .ZN(n5243) );
  OAI21_X1 U4218 ( .B1(n2589), .B2(n4101), .A(n4103), .ZN(n5242) );
  INV_X1 U4219 ( .A(n5242), .ZN(n3674) );
  INV_X1 U4220 ( .A(REG2_REG_11__SCAN_IN), .ZN(n3672) );
  OAI22_X1 U4221 ( .A1(n5208), .A2(n3672), .B1(n3689), .B2(n5210), .ZN(n3673)
         );
  AOI21_X1 U4222 ( .B1(n3674), .B2(n5328), .A(n3673), .ZN(n3682) );
  OAI211_X1 U4223 ( .C1(n3676), .C2(n4535), .A(n4096), .B(n5108), .ZN(n3680)
         );
  OAI22_X1 U4224 ( .A1(n4139), .A2(n5188), .B1(n3677), .B2(n5186), .ZN(n3678)
         );
  INV_X1 U4225 ( .A(n3678), .ZN(n3679) );
  OAI211_X1 U4226 ( .C1(n5319), .C2(n4101), .A(n3680), .B(n3679), .ZN(n5244)
         );
  NAND2_X1 U4227 ( .A1(n5244), .A2(n5208), .ZN(n3681) );
  OAI211_X1 U4228 ( .C1(n5243), .C2(n4962), .A(n3682), .B(n3681), .ZN(U3279)
         );
  XOR2_X1 U4229 ( .A(n3684), .B(n3683), .Z(n3685) );
  XNOR2_X1 U4230 ( .A(n3686), .B(n3685), .ZN(n3693) );
  AOI22_X1 U4231 ( .A1(n4399), .A2(n4585), .B1(n3687), .B2(n5276), .ZN(n3692)
         );
  OAI21_X1 U4232 ( .B1(n5287), .B2(n3689), .A(n3688), .ZN(n3690) );
  AOI21_X1 U4233 ( .B1(n4414), .B2(n4583), .A(n3690), .ZN(n3691) );
  OAI211_X1 U4234 ( .C1(n3693), .C2(n4417), .A(n3692), .B(n3691), .ZN(U3233)
         );
  XOR2_X1 U4235 ( .A(DATAI_29_), .B(keyinput_2), .Z(n3696) );
  XNOR2_X1 U4236 ( .A(DATAI_30_), .B(keyinput_1), .ZN(n3695) );
  XNOR2_X1 U4237 ( .A(DATAI_31_), .B(keyinput_0), .ZN(n3694) );
  NOR3_X1 U4238 ( .A1(n3696), .A2(n3695), .A3(n3694), .ZN(n3700) );
  XOR2_X1 U4239 ( .A(DATAI_28_), .B(keyinput_3), .Z(n3699) );
  XOR2_X1 U4240 ( .A(DATAI_27_), .B(keyinput_4), .Z(n3698) );
  XNOR2_X1 U4241 ( .A(DATAI_26_), .B(keyinput_5), .ZN(n3697) );
  OAI211_X1 U4242 ( .C1(n3700), .C2(n3699), .A(n3698), .B(n3697), .ZN(n3706)
         );
  XOR2_X1 U4243 ( .A(DATAI_25_), .B(keyinput_6), .Z(n3705) );
  XOR2_X1 U4244 ( .A(DATAI_22_), .B(keyinput_9), .Z(n3703) );
  XNOR2_X1 U4245 ( .A(DATAI_23_), .B(keyinput_8), .ZN(n3702) );
  XNOR2_X1 U4246 ( .A(DATAI_24_), .B(keyinput_7), .ZN(n3701) );
  NAND3_X1 U4247 ( .A1(n3703), .A2(n3702), .A3(n3701), .ZN(n3704) );
  AOI21_X1 U4248 ( .B1(n3706), .B2(n3705), .A(n3704), .ZN(n3718) );
  XNOR2_X1 U4249 ( .A(DATAI_21_), .B(keyinput_10), .ZN(n3717) );
  XNOR2_X1 U4250 ( .A(n3905), .B(keyinput_16), .ZN(n3711) );
  XOR2_X1 U4251 ( .A(DATAI_20_), .B(keyinput_11), .Z(n3710) );
  XNOR2_X1 U4252 ( .A(n3707), .B(keyinput_12), .ZN(n3709) );
  XNOR2_X1 U4253 ( .A(n3904), .B(keyinput_14), .ZN(n3708) );
  NAND4_X1 U4254 ( .A1(n3711), .A2(n3710), .A3(n3709), .A4(n3708), .ZN(n3715)
         );
  XNOR2_X1 U4255 ( .A(n3910), .B(keyinput_13), .ZN(n3714) );
  XNOR2_X1 U4256 ( .A(DATAI_14_), .B(keyinput_17), .ZN(n3713) );
  XNOR2_X1 U4257 ( .A(DATAI_16_), .B(keyinput_15), .ZN(n3712) );
  NOR4_X1 U4258 ( .A1(n3715), .A2(n3714), .A3(n3713), .A4(n3712), .ZN(n3716)
         );
  OAI21_X1 U4259 ( .B1(n3718), .B2(n3717), .A(n3716), .ZN(n3722) );
  XNOR2_X1 U4260 ( .A(n3719), .B(keyinput_18), .ZN(n3721) );
  XNOR2_X1 U4261 ( .A(DATAI_12_), .B(keyinput_19), .ZN(n3720) );
  AOI21_X1 U4262 ( .B1(n3722), .B2(n3721), .A(n3720), .ZN(n3728) );
  XOR2_X1 U4263 ( .A(DATAI_11_), .B(keyinput_20), .Z(n3727) );
  XOR2_X1 U4264 ( .A(DATAI_10_), .B(keyinput_21), .Z(n3725) );
  XNOR2_X1 U4265 ( .A(n3921), .B(keyinput_22), .ZN(n3724) );
  XNOR2_X1 U4266 ( .A(DATAI_8_), .B(keyinput_23), .ZN(n3723) );
  NOR3_X1 U4267 ( .A1(n3725), .A2(n3724), .A3(n3723), .ZN(n3726) );
  OAI21_X1 U4268 ( .B1(n3728), .B2(n3727), .A(n3726), .ZN(n3732) );
  XOR2_X1 U4269 ( .A(DATAI_7_), .B(keyinput_24), .Z(n3731) );
  XOR2_X1 U4270 ( .A(DATAI_5_), .B(keyinput_26), .Z(n3730) );
  XOR2_X1 U4271 ( .A(DATAI_6_), .B(keyinput_25), .Z(n3729) );
  AOI211_X1 U4272 ( .C1(n3732), .C2(n3731), .A(n3730), .B(n3729), .ZN(n3735)
         );
  XOR2_X1 U4273 ( .A(DATAI_4_), .B(keyinput_27), .Z(n3734) );
  XOR2_X1 U4274 ( .A(DATAI_3_), .B(keyinput_28), .Z(n3733) );
  NOR3_X1 U4275 ( .A1(n3735), .A2(n3734), .A3(n3733), .ZN(n3738) );
  XOR2_X1 U4276 ( .A(DATAI_1_), .B(keyinput_30), .Z(n3737) );
  XNOR2_X1 U4277 ( .A(DATAI_2_), .B(keyinput_29), .ZN(n3736) );
  NOR3_X1 U4278 ( .A1(n3738), .A2(n3737), .A3(n3736), .ZN(n3741) );
  XOR2_X1 U4279 ( .A(DATAI_0_), .B(keyinput_31), .Z(n3740) );
  XNOR2_X1 U4280 ( .A(U3149), .B(keyinput_32), .ZN(n3739) );
  NOR3_X1 U4281 ( .A1(n3741), .A2(n3740), .A3(n3739), .ZN(n3745) );
  XNOR2_X1 U4282 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput_33), .ZN(n3744) );
  XNOR2_X1 U4283 ( .A(n3742), .B(keyinput_34), .ZN(n3743) );
  OAI21_X1 U4284 ( .B1(n3745), .B2(n3744), .A(n3743), .ZN(n3753) );
  XNOR2_X1 U4285 ( .A(n3944), .B(keyinput_38), .ZN(n3750) );
  XOR2_X1 U4286 ( .A(REG3_REG_23__SCAN_IN), .B(keyinput_36), .Z(n3749) );
  INV_X1 U4287 ( .A(REG3_REG_14__SCAN_IN), .ZN(n4184) );
  XNOR2_X1 U4288 ( .A(n4184), .B(keyinput_35), .ZN(n3748) );
  XNOR2_X1 U4289 ( .A(n3746), .B(keyinput_37), .ZN(n3747) );
  NOR4_X1 U4290 ( .A1(n3750), .A2(n3749), .A3(n3748), .A4(n3747), .ZN(n3752)
         );
  XOR2_X1 U4291 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput_39), .Z(n3751) );
  AOI21_X1 U4292 ( .B1(n3753), .B2(n3752), .A(n3751), .ZN(n3756) );
  XOR2_X1 U4293 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput_41), .Z(n3755) );
  XNOR2_X1 U4294 ( .A(REG3_REG_28__SCAN_IN), .B(keyinput_40), .ZN(n3754) );
  NOR3_X1 U4295 ( .A1(n3756), .A2(n3755), .A3(n3754), .ZN(n3759) );
  XNOR2_X1 U4296 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_42), .ZN(n3758) );
  XNOR2_X1 U4297 ( .A(REG3_REG_21__SCAN_IN), .B(keyinput_43), .ZN(n3757) );
  OAI21_X1 U4298 ( .B1(n3759), .B2(n3758), .A(n3757), .ZN(n3762) );
  INV_X1 U4299 ( .A(REG3_REG_12__SCAN_IN), .ZN(n4114) );
  XNOR2_X1 U4300 ( .A(n4114), .B(keyinput_44), .ZN(n3761) );
  XOR2_X1 U4301 ( .A(REG3_REG_25__SCAN_IN), .B(keyinput_45), .Z(n3760) );
  AOI21_X1 U4302 ( .B1(n3762), .B2(n3761), .A(n3760), .ZN(n3769) );
  INV_X1 U4303 ( .A(REG3_REG_16__SCAN_IN), .ZN(n4333) );
  XNOR2_X1 U4304 ( .A(n4333), .B(keyinput_46), .ZN(n3768) );
  XOR2_X1 U4305 ( .A(REG3_REG_24__SCAN_IN), .B(keyinput_49), .Z(n3766) );
  XNOR2_X1 U4306 ( .A(n4367), .B(keyinput_50), .ZN(n3765) );
  XNOR2_X1 U4307 ( .A(REG3_REG_5__SCAN_IN), .B(keyinput_47), .ZN(n3764) );
  XNOR2_X1 U4308 ( .A(REG3_REG_17__SCAN_IN), .B(keyinput_48), .ZN(n3763) );
  NOR4_X1 U4309 ( .A1(n3766), .A2(n3765), .A3(n3764), .A4(n3763), .ZN(n3767)
         );
  OAI21_X1 U4310 ( .B1(n3769), .B2(n3768), .A(n3767), .ZN(n3773) );
  XOR2_X1 U4311 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_52), .Z(n3772) );
  XNOR2_X1 U4312 ( .A(n3770), .B(keyinput_51), .ZN(n3771) );
  NAND3_X1 U4313 ( .A1(n3773), .A2(n3772), .A3(n3771), .ZN(n3776) );
  XNOR2_X1 U4314 ( .A(REG3_REG_20__SCAN_IN), .B(keyinput_53), .ZN(n3775) );
  XNOR2_X1 U4315 ( .A(REG3_REG_13__SCAN_IN), .B(keyinput_54), .ZN(n3774) );
  NAND3_X1 U4316 ( .A1(n3776), .A2(n3775), .A3(n3774), .ZN(n3779) );
  XOR2_X1 U4317 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_55), .Z(n3778) );
  XOR2_X1 U4318 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_56), .Z(n3777) );
  NAND3_X1 U4319 ( .A1(n3779), .A2(n3778), .A3(n3777), .ZN(n3786) );
  XNOR2_X1 U4320 ( .A(n3780), .B(keyinput_57), .ZN(n3785) );
  XNOR2_X1 U4321 ( .A(n3980), .B(keyinput_59), .ZN(n3783) );
  XNOR2_X1 U4322 ( .A(n3977), .B(keyinput_58), .ZN(n3782) );
  XNOR2_X1 U4323 ( .A(IR_REG_5__SCAN_IN), .B(keyinput_60), .ZN(n3781) );
  NAND3_X1 U4324 ( .A1(n3783), .A2(n3782), .A3(n3781), .ZN(n3784) );
  AOI21_X1 U4325 ( .B1(n3786), .B2(n3785), .A(n3784), .ZN(n3791) );
  XNOR2_X1 U4326 ( .A(n3787), .B(keyinput_61), .ZN(n3790) );
  XNOR2_X1 U4327 ( .A(IR_REG_7__SCAN_IN), .B(keyinput_62), .ZN(n3789) );
  XNOR2_X1 U4328 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_63), .ZN(n3788) );
  NOR4_X1 U4329 ( .A1(n3791), .A2(n3790), .A3(n3789), .A4(n3788), .ZN(n3794)
         );
  XOR2_X1 U4330 ( .A(IR_REG_10__SCAN_IN), .B(keyinput_65), .Z(n3793) );
  XNOR2_X1 U4331 ( .A(IR_REG_9__SCAN_IN), .B(keyinput_64), .ZN(n3792) );
  NOR3_X1 U4332 ( .A1(n3794), .A2(n3793), .A3(n3792), .ZN(n3798) );
  XNOR2_X1 U4333 ( .A(n3795), .B(keyinput_66), .ZN(n3797) );
  XOR2_X1 U4334 ( .A(IR_REG_12__SCAN_IN), .B(keyinput_67), .Z(n3796) );
  NOR3_X1 U4335 ( .A1(n3798), .A2(n3797), .A3(n3796), .ZN(n3802) );
  XNOR2_X1 U4336 ( .A(n2754), .B(keyinput_68), .ZN(n3801) );
  XNOR2_X1 U4337 ( .A(n3996), .B(keyinput_69), .ZN(n3800) );
  XNOR2_X1 U4338 ( .A(IR_REG_15__SCAN_IN), .B(keyinput_70), .ZN(n3799) );
  OAI211_X1 U4339 ( .C1(n3802), .C2(n3801), .A(n3800), .B(n3799), .ZN(n3806)
         );
  XOR2_X1 U4340 ( .A(IR_REG_16__SCAN_IN), .B(keyinput_71), .Z(n3805) );
  XNOR2_X1 U4341 ( .A(n3803), .B(keyinput_72), .ZN(n3804) );
  NAND3_X1 U4342 ( .A1(n3806), .A2(n3805), .A3(n3804), .ZN(n3814) );
  XOR2_X1 U4343 ( .A(IR_REG_18__SCAN_IN), .B(keyinput_73), .Z(n3813) );
  XNOR2_X1 U4344 ( .A(n3807), .B(keyinput_75), .ZN(n3811) );
  XNOR2_X1 U4345 ( .A(n3808), .B(keyinput_76), .ZN(n3810) );
  XNOR2_X1 U4346 ( .A(IR_REG_19__SCAN_IN), .B(keyinput_74), .ZN(n3809) );
  NAND3_X1 U4347 ( .A1(n3811), .A2(n3810), .A3(n3809), .ZN(n3812) );
  AOI21_X1 U4348 ( .B1(n3814), .B2(n3813), .A(n3812), .ZN(n3823) );
  XNOR2_X1 U4349 ( .A(n2777), .B(keyinput_78), .ZN(n3819) );
  XNOR2_X1 U4350 ( .A(n4011), .B(keyinput_79), .ZN(n3818) );
  XNOR2_X1 U4351 ( .A(n3815), .B(keyinput_77), .ZN(n3817) );
  XNOR2_X1 U4352 ( .A(IR_REG_25__SCAN_IN), .B(keyinput_80), .ZN(n3816) );
  NAND4_X1 U4353 ( .A1(n3819), .A2(n3818), .A3(n3817), .A4(n3816), .ZN(n3822)
         );
  XNOR2_X1 U4354 ( .A(IR_REG_27__SCAN_IN), .B(keyinput_82), .ZN(n3821) );
  XNOR2_X1 U4355 ( .A(IR_REG_26__SCAN_IN), .B(keyinput_81), .ZN(n3820) );
  OAI211_X1 U4356 ( .C1(n3823), .C2(n3822), .A(n3821), .B(n3820), .ZN(n3826)
         );
  XNOR2_X1 U4357 ( .A(IR_REG_28__SCAN_IN), .B(keyinput_83), .ZN(n3825) );
  XOR2_X1 U4358 ( .A(IR_REG_29__SCAN_IN), .B(keyinput_84), .Z(n3824) );
  AOI21_X1 U4359 ( .B1(n3826), .B2(n3825), .A(n3824), .ZN(n3830) );
  XNOR2_X1 U4360 ( .A(n3827), .B(keyinput_85), .ZN(n3829) );
  XNOR2_X1 U4361 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_86), .ZN(n3828) );
  OAI21_X1 U4362 ( .B1(n3830), .B2(n3829), .A(n3828), .ZN(n3832) );
  XNOR2_X1 U4363 ( .A(D_REG_0__SCAN_IN), .B(keyinput_87), .ZN(n3831) );
  NAND2_X1 U4364 ( .A1(n3832), .A2(n3831), .ZN(n3836) );
  XOR2_X1 U4365 ( .A(D_REG_3__SCAN_IN), .B(keyinput_90), .Z(n3835) );
  XNOR2_X1 U4366 ( .A(D_REG_1__SCAN_IN), .B(keyinput_88), .ZN(n3834) );
  XNOR2_X1 U4367 ( .A(D_REG_2__SCAN_IN), .B(keyinput_89), .ZN(n3833) );
  NAND4_X1 U4368 ( .A1(n3836), .A2(n3835), .A3(n3834), .A4(n3833), .ZN(n3839)
         );
  INV_X1 U4369 ( .A(D_REG_4__SCAN_IN), .ZN(n5059) );
  XNOR2_X1 U4370 ( .A(n5059), .B(keyinput_91), .ZN(n3838) );
  XNOR2_X1 U4371 ( .A(D_REG_5__SCAN_IN), .B(keyinput_92), .ZN(n3837) );
  AOI21_X1 U4372 ( .B1(n3839), .B2(n3838), .A(n3837), .ZN(n3842) );
  XNOR2_X1 U4373 ( .A(D_REG_6__SCAN_IN), .B(keyinput_93), .ZN(n3841) );
  INV_X1 U4374 ( .A(D_REG_7__SCAN_IN), .ZN(n5062) );
  XNOR2_X1 U4375 ( .A(n5062), .B(keyinput_94), .ZN(n3840) );
  OAI21_X1 U4376 ( .B1(n3842), .B2(n3841), .A(n3840), .ZN(n3845) );
  INV_X1 U4377 ( .A(D_REG_9__SCAN_IN), .ZN(n5064) );
  XNOR2_X1 U4378 ( .A(n5064), .B(keyinput_96), .ZN(n3844) );
  XNOR2_X1 U4379 ( .A(D_REG_8__SCAN_IN), .B(keyinput_95), .ZN(n3843) );
  NAND3_X1 U4380 ( .A1(n3845), .A2(n3844), .A3(n3843), .ZN(n3848) );
  XNOR2_X1 U4381 ( .A(D_REG_10__SCAN_IN), .B(keyinput_97), .ZN(n3847) );
  INV_X1 U4382 ( .A(D_REG_11__SCAN_IN), .ZN(n5066) );
  XNOR2_X1 U4383 ( .A(n5066), .B(keyinput_98), .ZN(n3846) );
  AOI21_X1 U4384 ( .B1(n3848), .B2(n3847), .A(n3846), .ZN(n3851) );
  INV_X1 U4385 ( .A(D_REG_13__SCAN_IN), .ZN(n5068) );
  XNOR2_X1 U4386 ( .A(n5068), .B(keyinput_100), .ZN(n3850) );
  XNOR2_X1 U4387 ( .A(D_REG_12__SCAN_IN), .B(keyinput_99), .ZN(n3849) );
  NOR3_X1 U4388 ( .A1(n3851), .A2(n3850), .A3(n3849), .ZN(n3857) );
  INV_X1 U4389 ( .A(D_REG_14__SCAN_IN), .ZN(n5069) );
  XNOR2_X1 U4390 ( .A(n5069), .B(keyinput_101), .ZN(n3856) );
  INV_X1 U4391 ( .A(D_REG_15__SCAN_IN), .ZN(n5070) );
  XNOR2_X1 U4392 ( .A(n5070), .B(keyinput_102), .ZN(n3854) );
  INV_X1 U4393 ( .A(D_REG_17__SCAN_IN), .ZN(n5072) );
  XNOR2_X1 U4394 ( .A(n5072), .B(keyinput_104), .ZN(n3853) );
  INV_X1 U4395 ( .A(D_REG_16__SCAN_IN), .ZN(n5071) );
  XNOR2_X1 U4396 ( .A(n5071), .B(keyinput_103), .ZN(n3852) );
  NOR3_X1 U4397 ( .A1(n3854), .A2(n3853), .A3(n3852), .ZN(n3855) );
  OAI21_X1 U4398 ( .B1(n3857), .B2(n3856), .A(n3855), .ZN(n3860) );
  XNOR2_X1 U4399 ( .A(D_REG_18__SCAN_IN), .B(keyinput_105), .ZN(n3859) );
  INV_X1 U4400 ( .A(D_REG_19__SCAN_IN), .ZN(n5074) );
  XNOR2_X1 U4401 ( .A(n5074), .B(keyinput_106), .ZN(n3858) );
  AOI21_X1 U4402 ( .B1(n3860), .B2(n3859), .A(n3858), .ZN(n3863) );
  XNOR2_X1 U4403 ( .A(D_REG_20__SCAN_IN), .B(keyinput_107), .ZN(n3862) );
  XNOR2_X1 U4404 ( .A(D_REG_21__SCAN_IN), .B(keyinput_108), .ZN(n3861) );
  OAI21_X1 U4405 ( .B1(n3863), .B2(n3862), .A(n3861), .ZN(n3866) );
  INV_X1 U4406 ( .A(D_REG_22__SCAN_IN), .ZN(n5077) );
  XNOR2_X1 U4407 ( .A(n5077), .B(keyinput_109), .ZN(n3865) );
  INV_X1 U4408 ( .A(D_REG_23__SCAN_IN), .ZN(n5078) );
  XNOR2_X1 U4409 ( .A(n5078), .B(keyinput_110), .ZN(n3864) );
  NAND3_X1 U4410 ( .A1(n3866), .A2(n3865), .A3(n3864), .ZN(n3873) );
  INV_X1 U4411 ( .A(D_REG_27__SCAN_IN), .ZN(n5081) );
  XNOR2_X1 U4412 ( .A(n5081), .B(keyinput_114), .ZN(n3870) );
  INV_X1 U4413 ( .A(D_REG_26__SCAN_IN), .ZN(n5080) );
  XNOR2_X1 U4414 ( .A(n5080), .B(keyinput_113), .ZN(n3869) );
  XNOR2_X1 U4415 ( .A(D_REG_24__SCAN_IN), .B(keyinput_111), .ZN(n3868) );
  XNOR2_X1 U4416 ( .A(D_REG_25__SCAN_IN), .B(keyinput_112), .ZN(n3867) );
  NOR4_X1 U4417 ( .A1(n3870), .A2(n3869), .A3(n3868), .A4(n3867), .ZN(n3872)
         );
  INV_X1 U4418 ( .A(D_REG_28__SCAN_IN), .ZN(n5082) );
  XNOR2_X1 U4419 ( .A(n5082), .B(keyinput_115), .ZN(n3871) );
  AOI21_X1 U4420 ( .B1(n3873), .B2(n3872), .A(n3871), .ZN(n3879) );
  XNOR2_X1 U4421 ( .A(D_REG_29__SCAN_IN), .B(keyinput_116), .ZN(n3878) );
  XOR2_X1 U4422 ( .A(REG0_REG_0__SCAN_IN), .B(keyinput_119), .Z(n3876) );
  XNOR2_X1 U4423 ( .A(D_REG_30__SCAN_IN), .B(keyinput_117), .ZN(n3875) );
  XNOR2_X1 U4424 ( .A(D_REG_31__SCAN_IN), .B(keyinput_118), .ZN(n3874) );
  NOR3_X1 U4425 ( .A1(n3876), .A2(n3875), .A3(n3874), .ZN(n3877) );
  OAI21_X1 U4426 ( .B1(n3879), .B2(n3878), .A(n3877), .ZN(n3882) );
  XNOR2_X1 U4427 ( .A(REG0_REG_1__SCAN_IN), .B(keyinput_120), .ZN(n3881) );
  XOR2_X1 U4428 ( .A(REG0_REG_2__SCAN_IN), .B(keyinput_121), .Z(n3880) );
  AOI21_X1 U4429 ( .B1(n3882), .B2(n3881), .A(n3880), .ZN(n3885) );
  XOR2_X1 U4430 ( .A(REG0_REG_4__SCAN_IN), .B(keyinput_123), .Z(n3884) );
  XNOR2_X1 U4431 ( .A(REG0_REG_3__SCAN_IN), .B(keyinput_122), .ZN(n3883) );
  NOR3_X1 U4432 ( .A1(n3885), .A2(n3884), .A3(n3883), .ZN(n3889) );
  XOR2_X1 U4433 ( .A(REG0_REG_5__SCAN_IN), .B(keyinput_124), .Z(n3888) );
  XOR2_X1 U4434 ( .A(REG0_REG_7__SCAN_IN), .B(keyinput_126), .Z(n3887) );
  XNOR2_X1 U4435 ( .A(REG0_REG_6__SCAN_IN), .B(keyinput_125), .ZN(n3886) );
  NOR4_X1 U4436 ( .A1(n3889), .A2(n3888), .A3(n3887), .A4(n3886), .ZN(n4092)
         );
  XNOR2_X1 U4437 ( .A(REG0_REG_8__SCAN_IN), .B(keyinput_127), .ZN(n4091) );
  XOR2_X1 U4438 ( .A(REG0_REG_8__SCAN_IN), .B(keyinput_255), .Z(n4090) );
  XOR2_X1 U4439 ( .A(DATAI_21_), .B(keyinput_138), .Z(n3917) );
  XOR2_X1 U4440 ( .A(DATAI_30_), .B(keyinput_129), .Z(n3892) );
  XOR2_X1 U4441 ( .A(DATAI_31_), .B(keyinput_128), .Z(n3891) );
  XNOR2_X1 U4442 ( .A(DATAI_29_), .B(keyinput_130), .ZN(n3890) );
  NAND3_X1 U4443 ( .A1(n3892), .A2(n3891), .A3(n3890), .ZN(n3896) );
  XNOR2_X1 U4444 ( .A(DATAI_28_), .B(keyinput_131), .ZN(n3895) );
  XNOR2_X1 U4445 ( .A(DATAI_27_), .B(keyinput_132), .ZN(n3894) );
  XOR2_X1 U4446 ( .A(DATAI_26_), .B(keyinput_133), .Z(n3893) );
  AOI211_X1 U4447 ( .C1(n3896), .C2(n3895), .A(n3894), .B(n3893), .ZN(n3902)
         );
  XOR2_X1 U4448 ( .A(DATAI_25_), .B(keyinput_134), .Z(n3901) );
  XOR2_X1 U4449 ( .A(DATAI_24_), .B(keyinput_135), .Z(n3899) );
  XNOR2_X1 U4450 ( .A(DATAI_22_), .B(keyinput_137), .ZN(n3898) );
  XNOR2_X1 U4451 ( .A(DATAI_23_), .B(keyinput_136), .ZN(n3897) );
  NOR3_X1 U4452 ( .A1(n3899), .A2(n3898), .A3(n3897), .ZN(n3900) );
  OAI21_X1 U4453 ( .B1(n3902), .B2(n3901), .A(n3900), .ZN(n3916) );
  XNOR2_X1 U4454 ( .A(n3903), .B(keyinput_143), .ZN(n3909) );
  XOR2_X1 U4455 ( .A(DATAI_14_), .B(keyinput_145), .Z(n3908) );
  XNOR2_X1 U4456 ( .A(n3904), .B(keyinput_142), .ZN(n3907) );
  XNOR2_X1 U4457 ( .A(n3905), .B(keyinput_144), .ZN(n3906) );
  NOR4_X1 U4458 ( .A1(n3909), .A2(n3908), .A3(n3907), .A4(n3906), .ZN(n3914)
         );
  XNOR2_X1 U4459 ( .A(n3910), .B(keyinput_141), .ZN(n3913) );
  XNOR2_X1 U4460 ( .A(DATAI_20_), .B(keyinput_139), .ZN(n3912) );
  XNOR2_X1 U4461 ( .A(DATAI_19_), .B(keyinput_140), .ZN(n3911) );
  NAND4_X1 U4462 ( .A1(n3914), .A2(n3913), .A3(n3912), .A4(n3911), .ZN(n3915)
         );
  AOI21_X1 U4463 ( .B1(n3917), .B2(n3916), .A(n3915), .ZN(n3920) );
  XNOR2_X1 U4464 ( .A(DATAI_13_), .B(keyinput_146), .ZN(n3919) );
  XOR2_X1 U4465 ( .A(DATAI_12_), .B(keyinput_147), .Z(n3918) );
  OAI21_X1 U4466 ( .B1(n3920), .B2(n3919), .A(n3918), .ZN(n3927) );
  XNOR2_X1 U4467 ( .A(DATAI_11_), .B(keyinput_148), .ZN(n3926) );
  XOR2_X1 U4468 ( .A(DATAI_10_), .B(keyinput_149), .Z(n3924) );
  XNOR2_X1 U4469 ( .A(n3921), .B(keyinput_150), .ZN(n3923) );
  XNOR2_X1 U4470 ( .A(DATAI_8_), .B(keyinput_151), .ZN(n3922) );
  NAND3_X1 U4471 ( .A1(n3924), .A2(n3923), .A3(n3922), .ZN(n3925) );
  AOI21_X1 U4472 ( .B1(n3927), .B2(n3926), .A(n3925), .ZN(n3931) );
  XNOR2_X1 U4473 ( .A(DATAI_7_), .B(keyinput_152), .ZN(n3930) );
  XOR2_X1 U4474 ( .A(DATAI_5_), .B(keyinput_154), .Z(n3929) );
  XNOR2_X1 U4475 ( .A(DATAI_6_), .B(keyinput_153), .ZN(n3928) );
  OAI211_X1 U4476 ( .C1(n3931), .C2(n3930), .A(n3929), .B(n3928), .ZN(n3934)
         );
  XNOR2_X1 U4477 ( .A(DATAI_4_), .B(keyinput_155), .ZN(n3933) );
  XNOR2_X1 U4478 ( .A(DATAI_3_), .B(keyinput_156), .ZN(n3932) );
  NAND3_X1 U4479 ( .A1(n3934), .A2(n3933), .A3(n3932), .ZN(n3937) );
  XNOR2_X1 U4480 ( .A(DATAI_2_), .B(keyinput_157), .ZN(n3936) );
  XNOR2_X1 U4481 ( .A(DATAI_1_), .B(keyinput_158), .ZN(n3935) );
  NAND3_X1 U4482 ( .A1(n3937), .A2(n3936), .A3(n3935), .ZN(n3940) );
  XOR2_X1 U4483 ( .A(DATAI_0_), .B(keyinput_159), .Z(n3939) );
  XNOR2_X1 U4484 ( .A(U3149), .B(keyinput_160), .ZN(n3938) );
  NAND3_X1 U4485 ( .A1(n3940), .A2(n3939), .A3(n3938), .ZN(n3943) );
  XNOR2_X1 U4486 ( .A(REG3_REG_7__SCAN_IN), .B(keyinput_161), .ZN(n3942) );
  XNOR2_X1 U4487 ( .A(REG3_REG_27__SCAN_IN), .B(keyinput_162), .ZN(n3941) );
  AOI21_X1 U4488 ( .B1(n3943), .B2(n3942), .A(n3941), .ZN(n3951) );
  XOR2_X1 U4489 ( .A(REG3_REG_23__SCAN_IN), .B(keyinput_164), .Z(n3948) );
  XNOR2_X1 U4490 ( .A(n4184), .B(keyinput_163), .ZN(n3947) );
  XNOR2_X1 U4491 ( .A(n3944), .B(keyinput_166), .ZN(n3946) );
  XNOR2_X1 U4492 ( .A(REG3_REG_10__SCAN_IN), .B(keyinput_165), .ZN(n3945) );
  NAND4_X1 U4493 ( .A1(n3948), .A2(n3947), .A3(n3946), .A4(n3945), .ZN(n3950)
         );
  XOR2_X1 U4494 ( .A(REG3_REG_19__SCAN_IN), .B(keyinput_167), .Z(n3949) );
  OAI21_X1 U4495 ( .B1(n3951), .B2(n3950), .A(n3949), .ZN(n3954) );
  XNOR2_X1 U4496 ( .A(REG3_REG_28__SCAN_IN), .B(keyinput_168), .ZN(n3953) );
  XNOR2_X1 U4497 ( .A(REG3_REG_8__SCAN_IN), .B(keyinput_169), .ZN(n3952) );
  NAND3_X1 U4498 ( .A1(n3954), .A2(n3953), .A3(n3952), .ZN(n3957) );
  XNOR2_X1 U4499 ( .A(REG3_REG_1__SCAN_IN), .B(keyinput_170), .ZN(n3956) );
  XNOR2_X1 U4500 ( .A(REG3_REG_21__SCAN_IN), .B(keyinput_171), .ZN(n3955) );
  AOI21_X1 U4501 ( .B1(n3957), .B2(n3956), .A(n3955), .ZN(n3960) );
  XNOR2_X1 U4502 ( .A(n4114), .B(keyinput_172), .ZN(n3959) );
  XNOR2_X1 U4503 ( .A(REG3_REG_25__SCAN_IN), .B(keyinput_173), .ZN(n3958) );
  OAI21_X1 U4504 ( .B1(n3960), .B2(n3959), .A(n3958), .ZN(n3967) );
  XNOR2_X1 U4505 ( .A(REG3_REG_16__SCAN_IN), .B(keyinput_174), .ZN(n3966) );
  XOR2_X1 U4506 ( .A(REG3_REG_5__SCAN_IN), .B(keyinput_175), .Z(n3964) );
  XNOR2_X1 U4507 ( .A(REG3_REG_24__SCAN_IN), .B(keyinput_177), .ZN(n3963) );
  XNOR2_X1 U4508 ( .A(REG3_REG_4__SCAN_IN), .B(keyinput_178), .ZN(n3962) );
  XNOR2_X1 U4509 ( .A(REG3_REG_17__SCAN_IN), .B(keyinput_176), .ZN(n3961) );
  NAND4_X1 U4510 ( .A1(n3964), .A2(n3963), .A3(n3962), .A4(n3961), .ZN(n3965)
         );
  AOI21_X1 U4511 ( .B1(n3967), .B2(n3966), .A(n3965), .ZN(n3970) );
  XOR2_X1 U4512 ( .A(REG3_REG_0__SCAN_IN), .B(keyinput_180), .Z(n3969) );
  XNOR2_X1 U4513 ( .A(REG3_REG_9__SCAN_IN), .B(keyinput_179), .ZN(n3968) );
  NOR3_X1 U4514 ( .A1(n3970), .A2(n3969), .A3(n3968), .ZN(n3973) );
  XNOR2_X1 U4515 ( .A(REG3_REG_20__SCAN_IN), .B(keyinput_181), .ZN(n3972) );
  XNOR2_X1 U4516 ( .A(REG3_REG_13__SCAN_IN), .B(keyinput_182), .ZN(n3971) );
  NOR3_X1 U4517 ( .A1(n3973), .A2(n3972), .A3(n3971), .ZN(n3976) );
  XOR2_X1 U4518 ( .A(IR_REG_1__SCAN_IN), .B(keyinput_184), .Z(n3975) );
  XNOR2_X1 U4519 ( .A(IR_REG_0__SCAN_IN), .B(keyinput_183), .ZN(n3974) );
  NOR3_X1 U4520 ( .A1(n3976), .A2(n3975), .A3(n3974), .ZN(n3984) );
  XNOR2_X1 U4521 ( .A(IR_REG_2__SCAN_IN), .B(keyinput_185), .ZN(n3983) );
  XNOR2_X1 U4522 ( .A(n3977), .B(keyinput_186), .ZN(n3982) );
  OAI22_X1 U4523 ( .A1(n3980), .A2(keyinput_187), .B1(keyinput_188), .B2(
        IR_REG_5__SCAN_IN), .ZN(n3979) );
  AND2_X1 U4524 ( .A1(IR_REG_5__SCAN_IN), .A2(keyinput_188), .ZN(n3978) );
  AOI211_X1 U4525 ( .C1(keyinput_187), .C2(n3980), .A(n3979), .B(n3978), .ZN(
        n3981) );
  OAI211_X1 U4526 ( .C1(n3984), .C2(n3983), .A(n3982), .B(n3981), .ZN(n3992)
         );
  XNOR2_X1 U4527 ( .A(IR_REG_6__SCAN_IN), .B(keyinput_189), .ZN(n3987) );
  XNOR2_X1 U4528 ( .A(IR_REG_7__SCAN_IN), .B(keyinput_190), .ZN(n3986) );
  XNOR2_X1 U4529 ( .A(IR_REG_8__SCAN_IN), .B(keyinput_191), .ZN(n3985) );
  NOR3_X1 U4530 ( .A1(n3987), .A2(n3986), .A3(n3985), .ZN(n3991) );
  XNOR2_X1 U4531 ( .A(n3988), .B(keyinput_192), .ZN(n3990) );
  XOR2_X1 U4532 ( .A(IR_REG_10__SCAN_IN), .B(keyinput_193), .Z(n3989) );
  AOI211_X1 U4533 ( .C1(n3992), .C2(n3991), .A(n3990), .B(n3989), .ZN(n3995)
         );
  XNOR2_X1 U4534 ( .A(IR_REG_11__SCAN_IN), .B(keyinput_194), .ZN(n3994) );
  XNOR2_X1 U4535 ( .A(IR_REG_12__SCAN_IN), .B(keyinput_195), .ZN(n3993) );
  NOR3_X1 U4536 ( .A1(n3995), .A2(n3994), .A3(n3993), .ZN(n4001) );
  XNOR2_X1 U4537 ( .A(IR_REG_13__SCAN_IN), .B(keyinput_196), .ZN(n4000) );
  XNOR2_X1 U4538 ( .A(n3996), .B(keyinput_197), .ZN(n3999) );
  XNOR2_X1 U4539 ( .A(n3997), .B(keyinput_198), .ZN(n3998) );
  OAI211_X1 U4540 ( .C1(n4001), .C2(n4000), .A(n3999), .B(n3998), .ZN(n4004)
         );
  XOR2_X1 U4541 ( .A(IR_REG_16__SCAN_IN), .B(keyinput_199), .Z(n4003) );
  XNOR2_X1 U4542 ( .A(IR_REG_17__SCAN_IN), .B(keyinput_200), .ZN(n4002) );
  NAND3_X1 U4543 ( .A1(n4004), .A2(n4003), .A3(n4002), .ZN(n4010) );
  XNOR2_X1 U4544 ( .A(IR_REG_18__SCAN_IN), .B(keyinput_201), .ZN(n4009) );
  XNOR2_X1 U4545 ( .A(IR_REG_20__SCAN_IN), .B(keyinput_203), .ZN(n4007) );
  XNOR2_X1 U4546 ( .A(IR_REG_19__SCAN_IN), .B(keyinput_202), .ZN(n4006) );
  XNOR2_X1 U4547 ( .A(IR_REG_21__SCAN_IN), .B(keyinput_204), .ZN(n4005) );
  NAND3_X1 U4548 ( .A1(n4007), .A2(n4006), .A3(n4005), .ZN(n4008) );
  AOI21_X1 U4549 ( .B1(n4010), .B2(n4009), .A(n4008), .ZN(n4020) );
  XNOR2_X1 U4550 ( .A(n4011), .B(keyinput_207), .ZN(n4015) );
  XNOR2_X1 U4551 ( .A(IR_REG_23__SCAN_IN), .B(keyinput_206), .ZN(n4014) );
  XNOR2_X1 U4552 ( .A(IR_REG_22__SCAN_IN), .B(keyinput_205), .ZN(n4013) );
  XNOR2_X1 U4553 ( .A(IR_REG_25__SCAN_IN), .B(keyinput_208), .ZN(n4012) );
  NAND4_X1 U4554 ( .A1(n4015), .A2(n4014), .A3(n4013), .A4(n4012), .ZN(n4019)
         );
  XNOR2_X1 U4555 ( .A(n4016), .B(keyinput_210), .ZN(n4018) );
  XNOR2_X1 U4556 ( .A(IR_REG_26__SCAN_IN), .B(keyinput_209), .ZN(n4017) );
  OAI211_X1 U4557 ( .C1(n4020), .C2(n4019), .A(n4018), .B(n4017), .ZN(n4024)
         );
  XNOR2_X1 U4558 ( .A(n4021), .B(keyinput_211), .ZN(n4023) );
  XOR2_X1 U4559 ( .A(IR_REG_29__SCAN_IN), .B(keyinput_212), .Z(n4022) );
  AOI21_X1 U4560 ( .B1(n4024), .B2(n4023), .A(n4022), .ZN(n4027) );
  XNOR2_X1 U4561 ( .A(IR_REG_30__SCAN_IN), .B(keyinput_213), .ZN(n4026) );
  XNOR2_X1 U4562 ( .A(IR_REG_31__SCAN_IN), .B(keyinput_214), .ZN(n4025) );
  OAI21_X1 U4563 ( .B1(n4027), .B2(n4026), .A(n4025), .ZN(n4033) );
  XNOR2_X1 U4564 ( .A(D_REG_0__SCAN_IN), .B(keyinput_215), .ZN(n4032) );
  XOR2_X1 U4565 ( .A(D_REG_3__SCAN_IN), .B(keyinput_218), .Z(n4030) );
  XNOR2_X1 U4566 ( .A(D_REG_1__SCAN_IN), .B(keyinput_216), .ZN(n4029) );
  XNOR2_X1 U4567 ( .A(D_REG_2__SCAN_IN), .B(keyinput_217), .ZN(n4028) );
  NAND3_X1 U4568 ( .A1(n4030), .A2(n4029), .A3(n4028), .ZN(n4031) );
  AOI21_X1 U4569 ( .B1(n4033), .B2(n4032), .A(n4031), .ZN(n4036) );
  XNOR2_X1 U4570 ( .A(D_REG_4__SCAN_IN), .B(keyinput_219), .ZN(n4035) );
  XNOR2_X1 U4571 ( .A(D_REG_5__SCAN_IN), .B(keyinput_220), .ZN(n4034) );
  OAI21_X1 U4572 ( .B1(n4036), .B2(n4035), .A(n4034), .ZN(n4039) );
  XNOR2_X1 U4573 ( .A(D_REG_6__SCAN_IN), .B(keyinput_221), .ZN(n4038) );
  XNOR2_X1 U4574 ( .A(n5062), .B(keyinput_222), .ZN(n4037) );
  AOI21_X1 U4575 ( .B1(n4039), .B2(n4038), .A(n4037), .ZN(n4042) );
  XNOR2_X1 U4576 ( .A(n5064), .B(keyinput_224), .ZN(n4041) );
  XNOR2_X1 U4577 ( .A(D_REG_8__SCAN_IN), .B(keyinput_223), .ZN(n4040) );
  NOR3_X1 U4578 ( .A1(n4042), .A2(n4041), .A3(n4040), .ZN(n4045) );
  INV_X1 U4579 ( .A(D_REG_10__SCAN_IN), .ZN(n5065) );
  XNOR2_X1 U4580 ( .A(n5065), .B(keyinput_225), .ZN(n4044) );
  XNOR2_X1 U4581 ( .A(n5066), .B(keyinput_226), .ZN(n4043) );
  OAI21_X1 U4582 ( .B1(n4045), .B2(n4044), .A(n4043), .ZN(n4048) );
  XNOR2_X1 U4583 ( .A(D_REG_12__SCAN_IN), .B(keyinput_227), .ZN(n4047) );
  XNOR2_X1 U4584 ( .A(D_REG_13__SCAN_IN), .B(keyinput_228), .ZN(n4046) );
  NAND3_X1 U4585 ( .A1(n4048), .A2(n4047), .A3(n4046), .ZN(n4054) );
  XNOR2_X1 U4586 ( .A(n5069), .B(keyinput_229), .ZN(n4053) );
  XNOR2_X1 U4587 ( .A(D_REG_17__SCAN_IN), .B(keyinput_232), .ZN(n4051) );
  XNOR2_X1 U4588 ( .A(D_REG_16__SCAN_IN), .B(keyinput_231), .ZN(n4050) );
  XNOR2_X1 U4589 ( .A(D_REG_15__SCAN_IN), .B(keyinput_230), .ZN(n4049) );
  NAND3_X1 U4590 ( .A1(n4051), .A2(n4050), .A3(n4049), .ZN(n4052) );
  AOI21_X1 U4591 ( .B1(n4054), .B2(n4053), .A(n4052), .ZN(n4057) );
  INV_X1 U4592 ( .A(D_REG_18__SCAN_IN), .ZN(n5073) );
  XNOR2_X1 U4593 ( .A(n5073), .B(keyinput_233), .ZN(n4056) );
  XNOR2_X1 U4594 ( .A(D_REG_19__SCAN_IN), .B(keyinput_234), .ZN(n4055) );
  OAI21_X1 U4595 ( .B1(n4057), .B2(n4056), .A(n4055), .ZN(n4060) );
  XNOR2_X1 U4596 ( .A(D_REG_20__SCAN_IN), .B(keyinput_235), .ZN(n4059) );
  XNOR2_X1 U4597 ( .A(D_REG_21__SCAN_IN), .B(keyinput_236), .ZN(n4058) );
  AOI21_X1 U4598 ( .B1(n4060), .B2(n4059), .A(n4058), .ZN(n4063) );
  XNOR2_X1 U4599 ( .A(n5078), .B(keyinput_238), .ZN(n4062) );
  XNOR2_X1 U4600 ( .A(n5077), .B(keyinput_237), .ZN(n4061) );
  NOR3_X1 U4601 ( .A1(n4063), .A2(n4062), .A3(n4061), .ZN(n4071) );
  INV_X1 U4602 ( .A(keyinput_240), .ZN(n4064) );
  XNOR2_X1 U4603 ( .A(n4064), .B(D_REG_25__SCAN_IN), .ZN(n4068) );
  XNOR2_X1 U4604 ( .A(D_REG_27__SCAN_IN), .B(keyinput_242), .ZN(n4067) );
  XNOR2_X1 U4605 ( .A(D_REG_26__SCAN_IN), .B(keyinput_241), .ZN(n4066) );
  XNOR2_X1 U4606 ( .A(D_REG_24__SCAN_IN), .B(keyinput_239), .ZN(n4065) );
  NAND4_X1 U4607 ( .A1(n4068), .A2(n4067), .A3(n4066), .A4(n4065), .ZN(n4070)
         );
  XNOR2_X1 U4608 ( .A(D_REG_28__SCAN_IN), .B(keyinput_243), .ZN(n4069) );
  OAI21_X1 U4609 ( .B1(n4071), .B2(n4070), .A(n4069), .ZN(n4078) );
  INV_X1 U4610 ( .A(D_REG_29__SCAN_IN), .ZN(n5083) );
  XNOR2_X1 U4611 ( .A(n5083), .B(keyinput_244), .ZN(n4077) );
  INV_X1 U4612 ( .A(keyinput_247), .ZN(n4075) );
  XNOR2_X1 U4613 ( .A(D_REG_30__SCAN_IN), .B(keyinput_245), .ZN(n4074) );
  INV_X1 U4614 ( .A(REG0_REG_0__SCAN_IN), .ZN(n5112) );
  OAI22_X1 U4615 ( .A1(n5112), .A2(keyinput_247), .B1(D_REG_31__SCAN_IN), .B2(
        keyinput_246), .ZN(n4072) );
  AOI21_X1 U4616 ( .B1(D_REG_31__SCAN_IN), .B2(keyinput_246), .A(n4072), .ZN(
        n4073) );
  OAI211_X1 U4617 ( .C1(REG0_REG_0__SCAN_IN), .C2(n4075), .A(n4074), .B(n4073), 
        .ZN(n4076) );
  AOI21_X1 U4618 ( .B1(n4078), .B2(n4077), .A(n4076), .ZN(n4081) );
  XOR2_X1 U4619 ( .A(REG0_REG_1__SCAN_IN), .B(keyinput_248), .Z(n4080) );
  XNOR2_X1 U4620 ( .A(REG0_REG_2__SCAN_IN), .B(keyinput_249), .ZN(n4079) );
  OAI21_X1 U4621 ( .B1(n4081), .B2(n4080), .A(n4079), .ZN(n4084) );
  XOR2_X1 U4622 ( .A(REG0_REG_3__SCAN_IN), .B(keyinput_250), .Z(n4083) );
  XNOR2_X1 U4623 ( .A(REG0_REG_4__SCAN_IN), .B(keyinput_251), .ZN(n4082) );
  NAND3_X1 U4624 ( .A1(n4084), .A2(n4083), .A3(n4082), .ZN(n4088) );
  XOR2_X1 U4625 ( .A(REG0_REG_6__SCAN_IN), .B(keyinput_253), .Z(n4087) );
  XOR2_X1 U4626 ( .A(REG0_REG_7__SCAN_IN), .B(keyinput_254), .Z(n4086) );
  XNOR2_X1 U4627 ( .A(REG0_REG_5__SCAN_IN), .B(keyinput_252), .ZN(n4085) );
  NAND4_X1 U4628 ( .A1(n4088), .A2(n4087), .A3(n4086), .A4(n4085), .ZN(n4089)
         );
  OAI211_X1 U4629 ( .C1(n4092), .C2(n4091), .A(n4090), .B(n4089), .ZN(n4095)
         );
  MUX2_X1 U4630 ( .A(n4093), .B(DATAI_27_), .S(U3149), .Z(n4094) );
  XNOR2_X1 U4631 ( .A(n4095), .B(n4094), .ZN(U3325) );
  NAND2_X1 U4632 ( .A1(n4139), .A2(n4120), .ZN(n4461) );
  NAND2_X1 U4633 ( .A1(n4583), .A2(n4097), .ZN(n4134) );
  XNOR2_X1 U4634 ( .A(n4126), .B(n4536), .ZN(n4100) );
  OAI22_X1 U4635 ( .A1(n4102), .A2(n5186), .B1(n4128), .B2(n5188), .ZN(n4098)
         );
  AOI21_X1 U4636 ( .B1(n4120), .B2(n5191), .A(n4098), .ZN(n4099) );
  OAI21_X1 U4637 ( .B1(n4100), .B2(n5194), .A(n4099), .ZN(n5248) );
  INV_X1 U4638 ( .A(n5248), .ZN(n4110) );
  XNOR2_X1 U4639 ( .A(n4121), .B(n4536), .ZN(n5250) );
  NAND2_X1 U4640 ( .A1(n5250), .A2(n4935), .ZN(n4109) );
  NAND2_X1 U4641 ( .A1(n4103), .A2(n4120), .ZN(n4104) );
  NAND2_X1 U4642 ( .A1(n4104), .A2(n5333), .ZN(n4105) );
  NOR2_X1 U4643 ( .A1(n4149), .A2(n4105), .ZN(n5249) );
  INV_X1 U4644 ( .A(REG2_REG_12__SCAN_IN), .ZN(n4173) );
  INV_X1 U4645 ( .A(n4116), .ZN(n4106) );
  OAI22_X1 U4646 ( .A1(n5208), .A2(n4173), .B1(n4106), .B2(n5210), .ZN(n4107)
         );
  AOI21_X1 U4647 ( .B1(n5249), .B2(n4943), .A(n4107), .ZN(n4108) );
  OAI211_X1 U4648 ( .C1(n5330), .C2(n4110), .A(n4109), .B(n4108), .ZN(U3278)
         );
  NAND2_X1 U4649 ( .A1(n4111), .A2(n4157), .ZN(n4113) );
  XOR2_X1 U4650 ( .A(n4113), .B(n4112), .Z(n4119) );
  AOI22_X1 U4651 ( .A1(n4410), .A2(n4584), .B1(n4120), .B2(n5276), .ZN(n4118)
         );
  NOR2_X1 U4652 ( .A1(STATE_REG_SCAN_IN), .A2(n4114), .ZN(n4177) );
  NOR2_X1 U4653 ( .A1(n5271), .A2(n4128), .ZN(n4115) );
  AOI211_X1 U4654 ( .C1(n4345), .C2(n4116), .A(n4177), .B(n4115), .ZN(n4117)
         );
  OAI211_X1 U4655 ( .C1(n4119), .C2(n4417), .A(n4118), .B(n4117), .ZN(U3221)
         );
  INV_X1 U4656 ( .A(n4128), .ZN(n4582) );
  INV_X1 U4657 ( .A(n4148), .ZN(n4163) );
  AND2_X1 U4658 ( .A1(n4582), .A2(n4163), .ZN(n4143) );
  NAND2_X1 U4659 ( .A1(n5273), .A2(n4198), .ZN(n4507) );
  NAND2_X1 U4660 ( .A1(n4581), .A2(n4199), .ZN(n4442) );
  NAND2_X1 U4661 ( .A1(n4507), .A2(n4442), .ZN(n4191) );
  NAND2_X1 U4662 ( .A1(n4122), .A2(n4191), .ZN(n4201) );
  OAI21_X1 U4663 ( .B1(n4122), .B2(n4191), .A(n4201), .ZN(n4123) );
  INV_X1 U4664 ( .A(n4123), .ZN(n5265) );
  INV_X1 U4665 ( .A(n4203), .ZN(n4124) );
  AOI21_X1 U4666 ( .B1(n4198), .B2(n4150), .A(n4124), .ZN(n5262) );
  INV_X1 U4667 ( .A(REG2_REG_14__SCAN_IN), .ZN(n4623) );
  OAI22_X1 U4668 ( .A1(n5208), .A2(n4623), .B1(n4186), .B2(n5210), .ZN(n4125)
         );
  AOI21_X1 U4669 ( .B1(n5262), .B2(n5328), .A(n4125), .ZN(n4133) );
  NAND2_X1 U4670 ( .A1(n4582), .A2(n4148), .ZN(n4136) );
  AND2_X1 U4671 ( .A1(n4134), .A2(n4136), .ZN(n4458) );
  NAND2_X1 U4672 ( .A1(n4135), .A2(n4458), .ZN(n4127) );
  NAND2_X1 U4673 ( .A1(n4128), .A2(n4163), .ZN(n4457) );
  NAND2_X1 U4674 ( .A1(n4127), .A2(n4457), .ZN(n4192) );
  XNOR2_X1 U4675 ( .A(n4192), .B(n4191), .ZN(n4131) );
  OAI22_X1 U4676 ( .A1(n4128), .A2(n5186), .B1(n4223), .B2(n5188), .ZN(n4129)
         );
  AOI21_X1 U4677 ( .B1(n4198), .B2(n5191), .A(n4129), .ZN(n4130) );
  OAI21_X1 U4678 ( .B1(n4131), .B2(n5194), .A(n4130), .ZN(n5267) );
  NAND2_X1 U4679 ( .A1(n5267), .A2(n5208), .ZN(n4132) );
  OAI211_X1 U4680 ( .C1(n5265), .C2(n4962), .A(n4133), .B(n4132), .ZN(U3276)
         );
  NAND2_X1 U4681 ( .A1(n4135), .A2(n4134), .ZN(n4137) );
  NAND2_X1 U4682 ( .A1(n4457), .A2(n4136), .ZN(n4555) );
  XNOR2_X1 U4683 ( .A(n4137), .B(n4555), .ZN(n4138) );
  NAND2_X1 U4684 ( .A1(n4138), .A2(n5108), .ZN(n4142) );
  OAI22_X1 U4685 ( .A1(n5273), .A2(n5188), .B1(n4139), .B2(n5186), .ZN(n4140)
         );
  INV_X1 U4686 ( .A(n4140), .ZN(n4141) );
  OAI211_X1 U4687 ( .C1(n5319), .C2(n4148), .A(n4142), .B(n4141), .ZN(n5256)
         );
  INV_X1 U4688 ( .A(n5256), .ZN(n4156) );
  INV_X1 U4689 ( .A(n4143), .ZN(n4146) );
  INV_X1 U4690 ( .A(n4555), .ZN(n4145) );
  AOI22_X1 U4691 ( .A1(n4147), .A2(n4146), .B1(n4145), .B2(n4144), .ZN(n5258)
         );
  NOR2_X1 U4692 ( .A1(n4149), .A2(n4148), .ZN(n5255) );
  INV_X1 U4693 ( .A(n4150), .ZN(n5254) );
  NOR3_X1 U4694 ( .A1(n5255), .A2(n5254), .A3(n4904), .ZN(n4154) );
  INV_X1 U4695 ( .A(REG2_REG_13__SCAN_IN), .ZN(n4152) );
  INV_X1 U4696 ( .A(n4151), .ZN(n4166) );
  OAI22_X1 U4697 ( .A1(n5208), .A2(n4152), .B1(n4166), .B2(n5210), .ZN(n4153)
         );
  AOI211_X1 U4698 ( .C1(n5258), .C2(n4935), .A(n4154), .B(n4153), .ZN(n4155)
         );
  OAI21_X1 U4699 ( .B1(n5330), .B2(n4156), .A(n4155), .ZN(U3277) );
  NAND2_X1 U4700 ( .A1(n4158), .A2(n4157), .ZN(n4161) );
  INV_X1 U4701 ( .A(n4159), .ZN(n4160) );
  AOI21_X1 U4702 ( .B1(n4162), .B2(n4161), .A(n4160), .ZN(n4170) );
  AOI22_X1 U4703 ( .A1(n4399), .A2(n4583), .B1(n4163), .B2(n5276), .ZN(n4169)
         );
  NOR2_X1 U4704 ( .A1(n4164), .A2(STATE_REG_SCAN_IN), .ZN(n4610) );
  INV_X1 U4705 ( .A(n4610), .ZN(n4165) );
  OAI21_X1 U4706 ( .B1(n5287), .B2(n4166), .A(n4165), .ZN(n4167) );
  AOI21_X1 U4707 ( .B1(n4414), .B2(n4581), .A(n4167), .ZN(n4168) );
  OAI211_X1 U4708 ( .C1(n4170), .C2(n4417), .A(n4169), .B(n4168), .ZN(U3231)
         );
  INV_X1 U4709 ( .A(n5048), .ZN(n4601) );
  AOI211_X1 U4710 ( .C1(n4173), .C2(n4172), .A(n4603), .B(n5090), .ZN(n4181)
         );
  NAND2_X1 U4711 ( .A1(n5049), .A2(REG1_REG_11__SCAN_IN), .ZN(n4175) );
  NAND2_X1 U4712 ( .A1(REG1_REG_12__SCAN_IN), .A2(n4176), .ZN(n4595) );
  OAI211_X1 U4713 ( .C1(n4176), .C2(REG1_REG_12__SCAN_IN), .A(n5099), .B(n4595), .ZN(n4179) );
  AOI21_X1 U4714 ( .B1(n5088), .B2(ADDR_REG_12__SCAN_IN), .A(n4177), .ZN(n4178) );
  OAI211_X1 U4715 ( .C1(n5089), .C2(n4601), .A(n4179), .B(n4178), .ZN(n4180)
         );
  OR2_X1 U4716 ( .A1(n4181), .A2(n4180), .ZN(U3252) );
  XOR2_X1 U4717 ( .A(n4183), .B(n4182), .Z(n4190) );
  AOI22_X1 U4718 ( .A1(n4399), .A2(n4582), .B1(n4198), .B2(n5276), .ZN(n4189)
         );
  NOR2_X1 U4719 ( .A1(n4184), .A2(STATE_REG_SCAN_IN), .ZN(n4617) );
  INV_X1 U4720 ( .A(n4617), .ZN(n4185) );
  OAI21_X1 U4721 ( .B1(n5287), .B2(n4186), .A(n4185), .ZN(n4187) );
  AOI21_X1 U4722 ( .B1(n4414), .B2(n4950), .A(n4187), .ZN(n4188) );
  OAI211_X1 U4723 ( .C1(n4190), .C2(n4417), .A(n4189), .B(n4188), .ZN(U3212)
         );
  INV_X1 U4724 ( .A(n4191), .ZN(n4553) );
  NAND2_X1 U4725 ( .A1(n4192), .A2(n4553), .ZN(n4193) );
  INV_X1 U4726 ( .A(n4194), .ZN(n4195) );
  NAND2_X1 U4727 ( .A1(n4223), .A2(n5277), .ZN(n4509) );
  NAND2_X1 U4728 ( .A1(n4950), .A2(n4222), .ZN(n4443) );
  NAND2_X1 U4729 ( .A1(n4509), .A2(n4443), .ZN(n4202) );
  INV_X1 U4730 ( .A(n4202), .ZN(n4540) );
  OAI211_X1 U4731 ( .C1(n4195), .C2(n4540), .A(n5108), .B(n4234), .ZN(n4197)
         );
  AOI22_X1 U4732 ( .A1(n4581), .A2(n5157), .B1(n5154), .B2(n4929), .ZN(n4196)
         );
  OAI211_X1 U4733 ( .C1(n5319), .C2(n4222), .A(n4197), .B(n4196), .ZN(n5288)
         );
  INV_X1 U4734 ( .A(n5288), .ZN(n4209) );
  NAND2_X1 U4735 ( .A1(n4201), .A2(n4200), .ZN(n4224) );
  XNOR2_X1 U4736 ( .A(n4224), .B(n4202), .ZN(n5290) );
  NAND2_X1 U4737 ( .A1(n5290), .A2(n4935), .ZN(n4208) );
  NAND2_X1 U4738 ( .A1(n4203), .A2(n5277), .ZN(n4204) );
  NAND2_X1 U4739 ( .A1(n4204), .A2(n5333), .ZN(n4205) );
  NOR2_X1 U4740 ( .A1(n4954), .A2(n4205), .ZN(n5289) );
  INV_X1 U4741 ( .A(REG2_REG_15__SCAN_IN), .ZN(n4630) );
  OAI22_X1 U4742 ( .A1(n5208), .A2(n4630), .B1(n5286), .B2(n5210), .ZN(n4206)
         );
  AOI21_X1 U4743 ( .B1(n5289), .B2(n4943), .A(n4206), .ZN(n4207) );
  OAI211_X1 U4744 ( .C1(n5330), .C2(n4209), .A(n4208), .B(n4207), .ZN(U3275)
         );
  XNOR2_X1 U4745 ( .A(n4210), .B(n4538), .ZN(n5141) );
  XNOR2_X1 U4746 ( .A(n4211), .B(n4538), .ZN(n4215) );
  AOI22_X1 U4747 ( .A1(n5157), .A2(n4591), .B1(n4590), .B2(n5154), .ZN(n4212)
         );
  OAI21_X1 U4748 ( .B1(n4213), .B2(n5319), .A(n4212), .ZN(n4214) );
  AOI21_X1 U4749 ( .B1(n4215), .B2(n5108), .A(n4214), .ZN(n4216) );
  OAI21_X1 U4750 ( .B1(n5141), .B2(n4968), .A(n4216), .ZN(n5142) );
  NAND2_X1 U4751 ( .A1(n5142), .A2(n5208), .ZN(n4221) );
  AOI21_X1 U4752 ( .B1(n4218), .B2(n4217), .A(n5151), .ZN(n5144) );
  OAI22_X1 U4753 ( .A1(n5208), .A2(n3391), .B1(REG3_REG_3__SCAN_IN), .B2(n5210), .ZN(n4219) );
  AOI21_X1 U4754 ( .B1(n5144), .B2(n5328), .A(n4219), .ZN(n4220) );
  OAI211_X1 U4755 ( .C1(n5141), .C2(n4795), .A(n4221), .B(n4220), .ZN(U3287)
         );
  INV_X1 U4756 ( .A(n4953), .ZN(n4957) );
  NAND2_X1 U4757 ( .A1(n4224), .A2(n2536), .ZN(n4226) );
  AND2_X1 U4758 ( .A1(n4929), .A2(n4953), .ZN(n4470) );
  INV_X1 U4759 ( .A(n4929), .ZN(n5270) );
  NAND2_X1 U4760 ( .A1(n5270), .A2(n4957), .ZN(n4506) );
  AND2_X1 U4761 ( .A1(n4949), .A2(n4936), .ZN(n4471) );
  INV_X1 U4762 ( .A(n4936), .ZN(n4341) );
  NAND2_X1 U4763 ( .A1(n4227), .A2(n4341), .ZN(n4910) );
  NAND2_X1 U4764 ( .A1(n4236), .A2(n4910), .ZN(n4933) );
  NAND2_X1 U4765 ( .A1(n4932), .A2(n4228), .ZN(n4907) );
  INV_X1 U4766 ( .A(n4928), .ZN(n4343) );
  NAND2_X1 U4767 ( .A1(n4343), .A2(n4916), .ZN(n4238) );
  NAND2_X1 U4768 ( .A1(n4928), .A2(n4918), .ZN(n4890) );
  NAND2_X1 U4769 ( .A1(n4238), .A2(n4890), .ZN(n4889) );
  XNOR2_X1 U4770 ( .A(n4580), .B(n4898), .ZN(n4900) );
  NAND2_X1 U4771 ( .A1(n4892), .A2(n4376), .ZN(n4846) );
  INV_X1 U4772 ( .A(n4840), .ZN(n4877) );
  NOR2_X1 U4773 ( .A1(n4877), .A2(n4867), .ZN(n4847) );
  AND2_X1 U4774 ( .A1(n4579), .A2(n4385), .ZN(n4231) );
  AND2_X1 U4775 ( .A1(n4846), .A2(n2767), .ZN(n4233) );
  NAND2_X1 U4776 ( .A1(n4877), .A2(n4867), .ZN(n4848) );
  NAND2_X1 U4777 ( .A1(n4861), .A2(n4385), .ZN(n4478) );
  NAND2_X1 U4778 ( .A1(n4579), .A2(n4852), .ZN(n4480) );
  INV_X1 U4779 ( .A(n4850), .ZN(n4526) );
  AND2_X1 U4780 ( .A1(n4848), .A2(n4526), .ZN(n4230) );
  NOR2_X1 U4781 ( .A1(n4231), .A2(n4230), .ZN(n4232) );
  XNOR2_X1 U4782 ( .A(n4839), .B(n4716), .ZN(n4558) );
  XNOR2_X1 U4783 ( .A(n4719), .B(n4558), .ZN(n4998) );
  NAND2_X1 U4784 ( .A1(n4580), .A2(n4898), .ZN(n4237) );
  NAND2_X1 U4785 ( .A1(n4890), .A2(n4237), .ZN(n4469) );
  INV_X1 U4786 ( .A(n4580), .ZN(n4908) );
  AOI21_X1 U4787 ( .B1(n4238), .B2(n4910), .A(n4469), .ZN(n4239) );
  AOI21_X1 U4788 ( .B1(n4294), .B2(n4908), .A(n4239), .ZN(n4476) );
  NOR2_X1 U4789 ( .A1(n4862), .A2(n4376), .ZN(n4545) );
  INV_X1 U4790 ( .A(n4545), .ZN(n4240) );
  NAND2_X1 U4791 ( .A1(n4862), .A2(n4376), .ZN(n4475) );
  INV_X1 U4792 ( .A(n4475), .ZN(n4544) );
  INV_X1 U4793 ( .A(n4867), .ZN(n4314) );
  NAND2_X1 U4794 ( .A1(n4877), .A2(n4314), .ZN(n4474) );
  AND2_X1 U4795 ( .A1(n4840), .A2(n4867), .ZN(n4477) );
  AOI21_X1 U4796 ( .B1(n4860), .B2(n4474), .A(n4477), .ZN(n4838) );
  NAND2_X1 U4797 ( .A1(n4838), .A2(n4850), .ZN(n4837) );
  NAND2_X1 U4798 ( .A1(n4837), .A2(n4478), .ZN(n4242) );
  INV_X1 U4799 ( .A(n4558), .ZN(n4241) );
  XNOR2_X1 U4800 ( .A(n4242), .B(n4241), .ZN(n4245) );
  INV_X1 U4801 ( .A(n4720), .ZN(n4800) );
  NOR2_X1 U4802 ( .A1(n4800), .A2(n5188), .ZN(n4244) );
  OAI22_X1 U4803 ( .A1(n4861), .A2(n5186), .B1(n4716), .B2(n5319), .ZN(n4243)
         );
  AOI211_X1 U4804 ( .C1(n4245), .C2(n5108), .A(n4244), .B(n4243), .ZN(n4997)
         );
  INV_X1 U4805 ( .A(n4997), .ZN(n4249) );
  AOI21_X1 U4806 ( .B1(n2500), .B2(n4273), .A(n5264), .ZN(n4246) );
  NAND2_X1 U4807 ( .A1(n4246), .A2(n4828), .ZN(n4996) );
  AOI22_X1 U4808 ( .A1(n5330), .A2(REG2_REG_23__SCAN_IN), .B1(n4274), .B2(
        n5118), .ZN(n4247) );
  OAI21_X1 U4809 ( .B1(n4996), .B2(n4922), .A(n4247), .ZN(n4248) );
  AOI21_X1 U4810 ( .B1(n4249), .B2(n5208), .A(n4248), .ZN(n4250) );
  OAI21_X1 U4811 ( .B1(n4998), .B2(n4962), .A(n4250), .ZN(U3267) );
  AOI21_X1 U4812 ( .B1(n4252), .B2(n4251), .A(n4417), .ZN(n4254) );
  NAND2_X1 U4813 ( .A1(n4254), .A2(n4253), .ZN(n4261) );
  AOI22_X1 U4814 ( .A1(n4410), .A2(n4589), .B1(n4255), .B2(n5276), .ZN(n4260)
         );
  NOR2_X1 U4815 ( .A1(n5287), .A2(n4256), .ZN(n4257) );
  AOI211_X1 U4816 ( .C1(n4414), .C2(n4587), .A(n4258), .B(n4257), .ZN(n4259)
         );
  NAND3_X1 U4817 ( .A1(n4261), .A2(n4260), .A3(n4259), .ZN(U3210) );
  OAI211_X1 U4818 ( .C1(n4264), .C2(n4263), .A(n4262), .B(n5282), .ZN(n4268)
         );
  INV_X1 U4819 ( .A(n4770), .ZN(n4496) );
  AOI22_X1 U4820 ( .A1(n4410), .A2(n4809), .B1(n4496), .B2(n5276), .ZN(n4267)
         );
  AOI22_X1 U4821 ( .A1(n4345), .A2(n4772), .B1(REG3_REG_27__SCAN_IN), .B2(
        U3149), .ZN(n4266) );
  NAND2_X1 U4822 ( .A1(n4414), .A2(n4768), .ZN(n4265) );
  NAND4_X1 U4823 ( .A1(n4268), .A2(n4267), .A3(n4266), .A4(n4265), .ZN(U3211)
         );
  AOI21_X1 U4824 ( .B1(n4269), .B2(n4270), .A(n4417), .ZN(n4272) );
  NAND2_X1 U4825 ( .A1(n4272), .A2(n4271), .ZN(n4278) );
  AOI22_X1 U4826 ( .A1(n4410), .A2(n4579), .B1(n4273), .B2(n5276), .ZN(n4277)
         );
  AOI22_X1 U4827 ( .A1(n4345), .A2(n4274), .B1(REG3_REG_23__SCAN_IN), .B2(
        U3149), .ZN(n4276) );
  NAND2_X1 U4828 ( .A1(n4414), .A2(n4720), .ZN(n4275) );
  NAND4_X1 U4829 ( .A1(n4278), .A2(n4277), .A3(n4276), .A4(n4275), .ZN(U3213)
         );
  OAI211_X1 U4830 ( .C1(n4281), .C2(n4280), .A(n4279), .B(n5282), .ZN(n4289)
         );
  AOI22_X1 U4831 ( .A1(n4410), .A2(n4586), .B1(n4282), .B2(n5276), .ZN(n4288)
         );
  INV_X1 U4832 ( .A(n4283), .ZN(n4284) );
  OAI21_X1 U4833 ( .B1(n5287), .B2(n4285), .A(n4284), .ZN(n4286) );
  AOI21_X1 U4834 ( .B1(n4414), .B2(n4584), .A(n4286), .ZN(n4287) );
  NAND3_X1 U4835 ( .A1(n4289), .A2(n4288), .A3(n4287), .ZN(U3214) );
  OAI21_X1 U4836 ( .B1(n4292), .B2(n4291), .A(n4290), .ZN(n4293) );
  NAND2_X1 U4837 ( .A1(n4293), .A2(n5282), .ZN(n4299) );
  AOI22_X1 U4838 ( .A1(n4410), .A2(n4928), .B1(n4294), .B2(n5276), .ZN(n4298)
         );
  INV_X1 U4839 ( .A(REG3_REG_19__SCAN_IN), .ZN(n4295) );
  NOR2_X1 U4840 ( .A1(STATE_REG_SCAN_IN), .A2(n4295), .ZN(n4693) );
  AOI21_X1 U4841 ( .B1(n4345), .B2(n4901), .A(n4693), .ZN(n4297) );
  NAND2_X1 U4842 ( .A1(n4414), .A2(n4892), .ZN(n4296) );
  NAND4_X1 U4843 ( .A1(n4299), .A2(n4298), .A3(n4297), .A4(n4296), .ZN(U3216)
         );
  OAI211_X1 U4844 ( .C1(n4302), .C2(n4301), .A(n4300), .B(n5282), .ZN(n4307)
         );
  AOI22_X1 U4845 ( .A1(n5276), .A2(n4304), .B1(REG3_REG_1__SCAN_IN), .B2(n4303), .ZN(n4306) );
  AOI22_X1 U4846 ( .A1(n4410), .A2(n4593), .B1(n4414), .B2(n4591), .ZN(n4305)
         );
  NAND3_X1 U4847 ( .A1(n4307), .A2(n4306), .A3(n4305), .ZN(U3219) );
  OAI21_X1 U4848 ( .B1(n2750), .B2(n4310), .A(n4309), .ZN(n4312) );
  INV_X1 U4849 ( .A(n4309), .ZN(n4311) );
  AOI22_X1 U4850 ( .A1(n4313), .A2(n4312), .B1(n4311), .B2(n2750), .ZN(n4320)
         );
  AOI22_X1 U4851 ( .A1(n4410), .A2(n4892), .B1(n4314), .B2(n5276), .ZN(n4319)
         );
  INV_X1 U4852 ( .A(n4868), .ZN(n4316) );
  INV_X1 U4853 ( .A(REG3_REG_21__SCAN_IN), .ZN(n4315) );
  OAI22_X1 U4854 ( .A1(n5287), .A2(n4316), .B1(STATE_REG_SCAN_IN), .B2(n4315), 
        .ZN(n4317) );
  AOI21_X1 U4855 ( .B1(n4414), .B2(n4579), .A(n4317), .ZN(n4318) );
  OAI211_X1 U4856 ( .C1(n4320), .C2(n4417), .A(n4319), .B(n4318), .ZN(U3220)
         );
  AOI22_X1 U4857 ( .A1(n4410), .A2(n4720), .B1(n4724), .B2(n5276), .ZN(n4327)
         );
  INV_X1 U4858 ( .A(n4813), .ZN(n4324) );
  INV_X1 U4859 ( .A(REG3_REG_25__SCAN_IN), .ZN(n4323) );
  OAI22_X1 U4860 ( .A1(n5287), .A2(n4324), .B1(STATE_REG_SCAN_IN), .B2(n4323), 
        .ZN(n4325) );
  AOI21_X1 U4861 ( .B1(n4414), .B2(n4809), .A(n4325), .ZN(n4326) );
  OAI211_X1 U4862 ( .C1(n4328), .C2(n4417), .A(n4327), .B(n4326), .ZN(U3222)
         );
  XOR2_X1 U4863 ( .A(n4331), .B(n4330), .Z(n4332) );
  XNOR2_X1 U4864 ( .A(n4329), .B(n4332), .ZN(n4337) );
  AOI22_X1 U4865 ( .A1(n4399), .A2(n4950), .B1(n4957), .B2(n5276), .ZN(n4336)
         );
  NOR2_X1 U4866 ( .A1(STATE_REG_SCAN_IN), .A2(n4333), .ZN(n4652) );
  NOR2_X1 U4867 ( .A1(n5287), .A2(n4958), .ZN(n4334) );
  AOI211_X1 U4868 ( .C1(n4414), .C2(n4949), .A(n4652), .B(n4334), .ZN(n4335)
         );
  OAI211_X1 U4869 ( .C1(n4337), .C2(n4417), .A(n4336), .B(n4335), .ZN(U3223)
         );
  OR2_X1 U4870 ( .A1(n4338), .A2(n4340), .ZN(n4397) );
  INV_X1 U4871 ( .A(n4397), .ZN(n4339) );
  AOI21_X1 U4872 ( .B1(n4340), .B2(n4338), .A(n4339), .ZN(n4348) );
  AOI22_X1 U4873 ( .A1(n4399), .A2(n4929), .B1(n4341), .B2(n5276), .ZN(n4347)
         );
  NOR2_X1 U4874 ( .A1(STATE_REG_SCAN_IN), .A2(n4342), .ZN(n4668) );
  NOR2_X1 U4875 ( .A1(n5271), .A2(n4343), .ZN(n4344) );
  AOI211_X1 U4876 ( .C1(n4345), .C2(n4939), .A(n4668), .B(n4344), .ZN(n4346)
         );
  OAI211_X1 U4877 ( .C1(n4348), .C2(n4417), .A(n4347), .B(n4346), .ZN(U3225)
         );
  NAND2_X1 U4878 ( .A1(n2585), .A2(n4350), .ZN(n4352) );
  XNOR2_X1 U4879 ( .A(n4352), .B(n4351), .ZN(n4358) );
  AOI22_X1 U4880 ( .A1(n4414), .A2(n4725), .B1(n4827), .B2(n5276), .ZN(n4357)
         );
  INV_X1 U4881 ( .A(n4832), .ZN(n4354) );
  INV_X1 U4882 ( .A(REG3_REG_24__SCAN_IN), .ZN(n4353) );
  OAI22_X1 U4883 ( .A1(n5287), .A2(n4354), .B1(STATE_REG_SCAN_IN), .B2(n4353), 
        .ZN(n4355) );
  AOI21_X1 U4884 ( .B1(n4410), .B2(n4839), .A(n4355), .ZN(n4356) );
  OAI211_X1 U4885 ( .C1(n4358), .C2(n4417), .A(n4357), .B(n4356), .ZN(U3226)
         );
  INV_X1 U4886 ( .A(n4359), .ZN(n4360) );
  NAND2_X1 U4887 ( .A1(n4361), .A2(n4360), .ZN(n4362) );
  AND2_X1 U4888 ( .A1(n4363), .A2(n4362), .ZN(n4365) );
  AOI21_X1 U4889 ( .B1(n4365), .B2(n4364), .A(n4417), .ZN(n4366) );
  NAND2_X1 U4890 ( .A1(n4366), .A2(n2542), .ZN(n4371) );
  AOI22_X1 U4891 ( .A1(n4410), .A2(n5156), .B1(n5158), .B2(n5276), .ZN(n4370)
         );
  NOR2_X1 U4892 ( .A1(STATE_REG_SCAN_IN), .A2(n4367), .ZN(n5087) );
  NOR2_X1 U4893 ( .A1(n5287), .A2(n5177), .ZN(n4368) );
  AOI211_X1 U4894 ( .C1(n4414), .C2(n5155), .A(n5087), .B(n4368), .ZN(n4369)
         );
  NAND3_X1 U4895 ( .A1(n4371), .A2(n4370), .A3(n4369), .ZN(U3227) );
  NAND2_X1 U4896 ( .A1(n4373), .A2(n4372), .ZN(n4374) );
  XNOR2_X1 U4897 ( .A(n4375), .B(n4374), .ZN(n4382) );
  AOI22_X1 U4898 ( .A1(n4399), .A2(n4580), .B1(n4376), .B2(n5276), .ZN(n4381)
         );
  INV_X1 U4899 ( .A(n4884), .ZN(n4378) );
  INV_X1 U4900 ( .A(REG3_REG_20__SCAN_IN), .ZN(n4377) );
  OAI22_X1 U4901 ( .A1(n5287), .A2(n4378), .B1(STATE_REG_SCAN_IN), .B2(n4377), 
        .ZN(n4379) );
  AOI21_X1 U4902 ( .B1(n4414), .B2(n4840), .A(n4379), .ZN(n4380) );
  OAI211_X1 U4903 ( .C1(n4382), .C2(n4417), .A(n4381), .B(n4380), .ZN(U3230)
         );
  AOI21_X1 U4904 ( .B1(n4384), .B2(n4383), .A(n2768), .ZN(n4391) );
  AOI22_X1 U4905 ( .A1(n4410), .A2(n4840), .B1(n4385), .B2(n5276), .ZN(n4390)
         );
  INV_X1 U4906 ( .A(n4853), .ZN(n4387) );
  INV_X1 U4907 ( .A(REG3_REG_22__SCAN_IN), .ZN(n4386) );
  OAI22_X1 U4908 ( .A1(n5287), .A2(n4387), .B1(STATE_REG_SCAN_IN), .B2(n4386), 
        .ZN(n4388) );
  AOI21_X1 U4909 ( .B1(n4414), .B2(n4839), .A(n4388), .ZN(n4389) );
  OAI211_X1 U4910 ( .C1(n4391), .C2(n4417), .A(n4390), .B(n4389), .ZN(U3232)
         );
  INV_X1 U4911 ( .A(n4392), .ZN(n4393) );
  NOR2_X1 U4912 ( .A1(n4394), .A2(n4393), .ZN(n4398) );
  AOI21_X1 U4913 ( .B1(n4398), .B2(n4397), .A(n2529), .ZN(n4405) );
  AOI22_X1 U4914 ( .A1(n4399), .A2(n4949), .B1(n4916), .B2(n5276), .ZN(n4404)
         );
  INV_X1 U4915 ( .A(REG3_REG_18__SCAN_IN), .ZN(n4400) );
  NOR2_X1 U4916 ( .A1(n4400), .A2(STATE_REG_SCAN_IN), .ZN(n4677) );
  NOR2_X1 U4917 ( .A1(n5287), .A2(n4401), .ZN(n4402) );
  AOI211_X1 U4918 ( .C1(n4414), .C2(n4580), .A(n4677), .B(n4402), .ZN(n4403)
         );
  OAI211_X1 U4919 ( .C1(n4405), .C2(n4417), .A(n4404), .B(n4403), .ZN(U3235)
         );
  NAND2_X1 U4920 ( .A1(n2738), .A2(n4407), .ZN(n4408) );
  XNOR2_X1 U4921 ( .A(n4409), .B(n4408), .ZN(n4418) );
  INV_X1 U4922 ( .A(n4785), .ZN(n4791) );
  AOI22_X1 U4923 ( .A1(n4410), .A2(n4725), .B1(n4791), .B2(n5276), .ZN(n4416)
         );
  INV_X1 U4924 ( .A(n4411), .ZN(n4792) );
  INV_X1 U4925 ( .A(REG3_REG_26__SCAN_IN), .ZN(n4412) );
  OAI22_X1 U4926 ( .A1(n5287), .A2(n4792), .B1(STATE_REG_SCAN_IN), .B2(n4412), 
        .ZN(n4413) );
  AOI21_X1 U4927 ( .B1(n4414), .B2(n4787), .A(n4413), .ZN(n4415) );
  OAI211_X1 U4928 ( .C1(n4418), .C2(n4417), .A(n4416), .B(n4415), .ZN(U3237)
         );
  NOR2_X1 U4929 ( .A1(n4720), .A2(n4822), .ZN(n4700) );
  NOR2_X1 U4930 ( .A1(n4839), .A2(n4716), .ZN(n4698) );
  NOR2_X1 U4931 ( .A1(n4700), .A2(n4698), .ZN(n4516) );
  NOR2_X1 U4932 ( .A1(n2621), .A2(n5041), .ZN(n4531) );
  NOR2_X1 U4933 ( .A1(n4420), .A2(n4419), .ZN(n4525) );
  INV_X1 U4934 ( .A(n4525), .ZN(n5105) );
  NAND2_X1 U4935 ( .A1(n5105), .A2(n4421), .ZN(n4423) );
  OAI211_X1 U4936 ( .C1(n4531), .C2(n4423), .A(n4422), .B(n3483), .ZN(n4426)
         );
  NAND3_X1 U4937 ( .A1(n4426), .A2(n4425), .A3(n4424), .ZN(n4429) );
  NAND3_X1 U4938 ( .A1(n4429), .A2(n4428), .A3(n4427), .ZN(n4431) );
  NAND4_X1 U4939 ( .A1(n4432), .A2(n4431), .A3(n4451), .A4(n4430), .ZN(n4435)
         );
  NAND3_X1 U4940 ( .A1(n4435), .A2(n4434), .A3(n4433), .ZN(n4441) );
  AND2_X1 U4941 ( .A1(n4437), .A2(n4436), .ZN(n4453) );
  INV_X1 U4942 ( .A(n4438), .ZN(n4440) );
  AOI211_X1 U4943 ( .C1(n4441), .C2(n4453), .A(n4440), .B(n4439), .ZN(n4448)
         );
  INV_X1 U4944 ( .A(n4452), .ZN(n4447) );
  NAND2_X1 U4945 ( .A1(n4443), .A2(n4442), .ZN(n4510) );
  AND2_X1 U4946 ( .A1(n4445), .A2(n4444), .ZN(n4446) );
  NAND2_X1 U4947 ( .A1(n4458), .A2(n4446), .ZN(n4449) );
  NOR4_X1 U4948 ( .A1(n4448), .A2(n4447), .A3(n4510), .A4(n4449), .ZN(n4468)
         );
  INV_X1 U4949 ( .A(n4449), .ZN(n4465) );
  INV_X1 U4950 ( .A(n5155), .ZN(n4450) );
  NAND4_X1 U4951 ( .A1(n4452), .A2(n4451), .A3(n4450), .A4(n5192), .ZN(n4456)
         );
  INV_X1 U4952 ( .A(n4453), .ZN(n4455) );
  OAI21_X1 U4953 ( .B1(n4456), .B2(n4455), .A(n4454), .ZN(n4464) );
  NAND3_X1 U4954 ( .A1(n4507), .A2(n4509), .A3(n4457), .ZN(n4463) );
  INV_X1 U4955 ( .A(n4458), .ZN(n4459) );
  AOI21_X1 U4956 ( .B1(n4461), .B2(n4460), .A(n4459), .ZN(n4462) );
  AOI211_X1 U4957 ( .C1(n4465), .C2(n4464), .A(n4463), .B(n4462), .ZN(n4466)
         );
  AOI21_X1 U4958 ( .B1(n4509), .B2(n4510), .A(n4466), .ZN(n4467) );
  NOR2_X1 U4959 ( .A1(n4468), .A2(n4467), .ZN(n4473) );
  NOR4_X1 U4960 ( .A1(n4545), .A2(n4471), .A3(n4470), .A4(n4469), .ZN(n4514)
         );
  INV_X1 U4961 ( .A(n4514), .ZN(n4472) );
  AOI21_X1 U4962 ( .B1(n4473), .B2(n4506), .A(n4472), .ZN(n4484) );
  AND2_X1 U4963 ( .A1(n4478), .A2(n4474), .ZN(n4697) );
  OAI211_X1 U4964 ( .C1(n4545), .C2(n4476), .A(n4697), .B(n4475), .ZN(n4512)
         );
  NAND2_X1 U4965 ( .A1(n4478), .A2(n4477), .ZN(n4482) );
  NAND2_X1 U4966 ( .A1(n4839), .A2(n4716), .ZN(n4479) );
  AND2_X1 U4967 ( .A1(n4480), .A2(n4479), .ZN(n4481) );
  NAND2_X1 U4968 ( .A1(n4482), .A2(n4481), .ZN(n4696) );
  INV_X1 U4969 ( .A(n4696), .ZN(n4483) );
  OAI21_X1 U4970 ( .B1(n4484), .B2(n4512), .A(n4483), .ZN(n4485) );
  OR2_X1 U4971 ( .A1(n4823), .A2(n4724), .ZN(n4546) );
  NAND2_X1 U4972 ( .A1(n4720), .A2(n4822), .ZN(n4801) );
  NAND2_X1 U4973 ( .A1(n4546), .A2(n4801), .ZN(n4701) );
  AOI21_X1 U4974 ( .B1(n4516), .B2(n4485), .A(n4701), .ZN(n4487) );
  NAND2_X1 U4975 ( .A1(n4823), .A2(n4724), .ZN(n4781) );
  NAND2_X1 U4976 ( .A1(n4761), .A2(n4791), .ZN(n4529) );
  NAND2_X1 U4977 ( .A1(n4781), .A2(n4529), .ZN(n4703) );
  AND2_X1 U4978 ( .A1(n4787), .A2(n4770), .ZN(n4527) );
  AND2_X1 U4979 ( .A1(n4809), .A2(n4785), .ZN(n4702) );
  NAND2_X1 U4980 ( .A1(n4768), .A2(n4744), .ZN(n4523) );
  NAND2_X1 U4981 ( .A1(n2872), .A2(DATAI_29_), .ZN(n4732) );
  NAND2_X1 U4982 ( .A1(n4750), .A2(n4732), .ZN(n4486) );
  NAND2_X1 U4983 ( .A1(n4523), .A2(n4486), .ZN(n4497) );
  NOR3_X1 U4984 ( .A1(n4527), .A2(n4702), .A3(n4497), .ZN(n4518) );
  OAI21_X1 U4985 ( .B1(n4487), .B2(n4703), .A(n4518), .ZN(n4505) );
  INV_X1 U4986 ( .A(n4732), .ZN(n4734) );
  INV_X1 U4987 ( .A(n4750), .ZN(n4499) );
  NAND2_X1 U4988 ( .A1(n2865), .A2(REG1_REG_31__SCAN_IN), .ZN(n4490) );
  NAND2_X1 U4989 ( .A1(n3293), .A2(REG2_REG_31__SCAN_IN), .ZN(n4489) );
  NAND2_X1 U4990 ( .A1(n2497), .A2(REG0_REG_31__SCAN_IN), .ZN(n4488) );
  NAND3_X1 U4991 ( .A1(n4490), .A2(n4489), .A3(n4488), .ZN(n5310) );
  NAND2_X1 U4992 ( .A1(n4491), .A2(DATAI_31_), .ZN(n5320) );
  NAND2_X1 U4993 ( .A1(n5310), .A2(n5320), .ZN(n4503) );
  NAND2_X1 U4994 ( .A1(n2865), .A2(REG1_REG_30__SCAN_IN), .ZN(n4494) );
  NAND2_X1 U4995 ( .A1(n3293), .A2(REG2_REG_30__SCAN_IN), .ZN(n4493) );
  NAND2_X1 U4996 ( .A1(n2497), .A2(REG0_REG_30__SCAN_IN), .ZN(n4492) );
  NAND3_X1 U4997 ( .A1(n4494), .A2(n4493), .A3(n4492), .ZN(n4713) );
  NAND2_X1 U4998 ( .A1(n2872), .A2(DATAI_30_), .ZN(n5323) );
  OR2_X1 U4999 ( .A1(n4713), .A2(n5323), .ZN(n4495) );
  NAND2_X1 U5000 ( .A1(n4503), .A2(n4495), .ZN(n4524) );
  NAND2_X1 U5001 ( .A1(n4729), .A2(n4751), .ZN(n4706) );
  NAND2_X1 U5002 ( .A1(n4745), .A2(n4496), .ZN(n4704) );
  AOI21_X1 U5003 ( .B1(n4706), .B2(n4704), .A(n4497), .ZN(n4498) );
  AOI211_X1 U5004 ( .C1(n4734), .C2(n4499), .A(n4524), .B(n4498), .ZN(n4520)
         );
  INV_X1 U5005 ( .A(n5310), .ZN(n4500) );
  INV_X1 U5006 ( .A(n5320), .ZN(n5326) );
  NAND2_X1 U5007 ( .A1(n4500), .A2(n5326), .ZN(n4502) );
  NAND2_X1 U5008 ( .A1(n4713), .A2(n5323), .ZN(n4501) );
  AND2_X1 U5009 ( .A1(n4502), .A2(n4501), .ZN(n4557) );
  INV_X1 U5010 ( .A(n4557), .ZN(n4504) );
  AOI22_X1 U5011 ( .A1(n4505), .A2(n4520), .B1(n4504), .B2(n4503), .ZN(n4569)
         );
  INV_X1 U5012 ( .A(n4506), .ZN(n4515) );
  INV_X1 U5013 ( .A(n4507), .ZN(n4508) );
  NOR2_X1 U5014 ( .A1(n4192), .A2(n4508), .ZN(n4511) );
  OAI21_X1 U5015 ( .B1(n4511), .B2(n4510), .A(n4509), .ZN(n4513) );
  AOI221_X1 U5016 ( .B1(n4515), .B2(n4514), .C1(n4513), .C2(n4514), .A(n4512), 
        .ZN(n4517) );
  AOI221_X1 U5017 ( .B1(n4517), .B2(n4516), .C1(n4696), .C2(n4516), .A(n4701), 
        .ZN(n4519) );
  OAI21_X1 U5018 ( .B1(n4519), .B2(n4703), .A(n4518), .ZN(n4521) );
  OAI211_X1 U5019 ( .C1(n5310), .C2(n5323), .A(n4521), .B(n4520), .ZN(n4522)
         );
  OAI211_X1 U5020 ( .C1(n4557), .C2(n5320), .A(n4522), .B(n5041), .ZN(n4566)
         );
  INV_X1 U5021 ( .A(n4742), .ZN(n4747) );
  NOR4_X1 U5022 ( .A1(n4526), .A2(n4747), .A3(n4525), .A4(n4524), .ZN(n4532)
         );
  INV_X1 U5023 ( .A(n4527), .ZN(n4528) );
  NAND2_X1 U5024 ( .A1(n4528), .A2(n4704), .ZN(n4764) );
  INV_X1 U5025 ( .A(n4529), .ZN(n4530) );
  NAND4_X1 U5026 ( .A1(n4532), .A2(n2666), .A3(n4783), .A4(n4531), .ZN(n4543)
         );
  XNOR2_X1 U5027 ( .A(n4840), .B(n4867), .ZN(n4859) );
  NAND4_X1 U5028 ( .A1(n4536), .A2(n4535), .A3(n4534), .A4(n4533), .ZN(n4542)
         );
  INV_X1 U5029 ( .A(n3482), .ZN(n4539) );
  NAND4_X1 U5030 ( .A1(n4540), .A2(n4539), .A3(n4538), .A4(n4537), .ZN(n4541)
         );
  NOR4_X1 U5031 ( .A1(n4543), .A2(n4859), .A3(n4542), .A4(n4541), .ZN(n4564)
         );
  INV_X1 U5032 ( .A(n4900), .ZN(n4563) );
  INV_X1 U5033 ( .A(n5184), .ZN(n5179) );
  OR2_X1 U5034 ( .A1(n4545), .A2(n4544), .ZN(n4873) );
  INV_X1 U5035 ( .A(n4873), .ZN(n4875) );
  NAND2_X1 U5036 ( .A1(n4546), .A2(n4781), .ZN(n4804) );
  INV_X1 U5037 ( .A(n5153), .ZN(n4552) );
  INV_X1 U5038 ( .A(n4547), .ZN(n4549) );
  NOR4_X1 U5039 ( .A1(n4550), .A2(n4549), .A3(n4548), .A4(n4889), .ZN(n4551)
         );
  NAND3_X1 U5040 ( .A1(n4553), .A2(n4552), .A3(n4551), .ZN(n4554) );
  NOR4_X1 U5041 ( .A1(n4555), .A2(n4804), .A3(n4933), .A4(n4554), .ZN(n4556)
         );
  NAND4_X1 U5042 ( .A1(n4875), .A2(n4960), .A3(n4557), .A4(n4556), .ZN(n4561)
         );
  XOR2_X1 U5043 ( .A(n4732), .B(n4750), .Z(n4730) );
  INV_X1 U5044 ( .A(n4730), .ZN(n4560) );
  XNOR2_X1 U5045 ( .A(n4720), .B(n4827), .ZN(n4819) );
  INV_X1 U5046 ( .A(n4819), .ZN(n4559) );
  NOR4_X1 U5047 ( .A1(n4561), .A2(n4560), .A3(n4559), .A4(n4558), .ZN(n4562)
         );
  NAND4_X1 U5048 ( .A1(n4564), .A2(n4563), .A3(n5179), .A4(n4562), .ZN(n4565)
         );
  NAND2_X1 U5049 ( .A1(n4566), .A2(n4565), .ZN(n4568) );
  MUX2_X1 U5050 ( .A(n4569), .B(n4568), .S(n4567), .Z(n4570) );
  XNOR2_X1 U5051 ( .A(n4570), .B(n5114), .ZN(n4578) );
  INV_X1 U5052 ( .A(n4571), .ZN(n4574) );
  NOR3_X1 U5053 ( .A1(n4574), .A2(n4573), .A3(n4572), .ZN(n4576) );
  OAI21_X1 U5054 ( .B1(n4577), .B2(n5040), .A(B_REG_SCAN_IN), .ZN(n4575) );
  OAI22_X1 U5055 ( .A1(n4578), .A2(n4577), .B1(n4576), .B2(n4575), .ZN(U3239)
         );
  MUX2_X1 U5056 ( .A(n5310), .B(DATAO_REG_31__SCAN_IN), .S(n4592), .Z(U3581)
         );
  MUX2_X1 U5057 ( .A(n4713), .B(DATAO_REG_30__SCAN_IN), .S(n4592), .Z(U3580)
         );
  MUX2_X1 U5058 ( .A(n4750), .B(DATAO_REG_29__SCAN_IN), .S(n4592), .Z(U3579)
         );
  MUX2_X1 U5059 ( .A(DATAO_REG_28__SCAN_IN), .B(n4768), .S(U4043), .Z(U3578)
         );
  MUX2_X1 U5060 ( .A(n4787), .B(DATAO_REG_27__SCAN_IN), .S(n4592), .Z(U3577)
         );
  MUX2_X1 U5061 ( .A(n4809), .B(DATAO_REG_26__SCAN_IN), .S(n4592), .Z(U3576)
         );
  MUX2_X1 U5062 ( .A(DATAO_REG_25__SCAN_IN), .B(n4725), .S(U4043), .Z(U3575)
         );
  MUX2_X1 U5063 ( .A(n4720), .B(DATAO_REG_24__SCAN_IN), .S(n4592), .Z(U3574)
         );
  MUX2_X1 U5064 ( .A(n4839), .B(DATAO_REG_23__SCAN_IN), .S(n4592), .Z(U3573)
         );
  MUX2_X1 U5065 ( .A(DATAO_REG_22__SCAN_IN), .B(n4579), .S(U4043), .Z(U3572)
         );
  MUX2_X1 U5066 ( .A(n4840), .B(DATAO_REG_21__SCAN_IN), .S(n4592), .Z(U3571)
         );
  MUX2_X1 U5067 ( .A(DATAO_REG_20__SCAN_IN), .B(n4892), .S(U4043), .Z(U3570)
         );
  MUX2_X1 U5068 ( .A(n4580), .B(DATAO_REG_19__SCAN_IN), .S(n4592), .Z(U3569)
         );
  MUX2_X1 U5069 ( .A(n4928), .B(DATAO_REG_18__SCAN_IN), .S(n4592), .Z(U3568)
         );
  MUX2_X1 U5070 ( .A(n4949), .B(DATAO_REG_17__SCAN_IN), .S(n4592), .Z(U3567)
         );
  MUX2_X1 U5071 ( .A(n4929), .B(DATAO_REG_16__SCAN_IN), .S(n4592), .Z(U3566)
         );
  MUX2_X1 U5072 ( .A(DATAO_REG_15__SCAN_IN), .B(n4950), .S(U4043), .Z(U3565)
         );
  MUX2_X1 U5073 ( .A(DATAO_REG_14__SCAN_IN), .B(n4581), .S(U4043), .Z(U3564)
         );
  MUX2_X1 U5074 ( .A(DATAO_REG_13__SCAN_IN), .B(n4582), .S(U4043), .Z(U3563)
         );
  MUX2_X1 U5075 ( .A(DATAO_REG_12__SCAN_IN), .B(n4583), .S(U4043), .Z(U3562)
         );
  MUX2_X1 U5076 ( .A(DATAO_REG_11__SCAN_IN), .B(n4584), .S(U4043), .Z(U3561)
         );
  MUX2_X1 U5077 ( .A(DATAO_REG_10__SCAN_IN), .B(n4585), .S(U4043), .Z(U3560)
         );
  MUX2_X1 U5078 ( .A(DATAO_REG_9__SCAN_IN), .B(n4586), .S(U4043), .Z(U3559) );
  MUX2_X1 U5079 ( .A(n4587), .B(DATAO_REG_8__SCAN_IN), .S(n4592), .Z(U3558) );
  MUX2_X1 U5080 ( .A(DATAO_REG_7__SCAN_IN), .B(n4588), .S(U4043), .Z(U3557) );
  MUX2_X1 U5081 ( .A(n4589), .B(DATAO_REG_6__SCAN_IN), .S(n4592), .Z(U3556) );
  MUX2_X1 U5082 ( .A(n5155), .B(DATAO_REG_5__SCAN_IN), .S(n4592), .Z(U3555) );
  MUX2_X1 U5083 ( .A(DATAO_REG_4__SCAN_IN), .B(n4590), .S(U4043), .Z(U3554) );
  MUX2_X1 U5084 ( .A(n5156), .B(DATAO_REG_3__SCAN_IN), .S(n4592), .Z(U3553) );
  MUX2_X1 U5085 ( .A(DATAO_REG_2__SCAN_IN), .B(n4591), .S(U4043), .Z(U3552) );
  MUX2_X1 U5086 ( .A(DATAO_REG_1__SCAN_IN), .B(n3457), .S(U4043), .Z(U3551) );
  MUX2_X1 U5087 ( .A(n4593), .B(DATAO_REG_0__SCAN_IN), .S(n4592), .Z(U3550) );
  INV_X1 U5088 ( .A(REG1_REG_13__SCAN_IN), .ZN(n5259) );
  NOR2_X1 U5089 ( .A1(n4614), .A2(n5259), .ZN(n4597) );
  NAND2_X1 U5090 ( .A1(n5048), .A2(n4594), .ZN(n4596) );
  NAND2_X1 U5091 ( .A1(n4596), .A2(n4595), .ZN(n4598) );
  NOR2_X1 U5092 ( .A1(n4614), .A2(REG1_REG_13__SCAN_IN), .ZN(n4599) );
  AOI211_X1 U5093 ( .C1(n4614), .C2(REG1_REG_13__SCAN_IN), .A(n4599), .B(n4598), .ZN(n4600) );
  OR3_X1 U5094 ( .A1(n4615), .A2(n4600), .A3(n4671), .ZN(n4613) );
  NOR2_X1 U5095 ( .A1(n4602), .A2(n4601), .ZN(n4604) );
  INV_X1 U5096 ( .A(n4614), .ZN(n5047) );
  NAND2_X1 U5097 ( .A1(n5047), .A2(n4152), .ZN(n4606) );
  NAND2_X1 U5098 ( .A1(n4614), .A2(REG2_REG_13__SCAN_IN), .ZN(n4605) );
  AND2_X1 U5099 ( .A1(n4606), .A2(n4605), .ZN(n4608) );
  INV_X1 U5100 ( .A(n4620), .ZN(n4607) );
  AOI211_X1 U5101 ( .C1(n4609), .C2(n4608), .A(n4607), .B(n5090), .ZN(n4611)
         );
  AOI211_X1 U5102 ( .C1(n5088), .C2(ADDR_REG_13__SCAN_IN), .A(n4611), .B(n4610), .ZN(n4612) );
  OAI211_X1 U5103 ( .C1(n5089), .C2(n4614), .A(n4613), .B(n4612), .ZN(U3253)
         );
  XNOR2_X1 U5104 ( .A(n4634), .B(REG1_REG_14__SCAN_IN), .ZN(n4626) );
  AOI21_X1 U5105 ( .B1(n5088), .B2(ADDR_REG_14__SCAN_IN), .A(n4617), .ZN(n4618) );
  OAI21_X1 U5106 ( .B1(n2717), .B2(n5089), .A(n4618), .ZN(n4625) );
  NAND2_X1 U5107 ( .A1(n5047), .A2(REG2_REG_13__SCAN_IN), .ZN(n4619) );
  AOI211_X1 U5108 ( .C1(n4623), .C2(n4622), .A(n4628), .B(n5090), .ZN(n4624)
         );
  AOI211_X1 U5109 ( .C1(n5099), .C2(n4626), .A(n4625), .B(n4624), .ZN(n4627)
         );
  INV_X1 U5110 ( .A(n4627), .ZN(U3254) );
  AOI22_X1 U5111 ( .A1(n5045), .A2(n4630), .B1(REG2_REG_15__SCAN_IN), .B2(
        n4648), .ZN(n4631) );
  NOR2_X1 U5112 ( .A1(n4632), .A2(n4631), .ZN(n4644) );
  AOI211_X1 U5113 ( .C1(n4632), .C2(n4631), .A(n4644), .B(n5090), .ZN(n4643)
         );
  INV_X1 U5114 ( .A(REG1_REG_14__SCAN_IN), .ZN(n4633) );
  NOR2_X1 U5115 ( .A1(n5045), .A2(REG1_REG_15__SCAN_IN), .ZN(n4636) );
  AOI21_X1 U5116 ( .B1(REG1_REG_15__SCAN_IN), .B2(n5045), .A(n4636), .ZN(n4637) );
  NAND2_X1 U5117 ( .A1(n4637), .A2(n4638), .ZN(n4647) );
  OAI211_X1 U5118 ( .C1(n4638), .C2(n4637), .A(n5099), .B(n4647), .ZN(n4641)
         );
  NOR2_X1 U5119 ( .A1(STATE_REG_SCAN_IN), .A2(n4639), .ZN(n5275) );
  AOI21_X1 U5120 ( .B1(n5088), .B2(ADDR_REG_15__SCAN_IN), .A(n5275), .ZN(n4640) );
  OAI211_X1 U5121 ( .C1(n5089), .C2(n4648), .A(n4641), .B(n4640), .ZN(n4642)
         );
  OR2_X1 U5122 ( .A1(n4643), .A2(n4642), .ZN(U3255) );
  INV_X1 U5123 ( .A(REG2_REG_16__SCAN_IN), .ZN(n4959) );
  AOI221_X1 U5124 ( .B1(n4645), .B2(n4662), .C1(n4959), .C2(n4662), .A(n5090), 
        .ZN(n4646) );
  INV_X1 U5125 ( .A(n4646), .ZN(n4654) );
  INV_X1 U5126 ( .A(REG1_REG_15__SCAN_IN), .ZN(n5291) );
  OAI21_X1 U5127 ( .B1(n5291), .B2(n4648), .A(n4647), .ZN(n4655) );
  AOI21_X1 U5128 ( .B1(n4649), .B2(REG1_REG_16__SCAN_IN), .A(n4656), .ZN(n4650) );
  NOR2_X1 U5129 ( .A1(n4671), .A2(n4650), .ZN(n4651) );
  AOI211_X1 U5130 ( .C1(n5088), .C2(ADDR_REG_16__SCAN_IN), .A(n4652), .B(n4651), .ZN(n4653) );
  OAI211_X1 U5131 ( .C1(n5089), .C2(n4660), .A(n4654), .B(n4653), .ZN(U3256)
         );
  NOR2_X1 U5132 ( .A1(n5044), .A2(n4655), .ZN(n4657) );
  INV_X1 U5133 ( .A(REG1_REG_17__SCAN_IN), .ZN(n5306) );
  NOR2_X1 U5134 ( .A1(n5043), .A2(n5306), .ZN(n4658) );
  AOI21_X1 U5135 ( .B1(n5306), .B2(n5043), .A(n4658), .ZN(n4659) );
  AOI21_X1 U5136 ( .B1(n2513), .B2(n4659), .A(n4678), .ZN(n4672) );
  INV_X1 U5137 ( .A(REG2_REG_17__SCAN_IN), .ZN(n4941) );
  AOI22_X1 U5138 ( .A1(n5043), .A2(n4941), .B1(REG2_REG_17__SCAN_IN), .B2(
        n4679), .ZN(n4665) );
  NAND2_X1 U5139 ( .A1(n4661), .A2(n4660), .ZN(n4663) );
  NOR2_X1 U5140 ( .A1(n4665), .A2(n4664), .ZN(n4673) );
  AOI211_X1 U5141 ( .C1(n4665), .C2(n4664), .A(n4673), .B(n5090), .ZN(n4666)
         );
  INV_X1 U5142 ( .A(n4666), .ZN(n4670) );
  NOR2_X1 U5143 ( .A1(n5089), .A2(n4679), .ZN(n4667) );
  AOI211_X1 U5144 ( .C1(n5088), .C2(ADDR_REG_17__SCAN_IN), .A(n4668), .B(n4667), .ZN(n4669) );
  OAI211_X1 U5145 ( .C1(n4672), .C2(n4671), .A(n4670), .B(n4669), .ZN(U3257)
         );
  INV_X1 U5146 ( .A(REG2_REG_18__SCAN_IN), .ZN(n4674) );
  AOI22_X1 U5147 ( .A1(n5042), .A2(n4674), .B1(REG2_REG_18__SCAN_IN), .B2(
        n4684), .ZN(n4675) );
  AOI211_X1 U5148 ( .C1(n4676), .C2(n4675), .A(n4687), .B(n5090), .ZN(n4686)
         );
  AOI21_X1 U5149 ( .B1(n5088), .B2(ADDR_REG_18__SCAN_IN), .A(n4677), .ZN(n4683) );
  XNOR2_X1 U5150 ( .A(n4684), .B(REG1_REG_18__SCAN_IN), .ZN(n4681) );
  AOI21_X1 U5151 ( .B1(n4679), .B2(n5306), .A(n4678), .ZN(n4680) );
  OAI211_X1 U5152 ( .C1(n4681), .C2(n4680), .A(n5099), .B(n4690), .ZN(n4682)
         );
  OAI211_X1 U5153 ( .C1(n4684), .C2(n5089), .A(n4683), .B(n4682), .ZN(n4685)
         );
  OR2_X1 U5154 ( .A1(n4686), .A2(n4685), .ZN(U3258) );
  INV_X1 U5155 ( .A(REG2_REG_19__SCAN_IN), .ZN(n4688) );
  MUX2_X1 U5156 ( .A(n4688), .B(REG2_REG_19__SCAN_IN), .S(n5202), .Z(n4689) );
  INV_X1 U5157 ( .A(n5090), .ZN(n4691) );
  AOI21_X1 U5158 ( .B1(n5088), .B2(ADDR_REG_19__SCAN_IN), .A(n4693), .ZN(n4694) );
  OAI211_X1 U5159 ( .C1(n5202), .C2(n5089), .A(n4695), .B(n4694), .ZN(U3259)
         );
  INV_X1 U5160 ( .A(n4704), .ZN(n4705) );
  NOR2_X1 U5161 ( .A1(n4748), .A2(n4747), .ZN(n4746) );
  INV_X1 U5162 ( .A(n4706), .ZN(n4707) );
  NOR2_X1 U5163 ( .A1(n4746), .A2(n4707), .ZN(n4708) );
  XNOR2_X1 U5164 ( .A(n4708), .B(n4730), .ZN(n4715) );
  INV_X1 U5165 ( .A(B_REG_SCAN_IN), .ZN(n4709) );
  NOR2_X1 U5166 ( .A1(n4710), .A2(n4709), .ZN(n4711) );
  NOR2_X1 U5167 ( .A1(n5188), .A2(n4711), .ZN(n5309) );
  OAI22_X1 U5168 ( .A1(n4729), .A2(n5186), .B1(n4732), .B2(n5319), .ZN(n4712)
         );
  AOI21_X1 U5169 ( .B1(n5309), .B2(n4713), .A(n4712), .ZN(n4714) );
  OAI21_X1 U5170 ( .B1(n4715), .B2(n5194), .A(n4714), .ZN(n4971) );
  INV_X1 U5171 ( .A(n4971), .ZN(n4741) );
  NAND2_X1 U5172 ( .A1(n4821), .A2(n4716), .ZN(n4718) );
  NOR2_X1 U5173 ( .A1(n4821), .A2(n4716), .ZN(n4717) );
  AOI21_X2 U5174 ( .B1(n4719), .B2(n4718), .A(n4717), .ZN(n4818) );
  NAND2_X1 U5175 ( .A1(n4720), .A2(n4827), .ZN(n4721) );
  NAND2_X1 U5176 ( .A1(n4818), .A2(n4721), .ZN(n4723) );
  NAND2_X1 U5177 ( .A1(n4800), .A2(n4822), .ZN(n4722) );
  NAND2_X1 U5178 ( .A1(n4723), .A2(n4722), .ZN(n4799) );
  NOR2_X1 U5179 ( .A1(n4725), .A2(n4724), .ZN(n4727) );
  NAND2_X1 U5180 ( .A1(n4725), .A2(n4724), .ZN(n4726) );
  OAI21_X1 U5181 ( .B1(n4799), .B2(n4727), .A(n4726), .ZN(n4777) );
  NAND2_X1 U5182 ( .A1(n4761), .A2(n4785), .ZN(n4728) );
  XNOR2_X1 U5183 ( .A(n4731), .B(n4730), .ZN(n4969) );
  NAND2_X1 U5184 ( .A1(n4969), .A2(n4935), .ZN(n4740) );
  AND2_X2 U5185 ( .A1(n4830), .A2(n4810), .ZN(n4812) );
  AOI21_X1 U5186 ( .B1(n4752), .B2(n4734), .A(n5264), .ZN(n4735) );
  AND2_X1 U5187 ( .A1(n5325), .A2(n4735), .ZN(n4970) );
  INV_X1 U5188 ( .A(REG2_REG_29__SCAN_IN), .ZN(n4737) );
  OAI22_X1 U5189 ( .A1(n5208), .A2(n4737), .B1(n4736), .B2(n5210), .ZN(n4738)
         );
  AOI21_X1 U5190 ( .B1(n4970), .B2(n4943), .A(n4738), .ZN(n4739) );
  OAI211_X1 U5191 ( .C1(n4741), .C2(n5330), .A(n4740), .B(n4739), .ZN(U3354)
         );
  OAI22_X1 U5192 ( .A1(n4745), .A2(n5186), .B1(n5319), .B2(n4744), .ZN(n4749)
         );
  INV_X1 U5193 ( .A(n4980), .ZN(n4757) );
  AOI21_X1 U5194 ( .B1(n4769), .B2(n4751), .A(n5264), .ZN(n4753) );
  NAND2_X1 U5195 ( .A1(n4753), .A2(n4752), .ZN(n4979) );
  AOI22_X1 U5196 ( .A1(n5330), .A2(REG2_REG_28__SCAN_IN), .B1(n4754), .B2(
        n5118), .ZN(n4755) );
  OAI21_X1 U5197 ( .B1(n4979), .B2(n4922), .A(n4755), .ZN(n4756) );
  AOI21_X1 U5198 ( .B1(n4757), .B2(n5208), .A(n4756), .ZN(n4758) );
  OAI21_X1 U5199 ( .B1(n4981), .B2(n4962), .A(n4758), .ZN(U3262) );
  OAI21_X1 U5200 ( .B1(n4760), .B2(n4764), .A(n4759), .ZN(n4982) );
  OAI22_X1 U5201 ( .A1(n4761), .A2(n5186), .B1(n5319), .B2(n4770), .ZN(n4767)
         );
  AOI21_X1 U5202 ( .B1(n4764), .B2(n4763), .A(n4762), .ZN(n4765) );
  NOR2_X1 U5203 ( .A1(n4765), .A2(n5194), .ZN(n4766) );
  AOI211_X1 U5204 ( .C1(n5154), .C2(n4768), .A(n4767), .B(n4766), .ZN(n4983)
         );
  NOR2_X1 U5205 ( .A1(n4983), .A2(n5330), .ZN(n4775) );
  OAI21_X1 U5206 ( .B1(n4771), .B2(n4770), .A(n4769), .ZN(n4985) );
  AOI22_X1 U5207 ( .A1(n5330), .A2(REG2_REG_27__SCAN_IN), .B1(n4772), .B2(
        n5118), .ZN(n4773) );
  OAI21_X1 U5208 ( .B1(n4985), .B2(n4904), .A(n4773), .ZN(n4774) );
  AOI211_X1 U5209 ( .C1(n4982), .C2(n4935), .A(n4775), .B(n4774), .ZN(n4776)
         );
  INV_X1 U5210 ( .A(n4776), .ZN(U3263) );
  INV_X1 U5211 ( .A(n4777), .ZN(n4780) );
  INV_X1 U5212 ( .A(n4783), .ZN(n4779) );
  OAI21_X1 U5213 ( .B1(n4780), .B2(n4779), .A(n4778), .ZN(n4794) );
  INV_X1 U5214 ( .A(n4781), .ZN(n4782) );
  NOR2_X1 U5215 ( .A1(n2512), .A2(n4782), .ZN(n4784) );
  XNOR2_X1 U5216 ( .A(n4784), .B(n4783), .ZN(n4789) );
  OAI22_X1 U5217 ( .A1(n4823), .A2(n5186), .B1(n4785), .B2(n5319), .ZN(n4786)
         );
  AOI21_X1 U5218 ( .B1(n5154), .B2(n4787), .A(n4786), .ZN(n4788) );
  OAI21_X1 U5219 ( .B1(n4789), .B2(n5194), .A(n4788), .ZN(n4790) );
  AOI21_X1 U5220 ( .B1(n4794), .B2(n5163), .A(n4790), .ZN(n4988) );
  XNOR2_X1 U5221 ( .A(n4812), .B(n4791), .ZN(n4986) );
  INV_X1 U5222 ( .A(REG2_REG_26__SCAN_IN), .ZN(n4793) );
  OAI22_X1 U5223 ( .A1(n5208), .A2(n4793), .B1(n4792), .B2(n5210), .ZN(n4797)
         );
  INV_X1 U5224 ( .A(n4794), .ZN(n4989) );
  NOR2_X1 U5225 ( .A1(n4989), .A2(n4795), .ZN(n4796) );
  AOI211_X1 U5226 ( .C1(n5328), .C2(n4986), .A(n4797), .B(n4796), .ZN(n4798)
         );
  OAI21_X1 U5227 ( .B1(n5330), .B2(n4988), .A(n4798), .ZN(U3264) );
  XOR2_X1 U5228 ( .A(n4804), .B(n4799), .Z(n4992) );
  OAI22_X1 U5229 ( .A1(n4800), .A2(n5186), .B1(n4810), .B2(n5319), .ZN(n4808)
         );
  INV_X1 U5230 ( .A(n4801), .ZN(n4802) );
  NOR2_X1 U5231 ( .A1(n4803), .A2(n4802), .ZN(n4805) );
  XNOR2_X1 U5232 ( .A(n4805), .B(n4804), .ZN(n4806) );
  NOR2_X1 U5233 ( .A1(n4806), .A2(n5194), .ZN(n4807) );
  AOI211_X1 U5234 ( .C1(n5154), .C2(n4809), .A(n4808), .B(n4807), .ZN(n4991)
         );
  INV_X1 U5235 ( .A(n4991), .ZN(n4816) );
  OAI21_X1 U5236 ( .B1(n4830), .B2(n4810), .A(n5333), .ZN(n4811) );
  OR2_X1 U5237 ( .A1(n4812), .A2(n4811), .ZN(n4990) );
  AOI22_X1 U5238 ( .A1(n5330), .A2(REG2_REG_25__SCAN_IN), .B1(n4813), .B2(
        n5118), .ZN(n4814) );
  OAI21_X1 U5239 ( .B1(n4990), .B2(n4922), .A(n4814), .ZN(n4815) );
  AOI21_X1 U5240 ( .B1(n4816), .B2(n5208), .A(n4815), .ZN(n4817) );
  OAI21_X1 U5241 ( .B1(n4992), .B2(n4962), .A(n4817), .ZN(U3265) );
  XNOR2_X1 U5242 ( .A(n4818), .B(n4819), .ZN(n4995) );
  XNOR2_X1 U5243 ( .A(n4820), .B(n4819), .ZN(n4826) );
  NOR2_X1 U5244 ( .A1(n4821), .A2(n5186), .ZN(n4825) );
  OAI22_X1 U5245 ( .A1(n4823), .A2(n5188), .B1(n5319), .B2(n4822), .ZN(n4824)
         );
  AOI211_X1 U5246 ( .C1(n4826), .C2(n5108), .A(n4825), .B(n4824), .ZN(n4994)
         );
  INV_X1 U5247 ( .A(n4994), .ZN(n4835) );
  NAND2_X1 U5248 ( .A1(n4828), .A2(n4827), .ZN(n4829) );
  NAND2_X1 U5249 ( .A1(n4829), .A2(n5333), .ZN(n4831) );
  OR2_X1 U5250 ( .A1(n4831), .A2(n4830), .ZN(n4993) );
  AOI22_X1 U5251 ( .A1(n5330), .A2(REG2_REG_24__SCAN_IN), .B1(n4832), .B2(
        n5118), .ZN(n4833) );
  OAI21_X1 U5252 ( .B1(n4993), .B2(n4922), .A(n4833), .ZN(n4834) );
  AOI21_X1 U5253 ( .B1(n4835), .B2(n5208), .A(n4834), .ZN(n4836) );
  OAI21_X1 U5254 ( .B1(n4995), .B2(n4962), .A(n4836), .ZN(U3266) );
  OAI21_X1 U5255 ( .B1(n4850), .B2(n4838), .A(n4837), .ZN(n4844) );
  NAND2_X1 U5256 ( .A1(n4839), .A2(n5154), .ZN(n4842) );
  NAND2_X1 U5257 ( .A1(n4840), .A2(n5157), .ZN(n4841) );
  OAI211_X1 U5258 ( .C1(n5319), .C2(n4852), .A(n4842), .B(n4841), .ZN(n4843)
         );
  AOI21_X1 U5259 ( .B1(n4844), .B2(n5108), .A(n4843), .ZN(n5002) );
  NAND2_X1 U5260 ( .A1(n4845), .A2(n4846), .ZN(n4858) );
  OR2_X1 U5261 ( .A1(n4858), .A2(n4847), .ZN(n4849) );
  NAND2_X1 U5262 ( .A1(n4849), .A2(n4848), .ZN(n4851) );
  NAND2_X1 U5263 ( .A1(n4851), .A2(n4850), .ZN(n4999) );
  NAND3_X1 U5264 ( .A1(n5000), .A2(n4999), .A3(n4935), .ZN(n4857) );
  OAI211_X1 U5265 ( .C1(n2592), .C2(n4852), .A(n5333), .B(n2500), .ZN(n5001)
         );
  AOI22_X1 U5266 ( .A1(n5330), .A2(REG2_REG_22__SCAN_IN), .B1(n4853), .B2(
        n5118), .ZN(n4854) );
  OAI21_X1 U5267 ( .B1(n5001), .B2(n4922), .A(n4854), .ZN(n4855) );
  INV_X1 U5268 ( .A(n4855), .ZN(n4856) );
  OAI211_X1 U5269 ( .C1(n5330), .C2(n5002), .A(n4857), .B(n4856), .ZN(U3268)
         );
  XNOR2_X1 U5270 ( .A(n4858), .B(n4859), .ZN(n5006) );
  XNOR2_X1 U5271 ( .A(n4860), .B(n4859), .ZN(n4865) );
  NOR2_X1 U5272 ( .A1(n4861), .A2(n5188), .ZN(n4864) );
  OAI22_X1 U5273 ( .A1(n4862), .A2(n5186), .B1(n4867), .B2(n5319), .ZN(n4863)
         );
  AOI211_X1 U5274 ( .C1(n4865), .C2(n5108), .A(n4864), .B(n4863), .ZN(n5005)
         );
  INV_X1 U5275 ( .A(n5005), .ZN(n4871) );
  OAI211_X1 U5276 ( .C1(n4882), .C2(n4867), .A(n5333), .B(n4866), .ZN(n5004)
         );
  AOI22_X1 U5277 ( .A1(n5330), .A2(REG2_REG_21__SCAN_IN), .B1(n4868), .B2(
        n5118), .ZN(n4869) );
  OAI21_X1 U5278 ( .B1(n5004), .B2(n4922), .A(n4869), .ZN(n4870) );
  AOI21_X1 U5279 ( .B1(n4871), .B2(n5208), .A(n4870), .ZN(n4872) );
  OAI21_X1 U5280 ( .B1(n5006), .B2(n4962), .A(n4872), .ZN(U3269) );
  XNOR2_X1 U5281 ( .A(n4874), .B(n4873), .ZN(n5009) );
  XNOR2_X1 U5282 ( .A(n4876), .B(n4875), .ZN(n4880) );
  NOR2_X1 U5283 ( .A1(n4877), .A2(n5188), .ZN(n4879) );
  OAI22_X1 U5284 ( .A1(n4908), .A2(n5186), .B1(n4881), .B2(n5319), .ZN(n4878)
         );
  AOI211_X1 U5285 ( .C1(n4880), .C2(n5108), .A(n4879), .B(n4878), .ZN(n5008)
         );
  INV_X1 U5286 ( .A(n5008), .ZN(n4887) );
  OAI21_X1 U5287 ( .B1(n4896), .B2(n4881), .A(n5333), .ZN(n4883) );
  OR2_X1 U5288 ( .A1(n4883), .A2(n4882), .ZN(n5007) );
  AOI22_X1 U5289 ( .A1(n5330), .A2(REG2_REG_20__SCAN_IN), .B1(n4884), .B2(
        n5118), .ZN(n4885) );
  OAI21_X1 U5290 ( .B1(n5007), .B2(n4922), .A(n4885), .ZN(n4886) );
  AOI21_X1 U5291 ( .B1(n4887), .B2(n5208), .A(n4886), .ZN(n4888) );
  OAI21_X1 U5292 ( .B1(n5009), .B2(n4962), .A(n4888), .ZN(U3270) );
  NAND3_X1 U5293 ( .A1(n4911), .A2(n2653), .A3(n4910), .ZN(n4909) );
  NAND2_X1 U5294 ( .A1(n4909), .A2(n4890), .ZN(n4891) );
  XNOR2_X1 U5295 ( .A(n4891), .B(n4900), .ZN(n4895) );
  AOI22_X1 U5296 ( .A1(n4892), .A2(n5154), .B1(n5157), .B2(n4928), .ZN(n4893)
         );
  OAI21_X1 U5297 ( .B1(n4898), .B2(n5319), .A(n4893), .ZN(n4894) );
  AOI21_X1 U5298 ( .B1(n4895), .B2(n5108), .A(n4894), .ZN(n5012) );
  INV_X1 U5299 ( .A(n4917), .ZN(n4899) );
  INV_X1 U5300 ( .A(n4896), .ZN(n4897) );
  OAI21_X1 U5301 ( .B1(n4899), .B2(n4898), .A(n4897), .ZN(n5014) );
  OR2_X1 U5302 ( .A1(n2537), .A2(n4900), .ZN(n5011) );
  NAND3_X1 U5303 ( .A1(n5011), .A2(n5010), .A3(n4935), .ZN(n4903) );
  AOI22_X1 U5304 ( .A1(n5330), .A2(REG2_REG_19__SCAN_IN), .B1(n4901), .B2(
        n5118), .ZN(n4902) );
  OAI211_X1 U5305 ( .C1(n5014), .C2(n4904), .A(n4903), .B(n4902), .ZN(n4905)
         );
  INV_X1 U5306 ( .A(n4905), .ZN(n4906) );
  OAI21_X1 U5307 ( .B1(n5330), .B2(n5012), .A(n4906), .ZN(U3271) );
  XNOR2_X1 U5308 ( .A(n4907), .B(n2653), .ZN(n5017) );
  OAI22_X1 U5309 ( .A1(n4908), .A2(n5188), .B1(n4227), .B2(n5186), .ZN(n4915)
         );
  INV_X1 U5310 ( .A(n4909), .ZN(n4913) );
  AOI21_X1 U5311 ( .B1(n4911), .B2(n4910), .A(n2653), .ZN(n4912) );
  NOR3_X1 U5312 ( .A1(n4913), .A2(n4912), .A3(n5194), .ZN(n4914) );
  AOI211_X1 U5313 ( .C1(n5191), .C2(n4916), .A(n4915), .B(n4914), .ZN(n5016)
         );
  INV_X1 U5314 ( .A(n5016), .ZN(n4924) );
  INV_X1 U5315 ( .A(n4938), .ZN(n4919) );
  OAI211_X1 U5316 ( .C1(n4919), .C2(n4918), .A(n5333), .B(n4917), .ZN(n5015)
         );
  AOI22_X1 U5317 ( .A1(n5330), .A2(REG2_REG_18__SCAN_IN), .B1(n4920), .B2(
        n5118), .ZN(n4921) );
  OAI21_X1 U5318 ( .B1(n5015), .B2(n4922), .A(n4921), .ZN(n4923) );
  AOI21_X1 U5319 ( .B1(n4924), .B2(n5208), .A(n4923), .ZN(n4925) );
  OAI21_X1 U5320 ( .B1(n5017), .B2(n4962), .A(n4925), .ZN(U3272) );
  INV_X1 U5321 ( .A(n4933), .ZN(n4926) );
  XNOR2_X1 U5322 ( .A(n2535), .B(n4926), .ZN(n4927) );
  NAND2_X1 U5323 ( .A1(n4927), .A2(n5108), .ZN(n4931) );
  AOI22_X1 U5324 ( .A1(n5157), .A2(n4929), .B1(n4928), .B2(n5154), .ZN(n4930)
         );
  OAI211_X1 U5325 ( .C1(n5319), .C2(n4936), .A(n4931), .B(n4930), .ZN(n5302)
         );
  INV_X1 U5326 ( .A(n5302), .ZN(n4946) );
  OAI21_X1 U5327 ( .B1(n4934), .B2(n4933), .A(n4932), .ZN(n5305) );
  NAND2_X1 U5328 ( .A1(n5305), .A2(n4935), .ZN(n4945) );
  OR2_X1 U5329 ( .A1(n4955), .A2(n4936), .ZN(n4937) );
  AND3_X1 U5330 ( .A1(n4938), .A2(n4937), .A3(n5333), .ZN(n5303) );
  INV_X1 U5331 ( .A(n4939), .ZN(n4940) );
  OAI22_X1 U5332 ( .A1(n5208), .A2(n4941), .B1(n4940), .B2(n5210), .ZN(n4942)
         );
  AOI21_X1 U5333 ( .B1(n5303), .B2(n4943), .A(n4942), .ZN(n4944) );
  OAI211_X1 U5334 ( .C1(n5330), .C2(n4946), .A(n4945), .B(n4944), .ZN(U3273)
         );
  OAI211_X1 U5335 ( .C1(n4948), .C2(n4960), .A(n4947), .B(n5108), .ZN(n4952)
         );
  AOI22_X1 U5336 ( .A1(n4950), .A2(n5157), .B1(n5154), .B2(n4949), .ZN(n4951)
         );
  OAI211_X1 U5337 ( .C1(n5319), .C2(n4953), .A(n4952), .B(n4951), .ZN(n5298)
         );
  INV_X1 U5338 ( .A(n5298), .ZN(n4966) );
  INV_X1 U5339 ( .A(n4954), .ZN(n4956) );
  AOI21_X1 U5340 ( .B1(n4957), .B2(n4956), .A(n4955), .ZN(n5299) );
  OAI22_X1 U5341 ( .A1(n5208), .A2(n4959), .B1(n4958), .B2(n5210), .ZN(n4964)
         );
  AND2_X1 U5342 ( .A1(n4961), .A2(n4960), .ZN(n5295) );
  NOR3_X1 U5343 ( .A1(n5296), .A2(n5295), .A3(n4962), .ZN(n4963) );
  AOI211_X1 U5344 ( .C1(n5328), .C2(n5299), .A(n4964), .B(n4963), .ZN(n4965)
         );
  OAI21_X1 U5345 ( .B1(n5330), .B2(n4966), .A(n4965), .ZN(U3274) );
  NOR2_X1 U5346 ( .A1(n5202), .A2(n5040), .ZN(n4967) );
  NAND2_X1 U5347 ( .A1(n3286), .A2(n4967), .ZN(n5140) );
  NAND2_X1 U5348 ( .A1(n4969), .A2(n5304), .ZN(n4973) );
  NOR2_X1 U5349 ( .A1(n4971), .A2(n4970), .ZN(n4972) );
  NAND2_X1 U5350 ( .A1(n4973), .A2(n4972), .ZN(n5020) );
  NAND4_X1 U5351 ( .A1(n4977), .A2(n4976), .A3(n4975), .A4(n4974), .ZN(n5019)
         );
  MUX2_X1 U5352 ( .A(REG1_REG_29__SCAN_IN), .B(n5020), .S(n5337), .Z(U3547) );
  MUX2_X1 U5353 ( .A(REG1_REG_28__SCAN_IN), .B(n5021), .S(n5337), .Z(U3546) );
  NAND2_X1 U5354 ( .A1(n4982), .A2(n5304), .ZN(n4984) );
  OAI211_X1 U5355 ( .C1(n5264), .C2(n4985), .A(n4984), .B(n4983), .ZN(n5022)
         );
  MUX2_X1 U5356 ( .A(REG1_REG_27__SCAN_IN), .B(n5022), .S(n5337), .Z(U3545) );
  NAND2_X1 U5357 ( .A1(n4986), .A2(n5333), .ZN(n4987) );
  OAI211_X1 U5358 ( .C1(n4989), .C2(n5140), .A(n4988), .B(n4987), .ZN(n5023)
         );
  MUX2_X1 U5359 ( .A(REG1_REG_26__SCAN_IN), .B(n5023), .S(n5337), .Z(U3544) );
  OAI211_X1 U5360 ( .C1(n4992), .C2(n5294), .A(n4991), .B(n4990), .ZN(n5024)
         );
  MUX2_X1 U5361 ( .A(REG1_REG_25__SCAN_IN), .B(n5024), .S(n5337), .Z(U3543) );
  OAI211_X1 U5362 ( .C1(n4995), .C2(n5294), .A(n4994), .B(n4993), .ZN(n5025)
         );
  MUX2_X1 U5363 ( .A(REG1_REG_24__SCAN_IN), .B(n5025), .S(n5337), .Z(U3542) );
  OAI211_X1 U5364 ( .C1(n4998), .C2(n5294), .A(n4997), .B(n4996), .ZN(n5026)
         );
  MUX2_X1 U5365 ( .A(REG1_REG_23__SCAN_IN), .B(n5026), .S(n5337), .Z(U3541) );
  NAND3_X1 U5366 ( .A1(n5000), .A2(n4999), .A3(n5304), .ZN(n5003) );
  NAND3_X1 U5367 ( .A1(n5003), .A2(n5002), .A3(n5001), .ZN(n5027) );
  MUX2_X1 U5368 ( .A(REG1_REG_22__SCAN_IN), .B(n5027), .S(n5337), .Z(U3540) );
  OAI211_X1 U5369 ( .C1(n5006), .C2(n5294), .A(n5005), .B(n5004), .ZN(n5028)
         );
  MUX2_X1 U5370 ( .A(REG1_REG_21__SCAN_IN), .B(n5028), .S(n5337), .Z(U3539) );
  OAI211_X1 U5371 ( .C1(n5009), .C2(n5294), .A(n5008), .B(n5007), .ZN(n5029)
         );
  MUX2_X1 U5372 ( .A(REG1_REG_20__SCAN_IN), .B(n5029), .S(n5337), .Z(U3538) );
  NAND3_X1 U5373 ( .A1(n5011), .A2(n5010), .A3(n5304), .ZN(n5013) );
  OAI211_X1 U5374 ( .C1(n5264), .C2(n5014), .A(n5013), .B(n5012), .ZN(n5030)
         );
  MUX2_X1 U5375 ( .A(REG1_REG_19__SCAN_IN), .B(n5030), .S(n5337), .Z(U3537) );
  OAI211_X1 U5376 ( .C1(n5017), .C2(n5294), .A(n5016), .B(n5015), .ZN(n5031)
         );
  MUX2_X1 U5377 ( .A(REG1_REG_18__SCAN_IN), .B(n5031), .S(n5337), .Z(U3536) );
  MUX2_X1 U5378 ( .A(REG0_REG_29__SCAN_IN), .B(n5020), .S(n5341), .Z(U3515) );
  MUX2_X1 U5379 ( .A(REG0_REG_28__SCAN_IN), .B(n5021), .S(n5341), .Z(U3514) );
  MUX2_X1 U5380 ( .A(REG0_REG_27__SCAN_IN), .B(n5022), .S(n5341), .Z(U3513) );
  MUX2_X1 U5381 ( .A(REG0_REG_26__SCAN_IN), .B(n5023), .S(n5341), .Z(U3512) );
  MUX2_X1 U5382 ( .A(REG0_REG_25__SCAN_IN), .B(n5024), .S(n5341), .Z(U3511) );
  MUX2_X1 U5383 ( .A(REG0_REG_24__SCAN_IN), .B(n5025), .S(n5341), .Z(U3510) );
  MUX2_X1 U5384 ( .A(REG0_REG_23__SCAN_IN), .B(n5026), .S(n5341), .Z(U3509) );
  MUX2_X1 U5385 ( .A(REG0_REG_22__SCAN_IN), .B(n5027), .S(n5341), .Z(U3508) );
  MUX2_X1 U5386 ( .A(REG0_REG_21__SCAN_IN), .B(n5028), .S(n5341), .Z(U3507) );
  MUX2_X1 U5387 ( .A(REG0_REG_20__SCAN_IN), .B(n5029), .S(n5341), .Z(U3506) );
  MUX2_X1 U5388 ( .A(REG0_REG_19__SCAN_IN), .B(n5030), .S(n5341), .Z(U3505) );
  MUX2_X1 U5389 ( .A(REG0_REG_18__SCAN_IN), .B(n5031), .S(n5341), .Z(U3503) );
  MUX2_X1 U5390 ( .A(n5032), .B(D_REG_1__SCAN_IN), .S(n5086), .Z(U3459) );
  NOR3_X1 U5391 ( .A1(n5033), .A2(IR_REG_30__SCAN_IN), .A3(n3093), .ZN(n5034)
         );
  MUX2_X1 U5392 ( .A(n5034), .B(DATAI_31_), .S(U3149), .Z(U3321) );
  MUX2_X1 U5393 ( .A(n5035), .B(DATAI_30_), .S(U3149), .Z(U3322) );
  MUX2_X1 U5394 ( .A(n5036), .B(DATAI_29_), .S(U3149), .Z(U3323) );
  MUX2_X1 U5395 ( .A(DATAI_26_), .B(n5037), .S(STATE_REG_SCAN_IN), .Z(U3326)
         );
  MUX2_X1 U5396 ( .A(n5038), .B(DATAI_25_), .S(U3149), .Z(U3327) );
  MUX2_X1 U5397 ( .A(n5039), .B(DATAI_24_), .S(U3149), .Z(U3328) );
  MUX2_X1 U5398 ( .A(n5040), .B(DATAI_22_), .S(U3149), .Z(U3330) );
  MUX2_X1 U5399 ( .A(n5041), .B(DATAI_21_), .S(U3149), .Z(U3331) );
  MUX2_X1 U5400 ( .A(DATAI_19_), .B(n5114), .S(STATE_REG_SCAN_IN), .Z(U3333)
         );
  MUX2_X1 U5401 ( .A(DATAI_18_), .B(n5042), .S(STATE_REG_SCAN_IN), .Z(U3334)
         );
  MUX2_X1 U5402 ( .A(n5043), .B(DATAI_17_), .S(U3149), .Z(U3335) );
  MUX2_X1 U5403 ( .A(n5044), .B(DATAI_16_), .S(U3149), .Z(U3336) );
  MUX2_X1 U5404 ( .A(n5045), .B(DATAI_15_), .S(U3149), .Z(U3337) );
  MUX2_X1 U5405 ( .A(n5046), .B(DATAI_14_), .S(U3149), .Z(U3338) );
  MUX2_X1 U5406 ( .A(n5047), .B(DATAI_13_), .S(U3149), .Z(U3339) );
  MUX2_X1 U5407 ( .A(DATAI_12_), .B(n5048), .S(STATE_REG_SCAN_IN), .Z(U3340)
         );
  MUX2_X1 U5408 ( .A(n5049), .B(DATAI_11_), .S(U3149), .Z(U3341) );
  MUX2_X1 U5409 ( .A(n5050), .B(DATAI_10_), .S(U3149), .Z(U3342) );
  MUX2_X1 U5410 ( .A(DATAI_9_), .B(n5051), .S(STATE_REG_SCAN_IN), .Z(U3343) );
  MUX2_X1 U5411 ( .A(DATAI_8_), .B(n5052), .S(STATE_REG_SCAN_IN), .Z(U3344) );
  MUX2_X1 U5412 ( .A(DATAI_7_), .B(n5053), .S(STATE_REG_SCAN_IN), .Z(U3345) );
  MUX2_X1 U5413 ( .A(n5054), .B(DATAI_6_), .S(U3149), .Z(U3346) );
  MUX2_X1 U5414 ( .A(n5055), .B(DATAI_5_), .S(U3149), .Z(U3347) );
  MUX2_X1 U5415 ( .A(DATAI_4_), .B(n5096), .S(STATE_REG_SCAN_IN), .Z(U3348) );
  MUX2_X1 U5416 ( .A(n5056), .B(DATAI_3_), .S(U3149), .Z(U3349) );
  MUX2_X1 U5417 ( .A(n5057), .B(DATAI_2_), .S(U3149), .Z(U3350) );
  MUX2_X1 U5418 ( .A(n3347), .B(DATAI_1_), .S(U3149), .Z(U3351) );
  MUX2_X1 U5419 ( .A(DATAI_0_), .B(IR_REG_0__SCAN_IN), .S(STATE_REG_SCAN_IN), 
        .Z(U3352) );
  INV_X1 U5420 ( .A(D_REG_2__SCAN_IN), .ZN(n5058) );
  NOR2_X1 U5421 ( .A1(n5085), .A2(n5058), .ZN(U3320) );
  AND2_X1 U5422 ( .A1(n5086), .A2(D_REG_3__SCAN_IN), .ZN(U3319) );
  NOR2_X1 U5423 ( .A1(n5085), .A2(n5059), .ZN(U3318) );
  INV_X1 U5424 ( .A(D_REG_5__SCAN_IN), .ZN(n5060) );
  NOR2_X1 U5425 ( .A1(n5085), .A2(n5060), .ZN(U3317) );
  INV_X1 U5426 ( .A(D_REG_6__SCAN_IN), .ZN(n5061) );
  NOR2_X1 U5427 ( .A1(n5085), .A2(n5061), .ZN(U3316) );
  NOR2_X1 U5428 ( .A1(n5085), .A2(n5062), .ZN(U3315) );
  INV_X1 U5429 ( .A(D_REG_8__SCAN_IN), .ZN(n5063) );
  NOR2_X1 U5430 ( .A1(n5085), .A2(n5063), .ZN(U3314) );
  NOR2_X1 U5431 ( .A1(n5085), .A2(n5064), .ZN(U3313) );
  NOR2_X1 U5432 ( .A1(n5085), .A2(n5065), .ZN(U3312) );
  NOR2_X1 U5433 ( .A1(n5085), .A2(n5066), .ZN(U3311) );
  INV_X1 U5434 ( .A(D_REG_12__SCAN_IN), .ZN(n5067) );
  NOR2_X1 U5435 ( .A1(n5085), .A2(n5067), .ZN(U3310) );
  NOR2_X1 U5436 ( .A1(n5085), .A2(n5068), .ZN(U3309) );
  NOR2_X1 U5437 ( .A1(n5085), .A2(n5069), .ZN(U3308) );
  NOR2_X1 U5438 ( .A1(n5085), .A2(n5070), .ZN(U3307) );
  NOR2_X1 U5439 ( .A1(n5085), .A2(n5071), .ZN(U3306) );
  NOR2_X1 U5440 ( .A1(n5085), .A2(n5072), .ZN(U3305) );
  NOR2_X1 U5441 ( .A1(n5085), .A2(n5073), .ZN(U3304) );
  NOR2_X1 U5442 ( .A1(n5085), .A2(n5074), .ZN(U3303) );
  INV_X1 U5443 ( .A(D_REG_20__SCAN_IN), .ZN(n5075) );
  NOR2_X1 U5444 ( .A1(n5085), .A2(n5075), .ZN(U3302) );
  INV_X1 U5445 ( .A(D_REG_21__SCAN_IN), .ZN(n5076) );
  NOR2_X1 U5446 ( .A1(n5085), .A2(n5076), .ZN(U3301) );
  NOR2_X1 U5447 ( .A1(n5085), .A2(n5077), .ZN(U3300) );
  NOR2_X1 U5448 ( .A1(n5085), .A2(n5078), .ZN(U3299) );
  INV_X1 U5449 ( .A(D_REG_24__SCAN_IN), .ZN(n5079) );
  NOR2_X1 U5450 ( .A1(n5085), .A2(n5079), .ZN(U3298) );
  AND2_X1 U5451 ( .A1(n5086), .A2(D_REG_25__SCAN_IN), .ZN(U3297) );
  NOR2_X1 U5452 ( .A1(n5085), .A2(n5080), .ZN(U3296) );
  NOR2_X1 U5453 ( .A1(n5085), .A2(n5081), .ZN(U3295) );
  NOR2_X1 U5454 ( .A1(n5085), .A2(n5082), .ZN(U3294) );
  NOR2_X1 U5455 ( .A1(n5085), .A2(n5083), .ZN(U3293) );
  INV_X1 U5456 ( .A(D_REG_30__SCAN_IN), .ZN(n5084) );
  NOR2_X1 U5457 ( .A1(n5085), .A2(n5084), .ZN(U3292) );
  AND2_X1 U5458 ( .A1(n5086), .A2(D_REG_31__SCAN_IN), .ZN(U3291) );
  AOI21_X1 U5459 ( .B1(n5088), .B2(ADDR_REG_4__SCAN_IN), .A(n5087), .ZN(n5103)
         );
  INV_X1 U5460 ( .A(n5089), .ZN(n5097) );
  AOI211_X1 U5461 ( .C1(n5093), .C2(n5092), .A(n5091), .B(n5090), .ZN(n5095)
         );
  AOI211_X1 U5462 ( .C1(n5097), .C2(n5096), .A(n5095), .B(n5094), .ZN(n5102)
         );
  OAI211_X1 U5463 ( .C1(REG1_REG_4__SCAN_IN), .C2(n5100), .A(n5099), .B(n5098), 
        .ZN(n5101) );
  NAND3_X1 U5464 ( .A1(n5103), .A2(n5102), .A3(n5101), .ZN(U3244) );
  INV_X1 U5465 ( .A(n5140), .ZN(n5225) );
  NAND2_X1 U5466 ( .A1(n5105), .A2(n5104), .ZN(n5120) );
  NOR2_X1 U5467 ( .A1(n5107), .A2(n5106), .ZN(n5117) );
  OAI21_X1 U5468 ( .B1(n5163), .B2(n5108), .A(n5120), .ZN(n5109) );
  OAI21_X1 U5469 ( .B1(n5110), .B2(n5188), .A(n5109), .ZN(n5115) );
  AOI211_X1 U5470 ( .C1(n5225), .C2(n5120), .A(n5117), .B(n5115), .ZN(n5113)
         );
  AOI22_X1 U5471 ( .A1(n5337), .A2(n5113), .B1(n5111), .B2(n5335), .ZN(U3518)
         );
  AOI22_X1 U5472 ( .A1(n5341), .A2(n5113), .B1(n5112), .B2(n5338), .ZN(U3467)
         );
  NAND2_X1 U5473 ( .A1(n3286), .A2(n5114), .ZN(n5116) );
  AOI21_X1 U5474 ( .B1(n5117), .B2(n5116), .A(n5115), .ZN(n5123) );
  INV_X1 U5475 ( .A(REG2_REG_0__SCAN_IN), .ZN(n5122) );
  AOI22_X1 U5476 ( .A1(n5120), .A2(n5119), .B1(REG3_REG_0__SCAN_IN), .B2(n5118), .ZN(n5121) );
  OAI221_X1 U5477 ( .B1(n5330), .B2(n5123), .C1(n5208), .C2(n5122), .A(n5121), 
        .ZN(U3290) );
  INV_X1 U5478 ( .A(n5124), .ZN(n5129) );
  NOR3_X1 U5479 ( .A1(n5126), .A2(n5125), .A3(n5264), .ZN(n5128) );
  AOI211_X1 U5480 ( .C1(n5129), .C2(n5225), .A(n5128), .B(n5127), .ZN(n5132)
         );
  AOI22_X1 U5481 ( .A1(n5337), .A2(n5132), .B1(n5130), .B2(n5335), .ZN(U3519)
         );
  INV_X1 U5482 ( .A(REG0_REG_1__SCAN_IN), .ZN(n5131) );
  AOI22_X1 U5483 ( .A1(n5341), .A2(n5132), .B1(n5131), .B2(n5338), .ZN(U3469)
         );
  NOR2_X1 U5484 ( .A1(n5133), .A2(n5264), .ZN(n5135) );
  AOI211_X1 U5485 ( .C1(n5225), .C2(n5136), .A(n5135), .B(n5134), .ZN(n5139)
         );
  AOI22_X1 U5486 ( .A1(n5337), .A2(n5139), .B1(n5137), .B2(n5335), .ZN(U3520)
         );
  INV_X1 U5487 ( .A(REG0_REG_2__SCAN_IN), .ZN(n5138) );
  AOI22_X1 U5488 ( .A1(n5341), .A2(n5139), .B1(n5138), .B2(n5338), .ZN(U3471)
         );
  NOR2_X1 U5489 ( .A1(n5141), .A2(n5140), .ZN(n5143) );
  AOI211_X1 U5490 ( .C1(n5333), .C2(n5144), .A(n5143), .B(n5142), .ZN(n5147)
         );
  INV_X1 U5491 ( .A(REG1_REG_3__SCAN_IN), .ZN(n5145) );
  AOI22_X1 U5492 ( .A1(n5337), .A2(n5147), .B1(n5145), .B2(n5335), .ZN(U3521)
         );
  INV_X1 U5493 ( .A(REG0_REG_3__SCAN_IN), .ZN(n5146) );
  AOI22_X1 U5494 ( .A1(n5341), .A2(n5147), .B1(n5146), .B2(n5338), .ZN(U3473)
         );
  XOR2_X1 U5495 ( .A(n5148), .B(n5153), .Z(n5170) );
  INV_X1 U5496 ( .A(n5181), .ZN(n5149) );
  OAI211_X1 U5497 ( .C1(n5151), .C2(n5150), .A(n5149), .B(n5333), .ZN(n5171)
         );
  INV_X1 U5498 ( .A(n5171), .ZN(n5165) );
  XNOR2_X1 U5499 ( .A(n5153), .B(n5152), .ZN(n5161) );
  AOI22_X1 U5500 ( .A1(n5157), .A2(n5156), .B1(n5155), .B2(n5154), .ZN(n5160)
         );
  NAND2_X1 U5501 ( .A1(n5158), .A2(n5191), .ZN(n5159) );
  OAI211_X1 U5502 ( .C1(n5161), .C2(n5194), .A(n5160), .B(n5159), .ZN(n5162)
         );
  AOI21_X1 U5503 ( .B1(n5170), .B2(n5163), .A(n5162), .ZN(n5173) );
  INV_X1 U5504 ( .A(n5173), .ZN(n5164) );
  AOI211_X1 U5505 ( .C1(n5225), .C2(n5170), .A(n5165), .B(n5164), .ZN(n5168)
         );
  INV_X1 U5506 ( .A(REG1_REG_4__SCAN_IN), .ZN(n5166) );
  AOI22_X1 U5507 ( .A1(n5337), .A2(n5168), .B1(n5166), .B2(n5335), .ZN(U3522)
         );
  INV_X1 U5508 ( .A(REG0_REG_4__SCAN_IN), .ZN(n5167) );
  AOI22_X1 U5509 ( .A1(n5341), .A2(n5168), .B1(n5167), .B2(n5338), .ZN(U3475)
         );
  NAND2_X1 U5510 ( .A1(n5170), .A2(n5169), .ZN(n5172) );
  MUX2_X1 U5511 ( .A(n5172), .B(n5171), .S(n5202), .Z(n5174) );
  NAND3_X1 U5512 ( .A1(n5174), .A2(n5173), .A3(n5208), .ZN(n5175) );
  OAI21_X1 U5513 ( .B1(REG2_REG_4__SCAN_IN), .B2(n5208), .A(n5175), .ZN(n5176)
         );
  OAI21_X1 U5514 ( .B1(n5177), .B2(n5210), .A(n5176), .ZN(U3286) );
  XNOR2_X1 U5515 ( .A(n5178), .B(n5179), .ZN(n5200) );
  OR2_X1 U5516 ( .A1(n5181), .A2(n5180), .ZN(n5182) );
  AND3_X1 U5517 ( .A1(n5183), .A2(n5182), .A3(n5333), .ZN(n5203) );
  XNOR2_X1 U5518 ( .A(n5185), .B(n5184), .ZN(n5195) );
  OAI22_X1 U5519 ( .A1(n5189), .A2(n5188), .B1(n5187), .B2(n5186), .ZN(n5190)
         );
  AOI21_X1 U5520 ( .B1(n5192), .B2(n5191), .A(n5190), .ZN(n5193) );
  OAI21_X1 U5521 ( .B1(n5195), .B2(n5194), .A(n5193), .ZN(n5201) );
  AOI211_X1 U5522 ( .C1(n5200), .C2(n5304), .A(n5203), .B(n5201), .ZN(n5198)
         );
  AOI22_X1 U5523 ( .A1(n5337), .A2(n5198), .B1(n5196), .B2(n5335), .ZN(U3523)
         );
  INV_X1 U5524 ( .A(REG0_REG_5__SCAN_IN), .ZN(n5197) );
  AOI22_X1 U5525 ( .A1(n5341), .A2(n5198), .B1(n5197), .B2(n5338), .ZN(U3477)
         );
  INV_X1 U5526 ( .A(n5199), .ZN(n5206) );
  INV_X1 U5527 ( .A(n5200), .ZN(n5205) );
  AOI211_X1 U5528 ( .C1(n5203), .C2(n5202), .A(n5330), .B(n5201), .ZN(n5204)
         );
  OAI21_X1 U5529 ( .B1(n5206), .B2(n5205), .A(n5204), .ZN(n5207) );
  OAI21_X1 U5530 ( .B1(REG2_REG_5__SCAN_IN), .B2(n5208), .A(n5207), .ZN(n5209)
         );
  OAI21_X1 U5531 ( .B1(n5211), .B2(n5210), .A(n5209), .ZN(U3285) );
  AOI211_X1 U5532 ( .C1(n5304), .C2(n5214), .A(n5213), .B(n5212), .ZN(n5216)
         );
  AOI22_X1 U5533 ( .A1(n5337), .A2(n5216), .B1(n3367), .B2(n5335), .ZN(U3524)
         );
  INV_X1 U5534 ( .A(REG0_REG_6__SCAN_IN), .ZN(n5215) );
  AOI22_X1 U5535 ( .A1(n5341), .A2(n5216), .B1(n5215), .B2(n5338), .ZN(U3479)
         );
  AOI211_X1 U5536 ( .C1(n5219), .C2(n5304), .A(n5218), .B(n5217), .ZN(n5221)
         );
  AOI22_X1 U5537 ( .A1(n5337), .A2(n5221), .B1(n3369), .B2(n5335), .ZN(U3525)
         );
  INV_X1 U5538 ( .A(REG0_REG_7__SCAN_IN), .ZN(n5220) );
  AOI22_X1 U5539 ( .A1(n5341), .A2(n5221), .B1(n5220), .B2(n5338), .ZN(U3481)
         );
  INV_X1 U5540 ( .A(n5222), .ZN(n5224) );
  AOI211_X1 U5541 ( .C1(n5225), .C2(n5224), .A(n2539), .B(n5223), .ZN(n5228)
         );
  INV_X1 U5542 ( .A(REG1_REG_8__SCAN_IN), .ZN(n5226) );
  AOI22_X1 U5543 ( .A1(n5337), .A2(n5228), .B1(n5226), .B2(n5335), .ZN(U3526)
         );
  INV_X1 U5544 ( .A(REG0_REG_8__SCAN_IN), .ZN(n5227) );
  AOI22_X1 U5545 ( .A1(n5341), .A2(n5228), .B1(n5227), .B2(n5338), .ZN(U3483)
         );
  NOR2_X1 U5546 ( .A1(n5229), .A2(n5264), .ZN(n5231) );
  AOI211_X1 U5547 ( .C1(n5232), .C2(n5304), .A(n5231), .B(n5230), .ZN(n5234)
         );
  AOI22_X1 U5548 ( .A1(n5337), .A2(n5234), .B1(n3539), .B2(n5335), .ZN(U3527)
         );
  INV_X1 U5549 ( .A(REG0_REG_9__SCAN_IN), .ZN(n5233) );
  AOI22_X1 U5550 ( .A1(n5341), .A2(n5234), .B1(n5233), .B2(n5338), .ZN(U3485)
         );
  NOR3_X1 U5551 ( .A1(n5235), .A2(n2589), .A3(n5264), .ZN(n5237) );
  AOI211_X1 U5552 ( .C1(n5238), .C2(n5304), .A(n5237), .B(n5236), .ZN(n5241)
         );
  INV_X1 U5553 ( .A(REG1_REG_10__SCAN_IN), .ZN(n5239) );
  AOI22_X1 U5554 ( .A1(n5337), .A2(n5241), .B1(n5239), .B2(n5335), .ZN(U3528)
         );
  INV_X1 U5555 ( .A(REG0_REG_10__SCAN_IN), .ZN(n5240) );
  AOI22_X1 U5556 ( .A1(n5341), .A2(n5241), .B1(n5240), .B2(n5338), .ZN(U3487)
         );
  OAI22_X1 U5557 ( .A1(n5243), .A2(n5294), .B1(n5264), .B2(n5242), .ZN(n5245)
         );
  NOR2_X1 U5558 ( .A1(n5245), .A2(n5244), .ZN(n5247) );
  AOI22_X1 U5559 ( .A1(n5337), .A2(n5247), .B1(n3661), .B2(n5335), .ZN(U3529)
         );
  INV_X1 U5560 ( .A(REG0_REG_11__SCAN_IN), .ZN(n5246) );
  AOI22_X1 U5561 ( .A1(n5341), .A2(n5247), .B1(n5246), .B2(n5338), .ZN(U3489)
         );
  AOI211_X1 U5562 ( .C1(n5250), .C2(n5304), .A(n5249), .B(n5248), .ZN(n5253)
         );
  INV_X1 U5563 ( .A(REG1_REG_12__SCAN_IN), .ZN(n5251) );
  AOI22_X1 U5564 ( .A1(n5337), .A2(n5253), .B1(n5251), .B2(n5335), .ZN(U3530)
         );
  INV_X1 U5565 ( .A(REG0_REG_12__SCAN_IN), .ZN(n5252) );
  AOI22_X1 U5566 ( .A1(n5341), .A2(n5253), .B1(n5252), .B2(n5338), .ZN(U3491)
         );
  NOR3_X1 U5567 ( .A1(n5255), .A2(n5254), .A3(n5264), .ZN(n5257) );
  AOI211_X1 U5568 ( .C1(n5258), .C2(n5304), .A(n5257), .B(n5256), .ZN(n5261)
         );
  AOI22_X1 U5569 ( .A1(n5337), .A2(n5261), .B1(n5259), .B2(n5335), .ZN(U3531)
         );
  INV_X1 U5570 ( .A(REG0_REG_13__SCAN_IN), .ZN(n5260) );
  AOI22_X1 U5571 ( .A1(n5341), .A2(n5261), .B1(n5260), .B2(n5338), .ZN(U3493)
         );
  INV_X1 U5572 ( .A(n5262), .ZN(n5263) );
  OAI22_X1 U5573 ( .A1(n5265), .A2(n5294), .B1(n5264), .B2(n5263), .ZN(n5266)
         );
  NOR2_X1 U5574 ( .A1(n5267), .A2(n5266), .ZN(n5269) );
  AOI22_X1 U5575 ( .A1(n5337), .A2(n5269), .B1(n4633), .B2(n5335), .ZN(U3532)
         );
  INV_X1 U5576 ( .A(REG0_REG_14__SCAN_IN), .ZN(n5268) );
  AOI22_X1 U5577 ( .A1(n5341), .A2(n5269), .B1(n5268), .B2(n5338), .ZN(U3495)
         );
  OAI22_X1 U5578 ( .A1(n5273), .A2(n5272), .B1(n5271), .B2(n5270), .ZN(n5274)
         );
  AOI211_X1 U5579 ( .C1(n5277), .C2(n5276), .A(n5275), .B(n5274), .ZN(n5285)
         );
  NAND2_X1 U5580 ( .A1(n5279), .A2(n5278), .ZN(n5281) );
  XNOR2_X1 U5581 ( .A(n5281), .B(n5280), .ZN(n5283) );
  NAND2_X1 U5582 ( .A1(n5283), .A2(n5282), .ZN(n5284) );
  OAI211_X1 U5583 ( .C1(n5287), .C2(n5286), .A(n5285), .B(n5284), .ZN(U3238)
         );
  AOI211_X1 U5584 ( .C1(n5290), .C2(n5304), .A(n5289), .B(n5288), .ZN(n5293)
         );
  AOI22_X1 U5585 ( .A1(n5337), .A2(n5293), .B1(n5291), .B2(n5335), .ZN(U3533)
         );
  INV_X1 U5586 ( .A(REG0_REG_15__SCAN_IN), .ZN(n5292) );
  AOI22_X1 U5587 ( .A1(n5341), .A2(n5293), .B1(n5292), .B2(n5338), .ZN(U3497)
         );
  NOR3_X1 U5588 ( .A1(n5296), .A2(n5295), .A3(n5294), .ZN(n5297) );
  AOI211_X1 U5589 ( .C1(n5333), .C2(n5299), .A(n5298), .B(n5297), .ZN(n5301)
         );
  AOI22_X1 U5590 ( .A1(n5337), .A2(n5301), .B1(n2721), .B2(n5335), .ZN(U3534)
         );
  INV_X1 U5591 ( .A(REG0_REG_16__SCAN_IN), .ZN(n5300) );
  AOI22_X1 U5592 ( .A1(n5341), .A2(n5301), .B1(n5300), .B2(n5338), .ZN(U3499)
         );
  AOI211_X1 U5593 ( .C1(n5305), .C2(n5304), .A(n5303), .B(n5302), .ZN(n5308)
         );
  AOI22_X1 U5594 ( .A1(n5337), .A2(n5308), .B1(n5306), .B2(n5335), .ZN(U3535)
         );
  INV_X1 U5595 ( .A(REG0_REG_17__SCAN_IN), .ZN(n5307) );
  AOI22_X1 U5596 ( .A1(n5341), .A2(n5308), .B1(n5307), .B2(n5338), .ZN(U3501)
         );
  NAND2_X1 U5597 ( .A1(n5310), .A2(n5309), .ZN(n5322) );
  OR2_X1 U5598 ( .A1(n5323), .A2(n5319), .ZN(n5311) );
  AND2_X1 U5599 ( .A1(n5322), .A2(n5311), .ZN(n5313) );
  XNOR2_X1 U5600 ( .A(n5325), .B(n5323), .ZN(n5315) );
  AOI22_X1 U5601 ( .A1(n5315), .A2(n5328), .B1(REG2_REG_30__SCAN_IN), .B2(
        n5330), .ZN(n5312) );
  OAI21_X1 U5602 ( .B1(n5330), .B2(n5313), .A(n5312), .ZN(U3261) );
  INV_X1 U5603 ( .A(n5313), .ZN(n5314) );
  AOI21_X1 U5604 ( .B1(n5315), .B2(n5333), .A(n5314), .ZN(n5318) );
  INV_X1 U5605 ( .A(REG1_REG_30__SCAN_IN), .ZN(n5316) );
  AOI22_X1 U5606 ( .A1(n5337), .A2(n5318), .B1(n5316), .B2(n5335), .ZN(U3548)
         );
  INV_X1 U5607 ( .A(REG0_REG_30__SCAN_IN), .ZN(n5317) );
  AOI22_X1 U5608 ( .A1(n5341), .A2(n5318), .B1(n5317), .B2(n5338), .ZN(U3516)
         );
  OR2_X1 U5609 ( .A1(n5320), .A2(n5319), .ZN(n5321) );
  AND2_X1 U5610 ( .A1(n5322), .A2(n5321), .ZN(n5331) );
  INV_X1 U5611 ( .A(n5323), .ZN(n5324) );
  NOR2_X1 U5612 ( .A1(n5325), .A2(n5324), .ZN(n5327) );
  XNOR2_X1 U5613 ( .A(n5327), .B(n5326), .ZN(n5334) );
  AOI22_X1 U5614 ( .A1(n5334), .A2(n5328), .B1(n5330), .B2(
        REG2_REG_31__SCAN_IN), .ZN(n5329) );
  OAI21_X1 U5615 ( .B1(n5330), .B2(n5331), .A(n5329), .ZN(U3260) );
  INV_X1 U5616 ( .A(n5331), .ZN(n5332) );
  AOI21_X1 U5617 ( .B1(n5334), .B2(n5333), .A(n5332), .ZN(n5340) );
  INV_X1 U5618 ( .A(REG1_REG_31__SCAN_IN), .ZN(n5336) );
  AOI22_X1 U5619 ( .A1(n5337), .A2(n5340), .B1(n5336), .B2(n5335), .ZN(U3549)
         );
  INV_X1 U5620 ( .A(REG0_REG_31__SCAN_IN), .ZN(n5339) );
  AOI22_X1 U5621 ( .A1(n5341), .A2(n5340), .B1(n5339), .B2(n5338), .ZN(U3517)
         );
  INV_X2 U2542 ( .A(n3464), .ZN(n3252) );
endmodule

