

module b15_C_AntiSAT_k_128_8 ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1, 
        keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7, 
        keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13, 
        keyinput14, keyinput15, keyinput16, keyinput17, keyinput18, keyinput19, 
        keyinput20, keyinput21, keyinput22, keyinput23, keyinput24, keyinput25, 
        keyinput26, keyinput27, keyinput28, keyinput29, keyinput30, keyinput31, 
        keyinput32, keyinput33, keyinput34, keyinput35, keyinput36, keyinput37, 
        keyinput38, keyinput39, keyinput40, keyinput41, keyinput42, keyinput43, 
        keyinput44, keyinput45, keyinput46, keyinput47, keyinput48, keyinput49, 
        keyinput50, keyinput51, keyinput52, keyinput53, keyinput54, keyinput55, 
        keyinput56, keyinput57, keyinput58, keyinput59, keyinput60, keyinput61, 
        keyinput62, keyinput63, keyinput64, keyinput65, keyinput66, keyinput67, 
        keyinput68, keyinput69, keyinput70, keyinput71, keyinput72, keyinput73, 
        keyinput74, keyinput75, keyinput76, keyinput77, keyinput78, keyinput79, 
        keyinput80, keyinput81, keyinput82, keyinput83, keyinput84, keyinput85, 
        keyinput86, keyinput87, keyinput88, keyinput89, keyinput90, keyinput91, 
        keyinput92, keyinput93, keyinput94, keyinput95, keyinput96, keyinput97, 
        keyinput98, keyinput99, keyinput100, keyinput101, keyinput102, 
        keyinput103, keyinput104, keyinput105, keyinput106, keyinput107, 
        keyinput108, keyinput109, keyinput110, keyinput111, keyinput112, 
        keyinput113, keyinput114, keyinput115, keyinput116, keyinput117, 
        keyinput118, keyinput119, keyinput120, keyinput121, keyinput122, 
        keyinput123, keyinput124, keyinput125, keyinput126, keyinput127, U3445, 
        U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208, U3207, 
        U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198, U3197, 
        U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188, U3187, 
        U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180, U3179, 
        U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170, U3169, 
        U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160, U3159, 
        U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453, U3150, 
        U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141, U3140, 
        U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131, U3130, 
        U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121, U3120, 
        U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111, U3110, 
        U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101, U3100, 
        U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091, U3090, 
        U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081, U3080, 
        U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071, U3070, 
        U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061, U3060, 
        U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051, U3050, 
        U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041, U3040, 
        U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031, U3030, 
        U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021, U3020, 
        U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464, U3465, 
        U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010, U3009, 
        U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000, U2999, 
        U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990, U2989, 
        U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980, U2979, 
        U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970, U2969, 
        U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960, U2959, 
        U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950, U2949, 
        U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940, U2939, 
        U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930, U2929, 
        U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920, U2919, 
        U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910, U2909, 
        U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900, U2899, 
        U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890, U2889, 
        U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880, U2879, 
        U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870, U2869, 
        U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860, U2859, 
        U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850, U2849, 
        U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840, U2839, 
        U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830, U2829, 
        U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820, U2819, 
        U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810, U2809, 
        U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800, U2799, 
        U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793, U3471, 
        U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput0, keyinput1,
         keyinput2, keyinput3, keyinput4, keyinput5, keyinput6, keyinput7,
         keyinput8, keyinput9, keyinput10, keyinput11, keyinput12, keyinput13,
         keyinput14, keyinput15, keyinput16, keyinput17, keyinput18,
         keyinput19, keyinput20, keyinput21, keyinput22, keyinput23,
         keyinput24, keyinput25, keyinput26, keyinput27, keyinput28,
         keyinput29, keyinput30, keyinput31, keyinput32, keyinput33,
         keyinput34, keyinput35, keyinput36, keyinput37, keyinput38,
         keyinput39, keyinput40, keyinput41, keyinput42, keyinput43,
         keyinput44, keyinput45, keyinput46, keyinput47, keyinput48,
         keyinput49, keyinput50, keyinput51, keyinput52, keyinput53,
         keyinput54, keyinput55, keyinput56, keyinput57, keyinput58,
         keyinput59, keyinput60, keyinput61, keyinput62, keyinput63,
         keyinput64, keyinput65, keyinput66, keyinput67, keyinput68,
         keyinput69, keyinput70, keyinput71, keyinput72, keyinput73,
         keyinput74, keyinput75, keyinput76, keyinput77, keyinput78,
         keyinput79, keyinput80, keyinput81, keyinput82, keyinput83,
         keyinput84, keyinput85, keyinput86, keyinput87, keyinput88,
         keyinput89, keyinput90, keyinput91, keyinput92, keyinput93,
         keyinput94, keyinput95, keyinput96, keyinput97, keyinput98,
         keyinput99, keyinput100, keyinput101, keyinput102, keyinput103,
         keyinput104, keyinput105, keyinput106, keyinput107, keyinput108,
         keyinput109, keyinput110, keyinput111, keyinput112, keyinput113,
         keyinput114, keyinput115, keyinput116, keyinput117, keyinput118,
         keyinput119, keyinput120, keyinput121, keyinput122, keyinput123,
         keyinput124, keyinput125, keyinput126, keyinput127;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784;

  AND2_X1 U34470 ( .A1(n3259), .A2(n3271), .ZN(n5420) );
  CLKBUF_X2 U34480 ( .A(n3253), .Z(n3029) );
  BUF_X2 U3449 ( .A(n3204), .Z(n4258) );
  CLKBUF_X2 U3450 ( .A(n3393), .Z(n4239) );
  CLKBUF_X2 U34510 ( .A(n3399), .Z(n3033) );
  AND2_X2 U34520 ( .A1(n3291), .A2(n3290), .ZN(n6437) );
  CLKBUF_X2 U34530 ( .A(n3189), .Z(n4259) );
  CLKBUF_X2 U3454 ( .A(n3349), .Z(n4155) );
  CLKBUF_X2 U34550 ( .A(n3213), .Z(n4177) );
  CLKBUF_X2 U34560 ( .A(n3392), .Z(n4097) );
  AND2_X1 U3458 ( .A1(n3086), .A2(n4530), .ZN(n4149) );
  AND2_X2 U34590 ( .A1(n4367), .A2(n4530), .ZN(n3189) );
  AND2_X2 U34600 ( .A1(n4533), .A2(n3085), .ZN(n3036) );
  NOR2_X2 U34610 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4539) );
  INV_X1 U34630 ( .A(n3259), .ZN(n3635) );
  AND2_X2 U34640 ( .A1(n3055), .A2(n3054), .ZN(n4358) );
  INV_X1 U34650 ( .A(n3271), .ZN(n3348) );
  XNOR2_X2 U3466 ( .A(n3490), .B(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4498)
         );
  NOR2_X4 U3467 ( .A1(n5084), .A2(n3891), .ZN(n5083) );
  NOR2_X4 U34680 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3085) );
  NAND2_X1 U34700 ( .A1(n3777), .A2(n3037), .ZN(n5607) );
  INV_X4 U34710 ( .A(n5864), .ZN(n2999) );
  NAND2_X1 U34720 ( .A1(n4950), .A2(n4949), .ZN(n5529) );
  INV_X2 U34730 ( .A(n3273), .ZN(n4374) );
  BUF_X1 U34740 ( .A(n3032), .Z(n3026) );
  CLKBUF_X2 U3475 ( .A(n3398), .Z(n4233) );
  AND2_X1 U3476 ( .A1(n4539), .A2(n4324), .ZN(n3213) );
  INV_X1 U3477 ( .A(n3102), .ZN(n5620) );
  INV_X1 U3478 ( .A(n5607), .ZN(n5608) );
  OR2_X1 U3479 ( .A1(n3554), .A2(n3010), .ZN(n3557) );
  NOR2_X1 U3480 ( .A1(n3102), .A2(n3101), .ZN(n5475) );
  AOI211_X1 U3481 ( .C1(EBX_REG_27__SCAN_IN), .C2(n6042), .A(n5761), .B(n5760), 
        .ZN(n5763) );
  AOI211_X1 U3482 ( .C1(n5814), .C2(n6347), .A(n5441), .B(n5440), .ZN(n5442)
         );
  NAND2_X1 U3483 ( .A1(n5842), .A2(n5841), .ZN(n3777) );
  NAND2_X1 U3484 ( .A1(n3040), .A2(n5568), .ZN(n5759) );
  NAND2_X1 U3485 ( .A1(n5572), .A2(n3081), .ZN(n5560) );
  CLKBUF_X1 U3486 ( .A(n5854), .Z(n5855) );
  AOI21_X1 U3487 ( .B1(n5362), .B2(n5361), .A(n5360), .ZN(n6062) );
  NAND2_X1 U3488 ( .A1(n5197), .A2(n5273), .ZN(n5272) );
  NAND2_X1 U3489 ( .A1(n3515), .A2(n3514), .ZN(n4615) );
  OR2_X1 U3490 ( .A1(n3018), .A2(n4886), .ZN(n3017) );
  NOR2_X1 U3491 ( .A1(n3099), .A2(n3100), .ZN(n3096) );
  OR2_X1 U3492 ( .A1(n5313), .A2(n5316), .ZN(n5320) );
  INV_X1 U3493 ( .A(n4397), .ZN(n3822) );
  OR2_X1 U3494 ( .A1(n3043), .A2(n5061), .ZN(n3099) );
  NAND2_X1 U3495 ( .A1(n5638), .A2(n3556), .ZN(n3010) );
  NOR2_X1 U3496 ( .A1(n4459), .A2(n4399), .ZN(n3079) );
  AND2_X1 U3497 ( .A1(n5944), .A2(n5328), .ZN(n5523) );
  OR2_X1 U3498 ( .A1(n3517), .A2(n3448), .ZN(n3038) );
  AND2_X1 U3499 ( .A1(n4392), .A2(n3478), .ZN(n6138) );
  AND2_X1 U3500 ( .A1(n3484), .A2(n3493), .ZN(n3803) );
  NOR2_X1 U3501 ( .A1(n6342), .A2(n5163), .ZN(n4956) );
  NAND2_X1 U3502 ( .A1(n3329), .A2(n3328), .ZN(n4553) );
  NAND2_X1 U3503 ( .A1(n3409), .A2(n3408), .ZN(n3481) );
  NAND2_X1 U3504 ( .A1(n4478), .A2(n3794), .ZN(n4380) );
  OR2_X1 U3505 ( .A1(n6566), .A2(n4945), .ZN(n5281) );
  NAND2_X2 U3506 ( .A1(n6053), .A2(n3275), .ZN(n5589) );
  OR2_X1 U3507 ( .A1(n4476), .A2(n4475), .ZN(n4478) );
  NOR2_X1 U3508 ( .A1(n4876), .A2(n4875), .ZN(n4935) );
  NAND2_X1 U3509 ( .A1(n3378), .A2(n3076), .ZN(n3465) );
  NAND2_X2 U3510 ( .A1(n3614), .A2(n3613), .ZN(n5520) );
  NAND2_X1 U3511 ( .A1(n3789), .A2(n6596), .ZN(n3076) );
  AOI21_X1 U3512 ( .B1(n3310), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3307), 
        .ZN(n3389) );
  AND2_X1 U3513 ( .A1(n3377), .A2(n3376), .ZN(n3378) );
  OR2_X1 U3514 ( .A1(n3374), .A2(n3458), .ZN(n3377) );
  AOI21_X1 U3515 ( .B1(n3573), .B2(n3572), .A(n3571), .ZN(n3575) );
  AND3_X1 U3516 ( .A1(n3285), .A2(n3104), .A3(n3284), .ZN(n3286) );
  AND3_X1 U3517 ( .A1(n3264), .A2(n3618), .A3(n3619), .ZN(n3265) );
  AND2_X1 U3518 ( .A1(n3656), .A2(n3655), .ZN(n4508) );
  AND2_X1 U3519 ( .A1(n3263), .A2(n3471), .ZN(n3619) );
  NAND2_X1 U3520 ( .A1(n5415), .A2(n5486), .ZN(n5427) );
  OAI211_X1 U3521 ( .C1(n3599), .C2(n4719), .A(n3371), .B(n3449), .ZN(n3460)
         );
  NAND2_X2 U3522 ( .A1(n3646), .A2(n3271), .ZN(n5415) );
  NAND2_X1 U3523 ( .A1(n3567), .A2(n3566), .ZN(n3610) );
  NAND2_X1 U3524 ( .A1(n3348), .A2(n3259), .ZN(n4952) );
  AND2_X2 U3525 ( .A1(n3635), .A2(n3271), .ZN(n6436) );
  OR2_X1 U3526 ( .A1(n3370), .A2(n3369), .ZN(n3534) );
  NAND2_X1 U3527 ( .A1(n3274), .A2(n3259), .ZN(n5423) );
  OR2_X2 U3528 ( .A1(n3315), .A2(n6596), .ZN(n3599) );
  OR2_X2 U3529 ( .A1(n3188), .A2(n3187), .ZN(n3274) );
  NOR2_X2 U3530 ( .A1(n3271), .A2(n3259), .ZN(n5519) );
  OR2_X1 U3531 ( .A1(n3360), .A2(n3359), .ZN(n3470) );
  NAND2_X2 U3532 ( .A1(n3175), .A2(n3174), .ZN(n3203) );
  NAND4_X2 U3533 ( .A1(n3134), .A2(n3133), .A3(n3132), .A4(n3131), .ZN(n3273)
         );
  AND4_X1 U3534 ( .A1(n3168), .A2(n3167), .A3(n3166), .A4(n3165), .ZN(n3175)
         );
  AND4_X1 U3535 ( .A1(n3212), .A2(n3211), .A3(n3210), .A4(n3209), .ZN(n3224)
         );
  AND4_X1 U3536 ( .A1(n3217), .A2(n3216), .A3(n3215), .A4(n3214), .ZN(n3223)
         );
  AND4_X1 U3537 ( .A1(n3208), .A2(n3207), .A3(n3206), .A4(n3205), .ZN(n3225)
         );
  AND4_X1 U3538 ( .A1(n3142), .A2(n3141), .A3(n3140), .A4(n3139), .ZN(n3143)
         );
  AND4_X1 U3539 ( .A1(n3242), .A2(n3241), .A3(n3240), .A4(n3239), .ZN(n3243)
         );
  AND4_X1 U3540 ( .A1(n3237), .A2(n3236), .A3(n3235), .A4(n3234), .ZN(n3244)
         );
  AND4_X1 U3541 ( .A1(n3233), .A2(n3232), .A3(n3231), .A4(n3230), .ZN(n3245)
         );
  AND4_X1 U3542 ( .A1(n3229), .A2(n3228), .A3(n3227), .A4(n3226), .ZN(n3246)
         );
  AND4_X1 U3543 ( .A1(n3221), .A2(n3220), .A3(n3219), .A4(n3218), .ZN(n3222)
         );
  AND4_X1 U3544 ( .A1(n3116), .A2(n3115), .A3(n3114), .A4(n3113), .ZN(n3134)
         );
  AND4_X1 U3545 ( .A1(n3173), .A2(n3172), .A3(n3171), .A4(n3170), .ZN(n3174)
         );
  AND4_X1 U3546 ( .A1(n3120), .A2(n3119), .A3(n3118), .A4(n3117), .ZN(n3133)
         );
  AND4_X1 U3547 ( .A1(n3124), .A2(n3123), .A3(n3122), .A4(n3121), .ZN(n3132)
         );
  AND4_X1 U3548 ( .A1(n3130), .A2(n3129), .A3(n3128), .A4(n3127), .ZN(n3131)
         );
  CLKBUF_X3 U3549 ( .A(n4149), .Z(n4085) );
  BUF_X2 U3550 ( .A(n3182), .Z(n4264) );
  BUF_X2 U3551 ( .A(n3238), .Z(n3000) );
  AND2_X2 U3552 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4324) );
  INV_X1 U3553 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3055) );
  INV_X1 U3554 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3021) );
  NOR2_X2 U3555 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6354) );
  CLKBUF_X1 U3556 ( .A(n4484), .Z(n3001) );
  NAND2_X2 U3557 ( .A1(n4296), .A2(n3045), .ZN(n5213) );
  AND2_X1 U3558 ( .A1(n5560), .A2(n5559), .ZN(n5817) );
  NAND2_X2 U3559 ( .A1(n3802), .A2(n3801), .ZN(n4479) );
  NAND2_X1 U3560 ( .A1(n5213), .A2(n3005), .ZN(n3002) );
  AND2_X2 U3561 ( .A1(n3002), .A2(n3003), .ZN(n3549) );
  OR2_X1 U3562 ( .A1(n3004), .A2(n3046), .ZN(n3003) );
  INV_X1 U3563 ( .A(n3088), .ZN(n3004) );
  AND2_X1 U3564 ( .A1(n3545), .A2(n3088), .ZN(n3005) );
  INV_X1 U3565 ( .A(n3252), .ZN(n3293) );
  NAND2_X1 U3566 ( .A1(n5610), .A2(n5864), .ZN(n3006) );
  NAND2_X1 U3567 ( .A1(n5609), .A2(n2999), .ZN(n3007) );
  NAND2_X1 U3568 ( .A1(n3006), .A2(n3007), .ZN(n5613) );
  NOR2_X1 U3569 ( .A1(n5613), .A2(n5612), .ZN(n5614) );
  OR2_X2 U3570 ( .A1(n5847), .A2(n3009), .ZN(n5605) );
  XNOR2_X1 U3571 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .B(n3008), .ZN(n5463)
         );
  NAND2_X1 U3572 ( .A1(n5445), .A2(n3109), .ZN(n3008) );
  AND2_X1 U3573 ( .A1(n5864), .A2(n3773), .ZN(n3009) );
  AND2_X2 U3574 ( .A1(n3126), .A2(n4367), .ZN(n4154) );
  AND2_X4 U3575 ( .A1(n4339), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3126)
         );
  NAND3_X1 U3576 ( .A1(n4553), .A2(n3482), .A3(n3481), .ZN(n3493) );
  XNOR2_X1 U3577 ( .A(n3038), .B(n3525), .ZN(n3842) );
  NAND2_X4 U3578 ( .A1(n3144), .A2(n3143), .ZN(n4451) );
  XNOR2_X2 U3579 ( .A(n3347), .B(n3346), .ZN(n3789) );
  NAND2_X2 U3580 ( .A1(n3347), .A2(n3288), .ZN(n3331) );
  OAI21_X2 U3581 ( .B1(n3304), .B2(n3021), .A(n3268), .ZN(n3347) );
  NAND2_X2 U3582 ( .A1(n3309), .A2(n3308), .ZN(n4522) );
  NAND2_X1 U3583 ( .A1(n3012), .A2(n3785), .ZN(n3011) );
  NAND2_X1 U3584 ( .A1(n3035), .A2(n3983), .ZN(n3012) );
  BUF_X1 U3585 ( .A(n5197), .Z(n3013) );
  CLKBUF_X1 U3586 ( .A(n5199), .Z(n3014) );
  NAND2_X1 U3587 ( .A1(n3786), .A2(n3785), .ZN(n4381) );
  OR2_X1 U3588 ( .A1(n5438), .A2(n5498), .ZN(n5743) );
  OR2_X1 U3589 ( .A1(n5182), .A2(n3942), .ZN(n5273) );
  NOR2_X4 U3590 ( .A1(n5309), .A2(n5319), .ZN(n5648) );
  OAI21_X2 U3591 ( .B1(n5539), .B2(n6004), .A(n3065), .ZN(n3064) );
  NAND2_X2 U3592 ( .A1(n4044), .A2(n4043), .ZN(n5309) );
  NAND2_X1 U3593 ( .A1(n4928), .A2(n4929), .ZN(n3015) );
  NAND2_X1 U3594 ( .A1(n3523), .A2(n3019), .ZN(n3016) );
  AND2_X2 U3595 ( .A1(n3016), .A2(n3017), .ZN(n4928) );
  INV_X1 U3596 ( .A(n3533), .ZN(n3018) );
  AND2_X1 U3597 ( .A1(n3522), .A2(n3533), .ZN(n3019) );
  INV_X1 U3598 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3020) );
  NAND2_X1 U3599 ( .A1(n3266), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3022) );
  NAND2_X1 U3600 ( .A1(n4928), .A2(n4929), .ZN(n3540) );
  NAND2_X1 U3601 ( .A1(n3176), .A2(n4374), .ZN(n3270) );
  AND2_X1 U3602 ( .A1(n4539), .A2(n4324), .ZN(n3023) );
  AND4_X2 U3603 ( .A1(n3160), .A2(n3159), .A3(n3158), .A4(n3157), .ZN(n3161)
         );
  AND2_X1 U3604 ( .A1(n4358), .A2(n4530), .ZN(n3024) );
  AND2_X1 U3605 ( .A1(n4358), .A2(n4530), .ZN(n3025) );
  AND2_X1 U3606 ( .A1(n4358), .A2(n4530), .ZN(n3399) );
  NAND2_X1 U3607 ( .A1(n3475), .A2(n3474), .ZN(n4393) );
  BUF_X2 U3608 ( .A(n3252), .Z(n3176) );
  AND2_X1 U3609 ( .A1(n3125), .A2(n4358), .ZN(n3032) );
  NOR2_X2 U3610 ( .A1(n5443), .A2(n3051), .ZN(n5651) );
  NOR2_X2 U3611 ( .A1(n4871), .A2(n4977), .ZN(n4976) );
  NOR2_X2 U3612 ( .A1(n3549), .A2(n3039), .ZN(n5854) );
  AND2_X1 U3613 ( .A1(n3086), .A2(n4530), .ZN(n3027) );
  AND2_X1 U3614 ( .A1(n3086), .A2(n4530), .ZN(n3028) );
  XNOR2_X2 U3615 ( .A(n3332), .B(n3331), .ZN(n4357) );
  AND2_X2 U3616 ( .A1(n4324), .A2(n4530), .ZN(n3393) );
  AND3_X1 U3617 ( .A1(n3282), .A2(n4374), .A3(n4372), .ZN(n3250) );
  AND2_X4 U3618 ( .A1(n3126), .A2(n3086), .ZN(n3182) );
  NAND2_X2 U3619 ( .A1(n3176), .A2(n3248), .ZN(n3260) );
  INV_X1 U3620 ( .A(n5423), .ZN(n3253) );
  AOI21_X1 U3621 ( .B1(n3270), .B2(n3754), .A(n3272), .ZN(n3742) );
  NAND2_X2 U3622 ( .A1(n3251), .A2(n3250), .ZN(n3292) );
  NOR2_X2 U3623 ( .A1(n5455), .A2(n5542), .ZN(n5540) );
  OAI21_X2 U3624 ( .B1(n5175), .B2(n5176), .A(n3541), .ZN(n4298) );
  BUF_X1 U3625 ( .A(n3269), .Z(n3745) );
  OAI21_X2 U3626 ( .B1(n4499), .B2(n4498), .A(n3491), .ZN(n4516) );
  NAND4_X4 U3627 ( .A1(n3164), .A2(n3163), .A3(n3162), .A4(n3161), .ZN(n3252)
         );
  AND2_X1 U3628 ( .A1(n3126), .A2(n4367), .ZN(n3030) );
  AND2_X2 U3629 ( .A1(n3126), .A2(n4367), .ZN(n3031) );
  XNOR2_X2 U3630 ( .A(n4522), .B(n6253), .ZN(n4531) );
  BUF_X1 U3631 ( .A(n4404), .Z(n3034) );
  BUF_X4 U3632 ( .A(n4404), .Z(n3035) );
  XNOR2_X1 U3633 ( .A(n3467), .B(n3466), .ZN(n4404) );
  NAND2_X1 U3634 ( .A1(n3254), .A2(n3253), .ZN(n3281) );
  OAI211_X1 U3635 ( .C1(n3247), .C2(n3203), .A(n5519), .B(n3292), .ZN(n3269)
         );
  INV_X1 U3636 ( .A(n3464), .ZN(n3386) );
  OR2_X1 U3637 ( .A1(n3756), .A2(n5510), .ZN(n4300) );
  OR2_X1 U3638 ( .A1(n2999), .A2(n3692), .ZN(n3542) );
  OR2_X1 U3639 ( .A1(n4507), .A2(n3662), .ZN(n3061) );
  OR2_X1 U3640 ( .A1(n3756), .A2(n4532), .ZN(n5219) );
  AND2_X1 U3641 ( .A1(n3560), .A2(n3252), .ZN(n3573) );
  OR2_X1 U3642 ( .A1(n3565), .A2(n5519), .ZN(n3580) );
  INV_X1 U3643 ( .A(n5225), .ZN(n3091) );
  NAND2_X1 U3644 ( .A1(n3048), .A2(n3283), .ZN(n3284) );
  NAND2_X1 U3645 ( .A1(n5648), .A2(n3049), .ZN(n5455) );
  INV_X1 U3646 ( .A(n5456), .ZN(n4127) );
  AND2_X1 U3647 ( .A1(n3037), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n3103)
         );
  NOR2_X1 U3648 ( .A1(n3052), .A2(n3091), .ZN(n3089) );
  INV_X1 U3649 ( .A(n3539), .ZN(n3100) );
  AND2_X1 U3650 ( .A1(n3259), .A2(n3252), .ZN(n3566) );
  NAND2_X1 U3651 ( .A1(n3266), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3304) );
  INV_X1 U3652 ( .A(n3599), .ZN(n3567) );
  OR2_X1 U3653 ( .A1(n3342), .A2(n3341), .ZN(n3469) );
  NAND2_X1 U3654 ( .A1(n3388), .A2(n3387), .ZN(n3482) );
  NAND2_X1 U3655 ( .A1(n3465), .A2(n3386), .ZN(n3387) );
  OR2_X1 U3656 ( .A1(n3465), .A2(n3386), .ZN(n3384) );
  NAND2_X1 U3657 ( .A1(n4340), .A2(n6596), .ZN(n3409) );
  AND2_X2 U3658 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4530) );
  NAND2_X1 U3659 ( .A1(n3258), .A2(n4372), .ZN(n3289) );
  AND2_X1 U3660 ( .A1(n4374), .A2(n3275), .ZN(n3258) );
  AND2_X1 U3661 ( .A1(n3637), .A2(n3274), .ZN(n3471) );
  INV_X1 U3662 ( .A(n5529), .ZN(n5525) );
  INV_X1 U3663 ( .A(n3837), .ZN(n3838) );
  INV_X1 U3664 ( .A(n5281), .ZN(n5163) );
  INV_X1 U3665 ( .A(n5420), .ZN(n5426) );
  AND2_X1 U3666 ( .A1(n6342), .A2(STATEBS16_REG_SCAN_IN), .ZN(n4282) );
  AND2_X1 U3667 ( .A1(n3082), .A2(n4230), .ZN(n3081) );
  INV_X1 U3668 ( .A(n5558), .ZN(n4230) );
  AND2_X1 U3669 ( .A1(n4023), .A2(n5379), .ZN(n4024) );
  INV_X1 U3670 ( .A(n3805), .ZN(n3806) );
  NAND2_X1 U3671 ( .A1(n3806), .A2(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3816)
         );
  NOR2_X1 U3672 ( .A1(n5483), .A2(n3029), .ZN(n5489) );
  INV_X1 U3673 ( .A(n5227), .ZN(n3092) );
  OR2_X1 U3674 ( .A1(n2999), .A2(n3546), .ZN(n5225) );
  INV_X1 U3675 ( .A(n5216), .ZN(n3543) );
  OR2_X1 U3676 ( .A1(n2999), .A2(n6770), .ZN(n3541) );
  NAND2_X1 U3677 ( .A1(n4298), .A2(n4297), .ZN(n4296) );
  INV_X1 U3678 ( .A(n4300), .ZN(n6171) );
  OR2_X1 U3679 ( .A1(n3653), .A2(n3652), .ZN(n3654) );
  AND2_X1 U3680 ( .A1(n5219), .A2(n5229), .ZN(n4931) );
  AND2_X1 U3681 ( .A1(n3641), .A2(n3640), .ZN(n3756) );
  NAND2_X1 U3682 ( .A1(n3609), .A2(n3608), .ZN(n3614) );
  NOR2_X1 U3683 ( .A1(n5535), .A2(n3044), .ZN(n3065) );
  NOR2_X1 U3684 ( .A1(n3575), .A2(n3574), .ZN(n3589) );
  INV_X1 U3685 ( .A(n3580), .ZN(n3588) );
  NAND2_X1 U3686 ( .A1(n3422), .A2(n3047), .ZN(n3517) );
  OR2_X1 U3687 ( .A1(n3420), .A2(n3419), .ZN(n3494) );
  NAND2_X1 U3688 ( .A1(n3273), .A2(n3271), .ZN(n3315) );
  NOR2_X1 U3689 ( .A1(n3259), .A2(n3623), .ZN(n3295) );
  NAND2_X1 U3690 ( .A1(n3261), .A2(n3289), .ZN(n3618) );
  AND2_X1 U3691 ( .A1(n3260), .A2(n3271), .ZN(n3261) );
  OR2_X1 U3692 ( .A1(n3604), .A2(n3605), .ZN(n3629) );
  NAND2_X1 U3693 ( .A1(n3315), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3607) );
  NOR2_X1 U3694 ( .A1(n3274), .A2(n3203), .ZN(n4373) );
  NOR2_X1 U3695 ( .A1(n3083), .A2(n5567), .ZN(n3082) );
  INV_X1 U3696 ( .A(n5573), .ZN(n3083) );
  AND2_X1 U3697 ( .A1(n5396), .A2(n5647), .ZN(n3077) );
  INV_X1 U3698 ( .A(n4873), .ZN(n3843) );
  NAND2_X1 U3699 ( .A1(n5420), .A2(n5486), .ZN(n5411) );
  NAND2_X1 U3700 ( .A1(n4374), .A2(n3534), .ZN(n3449) );
  AND3_X2 U3701 ( .A1(n3745), .A2(n3287), .A3(n3286), .ZN(n3346) );
  AND2_X1 U3702 ( .A1(n3742), .A2(n3278), .ZN(n3287) );
  INV_X1 U3703 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3054) );
  NAND2_X1 U3704 ( .A1(n3314), .A2(n3313), .ZN(n6253) );
  INV_X1 U3705 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6415) );
  AOI22_X1 U3706 ( .A1(n4154), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3023), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3171) );
  AOI22_X1 U3707 ( .A1(n3177), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3238), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3168) );
  AOI22_X1 U3708 ( .A1(n3182), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3213), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3186) );
  AOI21_X1 U3709 ( .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6596), .A(n3602), 
        .ZN(n3609) );
  OAI22_X1 U3710 ( .A1(n3601), .A2(n3600), .B1(n3610), .B2(n3629), .ZN(n3602)
         );
  AND2_X1 U3711 ( .A1(n3599), .A2(n3598), .ZN(n3600) );
  AOI211_X1 U3712 ( .C1(n3593), .C2(n3592), .A(n3591), .B(n3590), .ZN(n3601)
         );
  INV_X1 U3713 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6421) );
  OR2_X1 U3714 ( .A1(n6554), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4287) );
  NOR2_X1 U3715 ( .A1(n5329), .A2(n5945), .ZN(n5802) );
  AND3_X1 U3716 ( .A1(n3271), .A2(n4956), .A3(n4948), .ZN(n4949) );
  NOR2_X1 U3717 ( .A1(n4251), .A2(n5747), .ZN(n4252) );
  AND2_X1 U3718 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n4208), .ZN(n4209)
         );
  AND2_X1 U3719 ( .A1(n4166), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4167)
         );
  AND2_X1 U3720 ( .A1(n4170), .A2(n4169), .ZN(n5579) );
  AND2_X1 U3722 ( .A1(n4123), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4166)
         );
  AND2_X1 U3723 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n4075), .ZN(n4076)
         );
  NOR2_X1 U3724 ( .A1(n4026), .A2(n4025), .ZN(n4027) );
  NAND2_X1 U3725 ( .A1(n4027), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4074)
         );
  INV_X1 U3726 ( .A(n5310), .ZN(n4043) );
  AND2_X1 U3727 ( .A1(n3960), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n4005)
         );
  NAND2_X1 U3728 ( .A1(n4005), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4026)
         );
  NOR2_X1 U3729 ( .A1(n3974), .A2(n3956), .ZN(n3960) );
  NAND2_X1 U3730 ( .A1(n4018), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3974)
         );
  OR2_X1 U3731 ( .A1(n5359), .A2(n5290), .ZN(n5361) );
  NAND2_X1 U3732 ( .A1(n3923), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3924)
         );
  AND2_X1 U3733 ( .A1(n5156), .A2(n5183), .ZN(n3080) );
  NOR2_X1 U3734 ( .A1(n3877), .A2(n3861), .ZN(n3902) );
  NAND2_X1 U3735 ( .A1(n3860), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3877)
         );
  INV_X1 U3736 ( .A(n3859), .ZN(n3860) );
  CLKBUF_X1 U3737 ( .A(n4871), .Z(n4872) );
  NAND2_X1 U3738 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n3831), .ZN(n3837)
         );
  NAND2_X1 U3739 ( .A1(n3824), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3830)
         );
  NAND2_X1 U3740 ( .A1(n3822), .A2(n3821), .ZN(n4460) );
  OAI21_X1 U3741 ( .B1(n4635), .B2(n4022), .A(n3811), .ZN(n4481) );
  NAND2_X1 U3742 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3805) );
  NAND2_X1 U3743 ( .A1(n3800), .A2(n3799), .ZN(n3801) );
  NAND2_X1 U3744 ( .A1(n3787), .A2(n3283), .ZN(n3788) );
  NAND2_X1 U3745 ( .A1(n3107), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n3101) );
  NAND2_X1 U3746 ( .A1(n5620), .A2(n3107), .ZN(n5433) );
  INV_X1 U3747 ( .A(n5605), .ZN(n5606) );
  OR2_X1 U3748 ( .A1(n5875), .A2(n5468), .ZN(n5663) );
  NOR2_X1 U3749 ( .A1(n5583), .A2(n5406), .ZN(n5587) );
  AND2_X1 U3750 ( .A1(n5587), .A2(n5574), .ZN(n5576) );
  NAND2_X1 U3751 ( .A1(n2999), .A2(n3775), .ZN(n3776) );
  NAND2_X1 U3752 ( .A1(n3072), .A2(n3071), .ZN(n5583) );
  NOR2_X1 U3753 ( .A1(n5448), .A2(n5449), .ZN(n3071) );
  INV_X1 U3754 ( .A(n5711), .ZN(n3072) );
  NOR2_X1 U3755 ( .A1(n5320), .A2(n3721), .ZN(n5709) );
  NAND2_X1 U3756 ( .A1(n5709), .A2(n5708), .ZN(n5711) );
  AND2_X1 U3757 ( .A1(n5350), .A2(n5349), .ZN(n5905) );
  AOI21_X1 U3758 ( .B1(n3090), .B2(n3089), .A(n3050), .ZN(n3088) );
  INV_X1 U3759 ( .A(n5261), .ZN(n3090) );
  NOR2_X1 U3760 ( .A1(n5263), .A2(n5264), .ZN(n5350) );
  NAND2_X1 U3761 ( .A1(n3057), .A2(n3056), .ZN(n5263) );
  INV_X1 U3762 ( .A(n5234), .ZN(n3056) );
  INV_X1 U3763 ( .A(n5200), .ZN(n3057) );
  AND2_X1 U3764 ( .A1(n5158), .A2(n4304), .ZN(n5202) );
  NAND2_X1 U3765 ( .A1(n3095), .A2(n3097), .ZN(n5175) );
  INV_X1 U3766 ( .A(n3098), .ZN(n3097) );
  NAND2_X1 U3767 ( .A1(n3096), .A2(n3540), .ZN(n3095) );
  NOR2_X1 U3768 ( .A1(n5159), .A2(n5160), .ZN(n5158) );
  INV_X1 U3769 ( .A(n4969), .ZN(n3685) );
  INV_X1 U3770 ( .A(n4968), .ZN(n3069) );
  NAND2_X1 U3771 ( .A1(n3068), .A2(n3067), .ZN(n5159) );
  INV_X1 U3772 ( .A(n5063), .ZN(n3067) );
  NOR2_X1 U3773 ( .A1(n2999), .A2(n5068), .ZN(n5061) );
  NAND2_X1 U3774 ( .A1(n3671), .A2(n3070), .ZN(n4876) );
  NOR2_X1 U3775 ( .A1(n4465), .A2(n4584), .ZN(n3070) );
  NAND2_X1 U3776 ( .A1(n3671), .A2(n3670), .ZN(n4585) );
  INV_X1 U3777 ( .A(n3662), .ZN(n3059) );
  NOR2_X1 U3778 ( .A1(n4507), .A2(n3053), .ZN(n3058) );
  OAI21_X1 U3779 ( .B1(n3787), .B2(n3586), .A(n3463), .ZN(n6144) );
  AND2_X1 U3780 ( .A1(n3383), .A2(n3382), .ZN(n3464) );
  NAND2_X1 U3781 ( .A1(n3343), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3344) );
  OR2_X1 U3782 ( .A1(n3282), .A2(n3615), .ZN(n6410) );
  INV_X1 U3783 ( .A(n3389), .ZN(n3308) );
  NOR2_X1 U3784 ( .A1(n4336), .A2(n4471), .ZN(n6409) );
  INV_X1 U3785 ( .A(n3787), .ZN(n4763) );
  AND2_X1 U3786 ( .A1(n4634), .A2(n3803), .ZN(n6298) );
  AOI22_X1 U3787 ( .A1(n3392), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3140) );
  OR2_X1 U3788 ( .A1(n3035), .A2(n3787), .ZN(n4733) );
  AND2_X1 U3789 ( .A1(n4413), .A2(n4412), .ZN(n4452) );
  AND2_X1 U3790 ( .A1(n3035), .A2(n3787), .ZN(n6218) );
  INV_X1 U3791 ( .A(n4630), .ZN(n6353) );
  INV_X1 U3792 ( .A(n3289), .ZN(n3291) );
  OR2_X1 U3793 ( .A1(n5516), .A2(n6451), .ZN(n5727) );
  INV_X1 U3794 ( .A(n6042), .ZN(n5974) );
  INV_X1 U3795 ( .A(n6004), .ZN(n5980) );
  INV_X1 U3796 ( .A(n6003), .ZN(n6031) );
  INV_X1 U3797 ( .A(n5987), .ZN(n6020) );
  AND2_X1 U3798 ( .A1(n4955), .A2(n4956), .ZN(n6042) );
  AND2_X1 U3799 ( .A1(n5281), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6003) );
  AOI21_X1 U3800 ( .B1(n5484), .B2(n5550), .A(n5489), .ZN(n5430) );
  INV_X1 U3801 ( .A(n5597), .ZN(n6049) );
  NAND2_X1 U3802 ( .A1(n6053), .A2(n5598), .ZN(n5597) );
  INV_X1 U3803 ( .A(n3275), .ZN(n5598) );
  INV_X2 U3804 ( .A(n5504), .ZN(n6063) );
  INV_X1 U3805 ( .A(n6061), .ZN(n5603) );
  AOI21_X1 U3806 ( .B1(n6105), .B2(n4387), .A(n6469), .ZN(n6089) );
  CLKBUF_X1 U3807 ( .A(n6095), .Z(n6569) );
  INV_X2 U3808 ( .A(n6104), .ZN(n6097) );
  OR2_X1 U3809 ( .A1(n6089), .A2(n6569), .ZN(n6104) );
  INV_X1 U3810 ( .A(n4690), .ZN(n6125) );
  OR2_X1 U3811 ( .A1(n4315), .A2(n3259), .ZN(n6105) );
  INV_X1 U3812 ( .A(n4283), .ZN(n4284) );
  INV_X1 U3813 ( .A(n5496), .ZN(n5497) );
  NAND2_X1 U3814 ( .A1(n6148), .A2(n6146), .ZN(n6143) );
  INV_X1 U3815 ( .A(n6143), .ZN(n5860) );
  INV_X1 U3816 ( .A(n6148), .ZN(n6134) );
  AND2_X1 U3817 ( .A1(n5446), .A2(n3767), .ZN(n5883) );
  INV_X1 U3818 ( .A(n5883), .ZN(n5696) );
  OAI21_X1 U3819 ( .B1(n5640), .B2(n3558), .A(n3557), .ZN(n3559) );
  NAND2_X1 U3820 ( .A1(n3092), .A2(n3052), .ZN(n3087) );
  NAND2_X1 U3821 ( .A1(n4296), .A2(n3542), .ZN(n5215) );
  INV_X1 U3822 ( .A(n3061), .ZN(n3060) );
  AND2_X1 U3823 ( .A1(n5219), .A2(n6188), .ZN(n4390) );
  NOR2_X1 U3824 ( .A1(n5217), .A2(n3763), .ZN(n5887) );
  CLKBUF_X1 U3825 ( .A(n3782), .Z(n5721) );
  INV_X1 U3826 ( .A(n3803), .ZN(n4635) );
  INV_X1 U3827 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6548) );
  INV_X1 U3828 ( .A(n6211), .ZN(n4865) );
  INV_X1 U3829 ( .A(n5046), .ZN(n6360) );
  INV_X1 U3830 ( .A(n5022), .ZN(n6366) );
  INV_X1 U3831 ( .A(n5038), .ZN(n6378) );
  INV_X1 U3832 ( .A(n5052), .ZN(n6384) );
  AND2_X1 U3833 ( .A1(n4894), .A2(n6218), .ZN(n6401) );
  INV_X1 U3834 ( .A(n5030), .ZN(n6397) );
  AND2_X1 U3835 ( .A1(n6548), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6443) );
  OAI211_X1 U3836 ( .C1(n3066), .C2(n5538), .A(n3063), .B(n3062), .ZN(U2796)
         );
  INV_X1 U3837 ( .A(n5536), .ZN(n3066) );
  NAND2_X1 U3838 ( .A1(n5472), .A2(n6013), .ZN(n3062) );
  INV_X1 U3839 ( .A(n3064), .ZN(n3063) );
  OAI22_X1 U3840 ( .A1(n3787), .A2(n6344), .B1(n6412), .B2(n5722), .ZN(n4560)
         );
  NAND2_X1 U3841 ( .A1(n3275), .A2(n3248), .ZN(n3282) );
  XNOR2_X1 U3842 ( .A(n5430), .B(n5429), .ZN(n5534) );
  OR2_X1 U3843 ( .A1(n5864), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n3037)
         );
  INV_X1 U3844 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3804) );
  AND2_X1 U3845 ( .A1(n2999), .A2(n5863), .ZN(n3039) );
  NAND2_X1 U3846 ( .A1(n5572), .A2(n3082), .ZN(n3040) );
  NAND2_X1 U3847 ( .A1(n5648), .A2(n3077), .ZN(n5395) );
  CLKBUF_X3 U3848 ( .A(n5423), .Z(n5486) );
  OR2_X1 U3849 ( .A1(n5561), .A2(n5563), .ZN(n3041) );
  NOR2_X1 U3850 ( .A1(n2999), .A2(n5348), .ZN(n5261) );
  INV_X1 U3851 ( .A(n3549), .ZN(n5344) );
  AND2_X1 U3852 ( .A1(n5648), .A2(n5647), .ZN(n3042) );
  NOR2_X1 U3853 ( .A1(n2999), .A2(n5067), .ZN(n3043) );
  AND3_X1 U3854 ( .A1(n5729), .A2(REIP_REG_30__SCAN_IN), .A3(n5538), .ZN(n3044) );
  INV_X1 U3855 ( .A(n4399), .ZN(n3821) );
  AND2_X1 U3856 ( .A1(n3543), .A2(n3542), .ZN(n3045) );
  NAND2_X1 U3857 ( .A1(n5576), .A2(n5569), .ZN(n5561) );
  NAND2_X1 U3858 ( .A1(n5572), .A2(n5573), .ZN(n5566) );
  AND2_X1 U3859 ( .A1(n3517), .A2(n3503), .ZN(n3823) );
  NOR2_X1 U3860 ( .A1(n5261), .A2(n3091), .ZN(n3046) );
  NAND2_X1 U3861 ( .A1(n5905), .A2(n5904), .ZN(n5313) );
  AND2_X1 U3862 ( .A1(n5083), .A2(n5156), .ZN(n5154) );
  NAND2_X1 U3863 ( .A1(n5420), .A2(n4958), .ZN(n6035) );
  INV_X1 U3864 ( .A(n6035), .ZN(n6013) );
  NAND2_X1 U3865 ( .A1(n3015), .A2(n3539), .ZN(n4966) );
  NAND2_X1 U3866 ( .A1(n3087), .A2(n5225), .ZN(n5260) );
  AND2_X1 U3867 ( .A1(n3822), .A2(n3079), .ZN(n4461) );
  AND2_X1 U3868 ( .A1(n3492), .A2(n3435), .ZN(n3047) );
  AND2_X1 U3869 ( .A1(n4373), .A2(n3348), .ZN(n3048) );
  INV_X1 U3870 ( .A(n3292), .ZN(n3753) );
  AND2_X1 U3871 ( .A1(n4127), .A2(n3077), .ZN(n3049) );
  AND2_X2 U3872 ( .A1(n3038), .A2(n3451), .ZN(n5864) );
  INV_X1 U3873 ( .A(n4553), .ZN(n4403) );
  INV_X1 U3874 ( .A(n3078), .ZN(n6406) );
  NOR2_X1 U3875 ( .A1(n6348), .A2(n3787), .ZN(n3078) );
  INV_X1 U3876 ( .A(n3203), .ZN(n3637) );
  AND2_X1 U3877 ( .A1(n2999), .A2(n5348), .ZN(n3050) );
  AND2_X1 U3878 ( .A1(n5864), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3051)
         );
  NAND2_X1 U3879 ( .A1(n3069), .A2(n3685), .ZN(n5064) );
  INV_X1 U3880 ( .A(n5064), .ZN(n3068) );
  NAND2_X1 U3881 ( .A1(n2999), .A2(n3546), .ZN(n3052) );
  INV_X1 U3882 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4339) );
  AND2_X1 U3883 ( .A1(n3668), .A2(n3667), .ZN(n3053) );
  INV_X1 U3884 ( .A(n4140), .ZN(n4275) );
  NOR3_X4 U3885 ( .A1(n6063), .A2(n5598), .A3(n3252), .ZN(n6064) );
  AOI21_X1 U3886 ( .B1(n3823), .B2(n3983), .A(n3828), .ZN(n4459) );
  NOR2_X2 U3887 ( .A1(n4451), .A2(n6342), .ZN(n3983) );
  AND2_X4 U3888 ( .A1(n3125), .A2(n4358), .ZN(n3194) );
  AND2_X2 U3889 ( .A1(n3804), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3125)
         );
  NAND2_X1 U3890 ( .A1(n3059), .A2(n3058), .ZN(n4464) );
  NAND2_X1 U3891 ( .A1(n3061), .A2(n3053), .ZN(n4400) );
  OR2_X1 U3892 ( .A1(n4510), .A2(n3060), .ZN(n6034) );
  NOR3_X2 U3893 ( .A1(n5561), .A2(n5563), .A3(n5551), .ZN(n5483) );
  NAND3_X1 U3894 ( .A1(n3259), .A2(n3271), .A3(n3648), .ZN(n3074) );
  NAND2_X1 U3895 ( .A1(n3649), .A2(n3073), .ZN(n3653) );
  NAND3_X1 U3896 ( .A1(n3075), .A2(n5486), .A3(n3074), .ZN(n3073) );
  NAND2_X1 U3897 ( .A1(n5415), .A2(n3647), .ZN(n3075) );
  NAND2_X1 U3898 ( .A1(n3076), .A2(n3460), .ZN(n3459) );
  NAND3_X1 U3899 ( .A1(n3822), .A2(n3079), .A3(n4582), .ZN(n4581) );
  INV_X1 U3900 ( .A(n4581), .ZN(n3844) );
  NAND2_X1 U3901 ( .A1(n5083), .A2(n3080), .ZN(n5182) );
  NAND2_X1 U3902 ( .A1(n5199), .A2(n5198), .ZN(n5197) );
  XNOR2_X2 U3903 ( .A(n5182), .B(n3941), .ZN(n5199) );
  NOR2_X2 U3904 ( .A1(n5560), .A2(n5437), .ZN(n5498) );
  NAND2_X1 U3905 ( .A1(n3084), .A2(n3331), .ZN(n3303) );
  NAND2_X1 U3906 ( .A1(n3084), .A2(n3330), .ZN(n3332) );
  NAND2_X1 U3907 ( .A1(n3300), .A2(n3110), .ZN(n3084) );
  AND2_X2 U3908 ( .A1(n4533), .A2(n3085), .ZN(n3169) );
  AND2_X2 U3909 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4533) );
  NAND2_X1 U3910 ( .A1(n5605), .A2(n3776), .ZN(n5842) );
  AND2_X2 U3911 ( .A1(n3086), .A2(n4539), .ZN(n3398) );
  AND2_X2 U3912 ( .A1(n3021), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3086)
         );
  OAI21_X1 U3913 ( .B1(n3015), .B2(n3094), .A(n3093), .ZN(n5058) );
  AOI21_X1 U3914 ( .B1(n3100), .B2(n4967), .A(n3043), .ZN(n3093) );
  INV_X1 U3915 ( .A(n4967), .ZN(n3094) );
  OAI21_X1 U3916 ( .B1(n3099), .B2(n4967), .A(n5059), .ZN(n3098) );
  NAND2_X1 U3917 ( .A1(n3777), .A2(n3103), .ZN(n3102) );
  NOR2_X1 U3918 ( .A1(n3292), .A2(n3271), .ZN(n4311) );
  NAND2_X1 U3919 ( .A1(n3422), .A2(n3492), .ZN(n3502) );
  OR2_X2 U3920 ( .A1(n3201), .A2(n3200), .ZN(n3275) );
  INV_X1 U3921 ( .A(n5311), .ZN(n4044) );
  XNOR2_X1 U3922 ( .A(n3482), .B(n3452), .ZN(n3782) );
  INV_X1 U3923 ( .A(n3481), .ZN(n3452) );
  XNOR2_X1 U3924 ( .A(n3559), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5637)
         );
  CLKBUF_X1 U3925 ( .A(n4397), .Z(n4480) );
  INV_X1 U3926 ( .A(n3022), .ZN(n3310) );
  OR2_X1 U3927 ( .A1(n4386), .A2(n5507), .ZN(n4315) );
  AOI21_X1 U3928 ( .B1(n3820), .B2(n3983), .A(n3819), .ZN(n4399) );
  CLKBUF_X1 U3929 ( .A(n5455), .Z(n5541) );
  OAI21_X1 U3930 ( .B1(n5847), .B2(n5848), .A(n3552), .ZN(n5655) );
  AOI21_X1 U3931 ( .B1(n3782), .B2(n3983), .A(n4282), .ZN(n3798) );
  OAI21_X1 U3932 ( .B1(n5434), .B2(n5608), .A(n5433), .ZN(n5435) );
  AOI21_X1 U3933 ( .B1(n3842), .B2(n3983), .A(n3841), .ZN(n4873) );
  NAND2_X1 U3934 ( .A1(n5498), .A2(n5496), .ZN(n4285) );
  NAND2_X1 U3935 ( .A1(n4451), .A2(n3275), .ZN(n3294) );
  INV_X1 U3936 ( .A(n4451), .ZN(n3248) );
  NAND2_X1 U3937 ( .A1(n3293), .A2(n4451), .ZN(n3249) );
  NAND2_X1 U3938 ( .A1(n3549), .A2(n3548), .ZN(n5857) );
  XNOR2_X1 U3939 ( .A(n3513), .B(n4493), .ZN(n4487) );
  NAND2_X1 U3940 ( .A1(n3512), .A2(n3511), .ZN(n3513) );
  AND2_X1 U3941 ( .A1(n3281), .A2(n3280), .ZN(n3104) );
  NOR2_X1 U3942 ( .A1(n6220), .A2(n4761), .ZN(n3105) );
  NOR2_X1 U3943 ( .A1(n3035), .A2(n5925), .ZN(n3106) );
  AND2_X1 U3944 ( .A1(n2999), .A2(n5665), .ZN(n3107) );
  AND2_X1 U3945 ( .A1(n3770), .A2(n3769), .ZN(n3108) );
  NAND2_X1 U3946 ( .A1(n5443), .A2(n5444), .ZN(n3109) );
  INV_X1 U3947 ( .A(n3790), .ZN(n3909) );
  OR2_X1 U3948 ( .A1(n3299), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3110)
         );
  AND3_X1 U3949 ( .A1(n4952), .A2(n3281), .A3(n3257), .ZN(n3111) );
  AND2_X1 U3950 ( .A1(n5871), .A2(n5870), .ZN(n3112) );
  OR2_X1 U3951 ( .A1(n3607), .A2(n3635), .ZN(n3560) );
  AOI211_X1 U3952 ( .C1(n3589), .C2(n3588), .A(n3607), .B(n3587), .ZN(n3590)
         );
  AND2_X1 U3953 ( .A1(n6769), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3577)
         );
  INV_X1 U3954 ( .A(n3407), .ZN(n3408) );
  INV_X1 U3955 ( .A(n3494), .ZN(n3504) );
  INV_X1 U3956 ( .A(n5076), .ZN(n3876) );
  OR2_X1 U3957 ( .A1(n3445), .A2(n3444), .ZN(n3527) );
  NOR2_X1 U3958 ( .A1(n4122), .A2(n5641), .ZN(n4123) );
  OAI21_X1 U3959 ( .B1(n5857), .B2(INSTADDRPOINTER_REG_18__SCAN_IN), .A(n5864), 
        .ZN(n3550) );
  INV_X1 U3960 ( .A(n5085), .ZN(n3891) );
  OAI21_X1 U3961 ( .B1(n3599), .B2(n4722), .A(n3421), .ZN(n3492) );
  INV_X1 U3962 ( .A(n4465), .ZN(n3670) );
  AND2_X1 U3963 ( .A1(n4957), .A2(n5530), .ZN(n4958) );
  INV_X1 U3964 ( .A(n3909), .ZN(n4277) );
  OR2_X1 U3965 ( .A1(n4291), .A2(n6597), .ZN(n4292) );
  NOR2_X1 U3966 ( .A1(n6744), .A2(n3924), .ZN(n4018) );
  NAND2_X1 U3967 ( .A1(n3902), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3907)
         );
  OR2_X1 U3968 ( .A1(n3748), .A2(n3294), .ZN(n3737) );
  OAI21_X1 U3969 ( .B1(n6572), .B2(n4558), .A(n6445), .ZN(n4412) );
  OR2_X1 U3970 ( .A1(n5527), .A2(n5757), .ZN(n5537) );
  INV_X1 U3971 ( .A(n4074), .ZN(n4075) );
  NAND2_X1 U3972 ( .A1(n5525), .A2(n5292), .ZN(n5945) );
  INV_X1 U3973 ( .A(n3830), .ZN(n3831) );
  INV_X1 U3974 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3815) );
  OAI211_X1 U3975 ( .C1(n3836), .C2(n4275), .A(n3835), .B(n3834), .ZN(n4582)
         );
  AND2_X1 U3976 ( .A1(n4078), .A2(n4077), .ZN(n5647) );
  AND2_X1 U3977 ( .A1(n5381), .A2(n5380), .ZN(n5872) );
  NOR2_X1 U3978 ( .A1(n3907), .A2(n3903), .ZN(n3923) );
  INV_X1 U3979 ( .A(n4976), .ZN(n5075) );
  NAND2_X1 U3980 ( .A1(n5619), .A2(n3778), .ZN(n3779) );
  AND2_X1 U3981 ( .A1(n5611), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5612)
         );
  INV_X1 U3982 ( .A(n5911), .ZN(n6579) );
  OR2_X1 U3983 ( .A1(n3479), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6136)
         );
  INV_X1 U3984 ( .A(n5054), .ZN(n5013) );
  INV_X1 U3985 ( .A(n6291), .ZN(n4824) );
  INV_X1 U3986 ( .A(n4531), .ZN(n6032) );
  NAND2_X1 U3987 ( .A1(n6596), .A2(n4412), .ZN(n4713) );
  NAND2_X1 U3988 ( .A1(n4209), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4251)
         );
  NOR2_X1 U3989 ( .A1(n5526), .A2(n5783), .ZN(n5766) );
  NAND2_X1 U3990 ( .A1(n4076), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4122)
         );
  NAND2_X1 U3991 ( .A1(n3838), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3859)
         );
  NOR2_X1 U3992 ( .A1(n3816), .A2(n3815), .ZN(n3824) );
  AND2_X1 U3993 ( .A1(n5281), .A2(n4963), .ZN(n5979) );
  INV_X1 U3994 ( .A(n5796), .ZN(n5832) );
  AND2_X1 U3995 ( .A1(n5504), .A2(n4473), .ZN(n6061) );
  INV_X1 U3996 ( .A(n6105), .ZN(n6129) );
  NAND2_X1 U3997 ( .A1(n4167), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4207)
         );
  NOR2_X1 U3998 ( .A1(n3112), .A2(n5872), .ZN(n6057) );
  NAND2_X1 U3999 ( .A1(n5520), .A2(n4469), .ZN(n4386) );
  AND2_X1 U4000 ( .A1(n6155), .A2(n5885), .ZN(n5911) );
  OR2_X1 U4001 ( .A1(n3756), .A2(n3739), .ZN(n6584) );
  NOR2_X1 U4002 ( .A1(n4931), .A2(n4390), .ZN(n6176) );
  INV_X1 U4003 ( .A(n6584), .ZN(n6170) );
  INV_X1 U4004 ( .A(n4713), .ZN(n4839) );
  OR2_X1 U4005 ( .A1(n4715), .A2(n4714), .ZN(n6203) );
  INV_X1 U4006 ( .A(n4834), .ZN(n4867) );
  NOR2_X1 U4007 ( .A1(n4414), .A2(n4595), .ZN(n5054) );
  INV_X1 U4008 ( .A(n6295), .ZN(n6274) );
  AND2_X1 U4009 ( .A1(n6298), .A2(n4727), .ZN(n6291) );
  INV_X1 U4010 ( .A(n6337), .ZN(n6320) );
  INV_X1 U4011 ( .A(n6323), .ZN(n6331) );
  OAI21_X1 U4012 ( .B1(n4899), .B2(n6761), .A(n4898), .ZN(n4921) );
  INV_X1 U4013 ( .A(n5042), .ZN(n6345) );
  INV_X1 U4014 ( .A(n5026), .ZN(n6372) );
  INV_X1 U4015 ( .A(n5034), .ZN(n6391) );
  NAND2_X1 U4016 ( .A1(n5520), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6445) );
  NAND2_X1 U4017 ( .A1(n4315), .A2(n5727), .ZN(n6566) );
  NAND2_X1 U4018 ( .A1(n5281), .A2(n4946), .ZN(n6004) );
  INV_X1 U4019 ( .A(n5979), .ZN(n6036) );
  NAND2_X1 U4020 ( .A1(n4472), .A2(n6133), .ZN(n5504) );
  INV_X1 U4021 ( .A(n6089), .ZN(n6103) );
  INV_X1 U4022 ( .A(n6130), .ZN(n4690) );
  NAND2_X1 U4023 ( .A1(n5926), .A2(n4288), .ZN(n6148) );
  XNOR2_X1 U4024 ( .A(n5480), .B(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5503)
         );
  OR2_X1 U4025 ( .A1(n3756), .A2(n3645), .ZN(n6589) );
  INV_X1 U4026 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6769) );
  INV_X1 U4027 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6425) );
  OR2_X1 U4028 ( .A1(n4590), .A2(n4733), .ZN(n5149) );
  INV_X1 U4029 ( .A(n6401), .ZN(n6389) );
  INV_X1 U4030 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6761) );
  NAND2_X1 U4031 ( .A1(n4149), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3116)
         );
  NAND2_X1 U4032 ( .A1(n3182), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n3115)
         );
  NAND2_X1 U4033 ( .A1(n4154), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3114) );
  AND2_X2 U4034 ( .A1(n4367), .A2(n4539), .ZN(n3204) );
  NAND2_X1 U4035 ( .A1(n3204), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3113) );
  AND2_X2 U4036 ( .A1(n4367), .A2(n3125), .ZN(n3392) );
  NAND2_X1 U4037 ( .A1(n3392), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3120) );
  NAND2_X1 U4038 ( .A1(n3398), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3119) );
  AND2_X2 U4039 ( .A1(n4358), .A2(n4539), .ZN(n3238) );
  NAND2_X1 U4040 ( .A1(n3238), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3118) );
  NAND2_X1 U4041 ( .A1(n3213), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3117) );
  NAND2_X1 U4042 ( .A1(n3194), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3124) );
  AND2_X2 U4043 ( .A1(n3126), .A2(n4358), .ZN(n3195) );
  NAND2_X1 U4044 ( .A1(n3195), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3123) );
  NAND2_X1 U4045 ( .A1(n3169), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3122) );
  NAND2_X1 U4046 ( .A1(n3393), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3121)
         );
  AND2_X2 U4047 ( .A1(n3125), .A2(n4324), .ZN(n3354) );
  NAND2_X1 U4048 ( .A1(n3354), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3130) );
  AND2_X2 U4049 ( .A1(n3126), .A2(n4324), .ZN(n3349) );
  NAND2_X1 U4050 ( .A1(n3349), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3129)
         );
  NAND2_X1 U4051 ( .A1(n3189), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3128)
         );
  NAND2_X1 U4052 ( .A1(n3025), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3127)
         );
  AOI22_X1 U4053 ( .A1(n3182), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n3138) );
  AOI22_X1 U4054 ( .A1(n3398), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3169), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n3137) );
  AOI22_X1 U4055 ( .A1(n4154), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3195), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3136) );
  AOI22_X1 U4056 ( .A1(n3194), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3204), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3135) );
  AND4_X2 U4057 ( .A1(n3138), .A2(n3137), .A3(n3136), .A4(n3135), .ZN(n3144)
         );
  AOI22_X1 U4058 ( .A1(n3025), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(
        INSTQUEUE_REG_0__6__SCAN_IN), .B2(n3238), .ZN(n3142) );
  AOI22_X1 U4059 ( .A1(n3028), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3141) );
  AOI22_X1 U4060 ( .A1(n3354), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3213), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3139) );
  NAND2_X1 U4061 ( .A1(n3392), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3148) );
  NAND2_X1 U4062 ( .A1(n3032), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3147) );
  NAND2_X1 U4063 ( .A1(n3204), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3146) );
  NAND2_X1 U4064 ( .A1(n3036), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3145) );
  AND4_X2 U4065 ( .A1(n3148), .A2(n3147), .A3(n3146), .A4(n3145), .ZN(n3164)
         );
  NAND2_X1 U4066 ( .A1(n3030), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3152) );
  NAND2_X1 U4067 ( .A1(n3027), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3151)
         );
  NAND2_X1 U4068 ( .A1(n3354), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3150) );
  NAND2_X1 U4069 ( .A1(n3195), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3149) );
  AND4_X2 U4070 ( .A1(n3152), .A2(n3151), .A3(n3150), .A4(n3149), .ZN(n3163)
         );
  NAND2_X1 U4071 ( .A1(n3182), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3156)
         );
  NAND2_X1 U4072 ( .A1(n3349), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3155)
         );
  NAND2_X1 U4073 ( .A1(n3213), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3154) );
  NAND2_X1 U4074 ( .A1(n3024), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3153)
         );
  AND4_X2 U4075 ( .A1(n3156), .A2(n3155), .A3(n3154), .A4(n3153), .ZN(n3162)
         );
  NAND2_X1 U4076 ( .A1(n3398), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3160) );
  NAND2_X1 U4077 ( .A1(n3189), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3159)
         );
  NAND2_X1 U4078 ( .A1(n3238), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3158) );
  NAND2_X1 U4079 ( .A1(n3393), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3157)
         );
  BUF_X4 U4080 ( .A(n3195), .Z(n3177) );
  AOI22_X1 U4081 ( .A1(n3354), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3349), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3167) );
  AOI22_X1 U4082 ( .A1(n4149), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3166) );
  AOI22_X1 U4083 ( .A1(n3398), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3165) );
  AOI22_X1 U4084 ( .A1(n3194), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3204), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3173) );
  AOI22_X1 U4085 ( .A1(n3182), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3172) );
  AOI22_X1 U4086 ( .A1(n3392), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3169), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3170) );
  OAI211_X1 U4087 ( .C1(n4374), .C2(n4451), .A(n3249), .B(n3637), .ZN(n3202)
         );
  AOI22_X1 U4088 ( .A1(n3398), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3181) );
  AOI22_X1 U4089 ( .A1(n4154), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3354), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3180) );
  AOI22_X1 U4090 ( .A1(n3177), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3238), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3179) );
  AOI22_X1 U4091 ( .A1(n4149), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3178) );
  NAND4_X1 U4092 ( .A1(n3181), .A2(n3180), .A3(n3179), .A4(n3178), .ZN(n3188)
         );
  AOI22_X1 U4093 ( .A1(n3349), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3185) );
  AOI22_X1 U4094 ( .A1(n3392), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3169), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3184) );
  AOI22_X1 U4095 ( .A1(n3204), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3183) );
  NAND4_X1 U4096 ( .A1(n3186), .A2(n3185), .A3(n3184), .A4(n3183), .ZN(n3187)
         );
  NAND2_X1 U4097 ( .A1(n3260), .A2(n3274), .ZN(n3279) );
  AOI22_X1 U4098 ( .A1(n4149), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3182), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3193) );
  AOI22_X1 U4099 ( .A1(n4154), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3204), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3192) );
  AOI22_X1 U4100 ( .A1(n3349), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3189), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3191) );
  AOI22_X1 U4101 ( .A1(n3354), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3190) );
  NAND4_X1 U4102 ( .A1(n3193), .A2(n3192), .A3(n3191), .A4(n3190), .ZN(n3201)
         );
  AOI22_X1 U4103 ( .A1(n3392), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3023), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3199) );
  AOI22_X1 U4104 ( .A1(n3398), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3238), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3198) );
  AOI22_X1 U4105 ( .A1(n3194), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3169), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3197) );
  AOI22_X1 U4106 ( .A1(n3195), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3196) );
  NAND4_X1 U4107 ( .A1(n3199), .A2(n3198), .A3(n3197), .A4(n3196), .ZN(n3200)
         );
  NAND3_X1 U4108 ( .A1(n3202), .A2(n3279), .A3(n3275), .ZN(n3247) );
  NAND2_X1 U4109 ( .A1(n4149), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3208)
         );
  NAND2_X1 U4110 ( .A1(n3182), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3207)
         );
  NAND2_X1 U4111 ( .A1(n4154), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3206) );
  NAND2_X1 U4112 ( .A1(n3204), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3205) );
  NAND2_X1 U4113 ( .A1(n3194), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3212) );
  NAND2_X1 U4114 ( .A1(n3195), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3211) );
  NAND2_X1 U4115 ( .A1(n3169), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3210) );
  NAND2_X1 U4116 ( .A1(n3393), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3209)
         );
  NAND2_X1 U4117 ( .A1(n3398), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3217) );
  NAND2_X1 U4118 ( .A1(n3392), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3216) );
  NAND2_X1 U4119 ( .A1(n3238), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3215) );
  NAND2_X1 U4120 ( .A1(n3023), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3214) );
  NAND2_X1 U4121 ( .A1(n3354), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3221) );
  NAND2_X1 U4122 ( .A1(n3349), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3220)
         );
  NAND2_X1 U4123 ( .A1(n3189), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3219)
         );
  NAND2_X1 U4124 ( .A1(n3025), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3218)
         );
  NAND4_X4 U4125 ( .A1(n3225), .A2(n3224), .A3(n3223), .A4(n3222), .ZN(n3271)
         );
  NAND2_X1 U4126 ( .A1(n3392), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3229) );
  NAND2_X1 U4127 ( .A1(n3349), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3228)
         );
  NAND2_X1 U4128 ( .A1(n3189), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3227)
         );
  NAND2_X1 U4129 ( .A1(n3025), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3226)
         );
  NAND2_X1 U4130 ( .A1(n3182), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3233)
         );
  NAND2_X1 U4131 ( .A1(n3354), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3232) );
  NAND2_X1 U4132 ( .A1(n4154), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3231) );
  NAND2_X1 U4133 ( .A1(n3204), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3230) );
  NAND2_X1 U4134 ( .A1(n3194), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3237) );
  NAND2_X1 U4135 ( .A1(n4149), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3236)
         );
  NAND2_X1 U4136 ( .A1(n3195), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3235) );
  NAND2_X1 U4137 ( .A1(n3023), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3234) );
  NAND2_X1 U4138 ( .A1(n3398), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3242) );
  NAND2_X1 U4139 ( .A1(n3238), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3241) );
  NAND2_X1 U4140 ( .A1(n3036), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3240) );
  NAND2_X1 U4141 ( .A1(n3393), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3239)
         );
  NAND4_X4 U4142 ( .A1(n3246), .A2(n3245), .A3(n3244), .A4(n3243), .ZN(n3259)
         );
  INV_X1 U4143 ( .A(n3247), .ZN(n3251) );
  BUF_X2 U4144 ( .A(n3249), .Z(n4372) );
  INV_X1 U4145 ( .A(n3270), .ZN(n3254) );
  NAND2_X1 U4146 ( .A1(STATE_REG_1__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n6464) );
  OAI21_X1 U4147 ( .B1(STATE_REG_2__SCAN_IN), .B2(STATE_REG_1__SCAN_IN), .A(
        n6464), .ZN(n3255) );
  INV_X1 U4148 ( .A(n3255), .ZN(n3623) );
  INV_X1 U4149 ( .A(n3295), .ZN(n3256) );
  NAND2_X1 U4150 ( .A1(n3256), .A2(n3293), .ZN(n3257) );
  NAND2_X1 U4151 ( .A1(n3289), .A2(n6436), .ZN(n3264) );
  NAND2_X1 U4152 ( .A1(n3270), .A2(n3275), .ZN(n3262) );
  NAND2_X1 U4153 ( .A1(n3262), .A2(n3294), .ZN(n3263) );
  NAND3_X1 U4154 ( .A1(n3269), .A2(n3111), .A3(n3265), .ZN(n3266) );
  INV_X1 U4155 ( .A(n6443), .ZN(n3297) );
  NAND2_X1 U4156 ( .A1(n6761), .A2(n6548), .ZN(n6554) );
  INV_X1 U4157 ( .A(n4287), .ZN(n3298) );
  MUX2_X1 U4158 ( .A(n3297), .B(n3298), .S(n6769), .Z(n3267) );
  INV_X1 U4159 ( .A(n3267), .ZN(n3268) );
  INV_X1 U4160 ( .A(n4952), .ZN(n3754) );
  AND2_X1 U4161 ( .A1(n3203), .A2(n3271), .ZN(n3272) );
  NAND2_X1 U4162 ( .A1(n3260), .A2(n3273), .ZN(n3276) );
  NAND4_X1 U4163 ( .A1(n4372), .A2(n3276), .A3(n3274), .A4(n3275), .ZN(n3277)
         );
  NAND2_X1 U4164 ( .A1(n3277), .A2(n3259), .ZN(n3278) );
  OAI21_X1 U4165 ( .B1(n3289), .B2(n3279), .A(n6436), .ZN(n3285) );
  OR2_X1 U4166 ( .A1(n6554), .A2(n6596), .ZN(n6452) );
  INV_X1 U4167 ( .A(n6452), .ZN(n3280) );
  INV_X1 U4168 ( .A(n3282), .ZN(n3283) );
  INV_X1 U4169 ( .A(n3346), .ZN(n3288) );
  AND2_X1 U4170 ( .A1(n3471), .A2(n3293), .ZN(n3290) );
  NAND2_X1 U4171 ( .A1(n6437), .A2(n3271), .ZN(n5507) );
  NAND2_X1 U4172 ( .A1(n3753), .A2(n5519), .ZN(n3643) );
  NAND3_X1 U4173 ( .A1(n4373), .A2(n3293), .A3(n5519), .ZN(n3748) );
  OAI211_X1 U4174 ( .C1(n3295), .C2(n5507), .A(n3643), .B(n3737), .ZN(n3296)
         );
  NAND2_X1 U4175 ( .A1(n3296), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3301) );
  INV_X1 U4176 ( .A(n3301), .ZN(n3300) );
  XNOR2_X1 U4177 ( .A(n6769), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6220)
         );
  AOI22_X1 U4178 ( .A1(n3298), .A2(n6220), .B1(n3297), .B2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3302) );
  INV_X1 U4179 ( .A(n3302), .ZN(n3299) );
  INV_X1 U4180 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4369) );
  OAI211_X1 U4181 ( .C1(n3022), .C2(n4369), .A(n3302), .B(n3301), .ZN(n3330)
         );
  NAND2_X1 U4182 ( .A1(n3303), .A2(n3330), .ZN(n3390) );
  INV_X1 U4183 ( .A(n3390), .ZN(n3309) );
  NAND2_X1 U4184 ( .A1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3305) );
  NAND2_X1 U4185 ( .A1(n3305), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3306) );
  NOR2_X1 U4186 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6415), .ZN(n5108)
         );
  NAND2_X1 U4187 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5108), .ZN(n6296) );
  AND2_X1 U4188 ( .A1(n3306), .A2(n6296), .ZN(n4716) );
  OAI22_X1 U4189 ( .A1(n4287), .A2(n4716), .B1(n6443), .B2(n6421), .ZN(n3307)
         );
  NAND2_X1 U4190 ( .A1(n3310), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3314) );
  NOR3_X1 U4191 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6421), .A3(n6415), 
        .ZN(n6257) );
  NAND2_X1 U4192 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6257), .ZN(n6252) );
  NAND2_X1 U4193 ( .A1(n6425), .A2(n6252), .ZN(n3311) );
  NAND3_X1 U4194 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n6343) );
  INV_X1 U4195 ( .A(n6343), .ZN(n6355) );
  NAND2_X1 U4196 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6355), .ZN(n6339) );
  NAND2_X1 U4197 ( .A1(n3311), .A2(n6339), .ZN(n4761) );
  OAI22_X1 U4198 ( .A1(n4287), .A2(n4761), .B1(n6443), .B2(n6425), .ZN(n3312)
         );
  INV_X1 U4199 ( .A(n3312), .ZN(n3313) );
  NAND2_X1 U4200 ( .A1(n4531), .A2(n6596), .ZN(n3329) );
  INV_X1 U4201 ( .A(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3326) );
  AOI22_X1 U4202 ( .A1(n4085), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3319) );
  AOI22_X1 U4203 ( .A1(n4154), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3318) );
  AOI22_X1 U4204 ( .A1(n4155), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3317) );
  INV_X1 U4205 ( .A(n3354), .ZN(n3414) );
  AOI22_X1 U4206 ( .A1(n4214), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3316) );
  NAND4_X1 U4207 ( .A1(n3319), .A2(n3318), .A3(n3317), .A4(n3316), .ZN(n3325)
         );
  AOI22_X1 U4208 ( .A1(n4233), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3323) );
  AOI22_X1 U4209 ( .A1(n4097), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3322) );
  AOI22_X1 U4210 ( .A1(n3026), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3321) );
  AOI22_X1 U4211 ( .A1(n3177), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3320) );
  NAND4_X1 U4212 ( .A1(n3323), .A2(n3322), .A3(n3321), .A4(n3320), .ZN(n3324)
         );
  NOR2_X1 U4213 ( .A1(n3325), .A2(n3324), .ZN(n3485) );
  OAI22_X1 U4214 ( .A1(n3599), .A2(n3326), .B1(n3607), .B2(n3485), .ZN(n3327)
         );
  INV_X1 U4215 ( .A(n3327), .ZN(n3328) );
  NAND2_X1 U4216 ( .A1(n4357), .A2(n6596), .ZN(n3345) );
  AOI22_X1 U4217 ( .A1(n4233), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3336) );
  AOI22_X1 U4218 ( .A1(n4214), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4155), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3335) );
  AOI22_X1 U4219 ( .A1(n3182), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3334) );
  AOI22_X1 U4220 ( .A1(n3194), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3333) );
  NAND4_X1 U4221 ( .A1(n3336), .A2(n3335), .A3(n3334), .A4(n3333), .ZN(n3342)
         );
  AOI22_X1 U4222 ( .A1(n4097), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3340) );
  AOI22_X1 U4223 ( .A1(n4154), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3339) );
  AOI22_X1 U4224 ( .A1(n4259), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3338) );
  AOI22_X1 U4225 ( .A1(n4085), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3337) );
  NAND4_X1 U4226 ( .A1(n3340), .A2(n3339), .A3(n3338), .A4(n3337), .ZN(n3341)
         );
  NAND2_X1 U4227 ( .A1(n4374), .A2(n3469), .ZN(n3343) );
  NAND2_X1 U4228 ( .A1(n3345), .A2(n3344), .ZN(n3467) );
  INV_X1 U4229 ( .A(n3467), .ZN(n3385) );
  INV_X1 U4230 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4719) );
  AOI22_X1 U4231 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n4085), .B1(n3194), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3353) );
  AOI22_X1 U4232 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n4097), .B1(n4154), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3352) );
  AOI22_X1 U4233 ( .A1(n3182), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4155), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3351) );
  AOI22_X1 U4234 ( .A1(n3398), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3169), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3350) );
  NAND4_X1 U4235 ( .A1(n3353), .A2(n3352), .A3(n3351), .A4(n3350), .ZN(n3360)
         );
  AOI22_X1 U4236 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n3354), .B1(n4259), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3358) );
  AOI22_X1 U4237 ( .A1(n3000), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3357) );
  AOI22_X1 U4238 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(n4258), .B1(n3033), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3356) );
  AOI22_X1 U4239 ( .A1(n3177), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3355) );
  NAND4_X1 U4240 ( .A1(n3358), .A2(n3357), .A3(n3356), .A4(n3355), .ZN(n3359)
         );
  AOI21_X1 U4241 ( .B1(n3348), .B2(n3470), .A(n6596), .ZN(n3371) );
  AOI22_X1 U4242 ( .A1(n3398), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3364) );
  AOI22_X1 U4243 ( .A1(n3182), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4154), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3363) );
  AOI22_X1 U4244 ( .A1(n4214), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4155), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3362) );
  AOI22_X1 U4245 ( .A1(n3204), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3361) );
  NAND4_X1 U4246 ( .A1(n3364), .A2(n3363), .A3(n3362), .A4(n3361), .ZN(n3370)
         );
  AOI22_X1 U4247 ( .A1(n4259), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3368) );
  AOI22_X1 U4248 ( .A1(n3177), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3399), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4249 ( .A1(n3194), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4250 ( .A1(n4097), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3393), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3365) );
  NAND4_X1 U4251 ( .A1(n3368), .A2(n3367), .A3(n3366), .A4(n3365), .ZN(n3369)
         );
  INV_X1 U4252 ( .A(n3460), .ZN(n3374) );
  INV_X1 U4253 ( .A(n3534), .ZN(n3524) );
  NAND2_X1 U4254 ( .A1(n3524), .A2(n4374), .ZN(n3380) );
  MUX2_X1 U4255 ( .A(n3449), .B(n3380), .S(n3470), .Z(n3372) );
  INV_X1 U4256 ( .A(n3372), .ZN(n3373) );
  NAND2_X1 U4257 ( .A1(n3373), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3458) );
  INV_X1 U4258 ( .A(n3449), .ZN(n3375) );
  NAND2_X1 U4259 ( .A1(n3375), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3376) );
  NAND2_X1 U4260 ( .A1(n3567), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3383) );
  NAND2_X1 U4261 ( .A1(n3348), .A2(n3469), .ZN(n3379) );
  NAND2_X1 U4262 ( .A1(n3380), .A2(n3379), .ZN(n3381) );
  NAND2_X1 U4263 ( .A1(n3381), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3382) );
  NAND2_X1 U4264 ( .A1(n3385), .A2(n3384), .ZN(n3388) );
  NAND2_X1 U4265 ( .A1(n3390), .A2(n3389), .ZN(n3391) );
  AND2_X2 U4266 ( .A1(n4522), .A2(n3391), .ZN(n4340) );
  INV_X1 U4267 ( .A(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3406) );
  AOI22_X1 U4268 ( .A1(n4264), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4097), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3397) );
  AOI22_X1 U4269 ( .A1(n4214), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4155), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3396) );
  AOI22_X1 U4270 ( .A1(n3194), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3169), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3395) );
  AOI22_X1 U4271 ( .A1(n4177), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3394) );
  NAND4_X1 U4272 ( .A1(n3397), .A2(n3396), .A3(n3395), .A4(n3394), .ZN(n3405)
         );
  AOI22_X1 U4273 ( .A1(n4233), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3403) );
  AOI22_X1 U4274 ( .A1(n4154), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3402) );
  AOI22_X1 U4275 ( .A1(n4085), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3401) );
  AOI22_X1 U4276 ( .A1(n4258), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3400) );
  NAND4_X1 U4277 ( .A1(n3403), .A2(n3402), .A3(n3401), .A4(n3400), .ZN(n3404)
         );
  NOR2_X1 U4278 ( .A1(n3405), .A2(n3404), .ZN(n3453) );
  OAI22_X1 U4279 ( .A1(n3599), .A2(n3406), .B1(n3607), .B2(n3453), .ZN(n3407)
         );
  INV_X1 U4280 ( .A(n3493), .ZN(n3422) );
  INV_X1 U4281 ( .A(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4722) );
  AOI22_X1 U4282 ( .A1(n4233), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3413) );
  AOI22_X1 U4283 ( .A1(n4085), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3412) );
  AOI22_X1 U4284 ( .A1(n4097), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3411) );
  AOI22_X1 U4285 ( .A1(n4155), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3410) );
  NAND4_X1 U4286 ( .A1(n3413), .A2(n3412), .A3(n3411), .A4(n3410), .ZN(n3420)
         );
  INV_X2 U4287 ( .A(n3414), .ZN(n4214) );
  AOI22_X1 U4288 ( .A1(n4214), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3418) );
  AOI22_X1 U4289 ( .A1(n3031), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3417) );
  AOI22_X1 U4290 ( .A1(n3177), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3169), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3416) );
  AOI22_X1 U4291 ( .A1(n3182), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3415) );
  NAND4_X1 U4292 ( .A1(n3418), .A2(n3417), .A3(n3416), .A4(n3415), .ZN(n3419)
         );
  OR2_X1 U4293 ( .A1(n3607), .A2(n3504), .ZN(n3421) );
  INV_X1 U4294 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3434) );
  AOI22_X1 U4295 ( .A1(n4085), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3426) );
  AOI22_X1 U4296 ( .A1(n3031), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3425) );
  AOI22_X1 U4297 ( .A1(n4155), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3424) );
  AOI22_X1 U4298 ( .A1(n4214), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3423) );
  NAND4_X1 U4299 ( .A1(n3426), .A2(n3425), .A3(n3424), .A4(n3423), .ZN(n3432)
         );
  AOI22_X1 U4300 ( .A1(n4233), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3430) );
  INV_X1 U4301 ( .A(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n6763) );
  AOI22_X1 U4302 ( .A1(n4097), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3429) );
  AOI22_X1 U4303 ( .A1(n3026), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3169), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3428) );
  AOI22_X1 U4304 ( .A1(n3177), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3427) );
  NAND4_X1 U4305 ( .A1(n3430), .A2(n3429), .A3(n3428), .A4(n3427), .ZN(n3431)
         );
  NOR2_X1 U4306 ( .A1(n3432), .A2(n3431), .ZN(n3508) );
  OR2_X1 U4307 ( .A1(n3607), .A2(n3508), .ZN(n3433) );
  OAI21_X1 U4308 ( .B1(n3599), .B2(n3434), .A(n3433), .ZN(n3435) );
  INV_X1 U4309 ( .A(n3435), .ZN(n3501) );
  INV_X1 U4310 ( .A(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4725) );
  AOI22_X1 U4311 ( .A1(n3031), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3439) );
  AOI22_X1 U4312 ( .A1(n4258), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3438) );
  AOI22_X1 U4313 ( .A1(n4233), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3169), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3437) );
  AOI22_X1 U4314 ( .A1(n4097), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3436) );
  NAND4_X1 U4315 ( .A1(n3439), .A2(n3438), .A3(n3437), .A4(n3436), .ZN(n3445)
         );
  AOI22_X1 U4316 ( .A1(n4214), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n4155), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3443) );
  AOI22_X1 U4317 ( .A1(n3194), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3442) );
  AOI22_X1 U4318 ( .A1(n4085), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3441) );
  AOI22_X1 U4319 ( .A1(n3182), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n3440) );
  NAND4_X1 U4320 ( .A1(n3443), .A2(n3442), .A3(n3441), .A4(n3440), .ZN(n3444)
         );
  INV_X1 U4321 ( .A(n3527), .ZN(n3446) );
  OR2_X1 U4322 ( .A1(n3607), .A2(n3446), .ZN(n3447) );
  OAI21_X1 U4323 ( .B1(n3599), .B2(n4725), .A(n3447), .ZN(n3516) );
  INV_X1 U4324 ( .A(n3516), .ZN(n3448) );
  NAND2_X1 U4325 ( .A1(n3566), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3450) );
  NOR2_X1 U4326 ( .A1(n3450), .A2(n3449), .ZN(n3451) );
  NAND2_X1 U4327 ( .A1(n3782), .A2(n3566), .ZN(n3457) );
  NAND2_X1 U4328 ( .A1(n3470), .A2(n3469), .ZN(n3468) );
  NAND2_X1 U4329 ( .A1(n3468), .A2(n3453), .ZN(n3486) );
  OAI21_X1 U4330 ( .B1(n3453), .B2(n3468), .A(n3486), .ZN(n3455) );
  NAND2_X1 U4331 ( .A1(n3348), .A2(n3274), .ZN(n3461) );
  INV_X1 U4332 ( .A(n3461), .ZN(n3454) );
  AOI21_X1 U4333 ( .B1(n3455), .B2(n6436), .A(n3454), .ZN(n3456) );
  NAND2_X1 U4334 ( .A1(n3457), .A2(n3456), .ZN(n3479) );
  NAND2_X1 U4335 ( .A1(n3479), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n6135)
         );
  MUX2_X2 U4336 ( .A(n3460), .B(n3459), .S(n3458), .Z(n3787) );
  INV_X1 U4337 ( .A(n3566), .ZN(n3586) );
  INV_X1 U4338 ( .A(n6436), .ZN(n6571) );
  OAI21_X1 U4339 ( .B1(n6571), .B2(n3470), .A(n3461), .ZN(n3462) );
  INV_X1 U4340 ( .A(n3462), .ZN(n3463) );
  NAND2_X1 U4341 ( .A1(n6144), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n3476)
         );
  XNOR2_X1 U4342 ( .A(n3476), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4394)
         );
  XNOR2_X1 U4343 ( .A(n3465), .B(n3464), .ZN(n3466) );
  NAND2_X1 U4344 ( .A1(n3034), .A2(n3566), .ZN(n3475) );
  OAI21_X1 U4345 ( .B1(n3470), .B2(n3469), .A(n3468), .ZN(n3472) );
  OAI211_X1 U4346 ( .C1(n3472), .C2(n6571), .A(n3471), .B(n3252), .ZN(n3473)
         );
  INV_X1 U4347 ( .A(n3473), .ZN(n3474) );
  NAND2_X1 U4348 ( .A1(n4394), .A2(n4393), .ZN(n4392) );
  INV_X1 U4349 ( .A(n3476), .ZN(n3477) );
  NAND2_X1 U4350 ( .A1(n3477), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3478)
         );
  NAND2_X1 U4351 ( .A1(n6135), .A2(n6138), .ZN(n3480) );
  NAND2_X1 U4352 ( .A1(n3480), .A2(n6136), .ZN(n4499) );
  NAND2_X1 U4353 ( .A1(n3482), .A2(n3481), .ZN(n3483) );
  NAND2_X1 U4354 ( .A1(n3483), .A2(n4403), .ZN(n3484) );
  NAND2_X1 U4355 ( .A1(n3803), .A2(n3566), .ZN(n3489) );
  INV_X1 U4356 ( .A(n3485), .ZN(n3487) );
  NAND2_X1 U4357 ( .A1(n3486), .A2(n3487), .ZN(n3505) );
  OAI211_X1 U4358 ( .C1(n3487), .C2(n3486), .A(n3505), .B(n6436), .ZN(n3488)
         );
  NAND2_X1 U4359 ( .A1(n3489), .A2(n3488), .ZN(n3490) );
  NAND2_X1 U4360 ( .A1(n3490), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3491)
         );
  XNOR2_X1 U4361 ( .A(n3493), .B(n3492), .ZN(n3820) );
  NAND2_X1 U4362 ( .A1(n3820), .A2(n3566), .ZN(n3497) );
  XNOR2_X1 U4363 ( .A(n3505), .B(n3494), .ZN(n3495) );
  NAND2_X1 U4364 ( .A1(n3495), .A2(n6436), .ZN(n3496) );
  NAND2_X1 U4365 ( .A1(n3497), .A2(n3496), .ZN(n3498) );
  INV_X1 U4366 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3663) );
  XNOR2_X1 U4367 ( .A(n3498), .B(n3663), .ZN(n4517) );
  NAND2_X1 U4368 ( .A1(n4516), .A2(n4517), .ZN(n3500) );
  NAND2_X1 U4369 ( .A1(n3498), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3499)
         );
  NAND2_X1 U4370 ( .A1(n3500), .A2(n3499), .ZN(n4486) );
  NAND2_X1 U4371 ( .A1(n3502), .A2(n3501), .ZN(n3503) );
  NAND2_X1 U4372 ( .A1(n3823), .A2(n3566), .ZN(n3512) );
  NOR2_X1 U4373 ( .A1(n3505), .A2(n3504), .ZN(n3507) );
  INV_X1 U4374 ( .A(n3508), .ZN(n3506) );
  NAND2_X1 U4375 ( .A1(n3507), .A2(n3506), .ZN(n3526) );
  INV_X1 U4376 ( .A(n3507), .ZN(n3509) );
  AOI21_X1 U4377 ( .B1(n3509), .B2(n3508), .A(n6571), .ZN(n3510) );
  NAND2_X1 U4378 ( .A1(n3526), .A2(n3510), .ZN(n3511) );
  INV_X1 U4379 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4493) );
  NAND2_X1 U4380 ( .A1(n4486), .A2(n4487), .ZN(n3515) );
  NAND2_X1 U4381 ( .A1(n3513), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3514)
         );
  NAND2_X1 U4382 ( .A1(n3517), .A2(n3448), .ZN(n3833) );
  NAND3_X1 U4383 ( .A1(n3038), .A2(n3566), .A3(n3833), .ZN(n3520) );
  XNOR2_X1 U4384 ( .A(n3526), .B(n3527), .ZN(n3518) );
  NAND2_X1 U4385 ( .A1(n3518), .A2(n6436), .ZN(n3519) );
  NAND2_X1 U4386 ( .A1(n3520), .A2(n3519), .ZN(n3521) );
  INV_X1 U4387 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3672) );
  XNOR2_X1 U4388 ( .A(n3521), .B(n3672), .ZN(n4616) );
  NAND2_X1 U4389 ( .A1(n4615), .A2(n4616), .ZN(n3523) );
  NAND2_X1 U4390 ( .A1(n3521), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3522)
         );
  NAND2_X1 U4391 ( .A1(n3523), .A2(n3522), .ZN(n4885) );
  INV_X1 U4392 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n6608) );
  OAI22_X1 U4393 ( .A1(n3599), .A2(n6608), .B1(n3607), .B2(n3524), .ZN(n3525)
         );
  NAND2_X1 U4394 ( .A1(n3842), .A2(n3566), .ZN(n3531) );
  INV_X1 U4395 ( .A(n3526), .ZN(n3528) );
  NAND2_X1 U4396 ( .A1(n3528), .A2(n3527), .ZN(n3536) );
  XNOR2_X1 U4397 ( .A(n3536), .B(n3534), .ZN(n3529) );
  NAND2_X1 U4398 ( .A1(n3529), .A2(n6436), .ZN(n3530) );
  NAND2_X1 U4399 ( .A1(n3531), .A2(n3530), .ZN(n3532) );
  INV_X1 U4400 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6723) );
  XNOR2_X1 U4401 ( .A(n3532), .B(n6723), .ZN(n4886) );
  NAND2_X1 U4402 ( .A1(n3532), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3533)
         );
  NAND2_X1 U4403 ( .A1(n6436), .A2(n3534), .ZN(n3535) );
  OR2_X1 U4404 ( .A1(n3536), .A2(n3535), .ZN(n3537) );
  NAND2_X1 U4405 ( .A1(n2999), .A2(n3537), .ZN(n3538) );
  INV_X1 U4406 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3679) );
  XNOR2_X1 U4407 ( .A(n3538), .B(n3679), .ZN(n4929) );
  NAND2_X1 U4408 ( .A1(n3538), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3539)
         );
  XNOR2_X1 U4409 ( .A(n2999), .B(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4967)
         );
  INV_X1 U4410 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5067) );
  INV_X1 U4411 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n5068) );
  NAND2_X1 U4412 ( .A1(n2999), .A2(n5068), .ZN(n5059) );
  INV_X1 U4413 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6770) );
  XNOR2_X1 U4414 ( .A(n2999), .B(n6770), .ZN(n5176) );
  XNOR2_X1 U4415 ( .A(n2999), .B(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4297)
         );
  INV_X1 U4416 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n3692) );
  INV_X1 U4417 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3544) );
  XNOR2_X1 U4418 ( .A(n2999), .B(n3544), .ZN(n5216) );
  NAND2_X1 U4419 ( .A1(n2999), .A2(n3544), .ZN(n3545) );
  NAND2_X1 U4420 ( .A1(n5213), .A2(n3545), .ZN(n5227) );
  INV_X1 U4421 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3546) );
  INV_X1 U4422 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5348) );
  INV_X1 U4423 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5863) );
  NAND2_X1 U4424 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5466) );
  INV_X1 U4425 ( .A(n5466), .ZN(n3547) );
  NAND2_X1 U4426 ( .A1(n5854), .A2(n3547), .ZN(n3551) );
  NOR2_X1 U4427 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3548) );
  NAND2_X1 U4428 ( .A1(n3551), .A2(n3550), .ZN(n5847) );
  INV_X1 U4429 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n3713) );
  XNOR2_X1 U4430 ( .A(n2999), .B(n3713), .ZN(n5848) );
  NAND2_X1 U4431 ( .A1(n2999), .A2(n3713), .ZN(n3552) );
  INV_X1 U4432 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n3553) );
  XNOR2_X1 U4433 ( .A(n2999), .B(n3553), .ZN(n5656) );
  NOR2_X1 U4434 ( .A1(n5655), .A2(n5656), .ZN(n5443) );
  XNOR2_X1 U4435 ( .A(n2999), .B(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5650)
         );
  NAND2_X1 U4436 ( .A1(n5651), .A2(n5650), .ZN(n3554) );
  OAI21_X1 U4437 ( .B1(INSTADDRPOINTER_REG_21__SCAN_IN), .B2(n5864), .A(n3554), 
        .ZN(n5640) );
  NAND3_X1 U4438 ( .A1(n2999), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3558) );
  INV_X1 U4439 ( .A(n3554), .ZN(n3555) );
  NOR2_X1 U4440 ( .A1(n2999), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5638)
         );
  NAND2_X1 U4441 ( .A1(n3555), .A2(n5638), .ZN(n5445) );
  INV_X1 U4442 ( .A(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3556) );
  XNOR2_X1 U4443 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3576) );
  INV_X1 U4444 ( .A(n3576), .ZN(n3561) );
  XNOR2_X1 U4445 ( .A(n3561), .B(n3577), .ZN(n3625) );
  NAND2_X1 U4446 ( .A1(n3625), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3572) );
  INV_X1 U4447 ( .A(n3577), .ZN(n3563) );
  NAND2_X1 U4448 ( .A1(n3020), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3562) );
  NAND2_X1 U4449 ( .A1(n3563), .A2(n3562), .ZN(n3568) );
  INV_X1 U4450 ( .A(n3568), .ZN(n3564) );
  AOI21_X1 U4451 ( .B1(n3270), .B2(n3564), .A(n3348), .ZN(n3570) );
  AND2_X1 U4452 ( .A1(n3635), .A2(n3252), .ZN(n3565) );
  OAI21_X1 U4453 ( .B1(n3607), .B2(n3568), .A(n3610), .ZN(n3569) );
  OAI21_X1 U4454 ( .B1(n3570), .B2(n3580), .A(n3569), .ZN(n3571) );
  AOI22_X1 U4455 ( .A1(n3573), .A2(n3625), .B1(n3610), .B2(n3572), .ZN(n3574)
         );
  INV_X1 U4456 ( .A(n3589), .ZN(n3593) );
  XNOR2_X1 U4457 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3581) );
  NAND2_X1 U4458 ( .A1(n3577), .A2(n3576), .ZN(n3579) );
  NAND2_X1 U4459 ( .A1(n6415), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3578) );
  NAND2_X1 U4460 ( .A1(n3579), .A2(n3578), .ZN(n3582) );
  XOR2_X1 U4461 ( .A(n3581), .B(n3582), .Z(n3624) );
  OAI21_X1 U4462 ( .B1(n3624), .B2(n3599), .A(n3588), .ZN(n3592) );
  NAND2_X1 U4463 ( .A1(n3582), .A2(n3581), .ZN(n3584) );
  NAND2_X1 U4464 ( .A1(n6421), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3583) );
  NAND2_X1 U4465 ( .A1(n3584), .A2(n3583), .ZN(n3595) );
  XNOR2_X1 U4466 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3594) );
  INV_X1 U4467 ( .A(n3594), .ZN(n3585) );
  XNOR2_X1 U4468 ( .A(n3595), .B(n3585), .ZN(n3626) );
  NOR2_X1 U4469 ( .A1(n3586), .A2(n3626), .ZN(n3591) );
  INV_X1 U4470 ( .A(n3624), .ZN(n3587) );
  NAND2_X1 U4471 ( .A1(n3595), .A2(n3594), .ZN(n3597) );
  NAND2_X1 U4472 ( .A1(n6425), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3596) );
  NAND2_X1 U4473 ( .A1(n3597), .A2(n3596), .ZN(n3604) );
  INV_X1 U4474 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4523) );
  NAND2_X1 U4475 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n4523), .ZN(n3605) );
  NAND2_X1 U4476 ( .A1(n3629), .A2(n3626), .ZN(n3598) );
  INV_X1 U4477 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n6191) );
  AND2_X1 U4478 ( .A1(n6191), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3603)
         );
  OR2_X1 U4479 ( .A1(n3604), .A2(n3603), .ZN(n3606) );
  NAND2_X1 U4480 ( .A1(n3606), .A2(n3605), .ZN(n3628) );
  OR2_X1 U4481 ( .A1(n3607), .A2(n3628), .ZN(n3608) );
  INV_X1 U4482 ( .A(n3610), .ZN(n3612) );
  INV_X1 U4483 ( .A(n3628), .ZN(n3611) );
  NAND2_X1 U4484 ( .A1(n3612), .A2(n3611), .ZN(n3613) );
  NAND2_X1 U4485 ( .A1(n3273), .A2(n3252), .ZN(n3615) );
  NOR2_X1 U4486 ( .A1(n6410), .A2(n3635), .ZN(n3750) );
  INV_X1 U4487 ( .A(n3750), .ZN(n3633) );
  INV_X1 U4488 ( .A(n4311), .ZN(n5514) );
  INV_X1 U4489 ( .A(n3260), .ZN(n3616) );
  NAND2_X1 U4490 ( .A1(n3616), .A2(n6436), .ZN(n3617) );
  NAND2_X1 U4491 ( .A1(n3618), .A2(n3617), .ZN(n3744) );
  INV_X1 U4492 ( .A(n3744), .ZN(n3621) );
  NAND2_X1 U4493 ( .A1(n6410), .A2(n3348), .ZN(n3620) );
  AND2_X1 U4494 ( .A1(n3619), .A2(n3620), .ZN(n3642) );
  NAND2_X1 U4495 ( .A1(n3621), .A2(n3642), .ZN(n3622) );
  NAND2_X1 U4496 ( .A1(n5514), .A2(n3622), .ZN(n4330) );
  INV_X1 U4497 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6474) );
  NAND2_X1 U4498 ( .A1(n3623), .A2(n6474), .ZN(n6469) );
  NAND2_X1 U4499 ( .A1(n3259), .A2(n6469), .ZN(n3631) );
  NAND3_X1 U4500 ( .A1(n3626), .A2(n3625), .A3(n3624), .ZN(n3627) );
  NAND2_X1 U4501 ( .A1(n3628), .A2(n3627), .ZN(n3630) );
  AND2_X1 U4502 ( .A1(n3630), .A2(n3629), .ZN(n4310) );
  NOR2_X1 U4503 ( .A1(READY_N), .A2(n4310), .ZN(n4333) );
  NAND3_X1 U4504 ( .A1(n3631), .A2(n4333), .A3(n3203), .ZN(n3632) );
  OAI211_X1 U4505 ( .C1(n5520), .C2(n3633), .A(n4330), .B(n3632), .ZN(n3634)
         );
  NAND2_X1 U4506 ( .A1(n6443), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6451) );
  INV_X1 U4507 ( .A(n6451), .ZN(n4469) );
  NAND2_X1 U4508 ( .A1(n3634), .A2(n4469), .ZN(n3641) );
  NAND2_X1 U4509 ( .A1(n3635), .A2(n6469), .ZN(n4950) );
  INV_X1 U4510 ( .A(READY_N), .ZN(n6568) );
  NAND3_X1 U4511 ( .A1(n6437), .A2(n4950), .A3(n6568), .ZN(n3636) );
  NAND3_X1 U4512 ( .A1(n3636), .A2(n3271), .A3(n3294), .ZN(n3638) );
  NAND2_X1 U4513 ( .A1(n3638), .A2(n3637), .ZN(n3639) );
  OR2_X1 U4514 ( .A1(n4386), .A2(n3639), .ZN(n3640) );
  AND2_X1 U4515 ( .A1(n3642), .A2(n5519), .ZN(n4332) );
  INV_X1 U4516 ( .A(n4332), .ZN(n4345) );
  NAND2_X1 U4517 ( .A1(n3642), .A2(n3254), .ZN(n6427) );
  NAND2_X1 U4518 ( .A1(n4345), .A2(n6427), .ZN(n5508) );
  NAND2_X1 U4519 ( .A1(n6437), .A2(n5420), .ZN(n4325) );
  OAI211_X1 U4520 ( .C1(n4374), .C2(n3737), .A(n3643), .B(n4325), .ZN(n3644)
         );
  NOR2_X1 U4521 ( .A1(n5508), .A2(n3644), .ZN(n3645) );
  INV_X1 U4522 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3648) );
  INV_X1 U4523 ( .A(n3274), .ZN(n3646) );
  INV_X1 U4524 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n3647) );
  NAND2_X1 U4525 ( .A1(n3029), .A2(n3648), .ZN(n3649) );
  NAND2_X1 U4526 ( .A1(n5415), .A2(EBX_REG_0__SCAN_IN), .ZN(n3651) );
  INV_X1 U4527 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4959) );
  NAND2_X1 U4528 ( .A1(n5486), .A2(n4959), .ZN(n3650) );
  NAND2_X1 U4529 ( .A1(n3651), .A2(n3650), .ZN(n4681) );
  XNOR2_X1 U4530 ( .A(n3653), .B(n4681), .ZN(n4382) );
  NAND2_X1 U4531 ( .A1(n4382), .A2(n5420), .ZN(n4384) );
  INV_X1 U4532 ( .A(n4681), .ZN(n3652) );
  NAND2_X1 U4533 ( .A1(n4384), .A2(n3654), .ZN(n4507) );
  MUX2_X1 U4534 ( .A(n5411), .B(n5486), .S(EBX_REG_3__SCAN_IN), .Z(n3656) );
  OR2_X1 U4535 ( .A1(n5427), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3655)
         );
  INV_X1 U4536 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n3657) );
  NAND2_X1 U4537 ( .A1(n5415), .A2(n3657), .ZN(n3659) );
  INV_X1 U4538 ( .A(EBX_REG_2__SCAN_IN), .ZN(n6052) );
  NAND2_X1 U4539 ( .A1(n5420), .A2(n6052), .ZN(n3658) );
  NAND3_X1 U4540 ( .A1(n3659), .A2(n5486), .A3(n3658), .ZN(n3661) );
  NAND2_X1 U4541 ( .A1(n3029), .A2(n6052), .ZN(n3660) );
  NAND2_X1 U4542 ( .A1(n3661), .A2(n3660), .ZN(n5000) );
  NAND2_X1 U4543 ( .A1(n4508), .A2(n5000), .ZN(n3662) );
  NAND2_X1 U4544 ( .A1(n5415), .A2(n3663), .ZN(n3665) );
  INV_X1 U4545 ( .A(EBX_REG_4__SCAN_IN), .ZN(n3666) );
  NAND2_X1 U4546 ( .A1(n5420), .A2(n3666), .ZN(n3664) );
  NAND3_X1 U4547 ( .A1(n3665), .A2(n5486), .A3(n3664), .ZN(n3668) );
  NAND2_X1 U4548 ( .A1(n3029), .A2(n3666), .ZN(n3667) );
  INV_X1 U4549 ( .A(n4464), .ZN(n3671) );
  MUX2_X1 U4550 ( .A(n5411), .B(n5486), .S(EBX_REG_5__SCAN_IN), .Z(n3669) );
  OAI21_X1 U4551 ( .B1(INSTADDRPOINTER_REG_5__SCAN_IN), .B2(n5427), .A(n3669), 
        .ZN(n4465) );
  NAND2_X1 U4552 ( .A1(n5415), .A2(n3672), .ZN(n3674) );
  INV_X1 U4553 ( .A(EBX_REG_6__SCAN_IN), .ZN(n3675) );
  NAND2_X1 U4554 ( .A1(n5420), .A2(n3675), .ZN(n3673) );
  NAND3_X1 U4555 ( .A1(n3674), .A2(n5486), .A3(n3673), .ZN(n3677) );
  NAND2_X1 U4556 ( .A1(n3029), .A2(n3675), .ZN(n3676) );
  AND2_X1 U4557 ( .A1(n3677), .A2(n3676), .ZN(n4584) );
  MUX2_X1 U4558 ( .A(n5411), .B(n5486), .S(EBX_REG_7__SCAN_IN), .Z(n3678) );
  OAI21_X1 U4559 ( .B1(INSTADDRPOINTER_REG_7__SCAN_IN), .B2(n5427), .A(n3678), 
        .ZN(n4875) );
  NAND2_X1 U4560 ( .A1(n5415), .A2(n3679), .ZN(n3681) );
  INV_X1 U4561 ( .A(EBX_REG_8__SCAN_IN), .ZN(n5975) );
  NAND2_X1 U4562 ( .A1(n5420), .A2(n5975), .ZN(n3680) );
  NAND3_X1 U4563 ( .A1(n3681), .A2(n5486), .A3(n3680), .ZN(n3683) );
  NAND2_X1 U4564 ( .A1(n3029), .A2(n5975), .ZN(n3682) );
  NAND2_X1 U4565 ( .A1(n3683), .A2(n3682), .ZN(n4934) );
  NAND2_X1 U4566 ( .A1(n4935), .A2(n4934), .ZN(n4968) );
  MUX2_X1 U4567 ( .A(n5411), .B(n5486), .S(EBX_REG_9__SCAN_IN), .Z(n3684) );
  OAI21_X1 U4568 ( .B1(INSTADDRPOINTER_REG_9__SCAN_IN), .B2(n5427), .A(n3684), 
        .ZN(n4969) );
  NAND2_X1 U4569 ( .A1(n5415), .A2(n5068), .ZN(n3687) );
  INV_X1 U4570 ( .A(EBX_REG_10__SCAN_IN), .ZN(n6621) );
  NAND2_X1 U4571 ( .A1(n5420), .A2(n6621), .ZN(n3686) );
  NAND3_X1 U4572 ( .A1(n3687), .A2(n5486), .A3(n3686), .ZN(n3689) );
  NAND2_X1 U4573 ( .A1(n3029), .A2(n6621), .ZN(n3688) );
  AND2_X1 U4574 ( .A1(n3689), .A2(n3688), .ZN(n5063) );
  NAND2_X1 U4575 ( .A1(n5486), .A2(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n3690) );
  OAI211_X1 U4576 ( .C1(n5426), .C2(EBX_REG_11__SCAN_IN), .A(n5415), .B(n3690), 
        .ZN(n3691) );
  OAI21_X1 U4577 ( .B1(n5411), .B2(EBX_REG_11__SCAN_IN), .A(n3691), .ZN(n5160)
         );
  NAND2_X1 U4578 ( .A1(n5415), .A2(n3692), .ZN(n3694) );
  INV_X1 U4579 ( .A(EBX_REG_12__SCAN_IN), .ZN(n3695) );
  NAND2_X1 U4580 ( .A1(n5420), .A2(n3695), .ZN(n3693) );
  NAND3_X1 U4581 ( .A1(n3694), .A2(n5486), .A3(n3693), .ZN(n3697) );
  NAND2_X1 U4582 ( .A1(n3029), .A2(n3695), .ZN(n3696) );
  NAND2_X1 U4583 ( .A1(n3697), .A2(n3696), .ZN(n4304) );
  MUX2_X1 U4584 ( .A(n5411), .B(n5486), .S(EBX_REG_13__SCAN_IN), .Z(n3699) );
  OR2_X1 U4585 ( .A1(n5427), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n3698)
         );
  AND2_X1 U4586 ( .A1(n3699), .A2(n3698), .ZN(n5201) );
  NAND2_X1 U4587 ( .A1(n5202), .A2(n5201), .ZN(n5200) );
  NAND2_X1 U4588 ( .A1(n5486), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n3700) );
  NAND2_X1 U4589 ( .A1(n5415), .A2(n3700), .ZN(n3703) );
  INV_X1 U4590 ( .A(EBX_REG_14__SCAN_IN), .ZN(n3701) );
  NAND2_X1 U4591 ( .A1(n5420), .A2(n3701), .ZN(n3702) );
  AOI22_X1 U4592 ( .A1(n3703), .A2(n3702), .B1(n3029), .B2(n3701), .ZN(n5234)
         );
  NAND2_X1 U4593 ( .A1(n5486), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n3704) );
  OAI211_X1 U4594 ( .C1(n5426), .C2(EBX_REG_15__SCAN_IN), .A(n5415), .B(n3704), 
        .ZN(n3705) );
  OAI21_X1 U4595 ( .B1(n5411), .B2(EBX_REG_15__SCAN_IN), .A(n3705), .ZN(n5264)
         );
  NAND2_X1 U4596 ( .A1(n5427), .A2(EBX_REG_16__SCAN_IN), .ZN(n3707) );
  NAND2_X1 U4597 ( .A1(n5426), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n3706) );
  NAND2_X1 U4598 ( .A1(n3707), .A2(n3706), .ZN(n3708) );
  XNOR2_X1 U4599 ( .A(n3708), .B(n5486), .ZN(n5349) );
  INV_X1 U4600 ( .A(n5411), .ZN(n3709) );
  INV_X1 U4601 ( .A(EBX_REG_17__SCAN_IN), .ZN(n6048) );
  NAND2_X1 U4602 ( .A1(n3709), .A2(n6048), .ZN(n3712) );
  NAND2_X1 U4603 ( .A1(n5486), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3710) );
  OAI211_X1 U4604 ( .C1(n5426), .C2(EBX_REG_17__SCAN_IN), .A(n5415), .B(n3710), 
        .ZN(n3711) );
  AND2_X1 U4605 ( .A1(n3712), .A2(n3711), .ZN(n5904) );
  NAND2_X1 U4606 ( .A1(n5415), .A2(n3713), .ZN(n3715) );
  INV_X1 U4607 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5800) );
  NAND2_X1 U4608 ( .A1(n5420), .A2(n5800), .ZN(n3714) );
  NAND3_X1 U4609 ( .A1(n3715), .A2(n5486), .A3(n3714), .ZN(n3717) );
  NAND2_X1 U4610 ( .A1(n3029), .A2(n5800), .ZN(n3716) );
  AND2_X1 U4611 ( .A1(n3717), .A2(n3716), .ZN(n5316) );
  OR2_X1 U4612 ( .A1(n5427), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n3718)
         );
  INV_X1 U4613 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5393) );
  NAND2_X1 U4614 ( .A1(n5420), .A2(n5393), .ZN(n5314) );
  AND2_X1 U4615 ( .A1(n3718), .A2(n5314), .ZN(n5321) );
  OAI22_X1 U4616 ( .A1(n5427), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .B1(
        EBX_REG_20__SCAN_IN), .B2(n5426), .ZN(n5323) );
  NAND2_X1 U4617 ( .A1(n5321), .A2(n5323), .ZN(n3720) );
  NAND2_X1 U4618 ( .A1(n3029), .A2(EBX_REG_20__SCAN_IN), .ZN(n3719) );
  OAI211_X1 U4619 ( .C1(n5321), .C2(n3029), .A(n3720), .B(n3719), .ZN(n3721)
         );
  MUX2_X1 U4620 ( .A(n5411), .B(n5486), .S(EBX_REG_21__SCAN_IN), .Z(n3723) );
  OR2_X1 U4621 ( .A1(n5427), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n3722)
         );
  AND2_X1 U4622 ( .A1(n3723), .A2(n3722), .ZN(n5708) );
  NAND2_X1 U4623 ( .A1(n5486), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3724) );
  NAND2_X1 U4624 ( .A1(n5415), .A2(n3724), .ZN(n3726) );
  INV_X1 U4625 ( .A(EBX_REG_22__SCAN_IN), .ZN(n3727) );
  NAND2_X1 U4626 ( .A1(n5420), .A2(n3727), .ZN(n3725) );
  NAND2_X1 U4627 ( .A1(n3726), .A2(n3725), .ZN(n3729) );
  NAND2_X1 U4628 ( .A1(n3029), .A2(n3727), .ZN(n3728) );
  AND2_X1 U4629 ( .A1(n3729), .A2(n3728), .ZN(n5449) );
  NAND2_X1 U4630 ( .A1(n5486), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3730) );
  OAI211_X1 U4631 ( .C1(n5426), .C2(EBX_REG_23__SCAN_IN), .A(n5415), .B(n3730), 
        .ZN(n3731) );
  OAI21_X1 U4632 ( .B1(n5411), .B2(EBX_REG_23__SCAN_IN), .A(n3731), .ZN(n5448)
         );
  NAND2_X1 U4633 ( .A1(n5486), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3732) );
  NAND2_X1 U4634 ( .A1(n5415), .A2(n3732), .ZN(n3734) );
  INV_X1 U4635 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5543) );
  NAND2_X1 U4636 ( .A1(n5420), .A2(n5543), .ZN(n3733) );
  NAND2_X1 U4637 ( .A1(n3734), .A2(n3733), .ZN(n3736) );
  NAND2_X1 U4638 ( .A1(n3029), .A2(n5543), .ZN(n3735) );
  NAND2_X1 U4639 ( .A1(n3736), .A2(n3735), .ZN(n5585) );
  XNOR2_X1 U4640 ( .A(n5583), .B(n5585), .ZN(n5591) );
  INV_X1 U4641 ( .A(n3737), .ZN(n3738) );
  AOI22_X1 U4642 ( .A1(n3738), .A2(n4374), .B1(n6437), .B2(n6436), .ZN(n3739)
         );
  INV_X2 U4643 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6342) );
  NAND2_X1 U4644 ( .A1(n6596), .A2(n6342), .ZN(n6457) );
  OR2_X1 U4645 ( .A1(n6554), .A2(n6457), .ZN(n5908) );
  INV_X1 U4646 ( .A(REIP_REG_24__SCAN_IN), .ZN(n3740) );
  NOR2_X1 U4647 ( .A1(n5908), .A2(n3740), .ZN(n5631) );
  AOI21_X1 U4648 ( .B1(n5591), .B2(n6170), .A(n5631), .ZN(n3770) );
  NAND2_X1 U4649 ( .A1(INSTADDRPOINTER_REG_8__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n5066) );
  NAND2_X1 U4650 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n5069) );
  NOR2_X1 U4651 ( .A1(n5066), .A2(n5069), .ZN(n3752) );
  NAND2_X1 U4652 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3751) );
  INV_X1 U4653 ( .A(n5427), .ZN(n3747) );
  NAND2_X1 U4654 ( .A1(n3294), .A2(n3203), .ZN(n3741) );
  OR2_X1 U4655 ( .A1(n4952), .A2(n3203), .ZN(n4329) );
  NAND3_X1 U4656 ( .A1(n3742), .A2(n3741), .A3(n4329), .ZN(n3743) );
  NOR2_X1 U4657 ( .A1(n3744), .A2(n3743), .ZN(n3746) );
  OAI211_X1 U4658 ( .C1(n3619), .C2(n3747), .A(n3746), .B(n3745), .ZN(n4344)
         );
  INV_X1 U4659 ( .A(n6410), .ZN(n4359) );
  NAND2_X1 U4660 ( .A1(n4359), .A2(n3048), .ZN(n4534) );
  OAI21_X1 U4661 ( .B1(n3748), .B2(n3282), .A(n4534), .ZN(n3749) );
  NOR2_X1 U4662 ( .A1(n4344), .A2(n3749), .ZN(n3755) );
  NAND2_X1 U4663 ( .A1(n3755), .A2(n3750), .ZN(n5510) );
  AOI21_X1 U4664 ( .B1(INSTADDRPOINTER_REG_1__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .ZN(n4505) );
  NAND2_X1 U4665 ( .A1(INSTADDRPOINTER_REG_4__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4683) );
  NOR2_X1 U4666 ( .A1(n4505), .A2(n4683), .ZN(n4617) );
  NAND2_X1 U4667 ( .A1(n6171), .A2(n4617), .ZN(n4492) );
  NOR2_X1 U4668 ( .A1(n3751), .A2(n4492), .ZN(n4933) );
  NAND2_X1 U4669 ( .A1(n3752), .A2(n4933), .ZN(n5228) );
  NOR2_X1 U4670 ( .A1(n3751), .A2(n4683), .ZN(n4937) );
  AND3_X1 U4671 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n4937), .ZN(n4930) );
  AND2_X1 U4672 ( .A1(n3752), .A2(n4930), .ZN(n3757) );
  NAND2_X1 U4673 ( .A1(n3753), .A2(n3754), .ZN(n4532) );
  OR2_X1 U4674 ( .A1(n3756), .A2(n3755), .ZN(n5229) );
  INV_X1 U4675 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6188) );
  NAND2_X1 U4676 ( .A1(n3757), .A2(n6176), .ZN(n4299) );
  NAND2_X1 U4677 ( .A1(n5228), .A2(n4299), .ZN(n6155) );
  NAND2_X1 U4678 ( .A1(INSTADDRPOINTER_REG_16__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5355) );
  NAND2_X1 U4679 ( .A1(INSTADDRPOINTER_REG_12__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n5220) );
  NOR2_X1 U4680 ( .A1(n3544), .A2(n5220), .ZN(n5232) );
  NAND2_X1 U4681 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5232), .ZN(n5346) );
  NOR2_X1 U4682 ( .A1(n5355), .A2(n5346), .ZN(n5885) );
  NAND2_X1 U4683 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5884) );
  NOR2_X1 U4684 ( .A1(n5466), .A2(n5884), .ZN(n3760) );
  NAND2_X1 U4685 ( .A1(n5911), .A2(n3760), .ZN(n5712) );
  NAND2_X1 U4686 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5447) );
  NOR3_X1 U4687 ( .A1(n5712), .A2(n5447), .A3(n3556), .ZN(n3768) );
  INV_X1 U4688 ( .A(n5228), .ZN(n3758) );
  NAND2_X1 U4689 ( .A1(n5908), .A2(n3756), .ZN(n3759) );
  NAND2_X1 U4690 ( .A1(n4300), .A2(n5229), .ZN(n5217) );
  NAND2_X1 U4691 ( .A1(n6188), .A2(n5217), .ZN(n6182) );
  NAND2_X1 U4692 ( .A1(n3759), .A2(n6182), .ZN(n4389) );
  NOR2_X1 U4693 ( .A1(n6171), .A2(n4389), .ZN(n4932) );
  OAI22_X1 U4694 ( .A1(n3758), .A2(n4932), .B1(n4931), .B2(n3757), .ZN(n5266)
         );
  AND2_X1 U4695 ( .A1(n3759), .A2(n5219), .ZN(n6189) );
  INV_X1 U4696 ( .A(n5217), .ZN(n3761) );
  AOI22_X1 U4697 ( .A1(n6189), .A2(n3761), .B1(n5885), .B2(n3760), .ZN(n3762)
         );
  OR2_X1 U4698 ( .A1(n5266), .A2(n3762), .ZN(n5706) );
  INV_X1 U4699 ( .A(n5219), .ZN(n3763) );
  INV_X1 U4700 ( .A(n5447), .ZN(n3764) );
  NOR2_X1 U4701 ( .A1(n5887), .A2(n3764), .ZN(n3765) );
  NOR2_X1 U4702 ( .A1(n5706), .A2(n3765), .ZN(n5446) );
  AND2_X1 U4703 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n3774) );
  INV_X1 U4704 ( .A(n3774), .ZN(n3766) );
  OAI21_X1 U4705 ( .B1(n6176), .B2(n6171), .A(n3766), .ZN(n3767) );
  OAI21_X1 U4706 ( .B1(INSTADDRPOINTER_REG_24__SCAN_IN), .B2(n3768), .A(n5696), 
        .ZN(n3769) );
  OAI21_X1 U4707 ( .B1(n5637), .B2(n6589), .A(n3108), .ZN(U2994) );
  NOR2_X1 U4708 ( .A1(INSTADDRPOINTER_REG_20__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n5894) );
  NOR2_X1 U4709 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3772) );
  INV_X1 U4710 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n3771) );
  INV_X1 U4711 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5717) );
  NAND4_X1 U4712 ( .A1(n5894), .A2(n3772), .A3(n3771), .A4(n5717), .ZN(n3773)
         );
  NOR2_X1 U4713 ( .A1(n5447), .A2(n5884), .ZN(n5444) );
  AND2_X1 U4714 ( .A1(n5444), .A2(n3774), .ZN(n5467) );
  INV_X1 U4715 ( .A(n5467), .ZN(n3775) );
  XNOR2_X1 U4716 ( .A(n2999), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5841)
         );
  INV_X1 U4717 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5611) );
  AND2_X1 U4718 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5665) );
  INV_X1 U4719 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5664) );
  NAND2_X1 U4720 ( .A1(n5475), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3780) );
  INV_X1 U4721 ( .A(n3777), .ZN(n5619) );
  OR2_X1 U4722 ( .A1(n2999), .A2(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5618)
         );
  INV_X1 U4723 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5414) );
  INV_X1 U4724 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5681) );
  NAND2_X1 U4725 ( .A1(n5414), .A2(n5681), .ZN(n5674) );
  NOR2_X1 U4726 ( .A1(n5618), .A2(n5674), .ZN(n5432) );
  NAND2_X1 U4727 ( .A1(n5432), .A2(n5664), .ZN(n5476) );
  NOR2_X1 U4728 ( .A1(n5476), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3778)
         );
  NAND2_X1 U4729 ( .A1(n3780), .A2(n3779), .ZN(n3781) );
  XNOR2_X1 U4730 ( .A(n3781), .B(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n5474)
         );
  OR2_X2 U4731 ( .A1(n4386), .A2(n6427), .ZN(n5926) );
  NAND2_X1 U4732 ( .A1(n3035), .A2(n3983), .ZN(n3786) );
  NOR2_X1 U4733 ( .A1(n3275), .A2(n6342), .ZN(n3790) );
  AOI22_X1 U4734 ( .A1(n3790), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6342), .ZN(n3784) );
  NOR2_X1 U4735 ( .A1(n3294), .A2(n6342), .ZN(n3812) );
  NAND2_X1 U4736 ( .A1(n3812), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3783) );
  AND2_X1 U4737 ( .A1(n3784), .A2(n3783), .ZN(n3785) );
  NAND2_X1 U4738 ( .A1(n3788), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4476) );
  INV_X1 U4739 ( .A(n3812), .ZN(n3809) );
  NAND2_X1 U4740 ( .A1(PHYADDRPOINTER_REG_0__SCAN_IN), .A2(n6342), .ZN(n3792)
         );
  NAND2_X1 U4741 ( .A1(n3790), .A2(EAX_REG_0__SCAN_IN), .ZN(n3791) );
  OAI211_X1 U4742 ( .C1(n3809), .C2(n3020), .A(n3792), .B(n3791), .ZN(n3793)
         );
  AOI21_X1 U4743 ( .B1(n3789), .B2(n3983), .A(n3793), .ZN(n4475) );
  NOR2_X1 U4744 ( .A1(STATE2_REG_2__SCAN_IN), .A2(STATEBS16_REG_SCAN_IN), .ZN(
        n4140) );
  NAND2_X1 U4745 ( .A1(n4475), .A2(n4140), .ZN(n3794) );
  NAND2_X1 U4746 ( .A1(n4381), .A2(n4380), .ZN(n4379) );
  NAND2_X1 U4747 ( .A1(n3798), .A2(n4379), .ZN(n4484) );
  INV_X1 U4748 ( .A(EAX_REG_2__SCAN_IN), .ZN(n3797) );
  NAND2_X1 U4749 ( .A1(n3812), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3796) );
  INV_X1 U4750 ( .A(n4275), .ZN(n4278) );
  OAI21_X1 U4751 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3805), .ZN(n6142) );
  AOI22_X1 U4752 ( .A1(n4278), .A2(n6142), .B1(n4282), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3795) );
  OAI211_X1 U4753 ( .C1(n3909), .C2(n3797), .A(n3796), .B(n3795), .ZN(n4483)
         );
  NAND2_X1 U4754 ( .A1(n4484), .A2(n4483), .ZN(n3802) );
  INV_X1 U4755 ( .A(n3798), .ZN(n3800) );
  INV_X1 U4756 ( .A(n4379), .ZN(n3799) );
  INV_X1 U4757 ( .A(n3983), .ZN(n4022) );
  OAI21_X1 U4758 ( .B1(n3806), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n3816), 
        .ZN(n6037) );
  AOI22_X1 U4759 ( .A1(n6037), .A2(n4140), .B1(n4282), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3808) );
  NAND2_X1 U4760 ( .A1(n4277), .A2(EAX_REG_3__SCAN_IN), .ZN(n3807) );
  OAI211_X1 U4761 ( .C1(n3809), .C2(n3804), .A(n3808), .B(n3807), .ZN(n3810)
         );
  INV_X1 U4762 ( .A(n3810), .ZN(n3811) );
  NAND2_X1 U4763 ( .A1(n4479), .A2(n4481), .ZN(n4397) );
  NAND2_X1 U4764 ( .A1(n3812), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n3818) );
  INV_X1 U4765 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n5925) );
  OAI21_X1 U4766 ( .B1(PHYADDRPOINTER_REG_4__SCAN_IN), .B2(n5925), .A(n6342), 
        .ZN(n3813) );
  INV_X1 U4767 ( .A(n3813), .ZN(n3814) );
  AOI21_X1 U4768 ( .B1(n4277), .B2(EAX_REG_4__SCAN_IN), .A(n3814), .ZN(n3817)
         );
  AOI21_X1 U4769 ( .B1(n3816), .B2(n3815), .A(n3824), .ZN(n4518) );
  AOI22_X1 U4770 ( .A1(n3818), .A2(n3817), .B1(n4278), .B2(n4518), .ZN(n3819)
         );
  INV_X1 U4771 ( .A(EAX_REG_5__SCAN_IN), .ZN(n3827) );
  OAI21_X1 U4772 ( .B1(n3824), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3830), 
        .ZN(n6027) );
  NAND2_X1 U4773 ( .A1(n6027), .A2(n4140), .ZN(n3826) );
  NAND2_X1 U4774 ( .A1(n4282), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3825)
         );
  OAI211_X1 U4775 ( .C1(n3909), .C2(n3827), .A(n3826), .B(n3825), .ZN(n3828)
         );
  INV_X1 U4776 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3829) );
  NAND2_X1 U4777 ( .A1(n3830), .A2(n3829), .ZN(n3832) );
  NAND2_X1 U4778 ( .A1(n3832), .A2(n3837), .ZN(n6012) );
  INV_X1 U4779 ( .A(n6012), .ZN(n3836) );
  NAND2_X1 U4780 ( .A1(n3833), .A2(n3983), .ZN(n3835) );
  AOI22_X1 U4781 ( .A1(n4277), .A2(EAX_REG_6__SCAN_IN), .B1(n4282), .B2(
        PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3834) );
  OAI21_X1 U4782 ( .B1(n3838), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3859), 
        .ZN(n5998) );
  NAND2_X1 U4783 ( .A1(n5998), .A2(n4140), .ZN(n3840) );
  AOI22_X1 U4784 ( .A1(n4277), .A2(EAX_REG_7__SCAN_IN), .B1(n4282), .B2(
        PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3839) );
  NAND2_X1 U4785 ( .A1(n3840), .A2(n3839), .ZN(n3841) );
  NAND2_X1 U4786 ( .A1(n3844), .A2(n3843), .ZN(n4871) );
  XNOR2_X1 U4787 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .B(n3859), .ZN(n5978) );
  INV_X1 U4788 ( .A(n5978), .ZN(n4995) );
  AOI22_X1 U4789 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n4085), .B1(n4259), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3848) );
  AOI22_X1 U4790 ( .A1(n3177), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3847) );
  AOI22_X1 U4791 ( .A1(n4233), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4792 ( .A1(n3000), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3845) );
  NAND4_X1 U4793 ( .A1(n3848), .A2(n3847), .A3(n3846), .A4(n3845), .ZN(n3854)
         );
  AOI22_X1 U4794 ( .A1(n4097), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3852) );
  AOI22_X1 U4795 ( .A1(n3182), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3031), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3851) );
  AOI22_X1 U4796 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4214), .B1(n4155), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3850) );
  AOI22_X1 U4797 ( .A1(n3026), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3849) );
  NAND4_X1 U4798 ( .A1(n3852), .A2(n3851), .A3(n3850), .A4(n3849), .ZN(n3853)
         );
  OAI21_X1 U4799 ( .B1(n3854), .B2(n3853), .A(n3983), .ZN(n3857) );
  NAND2_X1 U4800 ( .A1(n4277), .A2(EAX_REG_8__SCAN_IN), .ZN(n3856) );
  NAND2_X1 U4801 ( .A1(n4282), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3855)
         );
  NAND3_X1 U4802 ( .A1(n3857), .A2(n3856), .A3(n3855), .ZN(n3858) );
  AOI21_X1 U4803 ( .B1(n4995), .B2(n4278), .A(n3858), .ZN(n4977) );
  INV_X1 U4804 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3861) );
  XNOR2_X1 U4805 ( .A(n3877), .B(n3861), .ZN(n5965) );
  AOI22_X1 U4806 ( .A1(n4264), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4097), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3865) );
  AOI22_X1 U4807 ( .A1(n4085), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3864) );
  AOI22_X1 U4808 ( .A1(n3026), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3863) );
  AOI22_X1 U4809 ( .A1(n3177), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3169), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3862) );
  NAND4_X1 U4810 ( .A1(n3865), .A2(n3864), .A3(n3863), .A4(n3862), .ZN(n3871)
         );
  AOI22_X1 U4811 ( .A1(n4233), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3869) );
  AOI22_X1 U4812 ( .A1(n3031), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3868) );
  AOI22_X1 U4813 ( .A1(n4155), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3867) );
  AOI22_X1 U4814 ( .A1(n4258), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3866) );
  NAND4_X1 U4815 ( .A1(n3869), .A2(n3868), .A3(n3867), .A4(n3866), .ZN(n3870)
         );
  OAI21_X1 U4816 ( .B1(n3871), .B2(n3870), .A(n3983), .ZN(n3874) );
  NAND2_X1 U4817 ( .A1(n4277), .A2(EAX_REG_9__SCAN_IN), .ZN(n3873) );
  NAND2_X1 U4818 ( .A1(n4282), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3872)
         );
  NAND3_X1 U4819 ( .A1(n3874), .A2(n3873), .A3(n3872), .ZN(n3875) );
  AOI21_X1 U4820 ( .B1(n5965), .B2(n4140), .A(n3875), .ZN(n5076) );
  NAND2_X1 U4821 ( .A1(n4976), .A2(n3876), .ZN(n5084) );
  XOR2_X1 U4822 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .B(n3902), .Z(n5958) );
  AOI22_X1 U4823 ( .A1(n4097), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3881) );
  AOI22_X1 U4824 ( .A1(n4264), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4155), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3880) );
  AOI22_X1 U4825 ( .A1(n4238), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3169), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3879) );
  AOI22_X1 U4826 ( .A1(n4258), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3878) );
  NAND4_X1 U4827 ( .A1(n3881), .A2(n3880), .A3(n3879), .A4(n3878), .ZN(n3887)
         );
  AOI22_X1 U4828 ( .A1(n4085), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3194), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4829 ( .A1(n4233), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4830 ( .A1(n3000), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3883) );
  AOI22_X1 U4831 ( .A1(n3031), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3882) );
  NAND4_X1 U4832 ( .A1(n3885), .A2(n3884), .A3(n3883), .A4(n3882), .ZN(n3886)
         );
  OR2_X1 U4833 ( .A1(n3887), .A2(n3886), .ZN(n3888) );
  AOI22_X1 U4834 ( .A1(n3983), .A2(n3888), .B1(n4282), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3890) );
  NAND2_X1 U4835 ( .A1(n4277), .A2(EAX_REG_10__SCAN_IN), .ZN(n3889) );
  OAI211_X1 U4836 ( .C1(n5958), .C2(n4275), .A(n3890), .B(n3889), .ZN(n5085)
         );
  AOI22_X1 U4837 ( .A1(n3026), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3895) );
  AOI22_X1 U4838 ( .A1(n4214), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4155), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3894) );
  AOI22_X1 U4839 ( .A1(n3031), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n3893) );
  AOI22_X1 U4840 ( .A1(n4233), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3892) );
  NAND4_X1 U4841 ( .A1(n3895), .A2(n3894), .A3(n3893), .A4(n3892), .ZN(n3901)
         );
  AOI22_X1 U4842 ( .A1(n4264), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4097), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n3899) );
  AOI22_X1 U4843 ( .A1(n4238), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3898) );
  AOI22_X1 U4844 ( .A1(n4259), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3897) );
  AOI22_X1 U4845 ( .A1(n4085), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3896) );
  NAND4_X1 U4846 ( .A1(n3899), .A2(n3898), .A3(n3897), .A4(n3896), .ZN(n3900)
         );
  NOR2_X1 U4847 ( .A1(n3901), .A2(n3900), .ZN(n3906) );
  INV_X1 U4848 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3903) );
  XNOR2_X1 U4849 ( .A(n3907), .B(n3903), .ZN(n5177) );
  NAND2_X1 U4850 ( .A1(n5177), .A2(n4140), .ZN(n3905) );
  AOI22_X1 U4851 ( .A1(n4277), .A2(EAX_REG_11__SCAN_IN), .B1(n4282), .B2(
        PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3904) );
  OAI211_X1 U4852 ( .C1(n3906), .C2(n4022), .A(n3905), .B(n3904), .ZN(n5156)
         );
  XOR2_X1 U4853 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3923), .Z(n5210) );
  INV_X1 U4854 ( .A(EAX_REG_12__SCAN_IN), .ZN(n3908) );
  INV_X1 U4855 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5206) );
  OAI22_X1 U4856 ( .A1(n3909), .A2(n3908), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n5206), .ZN(n3921) );
  AOI22_X1 U4857 ( .A1(n4264), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4858 ( .A1(n3031), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4859 ( .A1(n4155), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4860 ( .A1(n4085), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3910) );
  NAND4_X1 U4861 ( .A1(n3913), .A2(n3912), .A3(n3911), .A4(n3910), .ZN(n3919)
         );
  AOI22_X1 U4862 ( .A1(n4233), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3917) );
  AOI22_X1 U4863 ( .A1(n4097), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3916) );
  AOI22_X1 U4864 ( .A1(n3194), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3915) );
  AOI22_X1 U4865 ( .A1(n4238), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3914) );
  NAND4_X1 U4866 ( .A1(n3917), .A2(n3916), .A3(n3915), .A4(n3914), .ZN(n3918)
         );
  OR2_X1 U4867 ( .A1(n3919), .A2(n3918), .ZN(n3920) );
  AOI22_X1 U4868 ( .A1(n3921), .A2(n4275), .B1(n3983), .B2(n3920), .ZN(n3922)
         );
  OAI21_X1 U4869 ( .B1(n5210), .B2(n4275), .A(n3922), .ZN(n5183) );
  INV_X1 U4870 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6744) );
  NAND2_X1 U4871 ( .A1(n3924), .A2(n6744), .ZN(n3926) );
  INV_X1 U4872 ( .A(n4018), .ZN(n3925) );
  NAND2_X1 U4873 ( .A1(n3926), .A2(n3925), .ZN(n5255) );
  NAND2_X1 U4874 ( .A1(n5255), .A2(n4140), .ZN(n3929) );
  INV_X1 U4875 ( .A(n4282), .ZN(n4143) );
  NOR2_X1 U4876 ( .A1(n4143), .A2(n6744), .ZN(n3927) );
  AOI21_X1 U4877 ( .B1(n4277), .B2(EAX_REG_13__SCAN_IN), .A(n3927), .ZN(n3928)
         );
  NAND2_X1 U4878 ( .A1(n3929), .A2(n3928), .ZN(n3941) );
  AOI22_X1 U4879 ( .A1(n4097), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3031), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3933) );
  AOI22_X1 U4880 ( .A1(n3026), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3932) );
  AOI22_X1 U4881 ( .A1(n4233), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3931) );
  AOI22_X1 U4882 ( .A1(n4238), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3930) );
  NAND4_X1 U4883 ( .A1(n3933), .A2(n3932), .A3(n3931), .A4(n3930), .ZN(n3939)
         );
  AOI22_X1 U4884 ( .A1(n4155), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3937) );
  AOI22_X1 U4885 ( .A1(n4085), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3936) );
  AOI22_X1 U4886 ( .A1(n4264), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4887 ( .A1(n4214), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3934) );
  NAND4_X1 U4888 ( .A1(n3937), .A2(n3936), .A3(n3935), .A4(n3934), .ZN(n3938)
         );
  OR2_X1 U4889 ( .A1(n3939), .A2(n3938), .ZN(n3940) );
  AND2_X1 U4890 ( .A1(n3983), .A2(n3940), .ZN(n5198) );
  INV_X1 U4891 ( .A(n3941), .ZN(n3942) );
  NAND2_X1 U4892 ( .A1(n4359), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4249) );
  NAND2_X1 U4893 ( .A1(n4249), .A2(n4275), .ZN(n4093) );
  AOI22_X1 U4894 ( .A1(n4264), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3948) );
  AOI22_X1 U4895 ( .A1(n3000), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3947) );
  AOI22_X1 U4896 ( .A1(n4097), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3946) );
  NAND2_X1 U4897 ( .A1(n4214), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3944)
         );
  AOI21_X1 U4898 ( .B1(n3169), .B2(INSTQUEUE_REG_9__2__SCAN_IN), .A(n4278), 
        .ZN(n3943) );
  AND2_X1 U4899 ( .A1(n3944), .A2(n3943), .ZN(n3945) );
  NAND4_X1 U4900 ( .A1(n3948), .A2(n3947), .A3(n3946), .A4(n3945), .ZN(n3954)
         );
  AOI22_X1 U4901 ( .A1(n4233), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3026), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3952) );
  AOI22_X1 U4902 ( .A1(n4085), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3951) );
  AOI22_X1 U4903 ( .A1(n4155), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3950) );
  AOI22_X1 U4904 ( .A1(n3031), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3949) );
  NAND4_X1 U4905 ( .A1(n3952), .A2(n3951), .A3(n3950), .A4(n3949), .ZN(n3953)
         );
  OR2_X1 U4906 ( .A1(n3954), .A2(n3953), .ZN(n3955) );
  NAND2_X1 U4907 ( .A1(n4093), .A2(n3955), .ZN(n3959) );
  AOI22_X1 U4908 ( .A1(n3790), .A2(EAX_REG_18__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_18__SCAN_IN), .B2(n6342), .ZN(n3958) );
  INV_X1 U4909 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3956) );
  XNOR2_X1 U4910 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .B(n4026), .ZN(n5859)
         );
  AND2_X1 U4911 ( .A1(n4278), .A2(n5859), .ZN(n3957) );
  AOI21_X1 U4912 ( .B1(n3959), .B2(n3958), .A(n3957), .ZN(n5382) );
  XNOR2_X1 U4913 ( .A(n3960), .B(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5373)
         );
  AOI22_X1 U4914 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n4097), .B1(n3031), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3964) );
  AOI22_X1 U4915 ( .A1(n4085), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3963) );
  AOI22_X1 U4916 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n4259), .B1(n4155), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3962) );
  AOI22_X1 U4917 ( .A1(n4258), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3961) );
  NAND4_X1 U4918 ( .A1(n3964), .A2(n3963), .A3(n3962), .A4(n3961), .ZN(n3970)
         );
  AOI22_X1 U4919 ( .A1(n3194), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3968) );
  AOI22_X1 U4920 ( .A1(n4238), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3967) );
  AOI22_X1 U4921 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n4214), .B1(n4177), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3966) );
  AOI22_X1 U4922 ( .A1(n4233), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3965) );
  NAND4_X1 U4923 ( .A1(n3968), .A2(n3967), .A3(n3966), .A4(n3965), .ZN(n3969)
         );
  NOR2_X1 U4924 ( .A1(n3970), .A2(n3969), .ZN(n3972) );
  AOI22_X1 U4925 ( .A1(n3790), .A2(EAX_REG_16__SCAN_IN), .B1(n4282), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3971) );
  OAI21_X1 U4926 ( .B1(n4249), .B2(n3972), .A(n3971), .ZN(n3973) );
  AOI21_X1 U4927 ( .B1(n5373), .B2(n4278), .A(n3973), .ZN(n5362) );
  XNOR2_X1 U4928 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .B(n3974), .ZN(n5338)
         );
  INV_X1 U4929 ( .A(n5338), .ZN(n3990) );
  AOI22_X1 U4930 ( .A1(n4264), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3978) );
  AOI22_X1 U4931 ( .A1(n3000), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3977) );
  AOI22_X1 U4932 ( .A1(n3026), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3169), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4933 ( .A1(n4085), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3975) );
  NAND4_X1 U4934 ( .A1(n3978), .A2(n3977), .A3(n3976), .A4(n3975), .ZN(n3985)
         );
  AOI22_X1 U4935 ( .A1(n4233), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3982) );
  AOI22_X1 U4936 ( .A1(n3031), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3981) );
  AOI22_X1 U4937 ( .A1(n4155), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3980) );
  AOI22_X1 U4938 ( .A1(n4097), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3979) );
  NAND4_X1 U4939 ( .A1(n3982), .A2(n3981), .A3(n3980), .A4(n3979), .ZN(n3984)
         );
  OAI21_X1 U4940 ( .B1(n3985), .B2(n3984), .A(n3983), .ZN(n3988) );
  NAND2_X1 U4941 ( .A1(n4277), .A2(EAX_REG_15__SCAN_IN), .ZN(n3987) );
  NAND2_X1 U4942 ( .A1(n4282), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3986)
         );
  NAND3_X1 U4943 ( .A1(n3988), .A2(n3987), .A3(n3986), .ZN(n3989) );
  AOI21_X1 U4944 ( .B1(n3990), .B2(n4140), .A(n3989), .ZN(n5290) );
  OR2_X1 U4945 ( .A1(n5362), .A2(n5290), .ZN(n5358) );
  AOI22_X1 U4946 ( .A1(n4085), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U4947 ( .A1(n4238), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U4948 ( .A1(n3000), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U4949 ( .A1(n4155), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3991) );
  NAND4_X1 U4950 ( .A1(n3994), .A2(n3993), .A3(n3992), .A4(n3991), .ZN(n4000)
         );
  AOI22_X1 U4951 ( .A1(n4233), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3998) );
  AOI22_X1 U4952 ( .A1(n3194), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3997) );
  AOI22_X1 U4953 ( .A1(n4097), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3996) );
  AOI22_X1 U4954 ( .A1(n3031), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3995) );
  NAND4_X1 U4955 ( .A1(n3998), .A2(n3997), .A3(n3996), .A4(n3995), .ZN(n3999)
         );
  NOR2_X1 U4956 ( .A1(n4000), .A2(n3999), .ZN(n4004) );
  NAND2_X1 U4957 ( .A1(n6342), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4001)
         );
  NAND2_X1 U4958 ( .A1(n4275), .A2(n4001), .ZN(n4002) );
  AOI21_X1 U4959 ( .B1(n4277), .B2(EAX_REG_17__SCAN_IN), .A(n4002), .ZN(n4003)
         );
  OAI21_X1 U4960 ( .B1(n4249), .B2(n4004), .A(n4003), .ZN(n4007) );
  OAI21_X1 U4961 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n4005), .A(n4026), 
        .ZN(n5953) );
  OR2_X1 U4962 ( .A1(n4275), .A2(n5953), .ZN(n4006) );
  NAND2_X1 U4963 ( .A1(n4007), .A2(n4006), .ZN(n5870) );
  NOR2_X1 U4964 ( .A1(n5358), .A2(n5870), .ZN(n5380) );
  AND2_X1 U4965 ( .A1(n5382), .A2(n5380), .ZN(n4023) );
  AOI22_X1 U4966 ( .A1(n4233), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4011) );
  AOI22_X1 U4967 ( .A1(n4264), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4155), 
        .B2(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U4968 ( .A1(n4085), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U4969 ( .A1(n4214), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4008) );
  NAND4_X1 U4970 ( .A1(n4011), .A2(n4010), .A3(n4009), .A4(n4008), .ZN(n4017)
         );
  AOI22_X1 U4971 ( .A1(n3194), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4015) );
  AOI22_X1 U4972 ( .A1(n3031), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4014) );
  AOI22_X1 U4973 ( .A1(n4238), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4013) );
  AOI22_X1 U4974 ( .A1(n4097), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4012) );
  NAND4_X1 U4975 ( .A1(n4015), .A2(n4014), .A3(n4013), .A4(n4012), .ZN(n4016)
         );
  NOR2_X1 U4976 ( .A1(n4017), .A2(n4016), .ZN(n4021) );
  XNOR2_X1 U4977 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .B(n4018), .ZN(n5299)
         );
  AOI22_X1 U4978 ( .A1(n4278), .A2(n5299), .B1(n4282), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n4020) );
  NAND2_X1 U4979 ( .A1(n3790), .A2(EAX_REG_14__SCAN_IN), .ZN(n4019) );
  OAI211_X1 U4980 ( .C1(n4022), .C2(n4021), .A(n4020), .B(n4019), .ZN(n5379)
         );
  NAND2_X1 U4981 ( .A1(n5272), .A2(n4024), .ZN(n5311) );
  INV_X1 U4982 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n4025) );
  OR2_X1 U4983 ( .A1(n4027), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4028)
         );
  NAND2_X1 U4984 ( .A1(n4028), .A2(n4074), .ZN(n5849) );
  AOI22_X1 U4985 ( .A1(n4233), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4085), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4032) );
  AOI22_X1 U4986 ( .A1(n4264), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4097), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n4031) );
  AOI22_X1 U4987 ( .A1(n4238), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n4030) );
  AOI22_X1 U4988 ( .A1(n4259), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4029) );
  NAND4_X1 U4989 ( .A1(n4032), .A2(n4031), .A3(n4030), .A4(n4029), .ZN(n4038)
         );
  AOI22_X1 U4990 ( .A1(n3194), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4036) );
  AOI22_X1 U4991 ( .A1(n3031), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4035) );
  AOI22_X1 U4992 ( .A1(n4155), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4034) );
  AOI22_X1 U4993 ( .A1(n4258), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4033) );
  NAND4_X1 U4994 ( .A1(n4036), .A2(n4035), .A3(n4034), .A4(n4033), .ZN(n4037)
         );
  NOR2_X1 U4995 ( .A1(n4038), .A2(n4037), .ZN(n4041) );
  OAI21_X1 U4996 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n5925), .A(n6342), 
        .ZN(n4040) );
  NAND2_X1 U4997 ( .A1(n3790), .A2(EAX_REG_19__SCAN_IN), .ZN(n4039) );
  OAI211_X1 U4998 ( .C1(n4249), .C2(n4041), .A(n4040), .B(n4039), .ZN(n4042)
         );
  OAI21_X1 U4999 ( .B1(n5849), .B2(n4275), .A(n4042), .ZN(n5310) );
  AOI22_X1 U5000 ( .A1(n4097), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4048) );
  AOI22_X1 U5001 ( .A1(n4258), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4047) );
  AOI22_X1 U5002 ( .A1(n3000), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4046) );
  AOI22_X1 U5003 ( .A1(n3026), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4045) );
  NAND4_X1 U5004 ( .A1(n4048), .A2(n4047), .A3(n4046), .A4(n4045), .ZN(n4056)
         );
  AOI22_X1 U5005 ( .A1(n4233), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n4054) );
  AOI22_X1 U5006 ( .A1(n4085), .A2(INSTQUEUE_REG_1__4__SCAN_IN), .B1(n4214), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4053) );
  AOI22_X1 U5007 ( .A1(n3031), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4052) );
  NAND2_X1 U5008 ( .A1(n4155), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4050)
         );
  AOI21_X1 U5009 ( .B1(n3169), .B2(INSTQUEUE_REG_9__4__SCAN_IN), .A(n4278), 
        .ZN(n4049) );
  AND2_X1 U5010 ( .A1(n4050), .A2(n4049), .ZN(n4051) );
  NAND4_X1 U5011 ( .A1(n4054), .A2(n4053), .A3(n4052), .A4(n4051), .ZN(n4055)
         );
  OAI21_X1 U5012 ( .B1(n4056), .B2(n4055), .A(n4093), .ZN(n4058) );
  AOI22_X1 U5013 ( .A1(n3790), .A2(EAX_REG_20__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_20__SCAN_IN), .B2(n6342), .ZN(n4057) );
  NAND2_X1 U5014 ( .A1(n4058), .A2(n4057), .ZN(n4060) );
  XNOR2_X1 U5015 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .B(n4074), .ZN(n5661)
         );
  NAND2_X1 U5016 ( .A1(n4278), .A2(n5661), .ZN(n4059) );
  NAND2_X1 U5017 ( .A1(n4060), .A2(n4059), .ZN(n5319) );
  AOI22_X1 U5018 ( .A1(n4233), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3026), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4064) );
  AOI22_X1 U5019 ( .A1(n4085), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n4063) );
  AOI22_X1 U5020 ( .A1(n4097), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4062) );
  AOI22_X1 U5021 ( .A1(n3031), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4061) );
  NAND4_X1 U5022 ( .A1(n4064), .A2(n4063), .A3(n4062), .A4(n4061), .ZN(n4070)
         );
  AOI22_X1 U5023 ( .A1(n4155), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4068) );
  AOI22_X1 U5024 ( .A1(n4214), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4067) );
  AOI22_X1 U5025 ( .A1(n3000), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4066) );
  AOI22_X1 U5026 ( .A1(n4258), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4065) );
  NAND4_X1 U5027 ( .A1(n4068), .A2(n4067), .A3(n4066), .A4(n4065), .ZN(n4069)
         );
  NOR2_X1 U5028 ( .A1(n4070), .A2(n4069), .ZN(n4073) );
  INV_X1 U5029 ( .A(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5792) );
  OAI21_X1 U5030 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5792), .A(n4275), .ZN(
        n4071) );
  AOI21_X1 U5031 ( .B1(n4277), .B2(EAX_REG_21__SCAN_IN), .A(n4071), .ZN(n4072)
         );
  OAI21_X1 U5032 ( .B1(n4249), .B2(n4073), .A(n4072), .ZN(n4078) );
  OAI21_X1 U5033 ( .B1(n4076), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n4122), 
        .ZN(n5799) );
  OR2_X1 U5034 ( .A1(n5799), .A2(n4275), .ZN(n4077) );
  AOI22_X1 U5035 ( .A1(n3194), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4084) );
  AOI22_X1 U5036 ( .A1(n3031), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4083) );
  AOI22_X1 U5037 ( .A1(n3182), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4082) );
  NAND2_X1 U5038 ( .A1(n4155), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4080)
         );
  AOI21_X1 U5039 ( .B1(n3169), .B2(INSTQUEUE_REG_9__6__SCAN_IN), .A(n4278), 
        .ZN(n4079) );
  AND2_X1 U5040 ( .A1(n4080), .A2(n4079), .ZN(n4081) );
  NAND4_X1 U5041 ( .A1(n4084), .A2(n4083), .A3(n4082), .A4(n4081), .ZN(n4091)
         );
  AOI22_X1 U5042 ( .A1(n4085), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4089) );
  AOI22_X1 U5043 ( .A1(n4097), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4088) );
  AOI22_X1 U5044 ( .A1(n4214), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4087) );
  AOI22_X1 U5045 ( .A1(n4233), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4086) );
  NAND4_X1 U5046 ( .A1(n4089), .A2(n4088), .A3(n4087), .A4(n4086), .ZN(n4090)
         );
  OR2_X1 U5047 ( .A1(n4091), .A2(n4090), .ZN(n4092) );
  NAND2_X1 U5048 ( .A1(n4093), .A2(n4092), .ZN(n4096) );
  AOI22_X1 U5049 ( .A1(n3790), .A2(EAX_REG_22__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_22__SCAN_IN), .B2(n6342), .ZN(n4095) );
  XNOR2_X1 U5050 ( .A(n4122), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5645)
         );
  AND2_X1 U5051 ( .A1(n5645), .A2(n4278), .ZN(n4094) );
  AOI21_X1 U5052 ( .B1(n4096), .B2(n4095), .A(n4094), .ZN(n5396) );
  AOI22_X1 U5053 ( .A1(n4233), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n4097), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4101) );
  AOI22_X1 U5054 ( .A1(n4214), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4100) );
  AOI22_X1 U5055 ( .A1(n3026), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4099) );
  AOI22_X1 U5056 ( .A1(n3000), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4098) );
  NAND4_X1 U5057 ( .A1(n4101), .A2(n4100), .A3(n4099), .A4(n4098), .ZN(n4107)
         );
  AOI22_X1 U5058 ( .A1(n4264), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3177), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4105) );
  AOI22_X1 U5059 ( .A1(n3031), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4104) );
  AOI22_X1 U5060 ( .A1(n4085), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4103) );
  AOI22_X1 U5061 ( .A1(n4155), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4102) );
  NAND4_X1 U5062 ( .A1(n4105), .A2(n4104), .A3(n4103), .A4(n4102), .ZN(n4106)
         );
  NOR2_X1 U5063 ( .A1(n4107), .A2(n4106), .ZN(n4128) );
  AOI22_X1 U5064 ( .A1(n4097), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4111) );
  AOI22_X1 U5065 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n4155), .B1(n4259), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n4110) );
  AOI22_X1 U5066 ( .A1(n4214), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4109) );
  AOI22_X1 U5067 ( .A1(n4233), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4108) );
  NAND4_X1 U5068 ( .A1(n4111), .A2(n4110), .A3(n4109), .A4(n4108), .ZN(n4117)
         );
  AOI22_X1 U5069 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n4264), .B1(n3031), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n4115) );
  AOI22_X1 U5070 ( .A1(n3026), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4114) );
  AOI22_X1 U5071 ( .A1(n4085), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4113) );
  AOI22_X1 U5072 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n3033), .B1(n4177), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4112) );
  NAND4_X1 U5073 ( .A1(n4115), .A2(n4114), .A3(n4113), .A4(n4112), .ZN(n4116)
         );
  NOR2_X1 U5074 ( .A1(n4117), .A2(n4116), .ZN(n4129) );
  XNOR2_X1 U5075 ( .A(n4128), .B(n4129), .ZN(n4121) );
  NAND2_X1 U5076 ( .A1(n6342), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4118)
         );
  NAND2_X1 U5077 ( .A1(n4275), .A2(n4118), .ZN(n4119) );
  AOI21_X1 U5078 ( .B1(n4277), .B2(EAX_REG_23__SCAN_IN), .A(n4119), .ZN(n4120)
         );
  OAI21_X1 U5079 ( .B1(n4249), .B2(n4121), .A(n4120), .ZN(n4126) );
  INV_X1 U5080 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5641) );
  NOR2_X1 U5081 ( .A1(n4123), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4124)
         );
  OR2_X1 U5082 ( .A1(n4166), .A2(n4124), .ZN(n5460) );
  INV_X1 U5083 ( .A(n5460), .ZN(n5787) );
  NAND2_X1 U5084 ( .A1(n5787), .A2(n4140), .ZN(n4125) );
  NAND2_X1 U5085 ( .A1(n4126), .A2(n4125), .ZN(n5456) );
  OR2_X1 U5086 ( .A1(n4129), .A2(n4128), .ZN(n4148) );
  AOI22_X1 U5087 ( .A1(n4233), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3031), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n4133) );
  AOI22_X1 U5088 ( .A1(n4258), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n4155), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n4132) );
  AOI22_X1 U5089 ( .A1(n4214), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4131) );
  AOI22_X1 U5090 ( .A1(n4259), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4130) );
  NAND4_X1 U5091 ( .A1(n4133), .A2(n4132), .A3(n4131), .A4(n4130), .ZN(n4139)
         );
  AOI22_X1 U5092 ( .A1(n4085), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4137) );
  AOI22_X1 U5093 ( .A1(n3026), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4136) );
  AOI22_X1 U5094 ( .A1(n4264), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4135) );
  AOI22_X1 U5095 ( .A1(n4097), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4134) );
  NAND4_X1 U5096 ( .A1(n4137), .A2(n4136), .A3(n4135), .A4(n4134), .ZN(n4138)
         );
  OR2_X1 U5097 ( .A1(n4139), .A2(n4138), .ZN(n4146) );
  XNOR2_X1 U5098 ( .A(n4148), .B(n4146), .ZN(n4145) );
  INV_X1 U5099 ( .A(n4249), .ZN(n4273) );
  INV_X1 U5100 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5544) );
  NAND2_X1 U5101 ( .A1(n4277), .A2(EAX_REG_24__SCAN_IN), .ZN(n4142) );
  XNOR2_X1 U5102 ( .A(n4166), .B(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n5633)
         );
  NAND2_X1 U5103 ( .A1(n5633), .A2(n4140), .ZN(n4141) );
  OAI211_X1 U5104 ( .C1(n5544), .C2(n4143), .A(n4142), .B(n4141), .ZN(n4144)
         );
  AOI21_X1 U5105 ( .B1(n4145), .B2(n4273), .A(n4144), .ZN(n5542) );
  INV_X1 U5106 ( .A(n4146), .ZN(n4147) );
  OR2_X1 U5107 ( .A1(n4148), .A2(n4147), .ZN(n4171) );
  AOI22_X1 U5108 ( .A1(n4214), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n4153) );
  AOI22_X1 U5109 ( .A1(n4085), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4152) );
  AOI22_X1 U5110 ( .A1(n4264), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4151) );
  AOI22_X1 U5111 ( .A1(n3026), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4150) );
  NAND4_X1 U5112 ( .A1(n4153), .A2(n4152), .A3(n4151), .A4(n4150), .ZN(n4161)
         );
  AOI22_X1 U5113 ( .A1(n4097), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3031), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n4159) );
  AOI22_X1 U5114 ( .A1(n4258), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n4155), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4158) );
  AOI22_X1 U5115 ( .A1(n4233), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4157) );
  AOI22_X1 U5116 ( .A1(n4238), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n4156) );
  NAND4_X1 U5117 ( .A1(n4159), .A2(n4158), .A3(n4157), .A4(n4156), .ZN(n4160)
         );
  NOR2_X1 U5118 ( .A1(n4161), .A2(n4160), .ZN(n4172) );
  XNOR2_X1 U5119 ( .A(n4171), .B(n4172), .ZN(n4165) );
  INV_X1 U5120 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4162) );
  AOI21_X1 U5121 ( .B1(n4162), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4163) );
  AOI21_X1 U5122 ( .B1(n4277), .B2(EAX_REG_25__SCAN_IN), .A(n4163), .ZN(n4164)
         );
  OAI21_X1 U5123 ( .B1(n4165), .B2(n4249), .A(n4164), .ZN(n4170) );
  OR2_X1 U5124 ( .A1(n4167), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4168)
         );
  NAND2_X1 U5125 ( .A1(n4168), .A2(n4207), .ZN(n5846) );
  INV_X1 U5126 ( .A(n5846), .ZN(n5779) );
  NAND2_X1 U5127 ( .A1(n5779), .A2(n4278), .ZN(n4169) );
  AND2_X2 U5128 ( .A1(n5540), .A2(n5579), .ZN(n5572) );
  NOR2_X1 U5129 ( .A1(n4172), .A2(n4171), .ZN(n4192) );
  AOI22_X1 U5130 ( .A1(n4085), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4176) );
  AOI22_X1 U5131 ( .A1(n3031), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4175) );
  AOI22_X1 U5132 ( .A1(n4155), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4174) );
  AOI22_X1 U5133 ( .A1(n4214), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4173) );
  NAND4_X1 U5134 ( .A1(n4176), .A2(n4175), .A3(n4174), .A4(n4173), .ZN(n4183)
         );
  AOI22_X1 U5135 ( .A1(n4233), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4181) );
  AOI22_X1 U5136 ( .A1(n4097), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4180) );
  AOI22_X1 U5137 ( .A1(n3026), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3169), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4179) );
  AOI22_X1 U5138 ( .A1(n4238), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4178) );
  NAND4_X1 U5139 ( .A1(n4181), .A2(n4180), .A3(n4179), .A4(n4178), .ZN(n4182)
         );
  OR2_X1 U5140 ( .A1(n4183), .A2(n4182), .ZN(n4191) );
  INV_X1 U5141 ( .A(n4191), .ZN(n4184) );
  XNOR2_X1 U5142 ( .A(n4192), .B(n4184), .ZN(n4185) );
  NAND2_X1 U5143 ( .A1(n4185), .A2(n4273), .ZN(n4190) );
  NAND2_X1 U5144 ( .A1(n6342), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4186)
         );
  NAND2_X1 U5145 ( .A1(n4275), .A2(n4186), .ZN(n4187) );
  AOI21_X1 U5146 ( .B1(n4277), .B2(EAX_REG_26__SCAN_IN), .A(n4187), .ZN(n4189)
         );
  XNOR2_X1 U5147 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .B(n4207), .ZN(n5765)
         );
  AND2_X1 U5148 ( .A1(n5765), .A2(n4278), .ZN(n4188) );
  AOI21_X1 U5149 ( .B1(n4190), .B2(n4189), .A(n4188), .ZN(n5573) );
  NAND2_X1 U5150 ( .A1(n4192), .A2(n4191), .ZN(n4212) );
  AOI22_X1 U5151 ( .A1(n4264), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n3026), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4196) );
  AOI22_X1 U5152 ( .A1(n3031), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4195) );
  AOI22_X1 U5153 ( .A1(n4155), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4194) );
  AOI22_X1 U5154 ( .A1(n4085), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4193) );
  NAND4_X1 U5155 ( .A1(n4196), .A2(n4195), .A3(n4194), .A4(n4193), .ZN(n4202)
         );
  AOI22_X1 U5156 ( .A1(n4097), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4238), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4200) );
  AOI22_X1 U5157 ( .A1(n4214), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4199) );
  AOI22_X1 U5158 ( .A1(n4258), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4198) );
  AOI22_X1 U5159 ( .A1(n4233), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4197) );
  NAND4_X1 U5160 ( .A1(n4200), .A2(n4199), .A3(n4198), .A4(n4197), .ZN(n4201)
         );
  NOR2_X1 U5161 ( .A1(n4202), .A2(n4201), .ZN(n4213) );
  XNOR2_X1 U5162 ( .A(n4212), .B(n4213), .ZN(n4206) );
  NAND2_X1 U5163 ( .A1(n6342), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4203)
         );
  NAND2_X1 U5164 ( .A1(n4275), .A2(n4203), .ZN(n4204) );
  AOI21_X1 U5165 ( .B1(n4277), .B2(EAX_REG_27__SCAN_IN), .A(n4204), .ZN(n4205)
         );
  OAI21_X1 U5166 ( .B1(n4206), .B2(n4249), .A(n4205), .ZN(n4211) );
  INV_X1 U5167 ( .A(n4207), .ZN(n4208) );
  OAI21_X1 U5168 ( .B1(n4209), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n4251), 
        .ZN(n5764) );
  OR2_X1 U5169 ( .A1(n5764), .A2(n4275), .ZN(n4210) );
  NAND2_X1 U5170 ( .A1(n4211), .A2(n4210), .ZN(n5567) );
  NOR2_X1 U5171 ( .A1(n4213), .A2(n4212), .ZN(n4232) );
  AOI22_X1 U5172 ( .A1(n4085), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4218) );
  AOI22_X1 U5173 ( .A1(n3031), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4217) );
  AOI22_X1 U5174 ( .A1(n4155), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4216) );
  AOI22_X1 U5175 ( .A1(n4214), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4215) );
  NAND4_X1 U5176 ( .A1(n4218), .A2(n4217), .A3(n4216), .A4(n4215), .ZN(n4224)
         );
  AOI22_X1 U5177 ( .A1(n4233), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4222) );
  AOI22_X1 U5178 ( .A1(n4097), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4221) );
  AOI22_X1 U5179 ( .A1(n3194), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3169), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n4220) );
  AOI22_X1 U5180 ( .A1(n4238), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4219) );
  NAND4_X1 U5181 ( .A1(n4222), .A2(n4221), .A3(n4220), .A4(n4219), .ZN(n4223)
         );
  OR2_X1 U5182 ( .A1(n4224), .A2(n4223), .ZN(n4231) );
  XNOR2_X1 U5183 ( .A(n4232), .B(n4231), .ZN(n4227) );
  INV_X1 U5184 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5747) );
  OAI21_X1 U5185 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n5747), .A(n4275), .ZN(
        n4225) );
  AOI21_X1 U5186 ( .B1(n4277), .B2(EAX_REG_28__SCAN_IN), .A(n4225), .ZN(n4226)
         );
  OAI21_X1 U5187 ( .B1(n4227), .B2(n4249), .A(n4226), .ZN(n4229) );
  XNOR2_X1 U5188 ( .A(n4251), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5751)
         );
  NAND2_X1 U5189 ( .A1(n5751), .A2(n4278), .ZN(n4228) );
  NAND2_X1 U5190 ( .A1(n4229), .A2(n4228), .ZN(n5558) );
  NAND2_X1 U5191 ( .A1(n4232), .A2(n4231), .ZN(n4256) );
  AOI22_X1 U5192 ( .A1(n4233), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3026), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4237) );
  AOI22_X1 U5193 ( .A1(n4214), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4236) );
  AOI22_X1 U5194 ( .A1(n4097), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3000), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n4235) );
  AOI22_X1 U5195 ( .A1(n4085), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n4177), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4234) );
  NAND4_X1 U5196 ( .A1(n4237), .A2(n4236), .A3(n4235), .A4(n4234), .ZN(n4245)
         );
  AOI22_X1 U5197 ( .A1(n3031), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4243) );
  AOI22_X1 U5198 ( .A1(n4155), .A2(INSTQUEUE_REG_15__6__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4242) );
  AOI22_X1 U5199 ( .A1(n4238), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3036), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4241) );
  AOI22_X1 U5200 ( .A1(n4264), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4240) );
  NAND4_X1 U5201 ( .A1(n4243), .A2(n4242), .A3(n4241), .A4(n4240), .ZN(n4244)
         );
  NOR2_X1 U5202 ( .A1(n4245), .A2(n4244), .ZN(n4257) );
  XNOR2_X1 U5203 ( .A(n4256), .B(n4257), .ZN(n4250) );
  NAND2_X1 U5204 ( .A1(n6342), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4246)
         );
  NAND2_X1 U5205 ( .A1(n4275), .A2(n4246), .ZN(n4247) );
  AOI21_X1 U5206 ( .B1(n4277), .B2(EAX_REG_29__SCAN_IN), .A(n4247), .ZN(n4248)
         );
  OAI21_X1 U5207 ( .B1(n4250), .B2(n4249), .A(n4248), .ZN(n4255) );
  NAND2_X1 U5208 ( .A1(n4252), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4291)
         );
  OR2_X1 U5209 ( .A1(n4252), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4253)
         );
  NAND2_X1 U5210 ( .A1(n4291), .A2(n4253), .ZN(n5739) );
  OR2_X1 U5211 ( .A1(n5739), .A2(n4275), .ZN(n4254) );
  NAND2_X1 U5212 ( .A1(n4255), .A2(n4254), .ZN(n5437) );
  NOR2_X1 U5213 ( .A1(n4257), .A2(n4256), .ZN(n4272) );
  AOI22_X1 U5214 ( .A1(n4238), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4258), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4263) );
  AOI22_X1 U5215 ( .A1(n4214), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4259), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4262) );
  AOI22_X1 U5216 ( .A1(n3000), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3169), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4261) );
  AOI22_X1 U5217 ( .A1(n4177), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3033), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4260) );
  NAND4_X1 U5218 ( .A1(n4263), .A2(n4262), .A3(n4261), .A4(n4260), .ZN(n4270)
         );
  AOI22_X1 U5219 ( .A1(n4233), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n4097), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n4268) );
  AOI22_X1 U5220 ( .A1(n4085), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .B1(n4264), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4267) );
  AOI22_X1 U5221 ( .A1(n3031), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4155), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4266) );
  AOI22_X1 U5222 ( .A1(n3026), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4239), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4265) );
  NAND4_X1 U5223 ( .A1(n4268), .A2(n4267), .A3(n4266), .A4(n4265), .ZN(n4269)
         );
  NOR2_X1 U5224 ( .A1(n4270), .A2(n4269), .ZN(n4271) );
  XNOR2_X1 U5225 ( .A(n4272), .B(n4271), .ZN(n4274) );
  NAND2_X1 U5226 ( .A1(n4274), .A2(n4273), .ZN(n4281) );
  INV_X1 U5227 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n6597) );
  OAI21_X1 U5228 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6597), .A(n4275), .ZN(
        n4276) );
  AOI21_X1 U5229 ( .B1(n4277), .B2(EAX_REG_30__SCAN_IN), .A(n4276), .ZN(n4280)
         );
  XNOR2_X1 U5230 ( .A(n4291), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5730)
         );
  AND2_X1 U5231 ( .A1(n5730), .A2(n4278), .ZN(n4279) );
  AOI21_X1 U5232 ( .B1(n4281), .B2(n4280), .A(n4279), .ZN(n5496) );
  AOI22_X1 U5233 ( .A1(n3790), .A2(EAX_REG_31__SCAN_IN), .B1(n4282), .B2(
        PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4283) );
  XNOR2_X2 U5234 ( .A(n4285), .B(n4284), .ZN(n5522) );
  NAND3_X1 U5235 ( .A1(n6596), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6458) );
  INV_X1 U5236 ( .A(n6458), .ZN(n4286) );
  NAND2_X1 U5237 ( .A1(n4286), .A2(n6354), .ZN(n5642) );
  INV_X1 U5238 ( .A(n5642), .ZN(n6347) );
  INV_X1 U5239 ( .A(n6354), .ZN(n6344) );
  NAND2_X1 U5240 ( .A1(n6344), .A2(n4287), .ZN(n6567) );
  NAND2_X1 U5241 ( .A1(n6567), .A2(n6596), .ZN(n4288) );
  NAND2_X1 U5242 ( .A1(n6596), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4290) );
  NAND2_X1 U5243 ( .A1(n5925), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4289) );
  NAND2_X1 U5244 ( .A1(n4290), .A2(n4289), .ZN(n6146) );
  INV_X1 U5245 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n5533) );
  XNOR2_X1 U5246 ( .A(n4292), .B(n5533), .ZN(n4962) );
  INV_X2 U5247 ( .A(n5908), .ZN(n6582) );
  NAND2_X1 U5248 ( .A1(n6582), .A2(REIP_REG_31__SCAN_IN), .ZN(n5470) );
  NAND2_X1 U5249 ( .A1(n6134), .A2(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4293)
         );
  OAI211_X1 U5250 ( .C1(n6143), .C2(n4962), .A(n5470), .B(n4293), .ZN(n4294)
         );
  AOI21_X1 U5251 ( .B1(n5522), .B2(n6347), .A(n4294), .ZN(n4295) );
  OAI21_X1 U5252 ( .B1(n5474), .B2(n5926), .A(n4295), .ZN(U2955) );
  OAI21_X1 U5253 ( .B1(n4298), .B2(n4297), .A(n4296), .ZN(n5212) );
  NOR2_X1 U5254 ( .A1(n5212), .A2(n6589), .ZN(n4308) );
  INV_X1 U5255 ( .A(n6155), .ZN(n5347) );
  NOR2_X1 U5256 ( .A1(n5347), .A2(n6770), .ZN(n4303) );
  NAND2_X1 U5257 ( .A1(n4300), .A2(n4299), .ZN(n5886) );
  AOI21_X1 U5258 ( .B1(n6770), .B2(n5886), .A(n5266), .ZN(n4301) );
  INV_X1 U5259 ( .A(n4301), .ZN(n4302) );
  MUX2_X1 U5260 ( .A(n4303), .B(n4302), .S(INSTADDRPOINTER_REG_12__SCAN_IN), 
        .Z(n4307) );
  NOR2_X1 U5261 ( .A1(n5158), .A2(n4304), .ZN(n4305) );
  OR2_X1 U5262 ( .A1(n5202), .A2(n4305), .ZN(n5184) );
  NAND2_X1 U5263 ( .A1(n6582), .A2(REIP_REG_12__SCAN_IN), .ZN(n5205) );
  OAI21_X1 U5264 ( .B1(n6584), .B2(n5184), .A(n5205), .ZN(n4306) );
  OR3_X1 U5265 ( .A1(n4308), .A2(n4307), .A3(n4306), .ZN(U3006) );
  AND2_X1 U5266 ( .A1(n6354), .A2(n6548), .ZN(n4984) );
  INV_X1 U5267 ( .A(n4984), .ZN(n4309) );
  NAND2_X1 U5268 ( .A1(n4315), .A2(n4309), .ZN(n5726) );
  NOR2_X1 U5269 ( .A1(n5726), .A2(READREQUEST_REG_SCAN_IN), .ZN(n4312) );
  INV_X1 U5270 ( .A(n4310), .ZN(n5515) );
  NAND2_X1 U5271 ( .A1(n4311), .A2(n5515), .ZN(n5516) );
  AND2_X1 U5272 ( .A1(n4312), .A2(n5727), .ZN(n4313) );
  NAND2_X1 U5273 ( .A1(n6571), .A2(n4952), .ZN(n5521) );
  OAI22_X1 U5274 ( .A1(n4313), .A2(n5521), .B1(n4312), .B2(n6566), .ZN(U3474)
         );
  INV_X1 U5275 ( .A(DATAI_2_), .ZN(n4317) );
  OR3_X2 U5276 ( .A1(n4386), .A2(READY_N), .A3(n4325), .ZN(n6133) );
  INV_X1 U5277 ( .A(UWORD_REG_2__SCAN_IN), .ZN(n4316) );
  INV_X1 U5278 ( .A(n4315), .ZN(n4314) );
  OAI21_X2 U5279 ( .B1(n6436), .B2(n6568), .A(n4314), .ZN(n6130) );
  INV_X1 U5280 ( .A(EAX_REG_18__SCAN_IN), .ZN(n4568) );
  OAI222_X1 U5281 ( .A1(n4317), .A2(n6133), .B1(n4316), .B2(n4690), .C1(n6105), 
        .C2(n4568), .ZN(U2926) );
  INV_X1 U5282 ( .A(DATAI_1_), .ZN(n4319) );
  INV_X1 U5283 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n4318) );
  INV_X1 U5284 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4570) );
  OAI222_X1 U5285 ( .A1(n4319), .A2(n6133), .B1(n4318), .B2(n4690), .C1(n6105), 
        .C2(n4570), .ZN(U2925) );
  INV_X1 U5286 ( .A(DATAI_3_), .ZN(n4321) );
  INV_X1 U5287 ( .A(UWORD_REG_3__SCAN_IN), .ZN(n4320) );
  INV_X1 U5288 ( .A(EAX_REG_19__SCAN_IN), .ZN(n4566) );
  OAI222_X1 U5289 ( .A1(n4321), .A2(n6133), .B1(n4320), .B2(n4690), .C1(n4566), 
        .C2(n6105), .ZN(U2927) );
  INV_X1 U5290 ( .A(DATAI_0_), .ZN(n4323) );
  INV_X1 U5291 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n4322) );
  INV_X1 U5292 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4572) );
  OAI222_X1 U5293 ( .A1(n4323), .A2(n6133), .B1(n4322), .B2(n4690), .C1(n6105), 
        .C2(n4572), .ZN(U2924) );
  INV_X1 U5294 ( .A(n6445), .ZN(n6544) );
  INV_X1 U5295 ( .A(n4324), .ZN(n4535) );
  OR2_X1 U5296 ( .A1(n5520), .A2(n5510), .ZN(n4377) );
  INV_X1 U5297 ( .A(n4325), .ZN(n4328) );
  INV_X1 U5298 ( .A(n6437), .ZN(n4326) );
  AOI21_X1 U5299 ( .B1(n4532), .B2(n4326), .A(n6469), .ZN(n4327) );
  OAI211_X1 U5300 ( .C1(n4328), .C2(n4327), .A(n5520), .B(n6568), .ZN(n4331)
         );
  NAND4_X1 U5301 ( .A1(n4377), .A2(n4331), .A3(n4330), .A4(n4329), .ZN(n4336)
         );
  NAND2_X1 U5302 ( .A1(n5520), .A2(n4332), .ZN(n4335) );
  INV_X1 U5303 ( .A(n3643), .ZN(n5916) );
  NAND2_X1 U5304 ( .A1(n5916), .A2(n4333), .ZN(n4334) );
  NAND2_X1 U5305 ( .A1(n4335), .A2(n4334), .ZN(n4471) );
  INV_X1 U5306 ( .A(n6409), .ZN(n4337) );
  NAND2_X1 U5307 ( .A1(n4337), .A2(n4469), .ZN(n5914) );
  NOR2_X1 U5308 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6761), .ZN(n4413) );
  INV_X1 U5309 ( .A(n4413), .ZN(n6539) );
  INV_X1 U5310 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5927) );
  NOR2_X1 U5311 ( .A1(n6548), .A2(n6342), .ZN(n4558) );
  NAND2_X1 U5312 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4558), .ZN(n6538) );
  OR2_X1 U5313 ( .A1(n5927), .A2(n6538), .ZN(n4338) );
  NAND3_X1 U5314 ( .A1(n5914), .A2(n6539), .A3(n4338), .ZN(n6552) );
  INV_X1 U5315 ( .A(n6552), .ZN(n4371) );
  AOI21_X1 U5316 ( .B1(n6544), .B2(n4535), .A(n4371), .ZN(n4354) );
  INV_X1 U5317 ( .A(n6554), .ZN(n6542) );
  INV_X1 U5318 ( .A(n4340), .ZN(n5723) );
  INV_X1 U5319 ( .A(n3748), .ZN(n4341) );
  NOR2_X1 U5320 ( .A1(n6437), .A2(n4341), .ZN(n4342) );
  NAND2_X1 U5321 ( .A1(n3643), .A2(n4342), .ZN(n4343) );
  NOR2_X1 U5322 ( .A1(n4344), .A2(n4343), .ZN(n6411) );
  NAND2_X1 U5323 ( .A1(n5510), .A2(n4345), .ZN(n4542) );
  XNOR2_X1 U5324 ( .A(n4324), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4348)
         );
  XNOR2_X1 U5325 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4346) );
  OAI22_X1 U5326 ( .A1(n4532), .A2(n4346), .B1(n4534), .B2(n4348), .ZN(n4347)
         );
  AOI21_X1 U5327 ( .B1(n4542), .B2(n4348), .A(n4347), .ZN(n4349) );
  OAI21_X1 U5328 ( .B1(n5723), .B2(n6411), .A(n4349), .ZN(n4545) );
  INV_X1 U5329 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4350) );
  AOI22_X1 U5330 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4350), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n3647), .ZN(n4363) );
  NAND2_X1 U5331 ( .A1(STATE2_REG_1__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4365) );
  NOR2_X1 U5332 ( .A1(n4363), .A2(n4365), .ZN(n4352) );
  NOR3_X1 U5333 ( .A1(n6445), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n4535), 
        .ZN(n4351) );
  AOI211_X1 U5334 ( .C1(n6542), .C2(n4545), .A(n4352), .B(n4351), .ZN(n4353)
         );
  OAI22_X1 U5335 ( .A1(n4354), .A2(n4339), .B1(n4371), .B2(n4353), .ZN(U3459)
         );
  INV_X1 U5336 ( .A(DATAI_15_), .ZN(n4356) );
  INV_X1 U5337 ( .A(EAX_REG_15__SCAN_IN), .ZN(n6072) );
  INV_X1 U5338 ( .A(LWORD_REG_15__SCAN_IN), .ZN(n4355) );
  OAI222_X1 U5339 ( .A1(n4356), .A2(n6133), .B1(n6105), .B2(n6072), .C1(n4355), 
        .C2(n4690), .ZN(U2954) );
  INV_X1 U5340 ( .A(n4357), .ZN(n5097) );
  INV_X1 U5341 ( .A(n6411), .ZN(n4362) );
  INV_X1 U5342 ( .A(n4358), .ZN(n4550) );
  NAND3_X1 U5343 ( .A1(n4359), .A2(n4550), .A3(n4535), .ZN(n4360) );
  OAI21_X1 U5344 ( .B1(n4532), .B2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A(n4360), 
        .ZN(n4361) );
  AOI21_X1 U5345 ( .B1(n5097), .B2(n4362), .A(n4361), .ZN(n6408) );
  INV_X1 U5346 ( .A(n4363), .ZN(n4364) );
  OAI22_X1 U5347 ( .A1(n6408), .A2(n6554), .B1(n4365), .B2(n4364), .ZN(n4366)
         );
  AOI21_X1 U5348 ( .B1(n6544), .B2(n4367), .A(n4366), .ZN(n4370) );
  OAI21_X1 U5349 ( .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6445), .A(n6552), 
        .ZN(n6550) );
  INV_X1 U5350 ( .A(n6550), .ZN(n4368) );
  OAI22_X1 U5351 ( .A1(n4371), .A2(n4370), .B1(n4369), .B2(n4368), .ZN(U3460)
         );
  INV_X1 U5352 ( .A(n4372), .ZN(n4375) );
  NAND4_X1 U5353 ( .A1(n4375), .A2(n4374), .A3(n5598), .A4(n4373), .ZN(n4468)
         );
  OR2_X1 U5354 ( .A1(n4468), .A2(n5426), .ZN(n4376) );
  NAND2_X1 U5355 ( .A1(n4377), .A2(n4376), .ZN(n4378) );
  AND2_X2 U5356 ( .A1(n4378), .A2(n4469), .ZN(n6053) );
  OAI21_X1 U5357 ( .B1(n3011), .B2(n4380), .A(n4379), .ZN(n5103) );
  OR2_X1 U5358 ( .A1(n4382), .A2(n5420), .ZN(n4383) );
  NAND2_X1 U5359 ( .A1(n4384), .A2(n4383), .ZN(n5091) );
  INV_X1 U5360 ( .A(n6053), .ZN(n5590) );
  AOI22_X1 U5361 ( .A1(n6049), .A2(n5091), .B1(EBX_REG_1__SCAN_IN), .B2(n5590), 
        .ZN(n4385) );
  OAI21_X1 U5362 ( .B1(n5589), .B2(n5103), .A(n4385), .ZN(U2858) );
  OR2_X1 U5363 ( .A1(n4386), .A2(n4532), .ZN(n4387) );
  NAND2_X1 U5364 ( .A1(n6596), .A2(n4558), .ZN(n6101) );
  INV_X1 U5365 ( .A(n6101), .ZN(n6095) );
  INV_X1 U5366 ( .A(DATAO_REG_21__SCAN_IN), .ZN(n6751) );
  NAND2_X1 U5367 ( .A1(n6089), .A2(n3271), .ZN(n6067) );
  INV_X1 U5368 ( .A(EAX_REG_21__SCAN_IN), .ZN(n4388) );
  INV_X1 U5369 ( .A(UWORD_REG_5__SCAN_IN), .ZN(n6745) );
  OAI222_X1 U5370 ( .A1(n6104), .A2(n6751), .B1(n6067), .B2(n4388), .C1(n6745), 
        .C2(n6101), .ZN(U2902) );
  INV_X1 U5371 ( .A(n4389), .ZN(n4488) );
  INV_X1 U5372 ( .A(REIP_REG_1__SCAN_IN), .ZN(n5099) );
  NOR2_X1 U5373 ( .A1(n5908), .A2(n5099), .ZN(n4881) );
  NOR3_X1 U5374 ( .A1(n5887), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n4390), 
        .ZN(n4391) );
  AOI211_X1 U5375 ( .C1(n6170), .C2(n5091), .A(n4881), .B(n4391), .ZN(n4396)
         );
  INV_X1 U5376 ( .A(n6589), .ZN(n6186) );
  OR2_X1 U5377 ( .A1(n4394), .A2(n4393), .ZN(n4882) );
  NAND3_X1 U5378 ( .A1(n6186), .A2(n4392), .A3(n4882), .ZN(n4395) );
  OAI211_X1 U5379 ( .C1(n4488), .C2(n3647), .A(n4396), .B(n4395), .ZN(U3017)
         );
  INV_X1 U5380 ( .A(n4460), .ZN(n4398) );
  AOI21_X1 U5381 ( .B1(n4399), .B2(n4480), .A(n4398), .ZN(n4982) );
  INV_X1 U5382 ( .A(n4982), .ZN(n4482) );
  NAND2_X1 U5383 ( .A1(n4464), .A2(n4400), .ZN(n4988) );
  INV_X1 U5384 ( .A(n4988), .ZN(n4401) );
  AOI22_X1 U5385 ( .A1(n6049), .A2(n4401), .B1(EBX_REG_4__SCAN_IN), .B2(n5590), 
        .ZN(n4402) );
  OAI21_X1 U5386 ( .B1(n4482), .B2(n5589), .A(n4402), .ZN(U2855) );
  NAND2_X1 U5387 ( .A1(n5721), .A2(n4403), .ZN(n4414) );
  INV_X1 U5388 ( .A(n4414), .ZN(n6219) );
  AOI21_X1 U5389 ( .B1(n6219), .B2(n3106), .A(n6344), .ZN(n4409) );
  AND2_X1 U5390 ( .A1(n4340), .A2(n4357), .ZN(n5010) );
  INV_X1 U5391 ( .A(n6253), .ZN(n4766) );
  NAND2_X1 U5392 ( .A1(n5010), .A2(n4766), .ZN(n5014) );
  INV_X1 U5393 ( .A(n3789), .ZN(n6412) );
  NAND3_X1 U5394 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6425), .A3(n6415), .ZN(n5012) );
  OR2_X1 U5395 ( .A1(n6769), .A2(n5012), .ZN(n4454) );
  OAI21_X1 U5396 ( .B1(n5014), .B2(n6412), .A(n4454), .ZN(n4405) );
  INV_X1 U5397 ( .A(n5012), .ZN(n4406) );
  AOI22_X1 U5398 ( .A1(n4409), .A2(n4405), .B1(STATE2_REG_2__SCAN_IN), .B2(
        n4406), .ZN(n4458) );
  NAND2_X1 U5399 ( .A1(n6548), .A2(n6342), .ZN(n6446) );
  INV_X1 U5400 ( .A(n6446), .ZN(n6572) );
  NOR2_X1 U5401 ( .A1(n4317), .A2(n4713), .ZN(n6367) );
  INV_X1 U5402 ( .A(n6367), .ZN(n5137) );
  OAI21_X1 U5403 ( .B1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(n6761), .A(n4839), 
        .ZN(n4630) );
  INV_X1 U5404 ( .A(n4405), .ZN(n4408) );
  NOR2_X1 U5405 ( .A1(n6354), .A2(n4406), .ZN(n4407) );
  AOI21_X1 U5406 ( .B1(n4409), .B2(n4408), .A(n4407), .ZN(n4410) );
  NAND2_X1 U5407 ( .A1(n6353), .A2(n4410), .ZN(n4449) );
  NAND2_X1 U5408 ( .A1(n4449), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n4418) );
  INV_X1 U5409 ( .A(DATAI_18_), .ZN(n4411) );
  OR2_X1 U5410 ( .A1(n5642), .A2(n4411), .ZN(n6315) );
  INV_X1 U5411 ( .A(n6315), .ZN(n6368) );
  NOR2_X2 U5412 ( .A1(n4414), .A2(n4733), .ZN(n6248) );
  NAND2_X1 U5413 ( .A1(n4452), .A2(n3203), .ZN(n5022) );
  OR2_X1 U5414 ( .A1(n3035), .A2(n4763), .ZN(n4595) );
  INV_X1 U5415 ( .A(DATAI_26_), .ZN(n4415) );
  OR2_X1 U5416 ( .A1(n5642), .A2(n4415), .ZN(n6371) );
  OAI22_X1 U5417 ( .A1(n5022), .A2(n4454), .B1(n5013), .B2(n6371), .ZN(n4416)
         );
  AOI21_X1 U5418 ( .B1(n6368), .B2(n6248), .A(n4416), .ZN(n4417) );
  OAI211_X1 U5419 ( .C1(n4458), .C2(n5137), .A(n4418), .B(n4417), .ZN(U3062)
         );
  NOR2_X1 U5420 ( .A1(n4323), .A2(n4713), .ZN(n6346) );
  INV_X1 U5421 ( .A(n6346), .ZN(n5119) );
  NAND2_X1 U5422 ( .A1(n4449), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n4423) );
  INV_X1 U5423 ( .A(DATAI_16_), .ZN(n4419) );
  OR2_X1 U5424 ( .A1(n5642), .A2(n4419), .ZN(n6359) );
  INV_X1 U5425 ( .A(n6359), .ZN(n5117) );
  NAND2_X1 U5426 ( .A1(n4452), .A2(n3271), .ZN(n5042) );
  INV_X1 U5427 ( .A(DATAI_24_), .ZN(n4420) );
  OR2_X1 U5428 ( .A1(n5642), .A2(n4420), .ZN(n5115) );
  OAI22_X1 U5429 ( .A1(n5042), .A2(n4454), .B1(n5013), .B2(n5115), .ZN(n4421)
         );
  AOI21_X1 U5430 ( .B1(n5117), .B2(n6248), .A(n4421), .ZN(n4422) );
  OAI211_X1 U5431 ( .C1(n4458), .C2(n5119), .A(n4423), .B(n4422), .ZN(U3060)
         );
  INV_X1 U5432 ( .A(DATAI_7_), .ZN(n6124) );
  NOR2_X1 U5433 ( .A1(n6124), .A2(n4713), .ZN(n6400) );
  INV_X1 U5434 ( .A(n6400), .ZN(n5133) );
  NAND2_X1 U5435 ( .A1(n4449), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4428) );
  INV_X1 U5436 ( .A(DATAI_23_), .ZN(n4424) );
  OR2_X1 U5437 ( .A1(n5642), .A2(n4424), .ZN(n6407) );
  INV_X1 U5438 ( .A(n6407), .ZN(n6330) );
  NAND2_X1 U5439 ( .A1(n4452), .A2(n3275), .ZN(n5030) );
  INV_X1 U5440 ( .A(DATAI_31_), .ZN(n4425) );
  OR2_X1 U5441 ( .A1(n5642), .A2(n4425), .ZN(n6338) );
  OAI22_X1 U5442 ( .A1(n5030), .A2(n4454), .B1(n5013), .B2(n6338), .ZN(n4426)
         );
  AOI21_X1 U5443 ( .B1(n6330), .B2(n6248), .A(n4426), .ZN(n4427) );
  OAI211_X1 U5444 ( .C1(n4458), .C2(n5133), .A(n4428), .B(n4427), .ZN(U3067)
         );
  NOR2_X1 U5445 ( .A1(n4319), .A2(n4713), .ZN(n6361) );
  INV_X1 U5446 ( .A(n6361), .ZN(n5141) );
  NAND2_X1 U5447 ( .A1(n4449), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n4433) );
  INV_X1 U5448 ( .A(DATAI_17_), .ZN(n4429) );
  OR2_X1 U5449 ( .A1(n5642), .A2(n4429), .ZN(n6267) );
  INV_X1 U5450 ( .A(n6267), .ZN(n6362) );
  NAND2_X1 U5451 ( .A1(n4452), .A2(n3259), .ZN(n5046) );
  INV_X1 U5452 ( .A(DATAI_25_), .ZN(n4430) );
  OR2_X1 U5453 ( .A1(n5642), .A2(n4430), .ZN(n6365) );
  OAI22_X1 U5454 ( .A1(n5046), .A2(n4454), .B1(n5013), .B2(n6365), .ZN(n4431)
         );
  AOI21_X1 U5455 ( .B1(n6362), .B2(n6248), .A(n4431), .ZN(n4432) );
  OAI211_X1 U5456 ( .C1(n4458), .C2(n5141), .A(n4433), .B(n4432), .ZN(U3061)
         );
  INV_X1 U5457 ( .A(DATAI_5_), .ZN(n6120) );
  NOR2_X1 U5458 ( .A1(n6120), .A2(n4713), .ZN(n6385) );
  INV_X1 U5459 ( .A(n6385), .ZN(n5152) );
  NAND2_X1 U5460 ( .A1(n4449), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n4438) );
  INV_X1 U5461 ( .A(DATAI_21_), .ZN(n4434) );
  OR2_X1 U5462 ( .A1(n5642), .A2(n4434), .ZN(n6243) );
  INV_X1 U5463 ( .A(n6243), .ZN(n6386) );
  NAND2_X1 U5464 ( .A1(n4452), .A2(n3252), .ZN(n5052) );
  INV_X1 U5465 ( .A(DATAI_29_), .ZN(n4435) );
  OR2_X1 U5466 ( .A1(n5642), .A2(n4435), .ZN(n6390) );
  OAI22_X1 U5467 ( .A1(n5052), .A2(n4454), .B1(n5013), .B2(n6390), .ZN(n4436)
         );
  AOI21_X1 U5468 ( .B1(n6386), .B2(n6248), .A(n4436), .ZN(n4437) );
  OAI211_X1 U5469 ( .C1(n4458), .C2(n5152), .A(n4438), .B(n4437), .ZN(U3065)
         );
  INV_X1 U5470 ( .A(DATAI_4_), .ZN(n6118) );
  NOR2_X1 U5471 ( .A1(n6118), .A2(n4713), .ZN(n6379) );
  INV_X1 U5472 ( .A(n6379), .ZN(n5125) );
  NAND2_X1 U5473 ( .A1(n4449), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n4443) );
  INV_X1 U5474 ( .A(DATAI_20_), .ZN(n4439) );
  OR2_X1 U5475 ( .A1(n5642), .A2(n4439), .ZN(n6383) );
  INV_X1 U5476 ( .A(n6383), .ZN(n5123) );
  NAND2_X1 U5477 ( .A1(n4452), .A2(n3273), .ZN(n5038) );
  INV_X1 U5478 ( .A(DATAI_28_), .ZN(n4440) );
  OR2_X1 U5479 ( .A1(n5642), .A2(n4440), .ZN(n5121) );
  OAI22_X1 U5480 ( .A1(n5038), .A2(n4454), .B1(n5013), .B2(n5121), .ZN(n4441)
         );
  AOI21_X1 U5481 ( .B1(n5123), .B2(n6248), .A(n4441), .ZN(n4442) );
  OAI211_X1 U5482 ( .C1(n4458), .C2(n5125), .A(n4443), .B(n4442), .ZN(U3064)
         );
  NOR2_X1 U5483 ( .A1(n4321), .A2(n4713), .ZN(n6373) );
  INV_X1 U5484 ( .A(n6373), .ZN(n5145) );
  NAND2_X1 U5485 ( .A1(n4449), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n4448) );
  INV_X1 U5486 ( .A(DATAI_19_), .ZN(n4444) );
  OR2_X1 U5487 ( .A1(n5642), .A2(n4444), .ZN(n6377) );
  INV_X1 U5488 ( .A(n6377), .ZN(n6316) );
  NAND2_X1 U5489 ( .A1(n4452), .A2(n3274), .ZN(n5026) );
  INV_X1 U5490 ( .A(DATAI_27_), .ZN(n4445) );
  OR2_X1 U5491 ( .A1(n5642), .A2(n4445), .ZN(n6319) );
  OAI22_X1 U5492 ( .A1(n5026), .A2(n4454), .B1(n5013), .B2(n6319), .ZN(n4446)
         );
  AOI21_X1 U5493 ( .B1(n6316), .B2(n6248), .A(n4446), .ZN(n4447) );
  OAI211_X1 U5494 ( .C1(n4458), .C2(n5145), .A(n4448), .B(n4447), .ZN(U3063)
         );
  INV_X1 U5495 ( .A(DATAI_6_), .ZN(n6122) );
  NOR2_X1 U5496 ( .A1(n6122), .A2(n4713), .ZN(n6392) );
  INV_X1 U5497 ( .A(n6392), .ZN(n5129) );
  NAND2_X1 U5498 ( .A1(n4449), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n4457) );
  INV_X1 U5499 ( .A(DATAI_22_), .ZN(n4450) );
  OR2_X1 U5500 ( .A1(n5642), .A2(n4450), .ZN(n6396) );
  INV_X1 U5501 ( .A(n6396), .ZN(n6326) );
  NAND2_X1 U5502 ( .A1(n4452), .A2(n4451), .ZN(n5034) );
  INV_X1 U5503 ( .A(DATAI_30_), .ZN(n4453) );
  OR2_X1 U5504 ( .A1(n5642), .A2(n4453), .ZN(n6329) );
  OAI22_X1 U5505 ( .A1(n5034), .A2(n4454), .B1(n5013), .B2(n6329), .ZN(n4455)
         );
  AOI21_X1 U5506 ( .B1(n6326), .B2(n6248), .A(n4455), .ZN(n4456) );
  OAI211_X1 U5507 ( .C1(n4458), .C2(n5129), .A(n4457), .B(n4456), .ZN(U3066)
         );
  AND2_X1 U5508 ( .A1(n4460), .A2(n4459), .ZN(n4462) );
  OR2_X1 U5509 ( .A1(n4462), .A2(n4461), .ZN(n4755) );
  INV_X1 U5510 ( .A(n4585), .ZN(n4463) );
  AOI21_X1 U5511 ( .B1(n4465), .B2(n4464), .A(n4463), .ZN(n6014) );
  AOI22_X1 U5512 ( .A1(n6049), .A2(n6014), .B1(EBX_REG_5__SCAN_IN), .B2(n5590), 
        .ZN(n4466) );
  OAI21_X1 U5513 ( .B1(n4755), .B2(n5589), .A(n4466), .ZN(U2854) );
  INV_X1 U5514 ( .A(n5519), .ZN(n4467) );
  NOR2_X1 U5515 ( .A1(n4468), .A2(n4467), .ZN(n4470) );
  OAI21_X1 U5516 ( .B1(n4471), .B2(n4470), .A(n4469), .ZN(n4472) );
  NAND2_X1 U5517 ( .A1(n3260), .A2(n3275), .ZN(n4473) );
  INV_X1 U5518 ( .A(n4473), .ZN(n4474) );
  NAND2_X1 U5519 ( .A1(n5504), .A2(n4474), .ZN(n5306) );
  INV_X1 U5520 ( .A(EAX_REG_1__SCAN_IN), .ZN(n6099) );
  OAI222_X1 U5521 ( .A1(n5103), .A2(n5603), .B1(n5306), .B2(n4319), .C1(n5504), 
        .C2(n6099), .ZN(U2890) );
  NAND2_X1 U5522 ( .A1(n4476), .A2(n4475), .ZN(n4477) );
  NAND2_X1 U5523 ( .A1(n4478), .A2(n4477), .ZN(n6152) );
  INV_X1 U5524 ( .A(EAX_REG_0__SCAN_IN), .ZN(n6102) );
  OAI222_X1 U5525 ( .A1(n6152), .A2(n5603), .B1(n5306), .B2(n4323), .C1(n5504), 
        .C2(n6102), .ZN(U2891) );
  OAI21_X1 U5526 ( .B1(n4479), .B2(n4481), .A(n4480), .ZN(n6039) );
  INV_X1 U5527 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6094) );
  OAI222_X1 U5528 ( .A1(n6039), .A2(n5603), .B1(n5306), .B2(n4321), .C1(n5504), 
        .C2(n6094), .ZN(U2888) );
  INV_X1 U5529 ( .A(EAX_REG_4__SCAN_IN), .ZN(n6092) );
  OAI222_X1 U5530 ( .A1(n4482), .A2(n5603), .B1(n5306), .B2(n6118), .C1(n5504), 
        .C2(n6092), .ZN(U2887) );
  NOR2_X1 U5531 ( .A1(n3001), .A2(n4483), .ZN(n4485) );
  NOR2_X1 U5532 ( .A1(n4479), .A2(n4485), .ZN(n6139) );
  INV_X1 U5533 ( .A(n6139), .ZN(n5007) );
  OAI222_X1 U5534 ( .A1(n5007), .A2(n5603), .B1(n5306), .B2(n4317), .C1(n5504), 
        .C2(n3797), .ZN(U2889) );
  XNOR2_X1 U5535 ( .A(n4487), .B(n4486), .ZN(n4760) );
  NOR2_X1 U5536 ( .A1(n3657), .A2(n3647), .ZN(n4504) );
  OAI22_X1 U5537 ( .A1(n6171), .A2(n4488), .B1(n4931), .B2(n4504), .ZN(n4489)
         );
  INV_X1 U5538 ( .A(n4489), .ZN(n6173) );
  INV_X1 U5539 ( .A(n4617), .ZN(n4490) );
  INV_X1 U5540 ( .A(n5887), .ZN(n5464) );
  OAI21_X1 U5541 ( .B1(n4493), .B2(n4490), .A(n5464), .ZN(n4491) );
  NAND2_X1 U5542 ( .A1(n6173), .A2(n4491), .ZN(n4623) );
  NAND3_X1 U5543 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n6176), .ZN(n4494) );
  OAI211_X1 U5544 ( .C1(n4683), .C2(n4494), .A(n4493), .B(n4492), .ZN(n4495)
         );
  NAND2_X1 U5545 ( .A1(n4623), .A2(n4495), .ZN(n4497) );
  INV_X1 U5546 ( .A(REIP_REG_5__SCAN_IN), .ZN(n6488) );
  NOR2_X1 U5547 ( .A1(n5908), .A2(n6488), .ZN(n4756) );
  AOI21_X1 U5548 ( .B1(n6170), .B2(n6014), .A(n4756), .ZN(n4496) );
  OAI211_X1 U5549 ( .C1(n4760), .C2(n6589), .A(n4497), .B(n4496), .ZN(U3013)
         );
  OAI222_X1 U5550 ( .A1(n4755), .A2(n5603), .B1(n5306), .B2(n6120), .C1(n5504), 
        .C2(n3827), .ZN(U2886) );
  XNOR2_X1 U5551 ( .A(n4499), .B(n4498), .ZN(n4515) );
  INV_X1 U5552 ( .A(n6039), .ZN(n4502) );
  INV_X1 U5553 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6484) );
  NOR2_X1 U5554 ( .A1(n5908), .A2(n6484), .ZN(n4511) );
  AOI21_X1 U5555 ( .B1(n6134), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n4511), 
        .ZN(n4500) );
  OAI21_X1 U5556 ( .B1(n6037), .B2(n6143), .A(n4500), .ZN(n4501) );
  AOI21_X1 U5557 ( .B1(n4502), .B2(n6347), .A(n4501), .ZN(n4503) );
  OAI21_X1 U5558 ( .B1(n4515), .B2(n5926), .A(n4503), .ZN(U2983) );
  NAND2_X1 U5559 ( .A1(n6171), .A2(n4505), .ZN(n6178) );
  NAND2_X1 U5560 ( .A1(n6173), .A2(n6178), .ZN(n4687) );
  AOI21_X1 U5561 ( .B1(n4504), .B2(n6176), .A(n6171), .ZN(n4619) );
  NOR2_X1 U5562 ( .A1(n4505), .A2(n4619), .ZN(n4936) );
  INV_X1 U5563 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4506) );
  AOI22_X1 U5564 ( .A1(INSTADDRPOINTER_REG_3__SCAN_IN), .A2(n4687), .B1(n4936), 
        .B2(n4506), .ZN(n4514) );
  INV_X1 U5565 ( .A(n4507), .ZN(n4509) );
  AOI21_X1 U5566 ( .B1(n4509), .B2(n5000), .A(n4508), .ZN(n4510) );
  INV_X1 U5567 ( .A(n6034), .ZN(n4512) );
  AOI21_X1 U5568 ( .B1(n6170), .B2(n4512), .A(n4511), .ZN(n4513) );
  OAI211_X1 U5569 ( .C1(n4515), .C2(n6589), .A(n4514), .B(n4513), .ZN(U3015)
         );
  XNOR2_X1 U5570 ( .A(n4516), .B(n4517), .ZN(n4689) );
  INV_X1 U5571 ( .A(n4518), .ZN(n4992) );
  AOI22_X1 U5572 ( .A1(n6134), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n6582), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n4519) );
  OAI21_X1 U5573 ( .B1(n4992), .B2(n6143), .A(n4519), .ZN(n4520) );
  AOI21_X1 U5574 ( .B1(n4982), .B2(n6347), .A(n4520), .ZN(n4521) );
  OAI21_X1 U5575 ( .B1(n5926), .B2(n4689), .A(n4521), .ZN(U2982) );
  NAND2_X1 U5576 ( .A1(n6409), .A2(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n4526) );
  NOR2_X1 U5577 ( .A1(n4522), .A2(n4766), .ZN(n4524) );
  XNOR2_X1 U5578 ( .A(n4524), .B(n4523), .ZN(n5915) );
  NAND2_X1 U5579 ( .A1(n5915), .A2(n5916), .ZN(n4525) );
  NAND2_X1 U5580 ( .A1(n4526), .A2(n4525), .ZN(n4529) );
  NAND2_X1 U5581 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5927), .ZN(n4549) );
  INV_X1 U5582 ( .A(n4549), .ZN(n4527) );
  AND2_X1 U5583 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n4527), .ZN(n4528)
         );
  AOI21_X1 U5584 ( .B1(n4529), .B2(n6548), .A(n4528), .ZN(n4546) );
  INV_X1 U5585 ( .A(n4546), .ZN(n4551) );
  INV_X1 U5586 ( .A(n4530), .ZN(n4548) );
  INV_X1 U5587 ( .A(n4532), .ZN(n6413) );
  XNOR2_X1 U5588 ( .A(n3804), .B(n4533), .ZN(n4538) );
  INV_X1 U5589 ( .A(n4534), .ZN(n4537) );
  OAI21_X1 U5590 ( .B1(n4535), .B2(n4339), .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .ZN(n4536) );
  NAND2_X1 U5591 ( .A1(n3414), .A2(n4536), .ZN(n6543) );
  AOI22_X1 U5592 ( .A1(n6413), .A2(n4538), .B1(n4537), .B2(n6543), .ZN(n4544)
         );
  INV_X1 U5593 ( .A(n4539), .ZN(n4540) );
  MUX2_X1 U5594 ( .A(n4540), .B(n3804), .S(n4324), .Z(n4541) );
  NAND3_X1 U5595 ( .A1(n4542), .A2(n4548), .A3(n4541), .ZN(n4543) );
  OAI211_X1 U5596 ( .C1(n6032), .C2(n6411), .A(n4544), .B(n4543), .ZN(n6541)
         );
  MUX2_X1 U5597 ( .A(n6541), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n6409), 
        .Z(n6426) );
  MUX2_X1 U5598 ( .A(n4545), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .S(n6409), 
        .Z(n6420) );
  NAND3_X1 U5599 ( .A1(n6426), .A2(n6420), .A3(n6548), .ZN(n4547) );
  OAI211_X1 U5600 ( .C1(n4549), .C2(n4548), .A(n4547), .B(n4546), .ZN(n6430)
         );
  OAI21_X1 U5601 ( .B1(n4551), .B2(n4550), .A(n6430), .ZN(n4559) );
  AOI21_X1 U5602 ( .B1(n4559), .B2(n5927), .A(n6538), .ZN(n4552) );
  OR2_X1 U5603 ( .A1(n4552), .A2(n4839), .ZN(n6190) );
  AND2_X1 U5604 ( .A1(n4553), .A2(n5721), .ZN(n4894) );
  NAND2_X1 U5605 ( .A1(n4894), .A2(n3106), .ZN(n4730) );
  INV_X1 U5606 ( .A(n4730), .ZN(n4554) );
  INV_X1 U5607 ( .A(n5721), .ZN(n4634) );
  NOR2_X1 U5608 ( .A1(n4554), .A2(n6298), .ZN(n4625) );
  AND2_X1 U5609 ( .A1(n3035), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6297) );
  NAND2_X1 U5610 ( .A1(n6219), .A2(n6297), .ZN(n6258) );
  AOI21_X1 U5611 ( .B1(n4625), .B2(n6258), .A(n6344), .ZN(n4556) );
  NAND2_X1 U5612 ( .A1(n6354), .A2(n5925), .ZN(n4835) );
  AND2_X1 U5613 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6761), .ZN(n5722) );
  OAI22_X1 U5614 ( .A1(n4635), .A2(n4835), .B1(n6032), .B2(n5722), .ZN(n4555)
         );
  OAI21_X1 U5615 ( .B1(n4556), .B2(n4555), .A(n6190), .ZN(n4557) );
  OAI21_X1 U5616 ( .B1(n6190), .B2(n6425), .A(n4557), .ZN(U3462) );
  NAND2_X1 U5617 ( .A1(n4559), .A2(n4558), .ZN(n6448) );
  INV_X1 U5618 ( .A(n6448), .ZN(n4561) );
  OAI21_X1 U5619 ( .B1(n4561), .B2(n4560), .A(n6190), .ZN(n4562) );
  OAI21_X1 U5620 ( .B1(n6190), .B2(n6769), .A(n4562), .ZN(U3465) );
  INV_X1 U5621 ( .A(EAX_REG_24__SCAN_IN), .ZN(n4704) );
  AOI22_X1 U5622 ( .A1(UWORD_REG_8__SCAN_IN), .A2(n6569), .B1(n6097), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4563) );
  OAI21_X1 U5623 ( .B1(n4704), .B2(n6067), .A(n4563), .ZN(U2899) );
  INV_X1 U5624 ( .A(EAX_REG_30__SCAN_IN), .ZN(n4696) );
  AOI22_X1 U5625 ( .A1(n6569), .A2(UWORD_REG_14__SCAN_IN), .B1(n6097), .B2(
        DATAO_REG_30__SCAN_IN), .ZN(n4564) );
  OAI21_X1 U5626 ( .B1(n4696), .B2(n6067), .A(n4564), .ZN(U2893) );
  AOI22_X1 U5627 ( .A1(n6095), .A2(UWORD_REG_3__SCAN_IN), .B1(n6097), .B2(
        DATAO_REG_19__SCAN_IN), .ZN(n4565) );
  OAI21_X1 U5628 ( .B1(n4566), .B2(n6067), .A(n4565), .ZN(U2904) );
  AOI22_X1 U5629 ( .A1(n6095), .A2(UWORD_REG_2__SCAN_IN), .B1(n6097), .B2(
        DATAO_REG_18__SCAN_IN), .ZN(n4567) );
  OAI21_X1 U5630 ( .B1(n4568), .B2(n6067), .A(n4567), .ZN(U2905) );
  AOI22_X1 U5631 ( .A1(n6569), .A2(UWORD_REG_1__SCAN_IN), .B1(n6097), .B2(
        DATAO_REG_17__SCAN_IN), .ZN(n4569) );
  OAI21_X1 U5632 ( .B1(n4570), .B2(n6067), .A(n4569), .ZN(U2906) );
  AOI22_X1 U5633 ( .A1(n6569), .A2(UWORD_REG_0__SCAN_IN), .B1(n6097), .B2(
        DATAO_REG_16__SCAN_IN), .ZN(n4571) );
  OAI21_X1 U5634 ( .B1(n4572), .B2(n6067), .A(n4571), .ZN(U2907) );
  INV_X1 U5635 ( .A(EAX_REG_27__SCAN_IN), .ZN(n4707) );
  AOI22_X1 U5636 ( .A1(n6095), .A2(UWORD_REG_11__SCAN_IN), .B1(n6097), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4573) );
  OAI21_X1 U5637 ( .B1(n4707), .B2(n6067), .A(n4573), .ZN(U2896) );
  INV_X1 U5638 ( .A(EAX_REG_26__SCAN_IN), .ZN(n4701) );
  AOI22_X1 U5639 ( .A1(n6095), .A2(UWORD_REG_10__SCAN_IN), .B1(n6097), .B2(
        DATAO_REG_26__SCAN_IN), .ZN(n4574) );
  OAI21_X1 U5640 ( .B1(n4701), .B2(n6067), .A(n4574), .ZN(U2897) );
  INV_X1 U5641 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4576) );
  AOI22_X1 U5642 ( .A1(n6095), .A2(UWORD_REG_9__SCAN_IN), .B1(n6097), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4575) );
  OAI21_X1 U5643 ( .B1(n4576), .B2(n6067), .A(n4575), .ZN(U2898) );
  INV_X1 U5644 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4578) );
  AOI22_X1 U5645 ( .A1(n6095), .A2(UWORD_REG_6__SCAN_IN), .B1(n6097), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4577) );
  OAI21_X1 U5646 ( .B1(n4578), .B2(n6067), .A(n4577), .ZN(U2901) );
  INV_X1 U5647 ( .A(EAX_REG_29__SCAN_IN), .ZN(n4580) );
  AOI22_X1 U5648 ( .A1(n6095), .A2(UWORD_REG_13__SCAN_IN), .B1(n6097), .B2(
        DATAO_REG_29__SCAN_IN), .ZN(n4579) );
  OAI21_X1 U5649 ( .B1(n4580), .B2(n6067), .A(n4579), .ZN(U2894) );
  OR2_X1 U5650 ( .A1(n4461), .A2(n4582), .ZN(n4583) );
  NAND2_X1 U5651 ( .A1(n4581), .A2(n4583), .ZN(n6005) );
  NAND2_X1 U5652 ( .A1(n4585), .A2(n4584), .ZN(n4586) );
  AND2_X1 U5653 ( .A1(n4876), .A2(n4586), .ZN(n6000) );
  AOI22_X1 U5654 ( .A1(n6049), .A2(n6000), .B1(EBX_REG_6__SCAN_IN), .B2(n5590), 
        .ZN(n4587) );
  OAI21_X1 U5655 ( .B1(n6005), .B2(n5589), .A(n4587), .ZN(U2853) );
  INV_X1 U5656 ( .A(EAX_REG_23__SCAN_IN), .ZN(n4589) );
  AOI22_X1 U5657 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n6095), .B1(
        DATAO_REG_23__SCAN_IN), .B2(n6097), .ZN(n4588) );
  OAI21_X1 U5658 ( .B1(n4589), .B2(n6067), .A(n4588), .ZN(U2900) );
  INV_X1 U5659 ( .A(n6298), .ZN(n4590) );
  NOR2_X1 U5660 ( .A1(n6032), .A2(n6412), .ZN(n6341) );
  NOR2_X1 U5661 ( .A1(n4340), .A2(n5097), .ZN(n4802) );
  NAND3_X1 U5662 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6421), .A3(n6415), .ZN(n4799) );
  NOR2_X1 U5663 ( .A1(n6769), .A2(n4799), .ZN(n4612) );
  AOI21_X1 U5664 ( .B1(n6341), .B2(n4802), .A(n4612), .ZN(n4594) );
  AOI21_X1 U5665 ( .B1(n6298), .B2(n3106), .A(n6344), .ZN(n4592) );
  AOI22_X1 U5666 ( .A1(n4594), .A2(n4592), .B1(n6344), .B2(n4799), .ZN(n4591)
         );
  NAND2_X1 U5667 ( .A1(n6353), .A2(n4591), .ZN(n4611) );
  INV_X1 U5668 ( .A(n4592), .ZN(n4593) );
  OAI22_X1 U5669 ( .A1(n4594), .A2(n4593), .B1(n6342), .B2(n4799), .ZN(n4610)
         );
  AOI22_X1 U5670 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n4611), .B1(n6346), 
        .B2(n4610), .ZN(n4597) );
  INV_X1 U5671 ( .A(n5115), .ZN(n6356) );
  INV_X1 U5672 ( .A(n4595), .ZN(n4727) );
  AOI22_X1 U5673 ( .A1(n6345), .A2(n4612), .B1(n6356), .B2(n6291), .ZN(n4596)
         );
  OAI211_X1 U5674 ( .C1(n6359), .C2(n5149), .A(n4597), .B(n4596), .ZN(U3092)
         );
  AOI22_X1 U5675 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n4611), .B1(n6367), 
        .B2(n4610), .ZN(n4599) );
  INV_X1 U5676 ( .A(n6371), .ZN(n6312) );
  AOI22_X1 U5677 ( .A1(n6366), .A2(n4612), .B1(n6312), .B2(n6291), .ZN(n4598)
         );
  OAI211_X1 U5678 ( .C1(n6315), .C2(n5149), .A(n4599), .B(n4598), .ZN(U3094)
         );
  AOI22_X1 U5679 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n4611), .B1(n6373), 
        .B2(n4610), .ZN(n4601) );
  INV_X1 U5680 ( .A(n6319), .ZN(n6374) );
  AOI22_X1 U5681 ( .A1(n6372), .A2(n4612), .B1(n6374), .B2(n6291), .ZN(n4600)
         );
  OAI211_X1 U5682 ( .C1(n6377), .C2(n5149), .A(n4601), .B(n4600), .ZN(U3095)
         );
  AOI22_X1 U5683 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n4611), .B1(n6361), 
        .B2(n4610), .ZN(n4603) );
  INV_X1 U5684 ( .A(n6365), .ZN(n6264) );
  AOI22_X1 U5685 ( .A1(n6360), .A2(n4612), .B1(n6264), .B2(n6291), .ZN(n4602)
         );
  OAI211_X1 U5686 ( .C1(n6267), .C2(n5149), .A(n4603), .B(n4602), .ZN(U3093)
         );
  AOI22_X1 U5687 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n4611), .B1(n6400), 
        .B2(n4610), .ZN(n4605) );
  INV_X1 U5688 ( .A(n6338), .ZN(n6402) );
  AOI22_X1 U5689 ( .A1(n6397), .A2(n4612), .B1(n6402), .B2(n6291), .ZN(n4604)
         );
  OAI211_X1 U5690 ( .C1(n6407), .C2(n5149), .A(n4605), .B(n4604), .ZN(U3099)
         );
  AOI22_X1 U5691 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n4611), .B1(n6392), 
        .B2(n4610), .ZN(n4607) );
  INV_X1 U5692 ( .A(n6329), .ZN(n6393) );
  AOI22_X1 U5693 ( .A1(n6391), .A2(n4612), .B1(n6393), .B2(n6291), .ZN(n4606)
         );
  OAI211_X1 U5694 ( .C1(n6396), .C2(n5149), .A(n4607), .B(n4606), .ZN(U3098)
         );
  AOI22_X1 U5695 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n4611), .B1(n6385), 
        .B2(n4610), .ZN(n4609) );
  INV_X1 U5696 ( .A(n6390), .ZN(n6240) );
  AOI22_X1 U5697 ( .A1(n6384), .A2(n4612), .B1(n6240), .B2(n6291), .ZN(n4608)
         );
  OAI211_X1 U5698 ( .C1(n6243), .C2(n5149), .A(n4609), .B(n4608), .ZN(U3097)
         );
  AOI22_X1 U5699 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4611), .B1(n6379), 
        .B2(n4610), .ZN(n4614) );
  INV_X1 U5700 ( .A(n5121), .ZN(n6380) );
  AOI22_X1 U5701 ( .A1(n6378), .A2(n4612), .B1(n6380), .B2(n6291), .ZN(n4613)
         );
  OAI211_X1 U5702 ( .C1(n6383), .C2(n5149), .A(n4614), .B(n4613), .ZN(U3096)
         );
  XNOR2_X1 U5703 ( .A(n4615), .B(n4616), .ZN(n4832) );
  NAND2_X1 U5704 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4617), .ZN(n4618)
         );
  NOR3_X1 U5705 ( .A1(INSTADDRPOINTER_REG_6__SCAN_IN), .A2(n4619), .A3(n4618), 
        .ZN(n4622) );
  INV_X1 U5706 ( .A(n6000), .ZN(n4620) );
  INV_X1 U5707 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6490) );
  OAI22_X1 U5708 ( .A1(n6584), .A2(n4620), .B1(n6490), .B2(n5908), .ZN(n4621)
         );
  AOI211_X1 U5709 ( .C1(n4623), .C2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n4622), 
        .B(n4621), .ZN(n4624) );
  OAI21_X1 U5710 ( .B1(n6589), .B2(n4832), .A(n4624), .ZN(U3012) );
  NAND3_X1 U5711 ( .A1(n4625), .A2(n6297), .A3(n4634), .ZN(n4626) );
  NAND2_X1 U5712 ( .A1(n4626), .A2(n6354), .ZN(n4633) );
  NOR2_X1 U5713 ( .A1(n4340), .A2(n4357), .ZN(n5105) );
  NAND2_X1 U5714 ( .A1(n5105), .A2(n6032), .ZN(n4836) );
  OR2_X1 U5715 ( .A1(n4836), .A2(n6412), .ZN(n4628) );
  INV_X1 U5716 ( .A(n6296), .ZN(n4627) );
  NAND2_X1 U5717 ( .A1(n4627), .A2(n6425), .ZN(n6206) );
  AND2_X1 U5718 ( .A1(n4628), .A2(n6206), .ZN(n4629) );
  NAND2_X1 U5719 ( .A1(n5108), .A2(n6425), .ZN(n4838) );
  OAI22_X1 U5720 ( .A1(n4633), .A2(n4629), .B1(n4838), .B2(n6342), .ZN(n6213)
         );
  INV_X1 U5721 ( .A(n6213), .ZN(n4651) );
  INV_X1 U5722 ( .A(n4629), .ZN(n4632) );
  AOI21_X1 U5723 ( .B1(n6344), .B2(n4838), .A(n4630), .ZN(n4631) );
  OAI21_X1 U5724 ( .B1(n4633), .B2(n4632), .A(n4631), .ZN(n6214) );
  NOR2_X1 U5725 ( .A1(n3803), .A2(n5721), .ZN(n4654) );
  AND2_X1 U5726 ( .A1(n4654), .A2(n6218), .ZN(n6211) );
  NOR2_X1 U5727 ( .A1(n4865), .A2(n6390), .ZN(n4637) );
  NAND4_X1 U5728 ( .A1(n4635), .A2(n4763), .A3(n4634), .A4(n3035), .ZN(n6217)
         );
  OAI22_X1 U5729 ( .A1(n5052), .A2(n6206), .B1(n6243), .B2(n6217), .ZN(n4636)
         );
  AOI211_X1 U5730 ( .C1(n6214), .C2(INSTQUEUE_REG_3__5__SCAN_IN), .A(n4637), 
        .B(n4636), .ZN(n4638) );
  OAI21_X1 U5731 ( .B1(n4651), .B2(n5152), .A(n4638), .ZN(U3049) );
  NOR2_X1 U5732 ( .A1(n4865), .A2(n6371), .ZN(n4640) );
  OAI22_X1 U5733 ( .A1(n5022), .A2(n6206), .B1(n6315), .B2(n6217), .ZN(n4639)
         );
  AOI211_X1 U5734 ( .C1(n6214), .C2(INSTQUEUE_REG_3__2__SCAN_IN), .A(n4640), 
        .B(n4639), .ZN(n4641) );
  OAI21_X1 U5735 ( .B1(n4651), .B2(n5137), .A(n4641), .ZN(U3046) );
  NOR2_X1 U5736 ( .A1(n4865), .A2(n6365), .ZN(n4643) );
  OAI22_X1 U5737 ( .A1(n5046), .A2(n6206), .B1(n6267), .B2(n6217), .ZN(n4642)
         );
  AOI211_X1 U5738 ( .C1(n6214), .C2(INSTQUEUE_REG_3__1__SCAN_IN), .A(n4643), 
        .B(n4642), .ZN(n4644) );
  OAI21_X1 U5739 ( .B1(n4651), .B2(n5141), .A(n4644), .ZN(U3045) );
  NOR2_X1 U5740 ( .A1(n4865), .A2(n6319), .ZN(n4646) );
  OAI22_X1 U5741 ( .A1(n5026), .A2(n6206), .B1(n6377), .B2(n6217), .ZN(n4645)
         );
  AOI211_X1 U5742 ( .C1(n6214), .C2(INSTQUEUE_REG_3__3__SCAN_IN), .A(n4646), 
        .B(n4645), .ZN(n4647) );
  OAI21_X1 U5743 ( .B1(n4651), .B2(n5145), .A(n4647), .ZN(U3047) );
  NOR2_X1 U5744 ( .A1(n4865), .A2(n6338), .ZN(n4649) );
  OAI22_X1 U5745 ( .A1(n5030), .A2(n6206), .B1(n6407), .B2(n6217), .ZN(n4648)
         );
  AOI211_X1 U5746 ( .C1(n6214), .C2(INSTQUEUE_REG_3__7__SCAN_IN), .A(n4649), 
        .B(n4648), .ZN(n4650) );
  OAI21_X1 U5747 ( .B1(n4651), .B2(n5133), .A(n4650), .ZN(U3051) );
  INV_X1 U5748 ( .A(EBX_REG_3__SCAN_IN), .ZN(n4652) );
  OAI222_X1 U5749 ( .A1(n6039), .A2(n5589), .B1(n4652), .B2(n6053), .C1(n5597), 
        .C2(n6034), .ZN(U2856) );
  INV_X1 U5750 ( .A(n3035), .ZN(n4653) );
  NAND2_X1 U5751 ( .A1(n4654), .A2(n4653), .ZN(n4661) );
  INV_X1 U5752 ( .A(n4661), .ZN(n4655) );
  NAND2_X1 U5753 ( .A1(n4655), .A2(n4763), .ZN(n4834) );
  INV_X1 U5754 ( .A(n4802), .ZN(n4801) );
  NOR2_X1 U5755 ( .A1(n4801), .A2(n4531), .ZN(n4709) );
  NAND3_X1 U5756 ( .A1(n6425), .A2(n6421), .A3(n6415), .ZN(n4711) );
  NOR2_X1 U5757 ( .A1(n6769), .A2(n4711), .ZN(n4678) );
  AOI21_X1 U5758 ( .B1(n4709), .B2(n3789), .A(n4678), .ZN(n4659) );
  OR2_X1 U5759 ( .A1(n4661), .A2(n5925), .ZN(n4656) );
  AND2_X1 U5760 ( .A1(n4656), .A2(n6354), .ZN(n4658) );
  AOI22_X1 U5761 ( .A1(n4659), .A2(n4658), .B1(n6344), .B2(n4711), .ZN(n4657)
         );
  NAND2_X1 U5762 ( .A1(n6353), .A2(n4657), .ZN(n4677) );
  INV_X1 U5763 ( .A(n4658), .ZN(n4660) );
  OAI22_X1 U5764 ( .A1(n4660), .A2(n4659), .B1(n6342), .B2(n4711), .ZN(n4676)
         );
  AOI22_X1 U5765 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n4677), .B1(n6367), 
        .B2(n4676), .ZN(n4663) );
  NOR2_X2 U5766 ( .A1(n4661), .A2(n4763), .ZN(n6202) );
  AOI22_X1 U5767 ( .A1(n6312), .A2(n6202), .B1(n6366), .B2(n4678), .ZN(n4662)
         );
  OAI211_X1 U5768 ( .C1(n6315), .C2(n4834), .A(n4663), .B(n4662), .ZN(U3030)
         );
  AOI22_X1 U5769 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n4677), .B1(n6385), 
        .B2(n4676), .ZN(n4665) );
  AOI22_X1 U5770 ( .A1(n6240), .A2(n6202), .B1(n6384), .B2(n4678), .ZN(n4664)
         );
  OAI211_X1 U5771 ( .C1(n6243), .C2(n4834), .A(n4665), .B(n4664), .ZN(U3033)
         );
  AOI22_X1 U5772 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n4677), .B1(n6346), 
        .B2(n4676), .ZN(n4667) );
  AOI22_X1 U5773 ( .A1(n6356), .A2(n6202), .B1(n6345), .B2(n4678), .ZN(n4666)
         );
  OAI211_X1 U5774 ( .C1(n6359), .C2(n4834), .A(n4667), .B(n4666), .ZN(U3028)
         );
  AOI22_X1 U5775 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n4677), .B1(n6373), 
        .B2(n4676), .ZN(n4669) );
  AOI22_X1 U5776 ( .A1(n6374), .A2(n6202), .B1(n6372), .B2(n4678), .ZN(n4668)
         );
  OAI211_X1 U5777 ( .C1(n6377), .C2(n4834), .A(n4669), .B(n4668), .ZN(U3031)
         );
  AOI22_X1 U5778 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n4677), .B1(n6392), 
        .B2(n4676), .ZN(n4671) );
  AOI22_X1 U5779 ( .A1(n6393), .A2(n6202), .B1(n6391), .B2(n4678), .ZN(n4670)
         );
  OAI211_X1 U5780 ( .C1(n6396), .C2(n4834), .A(n4671), .B(n4670), .ZN(U3034)
         );
  AOI22_X1 U5781 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n4677), .B1(n6361), 
        .B2(n4676), .ZN(n4673) );
  AOI22_X1 U5782 ( .A1(n6264), .A2(n6202), .B1(n6360), .B2(n4678), .ZN(n4672)
         );
  OAI211_X1 U5783 ( .C1(n6267), .C2(n4834), .A(n4673), .B(n4672), .ZN(U3029)
         );
  AOI22_X1 U5784 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4677), .B1(n6379), 
        .B2(n4676), .ZN(n4675) );
  AOI22_X1 U5785 ( .A1(n6380), .A2(n6202), .B1(n6378), .B2(n4678), .ZN(n4674)
         );
  OAI211_X1 U5786 ( .C1(n6383), .C2(n4834), .A(n4675), .B(n4674), .ZN(U3032)
         );
  AOI22_X1 U5787 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n4677), .B1(n6400), 
        .B2(n4676), .ZN(n4680) );
  AOI22_X1 U5788 ( .A1(n6402), .A2(n6202), .B1(n6397), .B2(n4678), .ZN(n4679)
         );
  OAI211_X1 U5789 ( .C1(n6407), .C2(n4834), .A(n4680), .B(n4679), .ZN(U3035)
         );
  INV_X1 U5790 ( .A(EAX_REG_6__SCAN_IN), .ZN(n6730) );
  OAI222_X1 U5791 ( .A1(n6005), .A2(n5603), .B1(n5306), .B2(n6122), .C1(n5504), 
        .C2(n6730), .ZN(U2885) );
  OR2_X1 U5792 ( .A1(n5427), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4682)
         );
  NAND2_X1 U5793 ( .A1(n4682), .A2(n4681), .ZN(n6183) );
  OAI222_X1 U5794 ( .A1(n6183), .A2(n5597), .B1(n4959), .B2(n6053), .C1(n6152), 
        .C2(n5589), .ZN(U2859) );
  INV_X1 U5795 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6486) );
  OAI22_X1 U5796 ( .A1(n6584), .A2(n4988), .B1(n6486), .B2(n5908), .ZN(n4686)
         );
  OAI211_X1 U5797 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_3__SCAN_IN), .A(n4936), .B(n4683), .ZN(n4684) );
  INV_X1 U5798 ( .A(n4684), .ZN(n4685) );
  AOI211_X1 U5799 ( .C1(INSTADDRPOINTER_REG_4__SCAN_IN), .C2(n4687), .A(n4686), 
        .B(n4685), .ZN(n4688) );
  OAI21_X1 U5800 ( .B1(n6589), .B2(n4689), .A(n4688), .ZN(U3014) );
  INV_X1 U5801 ( .A(EAX_REG_8__SCAN_IN), .ZN(n6085) );
  NAND2_X1 U5802 ( .A1(n6125), .A2(LWORD_REG_8__SCAN_IN), .ZN(n4691) );
  INV_X1 U5803 ( .A(n6133), .ZN(n4694) );
  NAND2_X1 U5804 ( .A1(n4694), .A2(DATAI_8_), .ZN(n4702) );
  OAI211_X1 U5805 ( .C1(n6085), .C2(n6105), .A(n4691), .B(n4702), .ZN(U2947)
         );
  INV_X1 U5806 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6079) );
  NAND2_X1 U5807 ( .A1(n6125), .A2(LWORD_REG_11__SCAN_IN), .ZN(n4692) );
  NAND2_X1 U5808 ( .A1(n4694), .A2(DATAI_11_), .ZN(n4705) );
  OAI211_X1 U5809 ( .C1(n6079), .C2(n6105), .A(n4692), .B(n4705), .ZN(U2950)
         );
  INV_X1 U5810 ( .A(EAX_REG_10__SCAN_IN), .ZN(n6081) );
  NAND2_X1 U5811 ( .A1(n6125), .A2(LWORD_REG_10__SCAN_IN), .ZN(n4693) );
  NAND2_X1 U5812 ( .A1(n4694), .A2(DATAI_10_), .ZN(n4699) );
  OAI211_X1 U5813 ( .C1(n6081), .C2(n6105), .A(n4693), .B(n4699), .ZN(U2949)
         );
  NAND2_X1 U5814 ( .A1(n6125), .A2(UWORD_REG_14__SCAN_IN), .ZN(n4695) );
  NAND2_X1 U5815 ( .A1(n4694), .A2(DATAI_14_), .ZN(n4697) );
  OAI211_X1 U5816 ( .C1(n4696), .C2(n6105), .A(n4695), .B(n4697), .ZN(U2938)
         );
  INV_X1 U5817 ( .A(EAX_REG_14__SCAN_IN), .ZN(n6074) );
  NAND2_X1 U5818 ( .A1(n6125), .A2(LWORD_REG_14__SCAN_IN), .ZN(n4698) );
  OAI211_X1 U5819 ( .C1(n6074), .C2(n6105), .A(n4698), .B(n4697), .ZN(U2953)
         );
  NAND2_X1 U5820 ( .A1(n6125), .A2(UWORD_REG_10__SCAN_IN), .ZN(n4700) );
  OAI211_X1 U5821 ( .C1(n4701), .C2(n6105), .A(n4700), .B(n4699), .ZN(U2934)
         );
  NAND2_X1 U5822 ( .A1(n6125), .A2(UWORD_REG_8__SCAN_IN), .ZN(n4703) );
  OAI211_X1 U5823 ( .C1(n4704), .C2(n6105), .A(n4703), .B(n4702), .ZN(U2932)
         );
  NAND2_X1 U5824 ( .A1(n6125), .A2(UWORD_REG_11__SCAN_IN), .ZN(n4706) );
  OAI211_X1 U5825 ( .C1(n4707), .C2(n6105), .A(n4706), .B(n4705), .ZN(U2935)
         );
  INV_X1 U5826 ( .A(n6202), .ZN(n4708) );
  NAND2_X1 U5827 ( .A1(n4894), .A2(n3035), .ZN(n6348) );
  NAND3_X1 U5828 ( .A1(n4708), .A2(n6354), .A3(n6406), .ZN(n4710) );
  AOI21_X1 U5829 ( .B1(n4710), .B2(n4835), .A(n4709), .ZN(n4715) );
  NOR2_X1 U5830 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4711), .ZN(n6200)
         );
  NOR2_X1 U5831 ( .A1(n4716), .A2(n6342), .ZN(n6221) );
  INV_X1 U5832 ( .A(n6221), .ZN(n4891) );
  INV_X1 U5833 ( .A(n4761), .ZN(n4712) );
  OR2_X1 U5834 ( .A1(n6220), .A2(n4712), .ZN(n5008) );
  AOI21_X1 U5835 ( .B1(n5008), .B2(STATE2_REG_2__SCAN_IN), .A(n4713), .ZN(
        n5017) );
  OAI211_X1 U5836 ( .C1(n6761), .C2(n6200), .A(n4891), .B(n5017), .ZN(n4714)
         );
  INV_X1 U5837 ( .A(n6203), .ZN(n4726) );
  AOI22_X1 U5838 ( .A1(n5117), .A2(n6202), .B1(n6345), .B2(n6200), .ZN(n4718)
         );
  NOR2_X1 U5839 ( .A1(n4531), .A2(n6344), .ZN(n5011) );
  INV_X1 U5840 ( .A(n5011), .ZN(n6223) );
  AND2_X1 U5841 ( .A1(n4716), .A2(STATE2_REG_2__SCAN_IN), .ZN(n6226) );
  INV_X1 U5842 ( .A(n6226), .ZN(n5106) );
  OAI22_X1 U5843 ( .A1(n6223), .A2(n4801), .B1(n5008), .B2(n5106), .ZN(n6201)
         );
  AOI22_X1 U5844 ( .A1(n6346), .A2(n6201), .B1(n6356), .B2(n3078), .ZN(n4717)
         );
  OAI211_X1 U5845 ( .C1(n4726), .C2(n4719), .A(n4718), .B(n4717), .ZN(U3020)
         );
  AOI22_X1 U5846 ( .A1(n5123), .A2(n6202), .B1(n6378), .B2(n6200), .ZN(n4721)
         );
  AOI22_X1 U5847 ( .A1(n6379), .A2(n6201), .B1(n6380), .B2(n3078), .ZN(n4720)
         );
  OAI211_X1 U5848 ( .C1(n4726), .C2(n4722), .A(n4721), .B(n4720), .ZN(U3024)
         );
  AOI22_X1 U5849 ( .A1(n6326), .A2(n6202), .B1(n6391), .B2(n6200), .ZN(n4724)
         );
  AOI22_X1 U5850 ( .A1(n6392), .A2(n6201), .B1(n6393), .B2(n3078), .ZN(n4723)
         );
  OAI211_X1 U5851 ( .C1(n4726), .C2(n4725), .A(n4724), .B(n4723), .ZN(U3026)
         );
  NAND2_X1 U5852 ( .A1(n4894), .A2(n4727), .ZN(n4793) );
  NAND3_X1 U5853 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6415), .ZN(n4762) );
  INV_X1 U5854 ( .A(n4762), .ZN(n4729) );
  NOR2_X1 U5855 ( .A1(n6769), .A2(n4762), .ZN(n4752) );
  AOI21_X1 U5856 ( .B1(n6341), .B2(n5010), .A(n4752), .ZN(n4732) );
  NAND3_X1 U5857 ( .A1(n6354), .A2(n4732), .A3(n4730), .ZN(n4728) );
  OAI211_X1 U5858 ( .C1(n6354), .C2(n4729), .A(n6353), .B(n4728), .ZN(n4750)
         );
  NAND2_X1 U5859 ( .A1(n6354), .A2(n4730), .ZN(n4731) );
  OAI22_X1 U5860 ( .A1(n4732), .A2(n4731), .B1(n6342), .B2(n4762), .ZN(n4749)
         );
  AOI22_X1 U5861 ( .A1(INSTQUEUE_REG_13__2__SCAN_IN), .A2(n4750), .B1(n6367), 
        .B2(n4749), .ZN(n4736) );
  INV_X1 U5862 ( .A(n4733), .ZN(n4734) );
  NAND2_X1 U5863 ( .A1(n4894), .A2(n4734), .ZN(n4922) );
  INV_X1 U5864 ( .A(n4922), .ZN(n4751) );
  AOI22_X1 U5865 ( .A1(n6366), .A2(n4752), .B1(n4751), .B2(n6368), .ZN(n4735)
         );
  OAI211_X1 U5866 ( .C1(n6371), .C2(n4793), .A(n4736), .B(n4735), .ZN(U3126)
         );
  AOI22_X1 U5867 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n4750), .B1(n6385), 
        .B2(n4749), .ZN(n4738) );
  AOI22_X1 U5868 ( .A1(n6384), .A2(n4752), .B1(n4751), .B2(n6386), .ZN(n4737)
         );
  OAI211_X1 U5869 ( .C1(n6390), .C2(n4793), .A(n4738), .B(n4737), .ZN(U3129)
         );
  AOI22_X1 U5870 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n4750), .B1(n6361), 
        .B2(n4749), .ZN(n4740) );
  AOI22_X1 U5871 ( .A1(n6360), .A2(n4752), .B1(n4751), .B2(n6362), .ZN(n4739)
         );
  OAI211_X1 U5872 ( .C1(n6365), .C2(n4793), .A(n4740), .B(n4739), .ZN(U3125)
         );
  AOI22_X1 U5873 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n4750), .B1(n6392), 
        .B2(n4749), .ZN(n4742) );
  AOI22_X1 U5874 ( .A1(n6391), .A2(n4752), .B1(n4751), .B2(n6326), .ZN(n4741)
         );
  OAI211_X1 U5875 ( .C1(n6329), .C2(n4793), .A(n4742), .B(n4741), .ZN(U3130)
         );
  AOI22_X1 U5876 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4750), .B1(n6379), 
        .B2(n4749), .ZN(n4744) );
  AOI22_X1 U5877 ( .A1(n6378), .A2(n4752), .B1(n4751), .B2(n5123), .ZN(n4743)
         );
  OAI211_X1 U5878 ( .C1(n5121), .C2(n4793), .A(n4744), .B(n4743), .ZN(U3128)
         );
  AOI22_X1 U5879 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n4750), .B1(n6400), 
        .B2(n4749), .ZN(n4746) );
  AOI22_X1 U5880 ( .A1(n6397), .A2(n4752), .B1(n4751), .B2(n6330), .ZN(n4745)
         );
  OAI211_X1 U5881 ( .C1(n6338), .C2(n4793), .A(n4746), .B(n4745), .ZN(U3131)
         );
  AOI22_X1 U5882 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(n4750), .B1(n6346), 
        .B2(n4749), .ZN(n4748) );
  AOI22_X1 U5883 ( .A1(n6345), .A2(n4752), .B1(n5117), .B2(n4751), .ZN(n4747)
         );
  OAI211_X1 U5884 ( .C1(n5115), .C2(n4793), .A(n4748), .B(n4747), .ZN(U3124)
         );
  AOI22_X1 U5885 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n4750), .B1(n6373), 
        .B2(n4749), .ZN(n4754) );
  AOI22_X1 U5886 ( .A1(n6372), .A2(n4752), .B1(n4751), .B2(n6316), .ZN(n4753)
         );
  OAI211_X1 U5887 ( .C1(n6319), .C2(n4793), .A(n4754), .B(n4753), .ZN(U3127)
         );
  INV_X1 U5888 ( .A(n4755), .ZN(n6025) );
  AOI21_X1 U5889 ( .B1(n6134), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n4756), 
        .ZN(n4757) );
  OAI21_X1 U5890 ( .B1(n6027), .B2(n6143), .A(n4757), .ZN(n4758) );
  AOI21_X1 U5891 ( .B1(n6025), .B2(n6347), .A(n4758), .ZN(n4759) );
  OAI21_X1 U5892 ( .B1(n5926), .B2(n4760), .A(n4759), .ZN(U2981) );
  NOR2_X1 U5893 ( .A1(n6032), .A2(n6344), .ZN(n4893) );
  AOI22_X1 U5894 ( .A1(n4893), .A2(n5010), .B1(n6221), .B2(n3105), .ZN(n4798)
         );
  NOR2_X1 U5895 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4762), .ZN(n4770)
         );
  AND2_X1 U5896 ( .A1(n3035), .A2(n4763), .ZN(n4803) );
  NAND2_X1 U5897 ( .A1(n6298), .A2(n4803), .ZN(n6323) );
  INV_X1 U5898 ( .A(n4793), .ZN(n4764) );
  NOR3_X1 U5899 ( .A1(n6331), .A2(n4764), .A3(n6344), .ZN(n4767) );
  INV_X1 U5900 ( .A(n4835), .ZN(n6350) );
  INV_X1 U5901 ( .A(n5010), .ZN(n4765) );
  OAI22_X1 U5902 ( .A1(n4767), .A2(n6350), .B1(n4766), .B2(n4765), .ZN(n4769)
         );
  OAI21_X1 U5903 ( .B1(n3105), .B2(n6342), .A(n4839), .ZN(n4800) );
  NOR2_X1 U5904 ( .A1(n6226), .A2(n4800), .ZN(n4768) );
  OAI211_X1 U5905 ( .C1(n4770), .C2(n6761), .A(n4769), .B(n4768), .ZN(n4792)
         );
  NAND2_X1 U5906 ( .A1(n4792), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4773)
         );
  INV_X1 U5907 ( .A(n4770), .ZN(n4794) );
  OAI22_X1 U5908 ( .A1(n5052), .A2(n4794), .B1(n6243), .B2(n4793), .ZN(n4771)
         );
  AOI21_X1 U5909 ( .B1(n6240), .B2(n6331), .A(n4771), .ZN(n4772) );
  OAI211_X1 U5910 ( .C1(n4798), .C2(n5152), .A(n4773), .B(n4772), .ZN(U3121)
         );
  NAND2_X1 U5911 ( .A1(n4792), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4776)
         );
  OAI22_X1 U5912 ( .A1(n5022), .A2(n4794), .B1(n6315), .B2(n4793), .ZN(n4774)
         );
  AOI21_X1 U5913 ( .B1(n6312), .B2(n6331), .A(n4774), .ZN(n4775) );
  OAI211_X1 U5914 ( .C1(n4798), .C2(n5137), .A(n4776), .B(n4775), .ZN(U3118)
         );
  NAND2_X1 U5915 ( .A1(n4792), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4779)
         );
  OAI22_X1 U5916 ( .A1(n5026), .A2(n4794), .B1(n6377), .B2(n4793), .ZN(n4777)
         );
  AOI21_X1 U5917 ( .B1(n6374), .B2(n6331), .A(n4777), .ZN(n4778) );
  OAI211_X1 U5918 ( .C1(n4798), .C2(n5145), .A(n4779), .B(n4778), .ZN(U3119)
         );
  NAND2_X1 U5919 ( .A1(n4792), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n4782)
         );
  OAI22_X1 U5920 ( .A1(n5030), .A2(n4794), .B1(n6407), .B2(n4793), .ZN(n4780)
         );
  AOI21_X1 U5921 ( .B1(n6402), .B2(n6331), .A(n4780), .ZN(n4781) );
  OAI211_X1 U5922 ( .C1(n4798), .C2(n5133), .A(n4782), .B(n4781), .ZN(U3123)
         );
  NAND2_X1 U5923 ( .A1(n4792), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4785)
         );
  OAI22_X1 U5924 ( .A1(n5038), .A2(n4794), .B1(n6383), .B2(n4793), .ZN(n4783)
         );
  AOI21_X1 U5925 ( .B1(n6380), .B2(n6331), .A(n4783), .ZN(n4784) );
  OAI211_X1 U5926 ( .C1(n4798), .C2(n5125), .A(n4785), .B(n4784), .ZN(U3120)
         );
  NAND2_X1 U5927 ( .A1(n4792), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n4788)
         );
  OAI22_X1 U5928 ( .A1(n5034), .A2(n4794), .B1(n6396), .B2(n4793), .ZN(n4786)
         );
  AOI21_X1 U5929 ( .B1(n6393), .B2(n6331), .A(n4786), .ZN(n4787) );
  OAI211_X1 U5930 ( .C1(n4798), .C2(n5129), .A(n4788), .B(n4787), .ZN(U3122)
         );
  NAND2_X1 U5931 ( .A1(n4792), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n4791)
         );
  OAI22_X1 U5932 ( .A1(n5042), .A2(n4794), .B1(n6359), .B2(n4793), .ZN(n4789)
         );
  AOI21_X1 U5933 ( .B1(n6356), .B2(n6331), .A(n4789), .ZN(n4790) );
  OAI211_X1 U5934 ( .C1(n4798), .C2(n5119), .A(n4791), .B(n4790), .ZN(U3116)
         );
  NAND2_X1 U5935 ( .A1(n4792), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n4797)
         );
  OAI22_X1 U5936 ( .A1(n5046), .A2(n4794), .B1(n6267), .B2(n4793), .ZN(n4795)
         );
  AOI21_X1 U5937 ( .B1(n6264), .B2(n6331), .A(n4795), .ZN(n4796) );
  OAI211_X1 U5938 ( .C1(n4798), .C2(n5141), .A(n4797), .B(n4796), .ZN(U3117)
         );
  AOI22_X1 U5939 ( .A1(n4893), .A2(n4802), .B1(n6226), .B2(n3105), .ZN(n6286)
         );
  NOR2_X1 U5940 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4799), .ZN(n6289)
         );
  INV_X1 U5941 ( .A(n6289), .ZN(n4823) );
  AOI211_X1 U5942 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n4823), .A(n6221), .B(
        n4800), .ZN(n4807) );
  NAND2_X1 U5943 ( .A1(n4801), .A2(n6350), .ZN(n4806) );
  NOR2_X1 U5944 ( .A1(n4802), .A2(n6344), .ZN(n4804) );
  NAND2_X1 U5945 ( .A1(n6219), .A2(n4803), .ZN(n6295) );
  OAI211_X1 U5946 ( .C1(n5011), .C2(n4804), .A(n4824), .B(n6295), .ZN(n4805)
         );
  NAND3_X1 U5947 ( .A1(n4807), .A2(n4806), .A3(n4805), .ZN(n6292) );
  NAND2_X1 U5948 ( .A1(n6292), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n4810) );
  OAI22_X1 U5949 ( .A1(n4824), .A2(n6315), .B1(n5022), .B2(n4823), .ZN(n4808)
         );
  AOI21_X1 U5950 ( .B1(n6312), .B2(n6274), .A(n4808), .ZN(n4809) );
  OAI211_X1 U5951 ( .C1(n6286), .C2(n5137), .A(n4810), .B(n4809), .ZN(U3086)
         );
  NAND2_X1 U5952 ( .A1(n6292), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n4813) );
  OAI22_X1 U5953 ( .A1(n4824), .A2(n6359), .B1(n5042), .B2(n4823), .ZN(n4811)
         );
  AOI21_X1 U5954 ( .B1(n6356), .B2(n6274), .A(n4811), .ZN(n4812) );
  OAI211_X1 U5955 ( .C1(n6286), .C2(n5119), .A(n4813), .B(n4812), .ZN(U3084)
         );
  NAND2_X1 U5956 ( .A1(n6292), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n4816) );
  OAI22_X1 U5957 ( .A1(n4824), .A2(n6243), .B1(n5052), .B2(n4823), .ZN(n4814)
         );
  AOI21_X1 U5958 ( .B1(n6240), .B2(n6274), .A(n4814), .ZN(n4815) );
  OAI211_X1 U5959 ( .C1(n6286), .C2(n5152), .A(n4816), .B(n4815), .ZN(U3089)
         );
  NAND2_X1 U5960 ( .A1(n6292), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n4819) );
  OAI22_X1 U5961 ( .A1(n4824), .A2(n6396), .B1(n5034), .B2(n4823), .ZN(n4817)
         );
  AOI21_X1 U5962 ( .B1(n6393), .B2(n6274), .A(n4817), .ZN(n4818) );
  OAI211_X1 U5963 ( .C1(n6286), .C2(n5129), .A(n4819), .B(n4818), .ZN(U3090)
         );
  NAND2_X1 U5964 ( .A1(n6292), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4822) );
  OAI22_X1 U5965 ( .A1(n4824), .A2(n6407), .B1(n5030), .B2(n4823), .ZN(n4820)
         );
  AOI21_X1 U5966 ( .B1(n6402), .B2(n6274), .A(n4820), .ZN(n4821) );
  OAI211_X1 U5967 ( .C1(n6286), .C2(n5133), .A(n4822), .B(n4821), .ZN(U3091)
         );
  NAND2_X1 U5968 ( .A1(n6292), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n4827) );
  OAI22_X1 U5969 ( .A1(n4824), .A2(n6383), .B1(n5038), .B2(n4823), .ZN(n4825)
         );
  AOI21_X1 U5970 ( .B1(n6380), .B2(n6274), .A(n4825), .ZN(n4826) );
  OAI211_X1 U5971 ( .C1(n6286), .C2(n5125), .A(n4827), .B(n4826), .ZN(U3088)
         );
  INV_X1 U5972 ( .A(n6005), .ZN(n4830) );
  AOI22_X1 U5973 ( .A1(n6134), .A2(PHYADDRPOINTER_REG_6__SCAN_IN), .B1(n6582), 
        .B2(REIP_REG_6__SCAN_IN), .ZN(n4828) );
  OAI21_X1 U5974 ( .B1(n6012), .B2(n6143), .A(n4828), .ZN(n4829) );
  AOI21_X1 U5975 ( .B1(n4830), .B2(n6347), .A(n4829), .ZN(n4831) );
  OAI21_X1 U5976 ( .B1(n5926), .B2(n4832), .A(n4831), .ZN(U2980) );
  NOR2_X1 U5977 ( .A1(n5106), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n4833)
         );
  AOI22_X1 U5978 ( .A1(n5011), .A2(n5105), .B1(n6220), .B2(n4833), .ZN(n4870)
         );
  OAI21_X1 U5979 ( .B1(n4867), .B2(n6211), .A(n4835), .ZN(n4837) );
  AOI21_X1 U5980 ( .B1(n4837), .B2(n4836), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n4840) );
  NOR2_X1 U5981 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n4838), .ZN(n4841)
         );
  OAI21_X1 U5982 ( .B1(n6220), .B2(n6342), .A(n4839), .ZN(n6225) );
  NOR2_X1 U5983 ( .A1(n6221), .A2(n6225), .ZN(n5113) );
  OAI21_X1 U5984 ( .B1(n4840), .B2(n4841), .A(n5113), .ZN(n4863) );
  NAND2_X1 U5985 ( .A1(n4863), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4844) );
  INV_X1 U5986 ( .A(n4841), .ZN(n4864) );
  OAI22_X1 U5987 ( .A1(n6377), .A2(n4865), .B1(n5026), .B2(n4864), .ZN(n4842)
         );
  AOI21_X1 U5988 ( .B1(n6374), .B2(n4867), .A(n4842), .ZN(n4843) );
  OAI211_X1 U5989 ( .C1(n4870), .C2(n5145), .A(n4844), .B(n4843), .ZN(U3039)
         );
  NAND2_X1 U5990 ( .A1(n4863), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4847) );
  OAI22_X1 U5991 ( .A1(n6315), .A2(n4865), .B1(n5022), .B2(n4864), .ZN(n4845)
         );
  AOI21_X1 U5992 ( .B1(n6312), .B2(n4867), .A(n4845), .ZN(n4846) );
  OAI211_X1 U5993 ( .C1(n4870), .C2(n5137), .A(n4847), .B(n4846), .ZN(U3038)
         );
  NAND2_X1 U5994 ( .A1(n4863), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4850) );
  OAI22_X1 U5995 ( .A1(n6243), .A2(n4865), .B1(n5052), .B2(n4864), .ZN(n4848)
         );
  AOI21_X1 U5996 ( .B1(n6240), .B2(n4867), .A(n4848), .ZN(n4849) );
  OAI211_X1 U5997 ( .C1(n4870), .C2(n5152), .A(n4850), .B(n4849), .ZN(U3041)
         );
  NAND2_X1 U5998 ( .A1(n4863), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n4853) );
  OAI22_X1 U5999 ( .A1(n6267), .A2(n4865), .B1(n5046), .B2(n4864), .ZN(n4851)
         );
  AOI21_X1 U6000 ( .B1(n6264), .B2(n4867), .A(n4851), .ZN(n4852) );
  OAI211_X1 U6001 ( .C1(n4870), .C2(n5141), .A(n4853), .B(n4852), .ZN(U3037)
         );
  NAND2_X1 U6002 ( .A1(n4863), .A2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4856) );
  OAI22_X1 U6003 ( .A1(n6407), .A2(n4865), .B1(n5030), .B2(n4864), .ZN(n4854)
         );
  AOI21_X1 U6004 ( .B1(n6402), .B2(n4867), .A(n4854), .ZN(n4855) );
  OAI211_X1 U6005 ( .C1(n4870), .C2(n5133), .A(n4856), .B(n4855), .ZN(U3043)
         );
  NAND2_X1 U6006 ( .A1(n4863), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4859) );
  OAI22_X1 U6007 ( .A1(n5042), .A2(n4864), .B1(n6359), .B2(n4865), .ZN(n4857)
         );
  AOI21_X1 U6008 ( .B1(n6356), .B2(n4867), .A(n4857), .ZN(n4858) );
  OAI211_X1 U6009 ( .C1(n4870), .C2(n5119), .A(n4859), .B(n4858), .ZN(U3036)
         );
  NAND2_X1 U6010 ( .A1(n4863), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4862) );
  OAI22_X1 U6011 ( .A1(n6383), .A2(n4865), .B1(n5038), .B2(n4864), .ZN(n4860)
         );
  AOI21_X1 U6012 ( .B1(n6380), .B2(n4867), .A(n4860), .ZN(n4861) );
  OAI211_X1 U6013 ( .C1(n4870), .C2(n5125), .A(n4862), .B(n4861), .ZN(U3040)
         );
  NAND2_X1 U6014 ( .A1(n4863), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4869) );
  OAI22_X1 U6015 ( .A1(n6396), .A2(n4865), .B1(n5034), .B2(n4864), .ZN(n4866)
         );
  AOI21_X1 U6016 ( .B1(n6393), .B2(n4867), .A(n4866), .ZN(n4868) );
  OAI211_X1 U6017 ( .C1(n4870), .C2(n5129), .A(n4869), .B(n4868), .ZN(U3042)
         );
  NAND2_X1 U6018 ( .A1(n4581), .A2(n4873), .ZN(n4874) );
  NAND2_X1 U6019 ( .A1(n4872), .A2(n4874), .ZN(n5994) );
  INV_X1 U6020 ( .A(EBX_REG_7__SCAN_IN), .ZN(n4878) );
  AND2_X1 U6021 ( .A1(n4876), .A2(n4875), .ZN(n4877) );
  OR2_X1 U6022 ( .A1(n4935), .A2(n4877), .ZN(n6162) );
  OAI222_X1 U6023 ( .A1(n5994), .A2(n5589), .B1(n4878), .B2(n6053), .C1(n6162), 
        .C2(n5597), .ZN(U2852) );
  INV_X1 U6024 ( .A(EAX_REG_7__SCAN_IN), .ZN(n6087) );
  OAI222_X1 U6025 ( .A1(n5994), .A2(n5603), .B1(n5306), .B2(n6124), .C1(n5504), 
        .C2(n6087), .ZN(U2884) );
  INV_X1 U6026 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n4879) );
  AND2_X1 U6027 ( .A1(n5860), .A2(n4879), .ZN(n4880) );
  AOI211_X1 U6028 ( .C1(n6134), .C2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n4881), 
        .B(n4880), .ZN(n4884) );
  INV_X1 U6029 ( .A(n5926), .ZN(n6150) );
  NAND3_X1 U6030 ( .A1(n4882), .A2(n6150), .A3(n4392), .ZN(n4883) );
  OAI211_X1 U6031 ( .C1(n5103), .C2(n5642), .A(n4884), .B(n4883), .ZN(U2985)
         );
  XOR2_X1 U6032 ( .A(n4886), .B(n4885), .Z(n6166) );
  NAND2_X1 U6033 ( .A1(n6166), .A2(n6150), .ZN(n4890) );
  NAND2_X1 U6034 ( .A1(n6582), .A2(REIP_REG_7__SCAN_IN), .ZN(n6161) );
  INV_X1 U6035 ( .A(n6161), .ZN(n4888) );
  NOR2_X1 U6036 ( .A1(n6143), .A2(n5998), .ZN(n4887) );
  AOI211_X1 U6037 ( .C1(n6134), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n4888), 
        .B(n4887), .ZN(n4889) );
  OAI211_X1 U6038 ( .C1(n5642), .C2(n5994), .A(n4890), .B(n4889), .ZN(U2979)
         );
  AND2_X1 U6039 ( .A1(n4340), .A2(n5097), .ZN(n6340) );
  NOR2_X1 U6040 ( .A1(n4891), .A2(n6425), .ZN(n4892) );
  AOI22_X1 U6041 ( .A1(n4893), .A2(n6340), .B1(n6220), .B2(n4892), .ZN(n4927)
         );
  NOR2_X1 U6042 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6343), .ZN(n4899)
         );
  AOI21_X1 U6043 ( .B1(n6389), .B2(n4922), .A(n5925), .ZN(n4896) );
  INV_X1 U6044 ( .A(n6340), .ZN(n6254) );
  NAND2_X1 U6045 ( .A1(n6254), .A2(n6354), .ZN(n4895) );
  NOR2_X1 U6046 ( .A1(n4896), .A2(n4895), .ZN(n4897) );
  NOR4_X1 U6047 ( .A1(n6425), .A2(n6226), .A3(n4897), .A4(n6225), .ZN(n4898)
         );
  NAND2_X1 U6048 ( .A1(n4921), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4902)
         );
  INV_X1 U6049 ( .A(n4899), .ZN(n4923) );
  OAI22_X1 U6050 ( .A1(n5042), .A2(n4923), .B1(n5115), .B2(n4922), .ZN(n4900)
         );
  AOI21_X1 U6051 ( .B1(n5117), .B2(n6401), .A(n4900), .ZN(n4901) );
  OAI211_X1 U6052 ( .C1(n4927), .C2(n5119), .A(n4902), .B(n4901), .ZN(U3132)
         );
  NAND2_X1 U6053 ( .A1(n4921), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n4905)
         );
  OAI22_X1 U6054 ( .A1(n5046), .A2(n4923), .B1(n4922), .B2(n6365), .ZN(n4903)
         );
  AOI21_X1 U6055 ( .B1(n6401), .B2(n6362), .A(n4903), .ZN(n4904) );
  OAI211_X1 U6056 ( .C1(n4927), .C2(n5141), .A(n4905), .B(n4904), .ZN(U3133)
         );
  NAND2_X1 U6057 ( .A1(n4921), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n4908)
         );
  OAI22_X1 U6058 ( .A1(n5026), .A2(n4923), .B1(n4922), .B2(n6319), .ZN(n4906)
         );
  AOI21_X1 U6059 ( .B1(n6401), .B2(n6316), .A(n4906), .ZN(n4907) );
  OAI211_X1 U6060 ( .C1(n4927), .C2(n5145), .A(n4908), .B(n4907), .ZN(U3135)
         );
  NAND2_X1 U6061 ( .A1(n4921), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4911)
         );
  OAI22_X1 U6062 ( .A1(n5034), .A2(n4923), .B1(n4922), .B2(n6329), .ZN(n4909)
         );
  AOI21_X1 U6063 ( .B1(n6401), .B2(n6326), .A(n4909), .ZN(n4910) );
  OAI211_X1 U6064 ( .C1(n4927), .C2(n5129), .A(n4911), .B(n4910), .ZN(U3138)
         );
  NAND2_X1 U6065 ( .A1(n4921), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n4914)
         );
  OAI22_X1 U6066 ( .A1(n5052), .A2(n4923), .B1(n4922), .B2(n6390), .ZN(n4912)
         );
  AOI21_X1 U6067 ( .B1(n6401), .B2(n6386), .A(n4912), .ZN(n4913) );
  OAI211_X1 U6068 ( .C1(n4927), .C2(n5152), .A(n4914), .B(n4913), .ZN(U3137)
         );
  NAND2_X1 U6069 ( .A1(n4921), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4917)
         );
  OAI22_X1 U6070 ( .A1(n5038), .A2(n4923), .B1(n4922), .B2(n5121), .ZN(n4915)
         );
  AOI21_X1 U6071 ( .B1(n6401), .B2(n5123), .A(n4915), .ZN(n4916) );
  OAI211_X1 U6072 ( .C1(n4927), .C2(n5125), .A(n4917), .B(n4916), .ZN(U3136)
         );
  NAND2_X1 U6073 ( .A1(n4921), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n4920)
         );
  OAI22_X1 U6074 ( .A1(n5022), .A2(n4923), .B1(n4922), .B2(n6371), .ZN(n4918)
         );
  AOI21_X1 U6075 ( .B1(n6401), .B2(n6368), .A(n4918), .ZN(n4919) );
  OAI211_X1 U6076 ( .C1(n4927), .C2(n5137), .A(n4920), .B(n4919), .ZN(U3134)
         );
  NAND2_X1 U6077 ( .A1(n4921), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4926)
         );
  OAI22_X1 U6078 ( .A1(n5030), .A2(n4923), .B1(n4922), .B2(n6338), .ZN(n4924)
         );
  AOI21_X1 U6079 ( .B1(n6401), .B2(n6330), .A(n4924), .ZN(n4925) );
  OAI211_X1 U6080 ( .C1(n4927), .C2(n5133), .A(n4926), .B(n4925), .ZN(U3139)
         );
  XNOR2_X1 U6081 ( .A(n4928), .B(n4929), .ZN(n4998) );
  OAI22_X1 U6082 ( .A1(n4933), .A2(n4932), .B1(n4931), .B2(n4930), .ZN(n6160)
         );
  OAI21_X1 U6083 ( .B1(n4935), .B2(n4934), .A(n4968), .ZN(n5976) );
  NAND2_X1 U6084 ( .A1(n6582), .A2(REIP_REG_8__SCAN_IN), .ZN(n4994) );
  OAI21_X1 U6085 ( .B1(n6584), .B2(n5976), .A(n4994), .ZN(n4940) );
  NAND2_X1 U6086 ( .A1(n4937), .A2(n4936), .ZN(n6163) );
  OAI21_X1 U6087 ( .B1(INSTADDRPOINTER_REG_8__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_7__SCAN_IN), .A(n5066), .ZN(n4938) );
  NOR2_X1 U6088 ( .A1(n6163), .A2(n4938), .ZN(n4939) );
  AOI211_X1 U6089 ( .C1(n6160), .C2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n4940), 
        .B(n4939), .ZN(n4941) );
  OAI21_X1 U6090 ( .B1(n6589), .B2(n4998), .A(n4941), .ZN(U3010) );
  NOR3_X1 U6091 ( .A1(STATEBS16_REG_SCAN_IN), .A2(n6457), .A3(n6548), .ZN(
        n6453) );
  INV_X1 U6092 ( .A(n6453), .ZN(n4942) );
  NAND2_X1 U6093 ( .A1(n5908), .A2(n4942), .ZN(n4944) );
  NOR3_X1 U6094 ( .A1(n6596), .A2(n6761), .A3(n6446), .ZN(n4943) );
  OR2_X1 U6095 ( .A1(n4944), .A2(n4943), .ZN(n4945) );
  NOR2_X1 U6096 ( .A1(n4962), .A2(n6548), .ZN(n4946) );
  NAND2_X1 U6097 ( .A1(n5519), .A2(n4956), .ZN(n4947) );
  NAND2_X1 U6098 ( .A1(n6004), .A2(n4947), .ZN(n6024) );
  INV_X1 U6099 ( .A(n6024), .ZN(n6038) );
  NAND2_X1 U6100 ( .A1(n6568), .A2(n5925), .ZN(n4957) );
  INV_X1 U6101 ( .A(n4957), .ZN(n4948) );
  NAND2_X1 U6102 ( .A1(n5281), .A2(n5529), .ZN(n5987) );
  INV_X1 U6103 ( .A(n4956), .ZN(n4951) );
  NOR2_X1 U6104 ( .A1(n4952), .A2(n4951), .ZN(n5096) );
  INV_X1 U6105 ( .A(n5096), .ZN(n6033) );
  NOR2_X1 U6106 ( .A1(n6412), .A2(n6033), .ZN(n4961) );
  NOR3_X1 U6107 ( .A1(READY_N), .A2(STATEBS16_REG_SCAN_IN), .A3(n6469), .ZN(
        n6435) );
  INV_X1 U6108 ( .A(n6435), .ZN(n4953) );
  NAND2_X1 U6109 ( .A1(n6436), .A2(n4953), .ZN(n5531) );
  INV_X1 U6110 ( .A(EBX_REG_31__SCAN_IN), .ZN(n5431) );
  NAND3_X1 U6111 ( .A1(n3271), .A2(n5431), .A3(n4957), .ZN(n4954) );
  NAND2_X1 U6112 ( .A1(n5531), .A2(n4954), .ZN(n4955) );
  AND2_X1 U6113 ( .A1(EBX_REG_31__SCAN_IN), .A2(n4956), .ZN(n5530) );
  OAI22_X1 U6114 ( .A1(n5974), .A2(n4959), .B1(n6183), .B2(n6035), .ZN(n4960)
         );
  AOI211_X1 U6115 ( .C1(n5987), .C2(REIP_REG_0__SCAN_IN), .A(n4961), .B(n4960), 
        .ZN(n4965) );
  AND2_X1 U6116 ( .A1(n4962), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4963) );
  OAI21_X1 U6117 ( .B1(n6003), .B2(n5979), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n4964) );
  OAI211_X1 U6118 ( .C1(n6038), .C2(n6152), .A(n4965), .B(n4964), .ZN(U2827)
         );
  XNOR2_X1 U6119 ( .A(n4966), .B(n4967), .ZN(n5081) );
  AOI21_X1 U6120 ( .B1(n4969), .B2(n4968), .A(n3068), .ZN(n5964) );
  NOR2_X1 U6121 ( .A1(n5066), .A2(n6163), .ZN(n4972) );
  INV_X1 U6122 ( .A(n5066), .ZN(n4970) );
  NOR2_X1 U6123 ( .A1(n5887), .A2(n4970), .ZN(n4971) );
  OR2_X1 U6124 ( .A1(n6160), .A2(n4971), .ZN(n5073) );
  MUX2_X1 U6125 ( .A(n4972), .B(n5073), .S(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .Z(n4974) );
  INV_X1 U6126 ( .A(REIP_REG_9__SCAN_IN), .ZN(n6495) );
  NOR2_X1 U6127 ( .A1(n5908), .A2(n6495), .ZN(n4973) );
  AOI211_X1 U6128 ( .C1(n6170), .C2(n5964), .A(n4974), .B(n4973), .ZN(n4975)
         );
  OAI21_X1 U6129 ( .B1(n5081), .B2(n6589), .A(n4975), .ZN(U3009) );
  AOI21_X1 U6130 ( .B1(n4977), .B2(n4872), .A(n4976), .ZN(n5981) );
  INV_X1 U6131 ( .A(n5981), .ZN(n4981) );
  INV_X1 U6132 ( .A(n5306), .ZN(n5276) );
  AOI22_X1 U6133 ( .A1(n5276), .A2(DATAI_8_), .B1(EAX_REG_8__SCAN_IN), .B2(
        n6063), .ZN(n4978) );
  OAI21_X1 U6134 ( .B1(n4981), .B2(n5603), .A(n4978), .ZN(U2883) );
  INV_X1 U6135 ( .A(n5976), .ZN(n4979) );
  AOI22_X1 U6136 ( .A1(n6049), .A2(n4979), .B1(EBX_REG_8__SCAN_IN), .B2(n5590), 
        .ZN(n4980) );
  OAI21_X1 U6137 ( .B1(n4981), .B2(n5589), .A(n4980), .ZN(U2851) );
  NAND2_X1 U6138 ( .A1(n4982), .A2(n6024), .ZN(n4991) );
  NAND2_X1 U6139 ( .A1(n5915), .A2(n5096), .ZN(n4987) );
  INV_X1 U6140 ( .A(REIP_REG_2__SCAN_IN), .ZN(n6482) );
  NOR3_X1 U6141 ( .A1(n5099), .A2(n6484), .A3(n6482), .ZN(n5162) );
  INV_X1 U6142 ( .A(n5162), .ZN(n4983) );
  OR2_X1 U6143 ( .A1(n5529), .A2(n4983), .ZN(n5168) );
  OAI21_X1 U6144 ( .B1(n5163), .B2(n4983), .A(n5987), .ZN(n6045) );
  NAND2_X1 U6145 ( .A1(n5281), .A2(n4984), .ZN(n6015) );
  OAI221_X1 U6146 ( .B1(REIP_REG_4__SCAN_IN), .B2(n5168), .C1(n6486), .C2(
        n6045), .A(n6015), .ZN(n4985) );
  AOI21_X1 U6147 ( .B1(n6042), .B2(EBX_REG_4__SCAN_IN), .A(n4985), .ZN(n4986)
         );
  OAI211_X1 U6148 ( .C1(n4988), .C2(n6035), .A(n4987), .B(n4986), .ZN(n4989)
         );
  AOI21_X1 U6149 ( .B1(n6003), .B2(PHYADDRPOINTER_REG_4__SCAN_IN), .A(n4989), 
        .ZN(n4990) );
  OAI211_X1 U6150 ( .C1(n4992), .C2(n6036), .A(n4991), .B(n4990), .ZN(U2823)
         );
  NAND2_X1 U6151 ( .A1(n6134), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n4993)
         );
  OAI211_X1 U6152 ( .C1(n6143), .C2(n4995), .A(n4994), .B(n4993), .ZN(n4996)
         );
  AOI21_X1 U6153 ( .B1(n5981), .B2(n6347), .A(n4996), .ZN(n4997) );
  OAI21_X1 U6154 ( .B1(n5926), .B2(n4998), .A(n4997), .ZN(U2978) );
  OR2_X1 U6155 ( .A1(n5529), .A2(REIP_REG_1__SCAN_IN), .ZN(n5093) );
  NAND2_X1 U6156 ( .A1(n5281), .A2(n5093), .ZN(n6028) );
  NOR3_X1 U6157 ( .A1(n5529), .A2(REIP_REG_2__SCAN_IN), .A3(n5099), .ZN(n4999)
         );
  AOI21_X1 U6158 ( .B1(n6042), .B2(EBX_REG_2__SCAN_IN), .A(n4999), .ZN(n5002)
         );
  XNOR2_X1 U6159 ( .A(n4507), .B(n5000), .ZN(n6169) );
  NAND2_X1 U6160 ( .A1(n6169), .A2(n6013), .ZN(n5001) );
  OAI211_X1 U6161 ( .C1(n5723), .C2(n6033), .A(n5002), .B(n5001), .ZN(n5003)
         );
  AOI21_X1 U6162 ( .B1(n6028), .B2(REIP_REG_2__SCAN_IN), .A(n5003), .ZN(n5006)
         );
  INV_X1 U6163 ( .A(n6142), .ZN(n5004) );
  AOI22_X1 U6164 ( .A1(n5004), .A2(n5979), .B1(n6003), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5005) );
  OAI211_X1 U6165 ( .C1(n5007), .C2(n6038), .A(n5006), .B(n5005), .ZN(U2825)
         );
  INV_X1 U6166 ( .A(n5008), .ZN(n5009) );
  AOI22_X1 U6167 ( .A1(n5011), .A2(n5010), .B1(n6221), .B2(n5009), .ZN(n5057)
         );
  NOR2_X1 U6168 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5012), .ZN(n5021)
         );
  AOI21_X1 U6169 ( .B1(n5013), .B2(n6217), .A(n5925), .ZN(n5016) );
  INV_X1 U6170 ( .A(n5014), .ZN(n5015) );
  NOR2_X1 U6171 ( .A1(n5016), .A2(n5015), .ZN(n5019) );
  INV_X1 U6172 ( .A(n5017), .ZN(n5018) );
  AOI211_X1 U6173 ( .C1(n6354), .C2(n5019), .A(n6226), .B(n5018), .ZN(n5020)
         );
  OAI21_X1 U6174 ( .B1(n5021), .B2(n6761), .A(n5020), .ZN(n5050) );
  NAND2_X1 U6175 ( .A1(n5050), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n5025) );
  INV_X1 U6176 ( .A(n5021), .ZN(n5051) );
  OAI22_X1 U6177 ( .A1(n5022), .A2(n5051), .B1(n6371), .B2(n6217), .ZN(n5023)
         );
  AOI21_X1 U6178 ( .B1(n6368), .B2(n5054), .A(n5023), .ZN(n5024) );
  OAI211_X1 U6179 ( .C1(n5057), .C2(n5137), .A(n5025), .B(n5024), .ZN(U3054)
         );
  NAND2_X1 U6180 ( .A1(n5050), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n5029) );
  OAI22_X1 U6181 ( .A1(n5026), .A2(n5051), .B1(n6319), .B2(n6217), .ZN(n5027)
         );
  AOI21_X1 U6182 ( .B1(n6316), .B2(n5054), .A(n5027), .ZN(n5028) );
  OAI211_X1 U6183 ( .C1(n5057), .C2(n5145), .A(n5029), .B(n5028), .ZN(U3055)
         );
  NAND2_X1 U6184 ( .A1(n5050), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n5033) );
  OAI22_X1 U6185 ( .A1(n5030), .A2(n5051), .B1(n6338), .B2(n6217), .ZN(n5031)
         );
  AOI21_X1 U6186 ( .B1(n6330), .B2(n5054), .A(n5031), .ZN(n5032) );
  OAI211_X1 U6187 ( .C1(n5057), .C2(n5133), .A(n5033), .B(n5032), .ZN(U3059)
         );
  NAND2_X1 U6188 ( .A1(n5050), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n5037) );
  OAI22_X1 U6189 ( .A1(n5034), .A2(n5051), .B1(n6329), .B2(n6217), .ZN(n5035)
         );
  AOI21_X1 U6190 ( .B1(n6326), .B2(n5054), .A(n5035), .ZN(n5036) );
  OAI211_X1 U6191 ( .C1(n5057), .C2(n5129), .A(n5037), .B(n5036), .ZN(U3058)
         );
  NAND2_X1 U6192 ( .A1(n5050), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n5041) );
  OAI22_X1 U6193 ( .A1(n5038), .A2(n5051), .B1(n5121), .B2(n6217), .ZN(n5039)
         );
  AOI21_X1 U6194 ( .B1(n5123), .B2(n5054), .A(n5039), .ZN(n5040) );
  OAI211_X1 U6195 ( .C1(n5057), .C2(n5125), .A(n5041), .B(n5040), .ZN(U3056)
         );
  NAND2_X1 U6196 ( .A1(n5050), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n5045) );
  OAI22_X1 U6197 ( .A1(n5042), .A2(n5051), .B1(n5115), .B2(n6217), .ZN(n5043)
         );
  AOI21_X1 U6198 ( .B1(n5117), .B2(n5054), .A(n5043), .ZN(n5044) );
  OAI211_X1 U6199 ( .C1(n5057), .C2(n5119), .A(n5045), .B(n5044), .ZN(U3052)
         );
  NAND2_X1 U6200 ( .A1(n5050), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n5049) );
  OAI22_X1 U6201 ( .A1(n5046), .A2(n5051), .B1(n6365), .B2(n6217), .ZN(n5047)
         );
  AOI21_X1 U6202 ( .B1(n6362), .B2(n5054), .A(n5047), .ZN(n5048) );
  OAI211_X1 U6203 ( .C1(n5057), .C2(n5141), .A(n5049), .B(n5048), .ZN(U3053)
         );
  NAND2_X1 U6204 ( .A1(n5050), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n5056) );
  OAI22_X1 U6205 ( .A1(n5052), .A2(n5051), .B1(n6390), .B2(n6217), .ZN(n5053)
         );
  AOI21_X1 U6206 ( .B1(n6386), .B2(n5054), .A(n5053), .ZN(n5055) );
  OAI211_X1 U6207 ( .C1(n5057), .C2(n5152), .A(n5056), .B(n5055), .ZN(U3057)
         );
  INV_X1 U6208 ( .A(n5059), .ZN(n5060) );
  NOR2_X1 U6209 ( .A1(n5061), .A2(n5060), .ZN(n5062) );
  XNOR2_X1 U6210 ( .A(n5058), .B(n5062), .ZN(n5196) );
  NAND2_X1 U6211 ( .A1(n5064), .A2(n5063), .ZN(n5065) );
  NAND2_X1 U6212 ( .A1(n5159), .A2(n5065), .ZN(n5955) );
  NAND2_X1 U6213 ( .A1(n6582), .A2(REIP_REG_10__SCAN_IN), .ZN(n5191) );
  AOI211_X1 U6214 ( .C1(n5068), .C2(n5067), .A(n5066), .B(n6163), .ZN(n5070)
         );
  NAND2_X1 U6215 ( .A1(n5070), .A2(n5069), .ZN(n5071) );
  OAI211_X1 U6216 ( .C1(n6584), .C2(n5955), .A(n5191), .B(n5071), .ZN(n5072)
         );
  AOI21_X1 U6217 ( .B1(n5073), .B2(INSTADDRPOINTER_REG_10__SCAN_IN), .A(n5072), 
        .ZN(n5074) );
  OAI21_X1 U6218 ( .B1(n5196), .B2(n6589), .A(n5074), .ZN(U3008) );
  XOR2_X1 U6219 ( .A(n5076), .B(n5075), .Z(n5967) );
  INV_X1 U6220 ( .A(n5967), .ZN(n5082) );
  AOI22_X1 U6221 ( .A1(n6049), .A2(n5964), .B1(EBX_REG_9__SCAN_IN), .B2(n5590), 
        .ZN(n5077) );
  OAI21_X1 U6222 ( .B1(n5082), .B2(n5589), .A(n5077), .ZN(U2850) );
  AOI22_X1 U6223 ( .A1(n6134), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .B1(n6582), 
        .B2(REIP_REG_9__SCAN_IN), .ZN(n5078) );
  OAI21_X1 U6224 ( .B1(n5965), .B2(n6143), .A(n5078), .ZN(n5079) );
  AOI21_X1 U6225 ( .B1(n5967), .B2(n6347), .A(n5079), .ZN(n5080) );
  OAI21_X1 U6226 ( .B1(n5081), .B2(n5926), .A(n5080), .ZN(U2977) );
  INV_X1 U6227 ( .A(DATAI_9_), .ZN(n6738) );
  INV_X1 U6228 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6083) );
  OAI222_X1 U6229 ( .A1(n5603), .A2(n5082), .B1(n5306), .B2(n6738), .C1(n5504), 
        .C2(n6083), .ZN(U2882) );
  INV_X1 U6230 ( .A(n5084), .ZN(n5086) );
  NOR2_X1 U6231 ( .A1(n5086), .A2(n5085), .ZN(n5087) );
  OR2_X1 U6232 ( .A1(n5083), .A2(n5087), .ZN(n5957) );
  AOI22_X1 U6233 ( .A1(n5276), .A2(DATAI_10_), .B1(EAX_REG_10__SCAN_IN), .B2(
        n6063), .ZN(n5088) );
  OAI21_X1 U6234 ( .B1(n5957), .B2(n5603), .A(n5088), .ZN(U2881) );
  INV_X1 U6235 ( .A(n5955), .ZN(n5089) );
  AOI22_X1 U6236 ( .A1(n6049), .A2(n5089), .B1(EBX_REG_10__SCAN_IN), .B2(n5590), .ZN(n5090) );
  OAI21_X1 U6237 ( .B1(n5957), .B2(n5589), .A(n5090), .ZN(U2849) );
  INV_X1 U6238 ( .A(n5091), .ZN(n5094) );
  NAND2_X1 U6239 ( .A1(n6042), .A2(EBX_REG_1__SCAN_IN), .ZN(n5092) );
  OAI211_X1 U6240 ( .C1(n5094), .C2(n6035), .A(n5093), .B(n5092), .ZN(n5095)
         );
  AOI21_X1 U6241 ( .B1(n5097), .B2(n5096), .A(n5095), .ZN(n5098) );
  OAI21_X1 U6242 ( .B1(n5281), .B2(n5099), .A(n5098), .ZN(n5101) );
  NOR2_X1 U6243 ( .A1(n6036), .A2(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5100)
         );
  AOI211_X1 U6244 ( .C1(n6003), .C2(PHYADDRPOINTER_REG_1__SCAN_IN), .A(n5101), 
        .B(n5100), .ZN(n5102) );
  OAI21_X1 U6245 ( .B1(n6038), .B2(n5103), .A(n5102), .ZN(U2826) );
  NAND2_X1 U6246 ( .A1(n6298), .A2(n6218), .ZN(n6337) );
  NAND2_X1 U6247 ( .A1(n6337), .A2(n5149), .ZN(n5104) );
  AOI21_X1 U6248 ( .B1(n5104), .B2(STATEBS16_REG_SCAN_IN), .A(n6344), .ZN(
        n5111) );
  AND2_X1 U6249 ( .A1(n5105), .A2(n4531), .ZN(n5109) );
  NOR2_X1 U6250 ( .A1(n5106), .A2(n6425), .ZN(n5107) );
  AOI22_X1 U6251 ( .A1(n5111), .A2(n5109), .B1(n6220), .B2(n5107), .ZN(n5153)
         );
  NAND2_X1 U6252 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n5108), .ZN(n6307) );
  NOR2_X1 U6253 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6307), .ZN(n5147)
         );
  INV_X1 U6254 ( .A(n5109), .ZN(n6300) );
  INV_X1 U6255 ( .A(n5147), .ZN(n5110) );
  AOI22_X1 U6256 ( .A1(n5111), .A2(n6300), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n5110), .ZN(n5112) );
  OAI211_X1 U6257 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6342), .A(n5113), .B(n5112), .ZN(n5146) );
  AOI22_X1 U6258 ( .A1(n6345), .A2(n5147), .B1(INSTQUEUE_REG_10__0__SCAN_IN), 
        .B2(n5146), .ZN(n5114) );
  OAI21_X1 U6259 ( .B1(n5115), .B2(n5149), .A(n5114), .ZN(n5116) );
  AOI21_X1 U6260 ( .B1(n5117), .B2(n6320), .A(n5116), .ZN(n5118) );
  OAI21_X1 U6261 ( .B1(n5153), .B2(n5119), .A(n5118), .ZN(U3100) );
  AOI22_X1 U6262 ( .A1(n6378), .A2(n5147), .B1(INSTQUEUE_REG_10__4__SCAN_IN), 
        .B2(n5146), .ZN(n5120) );
  OAI21_X1 U6263 ( .B1(n5121), .B2(n5149), .A(n5120), .ZN(n5122) );
  AOI21_X1 U6264 ( .B1(n5123), .B2(n6320), .A(n5122), .ZN(n5124) );
  OAI21_X1 U6265 ( .B1(n5153), .B2(n5125), .A(n5124), .ZN(U3104) );
  AOI22_X1 U6266 ( .A1(n6391), .A2(n5147), .B1(INSTQUEUE_REG_10__6__SCAN_IN), 
        .B2(n5146), .ZN(n5126) );
  OAI21_X1 U6267 ( .B1(n6329), .B2(n5149), .A(n5126), .ZN(n5127) );
  AOI21_X1 U6268 ( .B1(n6326), .B2(n6320), .A(n5127), .ZN(n5128) );
  OAI21_X1 U6269 ( .B1(n5153), .B2(n5129), .A(n5128), .ZN(U3106) );
  AOI22_X1 U6270 ( .A1(n6397), .A2(n5147), .B1(INSTQUEUE_REG_10__7__SCAN_IN), 
        .B2(n5146), .ZN(n5130) );
  OAI21_X1 U6271 ( .B1(n6338), .B2(n5149), .A(n5130), .ZN(n5131) );
  AOI21_X1 U6272 ( .B1(n6330), .B2(n6320), .A(n5131), .ZN(n5132) );
  OAI21_X1 U6273 ( .B1(n5153), .B2(n5133), .A(n5132), .ZN(U3107) );
  AOI22_X1 U6274 ( .A1(n6366), .A2(n5147), .B1(INSTQUEUE_REG_10__2__SCAN_IN), 
        .B2(n5146), .ZN(n5134) );
  OAI21_X1 U6275 ( .B1(n6371), .B2(n5149), .A(n5134), .ZN(n5135) );
  AOI21_X1 U6276 ( .B1(n6368), .B2(n6320), .A(n5135), .ZN(n5136) );
  OAI21_X1 U6277 ( .B1(n5153), .B2(n5137), .A(n5136), .ZN(U3102) );
  AOI22_X1 U6278 ( .A1(n6360), .A2(n5147), .B1(INSTQUEUE_REG_10__1__SCAN_IN), 
        .B2(n5146), .ZN(n5138) );
  OAI21_X1 U6279 ( .B1(n6365), .B2(n5149), .A(n5138), .ZN(n5139) );
  AOI21_X1 U6280 ( .B1(n6362), .B2(n6320), .A(n5139), .ZN(n5140) );
  OAI21_X1 U6281 ( .B1(n5153), .B2(n5141), .A(n5140), .ZN(U3101) );
  AOI22_X1 U6282 ( .A1(n6372), .A2(n5147), .B1(INSTQUEUE_REG_10__3__SCAN_IN), 
        .B2(n5146), .ZN(n5142) );
  OAI21_X1 U6283 ( .B1(n6319), .B2(n5149), .A(n5142), .ZN(n5143) );
  AOI21_X1 U6284 ( .B1(n6316), .B2(n6320), .A(n5143), .ZN(n5144) );
  OAI21_X1 U6285 ( .B1(n5153), .B2(n5145), .A(n5144), .ZN(U3103) );
  AOI22_X1 U6286 ( .A1(n6384), .A2(n5147), .B1(INSTQUEUE_REG_10__5__SCAN_IN), 
        .B2(n5146), .ZN(n5148) );
  OAI21_X1 U6287 ( .B1(n6390), .B2(n5149), .A(n5148), .ZN(n5150) );
  AOI21_X1 U6288 ( .B1(n6386), .B2(n6320), .A(n5150), .ZN(n5151) );
  OAI21_X1 U6289 ( .B1(n5153), .B2(n5152), .A(n5151), .ZN(U3105) );
  INV_X1 U6290 ( .A(n5154), .ZN(n5155) );
  OAI21_X1 U6291 ( .B1(n5083), .B2(n5156), .A(n5155), .ZN(n5181) );
  AOI22_X1 U6292 ( .A1(n5276), .A2(DATAI_11_), .B1(EAX_REG_11__SCAN_IN), .B2(
        n6063), .ZN(n5157) );
  OAI21_X1 U6293 ( .B1(n5181), .B2(n5603), .A(n5157), .ZN(U2880) );
  AOI21_X1 U6294 ( .B1(n5160), .B2(n5159), .A(n5158), .ZN(n6154) );
  AOI22_X1 U6295 ( .A1(n6049), .A2(n6154), .B1(EBX_REG_11__SCAN_IN), .B2(n5590), .ZN(n5161) );
  OAI21_X1 U6296 ( .B1(n5181), .B2(n5589), .A(n5161), .ZN(U2848) );
  INV_X1 U6297 ( .A(n5177), .ZN(n5172) );
  INV_X1 U6298 ( .A(EBX_REG_11__SCAN_IN), .ZN(n5167) );
  INV_X1 U6299 ( .A(n6015), .ZN(n5991) );
  AOI21_X1 U6300 ( .B1(n6003), .B2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n5991), 
        .ZN(n5166) );
  INV_X1 U6301 ( .A(REIP_REG_11__SCAN_IN), .ZN(n6499) );
  NAND2_X1 U6302 ( .A1(REIP_REG_10__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .ZN(
        n5169) );
  NOR2_X1 U6303 ( .A1(n6499), .A2(n5169), .ZN(n5241) );
  NAND2_X1 U6304 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .ZN(
        n5164) );
  NAND3_X1 U6305 ( .A1(REIP_REG_5__SCAN_IN), .A2(REIP_REG_4__SCAN_IN), .A3(
        n5162), .ZN(n5280) );
  NOR2_X1 U6306 ( .A1(n5163), .A2(n5280), .ZN(n6019) );
  NAND2_X1 U6307 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6019), .ZN(n5986) );
  OAI21_X1 U6308 ( .B1(n5164), .B2(n5986), .A(n5987), .ZN(n5984) );
  OAI21_X1 U6309 ( .B1(n6020), .B2(n5241), .A(n5984), .ZN(n5242) );
  AOI22_X1 U6310 ( .A1(n5242), .A2(REIP_REG_11__SCAN_IN), .B1(n6013), .B2(
        n6154), .ZN(n5165) );
  OAI211_X1 U6311 ( .C1(n5167), .C2(n5974), .A(n5166), .B(n5165), .ZN(n5171)
         );
  NOR2_X1 U6312 ( .A1(n5168), .A2(n6486), .ZN(n6018) );
  NAND2_X1 U6313 ( .A1(n6018), .A2(REIP_REG_5__SCAN_IN), .ZN(n5999) );
  NOR2_X1 U6314 ( .A1(n5999), .A2(n6490), .ZN(n5992) );
  NAND3_X1 U6315 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        n5992), .ZN(n5963) );
  NOR3_X1 U6316 ( .A1(REIP_REG_11__SCAN_IN), .A2(n5169), .A3(n5963), .ZN(n5170) );
  AOI211_X1 U6317 ( .C1(n5979), .C2(n5172), .A(n5171), .B(n5170), .ZN(n5173)
         );
  OAI21_X1 U6318 ( .B1(n6004), .B2(n5181), .A(n5173), .ZN(U2816) );
  NOR2_X1 U6319 ( .A1(n5175), .A2(n5176), .ZN(n5174) );
  AOI21_X1 U6320 ( .B1(n5176), .B2(n5175), .A(n5174), .ZN(n6156) );
  NAND2_X1 U6321 ( .A1(n6156), .A2(n6150), .ZN(n5180) );
  NOR2_X1 U6322 ( .A1(n5908), .A2(n6499), .ZN(n6153) );
  NOR2_X1 U6323 ( .A1(n6143), .A2(n5177), .ZN(n5178) );
  AOI211_X1 U6324 ( .C1(n6134), .C2(PHYADDRPOINTER_REG_11__SCAN_IN), .A(n6153), 
        .B(n5178), .ZN(n5179) );
  OAI211_X1 U6325 ( .C1(n5642), .C2(n5181), .A(n5180), .B(n5179), .ZN(U2975)
         );
  OAI21_X1 U6326 ( .B1(n5154), .B2(n5183), .A(n5182), .ZN(n5207) );
  INV_X1 U6327 ( .A(n5184), .ZN(n5186) );
  AOI22_X1 U6328 ( .A1(n6049), .A2(n5186), .B1(EBX_REG_12__SCAN_IN), .B2(n5590), .ZN(n5185) );
  OAI21_X1 U6329 ( .B1(n5207), .B2(n5589), .A(n5185), .ZN(U2847) );
  AOI22_X1 U6330 ( .A1(n5210), .A2(n5979), .B1(n6003), .B2(
        PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5188) );
  AOI22_X1 U6331 ( .A1(n5186), .A2(n6013), .B1(n6042), .B2(EBX_REG_12__SCAN_IN), .ZN(n5187) );
  NAND3_X1 U6332 ( .A1(n5188), .A2(n5187), .A3(n6015), .ZN(n5189) );
  INV_X1 U6333 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6500) );
  INV_X1 U6334 ( .A(n5963), .ZN(n5969) );
  AND3_X1 U6335 ( .A1(n6500), .A2(n5241), .A3(n5969), .ZN(n5243) );
  AOI211_X1 U6336 ( .C1(REIP_REG_12__SCAN_IN), .C2(n5242), .A(n5189), .B(n5243), .ZN(n5190) );
  OAI21_X1 U6337 ( .B1(n6004), .B2(n5207), .A(n5190), .ZN(U2815) );
  INV_X1 U6338 ( .A(DATAI_12_), .ZN(n6128) );
  OAI222_X1 U6339 ( .A1(n5207), .A2(n5603), .B1(n5306), .B2(n6128), .C1(n5504), 
        .C2(n3908), .ZN(U2879) );
  INV_X1 U6340 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5192) );
  OAI21_X1 U6341 ( .B1(n6148), .B2(n5192), .A(n5191), .ZN(n5194) );
  NOR2_X1 U6342 ( .A1(n5957), .A2(n5642), .ZN(n5193) );
  AOI211_X1 U6343 ( .C1(n5860), .C2(n5958), .A(n5194), .B(n5193), .ZN(n5195)
         );
  OAI21_X1 U6344 ( .B1(n5196), .B2(n5926), .A(n5195), .ZN(U2976) );
  OAI21_X1 U6345 ( .B1(n3014), .B2(n5198), .A(n3013), .ZN(n5240) );
  INV_X1 U6346 ( .A(DATAI_13_), .ZN(n6132) );
  INV_X1 U6347 ( .A(EAX_REG_13__SCAN_IN), .ZN(n6076) );
  OAI222_X1 U6348 ( .A1(n5240), .A2(n5603), .B1(n5306), .B2(n6132), .C1(n6076), 
        .C2(n5504), .ZN(U2878) );
  OR2_X1 U6349 ( .A1(n5202), .A2(n5201), .ZN(n5203) );
  NAND2_X1 U6350 ( .A1(n5200), .A2(n5203), .ZN(n5244) );
  INV_X1 U6351 ( .A(EBX_REG_13__SCAN_IN), .ZN(n5204) );
  OAI222_X1 U6352 ( .A1(n5244), .A2(n5597), .B1(n6053), .B2(n5204), .C1(n5240), 
        .C2(n5589), .ZN(U2846) );
  OAI21_X1 U6353 ( .B1(n6148), .B2(n5206), .A(n5205), .ZN(n5209) );
  NOR2_X1 U6354 ( .A1(n5207), .A2(n5642), .ZN(n5208) );
  AOI211_X1 U6355 ( .C1(n5860), .C2(n5210), .A(n5209), .B(n5208), .ZN(n5211)
         );
  OAI21_X1 U6356 ( .B1(n5926), .B2(n5212), .A(n5211), .ZN(U2974) );
  INV_X1 U6357 ( .A(n5213), .ZN(n5214) );
  AOI21_X1 U6358 ( .B1(n5216), .B2(n5215), .A(n5214), .ZN(n5259) );
  AOI21_X1 U6359 ( .B1(n5217), .B2(n5220), .A(n5266), .ZN(n5218) );
  OAI21_X1 U6360 ( .B1(n5232), .B2(n5219), .A(n5218), .ZN(n5230) );
  NOR2_X1 U6361 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n5220), .ZN(n5221)
         );
  NAND2_X1 U6362 ( .A1(n6155), .A2(n5221), .ZN(n5222) );
  NAND2_X1 U6363 ( .A1(n6582), .A2(REIP_REG_13__SCAN_IN), .ZN(n5254) );
  OAI211_X1 U6364 ( .C1(n6584), .C2(n5244), .A(n5222), .B(n5254), .ZN(n5223)
         );
  AOI21_X1 U6365 ( .B1(n5230), .B2(INSTADDRPOINTER_REG_13__SCAN_IN), .A(n5223), 
        .ZN(n5224) );
  OAI21_X1 U6366 ( .B1(n5259), .B2(n6589), .A(n5224), .ZN(U3005) );
  NAND2_X1 U6367 ( .A1(n3052), .A2(n5225), .ZN(n5226) );
  XNOR2_X1 U6368 ( .A(n5227), .B(n5226), .ZN(n5303) );
  AOI21_X1 U6369 ( .B1(n5229), .B2(n5228), .A(INSTADDRPOINTER_REG_13__SCAN_IN), 
        .ZN(n5231) );
  OAI21_X1 U6370 ( .B1(n5231), .B2(n5230), .A(INSTADDRPOINTER_REG_14__SCAN_IN), 
        .ZN(n5239) );
  INV_X1 U6371 ( .A(n5232), .ZN(n5233) );
  NOR3_X1 U6372 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5347), .A3(n5233), 
        .ZN(n5237) );
  NAND2_X1 U6373 ( .A1(n5200), .A2(n5234), .ZN(n5235) );
  NAND2_X1 U6374 ( .A1(n5263), .A2(n5235), .ZN(n5308) );
  INV_X1 U6375 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6717) );
  OAI22_X1 U6376 ( .A1(n5308), .A2(n6584), .B1(n6717), .B2(n5908), .ZN(n5236)
         );
  NOR2_X1 U6377 ( .A1(n5237), .A2(n5236), .ZN(n5238) );
  OAI211_X1 U6378 ( .C1(n5303), .C2(n6589), .A(n5239), .B(n5238), .ZN(U3004)
         );
  INV_X1 U6379 ( .A(n5240), .ZN(n5257) );
  NAND2_X1 U6380 ( .A1(REIP_REG_12__SCAN_IN), .A2(n5241), .ZN(n5279) );
  NOR3_X1 U6381 ( .A1(REIP_REG_13__SCAN_IN), .A2(n5279), .A3(n5963), .ZN(n5251) );
  OAI21_X1 U6382 ( .B1(n5243), .B2(n5242), .A(REIP_REG_13__SCAN_IN), .ZN(n5249) );
  INV_X1 U6383 ( .A(n5244), .ZN(n5245) );
  AOI22_X1 U6384 ( .A1(EBX_REG_13__SCAN_IN), .A2(n6042), .B1(n6013), .B2(n5245), .ZN(n5246) );
  OAI211_X1 U6385 ( .C1(n6031), .C2(n6744), .A(n5246), .B(n6015), .ZN(n5247)
         );
  INV_X1 U6386 ( .A(n5247), .ZN(n5248) );
  OAI211_X1 U6387 ( .C1(n6036), .C2(n5255), .A(n5249), .B(n5248), .ZN(n5250)
         );
  AOI211_X1 U6388 ( .C1(n5257), .C2(n5980), .A(n5251), .B(n5250), .ZN(n5252)
         );
  INV_X1 U6389 ( .A(n5252), .ZN(U2814) );
  NAND2_X1 U6390 ( .A1(n6134), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n5253)
         );
  OAI211_X1 U6391 ( .C1(n6143), .C2(n5255), .A(n5254), .B(n5253), .ZN(n5256)
         );
  AOI21_X1 U6392 ( .B1(n5257), .B2(n6347), .A(n5256), .ZN(n5258) );
  OAI21_X1 U6393 ( .B1(n5259), .B2(n5926), .A(n5258), .ZN(U2973) );
  NOR2_X1 U6394 ( .A1(n5261), .A2(n3050), .ZN(n5262) );
  XNOR2_X1 U6395 ( .A(n5260), .B(n5262), .ZN(n5342) );
  NOR2_X1 U6396 ( .A1(n5347), .A2(n5346), .ZN(n5270) );
  AOI21_X1 U6397 ( .B1(n5264), .B2(n5263), .A(n5350), .ZN(n5265) );
  INV_X1 U6398 ( .A(n5265), .ZN(n5304) );
  INV_X1 U6399 ( .A(n5346), .ZN(n5267) );
  INV_X1 U6400 ( .A(n5266), .ZN(n6159) );
  OAI21_X1 U6401 ( .B1(n5887), .B2(n5267), .A(n6159), .ZN(n5352) );
  NAND2_X1 U6402 ( .A1(n5352), .A2(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n5268) );
  NAND2_X1 U6403 ( .A1(n6582), .A2(REIP_REG_15__SCAN_IN), .ZN(n5336) );
  OAI211_X1 U6404 ( .C1(n6584), .C2(n5304), .A(n5268), .B(n5336), .ZN(n5269)
         );
  AOI21_X1 U6405 ( .B1(n5270), .B2(n5348), .A(n5269), .ZN(n5271) );
  OAI21_X1 U6406 ( .B1(n5342), .B2(n6589), .A(n5271), .ZN(U3003) );
  NAND2_X1 U6407 ( .A1(n5272), .A2(n5379), .ZN(n5359) );
  INV_X1 U6408 ( .A(n5379), .ZN(n5274) );
  NAND3_X1 U6409 ( .A1(n3013), .A2(n5274), .A3(n5273), .ZN(n5275) );
  AND2_X1 U6410 ( .A1(n5359), .A2(n5275), .ZN(n5301) );
  INV_X1 U6411 ( .A(n5301), .ZN(n5307) );
  AOI22_X1 U6412 ( .A1(n5276), .A2(DATAI_14_), .B1(EAX_REG_14__SCAN_IN), .B2(
        n6063), .ZN(n5277) );
  OAI21_X1 U6413 ( .B1(n5307), .B2(n5603), .A(n5277), .ZN(U2877) );
  NAND4_X1 U6414 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        REIP_REG_13__SCAN_IN), .A4(REIP_REG_6__SCAN_IN), .ZN(n5278) );
  OR3_X1 U6415 ( .A1(n5280), .A2(n5279), .A3(n5278), .ZN(n5284) );
  NOR2_X1 U6416 ( .A1(n6717), .A2(n5284), .ZN(n5292) );
  OR2_X1 U6417 ( .A1(n5292), .A2(n5529), .ZN(n5283) );
  NAND2_X1 U6418 ( .A1(n5281), .A2(n5283), .ZN(n5363) );
  AOI22_X1 U6419 ( .A1(EBX_REG_14__SCAN_IN), .A2(n6042), .B1(
        REIP_REG_14__SCAN_IN), .B2(n5363), .ZN(n5282) );
  OAI21_X1 U6420 ( .B1(n5284), .B2(n5283), .A(n5282), .ZN(n5288) );
  INV_X1 U6421 ( .A(n5299), .ZN(n5285) );
  AOI22_X1 U6422 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n6003), .B1(n5979), 
        .B2(n5285), .ZN(n5286) );
  OAI211_X1 U6423 ( .C1(n6035), .C2(n5308), .A(n5286), .B(n6015), .ZN(n5287)
         );
  AOI211_X1 U6424 ( .C1(n5301), .C2(n5980), .A(n5288), .B(n5287), .ZN(n5289)
         );
  INV_X1 U6425 ( .A(n5289), .ZN(U2813) );
  NAND2_X1 U6426 ( .A1(n5359), .A2(n5290), .ZN(n5291) );
  NAND2_X1 U6427 ( .A1(n5361), .A2(n5291), .ZN(n5339) );
  AOI22_X1 U6428 ( .A1(EBX_REG_15__SCAN_IN), .A2(n6042), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5363), .ZN(n5293) );
  OAI21_X1 U6429 ( .B1(REIP_REG_15__SCAN_IN), .B2(n5945), .A(n5293), .ZN(n5296) );
  AOI22_X1 U6430 ( .A1(PHYADDRPOINTER_REG_15__SCAN_IN), .A2(n6003), .B1(n5979), 
        .B2(n5338), .ZN(n5294) );
  OAI211_X1 U6431 ( .C1(n5304), .C2(n6035), .A(n5294), .B(n6015), .ZN(n5295)
         );
  NOR2_X1 U6432 ( .A1(n5296), .A2(n5295), .ZN(n5297) );
  OAI21_X1 U6433 ( .B1(n5339), .B2(n6004), .A(n5297), .ZN(U2812) );
  AOI22_X1 U6434 ( .A1(n6134), .A2(PHYADDRPOINTER_REG_14__SCAN_IN), .B1(n6582), 
        .B2(REIP_REG_14__SCAN_IN), .ZN(n5298) );
  OAI21_X1 U6435 ( .B1(n5299), .B2(n6143), .A(n5298), .ZN(n5300) );
  AOI21_X1 U6436 ( .B1(n5301), .B2(n6347), .A(n5300), .ZN(n5302) );
  OAI21_X1 U6437 ( .B1(n5303), .B2(n5926), .A(n5302), .ZN(U2972) );
  INV_X1 U6438 ( .A(EBX_REG_15__SCAN_IN), .ZN(n5305) );
  OAI222_X1 U6439 ( .A1(n5339), .A2(n5589), .B1(n5305), .B2(n6053), .C1(n5597), 
        .C2(n5304), .ZN(U2844) );
  OAI222_X1 U6440 ( .A1(n5339), .A2(n5603), .B1(n5306), .B2(n4356), .C1(n5504), 
        .C2(n6072), .ZN(U2876) );
  OAI222_X1 U6441 ( .A1(n5308), .A2(n5597), .B1(n6053), .B2(n3701), .C1(n5307), 
        .C2(n5589), .ZN(U2845) );
  NAND2_X1 U6442 ( .A1(n5311), .A2(n5310), .ZN(n5312) );
  AND2_X1 U6443 ( .A1(n5309), .A2(n5312), .ZN(n5850) );
  INV_X1 U6444 ( .A(n5589), .ZN(n6050) );
  INV_X1 U6445 ( .A(n5321), .ZN(n5315) );
  MUX2_X1 U6446 ( .A(n5315), .B(n5314), .S(n3029), .Z(n5383) );
  OR2_X1 U6447 ( .A1(n5313), .A2(n5383), .ZN(n5385) );
  XNOR2_X1 U6448 ( .A(n5385), .B(n5316), .ZN(n5897) );
  OAI22_X1 U6449 ( .A1(n5897), .A2(n5597), .B1(n5800), .B2(n6053), .ZN(n5317)
         );
  AOI21_X1 U6450 ( .B1(n5850), .B2(n6050), .A(n5317), .ZN(n5318) );
  INV_X1 U6451 ( .A(n5318), .ZN(U2840) );
  XNOR2_X1 U6452 ( .A(n5309), .B(n5319), .ZN(n5835) );
  MUX2_X1 U6453 ( .A(n5321), .B(n3029), .S(n5320), .Z(n5322) );
  XOR2_X1 U6454 ( .A(n5323), .B(n5322), .Z(n5888) );
  INV_X1 U6455 ( .A(n5888), .ZN(n5334) );
  INV_X1 U6456 ( .A(n5661), .ZN(n5324) );
  INV_X1 U6457 ( .A(EBX_REG_20__SCAN_IN), .ZN(n5343) );
  OAI22_X1 U6458 ( .A1(n6036), .A2(n5324), .B1(n5343), .B2(n5974), .ZN(n5333)
         );
  NAND3_X1 U6459 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .ZN(n5329) );
  INV_X1 U6460 ( .A(n5329), .ZN(n5325) );
  NOR2_X1 U6461 ( .A1(n5529), .A2(n5325), .ZN(n5326) );
  NOR2_X1 U6462 ( .A1(n5363), .A2(n5326), .ZN(n5944) );
  INV_X1 U6463 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6512) );
  NAND2_X1 U6464 ( .A1(REIP_REG_18__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .ZN(
        n5801) );
  NOR2_X1 U6465 ( .A1(n6512), .A2(n5801), .ZN(n5327) );
  OR2_X1 U6466 ( .A1(n5529), .A2(n5327), .ZN(n5328) );
  INV_X1 U6467 ( .A(n5801), .ZN(n5330) );
  AOI21_X1 U6468 ( .B1(n5330), .B2(n5802), .A(REIP_REG_20__SCAN_IN), .ZN(n5331) );
  INV_X1 U6469 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n5658) );
  OAI22_X1 U6470 ( .A1(n5523), .A2(n5331), .B1(n5658), .B2(n6031), .ZN(n5332)
         );
  AOI211_X1 U6471 ( .C1(n5334), .C2(n6013), .A(n5333), .B(n5332), .ZN(n5335)
         );
  OAI21_X1 U6472 ( .B1(n5835), .B2(n6004), .A(n5335), .ZN(U2807) );
  OAI21_X1 U6473 ( .B1(n6148), .B2(n3956), .A(n5336), .ZN(n5337) );
  AOI21_X1 U6474 ( .B1(n5860), .B2(n5338), .A(n5337), .ZN(n5341) );
  OR2_X1 U6475 ( .A1(n5339), .A2(n5642), .ZN(n5340) );
  OAI211_X1 U6476 ( .C1(n5342), .C2(n5926), .A(n5341), .B(n5340), .ZN(U2971)
         );
  OAI222_X1 U6477 ( .A1(n5835), .A2(n5589), .B1(n5343), .B2(n6053), .C1(n5597), 
        .C2(n5888), .ZN(U2839) );
  XNOR2_X1 U6478 ( .A(n2999), .B(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5345)
         );
  XNOR2_X1 U6479 ( .A(n5344), .B(n5345), .ZN(n5376) );
  AOI211_X1 U6480 ( .C1(n5863), .C2(n5348), .A(n5347), .B(n5346), .ZN(n5356)
         );
  NOR2_X1 U6481 ( .A1(n5350), .A2(n5349), .ZN(n5351) );
  OR2_X1 U6482 ( .A1(n5905), .A2(n5351), .ZN(n5378) );
  NAND2_X1 U6483 ( .A1(n5352), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5353) );
  NAND2_X1 U6484 ( .A1(n6582), .A2(REIP_REG_16__SCAN_IN), .ZN(n5372) );
  OAI211_X1 U6485 ( .C1(n6584), .C2(n5378), .A(n5353), .B(n5372), .ZN(n5354)
         );
  AOI21_X1 U6486 ( .B1(n5356), .B2(n5355), .A(n5354), .ZN(n5357) );
  OAI21_X1 U6487 ( .B1(n5376), .B2(n6589), .A(n5357), .ZN(U3002) );
  OR2_X1 U6488 ( .A1(n5359), .A2(n5358), .ZN(n5871) );
  INV_X1 U6489 ( .A(n5871), .ZN(n5360) );
  NAND2_X1 U6490 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n5946) );
  OAI21_X1 U6491 ( .B1(REIP_REG_16__SCAN_IN), .B2(REIP_REG_15__SCAN_IN), .A(
        n5946), .ZN(n5365) );
  AOI22_X1 U6492 ( .A1(EBX_REG_16__SCAN_IN), .A2(n6042), .B1(
        REIP_REG_16__SCAN_IN), .B2(n5363), .ZN(n5364) );
  OAI21_X1 U6493 ( .B1(n5945), .B2(n5365), .A(n5364), .ZN(n5369) );
  INV_X1 U6494 ( .A(n5373), .ZN(n5366) );
  AOI22_X1 U6495 ( .A1(n5366), .A2(n5979), .B1(n6003), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5367) );
  OAI211_X1 U6496 ( .C1(n5378), .C2(n6035), .A(n5367), .B(n6015), .ZN(n5368)
         );
  AOI211_X1 U6497 ( .C1(n6062), .C2(n5980), .A(n5369), .B(n5368), .ZN(n5370)
         );
  INV_X1 U6498 ( .A(n5370), .ZN(U2811) );
  NAND2_X1 U6499 ( .A1(n6134), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n5371)
         );
  OAI211_X1 U6500 ( .C1(n6143), .C2(n5373), .A(n5372), .B(n5371), .ZN(n5374)
         );
  AOI21_X1 U6501 ( .B1(n6062), .B2(n6347), .A(n5374), .ZN(n5375) );
  OAI21_X1 U6502 ( .B1(n5376), .B2(n5926), .A(n5375), .ZN(U2970) );
  INV_X1 U6503 ( .A(EBX_REG_16__SCAN_IN), .ZN(n6618) );
  INV_X1 U6504 ( .A(n6062), .ZN(n5377) );
  OAI222_X1 U6505 ( .A1(n5378), .A2(n5597), .B1(n6053), .B2(n6618), .C1(n5377), 
        .C2(n5589), .ZN(U2843) );
  AND2_X1 U6506 ( .A1(n5272), .A2(n5379), .ZN(n5381) );
  XOR2_X1 U6507 ( .A(n5382), .B(n5872), .Z(n6054) );
  INV_X1 U6508 ( .A(n6054), .ZN(n5394) );
  NAND2_X1 U6509 ( .A1(n5313), .A2(n5383), .ZN(n5384) );
  NAND2_X1 U6510 ( .A1(n5385), .A2(n5384), .ZN(n6585) );
  INV_X1 U6511 ( .A(n6585), .ZN(n5391) );
  INV_X1 U6512 ( .A(n5859), .ZN(n5387) );
  NAND2_X1 U6513 ( .A1(n6003), .A2(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5386)
         );
  OAI211_X1 U6514 ( .C1(n6036), .C2(n5387), .A(n6015), .B(n5386), .ZN(n5390)
         );
  INV_X1 U6515 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6508) );
  AOI22_X1 U6516 ( .A1(EBX_REG_18__SCAN_IN), .A2(n6042), .B1(n5802), .B2(n6508), .ZN(n5388) );
  OAI21_X1 U6517 ( .B1(n5944), .B2(n6508), .A(n5388), .ZN(n5389) );
  AOI211_X1 U6518 ( .C1(n5391), .C2(n6013), .A(n5390), .B(n5389), .ZN(n5392)
         );
  OAI21_X1 U6519 ( .B1(n5394), .B2(n6004), .A(n5392), .ZN(U2809) );
  OAI222_X1 U6520 ( .A1(n5394), .A2(n5589), .B1(n5393), .B2(n6053), .C1(n5597), 
        .C2(n6585), .ZN(U2841) );
  OR2_X1 U6521 ( .A1(n3042), .A2(n5396), .ZN(n5397) );
  NAND2_X1 U6522 ( .A1(n5395), .A2(n5397), .ZN(n5828) );
  INV_X1 U6523 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6516) );
  INV_X1 U6524 ( .A(REIP_REG_21__SCAN_IN), .ZN(n6514) );
  NOR2_X1 U6525 ( .A1(n6516), .A2(n6514), .ZN(n5784) );
  NAND4_X1 U6526 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .A3(
        REIP_REG_19__SCAN_IN), .A4(n5802), .ZN(n5783) );
  AOI211_X1 U6527 ( .C1(n6516), .C2(n6514), .A(n5784), .B(n5783), .ZN(n5401)
         );
  OAI22_X1 U6528 ( .A1(n5523), .A2(n6516), .B1(n5641), .B2(n6031), .ZN(n5400)
         );
  XOR2_X1 U6529 ( .A(n5449), .B(n5711), .Z(n5699) );
  INV_X1 U6530 ( .A(n5699), .ZN(n5596) );
  AOI22_X1 U6531 ( .A1(n5979), .A2(n5645), .B1(EBX_REG_22__SCAN_IN), .B2(n6042), .ZN(n5398) );
  OAI21_X1 U6532 ( .B1(n5596), .B2(n6035), .A(n5398), .ZN(n5399) );
  NOR3_X1 U6533 ( .A1(n5401), .A2(n5400), .A3(n5399), .ZN(n5402) );
  OAI21_X1 U6534 ( .B1(n5828), .B2(n6004), .A(n5402), .ZN(U2805) );
  AND2_X1 U6535 ( .A1(n5426), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5403)
         );
  AOI21_X1 U6536 ( .B1(n5427), .B2(EBX_REG_30__SCAN_IN), .A(n5403), .ZN(n5484)
         );
  MUX2_X1 U6537 ( .A(n5411), .B(n5486), .S(EBX_REG_25__SCAN_IN), .Z(n5405) );
  OR2_X1 U6538 ( .A1(n5427), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5404)
         );
  AND2_X1 U6539 ( .A1(n5405), .A2(n5404), .ZN(n5584) );
  NAND2_X1 U6540 ( .A1(n5584), .A2(n5585), .ZN(n5406) );
  NAND2_X1 U6541 ( .A1(n5415), .A2(n5611), .ZN(n5408) );
  INV_X1 U6542 ( .A(EBX_REG_26__SCAN_IN), .ZN(n5774) );
  NAND2_X1 U6543 ( .A1(n5420), .A2(n5774), .ZN(n5407) );
  NAND3_X1 U6544 ( .A1(n5408), .A2(n5486), .A3(n5407), .ZN(n5410) );
  NAND2_X1 U6545 ( .A1(n3029), .A2(n5774), .ZN(n5409) );
  NAND2_X1 U6546 ( .A1(n5410), .A2(n5409), .ZN(n5574) );
  MUX2_X1 U6547 ( .A(n5411), .B(n5486), .S(EBX_REG_27__SCAN_IN), .Z(n5413) );
  OR2_X1 U6548 ( .A1(n5427), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5412)
         );
  AND2_X1 U6549 ( .A1(n5413), .A2(n5412), .ZN(n5569) );
  NAND2_X1 U6550 ( .A1(n5415), .A2(n5414), .ZN(n5417) );
  INV_X1 U6551 ( .A(EBX_REG_28__SCAN_IN), .ZN(n5748) );
  NAND2_X1 U6552 ( .A1(n5420), .A2(n5748), .ZN(n5416) );
  NAND3_X1 U6553 ( .A1(n5417), .A2(n5486), .A3(n5416), .ZN(n5419) );
  NAND2_X1 U6554 ( .A1(n3029), .A2(n5748), .ZN(n5418) );
  AND2_X1 U6555 ( .A1(n5419), .A2(n5418), .ZN(n5563) );
  OR2_X1 U6556 ( .A1(n5427), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5422)
         );
  INV_X1 U6557 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5557) );
  NAND2_X1 U6558 ( .A1(n5420), .A2(n5557), .ZN(n5421) );
  NAND2_X1 U6559 ( .A1(n5422), .A2(n5421), .ZN(n5551) );
  NAND2_X1 U6560 ( .A1(n5483), .A2(n5423), .ZN(n5425) );
  INV_X1 U6561 ( .A(n3041), .ZN(n5562) );
  NOR2_X1 U6562 ( .A1(n5486), .A2(EBX_REG_29__SCAN_IN), .ZN(n5552) );
  NAND2_X1 U6563 ( .A1(n5562), .A2(n5552), .ZN(n5424) );
  NAND2_X1 U6564 ( .A1(n5425), .A2(n5424), .ZN(n5550) );
  AOI22_X1 U6565 ( .A1(n5427), .A2(EBX_REG_31__SCAN_IN), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5426), .ZN(n5428) );
  INV_X1 U6566 ( .A(n5428), .ZN(n5429) );
  OAI22_X1 U6567 ( .A1(n5534), .A2(n5597), .B1(n6053), .B2(n5431), .ZN(U2828)
         );
  INV_X1 U6568 ( .A(n5432), .ZN(n5434) );
  INV_X1 U6569 ( .A(n5435), .ZN(n5436) );
  XNOR2_X1 U6570 ( .A(n5436), .B(n5664), .ZN(n5671) );
  AND2_X1 U6571 ( .A1(n5560), .A2(n5437), .ZN(n5438) );
  INV_X1 U6572 ( .A(n5743), .ZN(n5814) );
  NOR2_X1 U6573 ( .A1(n6143), .A2(n5739), .ZN(n5441) );
  INV_X1 U6574 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5439) );
  NAND2_X1 U6575 ( .A1(n6582), .A2(REIP_REG_29__SCAN_IN), .ZN(n5667) );
  OAI21_X1 U6576 ( .B1(n6148), .B2(n5439), .A(n5667), .ZN(n5440) );
  OAI21_X1 U6577 ( .B1(n5671), .B2(n5926), .A(n5442), .ZN(U2957) );
  INV_X1 U6578 ( .A(n5446), .ZN(n5453) );
  NOR3_X1 U6579 ( .A1(n5712), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(n5447), 
        .ZN(n5452) );
  OAI21_X1 U6580 ( .B1(n5711), .B2(n5449), .A(n5448), .ZN(n5450) );
  NAND2_X1 U6581 ( .A1(n5450), .A2(n5583), .ZN(n5785) );
  NAND2_X1 U6582 ( .A1(n6582), .A2(REIP_REG_23__SCAN_IN), .ZN(n5459) );
  OAI21_X1 U6583 ( .B1(n5785), .B2(n6584), .A(n5459), .ZN(n5451) );
  AOI211_X1 U6584 ( .C1(n5453), .C2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n5452), .B(n5451), .ZN(n5454) );
  OAI21_X1 U6585 ( .B1(n5463), .B2(n6589), .A(n5454), .ZN(U2995) );
  NAND2_X1 U6586 ( .A1(n5395), .A2(n5456), .ZN(n5457) );
  AND2_X1 U6587 ( .A1(n5541), .A2(n5457), .ZN(n5825) );
  NAND2_X1 U6588 ( .A1(n6134), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5458)
         );
  OAI211_X1 U6589 ( .C1(n6143), .C2(n5460), .A(n5459), .B(n5458), .ZN(n5461)
         );
  AOI21_X1 U6590 ( .B1(n5825), .B2(n6347), .A(n5461), .ZN(n5462) );
  OAI21_X1 U6591 ( .B1(n5463), .B2(n5926), .A(n5462), .ZN(U2963) );
  INV_X1 U6592 ( .A(n5534), .ZN(n5472) );
  AND2_X1 U6593 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5690) );
  INV_X1 U6594 ( .A(n5690), .ZN(n5468) );
  AOI21_X1 U6595 ( .B1(n5464), .B2(n5468), .A(n5696), .ZN(n5672) );
  OAI21_X1 U6596 ( .B1(n5887), .B2(n5665), .A(n5672), .ZN(n5669) );
  AOI21_X1 U6597 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(
        INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5887), .ZN(n5465) );
  NOR2_X1 U6598 ( .A1(n5669), .A2(n5465), .ZN(n5481) );
  NOR2_X1 U6599 ( .A1(n5466), .A2(n6579), .ZN(n5895) );
  NAND2_X1 U6600 ( .A1(n5467), .A2(n5895), .ZN(n5875) );
  INV_X1 U6601 ( .A(n5665), .ZN(n5673) );
  NOR3_X1 U6602 ( .A1(n5663), .A2(n5673), .A3(n5664), .ZN(n5491) );
  NAND3_X1 U6603 ( .A1(n5491), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n4350), .ZN(n5469) );
  OAI211_X1 U6604 ( .C1(n5481), .C2(n4350), .A(n5470), .B(n5469), .ZN(n5471)
         );
  AOI21_X1 U6605 ( .B1(n5472), .B2(n6170), .A(n5471), .ZN(n5473) );
  OAI21_X1 U6606 ( .B1(n5474), .B2(n6589), .A(n5473), .ZN(U2987) );
  INV_X1 U6607 ( .A(n5475), .ZN(n5479) );
  INV_X1 U6608 ( .A(n5476), .ZN(n5477) );
  NAND2_X1 U6609 ( .A1(n5607), .A2(n5477), .ZN(n5478) );
  NAND2_X1 U6610 ( .A1(n5479), .A2(n5478), .ZN(n5480) );
  INV_X1 U6611 ( .A(n5481), .ZN(n5494) );
  INV_X1 U6612 ( .A(n5484), .ZN(n5482) );
  OAI21_X1 U6613 ( .B1(n5483), .B2(n3041), .A(n5482), .ZN(n5488) );
  INV_X1 U6614 ( .A(n5483), .ZN(n5485) );
  OAI211_X1 U6615 ( .C1(n5562), .C2(n5486), .A(n5485), .B(n5484), .ZN(n5487)
         );
  OAI21_X1 U6616 ( .B1(n5489), .B2(n5488), .A(n5487), .ZN(n5733) );
  NAND2_X1 U6617 ( .A1(n6582), .A2(REIP_REG_30__SCAN_IN), .ZN(n5499) );
  INV_X1 U6618 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n5490) );
  NAND2_X1 U6619 ( .A1(n5491), .A2(n5490), .ZN(n5492) );
  OAI211_X1 U6620 ( .C1(n5733), .C2(n6584), .A(n5499), .B(n5492), .ZN(n5493)
         );
  AOI21_X1 U6621 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5494), .A(n5493), 
        .ZN(n5495) );
  OAI21_X1 U6622 ( .B1(n5503), .B2(n6589), .A(n5495), .ZN(U2988) );
  XNOR2_X1 U6623 ( .A(n5498), .B(n5497), .ZN(n5811) );
  NAND2_X1 U6624 ( .A1(n5860), .A2(n5730), .ZN(n5500) );
  OAI211_X1 U6625 ( .C1(n6597), .C2(n6148), .A(n5500), .B(n5499), .ZN(n5501)
         );
  AOI21_X1 U6626 ( .B1(n5811), .B2(n6347), .A(n5501), .ZN(n5502) );
  OAI21_X1 U6627 ( .B1(n5503), .B2(n5926), .A(n5502), .ZN(U2956) );
  NAND3_X1 U6628 ( .A1(n5522), .A2(n5598), .A3(n5504), .ZN(n5506) );
  NOR2_X2 U6629 ( .A1(n6063), .A2(n3294), .ZN(n6060) );
  AOI22_X1 U6630 ( .A1(n6060), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n6063), .ZN(n5505) );
  NAND2_X1 U6631 ( .A1(n5506), .A2(n5505), .ZN(U2860) );
  INV_X1 U6632 ( .A(n5507), .ZN(n5518) );
  NOR2_X1 U6633 ( .A1(n5508), .A2(n5518), .ZN(n5509) );
  OR2_X1 U6634 ( .A1(n5520), .A2(n5509), .ZN(n5513) );
  INV_X1 U6635 ( .A(n5510), .ZN(n5511) );
  NAND2_X1 U6636 ( .A1(n5520), .A2(n5511), .ZN(n5512) );
  OAI211_X1 U6637 ( .C1(n5515), .C2(n5514), .A(n5513), .B(n5512), .ZN(n6428)
         );
  INV_X1 U6638 ( .A(n5516), .ZN(n5517) );
  OAI22_X1 U6639 ( .A1(n5520), .A2(n5519), .B1(n5518), .B2(n5517), .ZN(n5920)
         );
  AOI21_X1 U6640 ( .B1(n5521), .B2(n6469), .A(READY_N), .ZN(n6570) );
  NOR2_X1 U6641 ( .A1(n5920), .A2(n6570), .ZN(n6431) );
  NOR2_X1 U6642 ( .A1(n6431), .A2(n6451), .ZN(n5928) );
  MUX2_X1 U6643 ( .A(MORE_REG_SCAN_IN), .B(n6428), .S(n5928), .Z(U3471) );
  INV_X1 U6644 ( .A(n5522), .ZN(n5539) );
  NAND2_X1 U6645 ( .A1(REIP_REG_28__SCAN_IN), .A2(REIP_REG_27__SCAN_IN), .ZN(
        n5527) );
  INV_X1 U6646 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6519) );
  INV_X1 U6647 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6521) );
  NOR3_X1 U6648 ( .A1(n3740), .A2(n6519), .A3(n6521), .ZN(n5524) );
  NAND3_X1 U6649 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .ZN(n5526) );
  INV_X1 U6650 ( .A(n5523), .ZN(n5794) );
  AOI21_X1 U6651 ( .B1(n5525), .B2(n5526), .A(n5794), .ZN(n5791) );
  OAI21_X1 U6652 ( .B1(n5524), .B2(n6020), .A(n5791), .ZN(n5771) );
  AOI21_X1 U6653 ( .B1(n5525), .B2(n5527), .A(n5771), .ZN(n5755) );
  INV_X1 U6654 ( .A(n5755), .ZN(n5528) );
  NAND4_X1 U6655 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .A4(n5766), .ZN(n5757) );
  NOR2_X1 U6656 ( .A1(n5537), .A2(REIP_REG_29__SCAN_IN), .ZN(n5741) );
  NOR2_X1 U6657 ( .A1(n5528), .A2(n5741), .ZN(n5731) );
  OAI21_X1 U6658 ( .B1(REIP_REG_30__SCAN_IN), .B2(n5529), .A(n5731), .ZN(n5536) );
  INV_X1 U6659 ( .A(n5530), .ZN(n5532) );
  OAI22_X1 U6660 ( .A1(n6031), .A2(n5533), .B1(n5532), .B2(n5531), .ZN(n5535)
         );
  INV_X1 U6661 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6526) );
  NOR2_X1 U6662 ( .A1(n5537), .A2(n6526), .ZN(n5729) );
  INV_X1 U6663 ( .A(REIP_REG_31__SCAN_IN), .ZN(n5538) );
  AOI21_X1 U6664 ( .B1(n5542), .B2(n5541), .A(n5540), .ZN(n5635) );
  INV_X1 U6665 ( .A(n5635), .ZN(n5604) );
  OAI22_X1 U6666 ( .A1(n6036), .A2(n5633), .B1(n5543), .B2(n5974), .ZN(n5546)
         );
  OAI22_X1 U6667 ( .A1(n5791), .A2(n3740), .B1(n5544), .B2(n6031), .ZN(n5545)
         );
  AOI211_X1 U6668 ( .C1(n6013), .C2(n5591), .A(n5546), .B(n5545), .ZN(n5547)
         );
  NAND2_X1 U6669 ( .A1(n5766), .A2(n3740), .ZN(n5775) );
  OAI211_X1 U6670 ( .C1(n5604), .C2(n6004), .A(n5547), .B(n5775), .ZN(U2803)
         );
  INV_X1 U6671 ( .A(n5811), .ZN(n5549) );
  INV_X1 U6672 ( .A(EBX_REG_30__SCAN_IN), .ZN(n5548) );
  OAI222_X1 U6673 ( .A1(n5589), .A2(n5549), .B1(n5548), .B2(n6053), .C1(n5733), 
        .C2(n5597), .ZN(U2829) );
  INV_X1 U6674 ( .A(n5550), .ZN(n5556) );
  INV_X1 U6675 ( .A(n5551), .ZN(n5553) );
  AOI21_X1 U6676 ( .B1(n5553), .B2(n5486), .A(n5552), .ZN(n5554) );
  NAND2_X1 U6677 ( .A1(n3041), .A2(n5554), .ZN(n5555) );
  NAND2_X1 U6678 ( .A1(n5556), .A2(n5555), .ZN(n5742) );
  OAI222_X1 U6679 ( .A1(n5589), .A2(n5743), .B1(n5557), .B2(n6053), .C1(n5742), 
        .C2(n5597), .ZN(U2830) );
  NAND2_X1 U6680 ( .A1(n3040), .A2(n5558), .ZN(n5559) );
  INV_X1 U6681 ( .A(n5817), .ZN(n5565) );
  AOI21_X1 U6682 ( .B1(n5563), .B2(n5561), .A(n5562), .ZN(n5752) );
  AOI22_X1 U6683 ( .A1(n5752), .A2(n6049), .B1(EBX_REG_28__SCAN_IN), .B2(n5590), .ZN(n5564) );
  OAI21_X1 U6684 ( .B1(n5565), .B2(n5589), .A(n5564), .ZN(U2831) );
  NAND2_X1 U6685 ( .A1(n5566), .A2(n5567), .ZN(n5568) );
  INV_X1 U6686 ( .A(EBX_REG_27__SCAN_IN), .ZN(n5571) );
  OR2_X1 U6687 ( .A1(n5576), .A2(n5569), .ZN(n5570) );
  NAND2_X1 U6688 ( .A1(n5561), .A2(n5570), .ZN(n5758) );
  OAI222_X1 U6689 ( .A1(n5589), .A2(n5759), .B1(n6053), .B2(n5571), .C1(n5758), 
        .C2(n5597), .ZN(U2832) );
  OAI21_X1 U6690 ( .B1(n5580), .B2(n5573), .A(n5566), .ZN(n5768) );
  NOR2_X1 U6691 ( .A1(n5587), .A2(n5574), .ZN(n5575) );
  OR2_X1 U6692 ( .A1(n5576), .A2(n5575), .ZN(n5767) );
  OAI22_X1 U6693 ( .A1(n5767), .A2(n5597), .B1(n5774), .B2(n6053), .ZN(n5577)
         );
  INV_X1 U6694 ( .A(n5577), .ZN(n5578) );
  OAI21_X1 U6695 ( .B1(n5768), .B2(n5589), .A(n5578), .ZN(U2833) );
  INV_X1 U6696 ( .A(n5579), .ZN(n5582) );
  INV_X1 U6697 ( .A(n5540), .ZN(n5581) );
  AOI21_X1 U6698 ( .B1(n5582), .B2(n5581), .A(n5580), .ZN(n5843) );
  INV_X1 U6699 ( .A(n5843), .ZN(n5776) );
  INV_X1 U6700 ( .A(EBX_REG_25__SCAN_IN), .ZN(n6720) );
  INV_X1 U6701 ( .A(n5583), .ZN(n5586) );
  AOI21_X1 U6702 ( .B1(n5586), .B2(n5585), .A(n5584), .ZN(n5588) );
  OR2_X1 U6703 ( .A1(n5588), .A2(n5587), .ZN(n5877) );
  OAI222_X1 U6704 ( .A1(n5776), .A2(n5589), .B1(n6053), .B2(n6720), .C1(n5877), 
        .C2(n5597), .ZN(U2834) );
  AOI22_X1 U6705 ( .A1(n5591), .A2(n6049), .B1(EBX_REG_24__SCAN_IN), .B2(n5590), .ZN(n5592) );
  OAI21_X1 U6706 ( .B1(n5604), .B2(n5589), .A(n5592), .ZN(U2835) );
  INV_X1 U6707 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5593) );
  OAI22_X1 U6708 ( .A1(n5785), .A2(n5597), .B1(n5593), .B2(n6053), .ZN(n5594)
         );
  AOI21_X1 U6709 ( .B1(n5825), .B2(n6050), .A(n5594), .ZN(n5595) );
  INV_X1 U6710 ( .A(n5595), .ZN(U2836) );
  OAI222_X1 U6711 ( .A1(n5589), .A2(n5828), .B1(n6053), .B2(n3727), .C1(n5597), 
        .C2(n5596), .ZN(U2837) );
  AOI22_X1 U6712 ( .A1(n6064), .A2(DATAI_10_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n6063), .ZN(n5600) );
  NAND2_X1 U6713 ( .A1(n6060), .A2(DATAI_26_), .ZN(n5599) );
  OAI211_X1 U6714 ( .C1(n5768), .C2(n5603), .A(n5600), .B(n5599), .ZN(U2865)
         );
  AOI22_X1 U6715 ( .A1(n6060), .A2(DATAI_24_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n6063), .ZN(n5602) );
  NAND2_X1 U6716 ( .A1(n6064), .A2(DATAI_8_), .ZN(n5601) );
  OAI211_X1 U6717 ( .C1(n5604), .C2(n5603), .A(n5602), .B(n5601), .ZN(U2867)
         );
  NOR2_X1 U6718 ( .A1(INSTADDRPOINTER_REG_25__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5689) );
  NAND2_X1 U6719 ( .A1(n5606), .A2(n5689), .ZN(n5610) );
  NAND2_X1 U6720 ( .A1(n5608), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5609) );
  XNOR2_X1 U6721 ( .A(n5614), .B(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5680)
         );
  NAND2_X1 U6722 ( .A1(n5860), .A2(n5751), .ZN(n5615) );
  NAND2_X1 U6723 ( .A1(n6582), .A2(REIP_REG_28__SCAN_IN), .ZN(n5676) );
  OAI211_X1 U6724 ( .C1(n5747), .C2(n6148), .A(n5615), .B(n5676), .ZN(n5616)
         );
  AOI21_X1 U6725 ( .B1(n5817), .B2(n6347), .A(n5616), .ZN(n5617) );
  OAI21_X1 U6726 ( .B1(n5680), .B2(n5926), .A(n5617), .ZN(U2958) );
  INV_X1 U6727 ( .A(n5618), .ZN(n5625) );
  AOI22_X1 U6728 ( .A1(n5620), .A2(n2999), .B1(n5625), .B2(n5619), .ZN(n5621)
         );
  XNOR2_X1 U6729 ( .A(n5621), .B(n5681), .ZN(n5688) );
  INV_X1 U6730 ( .A(n5759), .ZN(n5820) );
  NAND2_X1 U6731 ( .A1(n6582), .A2(REIP_REG_27__SCAN_IN), .ZN(n5684) );
  NAND2_X1 U6732 ( .A1(n6134), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5622)
         );
  OAI211_X1 U6733 ( .C1(n6143), .C2(n5764), .A(n5684), .B(n5622), .ZN(n5623)
         );
  AOI21_X1 U6734 ( .B1(n5820), .B2(n6347), .A(n5623), .ZN(n5624) );
  OAI21_X1 U6735 ( .B1(n5688), .B2(n5926), .A(n5624), .ZN(U2959) );
  AOI21_X1 U6736 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n2999), .A(n5625), 
        .ZN(n5626) );
  XNOR2_X1 U6737 ( .A(n5607), .B(n5626), .ZN(n5698) );
  INV_X1 U6738 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n5627) );
  NAND2_X1 U6739 ( .A1(n6582), .A2(REIP_REG_26__SCAN_IN), .ZN(n5694) );
  OAI21_X1 U6740 ( .B1(n6148), .B2(n5627), .A(n5694), .ZN(n5629) );
  NOR2_X1 U6741 ( .A1(n5768), .A2(n5642), .ZN(n5628) );
  AOI211_X1 U6742 ( .C1(n5860), .C2(n5765), .A(n5629), .B(n5628), .ZN(n5630)
         );
  OAI21_X1 U6743 ( .B1(n5698), .B2(n5926), .A(n5630), .ZN(U2960) );
  AOI21_X1 U6744 ( .B1(n6134), .B2(PHYADDRPOINTER_REG_24__SCAN_IN), .A(n5631), 
        .ZN(n5632) );
  OAI21_X1 U6745 ( .B1(n5633), .B2(n6143), .A(n5632), .ZN(n5634) );
  AOI21_X1 U6746 ( .B1(n5635), .B2(n6347), .A(n5634), .ZN(n5636) );
  OAI21_X1 U6747 ( .B1(n5637), .B2(n5926), .A(n5636), .ZN(U2962) );
  AOI21_X1 U6748 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n2999), .A(n5638), 
        .ZN(n5639) );
  XNOR2_X1 U6749 ( .A(n5640), .B(n5639), .ZN(n5705) );
  NAND2_X1 U6750 ( .A1(n6582), .A2(REIP_REG_22__SCAN_IN), .ZN(n5700) );
  OAI21_X1 U6751 ( .B1(n6148), .B2(n5641), .A(n5700), .ZN(n5644) );
  NOR2_X1 U6752 ( .A1(n5828), .A2(n5642), .ZN(n5643) );
  AOI211_X1 U6753 ( .C1(n5860), .C2(n5645), .A(n5644), .B(n5643), .ZN(n5646)
         );
  OAI21_X1 U6754 ( .B1(n5705), .B2(n5926), .A(n5646), .ZN(U2964) );
  NOR2_X1 U6755 ( .A1(n5648), .A2(n5647), .ZN(n5649) );
  OR2_X1 U6756 ( .A1(n3042), .A2(n5649), .ZN(n5796) );
  OAI21_X1 U6757 ( .B1(n5651), .B2(n5650), .A(n3554), .ZN(n5707) );
  NAND2_X1 U6758 ( .A1(n5707), .A2(n6150), .ZN(n5654) );
  NOR2_X1 U6759 ( .A1(n5908), .A2(n6514), .ZN(n5714) );
  NOR2_X1 U6760 ( .A1(n6143), .A2(n5799), .ZN(n5652) );
  AOI211_X1 U6761 ( .C1(n6134), .C2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n5714), 
        .B(n5652), .ZN(n5653) );
  OAI211_X1 U6762 ( .C1(n5642), .C2(n5796), .A(n5654), .B(n5653), .ZN(U2965)
         );
  AOI21_X1 U6763 ( .B1(n5656), .B2(n5655), .A(n5443), .ZN(n5657) );
  INV_X1 U6764 ( .A(n5657), .ZN(n5889) );
  OAI22_X1 U6765 ( .A1(n6148), .A2(n5658), .B1(n5908), .B2(n6512), .ZN(n5660)
         );
  NOR2_X1 U6766 ( .A1(n5835), .A2(n5642), .ZN(n5659) );
  AOI211_X1 U6767 ( .C1(n5860), .C2(n5661), .A(n5660), .B(n5659), .ZN(n5662)
         );
  OAI21_X1 U6768 ( .B1(n5889), .B2(n5926), .A(n5662), .ZN(U2966) );
  INV_X1 U6769 ( .A(n5663), .ZN(n5682) );
  NAND3_X1 U6770 ( .A1(n5682), .A2(n5665), .A3(n5664), .ZN(n5666) );
  OAI211_X1 U6771 ( .C1(n5742), .C2(n6584), .A(n5667), .B(n5666), .ZN(n5668)
         );
  AOI21_X1 U6772 ( .B1(INSTADDRPOINTER_REG_29__SCAN_IN), .B2(n5669), .A(n5668), 
        .ZN(n5670) );
  OAI21_X1 U6773 ( .B1(n5671), .B2(n6589), .A(n5670), .ZN(U2989) );
  INV_X1 U6774 ( .A(n5672), .ZN(n5686) );
  INV_X1 U6775 ( .A(n5752), .ZN(n5677) );
  NAND3_X1 U6776 ( .A1(n5682), .A2(n5674), .A3(n5673), .ZN(n5675) );
  OAI211_X1 U6777 ( .C1(n5677), .C2(n6584), .A(n5676), .B(n5675), .ZN(n5678)
         );
  AOI21_X1 U6778 ( .B1(INSTADDRPOINTER_REG_28__SCAN_IN), .B2(n5686), .A(n5678), 
        .ZN(n5679) );
  OAI21_X1 U6779 ( .B1(n5680), .B2(n6589), .A(n5679), .ZN(U2990) );
  NAND2_X1 U6780 ( .A1(n5682), .A2(n5681), .ZN(n5683) );
  OAI211_X1 U6781 ( .C1(n5758), .C2(n6584), .A(n5684), .B(n5683), .ZN(n5685)
         );
  AOI21_X1 U6782 ( .B1(n5686), .B2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5685), 
        .ZN(n5687) );
  OAI21_X1 U6783 ( .B1(n5688), .B2(n6589), .A(n5687), .ZN(U2991) );
  INV_X1 U6784 ( .A(n5689), .ZN(n5692) );
  NOR2_X1 U6785 ( .A1(n5690), .A2(n5875), .ZN(n5691) );
  NAND2_X1 U6786 ( .A1(n5692), .A2(n5691), .ZN(n5693) );
  OAI211_X1 U6787 ( .C1(n5767), .C2(n6584), .A(n5694), .B(n5693), .ZN(n5695)
         );
  AOI21_X1 U6788 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n5696), .A(n5695), 
        .ZN(n5697) );
  OAI21_X1 U6789 ( .B1(n5698), .B2(n6589), .A(n5697), .ZN(U2992) );
  XNOR2_X1 U6790 ( .A(INSTADDRPOINTER_REG_22__SCAN_IN), .B(
        INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U6791 ( .A1(n5699), .A2(n6170), .ZN(n5701) );
  OAI211_X1 U6792 ( .C1(n5712), .C2(n5702), .A(n5701), .B(n5700), .ZN(n5703)
         );
  AOI21_X1 U6793 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5706), .A(n5703), 
        .ZN(n5704) );
  OAI21_X1 U6794 ( .B1(n5705), .B2(n6589), .A(n5704), .ZN(U2996) );
  INV_X1 U6795 ( .A(n5706), .ZN(n5718) );
  NAND2_X1 U6796 ( .A1(n5707), .A2(n6186), .ZN(n5716) );
  OR2_X1 U6797 ( .A1(n5709), .A2(n5708), .ZN(n5710) );
  AND2_X1 U6798 ( .A1(n5711), .A2(n5710), .ZN(n5808) );
  NOR2_X1 U6799 ( .A1(n5712), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5713)
         );
  AOI211_X1 U6800 ( .C1(n6170), .C2(n5808), .A(n5714), .B(n5713), .ZN(n5715)
         );
  OAI211_X1 U6801 ( .C1(n5718), .C2(n5717), .A(n5716), .B(n5715), .ZN(U2997)
         );
  OAI21_X1 U6802 ( .B1(n3035), .B2(STATEBS16_REG_SCAN_IN), .A(n6354), .ZN(
        n5719) );
  OAI22_X1 U6803 ( .A1(n5719), .A2(n6297), .B1(n4357), .B2(n5722), .ZN(n5720)
         );
  MUX2_X1 U6804 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5720), .S(n6190), 
        .Z(U3464) );
  XNOR2_X1 U6805 ( .A(n6297), .B(n5721), .ZN(n5724) );
  OAI22_X1 U6806 ( .A1(n5724), .A2(n6344), .B1(n5723), .B2(n5722), .ZN(n5725)
         );
  MUX2_X1 U6807 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B(n5725), .S(n6190), 
        .Z(U3463) );
  AND2_X1 U6808 ( .A1(n6097), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  AOI21_X1 U6809 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n5727), .A(n5726), .ZN(
        n5728) );
  INV_X1 U6810 ( .A(n5728), .ZN(U2788) );
  AOI22_X1 U6811 ( .A1(EBX_REG_30__SCAN_IN), .A2(n6042), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(n6003), .ZN(n5738) );
  INV_X1 U6812 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6533) );
  AOI22_X1 U6813 ( .A1(n5979), .A2(n5730), .B1(n5729), .B2(n6533), .ZN(n5737)
         );
  INV_X1 U6814 ( .A(n5731), .ZN(n5732) );
  AOI22_X1 U6815 ( .A1(n5811), .A2(n5980), .B1(REIP_REG_30__SCAN_IN), .B2(
        n5732), .ZN(n5736) );
  INV_X1 U6816 ( .A(n5733), .ZN(n5734) );
  NAND2_X1 U6817 ( .A1(n5734), .A2(n6013), .ZN(n5735) );
  NAND4_X1 U6818 ( .A1(n5738), .A2(n5737), .A3(n5736), .A4(n5735), .ZN(U2797)
         );
  OAI22_X1 U6819 ( .A1(n5439), .A2(n6031), .B1(n5739), .B2(n6036), .ZN(n5740)
         );
  AOI211_X1 U6820 ( .C1(EBX_REG_29__SCAN_IN), .C2(n6042), .A(n5741), .B(n5740), 
        .ZN(n5746) );
  OAI22_X1 U6821 ( .A1(n5743), .A2(n6004), .B1(n5742), .B2(n6035), .ZN(n5744)
         );
  INV_X1 U6822 ( .A(n5744), .ZN(n5745) );
  OAI211_X1 U6823 ( .C1(n5755), .C2(n6526), .A(n5746), .B(n5745), .ZN(U2798)
         );
  INV_X1 U6824 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6724) );
  INV_X1 U6825 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6523) );
  NOR3_X1 U6826 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6523), .A3(n5757), .ZN(n5750) );
  OAI22_X1 U6827 ( .A1(n5748), .A2(n5974), .B1(n5747), .B2(n6031), .ZN(n5749)
         );
  AOI211_X1 U6828 ( .C1(n5979), .C2(n5751), .A(n5750), .B(n5749), .ZN(n5754)
         );
  AOI22_X1 U6829 ( .A1(n5817), .A2(n5980), .B1(n5752), .B2(n6013), .ZN(n5753)
         );
  OAI211_X1 U6830 ( .C1(n5755), .C2(n6724), .A(n5754), .B(n5753), .ZN(U2799)
         );
  INV_X1 U6831 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5756) );
  OAI22_X1 U6832 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5757), .B1(n5756), .B2(
        n6031), .ZN(n5761) );
  OAI22_X1 U6833 ( .A1(n5759), .A2(n6004), .B1(n5758), .B2(n6035), .ZN(n5760)
         );
  NAND2_X1 U6834 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5771), .ZN(n5762) );
  OAI211_X1 U6835 ( .C1(n6036), .C2(n5764), .A(n5763), .B(n5762), .ZN(U2800)
         );
  AOI22_X1 U6836 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n6003), .B1(n5765), 
        .B2(n5979), .ZN(n5773) );
  NAND2_X1 U6837 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5766), .ZN(n5782) );
  OAI21_X1 U6838 ( .B1(n6521), .B2(n5782), .A(n6519), .ZN(n5770) );
  OAI22_X1 U6839 ( .A1(n5768), .A2(n6004), .B1(n6035), .B2(n5767), .ZN(n5769)
         );
  AOI21_X1 U6840 ( .B1(n5771), .B2(n5770), .A(n5769), .ZN(n5772) );
  OAI211_X1 U6841 ( .C1(n5774), .C2(n5974), .A(n5773), .B(n5772), .ZN(U2801)
         );
  AOI22_X1 U6842 ( .A1(EBX_REG_25__SCAN_IN), .A2(n6042), .B1(
        PHYADDRPOINTER_REG_25__SCAN_IN), .B2(n6003), .ZN(n5781) );
  AOI21_X1 U6843 ( .B1(n5791), .B2(n5775), .A(n6521), .ZN(n5778) );
  OAI22_X1 U6844 ( .A1(n5776), .A2(n6004), .B1(n6035), .B2(n5877), .ZN(n5777)
         );
  AOI211_X1 U6845 ( .C1(n5979), .C2(n5779), .A(n5778), .B(n5777), .ZN(n5780)
         );
  OAI211_X1 U6846 ( .C1(REIP_REG_25__SCAN_IN), .C2(n5782), .A(n5781), .B(n5780), .ZN(U2802) );
  INV_X1 U6847 ( .A(n5783), .ZN(n5795) );
  AOI21_X1 U6848 ( .B1(n5784), .B2(n5795), .A(REIP_REG_23__SCAN_IN), .ZN(n5790) );
  AOI22_X1 U6849 ( .A1(EBX_REG_23__SCAN_IN), .A2(n6042), .B1(
        PHYADDRPOINTER_REG_23__SCAN_IN), .B2(n6003), .ZN(n5789) );
  INV_X1 U6850 ( .A(n5785), .ZN(n5786) );
  AOI222_X1 U6851 ( .A1(n5825), .A2(n5980), .B1(n5787), .B2(n5979), .C1(n5786), 
        .C2(n6013), .ZN(n5788) );
  OAI211_X1 U6852 ( .C1(n5791), .C2(n5790), .A(n5789), .B(n5788), .ZN(U2804)
         );
  INV_X1 U6853 ( .A(EBX_REG_21__SCAN_IN), .ZN(n5810) );
  OAI22_X1 U6854 ( .A1(n5810), .A2(n5974), .B1(n5792), .B2(n6031), .ZN(n5793)
         );
  AOI221_X1 U6855 ( .B1(n5795), .B2(n6514), .C1(n5794), .C2(
        REIP_REG_21__SCAN_IN), .A(n5793), .ZN(n5798) );
  AOI22_X1 U6856 ( .A1(n5832), .A2(n5980), .B1(n6013), .B2(n5808), .ZN(n5797)
         );
  OAI211_X1 U6857 ( .C1(n5799), .C2(n6036), .A(n5798), .B(n5797), .ZN(U2806)
         );
  INV_X1 U6858 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6509) );
  OAI22_X1 U6859 ( .A1(n5944), .A2(n6509), .B1(n5800), .B2(n5974), .ZN(n5806)
         );
  OAI211_X1 U6860 ( .C1(REIP_REG_18__SCAN_IN), .C2(REIP_REG_19__SCAN_IN), .A(
        n5802), .B(n5801), .ZN(n5804) );
  AOI21_X1 U6861 ( .B1(n6003), .B2(PHYADDRPOINTER_REG_19__SCAN_IN), .A(n5991), 
        .ZN(n5803) );
  OAI211_X1 U6862 ( .C1(n5897), .C2(n6035), .A(n5804), .B(n5803), .ZN(n5805)
         );
  AOI211_X1 U6863 ( .C1(n5850), .C2(n5980), .A(n5806), .B(n5805), .ZN(n5807)
         );
  OAI21_X1 U6864 ( .B1(n5849), .B2(n6036), .A(n5807), .ZN(U2808) );
  AOI22_X1 U6865 ( .A1(n5832), .A2(n6050), .B1(n6049), .B2(n5808), .ZN(n5809)
         );
  OAI21_X1 U6866 ( .B1(n6053), .B2(n5810), .A(n5809), .ZN(U2838) );
  AOI22_X1 U6867 ( .A1(n5811), .A2(n6061), .B1(n6060), .B2(DATAI_30_), .ZN(
        n5813) );
  AOI22_X1 U6868 ( .A1(n6064), .A2(DATAI_14_), .B1(EAX_REG_30__SCAN_IN), .B2(
        n6063), .ZN(n5812) );
  NAND2_X1 U6869 ( .A1(n5813), .A2(n5812), .ZN(U2861) );
  AOI22_X1 U6870 ( .A1(n5814), .A2(n6061), .B1(n6060), .B2(DATAI_29_), .ZN(
        n5816) );
  AOI22_X1 U6871 ( .A1(n6064), .A2(DATAI_13_), .B1(EAX_REG_29__SCAN_IN), .B2(
        n6063), .ZN(n5815) );
  NAND2_X1 U6872 ( .A1(n5816), .A2(n5815), .ZN(U2862) );
  AOI22_X1 U6873 ( .A1(n5817), .A2(n6061), .B1(n6060), .B2(DATAI_28_), .ZN(
        n5819) );
  AOI22_X1 U6874 ( .A1(n6064), .A2(DATAI_12_), .B1(EAX_REG_28__SCAN_IN), .B2(
        n6063), .ZN(n5818) );
  NAND2_X1 U6875 ( .A1(n5819), .A2(n5818), .ZN(U2863) );
  AOI22_X1 U6876 ( .A1(n5820), .A2(n6061), .B1(n6060), .B2(DATAI_27_), .ZN(
        n5822) );
  AOI22_X1 U6877 ( .A1(n6064), .A2(DATAI_11_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n6063), .ZN(n5821) );
  NAND2_X1 U6878 ( .A1(n5822), .A2(n5821), .ZN(U2864) );
  AOI22_X1 U6879 ( .A1(n5843), .A2(n6061), .B1(n6060), .B2(DATAI_25_), .ZN(
        n5824) );
  AOI22_X1 U6880 ( .A1(n6064), .A2(DATAI_9_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n6063), .ZN(n5823) );
  NAND2_X1 U6881 ( .A1(n5824), .A2(n5823), .ZN(U2866) );
  AOI22_X1 U6882 ( .A1(n5825), .A2(n6061), .B1(n6060), .B2(DATAI_23_), .ZN(
        n5827) );
  AOI22_X1 U6883 ( .A1(n6064), .A2(DATAI_7_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n6063), .ZN(n5826) );
  NAND2_X1 U6884 ( .A1(n5827), .A2(n5826), .ZN(U2868) );
  INV_X1 U6885 ( .A(n5828), .ZN(n5829) );
  AOI22_X1 U6886 ( .A1(n5829), .A2(n6061), .B1(n6060), .B2(DATAI_22_), .ZN(
        n5831) );
  AOI22_X1 U6887 ( .A1(n6064), .A2(DATAI_6_), .B1(EAX_REG_22__SCAN_IN), .B2(
        n6063), .ZN(n5830) );
  NAND2_X1 U6888 ( .A1(n5831), .A2(n5830), .ZN(U2869) );
  AOI22_X1 U6889 ( .A1(n5832), .A2(n6061), .B1(n6060), .B2(DATAI_21_), .ZN(
        n5834) );
  AOI22_X1 U6890 ( .A1(n6064), .A2(DATAI_5_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n6063), .ZN(n5833) );
  NAND2_X1 U6891 ( .A1(n5834), .A2(n5833), .ZN(U2870) );
  INV_X1 U6892 ( .A(n5835), .ZN(n5836) );
  AOI22_X1 U6893 ( .A1(n5836), .A2(n6061), .B1(n6060), .B2(DATAI_20_), .ZN(
        n5838) );
  AOI22_X1 U6894 ( .A1(n6064), .A2(DATAI_4_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n6063), .ZN(n5837) );
  NAND2_X1 U6895 ( .A1(n5838), .A2(n5837), .ZN(U2871) );
  AOI22_X1 U6896 ( .A1(n5850), .A2(n6061), .B1(n6060), .B2(DATAI_19_), .ZN(
        n5840) );
  AOI22_X1 U6897 ( .A1(n6064), .A2(DATAI_3_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n6063), .ZN(n5839) );
  NAND2_X1 U6898 ( .A1(n5840), .A2(n5839), .ZN(U2872) );
  AOI22_X1 U6899 ( .A1(n6582), .A2(REIP_REG_25__SCAN_IN), .B1(n6134), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5845) );
  OAI21_X1 U6900 ( .B1(n5842), .B2(n5841), .A(n3777), .ZN(n5879) );
  AOI22_X1 U6901 ( .A1(n5843), .A2(n6347), .B1(n6150), .B2(n5879), .ZN(n5844)
         );
  OAI211_X1 U6902 ( .C1(n6143), .C2(n5846), .A(n5845), .B(n5844), .ZN(U2961)
         );
  INV_X1 U6903 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5853) );
  XNOR2_X1 U6904 ( .A(n5847), .B(n5848), .ZN(n5896) );
  INV_X1 U6905 ( .A(n5849), .ZN(n5851) );
  AOI222_X1 U6906 ( .A1(n5896), .A2(n6150), .B1(n5851), .B2(n5860), .C1(n6347), 
        .C2(n5850), .ZN(n5852) );
  NAND2_X1 U6907 ( .A1(n6582), .A2(REIP_REG_19__SCAN_IN), .ZN(n5901) );
  OAI211_X1 U6908 ( .C1(n5853), .C2(n6148), .A(n5852), .B(n5901), .ZN(U2967)
         );
  INV_X1 U6909 ( .A(n5855), .ZN(n5856) );
  INV_X1 U6910 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n6580) );
  NOR3_X1 U6911 ( .A1(n5856), .A2(n5864), .A3(n6580), .ZN(n5869) );
  NOR2_X1 U6912 ( .A1(n5857), .A2(n2999), .ZN(n5866) );
  NOR2_X1 U6913 ( .A1(n5869), .A2(n5866), .ZN(n5858) );
  XOR2_X1 U6914 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .B(n5858), .Z(n6590) );
  AOI22_X1 U6915 ( .A1(n6582), .A2(REIP_REG_18__SCAN_IN), .B1(n6134), .B2(
        PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n5862) );
  AOI22_X1 U6916 ( .A1(n6054), .A2(n6347), .B1(n5860), .B2(n5859), .ZN(n5861)
         );
  OAI211_X1 U6917 ( .C1(n6590), .C2(n5926), .A(n5862), .B(n5861), .ZN(U2968)
         );
  AOI22_X1 U6918 ( .A1(n6582), .A2(REIP_REG_17__SCAN_IN), .B1(n6134), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5874) );
  AOI21_X1 U6919 ( .B1(n5864), .B2(n5863), .A(n6580), .ZN(n5865) );
  OAI22_X1 U6920 ( .A1(n5855), .A2(n5865), .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n2999), .ZN(n5868) );
  INV_X1 U6921 ( .A(n5866), .ZN(n5867) );
  OAI21_X1 U6922 ( .B1(n5869), .B2(n5868), .A(n5867), .ZN(n5907) );
  AOI22_X1 U6923 ( .A1(n5907), .A2(n6150), .B1(n6347), .B2(n6057), .ZN(n5873)
         );
  OAI211_X1 U6924 ( .C1(n6143), .C2(n5953), .A(n5874), .B(n5873), .ZN(U2969)
         );
  INV_X1 U6925 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5882) );
  INV_X1 U6926 ( .A(n5875), .ZN(n5876) );
  AOI22_X1 U6927 ( .A1(REIP_REG_25__SCAN_IN), .A2(n6582), .B1(n5876), .B2(
        n5882), .ZN(n5881) );
  INV_X1 U6928 ( .A(n5877), .ZN(n5878) );
  AOI22_X1 U6929 ( .A1(n5879), .A2(n6186), .B1(n6170), .B2(n5878), .ZN(n5880)
         );
  OAI211_X1 U6930 ( .C1(n5883), .C2(n5882), .A(n5881), .B(n5880), .ZN(U2993)
         );
  NAND2_X1 U6931 ( .A1(n5895), .A2(n5884), .ZN(n5893) );
  OAI21_X1 U6932 ( .B1(n5885), .B2(n5887), .A(n6159), .ZN(n5910) );
  AOI21_X1 U6933 ( .B1(n6580), .B2(n5886), .A(n5910), .ZN(n6578) );
  OAI21_X1 U6934 ( .B1(INSTADDRPOINTER_REG_18__SCAN_IN), .B2(n5887), .A(n6578), 
        .ZN(n5900) );
  OAI22_X1 U6935 ( .A1(n5889), .A2(n6589), .B1(n6584), .B2(n5888), .ZN(n5890)
         );
  AOI21_X1 U6936 ( .B1(INSTADDRPOINTER_REG_20__SCAN_IN), .B2(n5900), .A(n5890), 
        .ZN(n5892) );
  NAND2_X1 U6937 ( .A1(n6582), .A2(REIP_REG_20__SCAN_IN), .ZN(n5891) );
  OAI211_X1 U6938 ( .C1(n5894), .C2(n5893), .A(n5892), .B(n5891), .ZN(U2998)
         );
  INV_X1 U6939 ( .A(n5895), .ZN(n5903) );
  INV_X1 U6940 ( .A(n5896), .ZN(n5898) );
  OAI22_X1 U6941 ( .A1(n5898), .A2(n6589), .B1(n5897), .B2(n6584), .ZN(n5899)
         );
  AOI21_X1 U6942 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5900), .A(n5899), 
        .ZN(n5902) );
  OAI211_X1 U6943 ( .C1(INSTADDRPOINTER_REG_19__SCAN_IN), .C2(n5903), .A(n5902), .B(n5901), .ZN(U2999) );
  OR2_X1 U6944 ( .A1(n5905), .A2(n5904), .ZN(n5906) );
  AND2_X1 U6945 ( .A1(n5313), .A2(n5906), .ZN(n6046) );
  AOI22_X1 U6946 ( .A1(n5907), .A2(n6186), .B1(n6170), .B2(n6046), .ZN(n5913)
         );
  INV_X1 U6947 ( .A(REIP_REG_17__SCAN_IN), .ZN(n6605) );
  NOR2_X1 U6948 ( .A1(n5908), .A2(n6605), .ZN(n5909) );
  AOI221_X1 U6949 ( .B1(n5911), .B2(n6580), .C1(n5910), .C2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .A(n5909), .ZN(n5912) );
  NAND2_X1 U6950 ( .A1(n5913), .A2(n5912), .ZN(U3001) );
  INV_X1 U6951 ( .A(n5914), .ZN(n5917) );
  NAND4_X1 U6952 ( .A1(n5917), .A2(n5916), .A3(n6542), .A4(n5915), .ZN(n5918)
         );
  OAI21_X1 U6953 ( .B1(n6552), .B2(n4523), .A(n5918), .ZN(U3455) );
  INV_X1 U6954 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6461) );
  AOI21_X1 U6955 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6461), .A(n6474), .ZN(n5923) );
  INV_X1 U6956 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5919) );
  AND2_X1 U6957 ( .A1(n6474), .A2(STATE_REG_1__SCAN_IN), .ZN(n6577) );
  AOI21_X1 U6958 ( .B1(n5923), .B2(n5919), .A(n6577), .ZN(U2789) );
  OAI21_X1 U6959 ( .B1(n5920), .B2(n6451), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5921) );
  OAI21_X1 U6960 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6452), .A(n5921), .ZN(
        U2790) );
  INV_X2 U6961 ( .A(n6577), .ZN(n6565) );
  NOR2_X1 U6962 ( .A1(STATE_REG_0__SCAN_IN), .A2(STATE_REG_2__SCAN_IN), .ZN(
        n5924) );
  OAI21_X1 U6963 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5924), .A(n6565), .ZN(n5922)
         );
  OAI21_X1 U6964 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6565), .A(n5922), .ZN(
        U2791) );
  NOR2_X1 U6965 ( .A1(n6577), .A2(n5923), .ZN(n6537) );
  OAI21_X1 U6966 ( .B1(BS16_N), .B2(n5924), .A(n6537), .ZN(n6535) );
  OAI21_X1 U6967 ( .B1(n6537), .B2(n5925), .A(n6535), .ZN(U2792) );
  OAI21_X1 U6968 ( .B1(n5928), .B2(n5927), .A(n5926), .ZN(U2793) );
  NOR4_X1 U6969 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_19__SCAN_IN), .A3(DATAWIDTH_REG_21__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n5932) );
  NOR4_X1 U6970 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(
        DATAWIDTH_REG_14__SCAN_IN), .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n5931) );
  NOR4_X1 U6971 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(
        DATAWIDTH_REG_28__SCAN_IN), .A3(DATAWIDTH_REG_29__SCAN_IN), .A4(
        DATAWIDTH_REG_31__SCAN_IN), .ZN(n5930) );
  NOR4_X1 U6972 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(
        DATAWIDTH_REG_24__SCAN_IN), .A3(DATAWIDTH_REG_25__SCAN_IN), .A4(
        DATAWIDTH_REG_26__SCAN_IN), .ZN(n5929) );
  NAND4_X1 U6973 ( .A1(n5932), .A2(n5931), .A3(n5930), .A4(n5929), .ZN(n5938)
         );
  NOR4_X1 U6974 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_6__SCAN_IN), .A4(
        DATAWIDTH_REG_2__SCAN_IN), .ZN(n5936) );
  AOI211_X1 U6975 ( .C1(DATAWIDTH_REG_1__SCAN_IN), .C2(
        DATAWIDTH_REG_0__SCAN_IN), .A(DATAWIDTH_REG_30__SCAN_IN), .B(
        DATAWIDTH_REG_8__SCAN_IN), .ZN(n5935) );
  NOR4_X1 U6976 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(DATAWIDTH_REG_10__SCAN_IN), .A3(DATAWIDTH_REG_11__SCAN_IN), .A4(DATAWIDTH_REG_12__SCAN_IN), .ZN(n5934)
         );
  NOR4_X1 U6977 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(DATAWIDTH_REG_4__SCAN_IN), 
        .A3(DATAWIDTH_REG_5__SCAN_IN), .A4(DATAWIDTH_REG_7__SCAN_IN), .ZN(
        n5933) );
  NAND4_X1 U6978 ( .A1(n5936), .A2(n5935), .A3(n5934), .A4(n5933), .ZN(n5937)
         );
  NOR2_X1 U6979 ( .A1(n5938), .A2(n5937), .ZN(n6564) );
  INV_X1 U6980 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5940) );
  NOR3_X1 U6981 ( .A1(REIP_REG_0__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .A3(DATAWIDTH_REG_0__SCAN_IN), .ZN(n5941) );
  OAI21_X1 U6982 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5941), .A(n6564), .ZN(n5939)
         );
  OAI21_X1 U6983 ( .B1(n6564), .B2(n5940), .A(n5939), .ZN(U2794) );
  INV_X1 U6984 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5943) );
  NOR2_X1 U6985 ( .A1(REIP_REG_1__SCAN_IN), .A2(DATAWIDTH_REG_1__SCAN_IN), 
        .ZN(n6558) );
  OAI21_X1 U6986 ( .B1(n5941), .B2(n6558), .A(n6564), .ZN(n5942) );
  OAI21_X1 U6987 ( .B1(n6564), .B2(n5943), .A(n5942), .ZN(U2795) );
  INV_X1 U6988 ( .A(n5944), .ZN(n5950) );
  OAI21_X1 U6989 ( .B1(n5946), .B2(n5945), .A(n6605), .ZN(n5949) );
  AOI22_X1 U6990 ( .A1(EBX_REG_17__SCAN_IN), .A2(n6042), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n6003), .ZN(n5947) );
  INV_X1 U6991 ( .A(n5947), .ZN(n5948) );
  AOI211_X1 U6992 ( .C1(n5950), .C2(n5949), .A(n5991), .B(n5948), .ZN(n5952)
         );
  AOI22_X1 U6993 ( .A1(n6057), .A2(n5980), .B1(n6013), .B2(n6046), .ZN(n5951)
         );
  OAI211_X1 U6994 ( .C1(n5953), .C2(n6036), .A(n5952), .B(n5951), .ZN(U2810)
         );
  INV_X1 U6995 ( .A(REIP_REG_10__SCAN_IN), .ZN(n6497) );
  NAND2_X1 U6996 ( .A1(REIP_REG_9__SCAN_IN), .A2(n6497), .ZN(n5962) );
  OAI21_X1 U6997 ( .B1(REIP_REG_9__SCAN_IN), .B2(n6020), .A(n5984), .ZN(n5968)
         );
  AOI22_X1 U6998 ( .A1(n6042), .A2(EBX_REG_10__SCAN_IN), .B1(
        REIP_REG_10__SCAN_IN), .B2(n5968), .ZN(n5954) );
  OAI21_X1 U6999 ( .B1(n5955), .B2(n6035), .A(n5954), .ZN(n5956) );
  AOI211_X1 U7000 ( .C1(n6003), .C2(PHYADDRPOINTER_REG_10__SCAN_IN), .A(n5991), 
        .B(n5956), .ZN(n5961) );
  INV_X1 U7001 ( .A(n5957), .ZN(n5959) );
  AOI22_X1 U7002 ( .A1(n5959), .A2(n5980), .B1(n5979), .B2(n5958), .ZN(n5960)
         );
  OAI211_X1 U7003 ( .C1(n5963), .C2(n5962), .A(n5961), .B(n5960), .ZN(U2817)
         );
  AOI22_X1 U7004 ( .A1(EBX_REG_9__SCAN_IN), .A2(n6042), .B1(
        PHYADDRPOINTER_REG_9__SCAN_IN), .B2(n6003), .ZN(n5973) );
  AOI21_X1 U7005 ( .B1(n6013), .B2(n5964), .A(n5991), .ZN(n5972) );
  INV_X1 U7006 ( .A(n5965), .ZN(n5966) );
  AOI22_X1 U7007 ( .A1(n5967), .A2(n5980), .B1(n5979), .B2(n5966), .ZN(n5971)
         );
  OAI21_X1 U7008 ( .B1(REIP_REG_9__SCAN_IN), .B2(n5969), .A(n5968), .ZN(n5970)
         );
  NAND4_X1 U7009 ( .A1(n5973), .A2(n5972), .A3(n5971), .A4(n5970), .ZN(U2818)
         );
  AOI21_X1 U7010 ( .B1(REIP_REG_7__SCAN_IN), .B2(n5992), .A(
        REIP_REG_8__SCAN_IN), .ZN(n5985) );
  OAI22_X1 U7011 ( .A1(n5976), .A2(n6035), .B1(n5975), .B2(n5974), .ZN(n5977)
         );
  AOI211_X1 U7012 ( .C1(n6003), .C2(PHYADDRPOINTER_REG_8__SCAN_IN), .A(n5991), 
        .B(n5977), .ZN(n5983) );
  AOI22_X1 U7013 ( .A1(n5981), .A2(n5980), .B1(n5979), .B2(n5978), .ZN(n5982)
         );
  OAI211_X1 U7014 ( .C1(n5985), .C2(n5984), .A(n5983), .B(n5982), .ZN(U2819)
         );
  INV_X1 U7015 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6492) );
  NAND2_X1 U7016 ( .A1(n5987), .A2(n5986), .ZN(n6009) );
  INV_X1 U7017 ( .A(n6162), .ZN(n5988) );
  AOI22_X1 U7018 ( .A1(n5988), .A2(n6013), .B1(n6042), .B2(EBX_REG_7__SCAN_IN), 
        .ZN(n5989) );
  OAI21_X1 U7019 ( .B1(n6492), .B2(n6009), .A(n5989), .ZN(n5990) );
  AOI211_X1 U7020 ( .C1(n6003), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n5991), 
        .B(n5990), .ZN(n5997) );
  INV_X1 U7021 ( .A(n5992), .ZN(n5993) );
  OAI22_X1 U7022 ( .A1(n5994), .A2(n6004), .B1(REIP_REG_7__SCAN_IN), .B2(n5993), .ZN(n5995) );
  INV_X1 U7023 ( .A(n5995), .ZN(n5996) );
  OAI211_X1 U7024 ( .C1(n5998), .C2(n6036), .A(n5997), .B(n5996), .ZN(U2820)
         );
  AND2_X1 U7025 ( .A1(n5999), .A2(n6490), .ZN(n6008) );
  AOI22_X1 U7026 ( .A1(n6000), .A2(n6013), .B1(n6042), .B2(EBX_REG_6__SCAN_IN), 
        .ZN(n6001) );
  NAND2_X1 U7027 ( .A1(n6015), .A2(n6001), .ZN(n6002) );
  AOI21_X1 U7028 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6003), .A(n6002), 
        .ZN(n6007) );
  OR2_X1 U7029 ( .A1(n6005), .A2(n6004), .ZN(n6006) );
  OAI211_X1 U7030 ( .C1(n6009), .C2(n6008), .A(n6007), .B(n6006), .ZN(n6010)
         );
  INV_X1 U7031 ( .A(n6010), .ZN(n6011) );
  OAI21_X1 U7032 ( .B1(n6012), .B2(n6036), .A(n6011), .ZN(U2821) );
  INV_X1 U7033 ( .A(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n6017) );
  AOI22_X1 U7034 ( .A1(n6014), .A2(n6013), .B1(n6042), .B2(EBX_REG_5__SCAN_IN), 
        .ZN(n6016) );
  OAI211_X1 U7035 ( .C1(n6031), .C2(n6017), .A(n6016), .B(n6015), .ZN(n6023)
         );
  INV_X1 U7036 ( .A(n6018), .ZN(n6021) );
  AOI211_X1 U7037 ( .C1(n6488), .C2(n6021), .A(n6020), .B(n6019), .ZN(n6022)
         );
  AOI211_X1 U7038 ( .C1(n6025), .C2(n6024), .A(n6023), .B(n6022), .ZN(n6026)
         );
  OAI21_X1 U7039 ( .B1(n6027), .B2(n6036), .A(n6026), .ZN(U2822) );
  INV_X1 U7040 ( .A(n6028), .ZN(n6029) );
  NAND2_X1 U7041 ( .A1(n6029), .A2(REIP_REG_2__SCAN_IN), .ZN(n6044) );
  INV_X1 U7042 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n6030) );
  OAI222_X1 U7043 ( .A1(n6035), .A2(n6034), .B1(n6033), .B2(n6032), .C1(n6031), 
        .C2(n6030), .ZN(n6041) );
  OAI22_X1 U7044 ( .A1(n6039), .A2(n6038), .B1(n6037), .B2(n6036), .ZN(n6040)
         );
  AOI211_X1 U7045 ( .C1(EBX_REG_3__SCAN_IN), .C2(n6042), .A(n6041), .B(n6040), 
        .ZN(n6043) );
  OAI221_X1 U7046 ( .B1(n6045), .B2(n6484), .C1(n6045), .C2(n6044), .A(n6043), 
        .ZN(U2824) );
  AOI22_X1 U7047 ( .A1(n6057), .A2(n6050), .B1(n6049), .B2(n6046), .ZN(n6047)
         );
  OAI21_X1 U7048 ( .B1(n6053), .B2(n6048), .A(n6047), .ZN(U2842) );
  AOI22_X1 U7049 ( .A1(n6139), .A2(n6050), .B1(n6049), .B2(n6169), .ZN(n6051)
         );
  OAI21_X1 U7050 ( .B1(n6053), .B2(n6052), .A(n6051), .ZN(U2857) );
  AOI22_X1 U7051 ( .A1(n6054), .A2(n6061), .B1(n6060), .B2(DATAI_18_), .ZN(
        n6056) );
  AOI22_X1 U7052 ( .A1(n6064), .A2(DATAI_2_), .B1(EAX_REG_18__SCAN_IN), .B2(
        n6063), .ZN(n6055) );
  NAND2_X1 U7053 ( .A1(n6056), .A2(n6055), .ZN(U2873) );
  AOI22_X1 U7054 ( .A1(n6057), .A2(n6061), .B1(n6060), .B2(DATAI_17_), .ZN(
        n6059) );
  AOI22_X1 U7055 ( .A1(n6064), .A2(DATAI_1_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n6063), .ZN(n6058) );
  NAND2_X1 U7056 ( .A1(n6059), .A2(n6058), .ZN(U2874) );
  AOI22_X1 U7057 ( .A1(n6062), .A2(n6061), .B1(n6060), .B2(DATAI_16_), .ZN(
        n6066) );
  AOI22_X1 U7058 ( .A1(n6064), .A2(DATAI_0_), .B1(EAX_REG_16__SCAN_IN), .B2(
        n6063), .ZN(n6065) );
  NAND2_X1 U7059 ( .A1(n6066), .A2(n6065), .ZN(U2875) );
  INV_X1 U7060 ( .A(UWORD_REG_12__SCAN_IN), .ZN(n6609) );
  INV_X1 U7061 ( .A(n6067), .ZN(n6069) );
  AOI22_X1 U7062 ( .A1(n6097), .A2(DATAO_REG_28__SCAN_IN), .B1(n6069), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n6068) );
  OAI21_X1 U7063 ( .B1(n6609), .B2(n6101), .A(n6068), .ZN(U2895) );
  INV_X1 U7064 ( .A(DATAO_REG_20__SCAN_IN), .ZN(n6767) );
  AOI22_X1 U7065 ( .A1(n6069), .A2(EAX_REG_20__SCAN_IN), .B1(n6569), .B2(
        UWORD_REG_4__SCAN_IN), .ZN(n6070) );
  OAI21_X1 U7066 ( .B1(n6767), .B2(n6104), .A(n6070), .ZN(U2903) );
  AOI22_X1 U7067 ( .A1(n6569), .A2(LWORD_REG_15__SCAN_IN), .B1(n6097), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n6071) );
  OAI21_X1 U7068 ( .B1(n6072), .B2(n6103), .A(n6071), .ZN(U2908) );
  AOI22_X1 U7069 ( .A1(n6569), .A2(LWORD_REG_14__SCAN_IN), .B1(n6097), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n6073) );
  OAI21_X1 U7070 ( .B1(n6074), .B2(n6103), .A(n6073), .ZN(U2909) );
  AOI22_X1 U7071 ( .A1(n6569), .A2(LWORD_REG_13__SCAN_IN), .B1(n6097), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n6075) );
  OAI21_X1 U7072 ( .B1(n6076), .B2(n6103), .A(n6075), .ZN(U2910) );
  AOI22_X1 U7073 ( .A1(n6569), .A2(LWORD_REG_12__SCAN_IN), .B1(n6097), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n6077) );
  OAI21_X1 U7074 ( .B1(n3908), .B2(n6103), .A(n6077), .ZN(U2911) );
  AOI22_X1 U7075 ( .A1(n6569), .A2(LWORD_REG_11__SCAN_IN), .B1(n6097), .B2(
        DATAO_REG_11__SCAN_IN), .ZN(n6078) );
  OAI21_X1 U7076 ( .B1(n6079), .B2(n6103), .A(n6078), .ZN(U2912) );
  AOI22_X1 U7077 ( .A1(n6569), .A2(LWORD_REG_10__SCAN_IN), .B1(n6097), .B2(
        DATAO_REG_10__SCAN_IN), .ZN(n6080) );
  OAI21_X1 U7078 ( .B1(n6081), .B2(n6103), .A(n6080), .ZN(U2913) );
  AOI22_X1 U7079 ( .A1(n6569), .A2(LWORD_REG_9__SCAN_IN), .B1(n6097), .B2(
        DATAO_REG_9__SCAN_IN), .ZN(n6082) );
  OAI21_X1 U7080 ( .B1(n6083), .B2(n6103), .A(n6082), .ZN(U2914) );
  AOI22_X1 U7081 ( .A1(n6569), .A2(LWORD_REG_8__SCAN_IN), .B1(n6097), .B2(
        DATAO_REG_8__SCAN_IN), .ZN(n6084) );
  OAI21_X1 U7082 ( .B1(n6085), .B2(n6103), .A(n6084), .ZN(U2915) );
  AOI22_X1 U7083 ( .A1(n6569), .A2(LWORD_REG_7__SCAN_IN), .B1(n6097), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n6086) );
  OAI21_X1 U7084 ( .B1(n6087), .B2(n6103), .A(n6086), .ZN(U2916) );
  AOI22_X1 U7085 ( .A1(n6569), .A2(LWORD_REG_6__SCAN_IN), .B1(n6097), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n6088) );
  OAI21_X1 U7086 ( .B1(n6730), .B2(n6103), .A(n6088), .ZN(U2917) );
  INV_X1 U7087 ( .A(LWORD_REG_5__SCAN_IN), .ZN(n6753) );
  AOI22_X1 U7088 ( .A1(EAX_REG_5__SCAN_IN), .A2(n6089), .B1(n6097), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n6090) );
  OAI21_X1 U7089 ( .B1(n6753), .B2(n6101), .A(n6090), .ZN(U2918) );
  AOI22_X1 U7090 ( .A1(n6569), .A2(LWORD_REG_4__SCAN_IN), .B1(n6097), .B2(
        DATAO_REG_4__SCAN_IN), .ZN(n6091) );
  OAI21_X1 U7091 ( .B1(n6092), .B2(n6103), .A(n6091), .ZN(U2919) );
  AOI22_X1 U7092 ( .A1(n6569), .A2(LWORD_REG_3__SCAN_IN), .B1(n6097), .B2(
        DATAO_REG_3__SCAN_IN), .ZN(n6093) );
  OAI21_X1 U7093 ( .B1(n6094), .B2(n6103), .A(n6093), .ZN(U2920) );
  AOI22_X1 U7094 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n6095), .B1(n6097), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n6096) );
  OAI21_X1 U7095 ( .B1(n3797), .B2(n6103), .A(n6096), .ZN(U2921) );
  AOI22_X1 U7096 ( .A1(n6569), .A2(LWORD_REG_1__SCAN_IN), .B1(n6097), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n6098) );
  OAI21_X1 U7097 ( .B1(n6099), .B2(n6103), .A(n6098), .ZN(U2922) );
  INV_X1 U7098 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n6715) );
  INV_X1 U7099 ( .A(LWORD_REG_0__SCAN_IN), .ZN(n6100) );
  OAI222_X1 U7100 ( .A1(n6104), .A2(n6715), .B1(n6103), .B2(n6102), .C1(n6101), 
        .C2(n6100), .ZN(U2923) );
  AOI22_X1 U7101 ( .A1(UWORD_REG_4__SCAN_IN), .A2(n6130), .B1(n6129), .B2(
        EAX_REG_20__SCAN_IN), .ZN(n6106) );
  OAI21_X1 U7102 ( .B1(n6133), .B2(n6118), .A(n6106), .ZN(U2928) );
  AOI22_X1 U7103 ( .A1(UWORD_REG_5__SCAN_IN), .A2(n6130), .B1(n6129), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n6107) );
  OAI21_X1 U7104 ( .B1(n6133), .B2(n6120), .A(n6107), .ZN(U2929) );
  AOI22_X1 U7105 ( .A1(UWORD_REG_6__SCAN_IN), .A2(n6130), .B1(n6129), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n6108) );
  OAI21_X1 U7106 ( .B1(n6133), .B2(n6122), .A(n6108), .ZN(U2930) );
  AOI22_X1 U7107 ( .A1(UWORD_REG_7__SCAN_IN), .A2(n6130), .B1(n6129), .B2(
        EAX_REG_23__SCAN_IN), .ZN(n6109) );
  OAI21_X1 U7108 ( .B1(n6133), .B2(n6124), .A(n6109), .ZN(U2931) );
  AOI22_X1 U7109 ( .A1(UWORD_REG_9__SCAN_IN), .A2(n6130), .B1(n6129), .B2(
        EAX_REG_25__SCAN_IN), .ZN(n6110) );
  OAI21_X1 U7110 ( .B1(n6133), .B2(n6738), .A(n6110), .ZN(U2933) );
  AOI22_X1 U7111 ( .A1(UWORD_REG_12__SCAN_IN), .A2(n6130), .B1(n6129), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n6111) );
  OAI21_X1 U7112 ( .B1(n6133), .B2(n6128), .A(n6111), .ZN(U2936) );
  AOI22_X1 U7113 ( .A1(UWORD_REG_13__SCAN_IN), .A2(n6130), .B1(n6129), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n6112) );
  OAI21_X1 U7114 ( .B1(n6133), .B2(n6132), .A(n6112), .ZN(U2937) );
  AOI22_X1 U7115 ( .A1(LWORD_REG_0__SCAN_IN), .A2(n6130), .B1(n6129), .B2(
        EAX_REG_0__SCAN_IN), .ZN(n6113) );
  OAI21_X1 U7116 ( .B1(n6133), .B2(n4323), .A(n6113), .ZN(U2939) );
  AOI22_X1 U7117 ( .A1(LWORD_REG_1__SCAN_IN), .A2(n6130), .B1(n6129), .B2(
        EAX_REG_1__SCAN_IN), .ZN(n6114) );
  OAI21_X1 U7118 ( .B1(n6133), .B2(n4319), .A(n6114), .ZN(U2940) );
  AOI22_X1 U7119 ( .A1(LWORD_REG_2__SCAN_IN), .A2(n6125), .B1(n6129), .B2(
        EAX_REG_2__SCAN_IN), .ZN(n6115) );
  OAI21_X1 U7120 ( .B1(n6133), .B2(n4317), .A(n6115), .ZN(U2941) );
  AOI22_X1 U7121 ( .A1(LWORD_REG_3__SCAN_IN), .A2(n6125), .B1(n6129), .B2(
        EAX_REG_3__SCAN_IN), .ZN(n6116) );
  OAI21_X1 U7122 ( .B1(n6133), .B2(n4321), .A(n6116), .ZN(U2942) );
  AOI22_X1 U7123 ( .A1(LWORD_REG_4__SCAN_IN), .A2(n6125), .B1(n6129), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n6117) );
  OAI21_X1 U7124 ( .B1(n6133), .B2(n6118), .A(n6117), .ZN(U2943) );
  AOI22_X1 U7125 ( .A1(LWORD_REG_5__SCAN_IN), .A2(n6125), .B1(n6129), .B2(
        EAX_REG_5__SCAN_IN), .ZN(n6119) );
  OAI21_X1 U7126 ( .B1(n6133), .B2(n6120), .A(n6119), .ZN(U2944) );
  AOI22_X1 U7127 ( .A1(LWORD_REG_6__SCAN_IN), .A2(n6125), .B1(n6129), .B2(
        EAX_REG_6__SCAN_IN), .ZN(n6121) );
  OAI21_X1 U7128 ( .B1(n6133), .B2(n6122), .A(n6121), .ZN(U2945) );
  AOI22_X1 U7129 ( .A1(LWORD_REG_7__SCAN_IN), .A2(n6125), .B1(n6129), .B2(
        EAX_REG_7__SCAN_IN), .ZN(n6123) );
  OAI21_X1 U7130 ( .B1(n6133), .B2(n6124), .A(n6123), .ZN(U2946) );
  AOI22_X1 U7131 ( .A1(LWORD_REG_9__SCAN_IN), .A2(n6125), .B1(n6129), .B2(
        EAX_REG_9__SCAN_IN), .ZN(n6126) );
  OAI21_X1 U7132 ( .B1(n6133), .B2(n6738), .A(n6126), .ZN(U2948) );
  AOI22_X1 U7133 ( .A1(LWORD_REG_12__SCAN_IN), .A2(n6130), .B1(n6129), .B2(
        EAX_REG_12__SCAN_IN), .ZN(n6127) );
  OAI21_X1 U7134 ( .B1(n6133), .B2(n6128), .A(n6127), .ZN(U2951) );
  AOI22_X1 U7135 ( .A1(LWORD_REG_13__SCAN_IN), .A2(n6130), .B1(n6129), .B2(
        EAX_REG_13__SCAN_IN), .ZN(n6131) );
  OAI21_X1 U7136 ( .B1(n6133), .B2(n6132), .A(n6131), .ZN(U2952) );
  AOI22_X1 U7137 ( .A1(n6582), .A2(REIP_REG_2__SCAN_IN), .B1(n6134), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n6141) );
  NAND2_X1 U7138 ( .A1(n6136), .A2(n6135), .ZN(n6137) );
  XOR2_X1 U7139 ( .A(n6138), .B(n6137), .Z(n6174) );
  AOI22_X1 U7140 ( .A1(n6174), .A2(n6150), .B1(n6139), .B2(n6347), .ZN(n6140)
         );
  OAI211_X1 U7141 ( .C1(n6143), .C2(n6142), .A(n6141), .B(n6140), .ZN(U2984)
         );
  OAI21_X1 U7142 ( .B1(n6144), .B2(INSTADDRPOINTER_REG_0__SCAN_IN), .A(n3476), 
        .ZN(n6145) );
  INV_X1 U7143 ( .A(n6145), .ZN(n6185) );
  INV_X1 U7144 ( .A(n6146), .ZN(n6147) );
  INV_X1 U7145 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n6737) );
  AOI21_X1 U7146 ( .B1(n6148), .B2(n6147), .A(n6737), .ZN(n6149) );
  AOI21_X1 U7147 ( .B1(n6185), .B2(n6150), .A(n6149), .ZN(n6151) );
  NAND2_X1 U7148 ( .A1(n6582), .A2(REIP_REG_0__SCAN_IN), .ZN(n6181) );
  OAI211_X1 U7149 ( .C1(n6152), .C2(n5642), .A(n6151), .B(n6181), .ZN(U2986)
         );
  AOI21_X1 U7150 ( .B1(n6170), .B2(n6154), .A(n6153), .ZN(n6158) );
  AOI22_X1 U7151 ( .A1(n6156), .A2(n6186), .B1(n6155), .B2(n6770), .ZN(n6157)
         );
  OAI211_X1 U7152 ( .C1(n6159), .C2(n6770), .A(n6158), .B(n6157), .ZN(U3007)
         );
  INV_X1 U7153 ( .A(n6160), .ZN(n6168) );
  OAI21_X1 U7154 ( .B1(n6584), .B2(n6162), .A(n6161), .ZN(n6165) );
  NOR2_X1 U7155 ( .A1(n6163), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n6164)
         );
  AOI211_X1 U7156 ( .C1(n6166), .C2(n6186), .A(n6165), .B(n6164), .ZN(n6167)
         );
  OAI21_X1 U7157 ( .B1(n6168), .B2(n6723), .A(n6167), .ZN(U3011) );
  AOI22_X1 U7158 ( .A1(n6170), .A2(n6169), .B1(n6582), .B2(REIP_REG_2__SCAN_IN), .ZN(n6180) );
  NAND3_X1 U7159 ( .A1(n6171), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n6172) );
  NAND2_X1 U7160 ( .A1(n6173), .A2(n6172), .ZN(n6175) );
  AOI22_X1 U7161 ( .A1(n6175), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .B1(n6186), 
        .B2(n6174), .ZN(n6179) );
  NAND3_X1 U7162 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n6176), .A3(n3657), 
        .ZN(n6177) );
  NAND4_X1 U7163 ( .A1(n6180), .A2(n6179), .A3(n6178), .A4(n6177), .ZN(U3016)
         );
  OAI211_X1 U7164 ( .C1(n6584), .C2(n6183), .A(n6182), .B(n6181), .ZN(n6184)
         );
  AOI21_X1 U7165 ( .B1(n6186), .B2(n6185), .A(n6184), .ZN(n6187) );
  OAI21_X1 U7166 ( .B1(n6189), .B2(n6188), .A(n6187), .ZN(U3018) );
  NOR2_X1 U7167 ( .A1(n6191), .A2(n6190), .ZN(U3019) );
  AOI22_X1 U7168 ( .A1(n6361), .A2(n6201), .B1(n6360), .B2(n6200), .ZN(n6193)
         );
  AOI22_X1 U7169 ( .A1(n6203), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .B1(n6362), 
        .B2(n6202), .ZN(n6192) );
  OAI211_X1 U7170 ( .C1(n6365), .C2(n6406), .A(n6193), .B(n6192), .ZN(U3021)
         );
  AOI22_X1 U7171 ( .A1(n6367), .A2(n6201), .B1(n6366), .B2(n6200), .ZN(n6195)
         );
  AOI22_X1 U7172 ( .A1(n6203), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n6368), 
        .B2(n6202), .ZN(n6194) );
  OAI211_X1 U7173 ( .C1(n6371), .C2(n6406), .A(n6195), .B(n6194), .ZN(U3022)
         );
  AOI22_X1 U7174 ( .A1(n6373), .A2(n6201), .B1(n6372), .B2(n6200), .ZN(n6197)
         );
  AOI22_X1 U7175 ( .A1(n6203), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n6316), 
        .B2(n6202), .ZN(n6196) );
  OAI211_X1 U7176 ( .C1(n6319), .C2(n6406), .A(n6197), .B(n6196), .ZN(U3023)
         );
  AOI22_X1 U7177 ( .A1(n6385), .A2(n6201), .B1(n6384), .B2(n6200), .ZN(n6199)
         );
  AOI22_X1 U7178 ( .A1(n6203), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n6386), 
        .B2(n6202), .ZN(n6198) );
  OAI211_X1 U7179 ( .C1(n6390), .C2(n6406), .A(n6199), .B(n6198), .ZN(U3025)
         );
  AOI22_X1 U7180 ( .A1(n6400), .A2(n6201), .B1(n6397), .B2(n6200), .ZN(n6205)
         );
  AOI22_X1 U7181 ( .A1(n6203), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n6330), 
        .B2(n6202), .ZN(n6204) );
  OAI211_X1 U7182 ( .C1(n6338), .C2(n6406), .A(n6205), .B(n6204), .ZN(U3027)
         );
  INV_X1 U7183 ( .A(n6206), .ZN(n6212) );
  AOI22_X1 U7184 ( .A1(n6345), .A2(n6212), .B1(n6356), .B2(n6211), .ZN(n6208)
         );
  AOI22_X1 U7185 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6214), .B1(n6346), 
        .B2(n6213), .ZN(n6207) );
  OAI211_X1 U7186 ( .C1(n6359), .C2(n6217), .A(n6208), .B(n6207), .ZN(U3044)
         );
  AOI22_X1 U7187 ( .A1(n6378), .A2(n6212), .B1(n6380), .B2(n6211), .ZN(n6210)
         );
  AOI22_X1 U7188 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6214), .B1(n6379), 
        .B2(n6213), .ZN(n6209) );
  OAI211_X1 U7189 ( .C1(n6383), .C2(n6217), .A(n6210), .B(n6209), .ZN(U3048)
         );
  AOI22_X1 U7190 ( .A1(n6391), .A2(n6212), .B1(n6393), .B2(n6211), .ZN(n6216)
         );
  AOI22_X1 U7191 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6214), .B1(n6392), 
        .B2(n6213), .ZN(n6215) );
  OAI211_X1 U7192 ( .C1(n6396), .C2(n6217), .A(n6216), .B(n6215), .ZN(U3050)
         );
  NAND2_X1 U7193 ( .A1(n6219), .A2(n6218), .ZN(n6277) );
  NAND3_X1 U7194 ( .A1(n6221), .A2(n6220), .A3(n6425), .ZN(n6222) );
  OAI21_X1 U7195 ( .B1(n6223), .B2(n6254), .A(n6222), .ZN(n6247) );
  INV_X1 U7196 ( .A(n6257), .ZN(n6259) );
  NOR2_X1 U7197 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6259), .ZN(n6246)
         );
  AOI22_X1 U7198 ( .A1(n6346), .A2(n6247), .B1(n6345), .B2(n6246), .ZN(n6231)
         );
  NOR2_X1 U7199 ( .A1(n6248), .A2(n6344), .ZN(n6224) );
  AOI21_X1 U7200 ( .B1(n6224), .B2(n6277), .A(n6350), .ZN(n6229) );
  INV_X1 U7201 ( .A(n6246), .ZN(n6227) );
  AOI211_X1 U7202 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6227), .A(n6226), .B(
        n6225), .ZN(n6228) );
  OAI211_X1 U7203 ( .C1(n6340), .C2(n6229), .A(n6228), .B(n6425), .ZN(n6249)
         );
  AOI22_X1 U7204 ( .A1(n6249), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n6356), 
        .B2(n6248), .ZN(n6230) );
  OAI211_X1 U7205 ( .C1(n6359), .C2(n6277), .A(n6231), .B(n6230), .ZN(U3068)
         );
  AOI22_X1 U7206 ( .A1(n6361), .A2(n6247), .B1(n6360), .B2(n6246), .ZN(n6233)
         );
  AOI22_X1 U7207 ( .A1(n6249), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n6264), 
        .B2(n6248), .ZN(n6232) );
  OAI211_X1 U7208 ( .C1(n6267), .C2(n6277), .A(n6233), .B(n6232), .ZN(U3069)
         );
  AOI22_X1 U7209 ( .A1(n6367), .A2(n6247), .B1(n6366), .B2(n6246), .ZN(n6235)
         );
  AOI22_X1 U7210 ( .A1(n6249), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n6312), 
        .B2(n6248), .ZN(n6234) );
  OAI211_X1 U7211 ( .C1(n6315), .C2(n6277), .A(n6235), .B(n6234), .ZN(U3070)
         );
  AOI22_X1 U7212 ( .A1(n6373), .A2(n6247), .B1(n6372), .B2(n6246), .ZN(n6237)
         );
  AOI22_X1 U7213 ( .A1(n6249), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n6374), 
        .B2(n6248), .ZN(n6236) );
  OAI211_X1 U7214 ( .C1(n6377), .C2(n6277), .A(n6237), .B(n6236), .ZN(U3071)
         );
  AOI22_X1 U7215 ( .A1(n6379), .A2(n6247), .B1(n6378), .B2(n6246), .ZN(n6239)
         );
  AOI22_X1 U7216 ( .A1(n6249), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n6380), 
        .B2(n6248), .ZN(n6238) );
  OAI211_X1 U7217 ( .C1(n6383), .C2(n6277), .A(n6239), .B(n6238), .ZN(U3072)
         );
  AOI22_X1 U7218 ( .A1(n6385), .A2(n6247), .B1(n6384), .B2(n6246), .ZN(n6242)
         );
  AOI22_X1 U7219 ( .A1(n6249), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n6240), 
        .B2(n6248), .ZN(n6241) );
  OAI211_X1 U7220 ( .C1(n6243), .C2(n6277), .A(n6242), .B(n6241), .ZN(U3073)
         );
  AOI22_X1 U7221 ( .A1(n6392), .A2(n6247), .B1(n6391), .B2(n6246), .ZN(n6245)
         );
  AOI22_X1 U7222 ( .A1(n6249), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n6393), 
        .B2(n6248), .ZN(n6244) );
  OAI211_X1 U7223 ( .C1(n6396), .C2(n6277), .A(n6245), .B(n6244), .ZN(U3074)
         );
  AOI22_X1 U7224 ( .A1(n6400), .A2(n6247), .B1(n6397), .B2(n6246), .ZN(n6251)
         );
  AOI22_X1 U7225 ( .A1(n6249), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n6402), 
        .B2(n6248), .ZN(n6250) );
  OAI211_X1 U7226 ( .C1(n6407), .C2(n6277), .A(n6251), .B(n6250), .ZN(U3075)
         );
  INV_X1 U7227 ( .A(n6252), .ZN(n6281) );
  INV_X1 U7228 ( .A(n6277), .ZN(n6280) );
  AOI22_X1 U7229 ( .A1(n6345), .A2(n6281), .B1(n6356), .B2(n6280), .ZN(n6263)
         );
  NOR3_X1 U7230 ( .A1(n6254), .A2(n6412), .A3(n6253), .ZN(n6255) );
  NOR2_X1 U7231 ( .A1(n6255), .A2(n6281), .ZN(n6261) );
  NAND3_X1 U7232 ( .A1(n6354), .A2(n6261), .A3(n6258), .ZN(n6256) );
  OAI211_X1 U7233 ( .C1(n6257), .C2(n6354), .A(n6353), .B(n6256), .ZN(n6283)
         );
  NAND2_X1 U7234 ( .A1(n6354), .A2(n6258), .ZN(n6260) );
  OAI22_X1 U7235 ( .A1(n6261), .A2(n6260), .B1(n6342), .B2(n6259), .ZN(n6282)
         );
  AOI22_X1 U7236 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6283), .B1(n6346), 
        .B2(n6282), .ZN(n6262) );
  OAI211_X1 U7237 ( .C1(n6359), .C2(n6295), .A(n6263), .B(n6262), .ZN(U3076)
         );
  AOI22_X1 U7238 ( .A1(n6360), .A2(n6281), .B1(n6264), .B2(n6280), .ZN(n6266)
         );
  AOI22_X1 U7239 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6283), .B1(n6361), 
        .B2(n6282), .ZN(n6265) );
  OAI211_X1 U7240 ( .C1(n6267), .C2(n6295), .A(n6266), .B(n6265), .ZN(U3077)
         );
  AOI22_X1 U7241 ( .A1(n6366), .A2(n6281), .B1(n6368), .B2(n6274), .ZN(n6269)
         );
  AOI22_X1 U7242 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6283), .B1(n6367), 
        .B2(n6282), .ZN(n6268) );
  OAI211_X1 U7243 ( .C1(n6371), .C2(n6277), .A(n6269), .B(n6268), .ZN(U3078)
         );
  AOI22_X1 U7244 ( .A1(n6372), .A2(n6281), .B1(n6316), .B2(n6274), .ZN(n6271)
         );
  AOI22_X1 U7245 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6283), .B1(n6373), 
        .B2(n6282), .ZN(n6270) );
  OAI211_X1 U7246 ( .C1(n6319), .C2(n6277), .A(n6271), .B(n6270), .ZN(U3079)
         );
  AOI22_X1 U7247 ( .A1(n6378), .A2(n6281), .B1(n6380), .B2(n6280), .ZN(n6273)
         );
  AOI22_X1 U7248 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6283), .B1(n6379), 
        .B2(n6282), .ZN(n6272) );
  OAI211_X1 U7249 ( .C1(n6383), .C2(n6295), .A(n6273), .B(n6272), .ZN(U3080)
         );
  AOI22_X1 U7250 ( .A1(n6384), .A2(n6281), .B1(n6386), .B2(n6274), .ZN(n6276)
         );
  AOI22_X1 U7251 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6283), .B1(n6385), 
        .B2(n6282), .ZN(n6275) );
  OAI211_X1 U7252 ( .C1(n6390), .C2(n6277), .A(n6276), .B(n6275), .ZN(U3081)
         );
  AOI22_X1 U7253 ( .A1(n6391), .A2(n6281), .B1(n6393), .B2(n6280), .ZN(n6279)
         );
  AOI22_X1 U7254 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6283), .B1(n6392), 
        .B2(n6282), .ZN(n6278) );
  OAI211_X1 U7255 ( .C1(n6396), .C2(n6295), .A(n6279), .B(n6278), .ZN(U3082)
         );
  AOI22_X1 U7256 ( .A1(n6397), .A2(n6281), .B1(n6402), .B2(n6280), .ZN(n6285)
         );
  AOI22_X1 U7257 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6283), .B1(n6400), 
        .B2(n6282), .ZN(n6284) );
  OAI211_X1 U7258 ( .C1(n6407), .C2(n6295), .A(n6285), .B(n6284), .ZN(U3083)
         );
  INV_X1 U7259 ( .A(n6286), .ZN(n6290) );
  AOI22_X1 U7260 ( .A1(n6361), .A2(n6290), .B1(n6360), .B2(n6289), .ZN(n6288)
         );
  AOI22_X1 U7261 ( .A1(n6292), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n6362), 
        .B2(n6291), .ZN(n6287) );
  OAI211_X1 U7262 ( .C1(n6365), .C2(n6295), .A(n6288), .B(n6287), .ZN(U3085)
         );
  AOI22_X1 U7263 ( .A1(n6373), .A2(n6290), .B1(n6372), .B2(n6289), .ZN(n6294)
         );
  AOI22_X1 U7264 ( .A1(n6292), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n6316), 
        .B2(n6291), .ZN(n6293) );
  OAI211_X1 U7265 ( .C1(n6319), .C2(n6295), .A(n6294), .B(n6293), .ZN(U3087)
         );
  NOR2_X1 U7266 ( .A1(n6425), .A2(n6296), .ZN(n6332) );
  AOI22_X1 U7267 ( .A1(n6345), .A2(n6332), .B1(n6320), .B2(n6356), .ZN(n6309)
         );
  INV_X1 U7268 ( .A(n6307), .ZN(n6303) );
  NAND2_X1 U7269 ( .A1(n6298), .A2(n6297), .ZN(n6305) );
  INV_X1 U7270 ( .A(n6332), .ZN(n6299) );
  OAI21_X1 U7271 ( .B1(n6300), .B2(n6412), .A(n6299), .ZN(n6304) );
  INV_X1 U7272 ( .A(n6304), .ZN(n6301) );
  NAND3_X1 U7273 ( .A1(n6305), .A2(n6354), .A3(n6301), .ZN(n6302) );
  OAI211_X1 U7274 ( .C1(n6354), .C2(n6303), .A(n6302), .B(n6353), .ZN(n6334)
         );
  NAND3_X1 U7275 ( .A1(n6305), .A2(n6354), .A3(n6304), .ZN(n6306) );
  OAI21_X1 U7276 ( .B1(n6307), .B2(n6342), .A(n6306), .ZN(n6333) );
  AOI22_X1 U7277 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6334), .B1(n6346), 
        .B2(n6333), .ZN(n6308) );
  OAI211_X1 U7278 ( .C1(n6359), .C2(n6323), .A(n6309), .B(n6308), .ZN(U3108)
         );
  AOI22_X1 U7279 ( .A1(n6360), .A2(n6332), .B1(n6331), .B2(n6362), .ZN(n6311)
         );
  AOI22_X1 U7280 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6334), .B1(n6361), 
        .B2(n6333), .ZN(n6310) );
  OAI211_X1 U7281 ( .C1(n6365), .C2(n6337), .A(n6311), .B(n6310), .ZN(U3109)
         );
  AOI22_X1 U7282 ( .A1(n6366), .A2(n6332), .B1(n6320), .B2(n6312), .ZN(n6314)
         );
  AOI22_X1 U7283 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6334), .B1(n6367), 
        .B2(n6333), .ZN(n6313) );
  OAI211_X1 U7284 ( .C1(n6315), .C2(n6323), .A(n6314), .B(n6313), .ZN(U3110)
         );
  AOI22_X1 U7285 ( .A1(n6372), .A2(n6332), .B1(n6331), .B2(n6316), .ZN(n6318)
         );
  AOI22_X1 U7286 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6334), .B1(n6373), 
        .B2(n6333), .ZN(n6317) );
  OAI211_X1 U7287 ( .C1(n6319), .C2(n6337), .A(n6318), .B(n6317), .ZN(U3111)
         );
  AOI22_X1 U7288 ( .A1(n6378), .A2(n6332), .B1(n6320), .B2(n6380), .ZN(n6322)
         );
  AOI22_X1 U7289 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6334), .B1(n6379), 
        .B2(n6333), .ZN(n6321) );
  OAI211_X1 U7290 ( .C1(n6383), .C2(n6323), .A(n6322), .B(n6321), .ZN(U3112)
         );
  AOI22_X1 U7291 ( .A1(n6384), .A2(n6332), .B1(n6331), .B2(n6386), .ZN(n6325)
         );
  AOI22_X1 U7292 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6334), .B1(n6385), 
        .B2(n6333), .ZN(n6324) );
  OAI211_X1 U7293 ( .C1(n6390), .C2(n6337), .A(n6325), .B(n6324), .ZN(U3113)
         );
  AOI22_X1 U7294 ( .A1(n6391), .A2(n6332), .B1(n6331), .B2(n6326), .ZN(n6328)
         );
  AOI22_X1 U7295 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6334), .B1(n6392), 
        .B2(n6333), .ZN(n6327) );
  OAI211_X1 U7296 ( .C1(n6329), .C2(n6337), .A(n6328), .B(n6327), .ZN(U3114)
         );
  AOI22_X1 U7297 ( .A1(n6397), .A2(n6332), .B1(n6331), .B2(n6330), .ZN(n6336)
         );
  AOI22_X1 U7298 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6334), .B1(n6400), 
        .B2(n6333), .ZN(n6335) );
  OAI211_X1 U7299 ( .C1(n6338), .C2(n6337), .A(n6336), .B(n6335), .ZN(U3115)
         );
  INV_X1 U7300 ( .A(n6339), .ZN(n6398) );
  AOI21_X1 U7301 ( .B1(n6341), .B2(n6340), .A(n6398), .ZN(n6349) );
  OAI22_X1 U7302 ( .A1(n6349), .A2(n6344), .B1(n6343), .B2(n6342), .ZN(n6399)
         );
  AOI22_X1 U7303 ( .A1(n6346), .A2(n6399), .B1(n6398), .B2(n6345), .ZN(n6358)
         );
  AND2_X1 U7304 ( .A1(n6348), .A2(n6347), .ZN(n6351) );
  OAI21_X1 U7305 ( .B1(n6351), .B2(n6350), .A(n6349), .ZN(n6352) );
  OAI211_X1 U7306 ( .C1(n6355), .C2(n6354), .A(n6353), .B(n6352), .ZN(n6403)
         );
  AOI22_X1 U7307 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n6403), .B1(n6356), 
        .B2(n6401), .ZN(n6357) );
  OAI211_X1 U7308 ( .C1(n6359), .C2(n6406), .A(n6358), .B(n6357), .ZN(U3140)
         );
  AOI22_X1 U7309 ( .A1(n6361), .A2(n6399), .B1(n6398), .B2(n6360), .ZN(n6364)
         );
  AOI22_X1 U7310 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n6403), .B1(n6362), 
        .B2(n3078), .ZN(n6363) );
  OAI211_X1 U7311 ( .C1(n6365), .C2(n6389), .A(n6364), .B(n6363), .ZN(U3141)
         );
  AOI22_X1 U7312 ( .A1(n6367), .A2(n6399), .B1(n6398), .B2(n6366), .ZN(n6370)
         );
  AOI22_X1 U7313 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(n6403), .B1(n6368), 
        .B2(n3078), .ZN(n6369) );
  OAI211_X1 U7314 ( .C1(n6371), .C2(n6389), .A(n6370), .B(n6369), .ZN(U3142)
         );
  AOI22_X1 U7315 ( .A1(n6373), .A2(n6399), .B1(n6398), .B2(n6372), .ZN(n6376)
         );
  AOI22_X1 U7316 ( .A1(INSTQUEUE_REG_15__3__SCAN_IN), .A2(n6403), .B1(n6374), 
        .B2(n6401), .ZN(n6375) );
  OAI211_X1 U7317 ( .C1(n6377), .C2(n6406), .A(n6376), .B(n6375), .ZN(U3143)
         );
  AOI22_X1 U7318 ( .A1(n6379), .A2(n6399), .B1(n6398), .B2(n6378), .ZN(n6382)
         );
  AOI22_X1 U7319 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n6403), .B1(n6380), 
        .B2(n6401), .ZN(n6381) );
  OAI211_X1 U7320 ( .C1(n6383), .C2(n6406), .A(n6382), .B(n6381), .ZN(U3144)
         );
  AOI22_X1 U7321 ( .A1(n6385), .A2(n6399), .B1(n6398), .B2(n6384), .ZN(n6388)
         );
  AOI22_X1 U7322 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n6403), .B1(n6386), 
        .B2(n3078), .ZN(n6387) );
  OAI211_X1 U7323 ( .C1(n6390), .C2(n6389), .A(n6388), .B(n6387), .ZN(U3145)
         );
  AOI22_X1 U7324 ( .A1(n6392), .A2(n6399), .B1(n6398), .B2(n6391), .ZN(n6395)
         );
  AOI22_X1 U7325 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n6403), .B1(n6393), 
        .B2(n6401), .ZN(n6394) );
  OAI211_X1 U7326 ( .C1(n6396), .C2(n6406), .A(n6395), .B(n6394), .ZN(U3146)
         );
  AOI22_X1 U7327 ( .A1(n6400), .A2(n6399), .B1(n6398), .B2(n6397), .ZN(n6405)
         );
  AOI22_X1 U7328 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n6403), .B1(n6402), 
        .B2(n6401), .ZN(n6404) );
  OAI211_X1 U7329 ( .C1(n6407), .C2(n6406), .A(n6405), .B(n6404), .ZN(U3147)
         );
  INV_X1 U7330 ( .A(n6420), .ZN(n6423) );
  NOR2_X1 U7331 ( .A1(n6409), .A2(n6408), .ZN(n6416) );
  INV_X1 U7332 ( .A(n6416), .ZN(n6418) );
  OAI22_X1 U7333 ( .A1(n6412), .A2(n6411), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6410), .ZN(n6547) );
  NAND2_X1 U7334 ( .A1(n6413), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6555) );
  NAND2_X1 U7335 ( .A1(n6555), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6414) );
  AOI211_X1 U7336 ( .C1(n6416), .C2(n6415), .A(n6547), .B(n6414), .ZN(n6417)
         );
  AOI21_X1 U7337 ( .B1(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B2(n6418), .A(n6417), 
        .ZN(n6419) );
  OAI21_X1 U7338 ( .B1(n6421), .B2(n6420), .A(n6419), .ZN(n6422) );
  OAI21_X1 U7339 ( .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6423), .A(n6422), 
        .ZN(n6424) );
  AOI222_X1 U7340 ( .A1(n6426), .A2(n6425), .B1(n6426), .B2(n6424), .C1(n6425), 
        .C2(n6424), .ZN(n6434) );
  INV_X1 U7341 ( .A(n6427), .ZN(n6429) );
  NOR3_X1 U7342 ( .A1(n6430), .A2(n6429), .A3(n6428), .ZN(n6433) );
  OAI21_X1 U7343 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6431), 
        .ZN(n6432) );
  OAI211_X1 U7344 ( .C1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .C2(n6434), .A(n6433), .B(n6432), .ZN(n6442) );
  NOR2_X1 U7345 ( .A1(n6761), .A2(n6446), .ZN(n6441) );
  NAND3_X1 U7346 ( .A1(n6437), .A2(n6436), .A3(n6435), .ZN(n6439) );
  OAI21_X1 U7347 ( .B1(n6568), .B2(n6548), .A(n6596), .ZN(n6438) );
  NAND3_X1 U7348 ( .A1(n6439), .A2(STATE2_REG_2__SCAN_IN), .A3(n6438), .ZN(
        n6444) );
  AOI221_X1 U7349 ( .B1(STATE2_REG_0__SCAN_IN), .B2(n6442), .C1(
        STATE2_REG_0__SCAN_IN), .C2(STATE2_REG_1__SCAN_IN), .A(n6444), .ZN(
        n6440) );
  INV_X1 U7350 ( .A(n6440), .ZN(n6540) );
  OAI21_X1 U7351 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6568), .A(n6540), .ZN(
        n6450) );
  AOI211_X1 U7352 ( .C1(n6443), .C2(n6442), .A(n6441), .B(n6450), .ZN(n6449)
         );
  OAI211_X1 U7353 ( .C1(n6446), .C2(n6445), .A(n6596), .B(n6444), .ZN(n6447)
         );
  OAI221_X1 U7354 ( .B1(n6596), .B2(n6449), .C1(n6596), .C2(n6448), .A(n6447), 
        .ZN(U3148) );
  NAND3_X1 U7355 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6457), .A3(n6450), .ZN(
        n6456) );
  OAI21_X1 U7356 ( .B1(READY_N), .B2(n6452), .A(n6451), .ZN(n6454) );
  AOI21_X1 U7357 ( .B1(n6454), .B2(n6540), .A(n6453), .ZN(n6455) );
  NAND2_X1 U7358 ( .A1(n6456), .A2(n6455), .ZN(U3149) );
  OAI211_X1 U7359 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6568), .A(n6457), .B(
        n6538), .ZN(n6459) );
  OAI21_X1 U7360 ( .B1(n6572), .B2(n6459), .A(n6458), .ZN(U3150) );
  INV_X1 U7361 ( .A(n6537), .ZN(n6460) );
  AND2_X1 U7362 ( .A1(DATAWIDTH_REG_31__SCAN_IN), .A2(n6460), .ZN(U3151) );
  INV_X1 U7363 ( .A(DATAWIDTH_REG_30__SCAN_IN), .ZN(n6632) );
  NOR2_X1 U7364 ( .A1(n6537), .A2(n6632), .ZN(U3152) );
  AND2_X1 U7365 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6460), .ZN(U3153) );
  AND2_X1 U7366 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6460), .ZN(U3154) );
  AND2_X1 U7367 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6460), .ZN(U3155) );
  AND2_X1 U7368 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6460), .ZN(U3156) );
  AND2_X1 U7369 ( .A1(DATAWIDTH_REG_25__SCAN_IN), .A2(n6460), .ZN(U3157) );
  AND2_X1 U7370 ( .A1(DATAWIDTH_REG_24__SCAN_IN), .A2(n6460), .ZN(U3158) );
  AND2_X1 U7371 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6460), .ZN(U3159) );
  AND2_X1 U7372 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6460), .ZN(U3160) );
  AND2_X1 U7373 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6460), .ZN(U3161) );
  AND2_X1 U7374 ( .A1(n6460), .A2(DATAWIDTH_REG_20__SCAN_IN), .ZN(U3162) );
  AND2_X1 U7375 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(n6460), .ZN(U3163) );
  AND2_X1 U7376 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6460), .ZN(U3164) );
  AND2_X1 U7377 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6460), .ZN(U3165) );
  INV_X1 U7378 ( .A(DATAWIDTH_REG_16__SCAN_IN), .ZN(n6766) );
  NOR2_X1 U7379 ( .A1(n6537), .A2(n6766), .ZN(U3166) );
  AND2_X1 U7380 ( .A1(DATAWIDTH_REG_15__SCAN_IN), .A2(n6460), .ZN(U3167) );
  AND2_X1 U7381 ( .A1(DATAWIDTH_REG_14__SCAN_IN), .A2(n6460), .ZN(U3168) );
  AND2_X1 U7382 ( .A1(DATAWIDTH_REG_13__SCAN_IN), .A2(n6460), .ZN(U3169) );
  AND2_X1 U7383 ( .A1(DATAWIDTH_REG_12__SCAN_IN), .A2(n6460), .ZN(U3170) );
  AND2_X1 U7384 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6460), .ZN(U3171) );
  AND2_X1 U7385 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(n6460), .ZN(U3172) );
  AND2_X1 U7386 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6460), .ZN(U3173) );
  INV_X1 U7387 ( .A(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6630) );
  NOR2_X1 U7388 ( .A1(n6537), .A2(n6630), .ZN(U3174) );
  AND2_X1 U7389 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6460), .ZN(U3175) );
  INV_X1 U7390 ( .A(DATAWIDTH_REG_6__SCAN_IN), .ZN(n6714) );
  NOR2_X1 U7391 ( .A1(n6537), .A2(n6714), .ZN(U3176) );
  AND2_X1 U7392 ( .A1(DATAWIDTH_REG_5__SCAN_IN), .A2(n6460), .ZN(U3177) );
  AND2_X1 U7393 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6460), .ZN(U3178) );
  AND2_X1 U7394 ( .A1(DATAWIDTH_REG_3__SCAN_IN), .A2(n6460), .ZN(U3179) );
  AND2_X1 U7395 ( .A1(DATAWIDTH_REG_2__SCAN_IN), .A2(n6460), .ZN(U3180) );
  NAND2_X1 U7396 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6467) );
  NAND2_X1 U7397 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6466) );
  NAND2_X1 U7398 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .ZN(n6473) );
  NAND2_X1 U7399 ( .A1(n6466), .A2(n6473), .ZN(n6463) );
  OAI211_X1 U7400 ( .C1(n6461), .C2(NA_N), .A(n6474), .B(n6464), .ZN(n6462) );
  INV_X1 U7401 ( .A(n6462), .ZN(n6479) );
  AOI21_X1 U7402 ( .B1(n6464), .B2(n6463), .A(n6479), .ZN(n6465) );
  OAI221_X1 U7403 ( .B1(n6577), .B2(REQUESTPENDING_REG_SCAN_IN), .C1(n6577), 
        .C2(n6467), .A(n6465), .ZN(U3181) );
  INV_X1 U7404 ( .A(n6466), .ZN(n6471) );
  INV_X1 U7405 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6475) );
  OAI21_X1 U7406 ( .B1(n6475), .B2(n6474), .A(n6467), .ZN(n6468) );
  INV_X1 U7407 ( .A(n6468), .ZN(n6470) );
  OAI211_X1 U7408 ( .C1(n6471), .C2(n6470), .A(n6469), .B(n6473), .ZN(U3182)
         );
  AOI221_X1 U7409 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6568), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6472) );
  AOI221_X1 U7410 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6472), .C2(HOLD), .A(n6474), .ZN(n6478) );
  OR4_X1 U7411 ( .A1(n6475), .A2(n6474), .A3(n6473), .A4(NA_N), .ZN(n6477) );
  NAND3_X1 U7412 ( .A1(READY_N), .A2(STATE_REG_2__SCAN_IN), .A3(
        STATE_REG_1__SCAN_IN), .ZN(n6476) );
  OAI211_X1 U7413 ( .C1(n6479), .C2(n6478), .A(n6477), .B(n6476), .ZN(U3183)
         );
  NAND2_X1 U7414 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6577), .ZN(n6532) );
  NOR2_X2 U7415 ( .A1(STATE_REG_2__SCAN_IN), .A2(n6565), .ZN(n6530) );
  AOI22_X1 U7416 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6530), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6565), .ZN(n6480) );
  OAI21_X1 U7417 ( .B1(n5099), .B2(n6532), .A(n6480), .ZN(U3184) );
  AOI22_X1 U7418 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6530), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6565), .ZN(n6481) );
  OAI21_X1 U7419 ( .B1(n6482), .B2(n6532), .A(n6481), .ZN(U3185) );
  AOI22_X1 U7420 ( .A1(REIP_REG_4__SCAN_IN), .A2(n6530), .B1(
        ADDRESS_REG_2__SCAN_IN), .B2(n6565), .ZN(n6483) );
  OAI21_X1 U7421 ( .B1(n6484), .B2(n6532), .A(n6483), .ZN(U3186) );
  AOI22_X1 U7422 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6530), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6565), .ZN(n6485) );
  OAI21_X1 U7423 ( .B1(n6486), .B2(n6532), .A(n6485), .ZN(U3187) );
  AOI22_X1 U7424 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6530), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6565), .ZN(n6487) );
  OAI21_X1 U7425 ( .B1(n6488), .B2(n6532), .A(n6487), .ZN(U3188) );
  AOI22_X1 U7426 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6530), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6565), .ZN(n6489) );
  OAI21_X1 U7427 ( .B1(n6490), .B2(n6532), .A(n6489), .ZN(U3189) );
  AOI22_X1 U7428 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6530), .B1(
        ADDRESS_REG_6__SCAN_IN), .B2(n6565), .ZN(n6491) );
  OAI21_X1 U7429 ( .B1(n6492), .B2(n6532), .A(n6491), .ZN(U3190) );
  INV_X1 U7430 ( .A(n6530), .ZN(n6529) );
  INV_X1 U7431 ( .A(n6532), .ZN(n6527) );
  AOI22_X1 U7432 ( .A1(REIP_REG_8__SCAN_IN), .A2(n6527), .B1(
        ADDRESS_REG_7__SCAN_IN), .B2(n6565), .ZN(n6493) );
  OAI21_X1 U7433 ( .B1(n6495), .B2(n6529), .A(n6493), .ZN(U3191) );
  AOI22_X1 U7434 ( .A1(REIP_REG_10__SCAN_IN), .A2(n6530), .B1(
        ADDRESS_REG_8__SCAN_IN), .B2(n6565), .ZN(n6494) );
  OAI21_X1 U7435 ( .B1(n6495), .B2(n6532), .A(n6494), .ZN(U3192) );
  AOI22_X1 U7436 ( .A1(REIP_REG_11__SCAN_IN), .A2(n6530), .B1(
        ADDRESS_REG_9__SCAN_IN), .B2(n6565), .ZN(n6496) );
  OAI21_X1 U7437 ( .B1(n6497), .B2(n6532), .A(n6496), .ZN(U3193) );
  AOI22_X1 U7438 ( .A1(REIP_REG_12__SCAN_IN), .A2(n6530), .B1(
        ADDRESS_REG_10__SCAN_IN), .B2(n6565), .ZN(n6498) );
  OAI21_X1 U7439 ( .B1(n6499), .B2(n6532), .A(n6498), .ZN(U3194) );
  INV_X1 U7440 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6502) );
  INV_X1 U7441 ( .A(ADDRESS_REG_11__SCAN_IN), .ZN(n6748) );
  OAI222_X1 U7442 ( .A1(n6529), .A2(n6502), .B1(n6748), .B2(n6577), .C1(n6500), 
        .C2(n6532), .ZN(U3195) );
  AOI22_X1 U7443 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6530), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6565), .ZN(n6501) );
  OAI21_X1 U7444 ( .B1(n6502), .B2(n6532), .A(n6501), .ZN(U3196) );
  AOI22_X1 U7445 ( .A1(REIP_REG_15__SCAN_IN), .A2(n6530), .B1(
        ADDRESS_REG_13__SCAN_IN), .B2(n6565), .ZN(n6503) );
  OAI21_X1 U7446 ( .B1(n6717), .B2(n6532), .A(n6503), .ZN(U3197) );
  INV_X1 U7447 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6505) );
  AOI22_X1 U7448 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6530), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6565), .ZN(n6504) );
  OAI21_X1 U7449 ( .B1(n6505), .B2(n6532), .A(n6504), .ZN(U3198) );
  AOI22_X1 U7450 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6527), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6565), .ZN(n6506) );
  OAI21_X1 U7451 ( .B1(n6605), .B2(n6529), .A(n6506), .ZN(U3199) );
  AOI22_X1 U7452 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6527), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6565), .ZN(n6507) );
  OAI21_X1 U7453 ( .B1(n6508), .B2(n6529), .A(n6507), .ZN(U3200) );
  INV_X1 U7454 ( .A(ADDRESS_REG_17__SCAN_IN), .ZN(n6620) );
  OAI222_X1 U7455 ( .A1(n6529), .A2(n6509), .B1(n6620), .B2(n6577), .C1(n6508), 
        .C2(n6532), .ZN(U3201) );
  AOI22_X1 U7456 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6527), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6565), .ZN(n6510) );
  OAI21_X1 U7457 ( .B1(n6512), .B2(n6529), .A(n6510), .ZN(U3202) );
  INV_X1 U7458 ( .A(ADDRESS_REG_19__SCAN_IN), .ZN(n6511) );
  OAI222_X1 U7459 ( .A1(n6532), .A2(n6512), .B1(n6511), .B2(n6577), .C1(n6514), 
        .C2(n6529), .ZN(U3203) );
  AOI22_X1 U7460 ( .A1(REIP_REG_22__SCAN_IN), .A2(n6530), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6565), .ZN(n6513) );
  OAI21_X1 U7461 ( .B1(n6514), .B2(n6532), .A(n6513), .ZN(U3204) );
  AOI22_X1 U7462 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6530), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6565), .ZN(n6515) );
  OAI21_X1 U7463 ( .B1(n6516), .B2(n6532), .A(n6515), .ZN(U3205) );
  AOI22_X1 U7464 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6527), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6565), .ZN(n6517) );
  OAI21_X1 U7465 ( .B1(n3740), .B2(n6529), .A(n6517), .ZN(U3206) );
  AOI22_X1 U7466 ( .A1(REIP_REG_24__SCAN_IN), .A2(n6527), .B1(
        ADDRESS_REG_23__SCAN_IN), .B2(n6565), .ZN(n6518) );
  OAI21_X1 U7467 ( .B1(n6521), .B2(n6529), .A(n6518), .ZN(U3207) );
  INV_X1 U7468 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n6520) );
  OAI222_X1 U7469 ( .A1(n6532), .A2(n6521), .B1(n6520), .B2(n6577), .C1(n6519), 
        .C2(n6529), .ZN(U3208) );
  AOI22_X1 U7470 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6527), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6565), .ZN(n6522) );
  OAI21_X1 U7471 ( .B1(n6523), .B2(n6529), .A(n6522), .ZN(U3209) );
  AOI22_X1 U7472 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6527), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6565), .ZN(n6524) );
  OAI21_X1 U7473 ( .B1(n6724), .B2(n6529), .A(n6524), .ZN(U3210) );
  AOI22_X1 U7474 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6527), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6565), .ZN(n6525) );
  OAI21_X1 U7475 ( .B1(n6526), .B2(n6529), .A(n6525), .ZN(U3211) );
  AOI22_X1 U7476 ( .A1(REIP_REG_29__SCAN_IN), .A2(n6527), .B1(
        ADDRESS_REG_28__SCAN_IN), .B2(n6565), .ZN(n6528) );
  OAI21_X1 U7477 ( .B1(n6533), .B2(n6529), .A(n6528), .ZN(U3212) );
  AOI22_X1 U7478 ( .A1(REIP_REG_31__SCAN_IN), .A2(n6530), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6565), .ZN(n6531) );
  OAI21_X1 U7479 ( .B1(n6533), .B2(n6532), .A(n6531), .ZN(U3213) );
  MUX2_X1 U7480 ( .A(BE_N_REG_3__SCAN_IN), .B(BYTEENABLE_REG_3__SCAN_IN), .S(
        n6577), .Z(U3445) );
  MUX2_X1 U7481 ( .A(BE_N_REG_2__SCAN_IN), .B(BYTEENABLE_REG_2__SCAN_IN), .S(
        n6577), .Z(U3446) );
  MUX2_X1 U7482 ( .A(BE_N_REG_1__SCAN_IN), .B(BYTEENABLE_REG_1__SCAN_IN), .S(
        n6577), .Z(U3447) );
  MUX2_X1 U7483 ( .A(BE_N_REG_0__SCAN_IN), .B(BYTEENABLE_REG_0__SCAN_IN), .S(
        n6577), .Z(U3448) );
  OAI21_X1 U7484 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6537), .A(n6535), .ZN(
        n6534) );
  INV_X1 U7485 ( .A(n6534), .ZN(U3451) );
  INV_X1 U7486 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6536) );
  OAI21_X1 U7487 ( .B1(n6537), .B2(n6536), .A(n6535), .ZN(U3452) );
  OAI211_X1 U7488 ( .C1(n6761), .C2(n6540), .A(n6539), .B(n6538), .ZN(U3453)
         );
  AOI22_X1 U7489 ( .A1(n6544), .A2(n6543), .B1(n6542), .B2(n6541), .ZN(n6545)
         );
  INV_X1 U7490 ( .A(n6545), .ZN(n6546) );
  MUX2_X1 U7491 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6546), .S(n6552), 
        .Z(U3456) );
  INV_X1 U7492 ( .A(n6547), .ZN(n6549) );
  OAI22_X1 U7493 ( .A1(n6549), .A2(n6554), .B1(INSTADDRPOINTER_REG_0__SCAN_IN), 
        .B2(n6548), .ZN(n6551) );
  OAI22_X1 U7494 ( .A1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A2(n6552), .B1(n6551), .B2(n6550), .ZN(n6553) );
  OAI21_X1 U7495 ( .B1(n6555), .B2(n6554), .A(n6553), .ZN(U3461) );
  INV_X1 U7496 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6557) );
  NOR3_X1 U7497 ( .A1(n6557), .A2(REIP_REG_0__SCAN_IN), .A3(
        REIP_REG_1__SCAN_IN), .ZN(n6556) );
  AOI221_X1 U7498 ( .B1(n6558), .B2(n6557), .C1(REIP_REG_1__SCAN_IN), .C2(
        REIP_REG_0__SCAN_IN), .A(n6556), .ZN(n6560) );
  INV_X1 U7499 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6559) );
  INV_X1 U7500 ( .A(n6564), .ZN(n6561) );
  AOI22_X1 U7501 ( .A1(n6564), .A2(n6560), .B1(n6559), .B2(n6561), .ZN(U3468)
         );
  NOR2_X1 U7502 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .ZN(
        n6563) );
  INV_X1 U7503 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6562) );
  AOI22_X1 U7504 ( .A1(n6564), .A2(n6563), .B1(n6562), .B2(n6561), .ZN(U3469)
         );
  INV_X1 U7505 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6734) );
  AOI22_X1 U7506 ( .A1(n6577), .A2(READREQUEST_REG_SCAN_IN), .B1(n6734), .B2(
        n6565), .ZN(U3470) );
  AOI211_X1 U7507 ( .C1(n6569), .C2(n6568), .A(n6567), .B(n6566), .ZN(n6576)
         );
  OAI211_X1 U7508 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6571), .A(n6570), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6573) );
  AOI21_X1 U7509 ( .B1(n6573), .B2(STATE2_REG_0__SCAN_IN), .A(n6572), .ZN(
        n6575) );
  NAND2_X1 U7510 ( .A1(n6576), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6574) );
  OAI21_X1 U7511 ( .B1(n6576), .B2(n6575), .A(n6574), .ZN(U3472) );
  MUX2_X1 U7512 ( .A(M_IO_N_REG_SCAN_IN), .B(MEMORYFETCH_REG_SCAN_IN), .S(
        n6577), .Z(U3473) );
  INV_X1 U7513 ( .A(n6578), .ZN(n6587) );
  NOR3_X1 U7514 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n6580), .A3(n6579), 
        .ZN(n6581) );
  AOI21_X1 U7515 ( .B1(n6582), .B2(REIP_REG_18__SCAN_IN), .A(n6581), .ZN(n6583) );
  OAI21_X1 U7516 ( .B1(n6585), .B2(n6584), .A(n6583), .ZN(n6586) );
  AOI21_X1 U7517 ( .B1(n6587), .B2(INSTADDRPOINTER_REG_18__SCAN_IN), .A(n6586), 
        .ZN(n6588) );
  OAI21_X1 U7518 ( .B1(n6590), .B2(n6589), .A(n6588), .ZN(n6784) );
  INV_X1 U7519 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n6592) );
  INV_X1 U7520 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6735) );
  AOI22_X1 U7521 ( .A1(n6592), .A2(keyinput85), .B1(keyinput122), .B2(n6735), 
        .ZN(n6591) );
  OAI221_X1 U7522 ( .B1(n6592), .B2(keyinput85), .C1(n6735), .C2(keyinput122), 
        .A(n6591), .ZN(n6601) );
  INV_X1 U7523 ( .A(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n6760) );
  AOI22_X1 U7524 ( .A1(n6760), .A2(keyinput71), .B1(n6763), .B2(keyinput104), 
        .ZN(n6593) );
  OAI221_X1 U7525 ( .B1(n6760), .B2(keyinput71), .C1(n6763), .C2(keyinput104), 
        .A(n6593), .ZN(n6600) );
  AOI22_X1 U7526 ( .A1(n6717), .A2(keyinput66), .B1(n3657), .B2(keyinput97), 
        .ZN(n6594) );
  OAI221_X1 U7527 ( .B1(n6717), .B2(keyinput66), .C1(n3657), .C2(keyinput97), 
        .A(n6594), .ZN(n6599) );
  AOI22_X1 U7528 ( .A1(n6597), .A2(keyinput89), .B1(n6596), .B2(keyinput90), 
        .ZN(n6595) );
  OAI221_X1 U7529 ( .B1(n6597), .B2(keyinput89), .C1(n6596), .C2(keyinput90), 
        .A(n6595), .ZN(n6598) );
  NOR4_X1 U7530 ( .A1(n6601), .A2(n6600), .A3(n6599), .A4(n6598), .ZN(n6640)
         );
  INV_X1 U7531 ( .A(LWORD_REG_2__SCAN_IN), .ZN(n6747) );
  AOI22_X1 U7532 ( .A1(n6747), .A2(keyinput77), .B1(keyinput73), .B2(n6714), 
        .ZN(n6602) );
  OAI221_X1 U7533 ( .B1(n6747), .B2(keyinput77), .C1(n6714), .C2(keyinput73), 
        .A(n6602), .ZN(n6613) );
  AOI22_X1 U7534 ( .A1(REIP_REG_13__SCAN_IN), .A2(keyinput82), .B1(n6761), 
        .B2(keyinput67), .ZN(n6603) );
  OAI221_X1 U7535 ( .B1(REIP_REG_13__SCAN_IN), .B2(keyinput82), .C1(n6761), 
        .C2(keyinput67), .A(n6603), .ZN(n6612) );
  INV_X1 U7536 ( .A(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n6606) );
  AOI22_X1 U7537 ( .A1(n6606), .A2(keyinput95), .B1(keyinput125), .B2(n6605), 
        .ZN(n6604) );
  OAI221_X1 U7538 ( .B1(n6606), .B2(keyinput95), .C1(n6605), .C2(keyinput125), 
        .A(n6604), .ZN(n6611) );
  AOI22_X1 U7539 ( .A1(n6609), .A2(keyinput96), .B1(n6608), .B2(keyinput103), 
        .ZN(n6607) );
  OAI221_X1 U7540 ( .B1(n6609), .B2(keyinput96), .C1(n6608), .C2(keyinput103), 
        .A(n6607), .ZN(n6610) );
  NOR4_X1 U7541 ( .A1(n6613), .A2(n6612), .A3(n6611), .A4(n6610), .ZN(n6639)
         );
  INV_X1 U7542 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n6615) );
  AOI22_X1 U7543 ( .A1(n6724), .A2(keyinput113), .B1(n6615), .B2(keyinput111), 
        .ZN(n6614) );
  OAI221_X1 U7544 ( .B1(n6724), .B2(keyinput113), .C1(n6615), .C2(keyinput111), 
        .A(n6614), .ZN(n6625) );
  AOI22_X1 U7545 ( .A1(n6737), .A2(keyinput126), .B1(keyinput99), .B2(n6767), 
        .ZN(n6616) );
  OAI221_X1 U7546 ( .B1(n6737), .B2(keyinput126), .C1(n6767), .C2(keyinput99), 
        .A(n6616), .ZN(n6624) );
  INV_X1 U7547 ( .A(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n6731) );
  AOI22_X1 U7548 ( .A1(n6618), .A2(keyinput75), .B1(n6731), .B2(keyinput118), 
        .ZN(n6617) );
  OAI221_X1 U7549 ( .B1(n6618), .B2(keyinput75), .C1(n6731), .C2(keyinput118), 
        .A(n6617), .ZN(n6623) );
  AOI22_X1 U7550 ( .A1(n6621), .A2(keyinput68), .B1(keyinput102), .B2(n6620), 
        .ZN(n6619) );
  OAI221_X1 U7551 ( .B1(n6621), .B2(keyinput68), .C1(n6620), .C2(keyinput102), 
        .A(n6619), .ZN(n6622) );
  NOR4_X1 U7552 ( .A1(n6625), .A2(n6624), .A3(n6623), .A4(n6622), .ZN(n6638)
         );
  INV_X1 U7553 ( .A(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n6754) );
  INV_X1 U7554 ( .A(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n6627) );
  AOI22_X1 U7555 ( .A1(n6754), .A2(keyinput78), .B1(keyinput84), .B2(n6627), 
        .ZN(n6626) );
  OAI221_X1 U7556 ( .B1(n6754), .B2(keyinput78), .C1(n6627), .C2(keyinput84), 
        .A(n6626), .ZN(n6636) );
  INV_X1 U7557 ( .A(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n6750) );
  AOI22_X1 U7558 ( .A1(n6750), .A2(keyinput87), .B1(keyinput98), .B2(n6744), 
        .ZN(n6628) );
  OAI221_X1 U7559 ( .B1(n6750), .B2(keyinput87), .C1(n6744), .C2(keyinput98), 
        .A(n6628), .ZN(n6635) );
  AOI22_X1 U7560 ( .A1(n6630), .A2(keyinput124), .B1(keyinput93), .B2(n4356), 
        .ZN(n6629) );
  OAI221_X1 U7561 ( .B1(n6630), .B2(keyinput124), .C1(n4356), .C2(keyinput93), 
        .A(n6629), .ZN(n6634) );
  AOI22_X1 U7562 ( .A1(n6632), .A2(keyinput69), .B1(n6723), .B2(keyinput65), 
        .ZN(n6631) );
  OAI221_X1 U7563 ( .B1(n6632), .B2(keyinput69), .C1(n6723), .C2(keyinput65), 
        .A(n6631), .ZN(n6633) );
  NOR4_X1 U7564 ( .A1(n6636), .A2(n6635), .A3(n6634), .A4(n6633), .ZN(n6637)
         );
  NAND4_X1 U7565 ( .A1(n6640), .A2(n6639), .A3(n6638), .A4(n6637), .ZN(n6782)
         );
  AOI22_X1 U7566 ( .A1(UWORD_REG_5__SCAN_IN), .A2(keyinput92), .B1(
        INSTADDRPOINTER_REG_19__SCAN_IN), .B2(keyinput127), .ZN(n6641) );
  OAI221_X1 U7567 ( .B1(UWORD_REG_5__SCAN_IN), .B2(keyinput92), .C1(
        INSTADDRPOINTER_REG_19__SCAN_IN), .C2(keyinput127), .A(n6641), .ZN(
        n6648) );
  AOI22_X1 U7568 ( .A1(UWORD_REG_8__SCAN_IN), .A2(keyinput80), .B1(
        EAX_REG_29__SCAN_IN), .B2(keyinput101), .ZN(n6642) );
  OAI221_X1 U7569 ( .B1(UWORD_REG_8__SCAN_IN), .B2(keyinput80), .C1(
        EAX_REG_29__SCAN_IN), .C2(keyinput101), .A(n6642), .ZN(n6647) );
  AOI22_X1 U7570 ( .A1(ADDRESS_REG_11__SCAN_IN), .A2(keyinput76), .B1(
        EBX_REG_25__SCAN_IN), .B2(keyinput74), .ZN(n6643) );
  OAI221_X1 U7571 ( .B1(ADDRESS_REG_11__SCAN_IN), .B2(keyinput76), .C1(
        EBX_REG_25__SCAN_IN), .C2(keyinput74), .A(n6643), .ZN(n6646) );
  AOI22_X1 U7572 ( .A1(DATAI_0_), .A2(keyinput86), .B1(FLUSH_REG_SCAN_IN), 
        .B2(keyinput70), .ZN(n6644) );
  OAI221_X1 U7573 ( .B1(DATAI_0_), .B2(keyinput86), .C1(FLUSH_REG_SCAN_IN), 
        .C2(keyinput70), .A(n6644), .ZN(n6645) );
  NOR4_X1 U7574 ( .A1(n6648), .A2(n6647), .A3(n6646), .A4(n6645), .ZN(n6676)
         );
  AOI22_X1 U7575 ( .A1(W_R_N_REG_SCAN_IN), .A2(keyinput88), .B1(
        INSTQUEUE_REG_13__2__SCAN_IN), .B2(keyinput123), .ZN(n6649) );
  OAI221_X1 U7576 ( .B1(W_R_N_REG_SCAN_IN), .B2(keyinput88), .C1(
        INSTQUEUE_REG_13__2__SCAN_IN), .C2(keyinput123), .A(n6649), .ZN(n6656)
         );
  AOI22_X1 U7577 ( .A1(EAX_REG_6__SCAN_IN), .A2(keyinput105), .B1(
        INSTQUEUE_REG_3__3__SCAN_IN), .B2(keyinput81), .ZN(n6650) );
  OAI221_X1 U7578 ( .B1(EAX_REG_6__SCAN_IN), .B2(keyinput105), .C1(
        INSTQUEUE_REG_3__3__SCAN_IN), .C2(keyinput81), .A(n6650), .ZN(n6655)
         );
  AOI22_X1 U7579 ( .A1(ADDRESS_REG_24__SCAN_IN), .A2(keyinput83), .B1(
        DATAO_REG_0__SCAN_IN), .B2(keyinput112), .ZN(n6651) );
  OAI221_X1 U7580 ( .B1(ADDRESS_REG_24__SCAN_IN), .B2(keyinput83), .C1(
        DATAO_REG_0__SCAN_IN), .C2(keyinput112), .A(n6651), .ZN(n6654) );
  AOI22_X1 U7581 ( .A1(DATAI_9_), .A2(keyinput72), .B1(
        DATAWIDTH_REG_16__SCAN_IN), .B2(keyinput79), .ZN(n6652) );
  OAI221_X1 U7582 ( .B1(DATAI_9_), .B2(keyinput72), .C1(
        DATAWIDTH_REG_16__SCAN_IN), .C2(keyinput79), .A(n6652), .ZN(n6653) );
  NOR4_X1 U7583 ( .A1(n6656), .A2(n6655), .A3(n6654), .A4(n6653), .ZN(n6675)
         );
  AOI22_X1 U7584 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(keyinput120), .B1(
        UWORD_REG_7__SCAN_IN), .B2(keyinput107), .ZN(n6657) );
  OAI221_X1 U7585 ( .B1(DATAWIDTH_REG_20__SCAN_IN), .B2(keyinput120), .C1(
        UWORD_REG_7__SCAN_IN), .C2(keyinput107), .A(n6657), .ZN(n6664) );
  AOI22_X1 U7586 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(keyinput119), .B1(
        INSTQUEUE_REG_0__4__SCAN_IN), .B2(keyinput100), .ZN(n6658) );
  OAI221_X1 U7587 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(keyinput119), .C1(
        INSTQUEUE_REG_0__4__SCAN_IN), .C2(keyinput100), .A(n6658), .ZN(n6663)
         );
  AOI22_X1 U7588 ( .A1(DATAO_REG_23__SCAN_IN), .A2(keyinput91), .B1(DATAI_13_), 
        .B2(keyinput121), .ZN(n6659) );
  OAI221_X1 U7589 ( .B1(DATAO_REG_23__SCAN_IN), .B2(keyinput91), .C1(DATAI_13_), .C2(keyinput121), .A(n6659), .ZN(n6662) );
  AOI22_X1 U7590 ( .A1(EAX_REG_30__SCAN_IN), .A2(keyinput64), .B1(
        INSTADDRPOINTER_REG_11__SCAN_IN), .B2(keyinput110), .ZN(n6660) );
  OAI221_X1 U7591 ( .B1(EAX_REG_30__SCAN_IN), .B2(keyinput64), .C1(
        INSTADDRPOINTER_REG_11__SCAN_IN), .C2(keyinput110), .A(n6660), .ZN(
        n6661) );
  NOR4_X1 U7592 ( .A1(n6664), .A2(n6663), .A3(n6662), .A4(n6661), .ZN(n6674)
         );
  AOI22_X1 U7593 ( .A1(LWORD_REG_5__SCAN_IN), .A2(keyinput109), .B1(
        INSTQUEUE_REG_5__0__SCAN_IN), .B2(keyinput106), .ZN(n6665) );
  OAI221_X1 U7594 ( .B1(LWORD_REG_5__SCAN_IN), .B2(keyinput109), .C1(
        INSTQUEUE_REG_5__0__SCAN_IN), .C2(keyinput106), .A(n6665), .ZN(n6672)
         );
  AOI22_X1 U7595 ( .A1(DATAO_REG_21__SCAN_IN), .A2(keyinput116), .B1(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .B2(keyinput117), .ZN(n6666) );
  OAI221_X1 U7596 ( .B1(DATAO_REG_21__SCAN_IN), .B2(keyinput116), .C1(
        INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .C2(keyinput117), .A(n6666), .ZN(
        n6671) );
  AOI22_X1 U7597 ( .A1(EAX_REG_12__SCAN_IN), .A2(keyinput115), .B1(
        INSTQUEUE_REG_5__1__SCAN_IN), .B2(keyinput94), .ZN(n6667) );
  OAI221_X1 U7598 ( .B1(EAX_REG_12__SCAN_IN), .B2(keyinput115), .C1(
        INSTQUEUE_REG_5__1__SCAN_IN), .C2(keyinput94), .A(n6667), .ZN(n6670)
         );
  AOI22_X1 U7599 ( .A1(ADDRESS_REG_19__SCAN_IN), .A2(keyinput108), .B1(
        INSTADDRPOINTER_REG_17__SCAN_IN), .B2(keyinput114), .ZN(n6668) );
  OAI221_X1 U7600 ( .B1(ADDRESS_REG_19__SCAN_IN), .B2(keyinput108), .C1(
        INSTADDRPOINTER_REG_17__SCAN_IN), .C2(keyinput114), .A(n6668), .ZN(
        n6669) );
  NOR4_X1 U7601 ( .A1(n6672), .A2(n6671), .A3(n6670), .A4(n6669), .ZN(n6673)
         );
  NAND4_X1 U7602 ( .A1(n6676), .A2(n6675), .A3(n6674), .A4(n6673), .ZN(n6781)
         );
  OAI22_X1 U7603 ( .A1(INSTQUEUE_REG_13__0__SCAN_IN), .A2(keyinput21), .B1(
        INSTADDRPOINTER_REG_19__SCAN_IN), .B2(keyinput63), .ZN(n6677) );
  AOI221_X1 U7604 ( .B1(INSTQUEUE_REG_13__0__SCAN_IN), .B2(keyinput21), .C1(
        keyinput63), .C2(INSTADDRPOINTER_REG_19__SCAN_IN), .A(n6677), .ZN(
        n6684) );
  OAI22_X1 U7605 ( .A1(INSTADDRPOINTER_REG_2__SCAN_IN), .A2(keyinput33), .B1(
        keyinput18), .B2(REIP_REG_13__SCAN_IN), .ZN(n6678) );
  AOI221_X1 U7606 ( .B1(INSTADDRPOINTER_REG_2__SCAN_IN), .B2(keyinput33), .C1(
        REIP_REG_13__SCAN_IN), .C2(keyinput18), .A(n6678), .ZN(n6683) );
  OAI22_X1 U7607 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(keyinput50), .B1(
        DATAI_15_), .B2(keyinput29), .ZN(n6679) );
  AOI221_X1 U7608 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(keyinput50), 
        .C1(keyinput29), .C2(DATAI_15_), .A(n6679), .ZN(n6682) );
  OAI22_X1 U7609 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(keyinput39), .B1(
        keyinput61), .B2(REIP_REG_17__SCAN_IN), .ZN(n6680) );
  AOI221_X1 U7610 ( .B1(INSTQUEUE_REG_0__7__SCAN_IN), .B2(keyinput39), .C1(
        REIP_REG_17__SCAN_IN), .C2(keyinput61), .A(n6680), .ZN(n6681) );
  NAND4_X1 U7611 ( .A1(n6684), .A2(n6683), .A3(n6682), .A4(n6681), .ZN(n6712)
         );
  OAI22_X1 U7612 ( .A1(DATAO_REG_23__SCAN_IN), .A2(keyinput27), .B1(
        DATAWIDTH_REG_30__SCAN_IN), .B2(keyinput5), .ZN(n6685) );
  AOI221_X1 U7613 ( .B1(DATAO_REG_23__SCAN_IN), .B2(keyinput27), .C1(keyinput5), .C2(DATAWIDTH_REG_30__SCAN_IN), .A(n6685), .ZN(n6692) );
  OAI22_X1 U7614 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(keyinput17), .B1(
        PHYADDRPOINTER_REG_30__SCAN_IN), .B2(keyinput25), .ZN(n6686) );
  AOI221_X1 U7615 ( .B1(INSTQUEUE_REG_3__3__SCAN_IN), .B2(keyinput17), .C1(
        keyinput25), .C2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n6686), .ZN(n6691) );
  OAI22_X1 U7616 ( .A1(EBX_REG_16__SCAN_IN), .A2(keyinput11), .B1(DATAI_0_), 
        .B2(keyinput22), .ZN(n6687) );
  AOI221_X1 U7617 ( .B1(EBX_REG_16__SCAN_IN), .B2(keyinput11), .C1(keyinput22), 
        .C2(DATAI_0_), .A(n6687), .ZN(n6690) );
  OAI22_X1 U7618 ( .A1(EBX_REG_10__SCAN_IN), .A2(keyinput4), .B1(keyinput43), 
        .B2(UWORD_REG_7__SCAN_IN), .ZN(n6688) );
  AOI221_X1 U7619 ( .B1(EBX_REG_10__SCAN_IN), .B2(keyinput4), .C1(
        UWORD_REG_7__SCAN_IN), .C2(keyinput43), .A(n6688), .ZN(n6689) );
  NAND4_X1 U7620 ( .A1(n6692), .A2(n6691), .A3(n6690), .A4(n6689), .ZN(n6711)
         );
  OAI22_X1 U7621 ( .A1(EAX_REG_30__SCAN_IN), .A2(keyinput0), .B1(keyinput60), 
        .B2(DATAWIDTH_REG_8__SCAN_IN), .ZN(n6693) );
  AOI221_X1 U7622 ( .B1(EAX_REG_30__SCAN_IN), .B2(keyinput0), .C1(
        DATAWIDTH_REG_8__SCAN_IN), .C2(keyinput60), .A(n6693), .ZN(n6700) );
  OAI22_X1 U7623 ( .A1(ADDRESS_REG_24__SCAN_IN), .A2(keyinput19), .B1(
        FLUSH_REG_SCAN_IN), .B2(keyinput6), .ZN(n6694) );
  AOI221_X1 U7624 ( .B1(ADDRESS_REG_24__SCAN_IN), .B2(keyinput19), .C1(
        keyinput6), .C2(FLUSH_REG_SCAN_IN), .A(n6694), .ZN(n6699) );
  OAI22_X1 U7625 ( .A1(ADDRESS_REG_19__SCAN_IN), .A2(keyinput44), .B1(
        keyinput57), .B2(DATAI_13_), .ZN(n6695) );
  AOI221_X1 U7626 ( .B1(ADDRESS_REG_19__SCAN_IN), .B2(keyinput44), .C1(
        DATAI_13_), .C2(keyinput57), .A(n6695), .ZN(n6698) );
  OAI22_X1 U7627 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(keyinput20), .B1(
        keyinput16), .B2(UWORD_REG_8__SCAN_IN), .ZN(n6696) );
  AOI221_X1 U7628 ( .B1(INSTQUEUE_REG_12__0__SCAN_IN), .B2(keyinput20), .C1(
        UWORD_REG_8__SCAN_IN), .C2(keyinput16), .A(n6696), .ZN(n6697) );
  NAND4_X1 U7629 ( .A1(n6700), .A2(n6699), .A3(n6698), .A4(n6697), .ZN(n6710)
         );
  OAI22_X1 U7630 ( .A1(EAX_REG_29__SCAN_IN), .A2(keyinput37), .B1(keyinput32), 
        .B2(UWORD_REG_12__SCAN_IN), .ZN(n6701) );
  AOI221_X1 U7631 ( .B1(EAX_REG_29__SCAN_IN), .B2(keyinput37), .C1(
        UWORD_REG_12__SCAN_IN), .C2(keyinput32), .A(n6701), .ZN(n6708) );
  OAI22_X1 U7632 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(keyinput36), .B1(
        EAX_REG_12__SCAN_IN), .B2(keyinput51), .ZN(n6702) );
  AOI221_X1 U7633 ( .B1(INSTQUEUE_REG_0__4__SCAN_IN), .B2(keyinput36), .C1(
        keyinput51), .C2(EAX_REG_12__SCAN_IN), .A(n6702), .ZN(n6707) );
  OAI22_X1 U7634 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(keyinput47), .B1(
        INSTQUEUE_REG_11__6__SCAN_IN), .B2(keyinput31), .ZN(n6703) );
  AOI221_X1 U7635 ( .B1(INSTQUEUE_REG_15__1__SCAN_IN), .B2(keyinput47), .C1(
        keyinput31), .C2(INSTQUEUE_REG_11__6__SCAN_IN), .A(n6703), .ZN(n6706)
         );
  OAI22_X1 U7636 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(keyinput55), .B1(
        keyinput38), .B2(ADDRESS_REG_17__SCAN_IN), .ZN(n6704) );
  AOI221_X1 U7637 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(keyinput55), .C1(
        ADDRESS_REG_17__SCAN_IN), .C2(keyinput38), .A(n6704), .ZN(n6705) );
  NAND4_X1 U7638 ( .A1(n6708), .A2(n6707), .A3(n6706), .A4(n6705), .ZN(n6709)
         );
  NOR4_X1 U7639 ( .A1(n6712), .A2(n6711), .A3(n6710), .A4(n6709), .ZN(n6780)
         );
  AOI22_X1 U7640 ( .A1(n6715), .A2(keyinput48), .B1(keyinput9), .B2(n6714), 
        .ZN(n6713) );
  OAI221_X1 U7641 ( .B1(n6715), .B2(keyinput48), .C1(n6714), .C2(keyinput9), 
        .A(n6713), .ZN(n6728) );
  INV_X1 U7642 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n6718) );
  AOI22_X1 U7643 ( .A1(n6718), .A2(keyinput59), .B1(keyinput2), .B2(n6717), 
        .ZN(n6716) );
  OAI221_X1 U7644 ( .B1(n6718), .B2(keyinput59), .C1(n6717), .C2(keyinput2), 
        .A(n6716), .ZN(n6727) );
  INV_X1 U7645 ( .A(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n6721) );
  AOI22_X1 U7646 ( .A1(n6721), .A2(keyinput42), .B1(keyinput10), .B2(n6720), 
        .ZN(n6719) );
  OAI221_X1 U7647 ( .B1(n6721), .B2(keyinput42), .C1(n6720), .C2(keyinput10), 
        .A(n6719), .ZN(n6726) );
  AOI22_X1 U7648 ( .A1(n6724), .A2(keyinput49), .B1(n6723), .B2(keyinput1), 
        .ZN(n6722) );
  OAI221_X1 U7649 ( .B1(n6724), .B2(keyinput49), .C1(n6723), .C2(keyinput1), 
        .A(n6722), .ZN(n6725) );
  NOR4_X1 U7650 ( .A1(n6728), .A2(n6727), .A3(n6726), .A4(n6725), .ZN(n6778)
         );
  AOI22_X1 U7651 ( .A1(n6731), .A2(keyinput54), .B1(keyinput41), .B2(n6730), 
        .ZN(n6729) );
  OAI221_X1 U7652 ( .B1(n6731), .B2(keyinput54), .C1(n6730), .C2(keyinput41), 
        .A(n6729), .ZN(n6742) );
  AOI22_X1 U7653 ( .A1(DATAWIDTH_REG_20__SCAN_IN), .A2(keyinput56), .B1(
        STATE2_REG_0__SCAN_IN), .B2(keyinput26), .ZN(n6732) );
  OAI221_X1 U7654 ( .B1(DATAWIDTH_REG_20__SCAN_IN), .B2(keyinput56), .C1(
        STATE2_REG_0__SCAN_IN), .C2(keyinput26), .A(n6732), .ZN(n6741) );
  AOI22_X1 U7655 ( .A1(n6735), .A2(keyinput58), .B1(n6734), .B2(keyinput24), 
        .ZN(n6733) );
  OAI221_X1 U7656 ( .B1(n6735), .B2(keyinput58), .C1(n6734), .C2(keyinput24), 
        .A(n6733), .ZN(n6740) );
  AOI22_X1 U7657 ( .A1(n6738), .A2(keyinput8), .B1(n6737), .B2(keyinput62), 
        .ZN(n6736) );
  OAI221_X1 U7658 ( .B1(n6738), .B2(keyinput8), .C1(n6737), .C2(keyinput62), 
        .A(n6736), .ZN(n6739) );
  NOR4_X1 U7659 ( .A1(n6742), .A2(n6741), .A3(n6740), .A4(n6739), .ZN(n6777)
         );
  AOI22_X1 U7660 ( .A1(n6745), .A2(keyinput28), .B1(n6744), .B2(keyinput34), 
        .ZN(n6743) );
  OAI221_X1 U7661 ( .B1(n6745), .B2(keyinput28), .C1(n6744), .C2(keyinput34), 
        .A(n6743), .ZN(n6758) );
  AOI22_X1 U7662 ( .A1(n6748), .A2(keyinput12), .B1(keyinput13), .B2(n6747), 
        .ZN(n6746) );
  OAI221_X1 U7663 ( .B1(n6748), .B2(keyinput12), .C1(n6747), .C2(keyinput13), 
        .A(n6746), .ZN(n6757) );
  AOI22_X1 U7664 ( .A1(n6751), .A2(keyinput52), .B1(n6750), .B2(keyinput23), 
        .ZN(n6749) );
  OAI221_X1 U7665 ( .B1(n6751), .B2(keyinput52), .C1(n6750), .C2(keyinput23), 
        .A(n6749), .ZN(n6756) );
  AOI22_X1 U7666 ( .A1(n6754), .A2(keyinput14), .B1(keyinput45), .B2(n6753), 
        .ZN(n6752) );
  OAI221_X1 U7667 ( .B1(n6754), .B2(keyinput14), .C1(n6753), .C2(keyinput45), 
        .A(n6752), .ZN(n6755) );
  NOR4_X1 U7668 ( .A1(n6758), .A2(n6757), .A3(n6756), .A4(n6755), .ZN(n6776)
         );
  AOI22_X1 U7669 ( .A1(n6761), .A2(keyinput3), .B1(n6760), .B2(keyinput7), 
        .ZN(n6759) );
  OAI221_X1 U7670 ( .B1(n6761), .B2(keyinput3), .C1(n6760), .C2(keyinput7), 
        .A(n6759), .ZN(n6774) );
  INV_X1 U7671 ( .A(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n6764) );
  AOI22_X1 U7672 ( .A1(n6764), .A2(keyinput30), .B1(keyinput40), .B2(n6763), 
        .ZN(n6762) );
  OAI221_X1 U7673 ( .B1(n6764), .B2(keyinput30), .C1(n6763), .C2(keyinput40), 
        .A(n6762), .ZN(n6773) );
  AOI22_X1 U7674 ( .A1(n6767), .A2(keyinput35), .B1(n6766), .B2(keyinput15), 
        .ZN(n6765) );
  OAI221_X1 U7675 ( .B1(n6767), .B2(keyinput35), .C1(n6766), .C2(keyinput15), 
        .A(n6765), .ZN(n6772) );
  AOI22_X1 U7676 ( .A1(n6770), .A2(keyinput46), .B1(n6769), .B2(keyinput53), 
        .ZN(n6768) );
  OAI221_X1 U7677 ( .B1(n6770), .B2(keyinput46), .C1(n6769), .C2(keyinput53), 
        .A(n6768), .ZN(n6771) );
  NOR4_X1 U7678 ( .A1(n6774), .A2(n6773), .A3(n6772), .A4(n6771), .ZN(n6775)
         );
  AND4_X1 U7679 ( .A1(n6778), .A2(n6777), .A3(n6776), .A4(n6775), .ZN(n6779)
         );
  OAI211_X1 U7680 ( .C1(n6782), .C2(n6781), .A(n6780), .B(n6779), .ZN(n6783)
         );
  XNOR2_X1 U7681 ( .A(n6784), .B(n6783), .ZN(U3000) );
  INV_X2 U3457 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6596) );
  CLKBUF_X1 U34620 ( .A(n3177), .Z(n4238) );
  CLKBUF_X1 U34690 ( .A(n5572), .Z(n5580) );
  AND2_X2 U3721 ( .A1(n4369), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4367)
         );
endmodule

