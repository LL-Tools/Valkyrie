

module b15_C_2inp_gates_syn ( DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, 
        DATAI_27_, DATAI_26_, DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, 
        DATAI_21_, DATAI_20_, DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, 
        DATAI_15_, DATAI_14_, DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, 
        DATAI_9_, DATAI_8_, DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, 
        DATAI_2_, DATAI_1_, DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, 
        READY_N, HOLD, READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, 
        CODEFETCH_REG_SCAN_IN, M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, 
        REQUESTPENDING_REG_SCAN_IN, STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, 
        FLUSH_REG_SCAN_IN, W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN, 
        BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN, 
        BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN, 
        REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN, 
        REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN, 
        REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN, 
        REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN, 
        REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN, 
        BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN, 
        ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN, 
        ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN, 
        ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN, 
        ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN, 
        ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN, 
        ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN, 
        ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN, 
        ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN, 
        ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN, 
        ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN, 
        ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN, ADDRESS_REG_7__SCAN_IN, 
        ADDRESS_REG_6__SCAN_IN, ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN, 
        ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN, ADDRESS_REG_1__SCAN_IN, 
        ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN, STATE_REG_1__SCAN_IN, 
        STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN, 
        DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN, 
        DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN, 
        DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN, 
        DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN, 
        DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN, 
        DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN, 
        DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN, 
        DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN, 
        DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN, 
        DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN, 
        DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN, 
        DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN, 
        DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN, 
        DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN, 
        DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN, 
        DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN, 
        STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN, 
        INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN, 
        INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN, 
        INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN, 
        INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN, 
        INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN, 
        INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN, 
        INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN, 
        INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN, 
        INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN, 
        INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN, 
        INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN, 
        INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN, 
        INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN, 
        INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN, 
        INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN, 
        INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN, 
        INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN, 
        INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN, 
        INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN, 
        INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN, 
        INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN, 
        INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN, 
        INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN, 
        INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN, 
        INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN, 
        INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN, 
        INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN, 
        INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN, 
        INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN, 
        INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN, 
        INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN, 
        INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN, 
        INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN, 
        INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN, 
        INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN, 
        INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN, 
        INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN, 
        INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN, 
        INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN, 
        INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN, 
        INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN, 
        INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN, 
        INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN, 
        INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN, 
        INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN, 
        INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN, 
        INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN, 
        INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN, 
        INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN, 
        INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN, 
        INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN, 
        INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN, 
        INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN, 
        INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN, 
        INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN, 
        INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN, 
        INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN, 
        INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN, 
        INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN, 
        INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN, 
        INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN, 
        INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN, 
        INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN, 
        INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN, 
        INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN, 
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN, 
        INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN, 
        INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN, 
        INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN, 
        INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN, 
        INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN, 
        INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN, 
        INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN, 
        INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN, 
        INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN, 
        INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN, 
        INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN, 
        INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN, 
        INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN, 
        INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN, 
        INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN, 
        INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN, 
        PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN, 
        PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN, 
        PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN, 
        PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN, 
        PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN, 
        PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN, 
        PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN, 
        PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN, 
        PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN, 
        PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN, 
        PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN, 
        PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN, 
        PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN, 
        PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN, 
        PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN, 
        PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN, 
        LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN, 
        LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN, 
        LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN, 
        LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN, 
        LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN, 
        LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN, 
        UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN, 
        UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN, 
        UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN, 
        UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN, 
        UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN, 
        DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN, 
        DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN, 
        DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN, 
        DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN, 
        DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN, 
        DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN, 
        DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN, 
        DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN, 
        DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN, 
        DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN, 
        EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN, 
        EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN, 
        EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN, 
        EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN, 
        EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN, 
        EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN, 
        EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN, 
        EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN, 
        EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN, 
        EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN, 
        EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN, 
        EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN, 
        EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN, 
        EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN, 
        EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN, 
        EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN, 
        EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN, 
        EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN, 
        EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN, 
        EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN, 
        EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN, 
        EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN, 
        REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN, 
        REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN, 
        REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN, 
        REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN, 
        REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, U3445, U3446, U3447, U3448, 
        U3213, U3212, U3211, U3210, U3209, U3208, U3207, U3206, U3205, U3204, 
        U3203, U3202, U3201, U3200, U3199, U3198, U3197, U3196, U3195, U3194, 
        U3193, U3192, U3191, U3190, U3189, U3188, U3187, U3186, U3185, U3184, 
        U3183, U3182, U3181, U3451, U3452, U3180, U3179, U3178, U3177, U3176, 
        U3175, U3174, U3173, U3172, U3171, U3170, U3169, U3168, U3167, U3166, 
        U3165, U3164, U3163, U3162, U3161, U3160, U3159, U3158, U3157, U3156, 
        U3155, U3154, U3153, U3152, U3151, U3453, U3150, U3149, U3148, U3147, 
        U3146, U3145, U3144, U3143, U3142, U3141, U3140, U3139, U3138, U3137, 
        U3136, U3135, U3134, U3133, U3132, U3131, U3130, U3129, U3128, U3127, 
        U3126, U3125, U3124, U3123, U3122, U3121, U3120, U3119, U3118, U3117, 
        U3116, U3115, U3114, U3113, U3112, U3111, U3110, U3109, U3108, U3107, 
        U3106, U3105, U3104, U3103, U3102, U3101, U3100, U3099, U3098, U3097, 
        U3096, U3095, U3094, U3093, U3092, U3091, U3090, U3089, U3088, U3087, 
        U3086, U3085, U3084, U3083, U3082, U3081, U3080, U3079, U3078, U3077, 
        U3076, U3075, U3074, U3073, U3072, U3071, U3070, U3069, U3068, U3067, 
        U3066, U3065, U3064, U3063, U3062, U3061, U3060, U3059, U3058, U3057, 
        U3056, U3055, U3054, U3053, U3052, U3051, U3050, U3049, U3048, U3047, 
        U3046, U3045, U3044, U3043, U3042, U3041, U3040, U3039, U3038, U3037, 
        U3036, U3035, U3034, U3033, U3032, U3031, U3030, U3029, U3028, U3027, 
        U3026, U3025, U3024, U3023, U3022, U3021, U3020, U3455, U3456, U3459, 
        U3460, U3461, U3019, U3462, U3463, U3464, U3465, U3018, U3017, U3016, 
        U3015, U3014, U3013, U3012, U3011, U3010, U3009, U3008, U3007, U3006, 
        U3005, U3004, U3003, U3002, U3001, U3000, U2999, U2998, U2997, U2996, 
        U2995, U2994, U2993, U2992, U2991, U2990, U2989, U2988, U2987, U2986, 
        U2985, U2984, U2983, U2982, U2981, U2980, U2979, U2978, U2977, U2976, 
        U2975, U2974, U2973, U2972, U2971, U2970, U2969, U2968, U2967, U2966, 
        U2965, U2964, U2963, U2962, U2961, U2960, U2959, U2958, U2957, U2956, 
        U2955, U2954, U2953, U2952, U2951, U2950, U2949, U2948, U2947, U2946, 
        U2945, U2944, U2943, U2942, U2941, U2940, U2939, U2938, U2937, U2936, 
        U2935, U2934, U2933, U2932, U2931, U2930, U2929, U2928, U2927, U2926, 
        U2925, U2924, U2923, U2922, U2921, U2920, U2919, U2918, U2917, U2916, 
        U2915, U2914, U2913, U2912, U2911, U2910, U2909, U2908, U2907, U2906, 
        U2905, U2904, U2903, U2902, U2901, U2900, U2899, U2898, U2897, U2896, 
        U2895, U2894, U2893, U2892, U2891, U2890, U2889, U2888, U2887, U2886, 
        U2885, U2884, U2883, U2882, U2881, U2880, U2879, U2878, U2877, U2876, 
        U2875, U2874, U2873, U2872, U2871, U2870, U2869, U2868, U2867, U2866, 
        U2865, U2864, U2863, U2862, U2861, U2860, U2859, U2858, U2857, U2856, 
        U2855, U2854, U2853, U2852, U2851, U2850, U2849, U2848, U2847, U2846, 
        U2845, U2844, U2843, U2842, U2841, U2840, U2839, U2838, U2837, U2836, 
        U2835, U2834, U2833, U2832, U2831, U2830, U2829, U2828, U2827, U2826, 
        U2825, U2824, U2823, U2822, U2821, U2820, U2819, U2818, U2817, U2816, 
        U2815, U2814, U2813, U2812, U2811, U2810, U2809, U2808, U2807, U2806, 
        U2805, U2804, U2803, U2802, U2801, U2800, U2799, U2798, U2797, U2796, 
        U2795, U3468, U2794, U3469, U3470, U2793, U3471, U2792, U3472, U2791, 
        U3473, U2790, U2789, U3474, U2788, keyinput127, keyinput126, 
        keyinput125, keyinput124, keyinput123, keyinput122, keyinput121, 
        keyinput120, keyinput119, keyinput118, keyinput117, keyinput116, 
        keyinput115, keyinput114, keyinput113, keyinput112, keyinput111, 
        keyinput110, keyinput109, keyinput108, keyinput107, keyinput106, 
        keyinput105, keyinput104, keyinput103, keyinput102, keyinput101, 
        keyinput100, keyinput99, keyinput98, keyinput97, keyinput96, 
        keyinput95, keyinput94, keyinput93, keyinput92, keyinput91, keyinput90, 
        keyinput89, keyinput88, keyinput87, keyinput86, keyinput85, keyinput84, 
        keyinput83, keyinput82, keyinput81, keyinput80, keyinput79, keyinput78, 
        keyinput77, keyinput76, keyinput75, keyinput74, keyinput73, keyinput72, 
        keyinput71, keyinput70, keyinput69, keyinput68, keyinput67, keyinput66, 
        keyinput65, keyinput64, keyinput63, keyinput62, keyinput61, keyinput60, 
        keyinput59, keyinput58, keyinput57, keyinput56, keyinput55, keyinput54, 
        keyinput53, keyinput52, keyinput51, keyinput50, keyinput49, keyinput48, 
        keyinput47, keyinput46, keyinput45, keyinput44, keyinput43, keyinput42, 
        keyinput41, keyinput40, keyinput39, keyinput38, keyinput37, keyinput36, 
        keyinput35, keyinput34, keyinput33, keyinput32, keyinput31, keyinput30, 
        keyinput29, keyinput28, keyinput27, keyinput26, keyinput25, keyinput24, 
        keyinput23, keyinput22, keyinput21, keyinput20, keyinput19, keyinput18, 
        keyinput17, keyinput16, keyinput15, keyinput14, keyinput13, keyinput12, 
        keyinput11, keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, 
        keyinput5, keyinput4, keyinput3, keyinput2, keyinput1, keyinput0 );
  input DATAI_31_, DATAI_30_, DATAI_29_, DATAI_28_, DATAI_27_, DATAI_26_,
         DATAI_25_, DATAI_24_, DATAI_23_, DATAI_22_, DATAI_21_, DATAI_20_,
         DATAI_19_, DATAI_18_, DATAI_17_, DATAI_16_, DATAI_15_, DATAI_14_,
         DATAI_13_, DATAI_12_, DATAI_11_, DATAI_10_, DATAI_9_, DATAI_8_,
         DATAI_7_, DATAI_6_, DATAI_5_, DATAI_4_, DATAI_3_, DATAI_2_, DATAI_1_,
         DATAI_0_, MEMORYFETCH_REG_SCAN_IN, NA_N, BS16_N, READY_N, HOLD,
         READREQUEST_REG_SCAN_IN, ADS_N_REG_SCAN_IN, CODEFETCH_REG_SCAN_IN,
         M_IO_N_REG_SCAN_IN, D_C_N_REG_SCAN_IN, REQUESTPENDING_REG_SCAN_IN,
         STATEBS16_REG_SCAN_IN, MORE_REG_SCAN_IN, FLUSH_REG_SCAN_IN,
         W_R_N_REG_SCAN_IN, BYTEENABLE_REG_0__SCAN_IN,
         BYTEENABLE_REG_1__SCAN_IN, BYTEENABLE_REG_2__SCAN_IN,
         BYTEENABLE_REG_3__SCAN_IN, REIP_REG_31__SCAN_IN, REIP_REG_30__SCAN_IN,
         REIP_REG_29__SCAN_IN, REIP_REG_28__SCAN_IN, REIP_REG_27__SCAN_IN,
         REIP_REG_26__SCAN_IN, REIP_REG_25__SCAN_IN, REIP_REG_24__SCAN_IN,
         REIP_REG_23__SCAN_IN, REIP_REG_22__SCAN_IN, REIP_REG_21__SCAN_IN,
         REIP_REG_20__SCAN_IN, REIP_REG_19__SCAN_IN, REIP_REG_18__SCAN_IN,
         REIP_REG_17__SCAN_IN, REIP_REG_16__SCAN_IN, BE_N_REG_3__SCAN_IN,
         BE_N_REG_2__SCAN_IN, BE_N_REG_1__SCAN_IN, BE_N_REG_0__SCAN_IN,
         ADDRESS_REG_29__SCAN_IN, ADDRESS_REG_28__SCAN_IN,
         ADDRESS_REG_27__SCAN_IN, ADDRESS_REG_26__SCAN_IN,
         ADDRESS_REG_25__SCAN_IN, ADDRESS_REG_24__SCAN_IN,
         ADDRESS_REG_23__SCAN_IN, ADDRESS_REG_22__SCAN_IN,
         ADDRESS_REG_21__SCAN_IN, ADDRESS_REG_20__SCAN_IN,
         ADDRESS_REG_19__SCAN_IN, ADDRESS_REG_18__SCAN_IN,
         ADDRESS_REG_17__SCAN_IN, ADDRESS_REG_16__SCAN_IN,
         ADDRESS_REG_15__SCAN_IN, ADDRESS_REG_14__SCAN_IN,
         ADDRESS_REG_13__SCAN_IN, ADDRESS_REG_12__SCAN_IN,
         ADDRESS_REG_11__SCAN_IN, ADDRESS_REG_10__SCAN_IN,
         ADDRESS_REG_9__SCAN_IN, ADDRESS_REG_8__SCAN_IN,
         ADDRESS_REG_7__SCAN_IN, ADDRESS_REG_6__SCAN_IN,
         ADDRESS_REG_5__SCAN_IN, ADDRESS_REG_4__SCAN_IN,
         ADDRESS_REG_3__SCAN_IN, ADDRESS_REG_2__SCAN_IN,
         ADDRESS_REG_1__SCAN_IN, ADDRESS_REG_0__SCAN_IN, STATE_REG_2__SCAN_IN,
         STATE_REG_1__SCAN_IN, STATE_REG_0__SCAN_IN, DATAWIDTH_REG_0__SCAN_IN,
         DATAWIDTH_REG_1__SCAN_IN, DATAWIDTH_REG_2__SCAN_IN,
         DATAWIDTH_REG_3__SCAN_IN, DATAWIDTH_REG_4__SCAN_IN,
         DATAWIDTH_REG_5__SCAN_IN, DATAWIDTH_REG_6__SCAN_IN,
         DATAWIDTH_REG_7__SCAN_IN, DATAWIDTH_REG_8__SCAN_IN,
         DATAWIDTH_REG_9__SCAN_IN, DATAWIDTH_REG_10__SCAN_IN,
         DATAWIDTH_REG_11__SCAN_IN, DATAWIDTH_REG_12__SCAN_IN,
         DATAWIDTH_REG_13__SCAN_IN, DATAWIDTH_REG_14__SCAN_IN,
         DATAWIDTH_REG_15__SCAN_IN, DATAWIDTH_REG_16__SCAN_IN,
         DATAWIDTH_REG_17__SCAN_IN, DATAWIDTH_REG_18__SCAN_IN,
         DATAWIDTH_REG_19__SCAN_IN, DATAWIDTH_REG_20__SCAN_IN,
         DATAWIDTH_REG_21__SCAN_IN, DATAWIDTH_REG_22__SCAN_IN,
         DATAWIDTH_REG_23__SCAN_IN, DATAWIDTH_REG_24__SCAN_IN,
         DATAWIDTH_REG_25__SCAN_IN, DATAWIDTH_REG_26__SCAN_IN,
         DATAWIDTH_REG_27__SCAN_IN, DATAWIDTH_REG_28__SCAN_IN,
         DATAWIDTH_REG_29__SCAN_IN, DATAWIDTH_REG_30__SCAN_IN,
         DATAWIDTH_REG_31__SCAN_IN, STATE2_REG_3__SCAN_IN,
         STATE2_REG_2__SCAN_IN, STATE2_REG_1__SCAN_IN, STATE2_REG_0__SCAN_IN,
         INSTQUEUE_REG_15__7__SCAN_IN, INSTQUEUE_REG_15__6__SCAN_IN,
         INSTQUEUE_REG_15__5__SCAN_IN, INSTQUEUE_REG_15__4__SCAN_IN,
         INSTQUEUE_REG_15__3__SCAN_IN, INSTQUEUE_REG_15__2__SCAN_IN,
         INSTQUEUE_REG_15__1__SCAN_IN, INSTQUEUE_REG_15__0__SCAN_IN,
         INSTQUEUE_REG_14__7__SCAN_IN, INSTQUEUE_REG_14__6__SCAN_IN,
         INSTQUEUE_REG_14__5__SCAN_IN, INSTQUEUE_REG_14__4__SCAN_IN,
         INSTQUEUE_REG_14__3__SCAN_IN, INSTQUEUE_REG_14__2__SCAN_IN,
         INSTQUEUE_REG_14__1__SCAN_IN, INSTQUEUE_REG_14__0__SCAN_IN,
         INSTQUEUE_REG_13__7__SCAN_IN, INSTQUEUE_REG_13__6__SCAN_IN,
         INSTQUEUE_REG_13__5__SCAN_IN, INSTQUEUE_REG_13__4__SCAN_IN,
         INSTQUEUE_REG_13__3__SCAN_IN, INSTQUEUE_REG_13__2__SCAN_IN,
         INSTQUEUE_REG_13__1__SCAN_IN, INSTQUEUE_REG_13__0__SCAN_IN,
         INSTQUEUE_REG_12__7__SCAN_IN, INSTQUEUE_REG_12__6__SCAN_IN,
         INSTQUEUE_REG_12__5__SCAN_IN, INSTQUEUE_REG_12__4__SCAN_IN,
         INSTQUEUE_REG_12__3__SCAN_IN, INSTQUEUE_REG_12__2__SCAN_IN,
         INSTQUEUE_REG_12__1__SCAN_IN, INSTQUEUE_REG_12__0__SCAN_IN,
         INSTQUEUE_REG_11__7__SCAN_IN, INSTQUEUE_REG_11__6__SCAN_IN,
         INSTQUEUE_REG_11__5__SCAN_IN, INSTQUEUE_REG_11__4__SCAN_IN,
         INSTQUEUE_REG_11__3__SCAN_IN, INSTQUEUE_REG_11__2__SCAN_IN,
         INSTQUEUE_REG_11__1__SCAN_IN, INSTQUEUE_REG_11__0__SCAN_IN,
         INSTQUEUE_REG_10__7__SCAN_IN, INSTQUEUE_REG_10__6__SCAN_IN,
         INSTQUEUE_REG_10__5__SCAN_IN, INSTQUEUE_REG_10__4__SCAN_IN,
         INSTQUEUE_REG_10__3__SCAN_IN, INSTQUEUE_REG_10__2__SCAN_IN,
         INSTQUEUE_REG_10__1__SCAN_IN, INSTQUEUE_REG_10__0__SCAN_IN,
         INSTQUEUE_REG_9__7__SCAN_IN, INSTQUEUE_REG_9__6__SCAN_IN,
         INSTQUEUE_REG_9__5__SCAN_IN, INSTQUEUE_REG_9__4__SCAN_IN,
         INSTQUEUE_REG_9__3__SCAN_IN, INSTQUEUE_REG_9__2__SCAN_IN,
         INSTQUEUE_REG_9__1__SCAN_IN, INSTQUEUE_REG_9__0__SCAN_IN,
         INSTQUEUE_REG_8__7__SCAN_IN, INSTQUEUE_REG_8__6__SCAN_IN,
         INSTQUEUE_REG_8__5__SCAN_IN, INSTQUEUE_REG_8__4__SCAN_IN,
         INSTQUEUE_REG_8__3__SCAN_IN, INSTQUEUE_REG_8__2__SCAN_IN,
         INSTQUEUE_REG_8__1__SCAN_IN, INSTQUEUE_REG_8__0__SCAN_IN,
         INSTQUEUE_REG_7__7__SCAN_IN, INSTQUEUE_REG_7__6__SCAN_IN,
         INSTQUEUE_REG_7__5__SCAN_IN, INSTQUEUE_REG_7__4__SCAN_IN,
         INSTQUEUE_REG_7__3__SCAN_IN, INSTQUEUE_REG_7__2__SCAN_IN,
         INSTQUEUE_REG_7__1__SCAN_IN, INSTQUEUE_REG_7__0__SCAN_IN,
         INSTQUEUE_REG_6__7__SCAN_IN, INSTQUEUE_REG_6__6__SCAN_IN,
         INSTQUEUE_REG_6__5__SCAN_IN, INSTQUEUE_REG_6__4__SCAN_IN,
         INSTQUEUE_REG_6__3__SCAN_IN, INSTQUEUE_REG_6__2__SCAN_IN,
         INSTQUEUE_REG_6__1__SCAN_IN, INSTQUEUE_REG_6__0__SCAN_IN,
         INSTQUEUE_REG_5__7__SCAN_IN, INSTQUEUE_REG_5__6__SCAN_IN,
         INSTQUEUE_REG_5__5__SCAN_IN, INSTQUEUE_REG_5__4__SCAN_IN,
         INSTQUEUE_REG_5__3__SCAN_IN, INSTQUEUE_REG_5__2__SCAN_IN,
         INSTQUEUE_REG_5__1__SCAN_IN, INSTQUEUE_REG_5__0__SCAN_IN,
         INSTQUEUE_REG_4__7__SCAN_IN, INSTQUEUE_REG_4__6__SCAN_IN,
         INSTQUEUE_REG_4__5__SCAN_IN, INSTQUEUE_REG_4__4__SCAN_IN,
         INSTQUEUE_REG_4__3__SCAN_IN, INSTQUEUE_REG_4__2__SCAN_IN,
         INSTQUEUE_REG_4__1__SCAN_IN, INSTQUEUE_REG_4__0__SCAN_IN,
         INSTQUEUE_REG_3__7__SCAN_IN, INSTQUEUE_REG_3__6__SCAN_IN,
         INSTQUEUE_REG_3__5__SCAN_IN, INSTQUEUE_REG_3__4__SCAN_IN,
         INSTQUEUE_REG_3__3__SCAN_IN, INSTQUEUE_REG_3__2__SCAN_IN,
         INSTQUEUE_REG_3__1__SCAN_IN, INSTQUEUE_REG_3__0__SCAN_IN,
         INSTQUEUE_REG_2__7__SCAN_IN, INSTQUEUE_REG_2__6__SCAN_IN,
         INSTQUEUE_REG_2__5__SCAN_IN, INSTQUEUE_REG_2__4__SCAN_IN,
         INSTQUEUE_REG_2__3__SCAN_IN, INSTQUEUE_REG_2__2__SCAN_IN,
         INSTQUEUE_REG_2__1__SCAN_IN, INSTQUEUE_REG_2__0__SCAN_IN,
         INSTQUEUE_REG_1__7__SCAN_IN, INSTQUEUE_REG_1__6__SCAN_IN,
         INSTQUEUE_REG_1__5__SCAN_IN, INSTQUEUE_REG_1__4__SCAN_IN,
         INSTQUEUE_REG_1__3__SCAN_IN, INSTQUEUE_REG_1__2__SCAN_IN,
         INSTQUEUE_REG_1__1__SCAN_IN, INSTQUEUE_REG_1__0__SCAN_IN,
         INSTQUEUE_REG_0__7__SCAN_IN, INSTQUEUE_REG_0__6__SCAN_IN,
         INSTQUEUE_REG_0__5__SCAN_IN, INSTQUEUE_REG_0__4__SCAN_IN,
         INSTQUEUE_REG_0__3__SCAN_IN, INSTQUEUE_REG_0__2__SCAN_IN,
         INSTQUEUE_REG_0__1__SCAN_IN, INSTQUEUE_REG_0__0__SCAN_IN,
         INSTQUEUERD_ADDR_REG_4__SCAN_IN, INSTQUEUERD_ADDR_REG_3__SCAN_IN,
         INSTQUEUERD_ADDR_REG_2__SCAN_IN, INSTQUEUERD_ADDR_REG_1__SCAN_IN,
         INSTQUEUERD_ADDR_REG_0__SCAN_IN, INSTQUEUEWR_ADDR_REG_4__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_3__SCAN_IN, INSTQUEUEWR_ADDR_REG_2__SCAN_IN,
         INSTQUEUEWR_ADDR_REG_1__SCAN_IN, INSTQUEUEWR_ADDR_REG_0__SCAN_IN,
         INSTADDRPOINTER_REG_0__SCAN_IN, INSTADDRPOINTER_REG_1__SCAN_IN,
         INSTADDRPOINTER_REG_2__SCAN_IN, INSTADDRPOINTER_REG_3__SCAN_IN,
         INSTADDRPOINTER_REG_4__SCAN_IN, INSTADDRPOINTER_REG_5__SCAN_IN,
         INSTADDRPOINTER_REG_6__SCAN_IN, INSTADDRPOINTER_REG_7__SCAN_IN,
         INSTADDRPOINTER_REG_8__SCAN_IN, INSTADDRPOINTER_REG_9__SCAN_IN,
         INSTADDRPOINTER_REG_10__SCAN_IN, INSTADDRPOINTER_REG_11__SCAN_IN,
         INSTADDRPOINTER_REG_12__SCAN_IN, INSTADDRPOINTER_REG_13__SCAN_IN,
         INSTADDRPOINTER_REG_14__SCAN_IN, INSTADDRPOINTER_REG_15__SCAN_IN,
         INSTADDRPOINTER_REG_16__SCAN_IN, INSTADDRPOINTER_REG_17__SCAN_IN,
         INSTADDRPOINTER_REG_18__SCAN_IN, INSTADDRPOINTER_REG_19__SCAN_IN,
         INSTADDRPOINTER_REG_20__SCAN_IN, INSTADDRPOINTER_REG_21__SCAN_IN,
         INSTADDRPOINTER_REG_22__SCAN_IN, INSTADDRPOINTER_REG_23__SCAN_IN,
         INSTADDRPOINTER_REG_24__SCAN_IN, INSTADDRPOINTER_REG_25__SCAN_IN,
         INSTADDRPOINTER_REG_26__SCAN_IN, INSTADDRPOINTER_REG_27__SCAN_IN,
         INSTADDRPOINTER_REG_28__SCAN_IN, INSTADDRPOINTER_REG_29__SCAN_IN,
         INSTADDRPOINTER_REG_30__SCAN_IN, INSTADDRPOINTER_REG_31__SCAN_IN,
         PHYADDRPOINTER_REG_0__SCAN_IN, PHYADDRPOINTER_REG_1__SCAN_IN,
         PHYADDRPOINTER_REG_2__SCAN_IN, PHYADDRPOINTER_REG_3__SCAN_IN,
         PHYADDRPOINTER_REG_4__SCAN_IN, PHYADDRPOINTER_REG_5__SCAN_IN,
         PHYADDRPOINTER_REG_6__SCAN_IN, PHYADDRPOINTER_REG_7__SCAN_IN,
         PHYADDRPOINTER_REG_8__SCAN_IN, PHYADDRPOINTER_REG_9__SCAN_IN,
         PHYADDRPOINTER_REG_10__SCAN_IN, PHYADDRPOINTER_REG_11__SCAN_IN,
         PHYADDRPOINTER_REG_12__SCAN_IN, PHYADDRPOINTER_REG_13__SCAN_IN,
         PHYADDRPOINTER_REG_14__SCAN_IN, PHYADDRPOINTER_REG_15__SCAN_IN,
         PHYADDRPOINTER_REG_16__SCAN_IN, PHYADDRPOINTER_REG_17__SCAN_IN,
         PHYADDRPOINTER_REG_18__SCAN_IN, PHYADDRPOINTER_REG_19__SCAN_IN,
         PHYADDRPOINTER_REG_20__SCAN_IN, PHYADDRPOINTER_REG_21__SCAN_IN,
         PHYADDRPOINTER_REG_22__SCAN_IN, PHYADDRPOINTER_REG_23__SCAN_IN,
         PHYADDRPOINTER_REG_24__SCAN_IN, PHYADDRPOINTER_REG_25__SCAN_IN,
         PHYADDRPOINTER_REG_26__SCAN_IN, PHYADDRPOINTER_REG_27__SCAN_IN,
         PHYADDRPOINTER_REG_28__SCAN_IN, PHYADDRPOINTER_REG_29__SCAN_IN,
         PHYADDRPOINTER_REG_30__SCAN_IN, PHYADDRPOINTER_REG_31__SCAN_IN,
         LWORD_REG_15__SCAN_IN, LWORD_REG_14__SCAN_IN, LWORD_REG_13__SCAN_IN,
         LWORD_REG_12__SCAN_IN, LWORD_REG_11__SCAN_IN, LWORD_REG_10__SCAN_IN,
         LWORD_REG_9__SCAN_IN, LWORD_REG_8__SCAN_IN, LWORD_REG_7__SCAN_IN,
         LWORD_REG_6__SCAN_IN, LWORD_REG_5__SCAN_IN, LWORD_REG_4__SCAN_IN,
         LWORD_REG_3__SCAN_IN, LWORD_REG_2__SCAN_IN, LWORD_REG_1__SCAN_IN,
         LWORD_REG_0__SCAN_IN, UWORD_REG_14__SCAN_IN, UWORD_REG_13__SCAN_IN,
         UWORD_REG_12__SCAN_IN, UWORD_REG_11__SCAN_IN, UWORD_REG_10__SCAN_IN,
         UWORD_REG_9__SCAN_IN, UWORD_REG_8__SCAN_IN, UWORD_REG_7__SCAN_IN,
         UWORD_REG_6__SCAN_IN, UWORD_REG_5__SCAN_IN, UWORD_REG_4__SCAN_IN,
         UWORD_REG_3__SCAN_IN, UWORD_REG_2__SCAN_IN, UWORD_REG_1__SCAN_IN,
         UWORD_REG_0__SCAN_IN, DATAO_REG_0__SCAN_IN, DATAO_REG_1__SCAN_IN,
         DATAO_REG_2__SCAN_IN, DATAO_REG_3__SCAN_IN, DATAO_REG_4__SCAN_IN,
         DATAO_REG_5__SCAN_IN, DATAO_REG_6__SCAN_IN, DATAO_REG_7__SCAN_IN,
         DATAO_REG_8__SCAN_IN, DATAO_REG_9__SCAN_IN, DATAO_REG_10__SCAN_IN,
         DATAO_REG_11__SCAN_IN, DATAO_REG_12__SCAN_IN, DATAO_REG_13__SCAN_IN,
         DATAO_REG_14__SCAN_IN, DATAO_REG_15__SCAN_IN, DATAO_REG_16__SCAN_IN,
         DATAO_REG_17__SCAN_IN, DATAO_REG_18__SCAN_IN, DATAO_REG_19__SCAN_IN,
         DATAO_REG_20__SCAN_IN, DATAO_REG_21__SCAN_IN, DATAO_REG_22__SCAN_IN,
         DATAO_REG_23__SCAN_IN, DATAO_REG_24__SCAN_IN, DATAO_REG_25__SCAN_IN,
         DATAO_REG_26__SCAN_IN, DATAO_REG_27__SCAN_IN, DATAO_REG_28__SCAN_IN,
         DATAO_REG_29__SCAN_IN, DATAO_REG_30__SCAN_IN, DATAO_REG_31__SCAN_IN,
         EAX_REG_0__SCAN_IN, EAX_REG_1__SCAN_IN, EAX_REG_2__SCAN_IN,
         EAX_REG_3__SCAN_IN, EAX_REG_4__SCAN_IN, EAX_REG_5__SCAN_IN,
         EAX_REG_6__SCAN_IN, EAX_REG_7__SCAN_IN, EAX_REG_8__SCAN_IN,
         EAX_REG_9__SCAN_IN, EAX_REG_10__SCAN_IN, EAX_REG_11__SCAN_IN,
         EAX_REG_12__SCAN_IN, EAX_REG_13__SCAN_IN, EAX_REG_14__SCAN_IN,
         EAX_REG_15__SCAN_IN, EAX_REG_16__SCAN_IN, EAX_REG_17__SCAN_IN,
         EAX_REG_18__SCAN_IN, EAX_REG_19__SCAN_IN, EAX_REG_20__SCAN_IN,
         EAX_REG_21__SCAN_IN, EAX_REG_22__SCAN_IN, EAX_REG_23__SCAN_IN,
         EAX_REG_24__SCAN_IN, EAX_REG_25__SCAN_IN, EAX_REG_26__SCAN_IN,
         EAX_REG_27__SCAN_IN, EAX_REG_28__SCAN_IN, EAX_REG_29__SCAN_IN,
         EAX_REG_30__SCAN_IN, EAX_REG_31__SCAN_IN, EBX_REG_0__SCAN_IN,
         EBX_REG_1__SCAN_IN, EBX_REG_2__SCAN_IN, EBX_REG_3__SCAN_IN,
         EBX_REG_4__SCAN_IN, EBX_REG_5__SCAN_IN, EBX_REG_6__SCAN_IN,
         EBX_REG_7__SCAN_IN, EBX_REG_8__SCAN_IN, EBX_REG_9__SCAN_IN,
         EBX_REG_10__SCAN_IN, EBX_REG_11__SCAN_IN, EBX_REG_12__SCAN_IN,
         EBX_REG_13__SCAN_IN, EBX_REG_14__SCAN_IN, EBX_REG_15__SCAN_IN,
         EBX_REG_16__SCAN_IN, EBX_REG_17__SCAN_IN, EBX_REG_18__SCAN_IN,
         EBX_REG_19__SCAN_IN, EBX_REG_20__SCAN_IN, EBX_REG_21__SCAN_IN,
         EBX_REG_22__SCAN_IN, EBX_REG_23__SCAN_IN, EBX_REG_24__SCAN_IN,
         EBX_REG_25__SCAN_IN, EBX_REG_26__SCAN_IN, EBX_REG_27__SCAN_IN,
         EBX_REG_28__SCAN_IN, EBX_REG_29__SCAN_IN, EBX_REG_30__SCAN_IN,
         EBX_REG_31__SCAN_IN, REIP_REG_0__SCAN_IN, REIP_REG_1__SCAN_IN,
         REIP_REG_2__SCAN_IN, REIP_REG_3__SCAN_IN, REIP_REG_4__SCAN_IN,
         REIP_REG_5__SCAN_IN, REIP_REG_6__SCAN_IN, REIP_REG_7__SCAN_IN,
         REIP_REG_8__SCAN_IN, REIP_REG_9__SCAN_IN, REIP_REG_10__SCAN_IN,
         REIP_REG_11__SCAN_IN, REIP_REG_12__SCAN_IN, REIP_REG_13__SCAN_IN,
         REIP_REG_14__SCAN_IN, REIP_REG_15__SCAN_IN, keyinput127, keyinput126,
         keyinput125, keyinput124, keyinput123, keyinput122, keyinput121,
         keyinput120, keyinput119, keyinput118, keyinput117, keyinput116,
         keyinput115, keyinput114, keyinput113, keyinput112, keyinput111,
         keyinput110, keyinput109, keyinput108, keyinput107, keyinput106,
         keyinput105, keyinput104, keyinput103, keyinput102, keyinput101,
         keyinput100, keyinput99, keyinput98, keyinput97, keyinput96,
         keyinput95, keyinput94, keyinput93, keyinput92, keyinput91,
         keyinput90, keyinput89, keyinput88, keyinput87, keyinput86,
         keyinput85, keyinput84, keyinput83, keyinput82, keyinput81,
         keyinput80, keyinput79, keyinput78, keyinput77, keyinput76,
         keyinput75, keyinput74, keyinput73, keyinput72, keyinput71,
         keyinput70, keyinput69, keyinput68, keyinput67, keyinput66,
         keyinput65, keyinput64, keyinput63, keyinput62, keyinput61,
         keyinput60, keyinput59, keyinput58, keyinput57, keyinput56,
         keyinput55, keyinput54, keyinput53, keyinput52, keyinput51,
         keyinput50, keyinput49, keyinput48, keyinput47, keyinput46,
         keyinput45, keyinput44, keyinput43, keyinput42, keyinput41,
         keyinput40, keyinput39, keyinput38, keyinput37, keyinput36,
         keyinput35, keyinput34, keyinput33, keyinput32, keyinput31,
         keyinput30, keyinput29, keyinput28, keyinput27, keyinput26,
         keyinput25, keyinput24, keyinput23, keyinput22, keyinput21,
         keyinput20, keyinput19, keyinput18, keyinput17, keyinput16,
         keyinput15, keyinput14, keyinput13, keyinput12, keyinput11,
         keyinput10, keyinput9, keyinput8, keyinput7, keyinput6, keyinput5,
         keyinput4, keyinput3, keyinput2, keyinput1, keyinput0;
  output U3445, U3446, U3447, U3448, U3213, U3212, U3211, U3210, U3209, U3208,
         U3207, U3206, U3205, U3204, U3203, U3202, U3201, U3200, U3199, U3198,
         U3197, U3196, U3195, U3194, U3193, U3192, U3191, U3190, U3189, U3188,
         U3187, U3186, U3185, U3184, U3183, U3182, U3181, U3451, U3452, U3180,
         U3179, U3178, U3177, U3176, U3175, U3174, U3173, U3172, U3171, U3170,
         U3169, U3168, U3167, U3166, U3165, U3164, U3163, U3162, U3161, U3160,
         U3159, U3158, U3157, U3156, U3155, U3154, U3153, U3152, U3151, U3453,
         U3150, U3149, U3148, U3147, U3146, U3145, U3144, U3143, U3142, U3141,
         U3140, U3139, U3138, U3137, U3136, U3135, U3134, U3133, U3132, U3131,
         U3130, U3129, U3128, U3127, U3126, U3125, U3124, U3123, U3122, U3121,
         U3120, U3119, U3118, U3117, U3116, U3115, U3114, U3113, U3112, U3111,
         U3110, U3109, U3108, U3107, U3106, U3105, U3104, U3103, U3102, U3101,
         U3100, U3099, U3098, U3097, U3096, U3095, U3094, U3093, U3092, U3091,
         U3090, U3089, U3088, U3087, U3086, U3085, U3084, U3083, U3082, U3081,
         U3080, U3079, U3078, U3077, U3076, U3075, U3074, U3073, U3072, U3071,
         U3070, U3069, U3068, U3067, U3066, U3065, U3064, U3063, U3062, U3061,
         U3060, U3059, U3058, U3057, U3056, U3055, U3054, U3053, U3052, U3051,
         U3050, U3049, U3048, U3047, U3046, U3045, U3044, U3043, U3042, U3041,
         U3040, U3039, U3038, U3037, U3036, U3035, U3034, U3033, U3032, U3031,
         U3030, U3029, U3028, U3027, U3026, U3025, U3024, U3023, U3022, U3021,
         U3020, U3455, U3456, U3459, U3460, U3461, U3019, U3462, U3463, U3464,
         U3465, U3018, U3017, U3016, U3015, U3014, U3013, U3012, U3011, U3010,
         U3009, U3008, U3007, U3006, U3005, U3004, U3003, U3002, U3001, U3000,
         U2999, U2998, U2997, U2996, U2995, U2994, U2993, U2992, U2991, U2990,
         U2989, U2988, U2987, U2986, U2985, U2984, U2983, U2982, U2981, U2980,
         U2979, U2978, U2977, U2976, U2975, U2974, U2973, U2972, U2971, U2970,
         U2969, U2968, U2967, U2966, U2965, U2964, U2963, U2962, U2961, U2960,
         U2959, U2958, U2957, U2956, U2955, U2954, U2953, U2952, U2951, U2950,
         U2949, U2948, U2947, U2946, U2945, U2944, U2943, U2942, U2941, U2940,
         U2939, U2938, U2937, U2936, U2935, U2934, U2933, U2932, U2931, U2930,
         U2929, U2928, U2927, U2926, U2925, U2924, U2923, U2922, U2921, U2920,
         U2919, U2918, U2917, U2916, U2915, U2914, U2913, U2912, U2911, U2910,
         U2909, U2908, U2907, U2906, U2905, U2904, U2903, U2902, U2901, U2900,
         U2899, U2898, U2897, U2896, U2895, U2894, U2893, U2892, U2891, U2890,
         U2889, U2888, U2887, U2886, U2885, U2884, U2883, U2882, U2881, U2880,
         U2879, U2878, U2877, U2876, U2875, U2874, U2873, U2872, U2871, U2870,
         U2869, U2868, U2867, U2866, U2865, U2864, U2863, U2862, U2861, U2860,
         U2859, U2858, U2857, U2856, U2855, U2854, U2853, U2852, U2851, U2850,
         U2849, U2848, U2847, U2846, U2845, U2844, U2843, U2842, U2841, U2840,
         U2839, U2838, U2837, U2836, U2835, U2834, U2833, U2832, U2831, U2830,
         U2829, U2828, U2827, U2826, U2825, U2824, U2823, U2822, U2821, U2820,
         U2819, U2818, U2817, U2816, U2815, U2814, U2813, U2812, U2811, U2810,
         U2809, U2808, U2807, U2806, U2805, U2804, U2803, U2802, U2801, U2800,
         U2799, U2798, U2797, U2796, U2795, U3468, U2794, U3469, U3470, U2793,
         U3471, U2792, U3472, U2791, U3473, U2790, U2789, U3474, U2788;
  wire   n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964;

  INV_X1 U3542 ( .A(n5200), .ZN(n5469) );
  OAI221_X1 U3543 ( .B1(n6706), .B2(keyinput70), .C1(n6705), .C2(keyinput95), 
        .A(n6704), .ZN(n6711) );
  NAND2_X1 U3544 ( .A1(n3822), .A2(n3821), .ZN(n4743) );
  CLKBUF_X2 U3545 ( .A(n3320), .Z(n3104) );
  NAND2_X1 U3546 ( .A1(n5906), .A2(n3393), .ZN(n3434) );
  NAND2_X1 U3547 ( .A1(n3481), .A2(n3479), .ZN(n3177) );
  AOI22_X1 U3548 ( .A1(n4823), .A2(keyinput63), .B1(n6740), .B2(keyinput97), 
        .ZN(n6739) );
  AOI22_X1 U3549 ( .A1(n6706), .A2(keyinput70), .B1(keyinput95), .B2(n6705), 
        .ZN(n6704) );
  NAND2_X1 U3550 ( .A1(n3409), .A2(n5888), .ZN(n4215) );
  INV_X1 U3551 ( .A(n4097), .ZN(n3409) );
  OAI221_X1 U3552 ( .B1(n4823), .B2(keyinput63), .C1(n6740), .C2(keyinput97), 
        .A(n6739), .ZN(n6741) );
  INV_X1 U3553 ( .A(n4122), .ZN(n4159) );
  AND2_X1 U3554 ( .A1(n3426), .A2(n3425), .ZN(n3481) );
  NAND2_X1 U3555 ( .A1(n4204), .A2(n4159), .ZN(n4468) );
  AND2_X1 U3556 ( .A1(n5687), .A2(n4821), .ZN(n5677) );
  INV_X1 U3557 ( .A(n4561), .ZN(n4178) );
  INV_X1 U3558 ( .A(n5164), .ZN(n5710) );
  INV_X1 U3559 ( .A(n5911), .ZN(n5768) );
  INV_X1 U3560 ( .A(n5631), .ZN(n5620) );
  INV_X1 U3561 ( .A(n5677), .ZN(n5691) );
  AND2_X1 U3562 ( .A1(n3341), .A2(n3338), .ZN(n3094) );
  XNOR2_X1 U3563 ( .A(n3523), .B(n3522), .ZN(n3600) );
  INV_X1 U3564 ( .A(n4428), .ZN(n3096) );
  INV_X8 U3565 ( .A(n3680), .ZN(n5245) );
  INV_X2 U3566 ( .A(n3680), .ZN(n5222) );
  INV_X4 U3567 ( .A(n3685), .ZN(n3680) );
  AOI21_X1 U3568 ( .B1(n3401), .B2(n3521), .A(n3400), .ZN(n3423) );
  AND2_X1 U3569 ( .A1(n3376), .A2(n4544), .ZN(n3427) );
  OR2_X1 U3570 ( .A1(n4220), .A2(n4108), .ZN(n4208) );
  INV_X1 U3571 ( .A(n4399), .ZN(n4453) );
  INV_X2 U3572 ( .A(n3397), .ZN(n3408) );
  INV_X1 U3573 ( .A(n3407), .ZN(n3095) );
  BUF_X2 U3574 ( .A(n4433), .Z(n4341) );
  CLKBUF_X2 U3575 ( .A(n3363), .Z(n4388) );
  BUF_X2 U3576 ( .A(n4364), .Z(n3110) );
  BUF_X2 U3577 ( .A(n4435), .Z(n3106) );
  CLKBUF_X2 U3578 ( .A(n3378), .Z(n3115) );
  INV_X2 U3579 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3777) );
  NOR2_X1 U3580 ( .A1(n4084), .A2(n3133), .ZN(n5207) );
  NAND2_X1 U3581 ( .A1(n3546), .A2(n3545), .ZN(n5863) );
  CLKBUF_X1 U3582 ( .A(n3390), .Z(n3719) );
  INV_X2 U3583 ( .A(n3435), .ZN(n3398) );
  AND2_X2 U3584 ( .A1(n3319), .A2(n3318), .ZN(n3435) );
  OR2_X1 U3585 ( .A1(n3373), .A2(n3372), .ZN(n5888) );
  AND2_X1 U3586 ( .A1(n3339), .A2(n3340), .ZN(n3129) );
  NAND4_X2 U3587 ( .A1(n3361), .A2(n3360), .A3(n3359), .A4(n3358), .ZN(n3407)
         );
  AND4_X1 U3588 ( .A1(n3317), .A2(n3316), .A3(n3315), .A4(n3314), .ZN(n3318)
         );
  AND4_X1 U3589 ( .A1(n3279), .A2(n3278), .A3(n3277), .A4(n3276), .ZN(n3295)
         );
  CLKBUF_X2 U3590 ( .A(n4359), .Z(n4427) );
  CLKBUF_X2 U3591 ( .A(n3465), .Z(n4434) );
  INV_X1 U3592 ( .A(STATE2_REG_1__SCAN_IN), .ZN(n6522) );
  AOI21_X1 U3593 ( .B1(n5195), .B2(n5768), .A(n5194), .ZN(n5196) );
  XNOR2_X1 U3594 ( .A(n5216), .B(n3699), .ZN(n5334) );
  OR2_X1 U3595 ( .A1(n5223), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n3167)
         );
  XNOR2_X1 U3596 ( .A(n3249), .B(n4455), .ZN(n5166) );
  OR2_X1 U3597 ( .A1(n5230), .A2(n5231), .ZN(n3172) );
  OR2_X1 U3598 ( .A1(n5230), .A2(n3168), .ZN(n5223) );
  OAI21_X1 U3599 ( .B1(n5124), .B2(n5117), .A(n5116), .ZN(n5416) );
  OAI22_X1 U3600 ( .A1(n5221), .A2(n5239), .B1(n5245), .B2(n5364), .ZN(n5230)
         );
  OR2_X1 U3601 ( .A1(n4084), .A2(n3134), .ZN(n5198) );
  AND2_X1 U3602 ( .A1(n5311), .A2(n5313), .ZN(n4084) );
  NAND2_X1 U3603 ( .A1(n5246), .A2(n3173), .ZN(n3695) );
  NAND2_X1 U3604 ( .A1(n5268), .A2(n3689), .ZN(n5246) );
  AND2_X1 U3605 ( .A1(n3155), .A2(n4882), .ZN(n3154) );
  NOR2_X1 U3606 ( .A1(n3165), .A2(n3164), .ZN(n3163) );
  INV_X1 U3607 ( .A(n4852), .ZN(n3918) );
  AOI21_X1 U3608 ( .B1(n3222), .B2(n3681), .A(n3225), .ZN(n3221) );
  NOR2_X1 U3609 ( .A1(n3226), .A2(n4836), .ZN(n3223) );
  NOR2_X1 U3610 ( .A1(n5258), .A2(n3220), .ZN(n3219) );
  NOR2_X1 U3611 ( .A1(n5245), .A2(n5534), .ZN(n3687) );
  OR2_X1 U3612 ( .A1(n5222), .A2(n4842), .ZN(n4837) );
  AOI21_X1 U3613 ( .B1(n3820), .B2(n3944), .A(n3819), .ZN(n4744) );
  OAI21_X1 U3614 ( .B1(n3801), .B2(n3851), .A(n3805), .ZN(n4704) );
  NAND2_X1 U3615 ( .A1(n3239), .A2(n3240), .ZN(n4649) );
  NAND3_X1 U3616 ( .A1(n3498), .A2(n3578), .A3(n3227), .ZN(n3580) );
  NAND2_X1 U3617 ( .A1(n5706), .A2(n5906), .ZN(n5162) );
  NAND2_X1 U3618 ( .A1(n6211), .A2(n6521), .ZN(n3546) );
  NAND2_X1 U3619 ( .A1(n3520), .A2(n3519), .ZN(n3523) );
  OR3_X1 U3620 ( .A1(n6626), .A2(n6516), .A3(n4457), .ZN(n5687) );
  AND2_X1 U3621 ( .A1(n3593), .A2(n3592), .ZN(n5868) );
  NAND2_X1 U3622 ( .A1(n3532), .A2(n3531), .ZN(n6020) );
  INV_X1 U3623 ( .A(n3098), .ZN(n4102) );
  NAND2_X1 U3624 ( .A1(n4159), .A2(n4561), .ZN(n4197) );
  NOR2_X1 U3625 ( .A1(n3744), .A2(n3399), .ZN(n3400) );
  OR2_X1 U3626 ( .A1(n3398), .A2(n6521), .ZN(n3533) );
  INV_X1 U3627 ( .A(n5888), .ZN(n4495) );
  AND4_X1 U3628 ( .A1(n3345), .A2(n3344), .A3(n3343), .A4(n3342), .ZN(n3361)
         );
  AND4_X1 U3629 ( .A1(n3357), .A2(n3356), .A3(n3355), .A4(n3354), .ZN(n3358)
         );
  AND4_X1 U3630 ( .A1(n3353), .A2(n3352), .A3(n3351), .A4(n3350), .ZN(n3359)
         );
  AND4_X1 U3631 ( .A1(n3332), .A2(n3331), .A3(n3330), .A4(n3329), .ZN(n3339)
         );
  AND4_X1 U3632 ( .A1(n3337), .A2(n3336), .A3(n3335), .A4(n3334), .ZN(n3338)
         );
  AND4_X1 U3633 ( .A1(n3328), .A2(n3327), .A3(n3326), .A4(n3325), .ZN(n3340)
         );
  AND4_X1 U3634 ( .A1(n3283), .A2(n3282), .A3(n3281), .A4(n3280), .ZN(n3294)
         );
  AND4_X1 U3635 ( .A1(n3324), .A2(n3323), .A3(n3322), .A4(n3321), .ZN(n3341)
         );
  AND4_X1 U3636 ( .A1(n3349), .A2(n3348), .A3(n3347), .A4(n3346), .ZN(n3360)
         );
  AND4_X1 U3637 ( .A1(n3287), .A2(n3286), .A3(n3285), .A4(n3284), .ZN(n3293)
         );
  NAND2_X2 U3638 ( .A1(n4071), .A2(n6419), .ZN(n5911) );
  AND2_X2 U3639 ( .A1(n4554), .A2(n3266), .ZN(n4433) );
  AND2_X2 U3640 ( .A1(n3258), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3266)
         );
  INV_X1 U3641 ( .A(STATE2_REG_3__SCAN_IN), .ZN(n6598) );
  NAND2_X1 U3642 ( .A1(n4496), .A2(n3252), .ZN(n3445) );
  AND2_X1 U3643 ( .A1(n3408), .A2(n3406), .ZN(n3097) );
  NOR2_X1 U3644 ( .A1(n3443), .A2(n3440), .ZN(n3098) );
  AND3_X1 U3645 ( .A1(n3396), .A2(n3429), .A3(n5906), .ZN(n3442) );
  AND2_X2 U3646 ( .A1(n3095), .A2(n3408), .ZN(n4812) );
  NAND2_X1 U3647 ( .A1(n3762), .A2(n3761), .ZN(n4608) );
  CLKBUF_X1 U3648 ( .A(n4651), .Z(n3119) );
  CLKBUF_X1 U3649 ( .A(n4649), .Z(n3099) );
  NAND2_X1 U3650 ( .A1(n3581), .A2(n3580), .ZN(n4688) );
  INV_X2 U3651 ( .A(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3258) );
  XNOR2_X1 U3652 ( .A(n3481), .B(n3480), .ZN(n6179) );
  NAND2_X2 U3653 ( .A1(n3580), .A2(n3498), .ZN(n3601) );
  AND4_X1 U3654 ( .A1(n3291), .A2(n3290), .A3(n3289), .A4(n3288), .ZN(n3292)
         );
  AND2_X2 U3655 ( .A1(n6659), .A2(n4549), .ZN(n4364) );
  NAND4_X1 U3656 ( .A1(n3361), .A2(n3360), .A3(n3359), .A4(n3358), .ZN(n3100)
         );
  NAND2_X1 U3657 ( .A1(n3407), .A2(n4495), .ZN(n4204) );
  OR2_X1 U3658 ( .A1(n3758), .A2(n3407), .ZN(n3440) );
  AND2_X1 U3659 ( .A1(n3268), .A2(n4550), .ZN(n3101) );
  AND2_X1 U3660 ( .A1(n3268), .A2(n4550), .ZN(n3320) );
  AND2_X2 U3661 ( .A1(n4693), .A2(n4704), .ZN(n4702) );
  AND2_X1 U3662 ( .A1(n6659), .A2(n4550), .ZN(n3362) );
  AND2_X1 U3663 ( .A1(n4550), .A2(n4660), .ZN(n3102) );
  AND2_X2 U3664 ( .A1(n4550), .A2(n4660), .ZN(n3103) );
  AND2_X2 U3665 ( .A1(n3268), .A2(n4549), .ZN(n3378) );
  AND2_X4 U3666 ( .A1(n3266), .A2(n3267), .ZN(n4359) );
  AND2_X1 U3667 ( .A1(n4554), .A2(n3266), .ZN(n3105) );
  AND2_X2 U3668 ( .A1(n3268), .A2(n3267), .ZN(n4435) );
  AND2_X4 U3669 ( .A1(n4554), .A2(n3268), .ZN(n3107) );
  AND2_X1 U3670 ( .A1(n3266), .A2(n4549), .ZN(n3117) );
  AND2_X1 U3671 ( .A1(n3266), .A2(n4549), .ZN(n3377) );
  AND2_X2 U3672 ( .A1(n3266), .A2(n4549), .ZN(n3116) );
  AND2_X2 U3673 ( .A1(n4549), .A2(n4660), .ZN(n3108) );
  AND2_X2 U3674 ( .A1(n4549), .A2(n4660), .ZN(n3109) );
  AND2_X2 U3675 ( .A1(n4549), .A2(n4660), .ZN(n4346) );
  AND2_X2 U3676 ( .A1(n3266), .A2(n4550), .ZN(n4428) );
  NAND2_X2 U3677 ( .A1(n3476), .A2(n3475), .ZN(n3498) );
  NAND2_X2 U3678 ( .A1(n4643), .A2(n4644), .ZN(n4642) );
  NAND2_X2 U3679 ( .A1(n3775), .A2(n3774), .ZN(n4643) );
  AND2_X1 U3680 ( .A1(n6659), .A2(n4554), .ZN(n3111) );
  AND2_X4 U3681 ( .A1(n6659), .A2(n4554), .ZN(n3112) );
  NAND2_X1 U3682 ( .A1(n3444), .A2(n3402), .ZN(n6475) );
  NAND2_X1 U3683 ( .A1(n3393), .A2(n3402), .ZN(n4604) );
  AND2_X1 U3684 ( .A1(n6659), .A2(n4550), .ZN(n3113) );
  AND2_X2 U3685 ( .A1(n6659), .A2(n4550), .ZN(n3114) );
  OR2_X2 U3686 ( .A1(n3389), .A2(n3388), .ZN(n4097) );
  NAND2_X4 U3687 ( .A1(n3129), .A2(n3094), .ZN(n3397) );
  NOR2_X1 U3688 ( .A1(n3434), .A2(n3435), .ZN(n3444) );
  NOR2_X4 U3689 ( .A1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3268) );
  NAND2_X2 U3690 ( .A1(n3410), .A2(n3390), .ZN(n4496) );
  INV_X2 U3691 ( .A(n3393), .ZN(n3410) );
  AND2_X2 U3692 ( .A1(n3404), .A2(n3403), .ZN(n4107) );
  NOR2_X2 U3693 ( .A1(n4952), .A2(n4966), .ZN(n4965) );
  NOR2_X2 U3694 ( .A1(n4983), .A2(n3235), .ZN(n5059) );
  NOR2_X2 U3695 ( .A1(n4070), .A2(n3241), .ZN(n5123) );
  XNOR2_X2 U3696 ( .A(n3905), .B(n3919), .ZN(n4910) );
  XNOR2_X2 U3697 ( .A(n5019), .B(n3250), .ZN(n5006) );
  AND2_X2 U3698 ( .A1(n5034), .A2(n3247), .ZN(n5019) );
  INV_X2 U3699 ( .A(n3096), .ZN(n3118) );
  XNOR2_X2 U3700 ( .A(n3601), .B(n3600), .ZN(n4687) );
  AND2_X1 U3701 ( .A1(n4554), .A2(n4660), .ZN(n3120) );
  AND2_X2 U3702 ( .A1(n4554), .A2(n4660), .ZN(n3121) );
  AND2_X4 U3703 ( .A1(n4554), .A2(n4660), .ZN(n3383) );
  AND2_X4 U3704 ( .A1(n4550), .A2(n4660), .ZN(n3333) );
  AND2_X4 U3705 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4550) );
  AND2_X4 U3706 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n4660) );
  NOR2_X4 U3707 ( .A1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4549) );
  NOR2_X1 U3708 ( .A1(n3122), .A2(n3135), .ZN(n3207) );
  INV_X1 U3709 ( .A(n3695), .ZN(n3208) );
  NAND2_X1 U3710 ( .A1(n3547), .A2(n3130), .ZN(n3622) );
  INV_X1 U3711 ( .A(n3619), .ZN(n3558) );
  OR2_X1 U3712 ( .A1(n3471), .A2(n3470), .ZN(n3671) );
  AND2_X1 U3713 ( .A1(n3100), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3714) );
  OR2_X1 U3714 ( .A1(n6475), .A2(n6521), .ZN(n4422) );
  INV_X1 U3715 ( .A(n3791), .ZN(n4448) );
  INV_X1 U3716 ( .A(n3683), .ZN(n3164) );
  NOR2_X1 U3717 ( .A1(n3157), .A2(n3158), .ZN(n3156) );
  INV_X1 U3718 ( .A(n3223), .ZN(n3157) );
  OR2_X1 U3719 ( .A1(n3491), .A2(n3490), .ZN(n3595) );
  INV_X1 U3720 ( .A(n3744), .ZN(n3707) );
  AOI21_X1 U3721 ( .B1(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B2(n6368), .A(n3743), 
        .ZN(n3739) );
  NAND2_X1 U3722 ( .A1(n3398), .A2(n3714), .ZN(n3744) );
  OR2_X1 U3723 ( .A1(n5222), .A2(n6828), .ZN(n5255) );
  NOR2_X1 U3724 ( .A1(n3174), .A2(n3136), .ZN(n3173) );
  INV_X1 U3725 ( .A(n3219), .ZN(n3174) );
  AND2_X1 U3726 ( .A1(n4113), .A2(n4112), .ZN(n4228) );
  OR2_X1 U3727 ( .A1(n4538), .A2(n4111), .ZN(n4112) );
  AND2_X1 U3728 ( .A1(n3707), .A2(n3706), .ZN(n3745) );
  NAND2_X1 U3729 ( .A1(n4197), .A2(n3180), .ZN(n3179) );
  AND2_X1 U3730 ( .A1(n5113), .A2(n3140), .ZN(n3188) );
  INV_X1 U3731 ( .A(n4467), .ZN(n3189) );
  NAND2_X1 U3732 ( .A1(n3238), .A2(n3253), .ZN(n3237) );
  INV_X1 U3733 ( .A(n5149), .ZN(n3238) );
  NAND2_X1 U3734 ( .A1(n3232), .A2(n4803), .ZN(n3231) );
  INV_X1 U3735 ( .A(n4774), .ZN(n3232) );
  INV_X1 U3736 ( .A(n3571), .ZN(n3569) );
  INV_X1 U3737 ( .A(n3763), .ZN(n3790) );
  NAND2_X1 U3738 ( .A1(n3202), .A2(n3201), .ZN(n3200) );
  INV_X1 U3739 ( .A(n4186), .ZN(n3202) );
  NOR2_X1 U3740 ( .A1(n3203), .A2(n5140), .ZN(n3201) );
  INV_X1 U3741 ( .A(n5135), .ZN(n3203) );
  INV_X1 U3742 ( .A(n4881), .ZN(n3158) );
  NAND2_X1 U3743 ( .A1(n4122), .A2(n4561), .ZN(n4199) );
  NOR2_X1 U3744 ( .A1(n3196), .A2(n3195), .ZN(n3194) );
  INV_X1 U3745 ( .A(n4705), .ZN(n3195) );
  NAND2_X1 U3746 ( .A1(n3198), .A2(n3197), .ZN(n3196) );
  INV_X1 U3747 ( .A(n4697), .ZN(n3197) );
  NAND2_X1 U3748 ( .A1(n3776), .A2(n3706), .ZN(n3152) );
  OAI211_X1 U3749 ( .C1(n3744), .C2(n3496), .A(n3495), .B(n3494), .ZN(n3589)
         );
  INV_X1 U3750 ( .A(n3671), .ZN(n3669) );
  INV_X1 U3751 ( .A(n3758), .ZN(n3374) );
  AND2_X1 U3752 ( .A1(n3504), .A2(n5980), .ZN(n5871) );
  OAI21_X1 U3753 ( .B1(n6631), .B2(n4680), .A(n6601), .ZN(n5866) );
  OR2_X1 U3754 ( .A1(n3407), .A2(n6521), .ZN(n3534) );
  AND2_X1 U3755 ( .A1(n5687), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4819) );
  INV_X1 U3756 ( .A(n4469), .ZN(n3186) );
  OR2_X1 U3757 ( .A1(n3188), .A2(n3187), .ZN(n3182) );
  NOR2_X1 U3758 ( .A1(n5023), .A2(n3191), .ZN(n3190) );
  INV_X1 U3759 ( .A(n4207), .ZN(n3191) );
  NOR2_X1 U3760 ( .A1(n5118), .A2(n5111), .ZN(n5113) );
  AND2_X1 U3761 ( .A1(n4162), .A2(n4161), .ZN(n4927) );
  INV_X1 U3762 ( .A(n3901), .ZN(n4452) );
  NOR2_X1 U3763 ( .A1(n4403), .A2(n5038), .ZN(n4404) );
  NAND2_X1 U3764 ( .A1(n4404), .A2(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n4459)
         );
  AND2_X1 U3765 ( .A1(n4338), .A2(n4337), .ZN(n5122) );
  OR2_X1 U3766 ( .A1(n5494), .A2(n3791), .ZN(n4337) );
  NAND2_X1 U3767 ( .A1(n5133), .A2(n3242), .ZN(n3241) );
  INV_X1 U3768 ( .A(n3243), .ZN(n3242) );
  NAND2_X1 U3769 ( .A1(n5233), .A2(n3251), .ZN(n4299) );
  AND2_X1 U3770 ( .A1(n4037), .A2(n4036), .ZN(n5061) );
  NOR2_X1 U3771 ( .A1(n3952), .A2(n3951), .ZN(n3982) );
  INV_X1 U3772 ( .A(n4863), .ZN(n3917) );
  NOR2_X1 U3773 ( .A1(n6716), .A2(n3823), .ZN(n3853) );
  OR2_X1 U3774 ( .A1(n3776), .A2(n3151), .ZN(n3144) );
  AOI21_X1 U3775 ( .B1(n3776), .B2(n3126), .A(n3146), .ZN(n3145) );
  NAND2_X1 U3776 ( .A1(n3608), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n5764)
         );
  NAND2_X1 U3777 ( .A1(n6513), .A2(n6518), .ZN(n4538) );
  INV_X1 U3778 ( .A(n4085), .ZN(n3213) );
  NAND2_X1 U3779 ( .A1(n5312), .A2(n3209), .ZN(n3211) );
  NOR2_X1 U3780 ( .A1(n3215), .A2(n4253), .ZN(n3209) );
  NAND2_X1 U3781 ( .A1(n5113), .A2(n4207), .ZN(n5022) );
  OR2_X1 U3782 ( .A1(n3133), .A2(n3216), .ZN(n3215) );
  NAND2_X1 U3783 ( .A1(n5205), .A2(n3217), .ZN(n3216) );
  INV_X1 U3784 ( .A(n5275), .ZN(n3217) );
  OR2_X1 U3785 ( .A1(n3128), .A2(n5120), .ZN(n5118) );
  NOR2_X1 U3786 ( .A1(n5215), .A2(n3170), .ZN(n3169) );
  INV_X1 U3787 ( .A(n3697), .ZN(n3170) );
  OR2_X1 U3788 ( .A1(n5231), .A2(n3171), .ZN(n3168) );
  INV_X1 U3789 ( .A(n5214), .ZN(n3171) );
  NAND2_X1 U3790 ( .A1(n5063), .A2(n4177), .ZN(n5345) );
  AND2_X1 U3791 ( .A1(n5255), .A2(n3693), .ZN(n3694) );
  NAND2_X1 U3792 ( .A1(n3218), .A2(n3162), .ZN(n3161) );
  NAND2_X1 U3793 ( .A1(n3684), .A2(n3163), .ZN(n3160) );
  INV_X1 U3794 ( .A(n3681), .ZN(n3226) );
  INV_X1 U3795 ( .A(n4837), .ZN(n3225) );
  NOR2_X1 U3796 ( .A1(n4736), .A2(n4735), .ZN(n4777) );
  NOR2_X1 U3797 ( .A1(n4076), .A2(STATE2_REG_2__SCAN_IN), .ZN(n5262) );
  CLKBUF_X1 U3798 ( .A(n4542), .Z(n4543) );
  INV_X1 U3799 ( .A(n5982), .ZN(n5979) );
  INV_X1 U3800 ( .A(n6177), .ZN(n6321) );
  AND2_X1 U3801 ( .A1(n4688), .A2(n5868), .ZN(n6108) );
  AND2_X1 U3802 ( .A1(n4687), .A2(n5863), .ZN(n6413) );
  AND2_X1 U3803 ( .A1(n6522), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3755) );
  NAND2_X1 U3804 ( .A1(n3534), .A2(n3533), .ZN(n3752) );
  AOI221_X1 U3805 ( .B1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .B2(n3739), .C1(
        n5548), .C2(n3739), .A(n3705), .ZN(n4095) );
  AND2_X1 U3806 ( .A1(n3746), .A2(n3744), .ZN(n3748) );
  OR2_X1 U3807 ( .A1(n5832), .A2(n6528), .ZN(n4457) );
  AND2_X1 U3808 ( .A1(n5164), .A2(n4979), .ZN(n5707) );
  AND2_X1 U3809 ( .A1(n5164), .A2(n4606), .ZN(n4956) );
  OR2_X1 U3810 ( .A1(n4538), .A2(n6496), .ZN(n5557) );
  INV_X1 U3811 ( .A(n5557), .ZN(n5774) );
  OR2_X1 U3812 ( .A1(n5307), .A2(n4247), .ZN(n5294) );
  INV_X1 U3813 ( .A(n3698), .ZN(n3699) );
  NAND2_X1 U3814 ( .A1(n3172), .A2(n3697), .ZN(n5216) );
  OR2_X1 U3815 ( .A1(n4228), .A2(n4210), .ZN(n5848) );
  OR2_X1 U3816 ( .A1(n4228), .A2(n4118), .ZN(n5824) );
  NAND2_X1 U3817 ( .A1(n6513), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6601) );
  AND2_X1 U3818 ( .A1(n6316), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3710)
         );
  NAND2_X1 U3819 ( .A1(n3408), .A2(n4088), .ZN(n3405) );
  OR2_X1 U3820 ( .A1(n3643), .A2(n3642), .ZN(n3651) );
  OR2_X1 U3821 ( .A1(n3458), .A2(n3457), .ZN(n3582) );
  OR2_X1 U3822 ( .A1(n3517), .A2(n3516), .ZN(n3573) );
  INV_X1 U3823 ( .A(n3533), .ZN(n3518) );
  INV_X1 U3824 ( .A(n3534), .ZN(n3521) );
  AND2_X1 U3825 ( .A1(n3421), .A2(n3423), .ZN(n3502) );
  AOI22_X1 U3826 ( .A1(n4359), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3465), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3270) );
  AND2_X1 U3827 ( .A1(n3741), .A2(n3740), .ZN(n3743) );
  INV_X1 U3828 ( .A(n4466), .ZN(n3187) );
  AND2_X1 U3829 ( .A1(n4979), .A2(STATE2_REG_2__SCAN_IN), .ZN(n3763) );
  NOR2_X1 U3830 ( .A1(n5020), .A2(n3248), .ZN(n3247) );
  INV_X1 U3831 ( .A(n5035), .ZN(n3248) );
  NAND2_X1 U3832 ( .A1(n3244), .A2(n3251), .ZN(n3243) );
  INV_X1 U3833 ( .A(n5139), .ZN(n3244) );
  NOR2_X1 U3834 ( .A1(n4955), .A2(n3234), .ZN(n3233) );
  INV_X1 U3835 ( .A(n4922), .ZN(n3234) );
  INV_X1 U3836 ( .A(n3764), .ZN(n4399) );
  OR2_X1 U3837 ( .A1(n3867), .A2(n5603), .ZN(n3882) );
  XNOR2_X1 U3838 ( .A(n3668), .B(n3661), .ZN(n3820) );
  NAND2_X1 U3839 ( .A1(n3127), .A2(n3147), .ZN(n3146) );
  NAND2_X1 U3840 ( .A1(n3150), .A2(n3148), .ZN(n3147) );
  NAND2_X1 U3841 ( .A1(n4608), .A2(n4607), .ZN(n3240) );
  INV_X1 U3842 ( .A(n3690), .ZN(n3220) );
  INV_X1 U3843 ( .A(n3686), .ZN(n3162) );
  NAND2_X1 U3844 ( .A1(n3179), .A2(n3178), .ZN(n4121) );
  NAND2_X1 U3845 ( .A1(n4159), .A2(EBX_REG_1__SCAN_IN), .ZN(n3178) );
  OR2_X1 U3846 ( .A1(n3544), .A2(n3543), .ZN(n3610) );
  AOI22_X1 U3847 ( .A1(n3111), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3113), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3296) );
  INV_X1 U3848 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6483) );
  INV_X1 U3849 ( .A(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n6489) );
  NAND2_X1 U3850 ( .A1(n3435), .A2(n3402), .ZN(n3758) );
  INV_X1 U3851 ( .A(n6480), .ZN(n4676) );
  OR2_X1 U3852 ( .A1(n6614), .A2(STATE2_REG_0__SCAN_IN), .ZN(n4076) );
  INV_X1 U3853 ( .A(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3951) );
  NOR2_X1 U3854 ( .A1(n3882), .A2(n4885), .ZN(n3897) );
  AND2_X1 U3855 ( .A1(n4206), .A2(n4205), .ZN(n4207) );
  INV_X1 U3856 ( .A(n3240), .ZN(n4610) );
  NOR2_X1 U3857 ( .A1(n3250), .A2(n3246), .ZN(n3245) );
  INV_X1 U3858 ( .A(n3247), .ZN(n3246) );
  INV_X1 U3859 ( .A(n5109), .ZN(n4383) );
  NAND2_X1 U3860 ( .A1(n4378), .A2(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n4403)
         );
  NAND2_X1 U3861 ( .A1(n4335), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4376)
         );
  AND2_X1 U3862 ( .A1(n4312), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4335)
         );
  NOR2_X1 U3863 ( .A1(n4293), .A2(n4292), .ZN(n4294) );
  INV_X1 U3864 ( .A(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n4292) );
  NAND2_X1 U3865 ( .A1(n4051), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4293)
         );
  INV_X1 U3866 ( .A(n4033), .ZN(n4034) );
  AND2_X1 U3867 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n4034), .ZN(n4051)
         );
  NAND2_X1 U3868 ( .A1(n5061), .A2(n3236), .ZN(n3235) );
  INV_X1 U3869 ( .A(n3237), .ZN(n3236) );
  NOR2_X1 U3870 ( .A1(n6705), .A2(n4000), .ZN(n4017) );
  AND2_X1 U3871 ( .A1(n3982), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3983)
         );
  NAND2_X1 U3872 ( .A1(n3983), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n4000)
         );
  NAND2_X1 U3873 ( .A1(n5246), .A2(n3690), .ZN(n5256) );
  AND2_X1 U3874 ( .A1(n3968), .A2(n3967), .ZN(n4966) );
  NOR2_X1 U3875 ( .A1(n6740), .A2(n3898), .ZN(n3932) );
  NOR2_X1 U3876 ( .A1(n3231), .A2(n3230), .ZN(n3229) );
  INV_X1 U3877 ( .A(n4853), .ZN(n3230) );
  NAND2_X1 U3878 ( .A1(n3853), .A2(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3867)
         );
  INV_X1 U3879 ( .A(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n5603) );
  AND2_X1 U3880 ( .A1(n3838), .A2(n3837), .ZN(n4774) );
  AND3_X1 U3881 ( .A1(n3836), .A2(n3835), .A3(n3834), .ZN(n3837) );
  NAND2_X1 U3882 ( .A1(n3815), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3823)
         );
  CLKBUF_X1 U3883 ( .A(n4710), .Z(n4711) );
  NOR2_X1 U3884 ( .A1(n3256), .A2(n3804), .ZN(n3805) );
  INV_X1 U3885 ( .A(n3803), .ZN(n3804) );
  AND2_X1 U3886 ( .A1(n3792), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3802)
         );
  AOI21_X1 U3887 ( .B1(n3800), .B2(n3944), .A(n3799), .ZN(n4695) );
  INV_X1 U3888 ( .A(n3798), .ZN(n3799) );
  CLKBUF_X1 U3889 ( .A(n4693), .Z(n4694) );
  NAND2_X1 U3890 ( .A1(PHYADDRPOINTER_REG_1__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3779) );
  INV_X1 U3891 ( .A(n5205), .ZN(n3214) );
  INV_X1 U3892 ( .A(n5127), .ZN(n3199) );
  AND2_X1 U3893 ( .A1(n4191), .A2(n4190), .ZN(n5135) );
  NOR2_X1 U3894 ( .A1(n5345), .A2(n3200), .ZN(n5137) );
  AND2_X1 U3895 ( .A1(n5346), .A2(n5335), .ZN(n5326) );
  NOR3_X1 U3896 ( .A1(n5345), .A2(n4186), .A3(n5140), .ZN(n5141) );
  AND2_X1 U3897 ( .A1(n4185), .A2(n4184), .ZN(n5051) );
  NAND2_X1 U3898 ( .A1(n5245), .A2(n5349), .ZN(n3697) );
  AND2_X1 U3899 ( .A1(n5078), .A2(n4172), .ZN(n5063) );
  OR2_X1 U3900 ( .A1(n5161), .A2(n4967), .ZN(n4987) );
  NOR2_X1 U3901 ( .A1(n4987), .A2(n4986), .ZN(n5078) );
  NOR2_X1 U3902 ( .A1(n4912), .A2(n4163), .ZN(n5159) );
  OR2_X1 U3903 ( .A1(n4228), .A2(n4225), .ZN(n5525) );
  NAND2_X1 U3904 ( .A1(n4847), .A2(n3204), .ZN(n4912) );
  AND2_X1 U3905 ( .A1(n3124), .A2(n3205), .ZN(n3204) );
  INV_X1 U3906 ( .A(n4878), .ZN(n3205) );
  OR2_X1 U3907 ( .A1(n4939), .A2(n4940), .ZN(n4942) );
  NAND2_X1 U3908 ( .A1(n4804), .A2(n3156), .ZN(n3153) );
  NAND2_X1 U3909 ( .A1(n4847), .A2(n3124), .ZN(n4877) );
  OR2_X1 U3910 ( .A1(n4804), .A2(n3678), .ZN(n3224) );
  AND2_X1 U3911 ( .A1(n4777), .A2(n4776), .ZN(n4847) );
  AND2_X1 U3912 ( .A1(n4903), .A2(n5859), .ZN(n5356) );
  AND2_X1 U3913 ( .A1(n4143), .A2(n4142), .ZN(n4735) );
  NAND2_X1 U3914 ( .A1(n3193), .A2(n3125), .ZN(n4736) );
  INV_X1 U3915 ( .A(n4715), .ZN(n3192) );
  NAND2_X1 U3916 ( .A1(n3193), .A2(n3194), .ZN(n4714) );
  NAND2_X1 U3917 ( .A1(n3193), .A2(n3198), .ZN(n4698) );
  NOR2_X1 U3918 ( .A1(n4826), .A2(n3196), .ZN(n4706) );
  NAND2_X1 U3919 ( .A1(n3618), .A2(n3617), .ZN(n4757) );
  NAND2_X1 U3920 ( .A1(n3152), .A2(n3614), .ZN(n3616) );
  OR2_X1 U3921 ( .A1(n4898), .A2(n5851), .ZN(n4241) );
  OR2_X1 U3922 ( .A1(n4228), .A2(n4653), .ZN(n4903) );
  AND2_X1 U3923 ( .A1(n5527), .A2(n6605), .ZN(n5851) );
  NAND2_X1 U3924 ( .A1(n5868), .A2(n3706), .ZN(n3598) );
  NOR2_X1 U3925 ( .A1(n4215), .A2(n3402), .ZN(n3404) );
  AOI21_X1 U3926 ( .B1(n3588), .B2(n3589), .A(n3497), .ZN(n3578) );
  INV_X1 U3927 ( .A(n4687), .ZN(n6149) );
  NAND2_X1 U3928 ( .A1(n3524), .A2(n3600), .ZN(n3609) );
  INV_X1 U3929 ( .A(n3525), .ZN(n3176) );
  NAND2_X1 U3930 ( .A1(n4687), .A2(n5398), .ZN(n6110) );
  NAND2_X1 U3931 ( .A1(n3776), .A2(n6149), .ZN(n6248) );
  INV_X1 U3932 ( .A(n6108), .ZN(n6244) );
  AND2_X1 U3933 ( .A1(n5867), .A2(n5866), .ZN(n5907) );
  NOR2_X1 U3934 ( .A1(n6522), .A2(n6511), .ZN(n4680) );
  NAND2_X1 U3935 ( .A1(n4525), .A2(n4505), .ZN(n6626) );
  NOR2_X1 U3936 ( .A1(STATE2_REG_1__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6631) );
  NOR2_X1 U3937 ( .A1(n5591), .A2(n4977), .ZN(n5579) );
  INV_X1 U3938 ( .A(PHYADDRPOINTER_REG_13__SCAN_IN), .ZN(n6740) );
  INV_X1 U3939 ( .A(n5693), .ZN(n5665) );
  NAND2_X1 U3940 ( .A1(n4819), .A2(n4475), .ZN(n5653) );
  INV_X1 U3941 ( .A(n5640), .ZN(n5651) );
  INV_X1 U3942 ( .A(n5674), .ZN(n5692) );
  AND2_X1 U3943 ( .A1(n4819), .A2(n4817), .ZN(n5693) );
  AND2_X1 U3944 ( .A1(n5620), .A2(n4813), .ZN(n5698) );
  NAND3_X1 U3945 ( .A1(n3184), .A2(n3183), .A3(n3181), .ZN(n5279) );
  NAND2_X1 U3946 ( .A1(n5113), .A2(n3190), .ZN(n5024) );
  NAND2_X1 U3947 ( .A1(n4500), .A2(n6518), .ZN(n5145) );
  NAND2_X1 U3948 ( .A1(n4556), .A2(n4499), .ZN(n4500) );
  INV_X1 U3949 ( .A(n5906), .ZN(n5165) );
  NAND2_X1 U3950 ( .A1(n4603), .A2(n4641), .ZN(n5164) );
  OAI21_X1 U3951 ( .B1(n4602), .B2(n4601), .A(n6518), .ZN(n4603) );
  INV_X1 U3952 ( .A(n4956), .ZN(n4951) );
  INV_X1 U3953 ( .A(n5714), .ZN(n5722) );
  AND2_X1 U3954 ( .A1(n4540), .A2(n4562), .ZN(n5739) );
  INV_X1 U3955 ( .A(n5749), .ZN(n5743) );
  OR3_X1 U3956 ( .A1(n4525), .A2(n3408), .A3(READY_N), .ZN(n4641) );
  OAI21_X1 U3957 ( .B1(n3428), .B2(n6628), .A(n4524), .ZN(n5753) );
  INV_X1 U3958 ( .A(n4641), .ZN(n5759) );
  XNOR2_X1 U3959 ( .A(n4461), .B(n4460), .ZN(n4820) );
  AOI21_X1 U3960 ( .B1(n5126), .B2(n5125), .A(n5124), .ZN(n5491) );
  INV_X1 U3961 ( .A(PHYADDRPOINTER_REG_18__SCAN_IN), .ZN(n6705) );
  INV_X1 U3962 ( .A(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n4885) );
  AND2_X1 U3963 ( .A1(n3149), .A2(n5765), .ZN(n4749) );
  OR2_X1 U3964 ( .A1(n5777), .A2(n4075), .ZN(n5773) );
  INV_X1 U3965 ( .A(n5777), .ZN(n5248) );
  AND2_X1 U3966 ( .A1(n4898), .A2(n4903), .ZN(n5852) );
  OAI21_X1 U3967 ( .B1(n5312), .B2(n3212), .A(n3211), .ZN(n3210) );
  NAND2_X1 U3968 ( .A1(n3213), .A2(n3143), .ZN(n3212) );
  NOR2_X1 U3969 ( .A1(n4084), .A2(n3215), .ZN(n4488) );
  NAND2_X1 U3970 ( .A1(n3167), .A2(n3166), .ZN(n5217) );
  NAND2_X1 U3971 ( .A1(n3172), .A2(n3169), .ZN(n3166) );
  AND2_X1 U3972 ( .A1(n5372), .A2(n5360), .ZN(n5346) );
  NOR2_X1 U3973 ( .A1(n4244), .A2(n5503), .ZN(n5372) );
  NAND2_X1 U3974 ( .A1(n3695), .A2(n3694), .ZN(n5370) );
  NAND2_X1 U3975 ( .A1(n4804), .A2(n3223), .ZN(n3159) );
  INV_X1 U3976 ( .A(n5262), .ZN(n5811) );
  INV_X1 U3977 ( .A(n5811), .ZN(n5832) );
  INV_X1 U3978 ( .A(n4903), .ZN(n5835) );
  INV_X1 U3979 ( .A(n5824), .ZN(n5854) );
  INV_X1 U3980 ( .A(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n6316) );
  INV_X1 U3981 ( .A(n6419), .ZN(n6410) );
  NOR2_X2 U3982 ( .A1(STATE2_REG_3__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6419) );
  OAI21_X1 U3983 ( .B1(n4679), .B2(n6596), .A(n6148), .ZN(n5860) );
  NAND2_X1 U3984 ( .A1(n6598), .A2(n6522), .ZN(n6614) );
  OAI21_X1 U3985 ( .B1(n5908), .B2(n6598), .A(n5873), .ZN(n5913) );
  OAI21_X1 U3986 ( .B1(n5972), .B2(n5957), .A(n6214), .ZN(n5975) );
  OAI211_X1 U3987 ( .C1(n6039), .C2(n6598), .A(n6024), .B(n6023), .ZN(n6042)
         );
  OAI211_X1 U3988 ( .C1(n6170), .C2(n6598), .A(n6290), .B(n6155), .ZN(n6173)
         );
  INV_X1 U3989 ( .A(n6357), .ZN(n6335) );
  NAND2_X1 U3990 ( .A1(n6413), .A2(n6321), .ZN(n6405) );
  INV_X1 U3991 ( .A(n6323), .ZN(n6411) );
  INV_X1 U3992 ( .A(n6333), .ZN(n6429) );
  INV_X1 U3993 ( .A(n6339), .ZN(n6435) );
  INV_X1 U3994 ( .A(n6347), .ZN(n6449) );
  INV_X1 U3995 ( .A(n6351), .ZN(n6456) );
  AND2_X1 U3996 ( .A1(n6413), .A2(n6370), .ZN(n6468) );
  AND2_X1 U3997 ( .A1(n3755), .A2(STATE2_REG_0__SCAN_IN), .ZN(n6518) );
  INV_X2 U3998 ( .A(STATE2_REG_0__SCAN_IN), .ZN(n6521) );
  AND2_X1 U3999 ( .A1(n3754), .A2(n3753), .ZN(n6513) );
  OAI21_X1 U4000 ( .B1(n5178), .B2(n5911), .A(n4078), .ZN(n4079) );
  AND2_X1 U4001 ( .A1(n4251), .A2(n4250), .ZN(n4252) );
  NAND2_X1 U4002 ( .A1(n3668), .A2(n3670), .ZN(n3685) );
  INV_X1 U4003 ( .A(n3407), .ZN(n3438) );
  AND2_X1 U4004 ( .A1(n3123), .A2(n3142), .ZN(n3122) );
  AND2_X1 U4005 ( .A1(n3694), .A2(n6854), .ZN(n3123) );
  INV_X1 U4006 ( .A(n4084), .ZN(n5312) );
  AND2_X1 U4007 ( .A1(n4152), .A2(n3139), .ZN(n3124) );
  AND2_X1 U4008 ( .A1(n3194), .A2(n3192), .ZN(n3125) );
  AND2_X1 U4009 ( .A1(n3706), .A2(n3615), .ZN(n3126) );
  OR2_X1 U4010 ( .A1(n3614), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3127)
         );
  OR3_X1 U4011 ( .A1(n5345), .A2(n3200), .A3(n3199), .ZN(n3128) );
  NAND2_X1 U4012 ( .A1(n5246), .A2(n3219), .ZN(n5244) );
  NOR2_X1 U4013 ( .A1(n4070), .A2(n3243), .ZN(n5132) );
  NAND2_X1 U4014 ( .A1(n4942), .A2(n3686), .ZN(n4958) );
  OAI22_X1 U4015 ( .A1(n3208), .A2(n3207), .B1(n3680), .B2(n4083), .ZN(n5311)
         );
  NAND2_X1 U4016 ( .A1(n3570), .A2(n3569), .ZN(n3646) );
  NAND2_X1 U4017 ( .A1(n3646), .A2(n3572), .ZN(n3801) );
  AND2_X1 U4018 ( .A1(n5863), .A2(n3558), .ZN(n3130) );
  AND2_X1 U4019 ( .A1(n3695), .A2(n3123), .ZN(n5369) );
  NAND2_X1 U4020 ( .A1(n3645), .A2(n3644), .ZN(n3668) );
  OR2_X1 U4021 ( .A1(n5868), .A2(n3434), .ZN(n3131) );
  NAND2_X1 U4022 ( .A1(n3498), .A2(n3227), .ZN(n3132) );
  NOR2_X1 U4023 ( .A1(n4983), .A2(n3237), .ZN(n5060) );
  AOI21_X1 U4024 ( .B1(n4940), .B2(n3686), .A(n3687), .ZN(n3218) );
  NAND2_X1 U4025 ( .A1(n5072), .A2(n3253), .ZN(n5071) );
  NAND2_X1 U4026 ( .A1(n3507), .A2(n3506), .ZN(n3526) );
  AND2_X1 U4027 ( .A1(n5245), .A2(n4192), .ZN(n3133) );
  AND2_X1 U4028 ( .A1(n3397), .A2(n3407), .ZN(n4561) );
  AND2_X1 U4029 ( .A1(n4107), .A2(n3407), .ZN(n4456) );
  INV_X1 U4030 ( .A(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3711) );
  NAND2_X1 U4031 ( .A1(n4923), .A2(n4922), .ZN(n4921) );
  NOR2_X1 U4032 ( .A1(n4743), .A2(n4774), .ZN(n4773) );
  NOR2_X1 U4033 ( .A1(n4743), .A2(n3231), .ZN(n4801) );
  INV_X1 U4034 ( .A(n4494), .ZN(n3250) );
  NAND2_X1 U4035 ( .A1(n3228), .A2(n3229), .ZN(n4852) );
  NAND2_X1 U4036 ( .A1(n3224), .A2(n3681), .ZN(n4835) );
  AND2_X1 U4037 ( .A1(n3397), .A2(n3402), .ZN(n3706) );
  INV_X1 U4038 ( .A(n3706), .ZN(n3148) );
  NAND2_X1 U4039 ( .A1(n3684), .A2(n3683), .ZN(n4939) );
  OR2_X1 U4040 ( .A1(n3133), .A2(n3214), .ZN(n3134) );
  AND2_X1 U4041 ( .A1(n3694), .A2(n5222), .ZN(n3135) );
  AND2_X1 U4042 ( .A1(n5245), .A2(n4244), .ZN(n3136) );
  OR2_X1 U4043 ( .A1(n5345), .A2(n4186), .ZN(n3137) );
  INV_X1 U4044 ( .A(n3151), .ZN(n3150) );
  NAND2_X1 U4045 ( .A1(n3614), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3151)
         );
  INV_X1 U4046 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3206) );
  AND2_X1 U4047 ( .A1(n4847), .A2(n4152), .ZN(n3138) );
  INV_X1 U4048 ( .A(n4826), .ZN(n3193) );
  NAND3_X1 U4049 ( .A1(n4154), .A2(n4180), .A3(n4153), .ZN(n3139) );
  AND2_X1 U4050 ( .A1(n3190), .A2(n3189), .ZN(n3140) );
  NOR2_X1 U4051 ( .A1(n3187), .A2(n4469), .ZN(n3141) );
  AND3_X1 U4052 ( .A1(n4082), .A2(n5336), .A3(n5364), .ZN(n3142) );
  NOR4_X1 U4053 ( .A1(INSTADDRPOINTER_REG_28__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_29__SCAN_IN), .A3(INSTADDRPOINTER_REG_26__SCAN_IN), 
        .A4(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n3143) );
  INV_X1 U4054 ( .A(EBX_REG_1__SCAN_IN), .ZN(n3180) );
  NAND3_X1 U4055 ( .A1(n3149), .A2(n5765), .A3(n4750), .ZN(n3618) );
  NAND2_X1 U4056 ( .A1(n3145), .A2(n3144), .ZN(n4750) );
  NAND2_X1 U4057 ( .A1(n5767), .A2(n5764), .ZN(n3149) );
  AND2_X1 U4058 ( .A1(n4786), .A2(n3599), .ZN(n5767) );
  OR2_X1 U4059 ( .A1(n3221), .A2(n3158), .ZN(n3155) );
  NAND2_X1 U4060 ( .A1(n3154), .A2(n3153), .ZN(n4891) );
  NAND2_X1 U4061 ( .A1(n3159), .A2(n3221), .ZN(n4880) );
  NAND3_X1 U4062 ( .A1(n3161), .A2(n3160), .A3(n3688), .ZN(n5268) );
  INV_X1 U4063 ( .A(n3218), .ZN(n3165) );
  INV_X1 U4064 ( .A(n3172), .ZN(n5229) );
  NAND2_X1 U4065 ( .A1(n3418), .A2(n3177), .ZN(n3175) );
  NAND2_X1 U4066 ( .A1(n3175), .A2(n3499), .ZN(n3525) );
  NAND2_X1 U4067 ( .A1(n3176), .A2(n3526), .ZN(n4674) );
  INV_X1 U4068 ( .A(n3177), .ZN(n3500) );
  NAND2_X1 U4069 ( .A1(n3418), .A2(n3499), .ZN(n3501) );
  NAND4_X1 U4070 ( .A1(n3409), .A2(n3719), .A3(n4495), .A4(n4812), .ZN(n4220)
         );
  NAND2_X1 U4071 ( .A1(n5888), .A2(n3397), .ZN(n4119) );
  NAND2_X1 U4072 ( .A1(n3182), .A2(n4469), .ZN(n3181) );
  OR2_X1 U4073 ( .A1(n4465), .A2(n3186), .ZN(n3183) );
  NAND3_X1 U4074 ( .A1(n4465), .A2(n3185), .A3(n3141), .ZN(n3184) );
  INV_X1 U4075 ( .A(n3188), .ZN(n3185) );
  INV_X1 U4076 ( .A(n4646), .ZN(n3198) );
  AND2_X4 U4077 ( .A1(n3206), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n4554)
         );
  NOR2_X1 U4078 ( .A1(n5312), .A2(n4085), .ZN(n4487) );
  INV_X1 U4079 ( .A(n3210), .ZN(n4489) );
  NAND2_X1 U4080 ( .A1(n3621), .A2(n3622), .ZN(n3787) );
  NAND2_X1 U4081 ( .A1(n3547), .A2(n5863), .ZN(n3620) );
  NOR2_X1 U4082 ( .A1(n4836), .A2(n3679), .ZN(n3222) );
  NAND2_X1 U4083 ( .A1(n3478), .A2(n3477), .ZN(n3227) );
  NAND3_X1 U4084 ( .A1(n3646), .A2(n3572), .A3(n3706), .ZN(n3577) );
  INV_X1 U4085 ( .A(n4743), .ZN(n3228) );
  NAND2_X1 U4086 ( .A1(n4923), .A2(n3233), .ZN(n4952) );
  NAND2_X2 U4087 ( .A1(n3921), .A2(n3920), .ZN(n4923) );
  NAND2_X1 U4088 ( .A1(n3770), .A2(n3901), .ZN(n3773) );
  INV_X1 U4089 ( .A(n3773), .ZN(n3239) );
  NAND2_X1 U4090 ( .A1(n4649), .A2(n4648), .ZN(n3775) );
  NAND2_X1 U4091 ( .A1(n5034), .A2(n5035), .ZN(n5018) );
  NAND2_X1 U4092 ( .A1(n5034), .A2(n3245), .ZN(n3249) );
  OR2_X1 U4093 ( .A1(n4610), .A2(n4609), .ZN(n4789) );
  NAND2_X1 U4094 ( .A1(n3103), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3308)
         );
  NOR4_X2 U4095 ( .A1(n5207), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_28__SCAN_IN), .A4(n5204), .ZN(n5181) );
  NAND2_X1 U4096 ( .A1(n5166), .A2(n5631), .ZN(n4486) );
  AND2_X1 U4097 ( .A1(n4069), .A2(n4068), .ZN(n3251) );
  NAND2_X1 U4098 ( .A1(n5164), .A2(n4605), .ZN(n5468) );
  AND2_X1 U4099 ( .A1(n5906), .A2(n3435), .ZN(n3252) );
  AND2_X1 U4100 ( .A1(n4002), .A2(n4001), .ZN(n3253) );
  AND2_X2 U4101 ( .A1(n5557), .A2(n4072), .ZN(n5777) );
  OR2_X1 U4102 ( .A1(n3424), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n3425)
         );
  INV_X1 U4103 ( .A(PHYADDRPOINTER_REG_6__SCAN_IN), .ZN(n3813) );
  OAI21_X1 U4104 ( .B1(n3695), .B2(n6854), .A(n5245), .ZN(n3691) );
  AND2_X1 U4105 ( .A1(n4266), .A2(n4265), .ZN(n3254) );
  NAND2_X1 U4106 ( .A1(n5706), .A2(n5165), .ZN(n5156) );
  INV_X1 U4107 ( .A(n5156), .ZN(n4502) );
  OR2_X1 U4108 ( .A1(n3416), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3255)
         );
  NAND2_X1 U4109 ( .A1(n6511), .A2(n6286), .ZN(n3791) );
  AND2_X1 U4110 ( .A1(n4453), .A2(EAX_REG_5__SCAN_IN), .ZN(n3256) );
  INV_X1 U4111 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .ZN(n5548) );
  INV_X1 U4112 ( .A(n4812), .ZN(n3717) );
  AND2_X1 U4113 ( .A1(n5245), .A2(n6828), .ZN(n5258) );
  NOR2_X1 U4114 ( .A1(n4863), .A2(n4876), .ZN(n3257) );
  NAND2_X1 U4115 ( .A1(n6521), .A2(n5866), .ZN(n6148) );
  INV_X1 U4116 ( .A(n3477), .ZN(n3475) );
  AOI21_X1 U4117 ( .B1(n3419), .B2(n6363), .A(n3413), .ZN(n3415) );
  OR2_X1 U4118 ( .A1(n3568), .A2(n3567), .ZN(n3648) );
  NAND2_X1 U4119 ( .A1(n3363), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3307) );
  OR2_X1 U4120 ( .A1(n3557), .A2(n3556), .ZN(n3624) );
  INV_X1 U4121 ( .A(n3440), .ZN(n3406) );
  AOI22_X1 U4122 ( .A1(n4364), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3320), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n3314) );
  NOR2_X1 U4123 ( .A1(n3148), .A2(n3669), .ZN(n3670) );
  INV_X1 U4124 ( .A(n3502), .ZN(n3527) );
  AND2_X1 U4125 ( .A1(n3441), .A2(n4213), .ZN(n3447) );
  AND2_X1 U4126 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n4377), .ZN(n4378)
         );
  NAND2_X1 U4127 ( .A1(n3897), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3898)
         );
  AND2_X1 U4128 ( .A1(PHYADDRPOINTER_REG_3__SCAN_IN), .A2(n3778), .ZN(n3792)
         );
  OR2_X1 U4129 ( .A1(n5405), .A2(n3791), .ZN(n4381) );
  AND2_X1 U4130 ( .A1(n4846), .A2(n4845), .ZN(n4152) );
  NAND2_X1 U4131 ( .A1(n4128), .A2(n4178), .ZN(n4180) );
  OR2_X1 U4132 ( .A1(n4459), .A2(n4458), .ZN(n4461) );
  AND2_X1 U4133 ( .A1(n4294), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4312)
         );
  NOR2_X1 U4134 ( .A1(n5906), .A2(n6511), .ZN(n3764) );
  NOR2_X1 U4135 ( .A1(n3814), .A2(n3813), .ZN(n3815) );
  INV_X1 U4136 ( .A(n3787), .ZN(n3800) );
  NOR2_X2 U4137 ( .A1(n3410), .A2(n6511), .ZN(n3944) );
  INV_X1 U4138 ( .A(n4197), .ZN(n4202) );
  OR2_X1 U4139 ( .A1(n6513), .A2(n4653), .ZN(n4556) );
  AND2_X1 U4140 ( .A1(n4521), .A2(n3098), .ZN(n4510) );
  NAND2_X1 U4141 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n3932), .ZN(n3952)
         );
  INV_X1 U4142 ( .A(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n6716) );
  AND2_X1 U4143 ( .A1(n4820), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4821) );
  AND3_X1 U4144 ( .A1(n4170), .A2(n4180), .A3(n4169), .ZN(n4986) );
  INV_X1 U4145 ( .A(n5587), .ZN(n5271) );
  NAND2_X1 U4146 ( .A1(n3802), .A2(PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3814)
         );
  OR2_X1 U4147 ( .A1(n3608), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n5765)
         );
  AND3_X1 U4148 ( .A1(n4237), .A2(n5358), .A3(n4236), .ZN(n5350) );
  AND2_X1 U4149 ( .A1(n5527), .A2(n5525), .ZN(n4898) );
  OR2_X1 U4150 ( .A1(n4228), .A2(n6478), .ZN(n5527) );
  INV_X1 U4151 ( .A(n6148), .ZN(n5956) );
  OR2_X1 U4152 ( .A1(n3776), .A2(n4687), .ZN(n5982) );
  INV_X1 U4153 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6368) );
  INV_X1 U4154 ( .A(n5868), .ZN(n5952) );
  AOI21_X1 U4155 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6316), .A(n6148), .ZN(
        n6418) );
  INV_X1 U4156 ( .A(n4456), .ZN(n4515) );
  NOR2_X1 U4157 ( .A1(n5073), .A2(n4481), .ZN(n5048) );
  NOR2_X1 U4158 ( .A1(n5602), .A2(n4914), .ZN(n4925) );
  NOR2_X1 U4159 ( .A1(n5653), .A2(n4480), .ZN(n5608) );
  AND2_X1 U4160 ( .A1(n5687), .A2(n4462), .ZN(n5631) );
  AND2_X1 U4161 ( .A1(n5687), .A2(STATE2_REG_3__SCAN_IN), .ZN(n5674) );
  AND2_X1 U4162 ( .A1(n4819), .A2(n4471), .ZN(n5690) );
  INV_X1 U4163 ( .A(n5162), .ZN(n5703) );
  INV_X1 U4164 ( .A(n5468), .ZN(n5708) );
  INV_X1 U4165 ( .A(n5746), .ZN(n5738) );
  INV_X1 U4166 ( .A(n4612), .ZN(n5760) );
  NAND2_X1 U4167 ( .A1(n4017), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4033)
         );
  INV_X1 U4168 ( .A(n5773), .ZN(n5250) );
  OR2_X1 U4169 ( .A1(n4116), .A2(n3758), .ZN(n6496) );
  INV_X1 U4170 ( .A(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4086) );
  OR2_X1 U4171 ( .A1(n5331), .A2(n4239), .ZN(n5318) );
  INV_X1 U4172 ( .A(n4241), .ZN(n5841) );
  INV_X1 U4173 ( .A(n5848), .ZN(n5834) );
  OR3_X1 U4174 ( .A1(n4570), .A2(n4602), .A3(n4569), .ZN(n6480) );
  INV_X1 U4175 ( .A(n5945), .ZN(n5912) );
  INV_X1 U4176 ( .A(n6011), .ZN(n5974) );
  INV_X1 U4177 ( .A(n6080), .ZN(n6041) );
  INV_X1 U4178 ( .A(n6144), .ZN(n6103) );
  INV_X1 U4179 ( .A(n6954), .ZN(n6172) );
  OR2_X1 U4180 ( .A1(n4688), .A2(n5868), .ZN(n6150) );
  OAI21_X1 U4181 ( .B1(n6217), .B2(n6249), .A(n6216), .ZN(n6240) );
  OR2_X1 U4182 ( .A1(n4688), .A2(n5952), .ZN(n6177) );
  OAI211_X1 U4183 ( .C1(n6293), .C2(n6292), .A(n6291), .B(n6290), .ZN(n6310)
         );
  INV_X1 U4184 ( .A(n6150), .ZN(n6285) );
  OAI211_X1 U4185 ( .C1(n6399), .C2(n6598), .A(n6375), .B(n6374), .ZN(n6402)
         );
  INV_X1 U4186 ( .A(n6951), .ZN(n6425) );
  INV_X1 U4187 ( .A(n6343), .ZN(n6442) );
  INV_X1 U4188 ( .A(n6356), .ZN(n6463) );
  INV_X2 U4189 ( .A(STATE2_REG_2__SCAN_IN), .ZN(n6511) );
  INV_X1 U4190 ( .A(n6589), .ZN(n6574) );
  INV_X1 U4191 ( .A(STATE_REG_0__SCAN_IN), .ZN(n6541) );
  OR2_X1 U4192 ( .A1(n4538), .A2(n4515), .ZN(n4525) );
  INV_X1 U4193 ( .A(STATEBS16_REG_SCAN_IN), .ZN(n6286) );
  NOR2_X1 U4194 ( .A1(n4484), .A2(n4483), .ZN(n4485) );
  INV_X1 U4195 ( .A(n5690), .ZN(n5681) );
  AOI21_X1 U4196 ( .B1(n4998), .B2(n4502), .A(n4501), .ZN(n4503) );
  INV_X2 U4197 ( .A(n5145), .ZN(n5706) );
  INV_X1 U4198 ( .A(n4946), .ZN(n4949) );
  INV_X1 U4199 ( .A(n5739), .ZN(n5748) );
  OR2_X1 U4200 ( .A1(n5739), .A2(n5738), .ZN(n5749) );
  INV_X1 U4201 ( .A(n5753), .ZN(n4612) );
  OR2_X1 U4202 ( .A1(n4538), .A2(n6507), .ZN(n5762) );
  INV_X1 U4203 ( .A(n4079), .ZN(n4080) );
  NAND2_X1 U4204 ( .A1(n5334), .A2(n5854), .ZN(n5342) );
  INV_X1 U4205 ( .A(n5533), .ZN(n5786) );
  AND2_X1 U4206 ( .A1(n4586), .A2(n4587), .ZN(n5859) );
  INV_X1 U4207 ( .A(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .ZN(n5861) );
  NAND2_X1 U4208 ( .A1(n5979), .A2(n6285), .ZN(n5945) );
  NAND2_X1 U4209 ( .A1(n5979), .A2(n6321), .ZN(n5978) );
  NAND2_X1 U4210 ( .A1(n5979), .A2(n6370), .ZN(n6011) );
  NAND2_X1 U4211 ( .A1(n5979), .A2(n6108), .ZN(n6045) );
  OR2_X1 U4212 ( .A1(n6150), .A2(n6110), .ZN(n6080) );
  OR2_X1 U4213 ( .A1(n6177), .A2(n6110), .ZN(n6107) );
  OR2_X1 U4214 ( .A1(n6110), .A2(n6207), .ZN(n6144) );
  OR2_X1 U4215 ( .A1(n6110), .A2(n6244), .ZN(n6176) );
  OR2_X1 U4216 ( .A1(n6248), .A2(n6150), .ZN(n6954) );
  OR2_X1 U4217 ( .A1(n6248), .A2(n6177), .ZN(n6961) );
  OR2_X1 U4218 ( .A1(n6248), .A2(n6207), .ZN(n6282) );
  OR2_X1 U4219 ( .A1(n6248), .A2(n6244), .ZN(n6313) );
  NAND2_X1 U4220 ( .A1(n6413), .A2(n6285), .ZN(n6357) );
  OR2_X1 U4221 ( .A1(n5911), .A2(n5862), .ZN(n6379) );
  OR2_X1 U4222 ( .A1(n5911), .A2(n5892), .ZN(n6444) );
  OR2_X1 U4223 ( .A1(n5911), .A2(n5878), .ZN(n6962) );
  NAND2_X1 U4224 ( .A1(n6413), .A2(n6108), .ZN(n6473) );
  INV_X1 U4225 ( .A(n6594), .ZN(n6533) );
  AND2_X1 U4226 ( .A1(n6541), .A2(STATE_REG_1__SCAN_IN), .ZN(n6625) );
  INV_X1 U4227 ( .A(n6587), .ZN(n6586) );
  NAND2_X1 U4228 ( .A1(n4486), .A2(n4485), .ZN(U2796) );
  OAI21_X1 U4229 ( .B1(n5197), .B2(n5824), .A(n4252), .ZN(U2990) );
  AND2_X4 U4230 ( .A1(n3777), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n6659)
         );
  AOI22_X1 U4231 ( .A1(n4433), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n4364), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3260) );
  AOI22_X1 U4232 ( .A1(n3362), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3259) );
  NAND2_X1 U4233 ( .A1(n3260), .A2(n3259), .ZN(n3264) );
  AOI22_X1 U4234 ( .A1(n4428), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3262) );
  AND2_X2 U4235 ( .A1(n3711), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3267)
         );
  AOI22_X1 U4236 ( .A1(n4435), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n3261) );
  NAND2_X1 U4237 ( .A1(n3262), .A2(n3261), .ZN(n3263) );
  NOR2_X1 U4238 ( .A1(n3264), .A2(n3263), .ZN(n3275) );
  AND2_X2 U4239 ( .A1(n6659), .A2(n3267), .ZN(n3363) );
  AND2_X4 U4240 ( .A1(n4554), .A2(n3268), .ZN(n4407) );
  AOI22_X1 U4241 ( .A1(n3363), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3274) );
  AOI22_X1 U4242 ( .A1(n3383), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3265) );
  INV_X1 U4243 ( .A(n3265), .ZN(n3272) );
  AND2_X2 U4244 ( .A1(n3267), .A2(n4660), .ZN(n3465) );
  AND2_X4 U4245 ( .A1(n6659), .A2(n4554), .ZN(n4277) );
  AOI22_X1 U4246 ( .A1(n3112), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3378), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3269) );
  NAND2_X1 U4247 ( .A1(n3270), .A2(n3269), .ZN(n3271) );
  NOR2_X1 U4248 ( .A1(n3272), .A2(n3271), .ZN(n3273) );
  AND3_X2 U4249 ( .A1(n3275), .A2(n3274), .A3(n3273), .ZN(n3393) );
  NAND2_X1 U4250 ( .A1(n3362), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n3279) );
  NAND2_X1 U4251 ( .A1(n4433), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3278) );
  NAND2_X1 U4252 ( .A1(n3112), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3277) );
  NAND2_X1 U4253 ( .A1(n3117), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3276) );
  NAND2_X1 U4254 ( .A1(n3107), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3283) );
  NAND2_X1 U4255 ( .A1(n3363), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n3282) );
  NAND2_X1 U4256 ( .A1(n4428), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n3281)
         );
  NAND2_X1 U4257 ( .A1(n3103), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3280)
         );
  NAND2_X1 U4258 ( .A1(n3121), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3287)
         );
  NAND2_X1 U4259 ( .A1(n4359), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3286)
         );
  NAND2_X1 U4260 ( .A1(n3465), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3285)
         );
  NAND2_X1 U4261 ( .A1(n4346), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3284)
         );
  NAND2_X1 U4262 ( .A1(n4364), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3291) );
  NAND2_X1 U4263 ( .A1(n4435), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3290) );
  NAND2_X1 U4264 ( .A1(n3378), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3289) );
  NAND2_X1 U4265 ( .A1(n3101), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n3288) );
  NAND4_X4 U4266 ( .A1(n3295), .A2(n3294), .A3(n3293), .A4(n3292), .ZN(n3402)
         );
  INV_X1 U4267 ( .A(n3402), .ZN(n3390) );
  AOI22_X1 U4268 ( .A1(n4407), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4428), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n3300) );
  AOI22_X1 U4269 ( .A1(n4364), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n4435), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3299) );
  AOI22_X1 U4270 ( .A1(n3377), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3102), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3297) );
  AND2_X1 U4271 ( .A1(n3297), .A2(n3296), .ZN(n3298) );
  NAND3_X1 U4272 ( .A1(n3300), .A2(n3299), .A3(n3298), .ZN(n3306) );
  AOI22_X1 U4273 ( .A1(n3383), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_12__7__SCAN_IN), .ZN(n3304) );
  AOI22_X1 U4274 ( .A1(n3378), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3101), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n3303) );
  AOI22_X1 U4275 ( .A1(n4433), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3302) );
  AOI22_X1 U4276 ( .A1(n4359), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3465), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3301) );
  NAND4_X1 U4277 ( .A1(n3304), .A2(n3303), .A3(n3302), .A4(n3301), .ZN(n3305)
         );
  OR2_X4 U4278 ( .A1(n3306), .A2(n3305), .ZN(n5906) );
  AOI22_X1 U4279 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n4407), .B1(n4428), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n3309) );
  NAND3_X1 U4280 ( .A1(n3309), .A2(n3308), .A3(n3307), .ZN(n3313) );
  AOI22_X1 U4281 ( .A1(n4359), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3465), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3311) );
  AOI22_X1 U4282 ( .A1(n3121), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3108), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3310) );
  NAND2_X1 U4283 ( .A1(n3311), .A2(n3310), .ZN(n3312) );
  NOR2_X1 U4284 ( .A1(n3313), .A2(n3312), .ZN(n3319) );
  AOI22_X1 U4285 ( .A1(n4435), .A2(INSTQUEUE_REG_2__4__SCAN_IN), .B1(n3378), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3317) );
  AOI22_X1 U4286 ( .A1(n4277), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3316) );
  AOI22_X1 U4287 ( .A1(n4433), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n3315) );
  NAND2_X1 U4288 ( .A1(n4277), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3324) );
  NAND2_X1 U4289 ( .A1(n4433), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3323) );
  NAND2_X1 U4290 ( .A1(n4364), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3322) );
  NAND2_X1 U4291 ( .A1(n3320), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n3321) );
  NAND2_X1 U4292 ( .A1(n3383), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3328)
         );
  NAND2_X1 U4293 ( .A1(n4428), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .ZN(n3327)
         );
  NAND2_X1 U4294 ( .A1(n4359), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3326)
         );
  NAND2_X1 U4295 ( .A1(n3465), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .ZN(n3325)
         );
  NAND2_X1 U4296 ( .A1(n3377), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3332) );
  NAND2_X1 U4297 ( .A1(n3362), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3331) );
  NAND2_X1 U4298 ( .A1(n4435), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3330) );
  NAND2_X1 U4299 ( .A1(n3378), .A2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3329) );
  NAND2_X1 U4300 ( .A1(n3363), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3337) );
  NAND2_X1 U4301 ( .A1(n3107), .A2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3336) );
  NAND2_X1 U4302 ( .A1(n3333), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3335)
         );
  NAND2_X1 U4303 ( .A1(n4346), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3334)
         );
  NAND2_X1 U4304 ( .A1(n4364), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3345) );
  NAND2_X1 U4305 ( .A1(n3112), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3344) );
  NAND2_X1 U4306 ( .A1(n3362), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n3343) );
  NAND2_X1 U4307 ( .A1(n3378), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3342) );
  NAND2_X1 U4308 ( .A1(n3107), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3349) );
  NAND2_X1 U4309 ( .A1(n4428), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n3348)
         );
  NAND2_X1 U4310 ( .A1(n4359), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3347)
         );
  NAND2_X1 U4311 ( .A1(n3109), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3346)
         );
  NAND2_X1 U4312 ( .A1(n3117), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3353) );
  NAND2_X1 U4313 ( .A1(n3383), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3352)
         );
  NAND2_X1 U4314 ( .A1(n3465), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3351)
         );
  NAND2_X1 U4315 ( .A1(n3333), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3350)
         );
  NAND2_X1 U4316 ( .A1(n4433), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3357) );
  NAND2_X1 U4317 ( .A1(n3363), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3356) );
  NAND2_X1 U4318 ( .A1(n4435), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3355) );
  NAND2_X1 U4319 ( .A1(n3320), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3354) );
  AND2_X4 U4320 ( .A1(n3408), .A2(n3100), .ZN(n3428) );
  NAND2_X1 U4321 ( .A1(n3445), .A2(n3428), .ZN(n3376) );
  AOI22_X1 U4322 ( .A1(n3362), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3363), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3367) );
  AOI22_X1 U4323 ( .A1(n3107), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n4428), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n3366) );
  AOI22_X1 U4324 ( .A1(n3105), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3320), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3365) );
  AOI22_X1 U4325 ( .A1(n3383), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3364) );
  NAND4_X1 U4326 ( .A1(n3367), .A2(n3366), .A3(n3365), .A4(n3364), .ZN(n3373)
         );
  AOI22_X1 U4327 ( .A1(n4277), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n4364), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3371) );
  AOI22_X1 U4328 ( .A1(n4359), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3465), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3370) );
  AOI22_X1 U4329 ( .A1(n4435), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3378), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3369) );
  AOI22_X1 U4330 ( .A1(n3377), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3368) );
  NAND4_X1 U4331 ( .A1(n3371), .A2(n3370), .A3(n3369), .A4(n3368), .ZN(n3372)
         );
  INV_X1 U4332 ( .A(n4119), .ZN(n3375) );
  NAND2_X1 U4333 ( .A1(n3375), .A2(n3374), .ZN(n4544) );
  OAI21_X1 U4334 ( .B1(n4604), .B2(n3398), .A(n5906), .ZN(n4212) );
  AOI22_X1 U4335 ( .A1(n3105), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3362), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3382) );
  AOI22_X1 U4336 ( .A1(n4277), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3117), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3381) );
  AOI22_X1 U4337 ( .A1(n4435), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3378), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3380) );
  AOI22_X1 U4338 ( .A1(n4364), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3320), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3379) );
  NAND4_X1 U4339 ( .A1(n3382), .A2(n3381), .A3(n3380), .A4(n3379), .ZN(n3389)
         );
  AOI22_X1 U4340 ( .A1(n3363), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3387) );
  AOI22_X1 U4341 ( .A1(n4359), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3465), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3386) );
  AOI22_X1 U4342 ( .A1(n4407), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n4428), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n3385) );
  AOI22_X1 U4343 ( .A1(n3120), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3384) );
  NAND4_X1 U4344 ( .A1(n3387), .A2(n3386), .A3(n3385), .A4(n3384), .ZN(n3388)
         );
  NOR2_X1 U4345 ( .A1(n4212), .A2(n4215), .ZN(n3757) );
  XNOR2_X1 U4346 ( .A(STATE_REG_1__SCAN_IN), .B(STATE_REG_2__SCAN_IN), .ZN(
        n4088) );
  NAND2_X1 U4347 ( .A1(n3405), .A2(n3719), .ZN(n3391) );
  NAND3_X1 U4348 ( .A1(n3427), .A2(n3757), .A3(n3391), .ZN(n3392) );
  NAND2_X1 U4349 ( .A1(n3392), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3421) );
  NAND2_X1 U4350 ( .A1(n3434), .A2(n4097), .ZN(n3395) );
  NAND2_X1 U4351 ( .A1(n3393), .A2(n3398), .ZN(n3394) );
  NAND3_X1 U4352 ( .A1(n3395), .A2(n4496), .A3(n3394), .ZN(n3396) );
  NAND2_X1 U4353 ( .A1(n4604), .A2(n5888), .ZN(n3429) );
  NAND2_X1 U4354 ( .A1(n3442), .A2(n3408), .ZN(n3401) );
  INV_X1 U4355 ( .A(n4604), .ZN(n3399) );
  INV_X1 U4356 ( .A(n3445), .ZN(n3403) );
  NAND2_X1 U4357 ( .A1(n4456), .A2(n3405), .ZN(n3411) );
  NAND2_X1 U4358 ( .A1(n3097), .A2(n3442), .ZN(n4114) );
  NAND2_X1 U4359 ( .A1(n3410), .A2(n5906), .ZN(n4108) );
  NAND3_X1 U4360 ( .A1(n3411), .A2(n4114), .A3(n4208), .ZN(n3412) );
  NAND2_X1 U4361 ( .A1(n3412), .A2(STATE2_REG_0__SCAN_IN), .ZN(n3414) );
  INV_X1 U4362 ( .A(n4076), .ZN(n3419) );
  XNOR2_X1 U4363 ( .A(n6316), .B(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6363)
         );
  INV_X1 U4364 ( .A(n3755), .ZN(n3420) );
  AND2_X1 U4365 ( .A1(n3420), .A2(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3413)
         );
  OAI211_X1 U4366 ( .C1(n3502), .C2(n3206), .A(n3414), .B(n3415), .ZN(n3499)
         );
  INV_X1 U4367 ( .A(n3414), .ZN(n3417) );
  INV_X1 U4368 ( .A(n3415), .ZN(n3416) );
  NAND2_X1 U4369 ( .A1(n3417), .A2(n3255), .ZN(n3418) );
  MUX2_X1 U4370 ( .A(n3420), .B(n3419), .S(n6316), .Z(n3424) );
  INV_X1 U4371 ( .A(n3424), .ZN(n3422) );
  NAND3_X1 U4372 ( .A1(n3423), .A2(n3422), .A3(n3421), .ZN(n3426) );
  INV_X1 U4373 ( .A(n3427), .ZN(n3433) );
  NAND2_X1 U4374 ( .A1(n3429), .A2(n3428), .ZN(n3431) );
  OR2_X1 U4375 ( .A1(n6614), .A2(n6521), .ZN(n6524) );
  INV_X1 U4376 ( .A(n6524), .ZN(n3430) );
  NAND2_X1 U4377 ( .A1(n3431), .A2(n3430), .ZN(n3432) );
  NOR2_X1 U4378 ( .A1(n3433), .A2(n3432), .ZN(n3448) );
  INV_X1 U4379 ( .A(n3444), .ZN(n3436) );
  NAND2_X1 U4380 ( .A1(n3436), .A2(n3408), .ZN(n3437) );
  NAND2_X1 U4381 ( .A1(n3437), .A2(n4495), .ZN(n3441) );
  NAND2_X1 U4382 ( .A1(n3095), .A2(n3397), .ZN(n4507) );
  NAND2_X1 U4383 ( .A1(n4507), .A2(n3409), .ZN(n3439) );
  NAND2_X1 U4384 ( .A1(n3440), .A2(n3439), .ZN(n4213) );
  INV_X1 U4385 ( .A(n3442), .ZN(n3443) );
  NAND2_X1 U4386 ( .A1(n3443), .A2(n4812), .ZN(n4219) );
  NAND3_X1 U4387 ( .A1(n6475), .A2(n3397), .A3(n3445), .ZN(n3446) );
  NAND4_X1 U4388 ( .A1(n3448), .A2(n3447), .A3(n4219), .A4(n3446), .ZN(n3479)
         );
  XNOR2_X1 U4389 ( .A(n3501), .B(n3500), .ZN(n4542) );
  NAND2_X1 U4390 ( .A1(n4542), .A2(n6521), .ZN(n3460) );
  AOI22_X1 U4391 ( .A1(n3112), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3110), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3452) );
  AOI22_X1 U4392 ( .A1(n3116), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n3451) );
  AOI22_X1 U4393 ( .A1(n3106), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n3450) );
  AOI22_X1 U4394 ( .A1(n4427), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3449) );
  NAND4_X1 U4395 ( .A1(n3452), .A2(n3451), .A3(n3450), .A4(n3449), .ZN(n3458)
         );
  AOI22_X1 U4396 ( .A1(n3114), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_12__1__SCAN_IN), .ZN(n3456) );
  AOI22_X1 U4397 ( .A1(n3121), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3465), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3455) );
  AOI22_X1 U4398 ( .A1(n4341), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3454) );
  AOI22_X1 U4399 ( .A1(n4407), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n4346), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3453) );
  NAND4_X1 U4400 ( .A1(n3456), .A2(n3455), .A3(n3454), .A4(n3453), .ZN(n3457)
         );
  NAND2_X1 U4401 ( .A1(n3518), .A2(n3582), .ZN(n3459) );
  NAND2_X1 U4402 ( .A1(n3460), .A2(n3459), .ZN(n3478) );
  INV_X1 U4403 ( .A(n3478), .ZN(n3476) );
  INV_X1 U4404 ( .A(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3474) );
  AOI22_X1 U4405 ( .A1(n4341), .A2(INSTQUEUE_REG_10__7__SCAN_IN), .B1(n3112), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n3464) );
  AOI22_X1 U4406 ( .A1(n3116), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3463) );
  AOI22_X1 U4407 ( .A1(n4435), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3378), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3462) );
  AOI22_X1 U4408 ( .A1(n4427), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n4346), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3461) );
  NAND4_X1 U4409 ( .A1(n3464), .A2(n3463), .A3(n3462), .A4(n3461), .ZN(n3471)
         );
  AOI22_X1 U4410 ( .A1(n3362), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n3469) );
  AOI22_X1 U4411 ( .A1(n3383), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3465), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n3468) );
  AOI22_X1 U4412 ( .A1(n3110), .A2(INSTQUEUE_REG_5__7__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n3467) );
  AOI22_X1 U4413 ( .A1(n3118), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3466) );
  NAND4_X1 U4414 ( .A1(n3469), .A2(n3468), .A3(n3467), .A4(n3466), .ZN(n3470)
         );
  NAND2_X1 U4415 ( .A1(n3518), .A2(n3669), .ZN(n3473) );
  NAND2_X1 U4416 ( .A1(n3521), .A2(n3582), .ZN(n3472) );
  OAI211_X1 U4417 ( .C1(n3744), .C2(n3474), .A(n3473), .B(n3472), .ZN(n3477)
         );
  INV_X1 U4418 ( .A(n3479), .ZN(n3480) );
  NAND2_X1 U4419 ( .A1(n6179), .A2(n6521), .ZN(n3493) );
  AOI22_X1 U4420 ( .A1(n3114), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3485) );
  AOI22_X1 U4421 ( .A1(n4388), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3107), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3484) );
  AOI22_X1 U4422 ( .A1(n4427), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3483) );
  AOI22_X1 U4423 ( .A1(n4341), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3482) );
  NAND4_X1 U4424 ( .A1(n3485), .A2(n3484), .A3(n3483), .A4(n3482), .ZN(n3491)
         );
  AOI22_X1 U4425 ( .A1(n4277), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3110), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3489) );
  AOI22_X1 U4426 ( .A1(n3106), .A2(INSTQUEUE_REG_3__0__SCAN_IN), .B1(n3378), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3488) );
  AOI22_X1 U4427 ( .A1(n3121), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n3487) );
  AOI22_X1 U4428 ( .A1(n3118), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3486) );
  NAND4_X1 U4429 ( .A1(n3489), .A2(n3488), .A3(n3487), .A4(n3486), .ZN(n3490)
         );
  XNOR2_X1 U4430 ( .A(n3669), .B(n3595), .ZN(n3492) );
  NAND2_X1 U4431 ( .A1(n3492), .A2(n3518), .ZN(n3591) );
  NAND2_X1 U4432 ( .A1(n3493), .A2(n3591), .ZN(n3588) );
  INV_X1 U4433 ( .A(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3496) );
  AOI21_X1 U4434 ( .B1(n3435), .B2(n3671), .A(n6521), .ZN(n3495) );
  NAND2_X1 U4435 ( .A1(n3438), .A2(n3595), .ZN(n3494) );
  NOR2_X1 U4436 ( .A1(n3669), .A2(n3533), .ZN(n3497) );
  INV_X1 U4437 ( .A(n3601), .ZN(n3524) );
  NAND2_X1 U4438 ( .A1(n3527), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3507) );
  NAND2_X1 U4439 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3503) );
  NAND2_X1 U4440 ( .A1(n3503), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3504) );
  NOR2_X1 U4441 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6483), .ZN(n6208)
         );
  NAND2_X1 U4442 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6208), .ZN(n5980) );
  OAI22_X1 U4443 ( .A1(n4076), .A2(n5871), .B1(n3755), .B2(n6489), .ZN(n3505)
         );
  INV_X1 U4444 ( .A(n3505), .ZN(n3506) );
  XNOR2_X1 U4445 ( .A(n3525), .B(n3526), .ZN(n4651) );
  NAND2_X1 U4446 ( .A1(n4651), .A2(n6521), .ZN(n3520) );
  AOI22_X1 U4447 ( .A1(n4341), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_8__2__SCAN_IN), .ZN(n3511) );
  AOI22_X1 U4448 ( .A1(n4277), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3510) );
  INV_X1 U4449 ( .A(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n6930) );
  AOI22_X1 U4450 ( .A1(n3106), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3509) );
  AOI22_X1 U4451 ( .A1(n3110), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3508) );
  NAND4_X1 U4452 ( .A1(n3511), .A2(n3510), .A3(n3509), .A4(n3508), .ZN(n3517)
         );
  AOI22_X1 U4453 ( .A1(n3107), .A2(INSTQUEUE_REG_2__2__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3515) );
  AOI22_X1 U4454 ( .A1(n4427), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3514) );
  AOI22_X1 U4455 ( .A1(n4388), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3513) );
  AOI22_X1 U4456 ( .A1(n3383), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3108), 
        .B2(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n3512) );
  NAND4_X1 U4457 ( .A1(n3515), .A2(n3514), .A3(n3513), .A4(n3512), .ZN(n3516)
         );
  NAND2_X1 U4458 ( .A1(n3518), .A2(n3573), .ZN(n3519) );
  AOI22_X1 U4459 ( .A1(n3707), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3521), 
        .B2(n3573), .ZN(n3522) );
  INV_X1 U4460 ( .A(n3609), .ZN(n3547) );
  NAND2_X1 U4461 ( .A1(n3527), .A2(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .ZN(n3532) );
  NAND3_X1 U4462 ( .A1(n6368), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A3(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n6115) );
  INV_X1 U4463 ( .A(n6115), .ZN(n3528) );
  NAND2_X1 U4464 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n3528), .ZN(n6138) );
  NAND2_X1 U4465 ( .A1(n6368), .A2(n6138), .ZN(n3529) );
  NOR3_X1 U4466 ( .A1(n6368), .A2(n6489), .A3(n6483), .ZN(n6420) );
  NAND2_X1 U4467 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6420), .ZN(n6406) );
  NAND2_X1 U4468 ( .A1(n3529), .A2(n6406), .ZN(n6145) );
  OAI22_X1 U4469 ( .A1(n4076), .A2(n6145), .B1(n3755), .B2(n6368), .ZN(n3530)
         );
  INV_X1 U4470 ( .A(n3530), .ZN(n3531) );
  XNOR2_X2 U4471 ( .A(n4674), .B(n6020), .ZN(n6211) );
  AOI22_X1 U4472 ( .A1(n4341), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3538) );
  AOI22_X1 U4473 ( .A1(n3112), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_9__3__SCAN_IN), .ZN(n3537) );
  AOI22_X1 U4474 ( .A1(n3106), .A2(INSTQUEUE_REG_3__3__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3536) );
  INV_X1 U4475 ( .A(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n6866) );
  AOI22_X1 U4476 ( .A1(n3110), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3535) );
  NAND4_X1 U4477 ( .A1(n3538), .A2(n3537), .A3(n3536), .A4(n3535), .ZN(n3544)
         );
  AOI22_X1 U4478 ( .A1(n4407), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3542) );
  AOI22_X1 U4479 ( .A1(n4427), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n3541) );
  AOI22_X1 U4480 ( .A1(n4388), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n3540) );
  AOI22_X1 U4481 ( .A1(n3121), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_13__3__SCAN_IN), .ZN(n3539) );
  NAND4_X1 U4482 ( .A1(n3542), .A2(n3541), .A3(n3540), .A4(n3539), .ZN(n3543)
         );
  AOI22_X1 U4483 ( .A1(n3707), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3752), 
        .B2(n3610), .ZN(n3545) );
  AOI22_X1 U4484 ( .A1(n4341), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3551) );
  AOI22_X1 U4485 ( .A1(n4277), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_9__4__SCAN_IN), .ZN(n3550) );
  AOI22_X1 U4486 ( .A1(n3106), .A2(INSTQUEUE_REG_3__4__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3549) );
  AOI22_X1 U4487 ( .A1(n3110), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n3548) );
  NAND4_X1 U4488 ( .A1(n3551), .A2(n3550), .A3(n3549), .A4(n3548), .ZN(n3557)
         );
  AOI22_X1 U4489 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n3107), .B1(n3118), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3555) );
  AOI22_X1 U4490 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n4427), .B1(n4434), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n3554) );
  AOI22_X1 U4491 ( .A1(n4388), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3553) );
  AOI22_X1 U4492 ( .A1(n3383), .A2(INSTQUEUE_REG_14__4__SCAN_IN), .B1(n4346), 
        .B2(INSTQUEUE_REG_13__4__SCAN_IN), .ZN(n3552) );
  NAND4_X1 U4493 ( .A1(n3555), .A2(n3554), .A3(n3553), .A4(n3552), .ZN(n3556)
         );
  AOI22_X1 U4494 ( .A1(n3707), .A2(INSTQUEUE_REG_0__4__SCAN_IN), .B1(n3752), 
        .B2(n3624), .ZN(n3619) );
  INV_X1 U4495 ( .A(n3622), .ZN(n3570) );
  AOI22_X1 U4496 ( .A1(n4341), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_8__5__SCAN_IN), .ZN(n3562) );
  AOI22_X1 U4497 ( .A1(n3112), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3561) );
  AOI22_X1 U4498 ( .A1(n3106), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3560) );
  AOI22_X1 U4499 ( .A1(n3110), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n3559) );
  NAND4_X1 U4500 ( .A1(n3562), .A2(n3561), .A3(n3560), .A4(n3559), .ZN(n3568)
         );
  AOI22_X1 U4501 ( .A1(n4407), .A2(INSTQUEUE_REG_2__5__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n3566) );
  AOI22_X1 U4502 ( .A1(n4427), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n3565) );
  AOI22_X1 U4503 ( .A1(n4388), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3564) );
  AOI22_X1 U4504 ( .A1(n3383), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3108), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3563) );
  NAND4_X1 U4505 ( .A1(n3566), .A2(n3565), .A3(n3564), .A4(n3563), .ZN(n3567)
         );
  AOI22_X1 U4506 ( .A1(n3707), .A2(INSTQUEUE_REG_0__5__SCAN_IN), .B1(n3752), 
        .B2(n3648), .ZN(n3571) );
  NAND2_X1 U4507 ( .A1(n3622), .A2(n3571), .ZN(n3572) );
  NAND2_X1 U4508 ( .A1(n3595), .A2(n3582), .ZN(n3602) );
  INV_X1 U4509 ( .A(n3573), .ZN(n3603) );
  NAND2_X1 U4510 ( .A1(n3602), .A2(n3603), .ZN(n3612) );
  NAND2_X1 U4511 ( .A1(n3612), .A2(n3610), .ZN(n3623) );
  INV_X1 U4512 ( .A(n3624), .ZN(n3574) );
  OR2_X1 U4513 ( .A1(n3623), .A2(n3574), .ZN(n3650) );
  XNOR2_X1 U4514 ( .A(n3650), .B(n3648), .ZN(n3575) );
  NAND2_X1 U4515 ( .A1(n3575), .A2(n3428), .ZN(n3576) );
  NAND2_X1 U4516 ( .A1(n3577), .A2(n3576), .ZN(n3631) );
  INV_X1 U4517 ( .A(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n4132) );
  XNOR2_X1 U4518 ( .A(n3631), .B(n4132), .ZN(n4725) );
  INV_X1 U4519 ( .A(n3578), .ZN(n3579) );
  NAND2_X1 U4520 ( .A1(n3132), .A2(n3579), .ZN(n3581) );
  NAND2_X1 U4521 ( .A1(n4688), .A2(n3706), .ZN(n3587) );
  OAI21_X1 U4522 ( .B1(n3595), .B2(n3582), .A(n3602), .ZN(n3584) );
  INV_X1 U4523 ( .A(n3428), .ZN(n6630) );
  INV_X1 U4524 ( .A(n4215), .ZN(n3583) );
  OAI211_X1 U4525 ( .C1(n3584), .C2(n6630), .A(n3583), .B(n3402), .ZN(n3585)
         );
  INV_X1 U4526 ( .A(n3585), .ZN(n3586) );
  NAND2_X1 U4527 ( .A1(n3587), .A2(n3586), .ZN(n4788) );
  NAND2_X1 U4528 ( .A1(n3588), .A2(n3589), .ZN(n3593) );
  INV_X1 U4529 ( .A(n3589), .ZN(n3590) );
  NAND2_X1 U4530 ( .A1(n3591), .A2(n3590), .ZN(n3592) );
  AND2_X1 U4531 ( .A1(n3438), .A2(n5888), .ZN(n3604) );
  INV_X1 U4532 ( .A(n3604), .ZN(n3594) );
  OAI21_X1 U4533 ( .B1(n6630), .B2(n3595), .A(n3594), .ZN(n3596) );
  INV_X1 U4534 ( .A(n3596), .ZN(n3597) );
  NAND2_X1 U4535 ( .A1(n3598), .A2(n3597), .ZN(n4580) );
  NAND2_X1 U4536 ( .A1(n4580), .A2(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n4581)
         );
  XNOR2_X1 U4537 ( .A(n4581), .B(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4787)
         );
  NAND2_X1 U4538 ( .A1(n4788), .A2(n4787), .ZN(n4786) );
  INV_X1 U4539 ( .A(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n5858) );
  OR2_X1 U4540 ( .A1(n4581), .A2(n5858), .ZN(n3599) );
  NAND2_X1 U4541 ( .A1(n4687), .A2(n3706), .ZN(n3607) );
  OAI21_X1 U4542 ( .B1(n3603), .B2(n3602), .A(n3612), .ZN(n3605) );
  AOI21_X1 U4543 ( .B1(n3605), .B2(n3428), .A(n3604), .ZN(n3606) );
  NAND2_X1 U4544 ( .A1(n3607), .A2(n3606), .ZN(n3608) );
  XNOR2_X2 U4545 ( .A(n3609), .B(n5863), .ZN(n3776) );
  INV_X1 U4546 ( .A(n3610), .ZN(n3611) );
  XNOR2_X1 U4547 ( .A(n3612), .B(n3611), .ZN(n3613) );
  NAND2_X1 U4548 ( .A1(n3613), .A2(n3428), .ZN(n3614) );
  INV_X1 U4549 ( .A(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3615) );
  NAND2_X1 U4550 ( .A1(n3616), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n3617)
         );
  NAND2_X1 U4551 ( .A1(n3620), .A2(n3619), .ZN(n3621) );
  INV_X1 U4552 ( .A(n3623), .ZN(n3625) );
  OAI211_X1 U4553 ( .C1(n3625), .C2(n3624), .A(n3428), .B(n3650), .ZN(n3626)
         );
  OAI21_X1 U4554 ( .B1(n3787), .B2(n3148), .A(n3626), .ZN(n3628) );
  INV_X1 U4555 ( .A(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3627) );
  XNOR2_X1 U4556 ( .A(n3628), .B(n3627), .ZN(n4756) );
  NAND2_X1 U4557 ( .A1(n4757), .A2(n4756), .ZN(n3630) );
  NAND2_X1 U4558 ( .A1(n3628), .A2(INSTADDRPOINTER_REG_4__SCAN_IN), .ZN(n3629)
         );
  NAND2_X1 U4559 ( .A1(n3630), .A2(n3629), .ZN(n4726) );
  NAND2_X1 U4560 ( .A1(n4725), .A2(n4726), .ZN(n3633) );
  NAND2_X1 U4561 ( .A1(n3631), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .ZN(n3632)
         );
  NAND2_X1 U4562 ( .A1(n3633), .A2(n3632), .ZN(n4768) );
  INV_X1 U4563 ( .A(n3646), .ZN(n3645) );
  AOI22_X1 U4564 ( .A1(n4277), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_8__6__SCAN_IN), .ZN(n3637) );
  AOI22_X1 U4565 ( .A1(n3116), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_12__6__SCAN_IN), .ZN(n3636) );
  AOI22_X1 U4566 ( .A1(n3107), .A2(INSTQUEUE_REG_2__6__SCAN_IN), .B1(n3383), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3635) );
  AOI22_X1 U4567 ( .A1(n4341), .A2(INSTQUEUE_REG_10__6__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n3634) );
  NAND4_X1 U4568 ( .A1(n3637), .A2(n3636), .A3(n3635), .A4(n3634), .ZN(n3643)
         );
  AOI22_X1 U4569 ( .A1(n3110), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n3641) );
  AOI22_X1 U4570 ( .A1(n4427), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3640) );
  AOI22_X1 U4571 ( .A1(n3106), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3639) );
  AOI22_X1 U4572 ( .A1(n4346), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3638) );
  NAND4_X1 U4573 ( .A1(n3641), .A2(n3640), .A3(n3639), .A4(n3638), .ZN(n3642)
         );
  AOI22_X1 U4574 ( .A1(n3707), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3752), 
        .B2(n3651), .ZN(n3647) );
  INV_X1 U4575 ( .A(n3647), .ZN(n3644) );
  NAND2_X1 U4576 ( .A1(n3646), .A2(n3647), .ZN(n3806) );
  NAND3_X1 U4577 ( .A1(n3668), .A2(n3706), .A3(n3806), .ZN(n3654) );
  INV_X1 U4578 ( .A(n3648), .ZN(n3649) );
  NOR2_X1 U4579 ( .A1(n3650), .A2(n3649), .ZN(n3652) );
  NAND2_X1 U4580 ( .A1(n3652), .A2(n3651), .ZN(n3673) );
  OAI211_X1 U4581 ( .C1(n3652), .C2(n3651), .A(n3673), .B(n3428), .ZN(n3653)
         );
  NAND2_X1 U4582 ( .A1(n3654), .A2(n3653), .ZN(n3656) );
  INV_X1 U4583 ( .A(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3655) );
  XNOR2_X1 U4584 ( .A(n3656), .B(n3655), .ZN(n4769) );
  NAND2_X1 U4585 ( .A1(n4768), .A2(n4769), .ZN(n3658) );
  NAND2_X1 U4586 ( .A1(n3656), .A2(INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n3657)
         );
  NAND2_X1 U4587 ( .A1(n3658), .A2(n3657), .ZN(n4731) );
  INV_X1 U4588 ( .A(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3660) );
  NAND2_X1 U4589 ( .A1(n3752), .A2(n3671), .ZN(n3659) );
  OAI21_X1 U4590 ( .B1(n3744), .B2(n3660), .A(n3659), .ZN(n3661) );
  NAND2_X1 U4591 ( .A1(n3820), .A2(n3706), .ZN(n3664) );
  XNOR2_X1 U4592 ( .A(n3673), .B(n3671), .ZN(n3662) );
  NAND2_X1 U4593 ( .A1(n3662), .A2(n3428), .ZN(n3663) );
  NAND2_X1 U4594 ( .A1(n3664), .A2(n3663), .ZN(n3665) );
  INV_X1 U4595 ( .A(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n4139) );
  XNOR2_X1 U4596 ( .A(n3665), .B(n4139), .ZN(n4732) );
  NAND2_X1 U4597 ( .A1(n4731), .A2(n4732), .ZN(n3667) );
  NAND2_X1 U4598 ( .A1(n3665), .A2(INSTADDRPOINTER_REG_7__SCAN_IN), .ZN(n3666)
         );
  NAND2_X1 U4599 ( .A1(n3667), .A2(n3666), .ZN(n4793) );
  NAND2_X1 U4600 ( .A1(n3428), .A2(n3671), .ZN(n3672) );
  OR2_X1 U4601 ( .A1(n3673), .A2(n3672), .ZN(n3674) );
  NAND2_X1 U4602 ( .A1(n3685), .A2(n3674), .ZN(n3675) );
  XNOR2_X1 U4603 ( .A(n3675), .B(n6759), .ZN(n4794) );
  NAND2_X1 U4604 ( .A1(n4793), .A2(n4794), .ZN(n3677) );
  NAND2_X1 U4605 ( .A1(n3675), .A2(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n3676)
         );
  NAND2_X1 U4606 ( .A1(n3677), .A2(n3676), .ZN(n4804) );
  INV_X1 U4607 ( .A(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n6751) );
  NOR2_X1 U4608 ( .A1(n5222), .A2(n6751), .ZN(n3678) );
  INV_X1 U4609 ( .A(n3678), .ZN(n3679) );
  NAND2_X1 U4610 ( .A1(n5245), .A2(n6751), .ZN(n3681) );
  INV_X1 U4611 ( .A(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4842) );
  AND2_X1 U4612 ( .A1(n5245), .A2(n4842), .ZN(n4836) );
  INV_X1 U4613 ( .A(INSTADDRPOINTER_REG_11__SCAN_IN), .ZN(n6798) );
  NAND2_X1 U4614 ( .A1(n5245), .A2(n6798), .ZN(n4881) );
  OR2_X1 U4615 ( .A1(n5222), .A2(n6798), .ZN(n4882) );
  INV_X1 U4616 ( .A(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6916) );
  NAND2_X1 U4617 ( .A1(n5245), .A2(n6916), .ZN(n3682) );
  NAND2_X1 U4618 ( .A1(n4891), .A2(n3682), .ZN(n3684) );
  OR2_X1 U4619 ( .A1(n5245), .A2(n6916), .ZN(n3683) );
  INV_X1 U4620 ( .A(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5545) );
  XNOR2_X1 U4621 ( .A(n5245), .B(n5545), .ZN(n4940) );
  NAND2_X1 U4622 ( .A1(n5222), .A2(n5545), .ZN(n3686) );
  INV_X1 U4623 ( .A(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n5534) );
  NAND2_X1 U4624 ( .A1(n5245), .A2(n5534), .ZN(n3688) );
  INV_X1 U4625 ( .A(INSTADDRPOINTER_REG_15__SCAN_IN), .ZN(n6844) );
  OR2_X1 U4626 ( .A1(n5245), .A2(n6844), .ZN(n3689) );
  NAND2_X1 U4627 ( .A1(n5245), .A2(n6844), .ZN(n3690) );
  INV_X1 U4628 ( .A(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6828) );
  NAND2_X1 U4629 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n4244) );
  INV_X1 U4630 ( .A(INSTADDRPOINTER_REG_19__SCAN_IN), .ZN(n6854) );
  NOR2_X1 U4631 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n3692) );
  OR2_X1 U4632 ( .A1(n5245), .A2(n3692), .ZN(n3693) );
  INV_X1 U4633 ( .A(n5369), .ZN(n3696) );
  NAND2_X1 U4634 ( .A1(n3691), .A2(n3696), .ZN(n5221) );
  INV_X1 U4635 ( .A(INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5364) );
  XNOR2_X1 U4636 ( .A(n5245), .B(n5364), .ZN(n5239) );
  INV_X1 U4637 ( .A(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n5349) );
  XNOR2_X1 U4638 ( .A(n5245), .B(n5349), .ZN(n5231) );
  NOR2_X1 U4639 ( .A1(n5222), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5214)
         );
  AOI21_X1 U4640 ( .B1(INSTADDRPOINTER_REG_22__SCAN_IN), .B2(n5222), .A(n5214), 
        .ZN(n3698) );
  XNOR2_X1 U4641 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .ZN(n3708) );
  NAND2_X1 U4642 ( .A1(n3710), .A2(n3708), .ZN(n3701) );
  NAND2_X1 U4643 ( .A1(n6483), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3700) );
  NAND2_X1 U4644 ( .A1(n3701), .A2(n3700), .ZN(n3732) );
  XNOR2_X1 U4645 ( .A(n3258), .B(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n3731)
         );
  INV_X1 U4646 ( .A(n3731), .ZN(n3702) );
  NAND2_X1 U4647 ( .A1(n3732), .A2(n3702), .ZN(n3704) );
  NAND2_X1 U4648 ( .A1(n6489), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n3703) );
  NAND2_X1 U4649 ( .A1(n3704), .A2(n3703), .ZN(n3741) );
  XNOR2_X1 U4650 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(
        INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n3740) );
  NOR2_X1 U4651 ( .A1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .A2(n5861), .ZN(n3705)
         );
  NAND2_X1 U4652 ( .A1(n4095), .A2(n3745), .ZN(n3751) );
  INV_X1 U4653 ( .A(n3708), .ZN(n3709) );
  XNOR2_X1 U4654 ( .A(n3709), .B(n3710), .ZN(n4092) );
  INV_X1 U4655 ( .A(n3745), .ZN(n3730) );
  INV_X1 U4656 ( .A(n3710), .ZN(n3713) );
  NAND2_X1 U4657 ( .A1(n3711), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .ZN(n3712) );
  NAND2_X1 U4658 ( .A1(n3713), .A2(n3712), .ZN(n3721) );
  INV_X1 U4659 ( .A(n3721), .ZN(n3716) );
  INV_X1 U4660 ( .A(n3714), .ZN(n3715) );
  AOI21_X1 U4661 ( .B1(n3758), .B2(n3716), .A(n3715), .ZN(n3725) );
  NAND2_X1 U4662 ( .A1(n3408), .A2(n3402), .ZN(n3718) );
  NAND2_X1 U4663 ( .A1(n3717), .A2(n3718), .ZN(n3733) );
  AOI21_X1 U4664 ( .B1(n3752), .B2(n3397), .A(n3719), .ZN(n3726) );
  INV_X1 U4665 ( .A(n4092), .ZN(n3720) );
  NAND2_X1 U4666 ( .A1(n3726), .A2(n3720), .ZN(n3724) );
  INV_X1 U4667 ( .A(n3752), .ZN(n3722) );
  OAI21_X1 U4668 ( .B1(n3722), .B2(n3721), .A(n3730), .ZN(n3723) );
  OAI211_X1 U4669 ( .C1(n3725), .C2(n3733), .A(n3724), .B(n3723), .ZN(n3729)
         );
  INV_X1 U4670 ( .A(n3726), .ZN(n3727) );
  NAND3_X1 U4671 ( .A1(n3727), .A2(STATE2_REG_0__SCAN_IN), .A3(n4092), .ZN(
        n3728) );
  OAI211_X1 U4672 ( .C1(n4092), .C2(n3730), .A(n3729), .B(n3728), .ZN(n3738)
         );
  XNOR2_X1 U4673 ( .A(n3732), .B(n3731), .ZN(n4091) );
  INV_X1 U4674 ( .A(n3733), .ZN(n3735) );
  NAND2_X1 U4675 ( .A1(n3752), .A2(n4091), .ZN(n3734) );
  OAI211_X1 U4676 ( .C1(n4091), .C2(n3744), .A(n3735), .B(n3734), .ZN(n3737)
         );
  NOR2_X1 U4677 ( .A1(n3735), .A2(n3734), .ZN(n3736) );
  AOI21_X1 U4678 ( .B1(n3738), .B2(n3737), .A(n3736), .ZN(n3749) );
  NAND3_X1 U4679 ( .A1(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A2(n3739), .A3(n5548), .ZN(n4093) );
  NOR2_X1 U4680 ( .A1(n3741), .A2(n3740), .ZN(n3742) );
  NOR2_X1 U4681 ( .A1(n3743), .A2(n3742), .ZN(n4090) );
  NAND2_X1 U4682 ( .A1(n4093), .A2(n4090), .ZN(n3746) );
  AOI22_X1 U4683 ( .A1(n3746), .A2(n3745), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n6521), .ZN(n3747) );
  OAI21_X1 U4684 ( .B1(n3749), .B2(n3748), .A(n3747), .ZN(n3750) );
  NAND2_X1 U4685 ( .A1(n3751), .A2(n3750), .ZN(n3754) );
  NAND2_X1 U4686 ( .A1(n4095), .A2(n3752), .ZN(n3753) );
  NAND2_X1 U4687 ( .A1(n6475), .A2(n3438), .ZN(n3756) );
  NAND2_X1 U4688 ( .A1(n3757), .A2(n3756), .ZN(n4116) );
  NAND2_X1 U4689 ( .A1(n5334), .A2(n5774), .ZN(n4081) );
  NAND2_X1 U4690 ( .A1(n4688), .A2(n3944), .ZN(n3762) );
  AOI22_X1 U4691 ( .A1(n4453), .A2(EAX_REG_1__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n6511), .ZN(n3760) );
  INV_X1 U4692 ( .A(n4108), .ZN(n4979) );
  NAND2_X1 U4693 ( .A1(n3763), .A2(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n3759) );
  AND2_X1 U4694 ( .A1(n3760), .A2(n3759), .ZN(n3761) );
  NAND2_X1 U4695 ( .A1(n3131), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4595) );
  NAND2_X1 U4696 ( .A1(n3764), .A2(EAX_REG_0__SCAN_IN), .ZN(n3766) );
  NAND2_X1 U4697 ( .A1(n6511), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n3765)
         );
  OAI211_X1 U4698 ( .C1(n3790), .C2(n3711), .A(n3766), .B(n3765), .ZN(n3767)
         );
  AOI21_X1 U4699 ( .B1(n6179), .B2(n3944), .A(n3767), .ZN(n3768) );
  OR2_X1 U4700 ( .A1(n4595), .A2(n3768), .ZN(n4596) );
  INV_X1 U4701 ( .A(n3768), .ZN(n4597) );
  OR2_X1 U4702 ( .A1(n4597), .A2(n3791), .ZN(n3769) );
  NAND2_X1 U4703 ( .A1(n4596), .A2(n3769), .ZN(n4607) );
  NAND2_X1 U4704 ( .A1(n4687), .A2(n3944), .ZN(n3770) );
  NAND2_X1 U4705 ( .A1(n6511), .A2(STATEBS16_REG_SCAN_IN), .ZN(n3901) );
  OAI21_X1 U4706 ( .B1(PHYADDRPOINTER_REG_1__SCAN_IN), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .A(n3779), .ZN(n5772) );
  AOI22_X1 U4707 ( .A1(n4448), .A2(n5772), .B1(n4452), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n3772) );
  NAND2_X1 U4708 ( .A1(n4453), .A2(EAX_REG_2__SCAN_IN), .ZN(n3771) );
  OAI211_X1 U4709 ( .C1(n3790), .C2(n3258), .A(n3772), .B(n3771), .ZN(n4648)
         );
  NAND2_X1 U4710 ( .A1(n3773), .A2(n4610), .ZN(n3774) );
  NAND2_X1 U4711 ( .A1(n3776), .A2(n3944), .ZN(n3786) );
  INV_X1 U4712 ( .A(n3779), .ZN(n3778) );
  INV_X1 U4713 ( .A(n3792), .ZN(n3793) );
  INV_X1 U4714 ( .A(PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3780) );
  NAND2_X1 U4715 ( .A1(n3780), .A2(n3779), .ZN(n3781) );
  NAND2_X1 U4716 ( .A1(n3793), .A2(n3781), .ZN(n5664) );
  AOI22_X1 U4717 ( .A1(n5664), .A2(n4448), .B1(n4452), .B2(
        PHYADDRPOINTER_REG_3__SCAN_IN), .ZN(n3783) );
  NAND2_X1 U4718 ( .A1(n4453), .A2(EAX_REG_3__SCAN_IN), .ZN(n3782) );
  OAI211_X1 U4719 ( .C1(n3790), .C2(n3777), .A(n3783), .B(n3782), .ZN(n3784)
         );
  INV_X1 U4720 ( .A(n3784), .ZN(n3785) );
  NAND2_X1 U4721 ( .A1(n3786), .A2(n3785), .ZN(n4644) );
  INV_X1 U4722 ( .A(n3944), .ZN(n3851) );
  NAND2_X1 U4723 ( .A1(n6511), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n3789)
         );
  NAND2_X1 U4724 ( .A1(n4453), .A2(EAX_REG_4__SCAN_IN), .ZN(n3788) );
  OAI211_X1 U4725 ( .C1(n3790), .C2(n5548), .A(n3789), .B(n3788), .ZN(n3797)
         );
  INV_X1 U4726 ( .A(n3802), .ZN(n3795) );
  INV_X1 U4727 ( .A(PHYADDRPOINTER_REG_4__SCAN_IN), .ZN(n6837) );
  NAND2_X1 U4728 ( .A1(n3793), .A2(n6837), .ZN(n3794) );
  NAND2_X1 U4729 ( .A1(n3795), .A2(n3794), .ZN(n5661) );
  AND2_X1 U4730 ( .A1(n5661), .A2(n4448), .ZN(n3796) );
  AOI21_X1 U4731 ( .B1(n3797), .B2(n3791), .A(n3796), .ZN(n3798) );
  NOR2_X2 U4732 ( .A1(n4642), .A2(n4695), .ZN(n4693) );
  OAI21_X1 U4733 ( .B1(n3802), .B2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n3814), 
        .ZN(n5642) );
  AOI22_X1 U4734 ( .A1(n5642), .A2(n4448), .B1(n4452), .B2(
        PHYADDRPOINTER_REG_5__SCAN_IN), .ZN(n3803) );
  NAND2_X1 U4735 ( .A1(n3806), .A2(n3944), .ZN(n3812) );
  INV_X1 U4736 ( .A(EAX_REG_6__SCAN_IN), .ZN(n3808) );
  OAI21_X1 U4737 ( .B1(PHYADDRPOINTER_REG_6__SCAN_IN), .B2(n6286), .A(n6511), 
        .ZN(n3807) );
  OAI21_X1 U4738 ( .B1(n4399), .B2(n3808), .A(n3807), .ZN(n3810) );
  XOR2_X1 U4739 ( .A(n3813), .B(n3814), .Z(n5630) );
  NAND2_X1 U4740 ( .A1(n5630), .A2(n4448), .ZN(n3809) );
  NAND2_X1 U4741 ( .A1(n3810), .A2(n3809), .ZN(n3811) );
  NAND2_X1 U4742 ( .A1(n3812), .A2(n3811), .ZN(n4712) );
  NAND2_X1 U4743 ( .A1(n4702), .A2(n4712), .ZN(n4710) );
  INV_X1 U4744 ( .A(n4710), .ZN(n3822) );
  OAI21_X1 U4745 ( .B1(n3815), .B2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n3823), 
        .ZN(n5619) );
  NAND2_X1 U4746 ( .A1(n5619), .A2(n4448), .ZN(n3818) );
  NAND2_X1 U4747 ( .A1(n4453), .A2(EAX_REG_7__SCAN_IN), .ZN(n3817) );
  NAND2_X1 U4748 ( .A1(n4452), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n3816)
         );
  NAND3_X1 U4749 ( .A1(n3818), .A2(n3817), .A3(n3816), .ZN(n3819) );
  INV_X1 U4750 ( .A(n4744), .ZN(n3821) );
  AOI21_X1 U4751 ( .B1(n6716), .B2(n3823), .A(n3853), .ZN(n4795) );
  OR2_X1 U4752 ( .A1(n4795), .A2(n3791), .ZN(n3838) );
  AOI22_X1 U4753 ( .A1(n3110), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n3827) );
  AOI22_X1 U4754 ( .A1(n4388), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3826) );
  AOI22_X1 U4755 ( .A1(n3383), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_12__0__SCAN_IN), .ZN(n3825) );
  AOI22_X1 U4756 ( .A1(n3115), .A2(INSTQUEUE_REG_2__0__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_5__0__SCAN_IN), .ZN(n3824) );
  NAND4_X1 U4757 ( .A1(n3827), .A2(n3826), .A3(n3825), .A4(n3824), .ZN(n3833)
         );
  AOI22_X1 U4758 ( .A1(n4277), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3831) );
  AOI22_X1 U4759 ( .A1(n4341), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3106), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n3830) );
  AOI22_X1 U4760 ( .A1(n3118), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3829) );
  AOI22_X1 U4761 ( .A1(n4434), .A2(INSTQUEUE_REG_0__0__SCAN_IN), .B1(n3108), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n3828) );
  NAND4_X1 U4762 ( .A1(n3831), .A2(n3830), .A3(n3829), .A4(n3828), .ZN(n3832)
         );
  OAI21_X1 U4763 ( .B1(n3833), .B2(n3832), .A(n3944), .ZN(n3836) );
  NAND2_X1 U4764 ( .A1(n4453), .A2(EAX_REG_8__SCAN_IN), .ZN(n3835) );
  NAND2_X1 U4765 ( .A1(n4452), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .ZN(n3834)
         );
  AOI22_X1 U4766 ( .A1(n3110), .A2(INSTQUEUE_REG_6__1__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3842) );
  AOI22_X1 U4767 ( .A1(n3112), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n3841) );
  AOI22_X1 U4768 ( .A1(n3106), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3840) );
  AOI22_X1 U4769 ( .A1(n3109), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3839) );
  NAND4_X1 U4770 ( .A1(n3842), .A2(n3841), .A3(n3840), .A4(n3839), .ZN(n3848)
         );
  AOI22_X1 U4771 ( .A1(n3116), .A2(INSTQUEUE_REG_10__1__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_13__1__SCAN_IN), .ZN(n3846) );
  AOI22_X1 U4772 ( .A1(n3107), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3845) );
  AOI22_X1 U4773 ( .A1(n4427), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3844) );
  AOI22_X1 U4774 ( .A1(n4341), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3843) );
  NAND4_X1 U4775 ( .A1(n3846), .A2(n3845), .A3(n3844), .A4(n3843), .ZN(n3847)
         );
  NOR2_X1 U4776 ( .A1(n3848), .A2(n3847), .ZN(n3852) );
  XNOR2_X1 U4777 ( .A(n3853), .B(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5087) );
  NAND2_X1 U4778 ( .A1(n5087), .A2(n4448), .ZN(n3850) );
  AOI22_X1 U4779 ( .A1(n4453), .A2(EAX_REG_9__SCAN_IN), .B1(n4452), .B2(
        PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n3849) );
  OAI211_X1 U4780 ( .C1(n3852), .C2(n3851), .A(n3850), .B(n3849), .ZN(n4803)
         );
  XOR2_X1 U4781 ( .A(n5603), .B(n3867), .Z(n5606) );
  AOI22_X1 U4782 ( .A1(n3114), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3857) );
  AOI22_X1 U4783 ( .A1(n3121), .A2(INSTQUEUE_REG_15__2__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n3856) );
  AOI22_X1 U4784 ( .A1(n3118), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3855) );
  AOI22_X1 U4785 ( .A1(n4407), .A2(INSTQUEUE_REG_3__2__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_14__2__SCAN_IN), .ZN(n3854) );
  NAND4_X1 U4786 ( .A1(n3857), .A2(n3856), .A3(n3855), .A4(n3854), .ZN(n3863)
         );
  AOI22_X1 U4787 ( .A1(n4341), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3112), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n3861) );
  AOI22_X1 U4788 ( .A1(n4388), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n3860) );
  AOI22_X1 U4789 ( .A1(n3106), .A2(INSTQUEUE_REG_4__2__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3859) );
  AOI22_X1 U4790 ( .A1(n3110), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n3858) );
  NAND4_X1 U4791 ( .A1(n3861), .A2(n3860), .A3(n3859), .A4(n3858), .ZN(n3862)
         );
  OR2_X1 U4792 ( .A1(n3863), .A2(n3862), .ZN(n3864) );
  AOI22_X1 U4793 ( .A1(n3944), .A2(n3864), .B1(n4452), .B2(
        PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n3866) );
  NAND2_X1 U4794 ( .A1(n4453), .A2(EAX_REG_10__SCAN_IN), .ZN(n3865) );
  OAI211_X1 U4795 ( .C1(n5606), .C2(n3791), .A(n3866), .B(n3865), .ZN(n4853)
         );
  XNOR2_X1 U4796 ( .A(n3882), .B(n4885), .ZN(n4865) );
  AOI22_X1 U4797 ( .A1(n4341), .A2(INSTQUEUE_REG_11__3__SCAN_IN), .B1(n3110), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n3871) );
  AOI22_X1 U4798 ( .A1(n3114), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3107), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n3870) );
  AOI22_X1 U4799 ( .A1(n3115), .A2(INSTQUEUE_REG_2__3__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_5__3__SCAN_IN), .ZN(n3869) );
  AOI22_X1 U4800 ( .A1(n4434), .A2(INSTQUEUE_REG_0__3__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_14__3__SCAN_IN), .ZN(n3868) );
  NAND4_X1 U4801 ( .A1(n3871), .A2(n3870), .A3(n3869), .A4(n3868), .ZN(n3877)
         );
  AOI22_X1 U4802 ( .A1(n3116), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_8__3__SCAN_IN), .ZN(n3875) );
  AOI22_X1 U4803 ( .A1(n3383), .A2(INSTQUEUE_REG_15__3__SCAN_IN), .B1(n4427), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n3874) );
  AOI22_X1 U4804 ( .A1(n4277), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3106), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n3873) );
  AOI22_X1 U4805 ( .A1(n3118), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n3872) );
  NAND4_X1 U4806 ( .A1(n3875), .A2(n3874), .A3(n3873), .A4(n3872), .ZN(n3876)
         );
  OAI21_X1 U4807 ( .B1(n3877), .B2(n3876), .A(n3944), .ZN(n3880) );
  NAND2_X1 U4808 ( .A1(n4453), .A2(EAX_REG_11__SCAN_IN), .ZN(n3879) );
  NAND2_X1 U4809 ( .A1(n4452), .A2(PHYADDRPOINTER_REG_11__SCAN_IN), .ZN(n3878)
         );
  NAND3_X1 U4810 ( .A1(n3880), .A2(n3879), .A3(n3878), .ZN(n3881) );
  AOI21_X1 U4811 ( .B1(n4865), .B2(n4448), .A(n3881), .ZN(n4863) );
  XOR2_X1 U4812 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .B(n3897), .Z(n5599) );
  INV_X1 U4813 ( .A(n5599), .ZN(n4894) );
  AOI22_X1 U4814 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n4277), .B1(n3110), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n3886) );
  AOI22_X1 U4815 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n4407), .B1(n4359), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n3885) );
  AOI22_X1 U4816 ( .A1(n3106), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_5__4__SCAN_IN), .ZN(n3884) );
  AOI22_X1 U4817 ( .A1(n3116), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n3883) );
  NAND4_X1 U4818 ( .A1(n3886), .A2(n3885), .A3(n3884), .A4(n3883), .ZN(n3892)
         );
  AOI22_X1 U4819 ( .A1(n3114), .A2(INSTQUEUE_REG_9__4__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_8__4__SCAN_IN), .ZN(n3890) );
  AOI22_X1 U4820 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n3120), .B1(n4434), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n3889) );
  AOI22_X1 U4821 ( .A1(n4341), .A2(INSTQUEUE_REG_11__4__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n3888) );
  AOI22_X1 U4822 ( .A1(n3118), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3108), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n3887) );
  NAND4_X1 U4823 ( .A1(n3890), .A2(n3889), .A3(n3888), .A4(n3887), .ZN(n3891)
         );
  OAI21_X1 U4824 ( .B1(n3892), .B2(n3891), .A(n3944), .ZN(n3895) );
  NAND2_X1 U4825 ( .A1(n4453), .A2(EAX_REG_12__SCAN_IN), .ZN(n3894) );
  NAND2_X1 U4826 ( .A1(n4452), .A2(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n3893)
         );
  NAND3_X1 U4827 ( .A1(n3895), .A2(n3894), .A3(n3893), .ZN(n3896) );
  AOI21_X1 U4828 ( .B1(n4894), .B2(n4448), .A(n3896), .ZN(n4876) );
  NAND2_X1 U4829 ( .A1(n3918), .A2(n3257), .ZN(n3905) );
  NAND2_X1 U4830 ( .A1(n3898), .A2(n6740), .ZN(n3900) );
  INV_X1 U4831 ( .A(n3932), .ZN(n3899) );
  NAND2_X1 U4832 ( .A1(n3900), .A2(n3899), .ZN(n4944) );
  NAND2_X1 U4833 ( .A1(n4944), .A2(n4448), .ZN(n3904) );
  NOR2_X1 U4834 ( .A1(n3901), .A2(n6740), .ZN(n3902) );
  AOI21_X1 U4835 ( .B1(n4453), .B2(EAX_REG_13__SCAN_IN), .A(n3902), .ZN(n3903)
         );
  NAND2_X1 U4836 ( .A1(n3904), .A2(n3903), .ZN(n3919) );
  AOI22_X1 U4837 ( .A1(n4341), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n3909) );
  AOI22_X1 U4838 ( .A1(n4277), .A2(INSTQUEUE_REG_7__5__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_10__5__SCAN_IN), .ZN(n3908) );
  AOI22_X1 U4839 ( .A1(n3106), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n3907) );
  AOI22_X1 U4840 ( .A1(n3110), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_5__5__SCAN_IN), .ZN(n3906) );
  NAND4_X1 U4841 ( .A1(n3909), .A2(n3908), .A3(n3907), .A4(n3906), .ZN(n3915)
         );
  AOI22_X1 U4842 ( .A1(n4407), .A2(INSTQUEUE_REG_3__5__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_13__5__SCAN_IN), .ZN(n3913) );
  AOI22_X1 U4843 ( .A1(n4427), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n3912) );
  AOI22_X1 U4844 ( .A1(n4388), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n3911) );
  AOI22_X1 U4845 ( .A1(n3121), .A2(INSTQUEUE_REG_15__5__SCAN_IN), .B1(n3108), 
        .B2(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n3910) );
  NAND4_X1 U4846 ( .A1(n3913), .A2(n3912), .A3(n3911), .A4(n3910), .ZN(n3914)
         );
  OR2_X1 U4847 ( .A1(n3915), .A2(n3914), .ZN(n3916) );
  AND2_X1 U4848 ( .A1(n3944), .A2(n3916), .ZN(n4911) );
  NAND2_X1 U4849 ( .A1(n4910), .A2(n4911), .ZN(n3921) );
  NAND2_X1 U4850 ( .A1(n3918), .A2(n3917), .ZN(n4862) );
  NOR2_X2 U4851 ( .A1(n4862), .A2(n4876), .ZN(n4875) );
  NAND2_X1 U4852 ( .A1(n4875), .A2(n3919), .ZN(n3920) );
  INV_X1 U4853 ( .A(EAX_REG_14__SCAN_IN), .ZN(n3935) );
  AOI22_X1 U4854 ( .A1(n4427), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n3925) );
  AOI22_X1 U4855 ( .A1(n3106), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n3924) );
  AOI22_X1 U4856 ( .A1(n3110), .A2(INSTQUEUE_REG_6__6__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_5__6__SCAN_IN), .ZN(n3923) );
  AOI22_X1 U4857 ( .A1(n4407), .A2(INSTQUEUE_REG_3__6__SCAN_IN), .B1(n4346), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n3922) );
  NAND4_X1 U4858 ( .A1(n3925), .A2(n3924), .A3(n3923), .A4(n3922), .ZN(n3931)
         );
  AOI22_X1 U4859 ( .A1(n4341), .A2(INSTQUEUE_REG_11__6__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_9__6__SCAN_IN), .ZN(n3929) );
  AOI22_X1 U4860 ( .A1(n3112), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n3928) );
  AOI22_X1 U4861 ( .A1(n3118), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3383), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n3927) );
  AOI22_X1 U4862 ( .A1(n4388), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n3926) );
  NAND4_X1 U4863 ( .A1(n3929), .A2(n3928), .A3(n3927), .A4(n3926), .ZN(n3930)
         );
  OAI21_X1 U4864 ( .B1(n3931), .B2(n3930), .A(n3944), .ZN(n3934) );
  OAI21_X1 U4865 ( .B1(PHYADDRPOINTER_REG_14__SCAN_IN), .B2(n3932), .A(n3952), 
        .ZN(n4960) );
  AOI22_X1 U4866 ( .A1(n4448), .A2(n4960), .B1(n4452), .B2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n3933) );
  OAI211_X1 U4867 ( .C1(n4399), .C2(n3935), .A(n3934), .B(n3933), .ZN(n4922)
         );
  XOR2_X1 U4868 ( .A(n3951), .B(n3952), .Z(n5587) );
  AOI22_X1 U4869 ( .A1(n3111), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_9__7__SCAN_IN), .ZN(n3939) );
  AOI22_X1 U4870 ( .A1(n3107), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_13__7__SCAN_IN), .ZN(n3938) );
  AOI22_X1 U4871 ( .A1(n4427), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n3937) );
  AOI22_X1 U4872 ( .A1(n4341), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n3936) );
  NAND4_X1 U4873 ( .A1(n3939), .A2(n3938), .A3(n3937), .A4(n3936), .ZN(n3946)
         );
  AOI22_X1 U4874 ( .A1(n3110), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n3943) );
  AOI22_X1 U4875 ( .A1(n3106), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n3942) );
  AOI22_X1 U4876 ( .A1(n3120), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3108), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n3941) );
  AOI22_X1 U4877 ( .A1(n4388), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n3940) );
  NAND4_X1 U4878 ( .A1(n3943), .A2(n3942), .A3(n3941), .A4(n3940), .ZN(n3945)
         );
  OAI21_X1 U4879 ( .B1(n3946), .B2(n3945), .A(n3944), .ZN(n3949) );
  NAND2_X1 U4880 ( .A1(n3764), .A2(EAX_REG_15__SCAN_IN), .ZN(n3948) );
  NAND2_X1 U4881 ( .A1(n4452), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .ZN(n3947)
         );
  NAND3_X1 U4882 ( .A1(n3949), .A2(n3948), .A3(n3947), .ZN(n3950) );
  AOI21_X1 U4883 ( .B1(n5271), .B2(n4448), .A(n3950), .ZN(n4955) );
  INV_X1 U4884 ( .A(PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3953) );
  XNOR2_X1 U4885 ( .A(n3982), .B(n3953), .ZN(n5261) );
  OR2_X1 U4886 ( .A1(n5261), .A2(n3791), .ZN(n3968) );
  AOI22_X1 U4887 ( .A1(n4341), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3111), 
        .B2(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n3957) );
  AOI22_X1 U4888 ( .A1(n3116), .A2(INSTQUEUE_REG_11__0__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n3956) );
  AOI22_X1 U4889 ( .A1(n4427), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_1__0__SCAN_IN), .ZN(n3955) );
  AOI22_X1 U4890 ( .A1(n3110), .A2(INSTQUEUE_REG_7__0__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n3954) );
  NAND4_X1 U4891 ( .A1(n3957), .A2(n3956), .A3(n3955), .A4(n3954), .ZN(n3963)
         );
  AOI22_X1 U4892 ( .A1(n3114), .A2(INSTQUEUE_REG_10__0__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_9__0__SCAN_IN), .ZN(n3961) );
  AOI22_X1 U4893 ( .A1(n3106), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n3960) );
  AOI22_X1 U4894 ( .A1(n4407), .A2(INSTQUEUE_REG_4__0__SCAN_IN), .B1(n3108), 
        .B2(INSTQUEUE_REG_15__0__SCAN_IN), .ZN(n3959) );
  AOI22_X1 U4895 ( .A1(n3118), .A2(INSTQUEUE_REG_14__0__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n3958) );
  NAND4_X1 U4896 ( .A1(n3961), .A2(n3960), .A3(n3959), .A4(n3958), .ZN(n3962)
         );
  NOR2_X1 U4897 ( .A1(n3963), .A2(n3962), .ZN(n3965) );
  AOI22_X1 U4898 ( .A1(n3764), .A2(EAX_REG_16__SCAN_IN), .B1(n4452), .B2(
        PHYADDRPOINTER_REG_16__SCAN_IN), .ZN(n3964) );
  OAI21_X1 U4899 ( .B1(n4422), .B2(n3965), .A(n3964), .ZN(n3966) );
  INV_X1 U4900 ( .A(n3966), .ZN(n3967) );
  AOI22_X1 U4901 ( .A1(n4277), .A2(INSTQUEUE_REG_8__1__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n3972) );
  AOI22_X1 U4902 ( .A1(n3116), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n3971) );
  AOI22_X1 U4903 ( .A1(n4341), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3106), 
        .B2(INSTQUEUE_REG_5__1__SCAN_IN), .ZN(n3970) );
  AOI22_X1 U4904 ( .A1(n3118), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n4346), 
        .B2(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n3969) );
  NAND4_X1 U4905 ( .A1(n3972), .A2(n3971), .A3(n3970), .A4(n3969), .ZN(n3978)
         );
  AOI22_X1 U4906 ( .A1(n3107), .A2(INSTQUEUE_REG_4__1__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n3976) );
  AOI22_X1 U4907 ( .A1(n4427), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n3975) );
  AOI22_X1 U4908 ( .A1(n3115), .A2(INSTQUEUE_REG_3__1__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n3974) );
  AOI22_X1 U4909 ( .A1(n3110), .A2(INSTQUEUE_REG_7__1__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_2__1__SCAN_IN), .ZN(n3973) );
  NAND4_X1 U4910 ( .A1(n3976), .A2(n3975), .A3(n3974), .A4(n3973), .ZN(n3977)
         );
  NOR2_X1 U4911 ( .A1(n3978), .A2(n3977), .ZN(n3979) );
  OR2_X1 U4912 ( .A1(n4422), .A2(n3979), .ZN(n3986) );
  NAND2_X1 U4913 ( .A1(n6511), .A2(PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n3980)
         );
  NAND2_X1 U4914 ( .A1(n3791), .A2(n3980), .ZN(n3981) );
  AOI21_X1 U4915 ( .B1(n3764), .B2(EAX_REG_17__SCAN_IN), .A(n3981), .ZN(n3985)
         );
  OAI21_X1 U4916 ( .B1(PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n3983), .A(n4000), 
        .ZN(n5575) );
  NOR2_X1 U4917 ( .A1(n5575), .A2(n3791), .ZN(n3984) );
  AOI21_X1 U4918 ( .B1(n3986), .B2(n3985), .A(n3984), .ZN(n4984) );
  NAND2_X1 U4919 ( .A1(n4965), .A2(n4984), .ZN(n4983) );
  AOI22_X1 U4920 ( .A1(n3112), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_10__2__SCAN_IN), .ZN(n3990) );
  AOI22_X1 U4921 ( .A1(n3116), .A2(INSTQUEUE_REG_11__2__SCAN_IN), .B1(n3107), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n3989) );
  AOI22_X1 U4922 ( .A1(n4427), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_1__2__SCAN_IN), .ZN(n3988) );
  AOI22_X1 U4923 ( .A1(n3106), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_6__2__SCAN_IN), .ZN(n3987) );
  NAND4_X1 U4924 ( .A1(n3990), .A2(n3989), .A3(n3988), .A4(n3987), .ZN(n3996)
         );
  AOI22_X1 U4925 ( .A1(n4341), .A2(INSTQUEUE_REG_12__2__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_9__2__SCAN_IN), .ZN(n3994) );
  AOI22_X1 U4926 ( .A1(n3110), .A2(INSTQUEUE_REG_7__2__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n3993) );
  AOI22_X1 U4927 ( .A1(n3383), .A2(INSTQUEUE_REG_0__2__SCAN_IN), .B1(n3108), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n3992) );
  AOI22_X1 U4928 ( .A1(n3118), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n3991) );
  NAND4_X1 U4929 ( .A1(n3994), .A2(n3993), .A3(n3992), .A4(n3991), .ZN(n3995)
         );
  NOR2_X1 U4930 ( .A1(n3996), .A2(n3995), .ZN(n3999) );
  OAI21_X1 U4931 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6705), .A(n3791), .ZN(
        n3997) );
  AOI21_X1 U4932 ( .B1(n3764), .B2(EAX_REG_18__SCAN_IN), .A(n3997), .ZN(n3998)
         );
  OAI21_X1 U4933 ( .B1(n4422), .B2(n3999), .A(n3998), .ZN(n4002) );
  AOI21_X1 U4934 ( .B1(n6705), .B2(n4000), .A(n4017), .ZN(n5251) );
  NAND2_X1 U4935 ( .A1(n5251), .A2(n4448), .ZN(n4001) );
  AOI22_X1 U4936 ( .A1(n4341), .A2(INSTQUEUE_REG_12__3__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_10__3__SCAN_IN), .ZN(n4006) );
  AOI22_X1 U4937 ( .A1(n3111), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4005) );
  AOI22_X1 U4938 ( .A1(n3110), .A2(INSTQUEUE_REG_7__3__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_6__3__SCAN_IN), .ZN(n4004) );
  AOI22_X1 U4939 ( .A1(n4388), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n4346), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4003) );
  NAND4_X1 U4940 ( .A1(n4006), .A2(n4005), .A3(n4004), .A4(n4003), .ZN(n4012)
         );
  AOI22_X1 U4941 ( .A1(n4407), .A2(INSTQUEUE_REG_4__3__SCAN_IN), .B1(n3121), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4010) );
  AOI22_X1 U4942 ( .A1(n4427), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_1__3__SCAN_IN), .ZN(n4009) );
  AOI22_X1 U4943 ( .A1(n3106), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4008) );
  AOI22_X1 U4944 ( .A1(n3118), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4007) );
  NAND4_X1 U4945 ( .A1(n4010), .A2(n4009), .A3(n4008), .A4(n4007), .ZN(n4011)
         );
  NOR2_X1 U4946 ( .A1(n4012), .A2(n4011), .ZN(n4016) );
  NAND2_X1 U4947 ( .A1(n6511), .A2(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n4013)
         );
  NAND2_X1 U4948 ( .A1(n3791), .A2(n4013), .ZN(n4014) );
  AOI21_X1 U4949 ( .B1(n3764), .B2(EAX_REG_19__SCAN_IN), .A(n4014), .ZN(n4015)
         );
  OAI21_X1 U4950 ( .B1(n4422), .B2(n4016), .A(n4015), .ZN(n4019) );
  OAI21_X1 U4951 ( .B1(PHYADDRPOINTER_REG_19__SCAN_IN), .B2(n4017), .A(n4033), 
        .ZN(n5499) );
  OR2_X1 U4952 ( .A1(n3791), .A2(n5499), .ZN(n4018) );
  NAND2_X1 U4953 ( .A1(n4019), .A2(n4018), .ZN(n5149) );
  AOI22_X1 U4954 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n4277), .B1(n3114), 
        .B2(INSTQUEUE_REG_10__4__SCAN_IN), .ZN(n4023) );
  AOI22_X1 U4955 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n4388), .B1(n3118), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4022) );
  AOI22_X1 U4956 ( .A1(n3106), .A2(INSTQUEUE_REG_5__4__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4021) );
  AOI22_X1 U4957 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n4427), .B1(n4346), 
        .B2(INSTQUEUE_REG_15__4__SCAN_IN), .ZN(n4020) );
  NAND4_X1 U4958 ( .A1(n4023), .A2(n4022), .A3(n4021), .A4(n4020), .ZN(n4029)
         );
  AOI22_X1 U4959 ( .A1(n4341), .A2(INSTQUEUE_REG_12__4__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4027) );
  AOI22_X1 U4960 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n3383), .B1(n4434), 
        .B2(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n4026) );
  AOI22_X1 U4961 ( .A1(n3110), .A2(INSTQUEUE_REG_7__4__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_6__4__SCAN_IN), .ZN(n4025) );
  AOI22_X1 U4962 ( .A1(n4407), .A2(INSTQUEUE_REG_4__4__SCAN_IN), .B1(n3102), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4024) );
  NAND4_X1 U4963 ( .A1(n4027), .A2(n4026), .A3(n4025), .A4(n4024), .ZN(n4028)
         );
  NOR2_X1 U4964 ( .A1(n4029), .A2(n4028), .ZN(n4032) );
  INV_X1 U4965 ( .A(PHYADDRPOINTER_REG_20__SCAN_IN), .ZN(n6690) );
  OAI21_X1 U4966 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6690), .A(n3791), .ZN(
        n4030) );
  AOI21_X1 U4967 ( .B1(n3764), .B2(EAX_REG_20__SCAN_IN), .A(n4030), .ZN(n4031)
         );
  OAI21_X1 U4968 ( .B1(n4422), .B2(n4032), .A(n4031), .ZN(n4037) );
  NOR2_X1 U4969 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(n4034), .ZN(n4035)
         );
  NOR2_X1 U4970 ( .A1(n4051), .A2(n4035), .ZN(n5242) );
  NAND2_X1 U4971 ( .A1(n5242), .A2(n4448), .ZN(n4036) );
  AOI22_X1 U4972 ( .A1(n3111), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3110), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4041) );
  AOI22_X1 U4973 ( .A1(n3118), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4040) );
  AOI22_X1 U4974 ( .A1(n4435), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n4039) );
  AOI22_X1 U4975 ( .A1(n3116), .A2(INSTQUEUE_REG_11__5__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4038) );
  NAND4_X1 U4976 ( .A1(n4041), .A2(n4040), .A3(n4039), .A4(n4038), .ZN(n4047)
         );
  AOI22_X1 U4977 ( .A1(n3114), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_9__5__SCAN_IN), .ZN(n4045) );
  AOI22_X1 U4978 ( .A1(n4427), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n4044) );
  AOI22_X1 U4979 ( .A1(n4341), .A2(INSTQUEUE_REG_12__5__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4043) );
  AOI22_X1 U4980 ( .A1(n4407), .A2(INSTQUEUE_REG_4__5__SCAN_IN), .B1(n3108), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4042) );
  NAND4_X1 U4981 ( .A1(n4045), .A2(n4044), .A3(n4043), .A4(n4042), .ZN(n4046)
         );
  NOR2_X1 U4982 ( .A1(n4047), .A2(n4046), .ZN(n4048) );
  OR2_X1 U4983 ( .A1(n4422), .A2(n4048), .ZN(n4054) );
  NAND2_X1 U4984 ( .A1(n6511), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n4049)
         );
  NAND2_X1 U4985 ( .A1(n3791), .A2(n4049), .ZN(n4050) );
  AOI21_X1 U4986 ( .B1(n4453), .B2(EAX_REG_21__SCAN_IN), .A(n4050), .ZN(n4053)
         );
  OAI21_X1 U4987 ( .B1(n4051), .B2(PHYADDRPOINTER_REG_21__SCAN_IN), .A(n4293), 
        .ZN(n5450) );
  NOR2_X1 U4988 ( .A1(n5450), .A2(n3791), .ZN(n4052) );
  AOI21_X1 U4989 ( .B1(n4054), .B2(n4053), .A(n4052), .ZN(n5232) );
  NAND2_X1 U4990 ( .A1(n5059), .A2(n5232), .ZN(n4070) );
  INV_X1 U4991 ( .A(n4070), .ZN(n5233) );
  AOI22_X1 U4992 ( .A1(n4341), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4058) );
  AOI22_X1 U4993 ( .A1(n3112), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4057) );
  AOI22_X1 U4994 ( .A1(n3106), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4056) );
  AOI22_X1 U4995 ( .A1(n3110), .A2(INSTQUEUE_REG_7__6__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4055) );
  NAND4_X1 U4996 ( .A1(n4058), .A2(n4057), .A3(n4056), .A4(n4055), .ZN(n4064)
         );
  AOI22_X1 U4997 ( .A1(n4407), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_14__6__SCAN_IN), .ZN(n4062) );
  AOI22_X1 U4998 ( .A1(n4427), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_1__6__SCAN_IN), .ZN(n4061) );
  AOI22_X1 U4999 ( .A1(n4388), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4060) );
  AOI22_X1 U5000 ( .A1(n3120), .A2(INSTQUEUE_REG_0__6__SCAN_IN), .B1(n3108), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4059) );
  NAND4_X1 U5001 ( .A1(n4062), .A2(n4061), .A3(n4060), .A4(n4059), .ZN(n4063)
         );
  NOR2_X1 U5002 ( .A1(n4064), .A2(n4063), .ZN(n4067) );
  AOI21_X1 U5003 ( .B1(n4292), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4065) );
  AOI21_X1 U5004 ( .B1(n4453), .B2(EAX_REG_22__SCAN_IN), .A(n4065), .ZN(n4066)
         );
  OAI21_X1 U5005 ( .B1(n4422), .B2(n4067), .A(n4066), .ZN(n4069) );
  XNOR2_X1 U5006 ( .A(n4293), .B(PHYADDRPOINTER_REG_22__SCAN_IN), .ZN(n5053)
         );
  NAND2_X1 U5007 ( .A1(n5053), .A2(n4448), .ZN(n4068) );
  OAI21_X1 U5008 ( .B1(n5233), .B2(n3251), .A(n4299), .ZN(n5178) );
  NAND3_X1 U5009 ( .A1(n6521), .A2(STATEBS16_REG_SCAN_IN), .A3(
        STATE2_REG_1__SCAN_IN), .ZN(n6530) );
  INV_X1 U5010 ( .A(n6530), .ZN(n4071) );
  NAND2_X1 U5011 ( .A1(n6410), .A2(n4076), .ZN(n6627) );
  NAND2_X1 U5012 ( .A1(n6627), .A2(n6521), .ZN(n4072) );
  NAND2_X1 U5013 ( .A1(n6521), .A2(STATE2_REG_2__SCAN_IN), .ZN(n4074) );
  NAND2_X1 U5014 ( .A1(n6286), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4073) );
  NAND2_X1 U5015 ( .A1(n4074), .A2(n4073), .ZN(n5776) );
  INV_X1 U5016 ( .A(n5776), .ZN(n4075) );
  AND2_X1 U5017 ( .A1(n5832), .A2(REIP_REG_22__SCAN_IN), .ZN(n5339) );
  NOR2_X1 U5018 ( .A1(n5248), .A2(n4292), .ZN(n4077) );
  AOI211_X1 U5019 ( .C1(n5250), .C2(n5053), .A(n5339), .B(n4077), .ZN(n4078)
         );
  NAND2_X1 U5020 ( .A1(n4081), .A2(n4080), .ZN(U2964) );
  NOR2_X1 U5021 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4082) );
  NOR2_X1 U5022 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5336) );
  AND2_X1 U5023 ( .A1(INSTADDRPOINTER_REG_19__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_20__SCAN_IN), .ZN(n5360) );
  AND2_X1 U5024 ( .A1(INSTADDRPOINTER_REG_21__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5335) );
  AND2_X1 U5025 ( .A1(INSTADDRPOINTER_REG_24__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n4245) );
  AND3_X1 U5026 ( .A1(n5360), .A2(n5335), .A3(n4245), .ZN(n4083) );
  XNOR2_X1 U5027 ( .A(n5245), .B(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5313)
         );
  INV_X1 U5028 ( .A(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4192) );
  INV_X1 U5029 ( .A(INSTADDRPOINTER_REG_26__SCAN_IN), .ZN(n5302) );
  NOR2_X1 U5030 ( .A1(n3680), .A2(n5302), .ZN(n5205) );
  INV_X1 U5031 ( .A(n5198), .ZN(n5182) );
  OR2_X1 U5032 ( .A1(n5245), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n4085)
         );
  OAI22_X1 U5033 ( .A1(n5182), .A2(n4487), .B1(INSTADDRPOINTER_REG_27__SCAN_IN), .B2(n5302), .ZN(n4087) );
  XNOR2_X1 U5034 ( .A(n4087), .B(n4086), .ZN(n5197) );
  NOR2_X1 U5035 ( .A1(n6475), .A2(n3408), .ZN(n4226) );
  INV_X1 U5036 ( .A(n4226), .ZN(n4105) );
  INV_X1 U5037 ( .A(n4088), .ZN(n4089) );
  NAND2_X1 U5038 ( .A1(n4089), .A2(n6541), .ZN(n6539) );
  NAND2_X1 U5039 ( .A1(n3397), .A2(n6539), .ZN(n4098) );
  AND3_X1 U5040 ( .A1(n4092), .A2(n4091), .A3(n4090), .ZN(n4094) );
  OAI21_X1 U5041 ( .B1(n4095), .B2(n4094), .A(n4093), .ZN(n4521) );
  INV_X1 U5042 ( .A(n4521), .ZN(n4096) );
  NOR2_X1 U5043 ( .A1(n4096), .A2(READY_N), .ZN(n4558) );
  NAND3_X1 U5044 ( .A1(n4098), .A2(n4558), .A3(n4097), .ZN(n4104) );
  NAND2_X1 U5045 ( .A1(n4604), .A2(n3407), .ZN(n4099) );
  NAND2_X1 U5046 ( .A1(n6630), .A2(n4099), .ZN(n4100) );
  NAND2_X1 U5047 ( .A1(n3445), .A2(n4100), .ZN(n4217) );
  INV_X1 U5048 ( .A(n4217), .ZN(n4101) );
  OR2_X1 U5049 ( .A1(n4116), .A2(n4101), .ZN(n4103) );
  NAND2_X1 U5050 ( .A1(n4103), .A2(n4102), .ZN(n4567) );
  OAI211_X1 U5051 ( .C1(n6513), .C2(n4105), .A(n4104), .B(n4567), .ZN(n4106)
         );
  NAND2_X1 U5052 ( .A1(n4106), .A2(n6518), .ZN(n4113) );
  NAND2_X1 U5053 ( .A1(n3408), .A2(n6539), .ZN(n4474) );
  NAND3_X1 U5054 ( .A1(n4107), .A2(n4474), .A3(n6628), .ZN(n4109) );
  NAND3_X1 U5055 ( .A1(n4109), .A2(n3407), .A3(n4108), .ZN(n4110) );
  NAND2_X1 U5056 ( .A1(n4110), .A2(n3409), .ZN(n4111) );
  INV_X1 U5057 ( .A(n4208), .ZN(n4115) );
  AOI22_X1 U5058 ( .A1(n4115), .A2(n3398), .B1(n4107), .B2(n4561), .ZN(n4117)
         );
  NOR2_X1 U5059 ( .A1(n4116), .A2(n3717), .ZN(n4557) );
  INV_X1 U5060 ( .A(n4557), .ZN(n4652) );
  AND4_X1 U5061 ( .A1(n4114), .A2(n4117), .A3(n4652), .A4(n6496), .ZN(n4118)
         );
  INV_X1 U5062 ( .A(n4119), .ZN(n4122) );
  OR2_X1 U5063 ( .A1(n4468), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .ZN(n4120)
         );
  NAND2_X1 U5064 ( .A1(n4121), .A2(n4120), .ZN(n4124) );
  INV_X1 U5065 ( .A(EBX_REG_0__SCAN_IN), .ZN(n4123) );
  OAI22_X1 U5066 ( .A1(n4204), .A2(n4123), .B1(n4159), .B2(EBX_REG_0__SCAN_IN), 
        .ZN(n4584) );
  XNOR2_X1 U5067 ( .A(n4124), .B(n4584), .ZN(n5675) );
  AOI21_X1 U5068 ( .B1(n5675), .B2(n4561), .A(n4124), .ZN(n4825) );
  INV_X1 U5069 ( .A(EBX_REG_2__SCAN_IN), .ZN(n5705) );
  NAND2_X1 U5070 ( .A1(n4202), .A2(n5705), .ZN(n4127) );
  NAND2_X1 U5071 ( .A1(n4159), .A2(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n4125)
         );
  OAI211_X1 U5072 ( .C1(n4178), .C2(EBX_REG_2__SCAN_IN), .A(n4204), .B(n4125), 
        .ZN(n4126) );
  AND2_X1 U5073 ( .A1(n4127), .A2(n4126), .ZN(n4824) );
  NAND2_X1 U5074 ( .A1(n4825), .A2(n4824), .ZN(n4826) );
  MUX2_X1 U5075 ( .A(n4199), .B(n4204), .S(EBX_REG_3__SCAN_IN), .Z(n4130) );
  INV_X1 U5076 ( .A(n4204), .ZN(n4128) );
  NAND2_X1 U5077 ( .A1(n4178), .A2(INSTADDRPOINTER_REG_3__SCAN_IN), .ZN(n4129)
         );
  AND3_X1 U5078 ( .A1(n4130), .A2(n4180), .A3(n4129), .ZN(n4646) );
  MUX2_X1 U5079 ( .A(n4197), .B(n4159), .S(EBX_REG_4__SCAN_IN), .Z(n4131) );
  OAI21_X1 U5080 ( .B1(INSTADDRPOINTER_REG_4__SCAN_IN), .B2(n4468), .A(n4131), 
        .ZN(n4697) );
  OR2_X1 U5081 ( .A1(n4199), .A2(EBX_REG_5__SCAN_IN), .ZN(n4137) );
  NAND2_X1 U5082 ( .A1(n4204), .A2(n4132), .ZN(n4135) );
  INV_X1 U5083 ( .A(EBX_REG_5__SCAN_IN), .ZN(n4133) );
  NAND2_X1 U5084 ( .A1(n4561), .A2(n4133), .ZN(n4134) );
  NAND3_X1 U5085 ( .A1(n4135), .A2(n4159), .A3(n4134), .ZN(n4136) );
  NAND2_X1 U5086 ( .A1(n4137), .A2(n4136), .ZN(n4705) );
  MUX2_X1 U5087 ( .A(n4197), .B(n4159), .S(EBX_REG_6__SCAN_IN), .Z(n4138) );
  OAI21_X1 U5088 ( .B1(n4468), .B2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n4138), 
        .ZN(n4715) );
  OR2_X1 U5089 ( .A1(n4199), .A2(EBX_REG_7__SCAN_IN), .ZN(n4143) );
  NAND2_X1 U5090 ( .A1(n4204), .A2(n4139), .ZN(n4141) );
  INV_X1 U5091 ( .A(EBX_REG_7__SCAN_IN), .ZN(n5625) );
  NAND2_X1 U5092 ( .A1(n4561), .A2(n5625), .ZN(n4140) );
  NAND3_X1 U5093 ( .A1(n4141), .A2(n4159), .A3(n4140), .ZN(n4142) );
  MUX2_X1 U5094 ( .A(n4197), .B(n4159), .S(EBX_REG_8__SCAN_IN), .Z(n4144) );
  OAI21_X1 U5095 ( .B1(n4468), .B2(INSTADDRPOINTER_REG_8__SCAN_IN), .A(n4144), 
        .ZN(n4145) );
  INV_X1 U5096 ( .A(n4145), .ZN(n4776) );
  MUX2_X1 U5097 ( .A(n4199), .B(n4204), .S(EBX_REG_9__SCAN_IN), .Z(n4148) );
  NAND2_X1 U5098 ( .A1(n4178), .A2(INSTADDRPOINTER_REG_9__SCAN_IN), .ZN(n4146)
         );
  AND2_X1 U5099 ( .A1(n4180), .A2(n4146), .ZN(n4147) );
  NAND2_X1 U5100 ( .A1(n4148), .A2(n4147), .ZN(n4846) );
  INV_X1 U5101 ( .A(EBX_REG_10__SCAN_IN), .ZN(n5702) );
  NAND2_X1 U5102 ( .A1(n4202), .A2(n5702), .ZN(n4151) );
  NAND2_X1 U5103 ( .A1(n4159), .A2(INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4149) );
  OAI211_X1 U5104 ( .C1(n4178), .C2(EBX_REG_10__SCAN_IN), .A(n4204), .B(n4149), 
        .ZN(n4150) );
  AND2_X1 U5105 ( .A1(n4151), .A2(n4150), .ZN(n4845) );
  MUX2_X1 U5106 ( .A(n4199), .B(n4204), .S(EBX_REG_11__SCAN_IN), .Z(n4154) );
  NAND2_X1 U5107 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(n4178), .ZN(n4153) );
  MUX2_X1 U5108 ( .A(n4197), .B(n4159), .S(EBX_REG_12__SCAN_IN), .Z(n4155) );
  OAI21_X1 U5109 ( .B1(INSTADDRPOINTER_REG_12__SCAN_IN), .B2(n4468), .A(n4155), 
        .ZN(n4878) );
  MUX2_X1 U5110 ( .A(n4199), .B(n4204), .S(EBX_REG_13__SCAN_IN), .Z(n4158) );
  NAND2_X1 U5111 ( .A1(INSTADDRPOINTER_REG_13__SCAN_IN), .A2(n4178), .ZN(n4156) );
  AND2_X1 U5112 ( .A1(n4180), .A2(n4156), .ZN(n4157) );
  NAND2_X1 U5113 ( .A1(n4158), .A2(n4157), .ZN(n4928) );
  INV_X1 U5114 ( .A(EBX_REG_14__SCAN_IN), .ZN(n6896) );
  NAND2_X1 U5115 ( .A1(n4202), .A2(n6896), .ZN(n4162) );
  NAND2_X1 U5116 ( .A1(n4159), .A2(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4160) );
  OAI211_X1 U5117 ( .C1(n4178), .C2(EBX_REG_14__SCAN_IN), .A(n4204), .B(n4160), 
        .ZN(n4161) );
  NAND2_X1 U5118 ( .A1(n4928), .A2(n4927), .ZN(n4163) );
  MUX2_X1 U5119 ( .A(n4199), .B(n4204), .S(EBX_REG_15__SCAN_IN), .Z(n4166) );
  NAND2_X1 U5120 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n4178), .ZN(n4164) );
  AND2_X1 U5121 ( .A1(n4180), .A2(n4164), .ZN(n4165) );
  NAND2_X1 U5122 ( .A1(n4166), .A2(n4165), .ZN(n5158) );
  NAND2_X1 U5123 ( .A1(n5159), .A2(n5158), .ZN(n5161) );
  NAND2_X1 U5124 ( .A1(n4159), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n4167) );
  OAI211_X1 U5125 ( .C1(n4178), .C2(EBX_REG_16__SCAN_IN), .A(n4204), .B(n4167), 
        .ZN(n4168) );
  OAI21_X1 U5126 ( .B1(n4197), .B2(EBX_REG_16__SCAN_IN), .A(n4168), .ZN(n4967)
         );
  MUX2_X1 U5127 ( .A(n4199), .B(n4204), .S(EBX_REG_17__SCAN_IN), .Z(n4170) );
  NAND2_X1 U5128 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n4178), .ZN(n4169) );
  MUX2_X1 U5129 ( .A(n4197), .B(n4159), .S(EBX_REG_19__SCAN_IN), .Z(n4171) );
  OAI21_X1 U5130 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n4468), .A(n4171), 
        .ZN(n5151) );
  INV_X1 U5131 ( .A(n5151), .ZN(n4172) );
  INV_X1 U5132 ( .A(n4468), .ZN(n4585) );
  NOR2_X1 U5133 ( .A1(n4178), .A2(EBX_REG_20__SCAN_IN), .ZN(n4173) );
  AOI21_X1 U5134 ( .B1(n4585), .B2(n5364), .A(n4173), .ZN(n5064) );
  OR2_X1 U5135 ( .A1(n4468), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n4174)
         );
  INV_X1 U5136 ( .A(EBX_REG_18__SCAN_IN), .ZN(n5157) );
  NAND2_X1 U5137 ( .A1(n4561), .A2(n5157), .ZN(n5074) );
  NAND2_X1 U5138 ( .A1(n4174), .A2(n5074), .ZN(n5075) );
  NOR2_X1 U5139 ( .A1(n5064), .A2(n5075), .ZN(n4176) );
  MUX2_X1 U5140 ( .A(n5075), .B(EBX_REG_20__SCAN_IN), .S(n4122), .Z(n4175) );
  NOR2_X1 U5141 ( .A1(n4176), .A2(n4175), .ZN(n4177) );
  MUX2_X1 U5142 ( .A(n4199), .B(n4204), .S(EBX_REG_21__SCAN_IN), .Z(n4182) );
  NAND2_X1 U5143 ( .A1(n4178), .A2(INSTADDRPOINTER_REG_21__SCAN_IN), .ZN(n4179) );
  AND2_X1 U5144 ( .A1(n4180), .A2(n4179), .ZN(n4181) );
  NAND2_X1 U5145 ( .A1(n4182), .A2(n4181), .ZN(n5344) );
  INV_X1 U5146 ( .A(EBX_REG_22__SCAN_IN), .ZN(n5049) );
  NAND2_X1 U5147 ( .A1(n4202), .A2(n5049), .ZN(n4185) );
  NAND2_X1 U5148 ( .A1(n4159), .A2(INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n4183) );
  OAI211_X1 U5149 ( .C1(n4178), .C2(EBX_REG_22__SCAN_IN), .A(n4204), .B(n4183), 
        .ZN(n4184) );
  NAND2_X1 U5150 ( .A1(n5344), .A2(n5051), .ZN(n4186) );
  NAND2_X1 U5151 ( .A1(INSTADDRPOINTER_REG_23__SCAN_IN), .A2(n4178), .ZN(n4188) );
  MUX2_X1 U5152 ( .A(n4199), .B(n4204), .S(EBX_REG_23__SCAN_IN), .Z(n4187) );
  AND2_X1 U5153 ( .A1(n4188), .A2(n4187), .ZN(n5140) );
  INV_X1 U5154 ( .A(EBX_REG_24__SCAN_IN), .ZN(n5138) );
  NAND2_X1 U5155 ( .A1(n4202), .A2(n5138), .ZN(n4191) );
  NAND2_X1 U5156 ( .A1(n4159), .A2(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n4189) );
  OAI211_X1 U5157 ( .C1(n4178), .C2(EBX_REG_24__SCAN_IN), .A(n4204), .B(n4189), 
        .ZN(n4190) );
  OR2_X1 U5158 ( .A1(n4199), .A2(EBX_REG_25__SCAN_IN), .ZN(n4196) );
  NAND2_X1 U5159 ( .A1(n4204), .A2(n4192), .ZN(n4194) );
  INV_X1 U5160 ( .A(EBX_REG_25__SCAN_IN), .ZN(n5129) );
  NAND2_X1 U5161 ( .A1(n4561), .A2(n5129), .ZN(n4193) );
  NAND3_X1 U5162 ( .A1(n4194), .A2(n4159), .A3(n4193), .ZN(n4195) );
  NAND2_X1 U5163 ( .A1(n4196), .A2(n4195), .ZN(n5127) );
  MUX2_X1 U5164 ( .A(n4197), .B(n4159), .S(EBX_REG_26__SCAN_IN), .Z(n4198) );
  OAI21_X1 U5165 ( .B1(INSTADDRPOINTER_REG_26__SCAN_IN), .B2(n4468), .A(n4198), 
        .ZN(n5120) );
  NAND2_X1 U5166 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(n4178), .ZN(n4201) );
  MUX2_X1 U5167 ( .A(n4199), .B(n4204), .S(EBX_REG_27__SCAN_IN), .Z(n4200) );
  AND2_X1 U5168 ( .A1(n4201), .A2(n4200), .ZN(n5111) );
  INV_X1 U5169 ( .A(EBX_REG_28__SCAN_IN), .ZN(n6885) );
  NAND2_X1 U5170 ( .A1(n4202), .A2(n6885), .ZN(n4206) );
  NAND2_X1 U5171 ( .A1(n4159), .A2(INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4203) );
  OAI211_X1 U5172 ( .C1(n4178), .C2(EBX_REG_28__SCAN_IN), .A(n4204), .B(n4203), 
        .ZN(n4205) );
  OAI21_X1 U5173 ( .B1(n5113), .B2(n4207), .A(n5022), .ZN(n5107) );
  INV_X1 U5174 ( .A(n5107), .ZN(n4211) );
  NAND2_X1 U5175 ( .A1(n4107), .A2(n3428), .ZN(n6507) );
  OAI21_X1 U5176 ( .B1(n4208), .B2(n3398), .A(n6507), .ZN(n4209) );
  INV_X1 U5177 ( .A(n4209), .ZN(n4210) );
  NAND2_X1 U5178 ( .A1(n4211), .A2(n5834), .ZN(n4251) );
  NAND2_X1 U5179 ( .A1(n3098), .A2(n3397), .ZN(n6478) );
  INV_X1 U5180 ( .A(n4212), .ZN(n4214) );
  AND2_X1 U5181 ( .A1(n4214), .A2(n4213), .ZN(n4218) );
  NOR2_X1 U5182 ( .A1(n4507), .A2(n4097), .ZN(n4565) );
  OAI21_X1 U5183 ( .B1(n4565), .B2(n4468), .A(n4215), .ZN(n4216) );
  NAND4_X1 U5184 ( .A1(n4219), .A2(n4218), .A3(n4217), .A4(n4216), .ZN(n4546)
         );
  NAND2_X1 U5185 ( .A1(n4495), .A2(n3438), .ZN(n4221) );
  OR3_X1 U5186 ( .A1(n6475), .A2(n4097), .A3(n4221), .ZN(n4665) );
  OAI21_X1 U5187 ( .B1(n4220), .B2(n3434), .A(n4665), .ZN(n4222) );
  NOR2_X1 U5188 ( .A1(n4546), .A2(n4222), .ZN(n4227) );
  INV_X1 U5189 ( .A(n4544), .ZN(n4223) );
  NAND2_X1 U5190 ( .A1(n4223), .A2(n3438), .ZN(n4224) );
  AND2_X1 U5191 ( .A1(n4227), .A2(n4224), .ZN(n4225) );
  NAND2_X1 U5192 ( .A1(n4227), .A2(n4226), .ZN(n4653) );
  INV_X1 U5193 ( .A(INSTADDRPOINTER_REG_0__SCAN_IN), .ZN(n6605) );
  NAND2_X1 U5194 ( .A1(n4903), .A2(n5525), .ZN(n5529) );
  NAND2_X1 U5195 ( .A1(n6605), .A2(n5529), .ZN(n4586) );
  NAND2_X1 U5196 ( .A1(n4228), .A2(n5811), .ZN(n4587) );
  NAND2_X1 U5197 ( .A1(n4898), .A2(n5356), .ZN(n4231) );
  INV_X1 U5198 ( .A(n4244), .ZN(n4229) );
  NAND2_X1 U5199 ( .A1(n4229), .A2(n5360), .ZN(n4230) );
  NAND2_X1 U5200 ( .A1(n4231), .A2(n4230), .ZN(n4237) );
  INV_X1 U5201 ( .A(INSTADDRPOINTER_REG_2__SCAN_IN), .ZN(n5840) );
  NOR2_X1 U5202 ( .A1(n5840), .A2(n5858), .ZN(n5836) );
  NOR2_X1 U5203 ( .A1(n3615), .A2(n3627), .ZN(n5818) );
  AND4_X1 U5204 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .A3(n5836), .A4(n5818), .ZN(n4734) );
  INV_X1 U5205 ( .A(INSTADDRPOINTER_REG_8__SCAN_IN), .ZN(n6759) );
  NOR2_X1 U5206 ( .A1(n4139), .A2(n6759), .ZN(n4841) );
  INV_X1 U5207 ( .A(n4841), .ZN(n5799) );
  NAND2_X1 U5208 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_10__SCAN_IN), .ZN(n4843) );
  NOR2_X1 U5209 ( .A1(n5799), .A2(n4843), .ZN(n4235) );
  NAND2_X1 U5210 ( .A1(n4734), .A2(n4235), .ZN(n4900) );
  NAND2_X1 U5211 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n6665) );
  NAND2_X1 U5212 ( .A1(INSTADDRPOINTER_REG_11__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n6661) );
  NOR2_X1 U5213 ( .A1(n5545), .A2(n6661), .ZN(n5535) );
  NAND2_X1 U5214 ( .A1(INSTADDRPOINTER_REG_14__SCAN_IN), .A2(n5535), .ZN(n5517) );
  OR2_X1 U5215 ( .A1(n6665), .A2(n5517), .ZN(n4243) );
  NOR2_X1 U5216 ( .A1(n4900), .A2(n4243), .ZN(n4232) );
  OR2_X1 U5217 ( .A1(n4898), .A2(n4232), .ZN(n5358) );
  NAND2_X1 U5218 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_6__SCAN_IN), .ZN(n4234) );
  OAI21_X1 U5219 ( .B1(n5858), .B2(n6605), .A(n5840), .ZN(n5820) );
  INV_X1 U5220 ( .A(n5820), .ZN(n5837) );
  INV_X1 U5221 ( .A(n5818), .ZN(n4233) );
  NOR2_X1 U5222 ( .A1(n5837), .A2(n4233), .ZN(n4739) );
  NAND2_X1 U5223 ( .A1(n5835), .A2(n4739), .ZN(n4717) );
  NOR2_X1 U5224 ( .A1(n4234), .A2(n4717), .ZN(n4733) );
  NAND2_X1 U5225 ( .A1(n4235), .A2(n4733), .ZN(n5526) );
  NOR2_X1 U5226 ( .A1(n4243), .A2(n5526), .ZN(n5354) );
  OR2_X1 U5227 ( .A1(n5356), .A2(n5354), .ZN(n4236) );
  OR2_X1 U5228 ( .A1(n5852), .A2(n5335), .ZN(n4238) );
  NAND2_X1 U5229 ( .A1(n5350), .A2(n4238), .ZN(n5331) );
  AOI21_X1 U5230 ( .B1(n4241), .B2(n4903), .A(n4245), .ZN(n4239) );
  AND2_X1 U5231 ( .A1(INSTADDRPOINTER_REG_26__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n4246) );
  NOR2_X1 U5232 ( .A1(n5852), .A2(n4246), .ZN(n4240) );
  NOR2_X1 U5233 ( .A1(n5318), .A2(n4240), .ZN(n4261) );
  INV_X1 U5234 ( .A(n4261), .ZN(n5297) );
  AND2_X1 U5235 ( .A1(n5262), .A2(REIP_REG_28__SCAN_IN), .ZN(n5191) );
  INV_X1 U5236 ( .A(n4900), .ZN(n4242) );
  NAND2_X1 U5237 ( .A1(n4242), .A2(n5841), .ZN(n4902) );
  NAND2_X1 U5238 ( .A1(n5526), .A2(n4902), .ZN(n5533) );
  NOR2_X1 U5239 ( .A1(n4243), .A2(n5786), .ZN(n5385) );
  INV_X1 U5240 ( .A(n5385), .ZN(n5503) );
  NAND2_X1 U5241 ( .A1(n5326), .A2(n4245), .ZN(n5307) );
  INV_X1 U5242 ( .A(n4246), .ZN(n4247) );
  XNOR2_X1 U5243 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .B(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n4248) );
  NOR2_X1 U5244 ( .A1(n5294), .A2(n4248), .ZN(n4249) );
  AOI211_X1 U5245 ( .C1(n5297), .C2(INSTADDRPOINTER_REG_28__SCAN_IN), .A(n5191), .B(n4249), .ZN(n4250) );
  NAND2_X1 U5246 ( .A1(n3680), .A2(n5302), .ZN(n5204) );
  INV_X1 U5247 ( .A(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5183) );
  AND2_X1 U5248 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_28__SCAN_IN), .ZN(n5284) );
  NAND2_X1 U5249 ( .A1(n5284), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n5275) );
  AOI21_X1 U5250 ( .B1(n5181), .B2(n5183), .A(n4488), .ZN(n4254) );
  INV_X1 U5251 ( .A(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4253) );
  XNOR2_X1 U5252 ( .A(n4254), .B(n4253), .ZN(n5008) );
  OR2_X1 U5253 ( .A1(n4468), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .ZN(n4256)
         );
  INV_X1 U5254 ( .A(EBX_REG_29__SCAN_IN), .ZN(n5106) );
  NAND2_X1 U5255 ( .A1(n4561), .A2(n5106), .ZN(n4255) );
  NAND2_X1 U5256 ( .A1(n4256), .A2(n4255), .ZN(n4463) );
  INV_X1 U5257 ( .A(n4463), .ZN(n4257) );
  NAND2_X1 U5258 ( .A1(n5022), .A2(n4159), .ZN(n4465) );
  OAI21_X1 U5259 ( .B1(n4257), .B2(n5022), .A(n4465), .ZN(n4260) );
  NAND2_X1 U5260 ( .A1(n4468), .A2(EBX_REG_30__SCAN_IN), .ZN(n4259) );
  NAND2_X1 U5261 ( .A1(n4178), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .ZN(n4258) );
  NAND2_X1 U5262 ( .A1(n4259), .A2(n4258), .ZN(n4467) );
  XNOR2_X1 U5263 ( .A(n4260), .B(n4467), .ZN(n4998) );
  NAND2_X1 U5264 ( .A1(n4998), .A2(n5834), .ZN(n4266) );
  INV_X1 U5265 ( .A(n5852), .ZN(n4262) );
  OAI21_X1 U5266 ( .B1(n5284), .B2(n5852), .A(n4261), .ZN(n5288) );
  AOI21_X1 U5267 ( .B1(n5183), .B2(n4262), .A(n5288), .ZN(n5274) );
  INV_X1 U5268 ( .A(n5274), .ZN(n4264) );
  AND2_X1 U5269 ( .A1(n5262), .A2(REIP_REG_30__SCAN_IN), .ZN(n5002) );
  NOR3_X1 U5270 ( .A1(n5294), .A2(INSTADDRPOINTER_REG_30__SCAN_IN), .A3(n5275), 
        .ZN(n4263) );
  AOI211_X1 U5271 ( .C1(n4264), .C2(INSTADDRPOINTER_REG_30__SCAN_IN), .A(n5002), .B(n4263), .ZN(n4265) );
  OAI21_X1 U5272 ( .B1(n5008), .B2(n5824), .A(n3254), .ZN(U2988) );
  AOI22_X1 U5273 ( .A1(n4341), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4270) );
  AOI22_X1 U5274 ( .A1(n4427), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_1__7__SCAN_IN), .ZN(n4269) );
  AOI22_X1 U5275 ( .A1(n3115), .A2(INSTQUEUE_REG_3__7__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_6__7__SCAN_IN), .ZN(n4268) );
  AOI22_X1 U5276 ( .A1(n3120), .A2(INSTQUEUE_REG_0__7__SCAN_IN), .B1(n3108), 
        .B2(INSTQUEUE_REG_15__7__SCAN_IN), .ZN(n4267) );
  NAND4_X1 U5277 ( .A1(n4270), .A2(n4269), .A3(n4268), .A4(n4267), .ZN(n4276)
         );
  AOI22_X1 U5278 ( .A1(n3112), .A2(INSTQUEUE_REG_8__7__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n4274) );
  AOI22_X1 U5279 ( .A1(n3107), .A2(INSTQUEUE_REG_4__7__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n4273) );
  AOI22_X1 U5280 ( .A1(n3110), .A2(INSTQUEUE_REG_7__7__SCAN_IN), .B1(n3106), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4272) );
  AOI22_X1 U5281 ( .A1(n4388), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4271) );
  NAND4_X1 U5282 ( .A1(n4274), .A2(n4273), .A3(n4272), .A4(n4271), .ZN(n4275)
         );
  NOR2_X1 U5283 ( .A1(n4276), .A2(n4275), .ZN(n4300) );
  AOI22_X1 U5284 ( .A1(n3112), .A2(INSTQUEUE_REG_9__0__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_11__0__SCAN_IN), .ZN(n4281) );
  AOI22_X1 U5285 ( .A1(n4407), .A2(INSTQUEUE_REG_5__0__SCAN_IN), .B1(n4359), 
        .B2(INSTQUEUE_REG_14__0__SCAN_IN), .ZN(n4280) );
  AOI22_X1 U5286 ( .A1(n3110), .A2(INSTQUEUE_REG_8__0__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_7__0__SCAN_IN), .ZN(n4279) );
  AOI22_X1 U5287 ( .A1(n3116), .A2(INSTQUEUE_REG_12__0__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_3__0__SCAN_IN), .ZN(n4278) );
  NAND4_X1 U5288 ( .A1(n4281), .A2(n4280), .A3(n4279), .A4(n4278), .ZN(n4287)
         );
  AOI22_X1 U5289 ( .A1(n4341), .A2(INSTQUEUE_REG_13__0__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n4285) );
  AOI22_X1 U5290 ( .A1(n3121), .A2(INSTQUEUE_REG_1__0__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n4284) );
  AOI22_X1 U5291 ( .A1(n3106), .A2(INSTQUEUE_REG_6__0__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__0__SCAN_IN), .ZN(n4283) );
  AOI22_X1 U5292 ( .A1(n3118), .A2(INSTQUEUE_REG_15__0__SCAN_IN), .B1(n4346), 
        .B2(INSTQUEUE_REG_0__0__SCAN_IN), .ZN(n4282) );
  NAND4_X1 U5293 ( .A1(n4285), .A2(n4284), .A3(n4283), .A4(n4282), .ZN(n4286)
         );
  NOR2_X1 U5294 ( .A1(n4287), .A2(n4286), .ZN(n4301) );
  XNOR2_X1 U5295 ( .A(n4300), .B(n4301), .ZN(n4291) );
  NAND2_X1 U5296 ( .A1(n6511), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4288)
         );
  NAND2_X1 U5297 ( .A1(n3791), .A2(n4288), .ZN(n4289) );
  AOI21_X1 U5298 ( .B1(n3764), .B2(EAX_REG_23__SCAN_IN), .A(n4289), .ZN(n4290)
         );
  OAI21_X1 U5299 ( .B1(n4422), .B2(n4291), .A(n4290), .ZN(n4298) );
  NOR2_X1 U5300 ( .A1(n4294), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n4295)
         );
  OR2_X1 U5301 ( .A1(n4312), .A2(n4295), .ZN(n5440) );
  INV_X1 U5302 ( .A(n5440), .ZN(n4296) );
  NAND2_X1 U5303 ( .A1(n4296), .A2(n4448), .ZN(n4297) );
  NAND2_X1 U5304 ( .A1(n4298), .A2(n4297), .ZN(n5139) );
  OR2_X1 U5305 ( .A1(n4301), .A2(n4300), .ZN(n4330) );
  AOI22_X1 U5306 ( .A1(n3118), .A2(INSTQUEUE_REG_15__1__SCAN_IN), .B1(n3120), 
        .B2(INSTQUEUE_REG_1__1__SCAN_IN), .ZN(n4305) );
  AOI22_X1 U5307 ( .A1(n4341), .A2(INSTQUEUE_REG_13__1__SCAN_IN), .B1(n3110), 
        .B2(INSTQUEUE_REG_8__1__SCAN_IN), .ZN(n4304) );
  AOI22_X1 U5308 ( .A1(n4277), .A2(INSTQUEUE_REG_9__1__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_10__1__SCAN_IN), .ZN(n4303) );
  AOI22_X1 U5309 ( .A1(n3116), .A2(INSTQUEUE_REG_12__1__SCAN_IN), .B1(n3106), 
        .B2(INSTQUEUE_REG_6__1__SCAN_IN), .ZN(n4302) );
  NAND4_X1 U5310 ( .A1(n4305), .A2(n4304), .A3(n4303), .A4(n4302), .ZN(n4311)
         );
  AOI22_X1 U5311 ( .A1(n3107), .A2(INSTQUEUE_REG_5__1__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_0__1__SCAN_IN), .ZN(n4309) );
  AOI22_X1 U5312 ( .A1(n3114), .A2(INSTQUEUE_REG_11__1__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n4308) );
  AOI22_X1 U5313 ( .A1(n4427), .A2(INSTQUEUE_REG_14__1__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n4307) );
  INV_X1 U5314 ( .A(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n6801) );
  AOI22_X1 U5315 ( .A1(n4434), .A2(INSTQUEUE_REG_2__1__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_3__1__SCAN_IN), .ZN(n4306) );
  NAND4_X1 U5316 ( .A1(n4309), .A2(n4308), .A3(n4307), .A4(n4306), .ZN(n4310)
         );
  NOR2_X1 U5317 ( .A1(n4311), .A2(n4310), .ZN(n4329) );
  XNOR2_X1 U5318 ( .A(n4330), .B(n4329), .ZN(n4318) );
  NOR2_X1 U5319 ( .A1(n4312), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4313)
         );
  NOR2_X1 U5320 ( .A1(n4335), .A2(n4313), .ZN(n5432) );
  NAND2_X1 U5321 ( .A1(n3764), .A2(EAX_REG_24__SCAN_IN), .ZN(n4315) );
  NAND2_X1 U5322 ( .A1(n4452), .A2(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n4314)
         );
  OAI211_X1 U5323 ( .C1(n5432), .C2(n3791), .A(n4315), .B(n4314), .ZN(n4316)
         );
  INV_X1 U5324 ( .A(n4316), .ZN(n4317) );
  OAI21_X1 U5325 ( .B1(n4422), .B2(n4318), .A(n4317), .ZN(n5133) );
  AOI22_X1 U5326 ( .A1(n4341), .A2(INSTQUEUE_REG_13__2__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_11__2__SCAN_IN), .ZN(n4322) );
  AOI22_X1 U5327 ( .A1(n3112), .A2(INSTQUEUE_REG_9__2__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_12__2__SCAN_IN), .ZN(n4321) );
  AOI22_X1 U5328 ( .A1(n3106), .A2(INSTQUEUE_REG_6__2__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__2__SCAN_IN), .ZN(n4320) );
  AOI22_X1 U5329 ( .A1(n3110), .A2(INSTQUEUE_REG_8__2__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_7__2__SCAN_IN), .ZN(n4319) );
  NAND4_X1 U5330 ( .A1(n4322), .A2(n4321), .A3(n4320), .A4(n4319), .ZN(n4328)
         );
  AOI22_X1 U5331 ( .A1(n3107), .A2(INSTQUEUE_REG_5__2__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n4326) );
  AOI22_X1 U5332 ( .A1(n4427), .A2(INSTQUEUE_REG_14__2__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_2__2__SCAN_IN), .ZN(n4325) );
  AOI22_X1 U5333 ( .A1(n4388), .A2(INSTQUEUE_REG_10__2__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_3__2__SCAN_IN), .ZN(n4324) );
  AOI22_X1 U5334 ( .A1(n3120), .A2(INSTQUEUE_REG_1__2__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_0__2__SCAN_IN), .ZN(n4323) );
  NAND4_X1 U5335 ( .A1(n4326), .A2(n4325), .A3(n4324), .A4(n4323), .ZN(n4327)
         );
  NOR2_X1 U5336 ( .A1(n4328), .A2(n4327), .ZN(n4340) );
  OR2_X1 U5337 ( .A1(n4330), .A2(n4329), .ZN(n4339) );
  XNOR2_X1 U5338 ( .A(n4340), .B(n4339), .ZN(n4334) );
  NAND2_X1 U5339 ( .A1(n6511), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4331)
         );
  NAND2_X1 U5340 ( .A1(n3791), .A2(n4331), .ZN(n4332) );
  AOI21_X1 U5341 ( .B1(n4453), .B2(EAX_REG_25__SCAN_IN), .A(n4332), .ZN(n4333)
         );
  OAI21_X1 U5342 ( .B1(n4334), .B2(n4422), .A(n4333), .ZN(n4338) );
  OR2_X1 U5343 ( .A1(n4335), .A2(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n4336)
         );
  NAND2_X1 U5344 ( .A1(n4336), .A2(n4376), .ZN(n5494) );
  NAND2_X1 U5345 ( .A1(n5123), .A2(n5122), .ZN(n5114) );
  NOR2_X1 U5346 ( .A1(n4340), .A2(n4339), .ZN(n4372) );
  AOI22_X1 U5347 ( .A1(n4341), .A2(INSTQUEUE_REG_13__3__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_11__3__SCAN_IN), .ZN(n4345) );
  AOI22_X1 U5348 ( .A1(n4277), .A2(INSTQUEUE_REG_9__3__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_12__3__SCAN_IN), .ZN(n4344) );
  AOI22_X1 U5349 ( .A1(n3106), .A2(INSTQUEUE_REG_6__3__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__3__SCAN_IN), .ZN(n4343) );
  AOI22_X1 U5350 ( .A1(n3110), .A2(INSTQUEUE_REG_8__3__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_7__3__SCAN_IN), .ZN(n4342) );
  NAND4_X1 U5351 ( .A1(n4345), .A2(n4344), .A3(n4343), .A4(n4342), .ZN(n4352)
         );
  AOI22_X1 U5352 ( .A1(n4407), .A2(INSTQUEUE_REG_5__3__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_15__3__SCAN_IN), .ZN(n4350) );
  AOI22_X1 U5353 ( .A1(n4427), .A2(INSTQUEUE_REG_14__3__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_2__3__SCAN_IN), .ZN(n4349) );
  AOI22_X1 U5354 ( .A1(n4388), .A2(INSTQUEUE_REG_10__3__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_3__3__SCAN_IN), .ZN(n4348) );
  AOI22_X1 U5355 ( .A1(n3120), .A2(INSTQUEUE_REG_1__3__SCAN_IN), .B1(n3108), 
        .B2(INSTQUEUE_REG_0__3__SCAN_IN), .ZN(n4347) );
  NAND4_X1 U5356 ( .A1(n4350), .A2(n4349), .A3(n4348), .A4(n4347), .ZN(n4351)
         );
  OR2_X1 U5357 ( .A1(n4352), .A2(n4351), .ZN(n4371) );
  XNOR2_X1 U5358 ( .A(n4372), .B(n4371), .ZN(n4356) );
  NAND2_X1 U5359 ( .A1(n6511), .A2(PHYADDRPOINTER_REG_26__SCAN_IN), .ZN(n4353)
         );
  NAND2_X1 U5360 ( .A1(n3791), .A2(n4353), .ZN(n4354) );
  AOI21_X1 U5361 ( .B1(n4453), .B2(EAX_REG_26__SCAN_IN), .A(n4354), .ZN(n4355)
         );
  OAI21_X1 U5362 ( .B1(n4356), .B2(n4422), .A(n4355), .ZN(n4358) );
  XNOR2_X1 U5363 ( .A(PHYADDRPOINTER_REG_26__SCAN_IN), .B(n4376), .ZN(n5413)
         );
  NAND2_X1 U5364 ( .A1(n4448), .A2(n5413), .ZN(n4357) );
  NAND2_X1 U5365 ( .A1(n4358), .A2(n4357), .ZN(n5115) );
  NOR2_X2 U5366 ( .A1(n5114), .A2(n5115), .ZN(n5108) );
  AOI22_X1 U5367 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n3111), .B1(n3114), 
        .B2(INSTQUEUE_REG_11__4__SCAN_IN), .ZN(n4363) );
  AOI22_X1 U5368 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n3107), .B1(n4359), 
        .B2(INSTQUEUE_REG_14__4__SCAN_IN), .ZN(n4362) );
  AOI22_X1 U5369 ( .A1(n3106), .A2(INSTQUEUE_REG_6__4__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_7__4__SCAN_IN), .ZN(n4361) );
  AOI22_X1 U5370 ( .A1(n3118), .A2(INSTQUEUE_REG_15__4__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_3__4__SCAN_IN), .ZN(n4360) );
  NAND4_X1 U5371 ( .A1(n4363), .A2(n4362), .A3(n4361), .A4(n4360), .ZN(n4370)
         );
  AOI22_X1 U5372 ( .A1(n4341), .A2(INSTQUEUE_REG_13__4__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_12__4__SCAN_IN), .ZN(n4368) );
  AOI22_X1 U5373 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n3120), .B1(n4434), 
        .B2(INSTQUEUE_REG_2__4__SCAN_IN), .ZN(n4367) );
  AOI22_X1 U5374 ( .A1(n3110), .A2(INSTQUEUE_REG_8__4__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__4__SCAN_IN), .ZN(n4366) );
  AOI22_X1 U5375 ( .A1(n4388), .A2(INSTQUEUE_REG_10__4__SCAN_IN), .B1(n3108), 
        .B2(INSTQUEUE_REG_0__4__SCAN_IN), .ZN(n4365) );
  NAND4_X1 U5376 ( .A1(n4368), .A2(n4367), .A3(n4366), .A4(n4365), .ZN(n4369)
         );
  NOR2_X1 U5377 ( .A1(n4370), .A2(n4369), .ZN(n4396) );
  NAND2_X1 U5378 ( .A1(n4372), .A2(n4371), .ZN(n4395) );
  XNOR2_X1 U5379 ( .A(n4396), .B(n4395), .ZN(n4375) );
  INV_X1 U5380 ( .A(PHYADDRPOINTER_REG_27__SCAN_IN), .ZN(n5406) );
  AOI21_X1 U5381 ( .B1(n5406), .B2(STATEBS16_REG_SCAN_IN), .A(
        STATE2_REG_2__SCAN_IN), .ZN(n4373) );
  AOI21_X1 U5382 ( .B1(n4453), .B2(EAX_REG_27__SCAN_IN), .A(n4373), .ZN(n4374)
         );
  OAI21_X1 U5383 ( .B1(n4375), .B2(n4422), .A(n4374), .ZN(n4382) );
  INV_X1 U5384 ( .A(n4376), .ZN(n4377) );
  INV_X1 U5385 ( .A(n4378), .ZN(n4379) );
  NAND2_X1 U5386 ( .A1(n4379), .A2(n5406), .ZN(n4380) );
  NAND2_X1 U5387 ( .A1(n4403), .A2(n4380), .ZN(n5405) );
  NAND2_X1 U5388 ( .A1(n4382), .A2(n4381), .ZN(n5109) );
  AND2_X2 U5389 ( .A1(n5108), .A2(n4383), .ZN(n5034) );
  XNOR2_X1 U5390 ( .A(n4403), .B(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5037)
         );
  AOI22_X1 U5391 ( .A1(n4341), .A2(INSTQUEUE_REG_13__5__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_11__5__SCAN_IN), .ZN(n4387) );
  AOI22_X1 U5392 ( .A1(n3111), .A2(INSTQUEUE_REG_9__5__SCAN_IN), .B1(n3116), 
        .B2(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n4386) );
  AOI22_X1 U5393 ( .A1(n3106), .A2(INSTQUEUE_REG_6__5__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__5__SCAN_IN), .ZN(n4385) );
  AOI22_X1 U5394 ( .A1(n3110), .A2(INSTQUEUE_REG_8__5__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_7__5__SCAN_IN), .ZN(n4384) );
  NAND4_X1 U5395 ( .A1(n4387), .A2(n4386), .A3(n4385), .A4(n4384), .ZN(n4394)
         );
  AOI22_X1 U5396 ( .A1(n3107), .A2(INSTQUEUE_REG_5__5__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n4392) );
  AOI22_X1 U5397 ( .A1(n4427), .A2(INSTQUEUE_REG_14__5__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_2__5__SCAN_IN), .ZN(n4391) );
  AOI22_X1 U5398 ( .A1(n4388), .A2(INSTQUEUE_REG_10__5__SCAN_IN), .B1(n3103), 
        .B2(INSTQUEUE_REG_3__5__SCAN_IN), .ZN(n4390) );
  AOI22_X1 U5399 ( .A1(n3121), .A2(INSTQUEUE_REG_1__5__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n4389) );
  NAND4_X1 U5400 ( .A1(n4392), .A2(n4391), .A3(n4390), .A4(n4389), .ZN(n4393)
         );
  OR2_X1 U5401 ( .A1(n4394), .A2(n4393), .ZN(n4418) );
  NOR2_X1 U5402 ( .A1(n4396), .A2(n4395), .ZN(n4419) );
  XOR2_X1 U5403 ( .A(n4418), .B(n4419), .Z(n4401) );
  INV_X1 U5404 ( .A(n4422), .ZN(n4444) );
  INV_X1 U5405 ( .A(EAX_REG_28__SCAN_IN), .ZN(n4398) );
  OAI21_X1 U5406 ( .B1(n6286), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n6511), 
        .ZN(n4397) );
  OAI21_X1 U5407 ( .B1(n4399), .B2(n4398), .A(n4397), .ZN(n4400) );
  AOI21_X1 U5408 ( .B1(n4401), .B2(n4444), .A(n4400), .ZN(n4402) );
  AOI21_X1 U5409 ( .B1(n4448), .B2(n5037), .A(n4402), .ZN(n5035) );
  INV_X1 U5410 ( .A(PHYADDRPOINTER_REG_28__SCAN_IN), .ZN(n5038) );
  INV_X1 U5411 ( .A(n4404), .ZN(n4405) );
  INV_X1 U5412 ( .A(PHYADDRPOINTER_REG_29__SCAN_IN), .ZN(n5021) );
  NAND2_X1 U5413 ( .A1(n4405), .A2(n5021), .ZN(n4406) );
  NAND2_X1 U5414 ( .A1(n4459), .A2(n4406), .ZN(n5186) );
  AOI22_X1 U5415 ( .A1(n4341), .A2(INSTQUEUE_REG_13__6__SCAN_IN), .B1(n3114), 
        .B2(INSTQUEUE_REG_11__6__SCAN_IN), .ZN(n4411) );
  AOI22_X1 U5416 ( .A1(n4277), .A2(INSTQUEUE_REG_9__6__SCAN_IN), .B1(n3118), 
        .B2(INSTQUEUE_REG_15__6__SCAN_IN), .ZN(n4410) );
  AOI22_X1 U5417 ( .A1(n3115), .A2(INSTQUEUE_REG_4__6__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n4409) );
  AOI22_X1 U5418 ( .A1(n3107), .A2(INSTQUEUE_REG_5__6__SCAN_IN), .B1(n4346), 
        .B2(INSTQUEUE_REG_0__6__SCAN_IN), .ZN(n4408) );
  NAND4_X1 U5419 ( .A1(n4411), .A2(n4410), .A3(n4409), .A4(n4408), .ZN(n4417)
         );
  AOI22_X1 U5420 ( .A1(n3110), .A2(INSTQUEUE_REG_8__6__SCAN_IN), .B1(n3106), 
        .B2(INSTQUEUE_REG_6__6__SCAN_IN), .ZN(n4415) );
  AOI22_X1 U5421 ( .A1(n3116), .A2(INSTQUEUE_REG_12__6__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_10__6__SCAN_IN), .ZN(n4414) );
  AOI22_X1 U5422 ( .A1(n4427), .A2(INSTQUEUE_REG_14__6__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_2__6__SCAN_IN), .ZN(n4413) );
  AOI22_X1 U5423 ( .A1(n3120), .A2(INSTQUEUE_REG_1__6__SCAN_IN), .B1(n3102), 
        .B2(INSTQUEUE_REG_3__6__SCAN_IN), .ZN(n4412) );
  NAND4_X1 U5424 ( .A1(n4415), .A2(n4414), .A3(n4413), .A4(n4412), .ZN(n4416)
         );
  NOR2_X1 U5425 ( .A1(n4417), .A2(n4416), .ZN(n4426) );
  NAND2_X1 U5426 ( .A1(n4419), .A2(n4418), .ZN(n4425) );
  XNOR2_X1 U5427 ( .A(n4426), .B(n4425), .ZN(n4423) );
  AOI21_X1 U5428 ( .B1(PHYADDRPOINTER_REG_29__SCAN_IN), .B2(n6511), .A(n4448), 
        .ZN(n4421) );
  NAND2_X1 U5429 ( .A1(n3764), .A2(EAX_REG_29__SCAN_IN), .ZN(n4420) );
  OAI211_X1 U5430 ( .C1(n4423), .C2(n4422), .A(n4421), .B(n4420), .ZN(n4424)
         );
  OAI21_X1 U5431 ( .B1(n3791), .B2(n5186), .A(n4424), .ZN(n5020) );
  NOR2_X1 U5432 ( .A1(n4426), .A2(n4425), .ZN(n4443) );
  AOI22_X1 U5433 ( .A1(n3116), .A2(INSTQUEUE_REG_12__7__SCAN_IN), .B1(n4388), 
        .B2(INSTQUEUE_REG_10__7__SCAN_IN), .ZN(n4432) );
  AOI22_X1 U5434 ( .A1(n3114), .A2(INSTQUEUE_REG_11__7__SCAN_IN), .B1(n3104), 
        .B2(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n4431) );
  AOI22_X1 U5435 ( .A1(n4427), .A2(INSTQUEUE_REG_14__7__SCAN_IN), .B1(n3109), 
        .B2(INSTQUEUE_REG_0__7__SCAN_IN), .ZN(n4430) );
  AOI22_X1 U5436 ( .A1(n3118), .A2(INSTQUEUE_REG_15__7__SCAN_IN), .B1(n3333), 
        .B2(INSTQUEUE_REG_3__7__SCAN_IN), .ZN(n4429) );
  NAND4_X1 U5437 ( .A1(n4432), .A2(n4431), .A3(n4430), .A4(n4429), .ZN(n4441)
         );
  AOI22_X1 U5438 ( .A1(n4341), .A2(INSTQUEUE_REG_13__7__SCAN_IN), .B1(n3110), 
        .B2(INSTQUEUE_REG_8__7__SCAN_IN), .ZN(n4439) );
  AOI22_X1 U5439 ( .A1(n3112), .A2(INSTQUEUE_REG_9__7__SCAN_IN), .B1(n4407), 
        .B2(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n4438) );
  AOI22_X1 U5440 ( .A1(n3383), .A2(INSTQUEUE_REG_1__7__SCAN_IN), .B1(n4434), 
        .B2(INSTQUEUE_REG_2__7__SCAN_IN), .ZN(n4437) );
  AOI22_X1 U5441 ( .A1(n3106), .A2(INSTQUEUE_REG_6__7__SCAN_IN), .B1(n3115), 
        .B2(INSTQUEUE_REG_4__7__SCAN_IN), .ZN(n4436) );
  NAND4_X1 U5442 ( .A1(n4439), .A2(n4438), .A3(n4437), .A4(n4436), .ZN(n4440)
         );
  NOR2_X1 U5443 ( .A1(n4441), .A2(n4440), .ZN(n4442) );
  XNOR2_X1 U5444 ( .A(n4443), .B(n4442), .ZN(n4445) );
  NAND2_X1 U5445 ( .A1(n4445), .A2(n4444), .ZN(n4451) );
  NAND2_X1 U5446 ( .A1(n6511), .A2(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4446)
         );
  NAND2_X1 U5447 ( .A1(n3791), .A2(n4446), .ZN(n4447) );
  AOI21_X1 U5448 ( .B1(n4453), .B2(EAX_REG_30__SCAN_IN), .A(n4447), .ZN(n4450)
         );
  XNOR2_X1 U5449 ( .A(n4459), .B(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n5001)
         );
  AND2_X1 U5450 ( .A1(n5001), .A2(n4448), .ZN(n4449) );
  AOI21_X1 U5451 ( .B1(n4451), .B2(n4450), .A(n4449), .ZN(n4494) );
  AOI22_X1 U5452 ( .A1(n4453), .A2(EAX_REG_31__SCAN_IN), .B1(
        PHYADDRPOINTER_REG_31__SCAN_IN), .B2(n4452), .ZN(n4454) );
  INV_X1 U5453 ( .A(n4454), .ZN(n4455) );
  NAND2_X1 U5454 ( .A1(n4510), .A2(n6518), .ZN(n4505) );
  INV_X1 U5455 ( .A(n6631), .ZN(n6529) );
  NOR3_X1 U5456 ( .A1(n6521), .A2(n6598), .A3(n6529), .ZN(n6516) );
  NOR3_X1 U5457 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n6522), .A3(n3791), .ZN(
        n6528) );
  INV_X1 U5458 ( .A(PHYADDRPOINTER_REG_30__SCAN_IN), .ZN(n4458) );
  INV_X1 U5459 ( .A(PHYADDRPOINTER_REG_31__SCAN_IN), .ZN(n4460) );
  NOR2_X1 U5460 ( .A1(n4820), .A2(n6522), .ZN(n4462) );
  NAND2_X1 U5461 ( .A1(n4463), .A2(n4159), .ZN(n4466) );
  NAND2_X1 U5462 ( .A1(n4122), .A2(EBX_REG_29__SCAN_IN), .ZN(n4464) );
  NAND2_X1 U5463 ( .A1(n4466), .A2(n4464), .ZN(n5023) );
  OAI22_X1 U5464 ( .A1(n4468), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .B1(
        EBX_REG_31__SCAN_IN), .B2(n4178), .ZN(n4469) );
  NAND2_X1 U5465 ( .A1(n6628), .A2(n6286), .ZN(n4814) );
  NAND2_X1 U5466 ( .A1(n4814), .A2(EBX_REG_31__SCAN_IN), .ZN(n4470) );
  NOR2_X1 U5467 ( .A1(n4178), .A2(n4470), .ZN(n4471) );
  OR2_X1 U5468 ( .A1(n6539), .A2(n4814), .ZN(n6506) );
  NAND2_X1 U5469 ( .A1(n3428), .A2(n6506), .ZN(n4816) );
  INV_X1 U5470 ( .A(EBX_REG_31__SCAN_IN), .ZN(n6734) );
  NOR2_X1 U5471 ( .A1(n4816), .A2(n6734), .ZN(n4472) );
  AOI22_X1 U5472 ( .A1(PHYADDRPOINTER_REG_31__SCAN_IN), .A2(n5674), .B1(n4819), 
        .B2(n4472), .ZN(n4479) );
  NAND3_X1 U5473 ( .A1(REIP_REG_20__SCAN_IN), .A2(REIP_REG_19__SCAN_IN), .A3(
        REIP_REG_18__SCAN_IN), .ZN(n4481) );
  INV_X1 U5474 ( .A(REIP_REG_14__SCAN_IN), .ZN(n6563) );
  NAND2_X1 U5475 ( .A1(REIP_REG_13__SCAN_IN), .A2(REIP_REG_12__SCAN_IN), .ZN(
        n4914) );
  INV_X1 U5476 ( .A(n5687), .ZN(n5649) );
  INV_X1 U5477 ( .A(REIP_REG_6__SCAN_IN), .ZN(n6557) );
  INV_X1 U5478 ( .A(REIP_REG_4__SCAN_IN), .ZN(n6929) );
  NAND3_X1 U5479 ( .A1(REIP_REG_2__SCAN_IN), .A2(REIP_REG_1__SCAN_IN), .A3(
        REIP_REG_3__SCAN_IN), .ZN(n5652) );
  NOR2_X1 U5480 ( .A1(n6929), .A2(n5652), .ZN(n5636) );
  NAND2_X1 U5481 ( .A1(REIP_REG_5__SCAN_IN), .A2(n5636), .ZN(n5618) );
  NOR2_X1 U5482 ( .A1(n6557), .A2(n5618), .ZN(n5097) );
  NAND3_X1 U5483 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_7__SCAN_IN), .A3(
        n5097), .ZN(n4480) );
  NOR2_X1 U5484 ( .A1(n5649), .A2(n4480), .ZN(n5089) );
  NAND4_X1 U5485 ( .A1(REIP_REG_11__SCAN_IN), .A2(REIP_REG_9__SCAN_IN), .A3(
        REIP_REG_10__SCAN_IN), .A4(n5089), .ZN(n4867) );
  NOR3_X1 U5486 ( .A1(n6563), .A2(n4914), .A3(n4867), .ZN(n4924) );
  NAND4_X1 U5487 ( .A1(REIP_REG_17__SCAN_IN), .A2(REIP_REG_16__SCAN_IN), .A3(
        REIP_REG_15__SCAN_IN), .A4(n4924), .ZN(n5081) );
  NOR2_X1 U5488 ( .A1(n4481), .A2(n5081), .ZN(n5045) );
  NAND4_X1 U5489 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5045), .ZN(n5427) );
  NAND3_X1 U5490 ( .A1(REIP_REG_24__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        REIP_REG_25__SCAN_IN), .ZN(n4482) );
  INV_X1 U5491 ( .A(n4814), .ZN(n4473) );
  AND3_X1 U5492 ( .A1(n4474), .A2(n4473), .A3(n3407), .ZN(n4475) );
  NAND2_X1 U5493 ( .A1(n5653), .A2(n5687), .ZN(n5688) );
  OAI21_X1 U5494 ( .B1(n5427), .B2(n4482), .A(n5688), .ZN(n5414) );
  INV_X1 U5495 ( .A(REIP_REG_28__SCAN_IN), .ZN(n6582) );
  INV_X1 U5496 ( .A(REIP_REG_27__SCAN_IN), .ZN(n6580) );
  NOR2_X1 U5497 ( .A1(n6582), .A2(n6580), .ZN(n4476) );
  OR2_X1 U5498 ( .A1(n5653), .A2(n4476), .ZN(n5036) );
  AND2_X1 U5499 ( .A1(n5036), .A2(REIP_REG_29__SCAN_IN), .ZN(n4477) );
  NAND2_X1 U5500 ( .A1(n5414), .A2(n4477), .ZN(n5030) );
  INV_X1 U5501 ( .A(REIP_REG_30__SCAN_IN), .ZN(n6584) );
  OAI211_X1 U5502 ( .C1(n5030), .C2(n6584), .A(REIP_REG_31__SCAN_IN), .B(n5688), .ZN(n4478) );
  OAI211_X1 U5503 ( .C1(n5279), .C2(n5681), .A(n4479), .B(n4478), .ZN(n4484)
         );
  NAND4_X1 U5504 ( .A1(n5608), .A2(REIP_REG_11__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .A4(REIP_REG_10__SCAN_IN), .ZN(n5602) );
  NAND2_X1 U5505 ( .A1(REIP_REG_14__SCAN_IN), .A2(n4925), .ZN(n5591) );
  NAND2_X1 U5506 ( .A1(REIP_REG_16__SCAN_IN), .A2(REIP_REG_15__SCAN_IN), .ZN(
        n4977) );
  NAND2_X1 U5507 ( .A1(REIP_REG_17__SCAN_IN), .A2(n5579), .ZN(n5073) );
  NAND4_X1 U5508 ( .A1(REIP_REG_23__SCAN_IN), .A2(REIP_REG_22__SCAN_IN), .A3(
        REIP_REG_21__SCAN_IN), .A4(n5048), .ZN(n5428) );
  NOR2_X1 U5509 ( .A1(n5428), .A2(n4482), .ZN(n5409) );
  NAND3_X1 U5510 ( .A1(n5409), .A2(REIP_REG_28__SCAN_IN), .A3(
        REIP_REG_27__SCAN_IN), .ZN(n5029) );
  INV_X1 U5511 ( .A(REIP_REG_29__SCAN_IN), .ZN(n6585) );
  NOR4_X1 U5512 ( .A1(n5029), .A2(REIP_REG_31__SCAN_IN), .A3(n6584), .A4(n6585), .ZN(n4483) );
  INV_X1 U5513 ( .A(INSTADDRPOINTER_REG_31__SCAN_IN), .ZN(n4553) );
  XNOR2_X1 U5514 ( .A(n4489), .B(n4553), .ZN(n5283) );
  AND2_X1 U5515 ( .A1(n5832), .A2(REIP_REG_31__SCAN_IN), .ZN(n5277) );
  AOI21_X1 U5516 ( .B1(n5777), .B2(PHYADDRPOINTER_REG_31__SCAN_IN), .A(n5277), 
        .ZN(n4490) );
  OAI21_X1 U5517 ( .B1(n5773), .B2(n4820), .A(n4490), .ZN(n4491) );
  INV_X1 U5518 ( .A(n4491), .ZN(n4493) );
  NAND2_X1 U5519 ( .A1(n5166), .A2(n5768), .ZN(n4492) );
  OAI211_X1 U5520 ( .C1(n5283), .C2(n5557), .A(n4493), .B(n4492), .ZN(U2955)
         );
  NAND4_X1 U5521 ( .A1(n3435), .A2(n4495), .A3(n5165), .A4(n3409), .ZN(n4599)
         );
  INV_X1 U5522 ( .A(n4599), .ZN(n4498) );
  INV_X1 U5523 ( .A(n4496), .ZN(n4497) );
  NAND3_X1 U5524 ( .A1(n4498), .A2(n4497), .A3(n4561), .ZN(n4499) );
  NAND2_X1 U5525 ( .A1(n5006), .A2(n5703), .ZN(n4504) );
  INV_X1 U5526 ( .A(EBX_REG_30__SCAN_IN), .ZN(n4995) );
  NOR2_X1 U5527 ( .A1(n5706), .A2(n4995), .ZN(n4501) );
  NAND2_X1 U5528 ( .A1(n4504), .A2(n4503), .ZN(U2829) );
  NOR2_X1 U5529 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6410), .ZN(n4866) );
  AOI21_X1 U5530 ( .B1(MEMORYFETCH_REG_SCAN_IN), .B2(n4505), .A(n4866), .ZN(
        n4506) );
  NAND2_X1 U5531 ( .A1(n4525), .A2(n4506), .ZN(U2788) );
  INV_X1 U5532 ( .A(n6626), .ZN(n4509) );
  INV_X1 U5533 ( .A(n4507), .ZN(n4818) );
  OR2_X1 U5534 ( .A1(n3428), .A2(n4818), .ZN(n4514) );
  OAI21_X1 U5535 ( .B1(n4866), .B2(READREQUEST_REG_SCAN_IN), .A(n4509), .ZN(
        n4508) );
  OAI21_X1 U5536 ( .B1(n4509), .B2(n4514), .A(n4508), .ZN(U3474) );
  OR2_X1 U5537 ( .A1(n6513), .A2(n4812), .ZN(n4513) );
  INV_X1 U5538 ( .A(n4510), .ZN(n4511) );
  NAND2_X1 U5539 ( .A1(n4511), .A2(n4515), .ZN(n4512) );
  NAND2_X1 U5540 ( .A1(n4513), .A2(n4512), .ZN(n5552) );
  AOI21_X1 U5541 ( .B1(n4514), .B2(n6539), .A(READY_N), .ZN(n6629) );
  NOR2_X1 U5542 ( .A1(n5552), .A2(n6629), .ZN(n6497) );
  INV_X1 U5543 ( .A(n6518), .ZN(n6525) );
  NOR2_X1 U5544 ( .A1(n6497), .A2(n6525), .ZN(n5559) );
  INV_X1 U5545 ( .A(MORE_REG_SCAN_IN), .ZN(n4523) );
  NAND2_X1 U5546 ( .A1(n6496), .A2(n4515), .ZN(n4516) );
  NOR2_X1 U5547 ( .A1(n4557), .A2(n4516), .ZN(n4517) );
  OR2_X1 U5548 ( .A1(n6513), .A2(n4517), .ZN(n4520) );
  INV_X1 U5549 ( .A(n4653), .ZN(n4518) );
  NAND2_X1 U5550 ( .A1(n6513), .A2(n4518), .ZN(n4519) );
  OAI211_X1 U5551 ( .C1(n4521), .C2(n4102), .A(n4520), .B(n4519), .ZN(n6499)
         );
  NAND2_X1 U5552 ( .A1(n5559), .A2(n6499), .ZN(n4522) );
  OAI21_X1 U5553 ( .B1(n5559), .B2(n4523), .A(n4522), .ZN(U3471) );
  INV_X1 U5554 ( .A(n4525), .ZN(n4524) );
  INV_X2 U5555 ( .A(n5762), .ZN(n5756) );
  AOI22_X1 U5556 ( .A1(n5753), .A2(LWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_7__SCAN_IN), .B2(n5756), .ZN(n4526) );
  NAND2_X1 U5557 ( .A1(n5759), .A2(DATAI_7_), .ZN(n4624) );
  NAND2_X1 U5558 ( .A1(n4526), .A2(n4624), .ZN(U2946) );
  AOI22_X1 U5559 ( .A1(n5753), .A2(LWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_14__SCAN_IN), .B2(n5756), .ZN(n4527) );
  NAND2_X1 U5560 ( .A1(n5759), .A2(DATAI_14_), .ZN(n4631) );
  NAND2_X1 U5561 ( .A1(n4527), .A2(n4631), .ZN(U2953) );
  AOI22_X1 U5562 ( .A1(n5753), .A2(UWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_21__SCAN_IN), .B2(n5756), .ZN(n4528) );
  NAND2_X1 U5563 ( .A1(n5759), .A2(DATAI_5_), .ZN(n4629) );
  NAND2_X1 U5564 ( .A1(n4528), .A2(n4629), .ZN(U2929) );
  AOI22_X1 U5565 ( .A1(n5753), .A2(LWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_12__SCAN_IN), .B2(n5756), .ZN(n4529) );
  NAND2_X1 U5566 ( .A1(n5759), .A2(DATAI_12_), .ZN(n4627) );
  NAND2_X1 U5567 ( .A1(n4529), .A2(n4627), .ZN(U2951) );
  AOI22_X1 U5568 ( .A1(n5753), .A2(UWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_19__SCAN_IN), .B2(n5756), .ZN(n4530) );
  NAND2_X1 U5569 ( .A1(n5759), .A2(DATAI_3_), .ZN(n4637) );
  NAND2_X1 U5570 ( .A1(n4530), .A2(n4637), .ZN(U2927) );
  AOI22_X1 U5571 ( .A1(n5753), .A2(UWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_20__SCAN_IN), .B2(n5756), .ZN(n4531) );
  NAND2_X1 U5572 ( .A1(n5759), .A2(DATAI_4_), .ZN(n4622) );
  NAND2_X1 U5573 ( .A1(n4531), .A2(n4622), .ZN(U2928) );
  AOI22_X1 U5574 ( .A1(n5753), .A2(UWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_22__SCAN_IN), .B2(n5756), .ZN(n4532) );
  NAND2_X1 U5575 ( .A1(n5759), .A2(DATAI_6_), .ZN(n4635) );
  NAND2_X1 U5576 ( .A1(n4532), .A2(n4635), .ZN(U2930) );
  INV_X1 U5577 ( .A(UWORD_REG_10__SCAN_IN), .ZN(n6879) );
  NAND2_X1 U5578 ( .A1(n5759), .A2(DATAI_10_), .ZN(n5757) );
  NAND2_X1 U5579 ( .A1(n5756), .A2(EAX_REG_26__SCAN_IN), .ZN(n4533) );
  OAI211_X1 U5580 ( .C1(n4612), .C2(n6879), .A(n5757), .B(n4533), .ZN(U2934)
         );
  INV_X1 U5581 ( .A(DATAI_0_), .ZN(n4535) );
  INV_X1 U5582 ( .A(UWORD_REG_0__SCAN_IN), .ZN(n6816) );
  INV_X1 U5583 ( .A(EAX_REG_16__SCAN_IN), .ZN(n4534) );
  OAI222_X1 U5584 ( .A1(n4535), .A2(n4641), .B1(n4612), .B2(n6816), .C1(n4534), 
        .C2(n5762), .ZN(U2924) );
  INV_X1 U5585 ( .A(DATAI_1_), .ZN(n4537) );
  INV_X1 U5586 ( .A(UWORD_REG_1__SCAN_IN), .ZN(n4541) );
  INV_X1 U5587 ( .A(EAX_REG_17__SCAN_IN), .ZN(n4536) );
  OAI222_X1 U5588 ( .A1(n4537), .A2(n4641), .B1(n4541), .B2(n4612), .C1(n4536), 
        .C2(n5762), .ZN(U2925) );
  OR2_X1 U5589 ( .A1(n4538), .A2(n6478), .ZN(n4539) );
  NAND2_X1 U5590 ( .A1(n5762), .A2(n4539), .ZN(n4540) );
  INV_X1 U5591 ( .A(n6539), .ZN(n4562) );
  NAND2_X1 U5592 ( .A1(n4680), .A2(n6521), .ZN(n5746) );
  INV_X1 U5593 ( .A(DATAO_REG_17__SCAN_IN), .ZN(n6766) );
  NAND2_X1 U5594 ( .A1(n5739), .A2(n3407), .ZN(n5714) );
  OAI222_X1 U5595 ( .A1(n5749), .A2(n6766), .B1(n5714), .B2(n4536), .C1(n5746), 
        .C2(n4541), .ZN(U2906) );
  NAND2_X1 U5596 ( .A1(n4220), .A2(n4544), .ZN(n4545) );
  NOR2_X1 U5597 ( .A1(n4107), .A2(n4545), .ZN(n4548) );
  INV_X1 U5598 ( .A(n4546), .ZN(n4547) );
  AND3_X1 U5599 ( .A1(n4114), .A2(n4548), .A3(n4547), .ZN(n6476) );
  INV_X1 U5600 ( .A(n6476), .ZN(n4659) );
  NAND2_X1 U5601 ( .A1(n4543), .A2(n4659), .ZN(n4552) );
  OR3_X1 U5602 ( .A1(n6475), .A2(n4549), .A3(n4550), .ZN(n4551) );
  OAI211_X1 U5603 ( .C1(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .C2(n6478), .A(n4552), .B(n4551), .ZN(n6481) );
  INV_X1 U5604 ( .A(n6614), .ZN(n6606) );
  NOR2_X1 U5605 ( .A1(n6522), .A2(n6605), .ZN(n4555) );
  AOI22_X1 U5606 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n4553), .B1(
        INSTADDRPOINTER_REG_31__SCAN_IN), .B2(n5858), .ZN(n5010) );
  INV_X1 U5607 ( .A(n6601), .ZN(n5009) );
  AOI222_X1 U5608 ( .A1(n6481), .A2(n6606), .B1(n4555), .B2(n5010), .C1(n4554), 
        .C2(n5009), .ZN(n4573) );
  INV_X1 U5609 ( .A(n4556), .ZN(n4570) );
  NAND2_X1 U5610 ( .A1(n6513), .A2(n4557), .ZN(n4560) );
  INV_X1 U5611 ( .A(n4114), .ZN(n5547) );
  NAND2_X1 U5612 ( .A1(n5547), .A2(n4558), .ZN(n4559) );
  NAND2_X1 U5613 ( .A1(n4560), .A2(n4559), .ZN(n4602) );
  OAI21_X1 U5614 ( .B1(n4562), .B2(n4561), .A(n4107), .ZN(n4563) );
  OAI21_X1 U5615 ( .B1(n6478), .B2(n6539), .A(n4563), .ZN(n4564) );
  NAND3_X1 U5616 ( .A1(n6513), .A2(n6628), .A3(n4564), .ZN(n4568) );
  INV_X1 U5617 ( .A(n4565), .ZN(n4566) );
  NAND3_X1 U5618 ( .A1(n4568), .A2(n4567), .A3(n4566), .ZN(n4569) );
  INV_X1 U5619 ( .A(FLUSH_REG_SCAN_IN), .ZN(n5558) );
  NAND2_X1 U5620 ( .A1(STATE2_REG_0__SCAN_IN), .A2(n4680), .ZN(n6596) );
  NOR2_X1 U5621 ( .A1(n5558), .A2(n6596), .ZN(n4571) );
  AOI21_X1 U5622 ( .B1(n6518), .B2(n6480), .A(n4571), .ZN(n5550) );
  NAND2_X1 U5623 ( .A1(n6521), .A2(STATE2_REG_3__SCAN_IN), .ZN(n6597) );
  NAND2_X1 U5624 ( .A1(n5550), .A2(n6597), .ZN(n6612) );
  INV_X1 U5625 ( .A(n6612), .ZN(n5015) );
  NOR2_X1 U5626 ( .A1(n6601), .A2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .ZN(n6608)
         );
  OAI21_X1 U5627 ( .B1(n5015), .B2(n6608), .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), 
        .ZN(n4572) );
  OAI21_X1 U5628 ( .B1(n4573), .B2(n5015), .A(n4572), .ZN(U3460) );
  INV_X1 U5629 ( .A(EAX_REG_24__SCAN_IN), .ZN(n5752) );
  AOI22_X1 U5630 ( .A1(n5738), .A2(UWORD_REG_8__SCAN_IN), .B1(n5743), .B2(
        DATAO_REG_24__SCAN_IN), .ZN(n4574) );
  OAI21_X1 U5631 ( .B1(n5752), .B2(n5714), .A(n4574), .ZN(U2899) );
  INV_X1 U5632 ( .A(EAX_REG_25__SCAN_IN), .ZN(n4576) );
  AOI22_X1 U5633 ( .A1(n5738), .A2(UWORD_REG_9__SCAN_IN), .B1(n5743), .B2(
        DATAO_REG_25__SCAN_IN), .ZN(n4575) );
  OAI21_X1 U5634 ( .B1(n4576), .B2(n5714), .A(n4575), .ZN(U2898) );
  INV_X1 U5635 ( .A(EAX_REG_20__SCAN_IN), .ZN(n4578) );
  AOI22_X1 U5636 ( .A1(n5738), .A2(UWORD_REG_4__SCAN_IN), .B1(n5743), .B2(
        DATAO_REG_20__SCAN_IN), .ZN(n4577) );
  OAI21_X1 U5637 ( .B1(n4578), .B2(n5714), .A(n4577), .ZN(U2903) );
  INV_X1 U5638 ( .A(EAX_REG_23__SCAN_IN), .ZN(n6880) );
  AOI22_X1 U5639 ( .A1(n5738), .A2(UWORD_REG_7__SCAN_IN), .B1(n5743), .B2(
        DATAO_REG_23__SCAN_IN), .ZN(n4579) );
  OAI21_X1 U5640 ( .B1(n6880), .B2(n5714), .A(n4579), .ZN(U2900) );
  INV_X1 U5641 ( .A(n4580), .ZN(n4583) );
  INV_X1 U5642 ( .A(n4581), .ZN(n4582) );
  AOI21_X1 U5643 ( .B1(n4583), .B2(n6605), .A(n4582), .ZN(n5775) );
  INV_X1 U5644 ( .A(n5775), .ZN(n4591) );
  AOI21_X1 U5645 ( .B1(n4585), .B2(n6605), .A(n4584), .ZN(n5689) );
  INV_X1 U5646 ( .A(REIP_REG_0__SCAN_IN), .ZN(n6622) );
  OAI21_X1 U5647 ( .B1(n5811), .B2(n6622), .A(n4586), .ZN(n4589) );
  AOI21_X1 U5648 ( .B1(n5527), .B2(n4587), .A(n6605), .ZN(n4588) );
  AOI211_X1 U5649 ( .C1(n5689), .C2(n5834), .A(n4589), .B(n4588), .ZN(n4590)
         );
  OAI21_X1 U5650 ( .B1(n4591), .B2(n5824), .A(n4590), .ZN(U3018) );
  INV_X1 U5651 ( .A(EAX_REG_22__SCAN_IN), .ZN(n4593) );
  AOI22_X1 U5652 ( .A1(n5738), .A2(UWORD_REG_6__SCAN_IN), .B1(n5743), .B2(
        DATAO_REG_22__SCAN_IN), .ZN(n4592) );
  OAI21_X1 U5653 ( .B1(n4593), .B2(n5714), .A(n4592), .ZN(U2901) );
  INV_X1 U5654 ( .A(EAX_REG_27__SCAN_IN), .ZN(n6902) );
  AOI22_X1 U5655 ( .A1(n5738), .A2(UWORD_REG_11__SCAN_IN), .B1(n5743), .B2(
        DATAO_REG_27__SCAN_IN), .ZN(n4594) );
  OAI21_X1 U5656 ( .B1(n6902), .B2(n5714), .A(n4594), .ZN(U2896) );
  INV_X1 U5657 ( .A(n4595), .ZN(n4598) );
  OAI21_X1 U5658 ( .B1(n4598), .B2(n4597), .A(n4596), .ZN(n5780) );
  OR2_X1 U5659 ( .A1(n4496), .A2(n3717), .ZN(n4600) );
  NOR2_X1 U5660 ( .A1(n4600), .A2(n4599), .ZN(n4601) );
  NAND2_X1 U5661 ( .A1(n4604), .A2(n5906), .ZN(n4605) );
  INV_X1 U5662 ( .A(n4605), .ZN(n4606) );
  INV_X1 U5663 ( .A(EAX_REG_0__SCAN_IN), .ZN(n5747) );
  OAI222_X1 U5664 ( .A1(n5780), .A2(n5468), .B1(n4951), .B2(n4535), .C1(n5164), 
        .C2(n5747), .ZN(U2891) );
  NOR2_X1 U5665 ( .A1(n4608), .A2(n4607), .ZN(n4609) );
  INV_X1 U5666 ( .A(EAX_REG_1__SCAN_IN), .ZN(n5745) );
  OAI222_X1 U5667 ( .A1(n4789), .A2(n5468), .B1(n4951), .B2(n4537), .C1(n5164), 
        .C2(n5745), .ZN(U2890) );
  INV_X1 U5668 ( .A(n5689), .ZN(n4611) );
  OAI222_X1 U5669 ( .A1(n4611), .A2(n5156), .B1(n4123), .B2(n5706), .C1(n5780), 
        .C2(n5162), .ZN(U2859) );
  XNOR2_X1 U5670 ( .A(n5675), .B(n4178), .ZN(n5847) );
  OAI222_X1 U5671 ( .A1(n4789), .A2(n5162), .B1(n3180), .B2(n5706), .C1(n5156), 
        .C2(n5847), .ZN(U2858) );
  AOI22_X1 U5672 ( .A1(n5760), .A2(LWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_9__SCAN_IN), .B2(n5756), .ZN(n4613) );
  INV_X1 U5673 ( .A(DATAI_9_), .ZN(n4811) );
  OR2_X1 U5674 ( .A1(n4641), .A2(n4811), .ZN(n4616) );
  NAND2_X1 U5675 ( .A1(n4613), .A2(n4616), .ZN(U2948) );
  AOI22_X1 U5676 ( .A1(n5760), .A2(LWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_11__SCAN_IN), .B2(n5756), .ZN(n4614) );
  INV_X1 U5677 ( .A(DATAI_11_), .ZN(n4873) );
  OR2_X1 U5678 ( .A1(n4641), .A2(n4873), .ZN(n4620) );
  NAND2_X1 U5679 ( .A1(n4614), .A2(n4620), .ZN(U2950) );
  AOI22_X1 U5680 ( .A1(n5760), .A2(LWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_13__SCAN_IN), .B2(n5756), .ZN(n4615) );
  INV_X1 U5681 ( .A(DATAI_13_), .ZN(n4950) );
  OR2_X1 U5682 ( .A1(n4641), .A2(n4950), .ZN(n4618) );
  NAND2_X1 U5683 ( .A1(n4615), .A2(n4618), .ZN(U2952) );
  AOI22_X1 U5684 ( .A1(n5760), .A2(UWORD_REG_9__SCAN_IN), .B1(
        EAX_REG_25__SCAN_IN), .B2(n5756), .ZN(n4617) );
  NAND2_X1 U5685 ( .A1(n4617), .A2(n4616), .ZN(U2933) );
  AOI22_X1 U5686 ( .A1(n5760), .A2(UWORD_REG_13__SCAN_IN), .B1(
        EAX_REG_29__SCAN_IN), .B2(n5756), .ZN(n4619) );
  NAND2_X1 U5687 ( .A1(n4619), .A2(n4618), .ZN(U2937) );
  AOI22_X1 U5688 ( .A1(n5760), .A2(UWORD_REG_11__SCAN_IN), .B1(
        EAX_REG_27__SCAN_IN), .B2(n5756), .ZN(n4621) );
  NAND2_X1 U5689 ( .A1(n4621), .A2(n4620), .ZN(U2935) );
  AOI22_X1 U5690 ( .A1(n5760), .A2(LWORD_REG_4__SCAN_IN), .B1(
        EAX_REG_4__SCAN_IN), .B2(n5756), .ZN(n4623) );
  NAND2_X1 U5691 ( .A1(n4623), .A2(n4622), .ZN(U2943) );
  AOI22_X1 U5692 ( .A1(n5760), .A2(UWORD_REG_7__SCAN_IN), .B1(
        EAX_REG_23__SCAN_IN), .B2(n5756), .ZN(n4625) );
  NAND2_X1 U5693 ( .A1(n4625), .A2(n4624), .ZN(U2931) );
  AOI22_X1 U5694 ( .A1(n5760), .A2(UWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_18__SCAN_IN), .B2(n5756), .ZN(n4626) );
  NAND2_X1 U5695 ( .A1(n5759), .A2(DATAI_2_), .ZN(n4633) );
  NAND2_X1 U5696 ( .A1(n4626), .A2(n4633), .ZN(U2926) );
  AOI22_X1 U5697 ( .A1(n5760), .A2(UWORD_REG_12__SCAN_IN), .B1(
        EAX_REG_28__SCAN_IN), .B2(n5756), .ZN(n4628) );
  NAND2_X1 U5698 ( .A1(n4628), .A2(n4627), .ZN(U2936) );
  AOI22_X1 U5699 ( .A1(n5760), .A2(LWORD_REG_5__SCAN_IN), .B1(
        EAX_REG_5__SCAN_IN), .B2(n5756), .ZN(n4630) );
  NAND2_X1 U5700 ( .A1(n4630), .A2(n4629), .ZN(U2944) );
  AOI22_X1 U5701 ( .A1(n5760), .A2(UWORD_REG_14__SCAN_IN), .B1(
        EAX_REG_30__SCAN_IN), .B2(n5756), .ZN(n4632) );
  NAND2_X1 U5702 ( .A1(n4632), .A2(n4631), .ZN(U2938) );
  AOI22_X1 U5703 ( .A1(n5760), .A2(LWORD_REG_2__SCAN_IN), .B1(
        EAX_REG_2__SCAN_IN), .B2(n5756), .ZN(n4634) );
  NAND2_X1 U5704 ( .A1(n4634), .A2(n4633), .ZN(U2941) );
  AOI22_X1 U5705 ( .A1(n5760), .A2(LWORD_REG_6__SCAN_IN), .B1(
        EAX_REG_6__SCAN_IN), .B2(n5756), .ZN(n4636) );
  NAND2_X1 U5706 ( .A1(n4636), .A2(n4635), .ZN(U2945) );
  AOI22_X1 U5707 ( .A1(n5760), .A2(LWORD_REG_3__SCAN_IN), .B1(
        EAX_REG_3__SCAN_IN), .B2(n5756), .ZN(n4638) );
  NAND2_X1 U5708 ( .A1(n4638), .A2(n4637), .ZN(U2942) );
  AOI22_X1 U5709 ( .A1(n5760), .A2(LWORD_REG_0__SCAN_IN), .B1(
        EAX_REG_0__SCAN_IN), .B2(n5756), .ZN(n4639) );
  OAI21_X1 U5710 ( .B1(n4535), .B2(n4641), .A(n4639), .ZN(U2939) );
  AOI22_X1 U5711 ( .A1(n5760), .A2(LWORD_REG_1__SCAN_IN), .B1(
        EAX_REG_1__SCAN_IN), .B2(n5756), .ZN(n4640) );
  OAI21_X1 U5712 ( .B1(n4537), .B2(n4641), .A(n4640), .ZN(U2940) );
  OR2_X1 U5713 ( .A1(n4643), .A2(n4644), .ZN(n4645) );
  NAND2_X1 U5714 ( .A1(n4642), .A2(n4645), .ZN(n5669) );
  INV_X1 U5715 ( .A(EBX_REG_3__SCAN_IN), .ZN(n6863) );
  NAND2_X1 U5716 ( .A1(n4826), .A2(n4646), .ZN(n4647) );
  NAND2_X1 U5717 ( .A1(n4698), .A2(n4647), .ZN(n5822) );
  OAI222_X1 U5718 ( .A1(n5669), .A2(n5162), .B1(n5706), .B2(n6863), .C1(n5822), 
        .C2(n5156), .ZN(U2856) );
  INV_X1 U5719 ( .A(DATAI_3_), .ZN(n5887) );
  INV_X1 U5720 ( .A(EAX_REG_3__SCAN_IN), .ZN(n6835) );
  OAI222_X1 U5721 ( .A1(n5669), .A2(n5468), .B1(n4951), .B2(n5887), .C1(n5164), 
        .C2(n6835), .ZN(U2888) );
  NOR2_X1 U5722 ( .A1(n3099), .A2(n4648), .ZN(n4650) );
  NOR2_X1 U5723 ( .A1(n4643), .A2(n4650), .ZN(n5769) );
  INV_X1 U5724 ( .A(n5769), .ZN(n4834) );
  INV_X1 U5725 ( .A(DATAI_2_), .ZN(n5882) );
  INV_X1 U5726 ( .A(EAX_REG_2__SCAN_IN), .ZN(n5742) );
  OAI222_X1 U5727 ( .A1(n4834), .A2(n5468), .B1(n4951), .B2(n5882), .C1(n5164), 
        .C2(n5742), .ZN(U2889) );
  INV_X1 U5728 ( .A(n3119), .ZN(n4686) );
  NAND2_X1 U5729 ( .A1(n4653), .A2(n4652), .ZN(n4669) );
  XNOR2_X1 U5730 ( .A(n4550), .B(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4656)
         );
  XNOR2_X1 U5731 ( .A(INSTQUEUERD_ADDR_REG_1__SCAN_IN), .B(
        INSTQUEUERD_ADDR_REG_2__SCAN_IN), .ZN(n4654) );
  OAI22_X1 U5732 ( .A1(n6478), .A2(n4654), .B1(n4665), .B2(n4656), .ZN(n4655)
         );
  AOI21_X1 U5733 ( .B1(n4669), .B2(n4656), .A(n4655), .ZN(n4657) );
  OAI21_X1 U5734 ( .B1(n4686), .B2(n6476), .A(n4657), .ZN(n5014) );
  NAND2_X1 U5735 ( .A1(n4676), .A2(n3258), .ZN(n4658) );
  OAI21_X1 U5736 ( .B1(n5014), .B2(n4676), .A(n4658), .ZN(n6486) );
  NOR2_X1 U5737 ( .A1(n6486), .A2(STATE2_REG_1__SCAN_IN), .ZN(n4673) );
  NAND2_X1 U5738 ( .A1(n6211), .A2(n4659), .ZN(n4671) );
  MUX2_X1 U5739 ( .A(n3268), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4550), 
        .Z(n4661) );
  NOR2_X1 U5740 ( .A1(n4661), .A2(n4660), .ZN(n4668) );
  NAND2_X1 U5741 ( .A1(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A2(
        INSTQUEUERD_ADDR_REG_1__SCAN_IN), .ZN(n4663) );
  INV_X1 U5742 ( .A(n4663), .ZN(n4662) );
  MUX2_X1 U5743 ( .A(n4663), .B(n4662), .S(INSTQUEUERD_ADDR_REG_3__SCAN_IN), 
        .Z(n4666) );
  AOI21_X1 U5744 ( .B1(n4550), .B2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A(n3777), 
        .ZN(n4664) );
  NOR2_X1 U5745 ( .A1(n3114), .A2(n4664), .ZN(n6602) );
  OAI22_X1 U5746 ( .A1(n6478), .A2(n4666), .B1(n6602), .B2(n4665), .ZN(n4667)
         );
  AOI21_X1 U5747 ( .B1(n4669), .B2(n4668), .A(n4667), .ZN(n4670) );
  NAND2_X1 U5748 ( .A1(n4671), .A2(n4670), .ZN(n6600) );
  MUX2_X1 U5749 ( .A(n6600), .B(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .S(n4676), 
        .Z(n6494) );
  NAND2_X1 U5750 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n5558), .ZN(n4677) );
  INV_X1 U5751 ( .A(n4677), .ZN(n4672) );
  AOI22_X1 U5752 ( .A1(n4673), .A2(n6494), .B1(n4660), .B2(n4672), .ZN(n6504)
         );
  NOR2_X1 U5753 ( .A1(n6504), .A2(n4549), .ZN(n4682) );
  INV_X1 U5754 ( .A(n6020), .ZN(n6082) );
  NOR2_X1 U5755 ( .A1(n4674), .A2(n6082), .ZN(n4675) );
  XOR2_X1 U5756 ( .A(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B(n4675), .Z(n5655) );
  AOI22_X1 U5757 ( .A1(n5655), .A2(n5547), .B1(INSTQUEUERD_ADDR_REG_4__SCAN_IN), .B2(n4676), .ZN(n4678) );
  OAI22_X1 U5758 ( .A1(n4678), .A2(STATE2_REG_1__SCAN_IN), .B1(n4677), .B2(
        n5548), .ZN(n6502) );
  NOR3_X1 U5759 ( .A1(n4682), .A2(n6502), .A3(FLUSH_REG_SCAN_IN), .ZN(n4679)
         );
  INV_X1 U5760 ( .A(n4680), .ZN(n4681) );
  OR3_X1 U5761 ( .A1(n4682), .A2(n6502), .A3(n4681), .ZN(n6520) );
  INV_X1 U5762 ( .A(n6520), .ZN(n4684) );
  INV_X1 U5763 ( .A(n6179), .ZN(n6477) );
  NAND2_X1 U5764 ( .A1(STATE2_REG_1__SCAN_IN), .A2(n6598), .ZN(n5400) );
  INV_X1 U5765 ( .A(n5400), .ZN(n5396) );
  OAI22_X1 U5766 ( .A1(n5952), .A2(n6410), .B1(n6477), .B2(n5396), .ZN(n4683)
         );
  OAI21_X1 U5767 ( .B1(n4684), .B2(n4683), .A(n5860), .ZN(n4685) );
  OAI21_X1 U5768 ( .B1(n5860), .B2(n6316), .A(n4685), .ZN(U3465) );
  INV_X1 U5769 ( .A(n5860), .ZN(n4692) );
  NAND2_X1 U5770 ( .A1(n4688), .A2(STATEBS16_REG_SCAN_IN), .ZN(n6247) );
  OAI21_X1 U5771 ( .B1(n6149), .B2(n6247), .A(n6419), .ZN(n5402) );
  AOI21_X1 U5772 ( .B1(n6149), .B2(n6247), .A(n5402), .ZN(n4689) );
  AOI21_X1 U5773 ( .B1(n5400), .B2(n3119), .A(n4689), .ZN(n4691) );
  NAND2_X1 U5774 ( .A1(n4692), .A2(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .ZN(n4690) );
  OAI21_X1 U5775 ( .B1(n4692), .B2(n4691), .A(n4690), .ZN(U3463) );
  AOI21_X1 U5776 ( .B1(n4695), .B2(n4642), .A(n4694), .ZN(n5658) );
  INV_X1 U5777 ( .A(n5658), .ZN(n4701) );
  AOI22_X1 U5778 ( .A1(n4956), .A2(DATAI_4_), .B1(n5710), .B2(
        EAX_REG_4__SCAN_IN), .ZN(n4696) );
  OAI21_X1 U5779 ( .B1(n4701), .B2(n5468), .A(n4696), .ZN(U2887) );
  INV_X1 U5780 ( .A(EBX_REG_4__SCAN_IN), .ZN(n4700) );
  AND2_X1 U5781 ( .A1(n4698), .A2(n4697), .ZN(n4699) );
  OR2_X1 U5782 ( .A1(n4699), .A2(n4706), .ZN(n5812) );
  OAI222_X1 U5783 ( .A1(n4701), .A2(n5162), .B1(n4700), .B2(n5706), .C1(n5156), 
        .C2(n5812), .ZN(U2855) );
  INV_X1 U5784 ( .A(n4702), .ZN(n4703) );
  OAI21_X1 U5785 ( .B1(n4694), .B2(n4704), .A(n4703), .ZN(n5643) );
  OR2_X1 U5786 ( .A1(n4706), .A2(n4705), .ZN(n4707) );
  NAND2_X1 U5787 ( .A1(n4714), .A2(n4707), .ZN(n5641) );
  INV_X1 U5788 ( .A(n5641), .ZN(n4708) );
  AOI22_X1 U5789 ( .A1(n4502), .A2(n4708), .B1(EBX_REG_5__SCAN_IN), .B2(n5145), 
        .ZN(n4709) );
  OAI21_X1 U5790 ( .B1(n5643), .B2(n5162), .A(n4709), .ZN(U2854) );
  OAI21_X1 U5791 ( .B1(n4702), .B2(n4712), .A(n4711), .ZN(n5629) );
  INV_X1 U5792 ( .A(n4736), .ZN(n4713) );
  AOI21_X1 U5793 ( .B1(n4715), .B2(n4714), .A(n4713), .ZN(n5803) );
  AOI22_X1 U5794 ( .A1(n5803), .A2(n4502), .B1(EBX_REG_6__SCAN_IN), .B2(n5145), 
        .ZN(n4716) );
  OAI21_X1 U5795 ( .B1(n5629), .B2(n5162), .A(n4716), .ZN(U2853) );
  INV_X1 U5796 ( .A(DATAI_5_), .ZN(n6785) );
  INV_X1 U5797 ( .A(EAX_REG_5__SCAN_IN), .ZN(n5736) );
  OAI222_X1 U5798 ( .A1(n5643), .A2(n5468), .B1(n4951), .B2(n6785), .C1(n5164), 
        .C2(n5736), .ZN(U2886) );
  INV_X1 U5799 ( .A(DATAI_6_), .ZN(n5901) );
  OAI222_X1 U5800 ( .A1(n5629), .A2(n5468), .B1(n4951), .B2(n5901), .C1(n5164), 
        .C2(n3808), .ZN(U2885) );
  NAND2_X1 U5801 ( .A1(n5836), .A2(n5841), .ZN(n4738) );
  INV_X1 U5802 ( .A(n4738), .ZN(n4719) );
  INV_X1 U5803 ( .A(n4717), .ZN(n4718) );
  AOI211_X1 U5804 ( .C1(n5818), .C2(n4719), .A(INSTADDRPOINTER_REG_5__SCAN_IN), 
        .B(n4718), .ZN(n4730) );
  AND2_X1 U5805 ( .A1(INSTADDRPOINTER_REG_5__SCAN_IN), .A2(n4739), .ZN(n4720)
         );
  OR2_X1 U5806 ( .A1(n5852), .A2(n4720), .ZN(n4724) );
  OR2_X1 U5807 ( .A1(n4898), .A2(n5836), .ZN(n4723) );
  INV_X1 U5808 ( .A(n5859), .ZN(n4721) );
  NAND2_X1 U5809 ( .A1(n4903), .A2(n4721), .ZN(n4722) );
  AND2_X1 U5810 ( .A1(n4723), .A2(n4722), .ZN(n5810) );
  AND2_X1 U5811 ( .A1(n4724), .A2(n5810), .ZN(n5809) );
  XOR2_X1 U5812 ( .A(n4726), .B(n4725), .Z(n4780) );
  NAND2_X1 U5813 ( .A1(n4780), .A2(n5854), .ZN(n4729) );
  NAND2_X1 U5814 ( .A1(n5262), .A2(REIP_REG_5__SCAN_IN), .ZN(n4781) );
  OAI21_X1 U5815 ( .B1(n5848), .B2(n5641), .A(n4781), .ZN(n4727) );
  INV_X1 U5816 ( .A(n4727), .ZN(n4728) );
  OAI211_X1 U5817 ( .C1(n4730), .C2(n5809), .A(n4729), .B(n4728), .ZN(U3013)
         );
  XNOR2_X1 U5818 ( .A(n4731), .B(n4732), .ZN(n4767) );
  OAI22_X1 U5819 ( .A1(n4898), .A2(n4734), .B1(n5356), .B2(n4733), .ZN(n4840)
         );
  AND2_X1 U5820 ( .A1(n4736), .A2(n4735), .ZN(n4737) );
  OR2_X1 U5821 ( .A1(n4737), .A2(n4777), .ZN(n5613) );
  NAND2_X1 U5822 ( .A1(n5832), .A2(REIP_REG_7__SCAN_IN), .ZN(n4762) );
  NAND2_X1 U5823 ( .A1(n4903), .A2(n4738), .ZN(n5819) );
  NAND3_X1 U5824 ( .A1(n4739), .A2(INSTADDRPOINTER_REG_5__SCAN_IN), .A3(n5819), 
        .ZN(n5805) );
  NOR2_X1 U5825 ( .A1(n3655), .A2(n5805), .ZN(n5800) );
  NAND2_X1 U5826 ( .A1(n4139), .A2(n5800), .ZN(n4740) );
  OAI211_X1 U5827 ( .C1(n5613), .C2(n5848), .A(n4762), .B(n4740), .ZN(n4741)
         );
  AOI21_X1 U5828 ( .B1(n4840), .B2(INSTADDRPOINTER_REG_7__SCAN_IN), .A(n4741), 
        .ZN(n4742) );
  OAI21_X1 U5829 ( .B1(n4767), .B2(n5824), .A(n4742), .ZN(U3011) );
  NAND2_X1 U5830 ( .A1(n4711), .A2(n4744), .ZN(n4745) );
  AND2_X1 U5831 ( .A1(n4743), .A2(n4745), .ZN(n4765) );
  OAI22_X1 U5832 ( .A1(n5613), .A2(n5156), .B1(n5625), .B2(n5706), .ZN(n4746)
         );
  AOI21_X1 U5833 ( .B1(n4765), .B2(n5703), .A(n4746), .ZN(n4747) );
  INV_X1 U5834 ( .A(n4747), .ZN(U2852) );
  INV_X1 U5835 ( .A(n4765), .ZN(n5621) );
  INV_X1 U5836 ( .A(DATAI_7_), .ZN(n6731) );
  INV_X1 U5837 ( .A(EAX_REG_7__SCAN_IN), .ZN(n4748) );
  OAI222_X1 U5838 ( .A1(n5621), .A2(n5468), .B1(n4951), .B2(n6731), .C1(n5164), 
        .C2(n4748), .ZN(U2884) );
  XNOR2_X1 U5839 ( .A(n4750), .B(n4749), .ZN(n5825) );
  INV_X1 U5840 ( .A(n5669), .ZN(n4754) );
  NAND2_X1 U5841 ( .A1(n5832), .A2(REIP_REG_3__SCAN_IN), .ZN(n5821) );
  INV_X1 U5842 ( .A(n5821), .ZN(n4751) );
  AOI21_X1 U5843 ( .B1(n5777), .B2(PHYADDRPOINTER_REG_3__SCAN_IN), .A(n4751), 
        .ZN(n4752) );
  OAI21_X1 U5844 ( .B1(n5773), .B2(n5664), .A(n4752), .ZN(n4753) );
  AOI21_X1 U5845 ( .B1(n4754), .B2(n5768), .A(n4753), .ZN(n4755) );
  OAI21_X1 U5846 ( .B1(n5825), .B2(n5557), .A(n4755), .ZN(U2983) );
  XOR2_X1 U5847 ( .A(n4756), .B(n4757), .Z(n5815) );
  INV_X1 U5848 ( .A(n5815), .ZN(n4761) );
  AOI22_X1 U5849 ( .A1(n5777), .A2(PHYADDRPOINTER_REG_4__SCAN_IN), .B1(n5262), 
        .B2(REIP_REG_4__SCAN_IN), .ZN(n4758) );
  OAI21_X1 U5850 ( .B1(n5773), .B2(n5661), .A(n4758), .ZN(n4759) );
  AOI21_X1 U5851 ( .B1(n5658), .B2(n5768), .A(n4759), .ZN(n4760) );
  OAI21_X1 U5852 ( .B1(n4761), .B2(n5557), .A(n4760), .ZN(U2982) );
  NAND2_X1 U5853 ( .A1(n5777), .A2(PHYADDRPOINTER_REG_7__SCAN_IN), .ZN(n4763)
         );
  OAI211_X1 U5854 ( .C1(n5773), .C2(n5619), .A(n4763), .B(n4762), .ZN(n4764)
         );
  AOI21_X1 U5855 ( .B1(n4765), .B2(n5768), .A(n4764), .ZN(n4766) );
  OAI21_X1 U5856 ( .B1(n4767), .B2(n5557), .A(n4766), .ZN(U2979) );
  XOR2_X1 U5857 ( .A(n4768), .B(n4769), .Z(n5807) );
  NAND2_X1 U5858 ( .A1(n5807), .A2(n5774), .ZN(n4772) );
  OAI22_X1 U5859 ( .A1(n5248), .A2(n3813), .B1(n5811), .B2(n6557), .ZN(n4770)
         );
  AOI21_X1 U5860 ( .B1(n5630), .B2(n5250), .A(n4770), .ZN(n4771) );
  OAI211_X1 U5861 ( .C1(n5911), .C2(n5629), .A(n4772), .B(n4771), .ZN(U2980)
         );
  AOI21_X1 U5862 ( .B1(n4774), .B2(n4743), .A(n4773), .ZN(n4798) );
  INV_X1 U5863 ( .A(n4798), .ZN(n5105) );
  AOI22_X1 U5864 ( .A1(n4956), .A2(DATAI_8_), .B1(n5710), .B2(
        EAX_REG_8__SCAN_IN), .ZN(n4775) );
  OAI21_X1 U5865 ( .B1(n5105), .B2(n5468), .A(n4775), .ZN(U2883) );
  INV_X1 U5866 ( .A(EBX_REG_8__SCAN_IN), .ZN(n4779) );
  NOR2_X1 U5867 ( .A1(n4777), .A2(n4776), .ZN(n4778) );
  OR2_X1 U5868 ( .A1(n4847), .A2(n4778), .ZN(n5795) );
  OAI222_X1 U5869 ( .A1(n5105), .A2(n5162), .B1(n5706), .B2(n4779), .C1(n5795), 
        .C2(n5156), .ZN(U2851) );
  NAND2_X1 U5870 ( .A1(n4780), .A2(n5774), .ZN(n4785) );
  INV_X1 U5871 ( .A(n4781), .ZN(n4783) );
  NOR2_X1 U5872 ( .A1(n5773), .A2(n5642), .ZN(n4782) );
  AOI211_X1 U5873 ( .C1(n5777), .C2(PHYADDRPOINTER_REG_5__SCAN_IN), .A(n4783), 
        .B(n4782), .ZN(n4784) );
  OAI211_X1 U5874 ( .C1(n5911), .C2(n5643), .A(n4785), .B(n4784), .ZN(U2981)
         );
  OAI21_X1 U5875 ( .B1(n4788), .B2(n4787), .A(n4786), .ZN(n5850) );
  INV_X1 U5876 ( .A(n4789), .ZN(n5684) );
  INV_X1 U5877 ( .A(PHYADDRPOINTER_REG_1__SCAN_IN), .ZN(n5676) );
  NAND2_X1 U5878 ( .A1(n5250), .A2(n5676), .ZN(n4790) );
  NAND2_X1 U5879 ( .A1(n5832), .A2(REIP_REG_1__SCAN_IN), .ZN(n5846) );
  OAI211_X1 U5880 ( .C1(n5248), .C2(n5676), .A(n4790), .B(n5846), .ZN(n4791)
         );
  AOI21_X1 U5881 ( .B1(n5684), .B2(n5768), .A(n4791), .ZN(n4792) );
  OAI21_X1 U5882 ( .B1(n5557), .B2(n5850), .A(n4792), .ZN(U2985) );
  XOR2_X1 U5883 ( .A(n4793), .B(n4794), .Z(n5798) );
  INV_X1 U5884 ( .A(n5798), .ZN(n4800) );
  INV_X1 U5885 ( .A(n4795), .ZN(n5100) );
  AOI22_X1 U5886 ( .A1(n5777), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .B1(n5262), 
        .B2(REIP_REG_8__SCAN_IN), .ZN(n4796) );
  OAI21_X1 U5887 ( .B1(n5773), .B2(n5100), .A(n4796), .ZN(n4797) );
  AOI21_X1 U5888 ( .B1(n4798), .B2(n5768), .A(n4797), .ZN(n4799) );
  OAI21_X1 U5889 ( .B1(n4800), .B2(n5557), .A(n4799), .ZN(U2978) );
  INV_X1 U5890 ( .A(n4801), .ZN(n4802) );
  OAI21_X1 U5891 ( .B1(n4773), .B2(n4803), .A(n4802), .ZN(n5096) );
  XNOR2_X1 U5892 ( .A(n5245), .B(n6751), .ZN(n4805) );
  XNOR2_X1 U5893 ( .A(n4804), .B(n4805), .ZN(n5790) );
  NAND2_X1 U5894 ( .A1(n5790), .A2(n5774), .ZN(n4809) );
  INV_X1 U5895 ( .A(REIP_REG_9__SCAN_IN), .ZN(n4806) );
  NOR2_X1 U5896 ( .A1(n5811), .A2(n4806), .ZN(n5787) );
  NOR2_X1 U5897 ( .A1(n5773), .A2(n5087), .ZN(n4807) );
  AOI211_X1 U5898 ( .C1(n5777), .C2(PHYADDRPOINTER_REG_9__SCAN_IN), .A(n5787), 
        .B(n4807), .ZN(n4808) );
  OAI211_X1 U5899 ( .C1(n5911), .C2(n5096), .A(n4809), .B(n4808), .ZN(U2977)
         );
  INV_X1 U5900 ( .A(EBX_REG_9__SCAN_IN), .ZN(n4810) );
  XNOR2_X1 U5901 ( .A(n4847), .B(n4846), .ZN(n5086) );
  OAI222_X1 U5902 ( .A1(n5096), .A2(n5162), .B1(n4810), .B2(n5706), .C1(n5156), 
        .C2(n5086), .ZN(U2850) );
  INV_X1 U5903 ( .A(EAX_REG_9__SCAN_IN), .ZN(n6692) );
  OAI222_X1 U5904 ( .A1(n5096), .A2(n5468), .B1(n4951), .B2(n4811), .C1(n5164), 
        .C2(n6692), .ZN(U2882) );
  NAND2_X1 U5905 ( .A1(n4819), .A2(n4812), .ZN(n4813) );
  OR2_X1 U5906 ( .A1(n5653), .A2(REIP_REG_1__SCAN_IN), .ZN(n5678) );
  NAND2_X1 U5907 ( .A1(n5678), .A2(n5687), .ZN(n5662) );
  NAND3_X1 U5908 ( .A1(n3407), .A2(n6734), .A3(n4814), .ZN(n4815) );
  NAND2_X1 U5909 ( .A1(n4816), .A2(n4815), .ZN(n4817) );
  AND2_X1 U5910 ( .A1(n4819), .A2(n4818), .ZN(n5694) );
  AOI22_X1 U5911 ( .A1(EBX_REG_2__SCAN_IN), .A2(n5693), .B1(n5694), .B2(n3119), 
        .ZN(n4831) );
  INV_X1 U5912 ( .A(n5772), .ZN(n4822) );
  AOI22_X1 U5913 ( .A1(n4822), .A2(n5677), .B1(n5674), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n4830) );
  INV_X1 U5914 ( .A(n5653), .ZN(n5098) );
  INV_X1 U5915 ( .A(REIP_REG_2__SCAN_IN), .ZN(n4823) );
  NAND3_X1 U5916 ( .A1(n5098), .A2(REIP_REG_1__SCAN_IN), .A3(n4823), .ZN(n4829) );
  OR2_X1 U5917 ( .A1(n4825), .A2(n4824), .ZN(n4827) );
  AND2_X1 U5918 ( .A1(n4827), .A2(n4826), .ZN(n5833) );
  NAND2_X1 U5919 ( .A1(n5690), .A2(n5833), .ZN(n4828) );
  NAND4_X1 U5920 ( .A1(n4831), .A2(n4830), .A3(n4829), .A4(n4828), .ZN(n4832)
         );
  AOI21_X1 U5921 ( .B1(REIP_REG_2__SCAN_IN), .B2(n5662), .A(n4832), .ZN(n4833)
         );
  OAI21_X1 U5922 ( .B1(n4834), .B2(n5698), .A(n4833), .ZN(U2825) );
  INV_X1 U5923 ( .A(n4836), .ZN(n4838) );
  NAND2_X1 U5924 ( .A1(n4838), .A2(n4837), .ZN(n4839) );
  XNOR2_X1 U5925 ( .A(n4835), .B(n4839), .ZN(n4861) );
  INV_X1 U5926 ( .A(n4840), .ZN(n5794) );
  OAI21_X1 U5927 ( .B1(n5852), .B2(n4841), .A(n5794), .ZN(n5789) );
  NAND2_X1 U5928 ( .A1(n4841), .A2(n5800), .ZN(n5793) );
  AOI21_X1 U5929 ( .B1(n6751), .B2(n4842), .A(n5793), .ZN(n4844) );
  AOI22_X1 U5930 ( .A1(INSTADDRPOINTER_REG_10__SCAN_IN), .A2(n5789), .B1(n4844), .B2(n4843), .ZN(n4851) );
  AOI21_X1 U5931 ( .B1(n4847), .B2(n4846), .A(n4845), .ZN(n4848) );
  NOR2_X1 U5932 ( .A1(n3138), .A2(n4848), .ZN(n5699) );
  INV_X1 U5933 ( .A(REIP_REG_10__SCAN_IN), .ZN(n4849) );
  NOR2_X1 U5934 ( .A1(n5811), .A2(n4849), .ZN(n4858) );
  AOI21_X1 U5935 ( .B1(n5699), .B2(n5834), .A(n4858), .ZN(n4850) );
  OAI211_X1 U5936 ( .C1(n4861), .C2(n5824), .A(n4851), .B(n4850), .ZN(U3008)
         );
  OR2_X1 U5937 ( .A1(n4801), .A2(n4853), .ZN(n4854) );
  AND2_X1 U5938 ( .A1(n4852), .A2(n4854), .ZN(n5700) );
  INV_X1 U5939 ( .A(n5700), .ZN(n4856) );
  AOI22_X1 U5940 ( .A1(n4956), .A2(DATAI_10_), .B1(n5710), .B2(
        EAX_REG_10__SCAN_IN), .ZN(n4855) );
  OAI21_X1 U5941 ( .B1(n4856), .B2(n5468), .A(n4855), .ZN(U2881) );
  AND2_X1 U5942 ( .A1(n5777), .A2(PHYADDRPOINTER_REG_10__SCAN_IN), .ZN(n4857)
         );
  AOI211_X1 U5943 ( .C1(n5250), .C2(n5606), .A(n4858), .B(n4857), .ZN(n4860)
         );
  NAND2_X1 U5944 ( .A1(n5700), .A2(n5768), .ZN(n4859) );
  OAI211_X1 U5945 ( .C1(n4861), .C2(n5557), .A(n4860), .B(n4859), .ZN(U2976)
         );
  NAND2_X1 U5946 ( .A1(n4852), .A2(n4863), .ZN(n4864) );
  NAND2_X1 U5947 ( .A1(n4862), .A2(n4864), .ZN(n4890) );
  INV_X1 U5948 ( .A(n4865), .ZN(n4887) );
  OAI21_X1 U5949 ( .B1(n3138), .B2(n3139), .A(n4877), .ZN(n5781) );
  NAND2_X1 U5950 ( .A1(n4866), .A2(n5687), .ZN(n5640) );
  NAND2_X1 U5951 ( .A1(n5688), .A2(n4867), .ZN(n5601) );
  OAI22_X1 U5952 ( .A1(n4885), .A2(n5692), .B1(n4884), .B2(n5601), .ZN(n4868)
         );
  AOI211_X1 U5953 ( .C1(n5693), .C2(EBX_REG_11__SCAN_IN), .A(n5651), .B(n4868), 
        .ZN(n4870) );
  NAND4_X1 U5954 ( .A1(n5608), .A2(REIP_REG_9__SCAN_IN), .A3(
        REIP_REG_10__SCAN_IN), .A4(n4884), .ZN(n4869) );
  OAI211_X1 U5955 ( .C1(n5781), .C2(n5681), .A(n4870), .B(n4869), .ZN(n4871)
         );
  AOI21_X1 U5956 ( .B1(n5677), .B2(n4887), .A(n4871), .ZN(n4872) );
  OAI21_X1 U5957 ( .B1(n4890), .B2(n5620), .A(n4872), .ZN(U2816) );
  INV_X1 U5958 ( .A(EAX_REG_11__SCAN_IN), .ZN(n6757) );
  OAI222_X1 U5959 ( .A1(n4890), .A2(n5468), .B1(n4951), .B2(n4873), .C1(n5164), 
        .C2(n6757), .ZN(U2880) );
  INV_X1 U5960 ( .A(EBX_REG_11__SCAN_IN), .ZN(n4874) );
  OAI222_X1 U5961 ( .A1(n4890), .A2(n5162), .B1(n5706), .B2(n4874), .C1(n5781), 
        .C2(n5156), .ZN(U2848) );
  AOI21_X1 U5962 ( .B1(n4876), .B2(n4862), .A(n4875), .ZN(n4896) );
  INV_X1 U5963 ( .A(n4896), .ZN(n5597) );
  INV_X1 U5964 ( .A(n4912), .ZN(n4929) );
  AOI21_X1 U5965 ( .B1(n4878), .B2(n4877), .A(n4929), .ZN(n5594) );
  AOI22_X1 U5966 ( .A1(n5594), .A2(n4502), .B1(EBX_REG_12__SCAN_IN), .B2(n5145), .ZN(n4879) );
  OAI21_X1 U5967 ( .B1(n5597), .B2(n5162), .A(n4879), .ZN(U2847) );
  INV_X1 U5968 ( .A(DATAI_12_), .ZN(n6737) );
  INV_X1 U5969 ( .A(EAX_REG_12__SCAN_IN), .ZN(n5729) );
  OAI222_X1 U5970 ( .A1(n5597), .A2(n5468), .B1(n4951), .B2(n6737), .C1(n5164), 
        .C2(n5729), .ZN(U2879) );
  NAND2_X1 U5971 ( .A1(n4882), .A2(n4881), .ZN(n4883) );
  XNOR2_X1 U5972 ( .A(n4880), .B(n4883), .ZN(n5783) );
  NAND2_X1 U5973 ( .A1(n5783), .A2(n5774), .ZN(n4889) );
  INV_X1 U5974 ( .A(REIP_REG_11__SCAN_IN), .ZN(n4884) );
  OAI22_X1 U5975 ( .A1(n5248), .A2(n4885), .B1(n5811), .B2(n4884), .ZN(n4886)
         );
  AOI21_X1 U5976 ( .B1(n5250), .B2(n4887), .A(n4886), .ZN(n4888) );
  OAI211_X1 U5977 ( .C1(n5911), .C2(n4890), .A(n4889), .B(n4888), .ZN(U2975)
         );
  XNOR2_X1 U5978 ( .A(n5245), .B(INSTADDRPOINTER_REG_12__SCAN_IN), .ZN(n4892)
         );
  XNOR2_X1 U5979 ( .A(n4891), .B(n4892), .ZN(n4909) );
  NOR2_X1 U5980 ( .A1(n5811), .A2(n6560), .ZN(n4906) );
  AOI21_X1 U5981 ( .B1(n5777), .B2(PHYADDRPOINTER_REG_12__SCAN_IN), .A(n4906), 
        .ZN(n4893) );
  OAI21_X1 U5982 ( .B1(n5773), .B2(n4894), .A(n4893), .ZN(n4895) );
  AOI21_X1 U5983 ( .B1(n4896), .B2(n5768), .A(n4895), .ZN(n4897) );
  OAI21_X1 U5984 ( .B1(n4909), .B2(n5557), .A(n4897), .ZN(U2974) );
  INV_X1 U5985 ( .A(n4898), .ZN(n4901) );
  INV_X1 U5986 ( .A(n5356), .ZN(n4899) );
  AOI22_X1 U5987 ( .A1(n4901), .A2(n4900), .B1(n4899), .B2(n5526), .ZN(n5785)
         );
  OAI221_X1 U5988 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n4903), .C1(
        INSTADDRPOINTER_REG_11__SCAN_IN), .C2(n4902), .A(n5785), .ZN(n4905) );
  OAI21_X1 U5989 ( .B1(n6798), .B2(n5786), .A(n6916), .ZN(n4904) );
  OAI21_X1 U5990 ( .B1(n6916), .B2(n4905), .A(n4904), .ZN(n4908) );
  AOI21_X1 U5991 ( .B1(n5594), .B2(n5834), .A(n4906), .ZN(n4907) );
  OAI211_X1 U5992 ( .C1(n4909), .C2(n5824), .A(n4908), .B(n4907), .ZN(U3006)
         );
  XOR2_X1 U5993 ( .A(n4911), .B(n4910), .Z(n4946) );
  XNOR2_X1 U5994 ( .A(n4912), .B(n4928), .ZN(n5539) );
  AOI22_X1 U5995 ( .A1(n5539), .A2(n4502), .B1(EBX_REG_13__SCAN_IN), .B2(n5145), .ZN(n4913) );
  OAI21_X1 U5996 ( .B1(n4949), .B2(n5162), .A(n4913), .ZN(U2846) );
  INV_X1 U5997 ( .A(n4944), .ZN(n4919) );
  OAI21_X1 U5998 ( .B1(REIP_REG_13__SCAN_IN), .B2(REIP_REG_12__SCAN_IN), .A(
        n4914), .ZN(n4915) );
  INV_X1 U5999 ( .A(REIP_REG_13__SCAN_IN), .ZN(n6562) );
  OAI22_X1 U6000 ( .A1(n5602), .A2(n4915), .B1(n6562), .B2(n5601), .ZN(n4918)
         );
  AOI22_X1 U6001 ( .A1(EBX_REG_13__SCAN_IN), .A2(n5693), .B1(n5690), .B2(n5539), .ZN(n4916) );
  OAI211_X1 U6002 ( .C1(n5692), .C2(n6740), .A(n4916), .B(n5640), .ZN(n4917)
         );
  AOI211_X1 U6003 ( .C1(n5677), .C2(n4919), .A(n4918), .B(n4917), .ZN(n4920)
         );
  OAI21_X1 U6004 ( .B1(n4949), .B2(n5620), .A(n4920), .ZN(U2814) );
  OAI21_X1 U6005 ( .B1(n4923), .B2(n4922), .A(n4921), .ZN(n4964) );
  INV_X1 U6006 ( .A(n5688), .ZN(n5090) );
  NOR2_X1 U6007 ( .A1(n5090), .A2(n4924), .ZN(n5583) );
  OAI21_X1 U6008 ( .B1(REIP_REG_14__SCAN_IN), .B2(n4925), .A(n5583), .ZN(n4926) );
  OAI21_X1 U6009 ( .B1(n4960), .B2(n5691), .A(n4926), .ZN(n4933) );
  AOI21_X1 U6010 ( .B1(n4929), .B2(n4928), .A(n4927), .ZN(n4930) );
  OR2_X1 U6011 ( .A1(n4930), .A2(n5159), .ZN(n4935) );
  INV_X1 U6012 ( .A(n4935), .ZN(n5524) );
  AOI22_X1 U6013 ( .A1(PHYADDRPOINTER_REG_14__SCAN_IN), .A2(n5674), .B1(n5690), 
        .B2(n5524), .ZN(n4931) );
  OAI211_X1 U6014 ( .C1(n5665), .C2(n6896), .A(n4931), .B(n5640), .ZN(n4932)
         );
  NOR2_X1 U6015 ( .A1(n4933), .A2(n4932), .ZN(n4934) );
  OAI21_X1 U6016 ( .B1(n4964), .B2(n5620), .A(n4934), .ZN(U2813) );
  OAI22_X1 U6017 ( .A1(n4935), .A2(n5156), .B1(n6896), .B2(n5706), .ZN(n4936)
         );
  INV_X1 U6018 ( .A(n4936), .ZN(n4937) );
  OAI21_X1 U6019 ( .B1(n4964), .B2(n5162), .A(n4937), .ZN(U2845) );
  AOI22_X1 U6020 ( .A1(n4956), .A2(DATAI_14_), .B1(n5710), .B2(
        EAX_REG_14__SCAN_IN), .ZN(n4938) );
  OAI21_X1 U6021 ( .B1(n4964), .B2(n5468), .A(n4938), .ZN(U2877) );
  NAND2_X1 U6022 ( .A1(n4939), .A2(n4940), .ZN(n4941) );
  NAND2_X1 U6023 ( .A1(n4942), .A2(n4941), .ZN(n5543) );
  INV_X1 U6024 ( .A(n5543), .ZN(n4948) );
  AOI22_X1 U6025 ( .A1(n5777), .A2(PHYADDRPOINTER_REG_13__SCAN_IN), .B1(n5262), 
        .B2(REIP_REG_13__SCAN_IN), .ZN(n4943) );
  OAI21_X1 U6026 ( .B1(n5773), .B2(n4944), .A(n4943), .ZN(n4945) );
  AOI21_X1 U6027 ( .B1(n4946), .B2(n5768), .A(n4945), .ZN(n4947) );
  OAI21_X1 U6028 ( .B1(n4948), .B2(n5557), .A(n4947), .ZN(U2973) );
  INV_X1 U6029 ( .A(EAX_REG_13__SCAN_IN), .ZN(n5727) );
  OAI222_X1 U6030 ( .A1(n5164), .A2(n5727), .B1(n4951), .B2(n4950), .C1(n5468), 
        .C2(n4949), .ZN(U2878) );
  INV_X1 U6032 ( .A(n4953), .ZN(n4954) );
  AOI21_X1 U6033 ( .B1(n4955), .B2(n4921), .A(n4954), .ZN(n5588) );
  INV_X1 U6034 ( .A(n5588), .ZN(n5163) );
  AOI22_X1 U6035 ( .A1(n4956), .A2(DATAI_15_), .B1(n5710), .B2(
        EAX_REG_15__SCAN_IN), .ZN(n4957) );
  OAI21_X1 U6036 ( .B1(n5163), .B2(n5468), .A(n4957), .ZN(U2876) );
  XNOR2_X1 U6037 ( .A(n5245), .B(INSTADDRPOINTER_REG_14__SCAN_IN), .ZN(n4959)
         );
  XNOR2_X1 U6038 ( .A(n4958), .B(n4959), .ZN(n5532) );
  NAND2_X1 U6039 ( .A1(n5532), .A2(n5774), .ZN(n4963) );
  NOR2_X1 U6040 ( .A1(n5811), .A2(n6563), .ZN(n5523) );
  NOR2_X1 U6041 ( .A1(n5773), .A2(n4960), .ZN(n4961) );
  AOI211_X1 U6042 ( .C1(n5777), .C2(PHYADDRPOINTER_REG_14__SCAN_IN), .A(n5523), 
        .B(n4961), .ZN(n4962) );
  OAI211_X1 U6043 ( .C1(n5911), .C2(n4964), .A(n4963), .B(n4962), .ZN(U2972)
         );
  AOI21_X1 U6044 ( .B1(n4966), .B2(n4953), .A(n4965), .ZN(n5266) );
  NAND2_X1 U6045 ( .A1(n5161), .A2(n4967), .ZN(n4968) );
  NAND2_X1 U6046 ( .A1(n4987), .A2(n4968), .ZN(n5512) );
  INV_X1 U6047 ( .A(EBX_REG_16__SCAN_IN), .ZN(n4973) );
  OAI22_X1 U6048 ( .A1(n5512), .A2(n5156), .B1(n4973), .B2(n5706), .ZN(n4969)
         );
  AOI21_X1 U6049 ( .B1(n5266), .B2(n5703), .A(n4969), .ZN(n4970) );
  INV_X1 U6050 ( .A(n4970), .ZN(U2843) );
  INV_X1 U6051 ( .A(n5266), .ZN(n4982) );
  INV_X1 U6052 ( .A(REIP_REG_16__SCAN_IN), .ZN(n6869) );
  INV_X1 U6053 ( .A(REIP_REG_15__SCAN_IN), .ZN(n6565) );
  AOI21_X1 U6054 ( .B1(n6869), .B2(n6565), .A(n5591), .ZN(n4976) );
  AOI21_X1 U6055 ( .B1(n5674), .B2(PHYADDRPOINTER_REG_16__SCAN_IN), .A(n5651), 
        .ZN(n4971) );
  OAI21_X1 U6056 ( .B1(n5512), .B2(n5681), .A(n4971), .ZN(n4975) );
  AOI22_X1 U6057 ( .A1(n5261), .A2(n5677), .B1(REIP_REG_16__SCAN_IN), .B2(
        n5583), .ZN(n4972) );
  OAI21_X1 U6058 ( .B1(n4973), .B2(n5665), .A(n4972), .ZN(n4974) );
  AOI211_X1 U6059 ( .C1(n4977), .C2(n4976), .A(n4975), .B(n4974), .ZN(n4978)
         );
  OAI21_X1 U6060 ( .B1(n4982), .B2(n5620), .A(n4978), .ZN(U2811) );
  AOI22_X1 U6061 ( .A1(n5707), .A2(DATAI_16_), .B1(n5710), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n4981) );
  NOR3_X4 U6062 ( .A1(n5710), .A2(n5165), .A3(n3402), .ZN(n5711) );
  NAND2_X1 U6063 ( .A1(n5711), .A2(DATAI_0_), .ZN(n4980) );
  OAI211_X1 U6064 ( .C1(n4982), .C2(n5468), .A(n4981), .B(n4980), .ZN(U2875)
         );
  OR2_X1 U6065 ( .A1(n4965), .A2(n4984), .ZN(n4985) );
  AND2_X1 U6066 ( .A1(n4983), .A2(n4985), .ZN(n5709) );
  INV_X1 U6067 ( .A(n5709), .ZN(n4990) );
  INV_X1 U6068 ( .A(EBX_REG_17__SCAN_IN), .ZN(n4989) );
  AND2_X1 U6069 ( .A1(n4987), .A2(n4986), .ZN(n4988) );
  OR2_X1 U6070 ( .A1(n4988), .A2(n5078), .ZN(n5582) );
  OAI222_X1 U6071 ( .A1(n4990), .A2(n5162), .B1(n4989), .B2(n5706), .C1(n5156), 
        .C2(n5582), .ZN(U2842) );
  INV_X1 U6072 ( .A(n5006), .ZN(n5000) );
  AOI22_X1 U6073 ( .A1(n5707), .A2(DATAI_30_), .B1(n5710), .B2(
        EAX_REG_30__SCAN_IN), .ZN(n4992) );
  NAND2_X1 U6074 ( .A1(n5711), .A2(DATAI_14_), .ZN(n4991) );
  OAI211_X1 U6075 ( .C1(n5000), .C2(n5468), .A(n4992), .B(n4991), .ZN(U2861)
         );
  NAND3_X1 U6076 ( .A1(n5030), .A2(REIP_REG_30__SCAN_IN), .A3(n5688), .ZN(
        n4994) );
  AOI22_X1 U6077 ( .A1(PHYADDRPOINTER_REG_30__SCAN_IN), .A2(n5674), .B1(n5677), 
        .B2(n5001), .ZN(n4993) );
  OAI211_X1 U6078 ( .C1(n4995), .C2(n5665), .A(n4994), .B(n4993), .ZN(n4997)
         );
  NOR3_X1 U6079 ( .A1(n5029), .A2(REIP_REG_30__SCAN_IN), .A3(n6585), .ZN(n4996) );
  AOI211_X1 U6080 ( .C1(n5690), .C2(n4998), .A(n4997), .B(n4996), .ZN(n4999)
         );
  OAI21_X1 U6081 ( .B1(n5000), .B2(n5620), .A(n4999), .ZN(U2797) );
  INV_X1 U6082 ( .A(n5001), .ZN(n5004) );
  AOI21_X1 U6083 ( .B1(n5777), .B2(PHYADDRPOINTER_REG_30__SCAN_IN), .A(n5002), 
        .ZN(n5003) );
  OAI21_X1 U6084 ( .B1(n5773), .B2(n5004), .A(n5003), .ZN(n5005) );
  AOI21_X1 U6085 ( .B1(n5006), .B2(n5768), .A(n5005), .ZN(n5007) );
  OAI21_X1 U6086 ( .B1(n5008), .B2(n5557), .A(n5007), .ZN(U2956) );
  INV_X1 U6087 ( .A(n4550), .ZN(n5011) );
  AOI21_X1 U6088 ( .B1(n5009), .B2(n5011), .A(n5015), .ZN(n5017) );
  NOR3_X1 U6089 ( .A1(n6522), .A2(n6605), .A3(n5010), .ZN(n5013) );
  NOR3_X1 U6090 ( .A1(n6601), .A2(INSTQUEUERD_ADDR_REG_2__SCAN_IN), .A3(n5011), 
        .ZN(n5012) );
  AOI211_X1 U6091 ( .C1(n5014), .C2(n6606), .A(n5013), .B(n5012), .ZN(n5016)
         );
  OAI22_X1 U6092 ( .A1(n5017), .A2(n3258), .B1(n5016), .B2(n5015), .ZN(U3459)
         );
  AOI21_X1 U6093 ( .B1(n5020), .B2(n5018), .A(n5019), .ZN(n5188) );
  INV_X1 U6094 ( .A(n5188), .ZN(n5171) );
  OAI22_X1 U6095 ( .A1(n5021), .A2(n5692), .B1(n5691), .B2(n5186), .ZN(n5028)
         );
  INV_X1 U6096 ( .A(n5022), .ZN(n5026) );
  INV_X1 U6097 ( .A(n5023), .ZN(n5025) );
  OAI21_X1 U6098 ( .B1(n5026), .B2(n5025), .A(n5024), .ZN(n5289) );
  NOR2_X1 U6099 ( .A1(n5289), .A2(n5681), .ZN(n5027) );
  AOI211_X1 U6100 ( .C1(n5693), .C2(EBX_REG_29__SCAN_IN), .A(n5028), .B(n5027), 
        .ZN(n5033) );
  INV_X1 U6101 ( .A(n5029), .ZN(n5031) );
  OAI21_X1 U6102 ( .B1(n5031), .B2(REIP_REG_29__SCAN_IN), .A(n5030), .ZN(n5032) );
  OAI211_X1 U6103 ( .C1(n5171), .C2(n5620), .A(n5033), .B(n5032), .ZN(U2798)
         );
  OAI21_X1 U6104 ( .B1(n5034), .B2(n5035), .A(n5018), .ZN(n5190) );
  NAND3_X1 U6105 ( .A1(REIP_REG_27__SCAN_IN), .A2(n5409), .A3(n6582), .ZN(
        n5044) );
  NAND2_X1 U6106 ( .A1(n5414), .A2(n5036), .ZN(n5042) );
  INV_X1 U6107 ( .A(n5037), .ZN(n5193) );
  OAI22_X1 U6108 ( .A1(n5038), .A2(n5692), .B1(n5691), .B2(n5193), .ZN(n5039)
         );
  AOI21_X1 U6109 ( .B1(n5693), .B2(EBX_REG_28__SCAN_IN), .A(n5039), .ZN(n5040)
         );
  OAI21_X1 U6110 ( .B1(n5107), .B2(n5681), .A(n5040), .ZN(n5041) );
  AOI21_X1 U6111 ( .B1(REIP_REG_28__SCAN_IN), .B2(n5042), .A(n5041), .ZN(n5043) );
  OAI211_X1 U6112 ( .C1(n5190), .C2(n5620), .A(n5044), .B(n5043), .ZN(U2799)
         );
  NOR2_X1 U6113 ( .A1(n5090), .A2(n5045), .ZN(n5451) );
  INV_X1 U6114 ( .A(REIP_REG_21__SCAN_IN), .ZN(n5046) );
  NAND2_X1 U6115 ( .A1(n5046), .A2(n5048), .ZN(n5453) );
  INV_X1 U6116 ( .A(n5453), .ZN(n5047) );
  OAI21_X1 U6117 ( .B1(n5451), .B2(n5047), .A(REIP_REG_22__SCAN_IN), .ZN(n5058) );
  NAND2_X1 U6118 ( .A1(REIP_REG_21__SCAN_IN), .A2(n5048), .ZN(n5444) );
  OAI22_X1 U6119 ( .A1(REIP_REG_22__SCAN_IN), .A2(n5444), .B1(n5049), .B2(
        n5665), .ZN(n5056) );
  INV_X1 U6120 ( .A(n5344), .ZN(n5050) );
  NOR2_X1 U6121 ( .A1(n5345), .A2(n5050), .ZN(n5052) );
  OAI21_X1 U6122 ( .B1(n5052), .B2(n5051), .A(n3137), .ZN(n5343) );
  AOI22_X1 U6123 ( .A1(PHYADDRPOINTER_REG_22__SCAN_IN), .A2(n5674), .B1(n5053), 
        .B2(n5677), .ZN(n5054) );
  OAI21_X1 U6124 ( .B1(n5343), .B2(n5681), .A(n5054), .ZN(n5055) );
  NOR2_X1 U6125 ( .A1(n5056), .A2(n5055), .ZN(n5057) );
  OAI211_X1 U6126 ( .C1(n5178), .C2(n5620), .A(n5058), .B(n5057), .ZN(U2805)
         );
  NOR2_X1 U6127 ( .A1(n5060), .A2(n5061), .ZN(n5062) );
  OR2_X1 U6128 ( .A1(n5059), .A2(n5062), .ZN(n5484) );
  NAND2_X1 U6129 ( .A1(REIP_REG_19__SCAN_IN), .A2(REIP_REG_18__SCAN_IN), .ZN(
        n5461) );
  INV_X1 U6130 ( .A(REIP_REG_20__SCAN_IN), .ZN(n6572) );
  OAI21_X1 U6131 ( .B1(n5073), .B2(n5461), .A(n6572), .ZN(n5069) );
  MUX2_X1 U6132 ( .A(n4159), .B(n5075), .S(n5063), .Z(n5065) );
  XNOR2_X1 U6133 ( .A(n5065), .B(n5064), .ZN(n5366) );
  INV_X1 U6134 ( .A(n5366), .ZN(n5148) );
  INV_X1 U6135 ( .A(EBX_REG_20__SCAN_IN), .ZN(n6935) );
  OAI22_X1 U6136 ( .A1(n6935), .A2(n5665), .B1(n6690), .B2(n5692), .ZN(n5066)
         );
  AOI21_X1 U6137 ( .B1(n5677), .B2(n5242), .A(n5066), .ZN(n5067) );
  OAI21_X1 U6138 ( .B1(n5148), .B2(n5681), .A(n5067), .ZN(n5068) );
  AOI21_X1 U6139 ( .B1(n5069), .B2(n5451), .A(n5068), .ZN(n5070) );
  OAI21_X1 U6140 ( .B1(n5484), .B2(n5620), .A(n5070), .ZN(U2807) );
  INV_X1 U6141 ( .A(n4983), .ZN(n5072) );
  OAI21_X1 U6142 ( .B1(n5072), .B2(n3253), .A(n5071), .ZN(n5254) );
  INV_X1 U6143 ( .A(n5073), .ZN(n5462) );
  INV_X1 U6144 ( .A(REIP_REG_18__SCAN_IN), .ZN(n6569) );
  MUX2_X1 U6145 ( .A(n5075), .B(n5074), .S(n4122), .Z(n5076) );
  INV_X1 U6146 ( .A(n5076), .ZN(n5077) );
  NAND2_X1 U6147 ( .A1(n5078), .A2(n5077), .ZN(n5152) );
  OR2_X1 U6148 ( .A1(n5078), .A2(n5077), .ZN(n5079) );
  AND2_X1 U6149 ( .A1(n5152), .A2(n5079), .ZN(n5506) );
  INV_X1 U6150 ( .A(n5506), .ZN(n5155) );
  AOI21_X1 U6151 ( .B1(n5674), .B2(PHYADDRPOINTER_REG_18__SCAN_IN), .A(n5651), 
        .ZN(n5080) );
  OAI21_X1 U6152 ( .B1(n5155), .B2(n5681), .A(n5080), .ZN(n5084) );
  NAND2_X1 U6153 ( .A1(n5688), .A2(n5081), .ZN(n5577) );
  AOI22_X1 U6154 ( .A1(EBX_REG_18__SCAN_IN), .A2(n5693), .B1(n5251), .B2(n5677), .ZN(n5082) );
  OAI21_X1 U6155 ( .B1(n6569), .B2(n5577), .A(n5082), .ZN(n5083) );
  AOI211_X1 U6156 ( .C1(n5462), .C2(n6569), .A(n5084), .B(n5083), .ZN(n5085)
         );
  OAI21_X1 U6157 ( .B1(n5254), .B2(n5620), .A(n5085), .ZN(U2809) );
  INV_X1 U6158 ( .A(n5086), .ZN(n5788) );
  INV_X1 U6159 ( .A(n5608), .ZN(n5088) );
  OAI22_X1 U6160 ( .A1(n5088), .A2(REIP_REG_9__SCAN_IN), .B1(n5087), .B2(n5691), .ZN(n5094) );
  INV_X1 U6161 ( .A(PHYADDRPOINTER_REG_9__SCAN_IN), .ZN(n5092) );
  NOR2_X1 U6162 ( .A1(n5090), .A2(n5089), .ZN(n5605) );
  AOI22_X1 U6163 ( .A1(EBX_REG_9__SCAN_IN), .A2(n5693), .B1(
        REIP_REG_9__SCAN_IN), .B2(n5605), .ZN(n5091) );
  OAI211_X1 U6164 ( .C1(n5692), .C2(n5092), .A(n5091), .B(n5640), .ZN(n5093)
         );
  AOI211_X1 U6165 ( .C1(n5690), .C2(n5788), .A(n5094), .B(n5093), .ZN(n5095)
         );
  OAI21_X1 U6166 ( .B1(n5620), .B2(n5096), .A(n5095), .ZN(U2818) );
  INV_X1 U6167 ( .A(REIP_REG_7__SCAN_IN), .ZN(n6558) );
  NAND2_X1 U6168 ( .A1(n5098), .A2(n5097), .ZN(n5614) );
  INV_X1 U6169 ( .A(REIP_REG_8__SCAN_IN), .ZN(n6767) );
  OAI21_X1 U6170 ( .B1(n6558), .B2(n5614), .A(n6767), .ZN(n5103) );
  NAND2_X1 U6171 ( .A1(n5693), .A2(EBX_REG_8__SCAN_IN), .ZN(n5099) );
  OAI211_X1 U6172 ( .C1(n5691), .C2(n5100), .A(n5099), .B(n5640), .ZN(n5102)
         );
  OAI22_X1 U6173 ( .A1(n6716), .A2(n5692), .B1(n5681), .B2(n5795), .ZN(n5101)
         );
  AOI211_X1 U6174 ( .C1(n5605), .C2(n5103), .A(n5102), .B(n5101), .ZN(n5104)
         );
  OAI21_X1 U6175 ( .B1(n5105), .B2(n5620), .A(n5104), .ZN(U2819) );
  OAI22_X1 U6176 ( .A1(n5279), .A2(n5156), .B1(n5706), .B2(n6734), .ZN(U2828)
         );
  OAI222_X1 U6177 ( .A1(n5162), .A2(n5171), .B1(n5106), .B2(n5706), .C1(n5289), 
        .C2(n5156), .ZN(U2830) );
  OAI222_X1 U6178 ( .A1(n5162), .A2(n5190), .B1(n6885), .B2(n5706), .C1(n5107), 
        .C2(n5156), .ZN(U2831) );
  INV_X1 U6179 ( .A(n5108), .ZN(n5116) );
  AND2_X1 U6180 ( .A1(n5116), .A2(n5109), .ZN(n5110) );
  OR2_X1 U6181 ( .A1(n5034), .A2(n5110), .ZN(n5200) );
  INV_X1 U6182 ( .A(EBX_REG_27__SCAN_IN), .ZN(n6814) );
  AND2_X1 U6183 ( .A1(n5118), .A2(n5111), .ZN(n5112) );
  OR2_X1 U6184 ( .A1(n5113), .A2(n5112), .ZN(n5412) );
  OAI222_X1 U6185 ( .A1(n5162), .A2(n5200), .B1(n5706), .B2(n6814), .C1(n5412), 
        .C2(n5156), .ZN(U2832) );
  INV_X1 U6186 ( .A(n5114), .ZN(n5124) );
  INV_X1 U6187 ( .A(n5115), .ZN(n5117) );
  INV_X1 U6188 ( .A(EBX_REG_26__SCAN_IN), .ZN(n6868) );
  INV_X1 U6189 ( .A(n5118), .ZN(n5119) );
  AOI21_X1 U6190 ( .B1(n5120), .B2(n3128), .A(n5119), .ZN(n5418) );
  INV_X1 U6191 ( .A(n5418), .ZN(n5121) );
  OAI222_X1 U6192 ( .A1(n5162), .A2(n5416), .B1(n5706), .B2(n6868), .C1(n5121), 
        .C2(n5156), .ZN(U2833) );
  INV_X1 U6193 ( .A(n5122), .ZN(n5126) );
  INV_X1 U6194 ( .A(n5123), .ZN(n5125) );
  OR2_X1 U6195 ( .A1(n5137), .A2(n5127), .ZN(n5128) );
  NAND2_X1 U6196 ( .A1(n3128), .A2(n5128), .ZN(n5431) );
  OAI22_X1 U6197 ( .A1(n5431), .A2(n5156), .B1(n5129), .B2(n5706), .ZN(n5130)
         );
  AOI21_X1 U6198 ( .B1(n5491), .B2(n5703), .A(n5130), .ZN(n5131) );
  INV_X1 U6199 ( .A(n5131), .ZN(U2834) );
  NOR2_X1 U6200 ( .A1(n5132), .A2(n5133), .ZN(n5134) );
  OR2_X1 U6201 ( .A1(n5123), .A2(n5134), .ZN(n5474) );
  NOR2_X1 U6202 ( .A1(n5141), .A2(n5135), .ZN(n5136) );
  OR2_X1 U6203 ( .A1(n5137), .A2(n5136), .ZN(n5433) );
  OAI222_X1 U6204 ( .A1(n5162), .A2(n5474), .B1(n5138), .B2(n5706), .C1(n5433), 
        .C2(n5156), .ZN(U2835) );
  AOI21_X1 U6205 ( .B1(n5139), .B2(n4299), .A(n5132), .ZN(n5478) );
  INV_X1 U6206 ( .A(n5478), .ZN(n5144) );
  INV_X1 U6207 ( .A(EBX_REG_23__SCAN_IN), .ZN(n5143) );
  AND2_X1 U6208 ( .A1(n3137), .A2(n5140), .ZN(n5142) );
  OR2_X1 U6209 ( .A1(n5142), .A2(n5141), .ZN(n5449) );
  OAI222_X1 U6210 ( .A1(n5162), .A2(n5144), .B1(n5143), .B2(n5706), .C1(n5449), 
        .C2(n5156), .ZN(U2836) );
  INV_X1 U6211 ( .A(n5343), .ZN(n5146) );
  AOI22_X1 U6212 ( .A1(n5146), .A2(n4502), .B1(EBX_REG_22__SCAN_IN), .B2(n5145), .ZN(n5147) );
  OAI21_X1 U6213 ( .B1(n5178), .B2(n5162), .A(n5147), .ZN(U2837) );
  OAI222_X1 U6214 ( .A1(n5484), .A2(n5162), .B1(n5706), .B2(n6935), .C1(n5148), 
        .C2(n5156), .ZN(U2839) );
  AND2_X1 U6215 ( .A1(n5071), .A2(n5149), .ZN(n5150) );
  NOR2_X1 U6216 ( .A1(n5060), .A2(n5150), .ZN(n5495) );
  INV_X1 U6217 ( .A(n5495), .ZN(n5154) );
  INV_X1 U6218 ( .A(EBX_REG_19__SCAN_IN), .ZN(n5153) );
  XNOR2_X1 U6219 ( .A(n5152), .B(n5151), .ZN(n5465) );
  OAI222_X1 U6220 ( .A1(n5154), .A2(n5162), .B1(n5153), .B2(n5706), .C1(n5156), 
        .C2(n5465), .ZN(U2840) );
  OAI222_X1 U6221 ( .A1(n5254), .A2(n5162), .B1(n5157), .B2(n5706), .C1(n5156), 
        .C2(n5155), .ZN(U2841) );
  OR2_X1 U6222 ( .A1(n5159), .A2(n5158), .ZN(n5160) );
  NAND2_X1 U6223 ( .A1(n5161), .A2(n5160), .ZN(n5585) );
  INV_X1 U6224 ( .A(EBX_REG_15__SCAN_IN), .ZN(n6845) );
  OAI222_X1 U6225 ( .A1(n5585), .A2(n5156), .B1(n5706), .B2(n6845), .C1(n5163), 
        .C2(n5162), .ZN(U2844) );
  NAND3_X1 U6226 ( .A1(n5166), .A2(n5165), .A3(n5164), .ZN(n5168) );
  AOI22_X1 U6227 ( .A1(n5707), .A2(DATAI_31_), .B1(EAX_REG_31__SCAN_IN), .B2(
        n5710), .ZN(n5167) );
  NAND2_X1 U6228 ( .A1(n5168), .A2(n5167), .ZN(U2860) );
  AOI22_X1 U6229 ( .A1(n5707), .A2(DATAI_29_), .B1(n5710), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5170) );
  NAND2_X1 U6230 ( .A1(n5711), .A2(DATAI_13_), .ZN(n5169) );
  OAI211_X1 U6231 ( .C1(n5171), .C2(n5468), .A(n5170), .B(n5169), .ZN(U2862)
         );
  AOI22_X1 U6232 ( .A1(n5707), .A2(DATAI_28_), .B1(n5710), .B2(
        EAX_REG_28__SCAN_IN), .ZN(n5173) );
  NAND2_X1 U6233 ( .A1(n5711), .A2(DATAI_12_), .ZN(n5172) );
  OAI211_X1 U6234 ( .C1(n5190), .C2(n5468), .A(n5173), .B(n5172), .ZN(U2863)
         );
  AOI22_X1 U6235 ( .A1(n5711), .A2(DATAI_10_), .B1(EAX_REG_26__SCAN_IN), .B2(
        n5710), .ZN(n5175) );
  NAND2_X1 U6236 ( .A1(n5707), .A2(DATAI_26_), .ZN(n5174) );
  OAI211_X1 U6237 ( .C1(n5416), .C2(n5468), .A(n5175), .B(n5174), .ZN(U2865)
         );
  AOI22_X1 U6238 ( .A1(n5707), .A2(DATAI_22_), .B1(n5710), .B2(
        EAX_REG_22__SCAN_IN), .ZN(n5177) );
  NAND2_X1 U6239 ( .A1(n5711), .A2(DATAI_6_), .ZN(n5176) );
  OAI211_X1 U6240 ( .C1(n5178), .C2(n5468), .A(n5177), .B(n5176), .ZN(U2869)
         );
  AOI22_X1 U6241 ( .A1(n5707), .A2(DATAI_18_), .B1(n5710), .B2(
        EAX_REG_18__SCAN_IN), .ZN(n5180) );
  NAND2_X1 U6242 ( .A1(n5711), .A2(DATAI_2_), .ZN(n5179) );
  OAI211_X1 U6243 ( .C1(n5254), .C2(n5468), .A(n5180), .B(n5179), .ZN(U2873)
         );
  AOI21_X1 U6244 ( .B1(n5284), .B2(n5182), .A(n5181), .ZN(n5184) );
  XNOR2_X1 U6245 ( .A(n5184), .B(n5183), .ZN(n5293) );
  AND2_X1 U6246 ( .A1(n5262), .A2(REIP_REG_29__SCAN_IN), .ZN(n5287) );
  AOI21_X1 U6247 ( .B1(n5777), .B2(PHYADDRPOINTER_REG_29__SCAN_IN), .A(n5287), 
        .ZN(n5185) );
  OAI21_X1 U6248 ( .B1(n5773), .B2(n5186), .A(n5185), .ZN(n5187) );
  AOI21_X1 U6249 ( .B1(n5188), .B2(n5768), .A(n5187), .ZN(n5189) );
  OAI21_X1 U6250 ( .B1(n5293), .B2(n5557), .A(n5189), .ZN(U2957) );
  INV_X1 U6251 ( .A(n5190), .ZN(n5195) );
  AOI21_X1 U6252 ( .B1(n5777), .B2(PHYADDRPOINTER_REG_28__SCAN_IN), .A(n5191), 
        .ZN(n5192) );
  OAI21_X1 U6253 ( .B1(n5773), .B2(n5193), .A(n5192), .ZN(n5194) );
  OAI21_X1 U6254 ( .B1(n5197), .B2(n5557), .A(n5196), .ZN(U2958) );
  OAI21_X1 U6255 ( .B1(n5312), .B2(n5204), .A(n5198), .ZN(n5199) );
  XNOR2_X1 U6256 ( .A(n5199), .B(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5301)
         );
  AND2_X1 U6257 ( .A1(n5262), .A2(REIP_REG_27__SCAN_IN), .ZN(n5296) );
  AOI21_X1 U6258 ( .B1(n5777), .B2(PHYADDRPOINTER_REG_27__SCAN_IN), .A(n5296), 
        .ZN(n5201) );
  OAI21_X1 U6259 ( .B1(n5773), .B2(n5405), .A(n5201), .ZN(n5202) );
  AOI21_X1 U6260 ( .B1(n5469), .B2(n5768), .A(n5202), .ZN(n5203) );
  OAI21_X1 U6261 ( .B1(n5301), .B2(n5557), .A(n5203), .ZN(U2959) );
  INV_X1 U6262 ( .A(n5204), .ZN(n5206) );
  NOR2_X1 U6263 ( .A1(n5206), .A2(n5205), .ZN(n5208) );
  XOR2_X1 U6264 ( .A(n5208), .B(n5207), .Z(n5310) );
  INV_X1 U6265 ( .A(n5416), .ZN(n5212) );
  INV_X1 U6266 ( .A(n5413), .ZN(n5210) );
  AND2_X1 U6267 ( .A1(n5262), .A2(REIP_REG_26__SCAN_IN), .ZN(n5303) );
  AOI21_X1 U6268 ( .B1(n5777), .B2(PHYADDRPOINTER_REG_26__SCAN_IN), .A(n5303), 
        .ZN(n5209) );
  OAI21_X1 U6269 ( .B1(n5773), .B2(n5210), .A(n5209), .ZN(n5211) );
  AOI21_X1 U6270 ( .B1(n5212), .B2(n5768), .A(n5211), .ZN(n5213) );
  OAI21_X1 U6271 ( .B1(n5310), .B2(n5557), .A(n5213), .ZN(U2960) );
  NAND3_X1 U6272 ( .A1(n5222), .A2(INSTADDRPOINTER_REG_23__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_22__SCAN_IN), .ZN(n5215) );
  XNOR2_X1 U6273 ( .A(n5217), .B(INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5325)
         );
  INV_X1 U6274 ( .A(PHYADDRPOINTER_REG_24__SCAN_IN), .ZN(n6887) );
  NAND2_X1 U6275 ( .A1(n5262), .A2(REIP_REG_24__SCAN_IN), .ZN(n5319) );
  OAI21_X1 U6276 ( .B1(n5248), .B2(n6887), .A(n5319), .ZN(n5219) );
  NOR2_X1 U6277 ( .A1(n5474), .A2(n5911), .ZN(n5218) );
  AOI211_X1 U6278 ( .C1(n5250), .C2(n5432), .A(n5219), .B(n5218), .ZN(n5220)
         );
  OAI21_X1 U6279 ( .B1(n5325), .B2(n5557), .A(n5220), .ZN(U2962) );
  NAND3_X1 U6280 ( .A1(n5222), .A2(INSTADDRPOINTER_REG_20__SCAN_IN), .A3(n5335), .ZN(n5224) );
  OAI21_X1 U6281 ( .B1(n5221), .B2(n5224), .A(n5223), .ZN(n5225) );
  XNOR2_X1 U6282 ( .A(n5225), .B(INSTADDRPOINTER_REG_23__SCAN_IN), .ZN(n5333)
         );
  NAND2_X1 U6283 ( .A1(n5832), .A2(REIP_REG_23__SCAN_IN), .ZN(n5327) );
  NAND2_X1 U6284 ( .A1(n5777), .A2(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5226)
         );
  OAI211_X1 U6285 ( .C1(n5773), .C2(n5440), .A(n5327), .B(n5226), .ZN(n5227)
         );
  AOI21_X1 U6286 ( .B1(n5478), .B2(n5768), .A(n5227), .ZN(n5228) );
  OAI21_X1 U6287 ( .B1(n5333), .B2(n5557), .A(n5228), .ZN(U2963) );
  AOI21_X1 U6288 ( .B1(n5231), .B2(n5230), .A(n5229), .ZN(n5353) );
  INV_X1 U6289 ( .A(n5232), .ZN(n5235) );
  INV_X1 U6290 ( .A(n5059), .ZN(n5234) );
  AOI21_X1 U6291 ( .B1(n5235), .B2(n5234), .A(n5233), .ZN(n5481) );
  NAND2_X1 U6292 ( .A1(n5832), .A2(REIP_REG_21__SCAN_IN), .ZN(n5348) );
  NAND2_X1 U6293 ( .A1(n5777), .A2(PHYADDRPOINTER_REG_21__SCAN_IN), .ZN(n5236)
         );
  OAI211_X1 U6294 ( .C1(n5773), .C2(n5450), .A(n5348), .B(n5236), .ZN(n5237)
         );
  AOI21_X1 U6295 ( .B1(n5481), .B2(n5768), .A(n5237), .ZN(n5238) );
  OAI21_X1 U6296 ( .B1(n5353), .B2(n5557), .A(n5238), .ZN(U2965) );
  XNOR2_X1 U6297 ( .A(n5221), .B(n5239), .ZN(n5368) );
  NAND2_X1 U6298 ( .A1(n5262), .A2(REIP_REG_20__SCAN_IN), .ZN(n5363) );
  OAI21_X1 U6299 ( .B1(n5248), .B2(n6690), .A(n5363), .ZN(n5241) );
  NOR2_X1 U6300 ( .A1(n5484), .A2(n5911), .ZN(n5240) );
  AOI211_X1 U6301 ( .C1(n5250), .C2(n5242), .A(n5241), .B(n5240), .ZN(n5243)
         );
  OAI21_X1 U6302 ( .B1(n5557), .B2(n5368), .A(n5243), .ZN(U2966) );
  INV_X1 U6303 ( .A(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5504) );
  NOR3_X1 U6304 ( .A1(n5244), .A2(n3680), .A3(n5504), .ZN(n5383) );
  OR2_X1 U6305 ( .A1(n5245), .A2(INSTADDRPOINTER_REG_16__SCAN_IN), .ZN(n5380)
         );
  NOR3_X1 U6306 ( .A1(n5246), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .A3(n5380), 
        .ZN(n5381) );
  NOR2_X1 U6307 ( .A1(n5383), .A2(n5381), .ZN(n5247) );
  XNOR2_X1 U6308 ( .A(n5247), .B(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5507)
         );
  NAND2_X1 U6309 ( .A1(n5507), .A2(n5774), .ZN(n5253) );
  OAI22_X1 U6310 ( .A1(n5248), .A2(n6705), .B1(n5811), .B2(n6569), .ZN(n5249)
         );
  AOI21_X1 U6311 ( .B1(n5251), .B2(n5250), .A(n5249), .ZN(n5252) );
  OAI211_X1 U6312 ( .C1(n5911), .C2(n5254), .A(n5253), .B(n5252), .ZN(U2968)
         );
  INV_X1 U6313 ( .A(n5255), .ZN(n5257) );
  OR2_X1 U6314 ( .A1(n5244), .A2(n5257), .ZN(n5260) );
  OAI21_X1 U6315 ( .B1(n5258), .B2(n5257), .A(n5256), .ZN(n5259) );
  NAND2_X1 U6316 ( .A1(n5260), .A2(n5259), .ZN(n5513) );
  INV_X1 U6317 ( .A(n5261), .ZN(n5264) );
  AOI22_X1 U6318 ( .A1(n5777), .A2(PHYADDRPOINTER_REG_16__SCAN_IN), .B1(n5262), 
        .B2(REIP_REG_16__SCAN_IN), .ZN(n5263) );
  OAI21_X1 U6319 ( .B1(n5773), .B2(n5264), .A(n5263), .ZN(n5265) );
  AOI21_X1 U6320 ( .B1(n5266), .B2(n5768), .A(n5265), .ZN(n5267) );
  OAI21_X1 U6321 ( .B1(n5513), .B2(n5557), .A(n5267), .ZN(U2970) );
  XNOR2_X1 U6322 ( .A(n3685), .B(n6844), .ZN(n5269) );
  XNOR2_X1 U6323 ( .A(n5268), .B(n5269), .ZN(n5394) );
  AOI22_X1 U6324 ( .A1(n5777), .A2(PHYADDRPOINTER_REG_15__SCAN_IN), .B1(n5832), 
        .B2(REIP_REG_15__SCAN_IN), .ZN(n5270) );
  OAI21_X1 U6325 ( .B1(n5773), .B2(n5271), .A(n5270), .ZN(n5272) );
  AOI21_X1 U6326 ( .B1(n5588), .B2(n5768), .A(n5272), .ZN(n5273) );
  OAI21_X1 U6327 ( .B1(n5557), .B2(n5394), .A(n5273), .ZN(U2971) );
  OAI21_X1 U6328 ( .B1(INSTADDRPOINTER_REG_30__SCAN_IN), .B2(n5852), .A(n5274), 
        .ZN(n5278) );
  NOR4_X1 U6329 ( .A1(n5294), .A2(INSTADDRPOINTER_REG_31__SCAN_IN), .A3(n5275), 
        .A4(n4253), .ZN(n5276) );
  AOI211_X1 U6330 ( .C1(n5278), .C2(INSTADDRPOINTER_REG_31__SCAN_IN), .A(n5277), .B(n5276), .ZN(n5282) );
  INV_X1 U6331 ( .A(n5279), .ZN(n5280) );
  NAND2_X1 U6332 ( .A1(n5280), .A2(n5834), .ZN(n5281) );
  OAI211_X1 U6333 ( .C1(n5283), .C2(n5824), .A(n5282), .B(n5281), .ZN(U2987)
         );
  INV_X1 U6334 ( .A(n5284), .ZN(n5285) );
  NOR3_X1 U6335 ( .A1(n5294), .A2(INSTADDRPOINTER_REG_29__SCAN_IN), .A3(n5285), 
        .ZN(n5286) );
  AOI211_X1 U6336 ( .C1(n5288), .C2(INSTADDRPOINTER_REG_29__SCAN_IN), .A(n5287), .B(n5286), .ZN(n5292) );
  INV_X1 U6337 ( .A(n5289), .ZN(n5290) );
  NAND2_X1 U6338 ( .A1(n5290), .A2(n5834), .ZN(n5291) );
  OAI211_X1 U6339 ( .C1(n5293), .C2(n5824), .A(n5292), .B(n5291), .ZN(U2989)
         );
  NOR2_X1 U6340 ( .A1(n5294), .A2(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n5295)
         );
  AOI211_X1 U6341 ( .C1(n5297), .C2(INSTADDRPOINTER_REG_27__SCAN_IN), .A(n5296), .B(n5295), .ZN(n5300) );
  INV_X1 U6342 ( .A(n5412), .ZN(n5298) );
  NAND2_X1 U6343 ( .A1(n5298), .A2(n5834), .ZN(n5299) );
  OAI211_X1 U6344 ( .C1(n5301), .C2(n5824), .A(n5300), .B(n5299), .ZN(U2991)
         );
  NAND2_X1 U6345 ( .A1(n5302), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5306) );
  NOR2_X1 U6346 ( .A1(n5307), .A2(INSTADDRPOINTER_REG_25__SCAN_IN), .ZN(n5315)
         );
  OAI21_X1 U6347 ( .B1(n5318), .B2(n5315), .A(INSTADDRPOINTER_REG_26__SCAN_IN), 
        .ZN(n5305) );
  INV_X1 U6348 ( .A(n5303), .ZN(n5304) );
  OAI211_X1 U6349 ( .C1(n5307), .C2(n5306), .A(n5305), .B(n5304), .ZN(n5308)
         );
  AOI21_X1 U6350 ( .B1(n5418), .B2(n5834), .A(n5308), .ZN(n5309) );
  OAI21_X1 U6351 ( .B1(n5310), .B2(n5824), .A(n5309), .ZN(U2992) );
  OAI21_X1 U6352 ( .B1(n5313), .B2(n5311), .A(n5312), .ZN(n5490) );
  NAND2_X1 U6353 ( .A1(n5490), .A2(n5854), .ZN(n5317) );
  AND2_X1 U6354 ( .A1(n5832), .A2(REIP_REG_25__SCAN_IN), .ZN(n5314) );
  AOI211_X1 U6355 ( .C1(n5318), .C2(INSTADDRPOINTER_REG_25__SCAN_IN), .A(n5315), .B(n5314), .ZN(n5316) );
  OAI211_X1 U6356 ( .C1(n5848), .C2(n5431), .A(n5317), .B(n5316), .ZN(U2993)
         );
  INV_X1 U6357 ( .A(n5433), .ZN(n5323) );
  INV_X1 U6358 ( .A(n5318), .ZN(n5321) );
  AOI21_X1 U6359 ( .B1(n5326), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(
        INSTADDRPOINTER_REG_24__SCAN_IN), .ZN(n5320) );
  OAI21_X1 U6360 ( .B1(n5321), .B2(n5320), .A(n5319), .ZN(n5322) );
  AOI21_X1 U6361 ( .B1(n5323), .B2(n5834), .A(n5322), .ZN(n5324) );
  OAI21_X1 U6362 ( .B1(n5325), .B2(n5824), .A(n5324), .ZN(U2994) );
  INV_X1 U6363 ( .A(n5326), .ZN(n5328) );
  OAI21_X1 U6364 ( .B1(n5328), .B2(INSTADDRPOINTER_REG_23__SCAN_IN), .A(n5327), 
        .ZN(n5330) );
  NOR2_X1 U6365 ( .A1(n5449), .A2(n5848), .ZN(n5329) );
  AOI211_X1 U6366 ( .C1(INSTADDRPOINTER_REG_23__SCAN_IN), .C2(n5331), .A(n5330), .B(n5329), .ZN(n5332) );
  OAI21_X1 U6367 ( .B1(n5333), .B2(n5824), .A(n5332), .ZN(U2995) );
  INV_X1 U6368 ( .A(n5350), .ZN(n5340) );
  INV_X1 U6369 ( .A(n5346), .ZN(n5337) );
  NOR3_X1 U6370 ( .A1(n5337), .A2(n5336), .A3(n5335), .ZN(n5338) );
  AOI211_X1 U6371 ( .C1(n5340), .C2(INSTADDRPOINTER_REG_22__SCAN_IN), .A(n5339), .B(n5338), .ZN(n5341) );
  OAI211_X1 U6372 ( .C1(n5848), .C2(n5343), .A(n5342), .B(n5341), .ZN(U2996)
         );
  XNOR2_X1 U6373 ( .A(n5345), .B(n5344), .ZN(n5466) );
  NAND2_X1 U6374 ( .A1(n5346), .A2(n5349), .ZN(n5347) );
  OAI211_X1 U6375 ( .C1(n5350), .C2(n5349), .A(n5348), .B(n5347), .ZN(n5351)
         );
  AOI21_X1 U6376 ( .B1(n5466), .B2(n5834), .A(n5351), .ZN(n5352) );
  OAI21_X1 U6377 ( .B1(n5353), .B2(n5824), .A(n5352), .ZN(U2997) );
  OR2_X1 U6378 ( .A1(n5852), .A2(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5359)
         );
  AND2_X1 U6379 ( .A1(INSTADDRPOINTER_REG_17__SCAN_IN), .A2(n5354), .ZN(n5355)
         );
  OR2_X1 U6380 ( .A1(n5356), .A2(n5355), .ZN(n5357) );
  NAND2_X1 U6381 ( .A1(n5358), .A2(n5357), .ZN(n5386) );
  AOI21_X1 U6382 ( .B1(n5841), .B2(n5504), .A(n5386), .ZN(n5511) );
  AND2_X1 U6383 ( .A1(n5359), .A2(n5511), .ZN(n5374) );
  AOI21_X1 U6384 ( .B1(n6854), .B2(n5364), .A(n5360), .ZN(n5361) );
  NAND2_X1 U6385 ( .A1(n5372), .A2(n5361), .ZN(n5362) );
  OAI211_X1 U6386 ( .C1(n5374), .C2(n5364), .A(n5363), .B(n5362), .ZN(n5365)
         );
  AOI21_X1 U6387 ( .B1(n5366), .B2(n5834), .A(n5365), .ZN(n5367) );
  OAI21_X1 U6388 ( .B1(n5368), .B2(n5824), .A(n5367), .ZN(U2998) );
  AOI21_X1 U6389 ( .B1(INSTADDRPOINTER_REG_19__SCAN_IN), .B2(n5370), .A(n5369), 
        .ZN(n5371) );
  XNOR2_X1 U6390 ( .A(n5371), .B(n3685), .ZN(n5496) );
  INV_X1 U6391 ( .A(n5496), .ZN(n5378) );
  INV_X1 U6392 ( .A(n5465), .ZN(n5376) );
  AOI22_X1 U6393 ( .A1(n5832), .A2(REIP_REG_19__SCAN_IN), .B1(n5372), .B2(
        n6854), .ZN(n5373) );
  OAI21_X1 U6394 ( .B1(n5374), .B2(n6854), .A(n5373), .ZN(n5375) );
  AOI21_X1 U6395 ( .B1(n5376), .B2(n5834), .A(n5375), .ZN(n5377) );
  OAI21_X1 U6396 ( .B1(n5378), .B2(n5824), .A(n5377), .ZN(U2999) );
  AOI21_X1 U6397 ( .B1(n3680), .B2(n5504), .A(n5244), .ZN(n5379) );
  AOI21_X1 U6398 ( .B1(INSTADDRPOINTER_REG_17__SCAN_IN), .B2(n5380), .A(n5379), 
        .ZN(n5384) );
  INV_X1 U6399 ( .A(n5381), .ZN(n5382) );
  OAI21_X1 U6400 ( .B1(n5384), .B2(n5383), .A(n5382), .ZN(n5500) );
  AOI22_X1 U6401 ( .A1(n5832), .A2(REIP_REG_17__SCAN_IN), .B1(n5385), .B2(
        n5504), .ZN(n5388) );
  NAND2_X1 U6402 ( .A1(n5386), .A2(INSTADDRPOINTER_REG_17__SCAN_IN), .ZN(n5387) );
  OAI211_X1 U6403 ( .C1(n5582), .C2(n5848), .A(n5388), .B(n5387), .ZN(n5389)
         );
  AOI21_X1 U6404 ( .B1(n5500), .B2(n5854), .A(n5389), .ZN(n5390) );
  INV_X1 U6405 ( .A(n5390), .ZN(U3001) );
  INV_X1 U6406 ( .A(n5517), .ZN(n5391) );
  OAI21_X1 U6407 ( .B1(n5391), .B2(n5852), .A(n5785), .ZN(n5515) );
  OAI22_X1 U6408 ( .A1(n5585), .A2(n5848), .B1(n6565), .B2(n5811), .ZN(n5392)
         );
  NOR3_X1 U6409 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n5786), .A3(n5517), 
        .ZN(n5516) );
  AOI211_X1 U6410 ( .C1(n5515), .C2(INSTADDRPOINTER_REG_15__SCAN_IN), .A(n5392), .B(n5516), .ZN(n5393) );
  OAI21_X1 U6411 ( .B1(n5394), .B2(n5824), .A(n5393), .ZN(U3003) );
  INV_X1 U6412 ( .A(n4543), .ZN(n6017) );
  OAI211_X1 U6413 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n4688), .A(n6247), .B(
        n6419), .ZN(n5395) );
  OAI21_X1 U6414 ( .B1(n5396), .B2(n6017), .A(n5395), .ZN(n5397) );
  MUX2_X1 U6415 ( .A(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), .B(n5397), .S(n5860), 
        .Z(U3464) );
  INV_X1 U6416 ( .A(n3776), .ZN(n5403) );
  INV_X1 U6417 ( .A(n5863), .ZN(n5398) );
  NOR3_X1 U6418 ( .A1(n6110), .A2(n6410), .A3(n6247), .ZN(n5399) );
  AOI21_X1 U6419 ( .B1(n5400), .B2(n6211), .A(n5399), .ZN(n5401) );
  OAI21_X1 U6420 ( .B1(n5403), .B2(n5402), .A(n5401), .ZN(n5404) );
  MUX2_X1 U6421 ( .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .B(n5404), .S(n5860), 
        .Z(U3462) );
  AND2_X1 U6422 ( .A1(n5743), .A2(DATAO_REG_31__SCAN_IN), .ZN(U2892) );
  NOR2_X1 U6423 ( .A1(n5405), .A2(n5691), .ZN(n5408) );
  OAI22_X1 U6424 ( .A1(n5406), .A2(n5692), .B1(n6580), .B2(n5414), .ZN(n5407)
         );
  AOI211_X1 U6425 ( .C1(n5693), .C2(EBX_REG_27__SCAN_IN), .A(n5408), .B(n5407), 
        .ZN(n5411) );
  AOI22_X1 U6426 ( .A1(n5469), .A2(n5631), .B1(n5409), .B2(n6580), .ZN(n5410)
         );
  OAI211_X1 U6427 ( .C1(n5412), .C2(n5681), .A(n5411), .B(n5410), .ZN(U2800)
         );
  AOI22_X1 U6428 ( .A1(PHYADDRPOINTER_REG_26__SCAN_IN), .A2(n5674), .B1(n5413), 
        .B2(n5677), .ZN(n5420) );
  INV_X1 U6429 ( .A(REIP_REG_24__SCAN_IN), .ZN(n6578) );
  NOR2_X1 U6430 ( .A1(n6578), .A2(n5428), .ZN(n5421) );
  AOI21_X1 U6431 ( .B1(REIP_REG_25__SCAN_IN), .B2(n5421), .A(
        REIP_REG_26__SCAN_IN), .ZN(n5415) );
  OAI22_X1 U6432 ( .A1(n5416), .A2(n5620), .B1(n5415), .B2(n5414), .ZN(n5417)
         );
  AOI21_X1 U6433 ( .B1(n5418), .B2(n5690), .A(n5417), .ZN(n5419) );
  OAI211_X1 U6434 ( .C1(n6868), .C2(n5665), .A(n5420), .B(n5419), .ZN(U2801)
         );
  INV_X1 U6435 ( .A(n5421), .ZN(n5425) );
  INV_X1 U6436 ( .A(PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5422) );
  OAI22_X1 U6437 ( .A1(n5422), .A2(n5692), .B1(n5691), .B2(n5494), .ZN(n5423)
         );
  AOI21_X1 U6438 ( .B1(n5693), .B2(EBX_REG_25__SCAN_IN), .A(n5423), .ZN(n5424)
         );
  OAI21_X1 U6439 ( .B1(n5425), .B2(REIP_REG_25__SCAN_IN), .A(n5424), .ZN(n5426) );
  AOI21_X1 U6440 ( .B1(n5491), .B2(n5631), .A(n5426), .ZN(n5430) );
  AND2_X1 U6441 ( .A1(n5427), .A2(n5688), .ZN(n5446) );
  NOR2_X1 U6442 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5428), .ZN(n5435) );
  OAI21_X1 U6443 ( .B1(n5446), .B2(n5435), .A(REIP_REG_25__SCAN_IN), .ZN(n5429) );
  OAI211_X1 U6444 ( .C1(n5431), .C2(n5681), .A(n5430), .B(n5429), .ZN(U2802)
         );
  AOI22_X1 U6445 ( .A1(EBX_REG_24__SCAN_IN), .A2(n5693), .B1(
        PHYADDRPOINTER_REG_24__SCAN_IN), .B2(n5674), .ZN(n5439) );
  AOI22_X1 U6446 ( .A1(REIP_REG_24__SCAN_IN), .A2(n5446), .B1(n5432), .B2(
        n5677), .ZN(n5438) );
  OAI22_X1 U6447 ( .A1(n5474), .A2(n5620), .B1(n5433), .B2(n5681), .ZN(n5434)
         );
  INV_X1 U6448 ( .A(n5434), .ZN(n5437) );
  INV_X1 U6449 ( .A(n5435), .ZN(n5436) );
  NAND4_X1 U6450 ( .A1(n5439), .A2(n5438), .A3(n5437), .A4(n5436), .ZN(U2803)
         );
  INV_X1 U6451 ( .A(PHYADDRPOINTER_REG_23__SCAN_IN), .ZN(n5441) );
  OAI22_X1 U6452 ( .A1(n5441), .A2(n5692), .B1(n5440), .B2(n5691), .ZN(n5442)
         );
  AOI21_X1 U6453 ( .B1(EBX_REG_23__SCAN_IN), .B2(n5693), .A(n5442), .ZN(n5448)
         );
  INV_X1 U6454 ( .A(REIP_REG_22__SCAN_IN), .ZN(n6576) );
  INV_X1 U6455 ( .A(REIP_REG_23__SCAN_IN), .ZN(n5443) );
  OAI21_X1 U6456 ( .B1(n6576), .B2(n5444), .A(n5443), .ZN(n5445) );
  AOI22_X1 U6457 ( .A1(n5478), .A2(n5631), .B1(n5446), .B2(n5445), .ZN(n5447)
         );
  OAI211_X1 U6458 ( .C1(n5449), .C2(n5681), .A(n5448), .B(n5447), .ZN(U2804)
         );
  AOI22_X1 U6459 ( .A1(EBX_REG_21__SCAN_IN), .A2(n5693), .B1(
        PHYADDRPOINTER_REG_21__SCAN_IN), .B2(n5674), .ZN(n5456) );
  INV_X1 U6460 ( .A(n5450), .ZN(n5452) );
  AOI22_X1 U6461 ( .A1(n5452), .A2(n5677), .B1(REIP_REG_21__SCAN_IN), .B2(
        n5451), .ZN(n5455) );
  AOI22_X1 U6462 ( .A1(n5481), .A2(n5631), .B1(n5690), .B2(n5466), .ZN(n5454)
         );
  NAND4_X1 U6463 ( .A1(n5456), .A2(n5455), .A3(n5454), .A4(n5453), .ZN(U2806)
         );
  INV_X1 U6464 ( .A(PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5459) );
  INV_X1 U6465 ( .A(REIP_REG_19__SCAN_IN), .ZN(n6738) );
  OAI22_X1 U6466 ( .A1(n5499), .A2(n5691), .B1(n6738), .B2(n5577), .ZN(n5457)
         );
  AOI21_X1 U6467 ( .B1(EBX_REG_19__SCAN_IN), .B2(n5693), .A(n5457), .ZN(n5458)
         );
  OAI211_X1 U6468 ( .C1(n5459), .C2(n5692), .A(n5458), .B(n5640), .ZN(n5460)
         );
  AOI21_X1 U6469 ( .B1(n5495), .B2(n5631), .A(n5460), .ZN(n5464) );
  OAI211_X1 U6470 ( .C1(REIP_REG_19__SCAN_IN), .C2(REIP_REG_18__SCAN_IN), .A(
        n5462), .B(n5461), .ZN(n5463) );
  OAI211_X1 U6471 ( .C1(n5465), .C2(n5681), .A(n5464), .B(n5463), .ZN(U2808)
         );
  INV_X1 U6472 ( .A(EBX_REG_21__SCAN_IN), .ZN(n6722) );
  AOI22_X1 U6473 ( .A1(n5481), .A2(n5703), .B1(n4502), .B2(n5466), .ZN(n5467)
         );
  OAI21_X1 U6474 ( .B1(n5706), .B2(n6722), .A(n5467), .ZN(U2838) );
  AOI22_X1 U6475 ( .A1(n5469), .A2(n5708), .B1(n5707), .B2(DATAI_27_), .ZN(
        n5471) );
  AOI22_X1 U6476 ( .A1(n5711), .A2(DATAI_11_), .B1(EAX_REG_27__SCAN_IN), .B2(
        n5710), .ZN(n5470) );
  NAND2_X1 U6477 ( .A1(n5471), .A2(n5470), .ZN(U2864) );
  AOI22_X1 U6478 ( .A1(n5491), .A2(n5708), .B1(n5707), .B2(DATAI_25_), .ZN(
        n5473) );
  AOI22_X1 U6479 ( .A1(n5711), .A2(DATAI_9_), .B1(EAX_REG_25__SCAN_IN), .B2(
        n5710), .ZN(n5472) );
  NAND2_X1 U6480 ( .A1(n5473), .A2(n5472), .ZN(U2866) );
  INV_X1 U6481 ( .A(n5474), .ZN(n5475) );
  AOI22_X1 U6482 ( .A1(n5475), .A2(n5708), .B1(n5707), .B2(DATAI_24_), .ZN(
        n5477) );
  AOI22_X1 U6483 ( .A1(n5711), .A2(DATAI_8_), .B1(EAX_REG_24__SCAN_IN), .B2(
        n5710), .ZN(n5476) );
  NAND2_X1 U6484 ( .A1(n5477), .A2(n5476), .ZN(U2867) );
  AOI22_X1 U6485 ( .A1(n5478), .A2(n5708), .B1(n5707), .B2(DATAI_23_), .ZN(
        n5480) );
  AOI22_X1 U6486 ( .A1(n5711), .A2(DATAI_7_), .B1(EAX_REG_23__SCAN_IN), .B2(
        n5710), .ZN(n5479) );
  NAND2_X1 U6487 ( .A1(n5480), .A2(n5479), .ZN(U2868) );
  AOI22_X1 U6488 ( .A1(n5481), .A2(n5708), .B1(n5707), .B2(DATAI_21_), .ZN(
        n5483) );
  AOI22_X1 U6489 ( .A1(n5711), .A2(DATAI_5_), .B1(EAX_REG_21__SCAN_IN), .B2(
        n5710), .ZN(n5482) );
  NAND2_X1 U6490 ( .A1(n5483), .A2(n5482), .ZN(U2870) );
  INV_X1 U6491 ( .A(n5484), .ZN(n5485) );
  AOI22_X1 U6492 ( .A1(n5485), .A2(n5708), .B1(n5707), .B2(DATAI_20_), .ZN(
        n5487) );
  AOI22_X1 U6493 ( .A1(n5711), .A2(DATAI_4_), .B1(EAX_REG_20__SCAN_IN), .B2(
        n5710), .ZN(n5486) );
  NAND2_X1 U6494 ( .A1(n5487), .A2(n5486), .ZN(U2871) );
  AOI22_X1 U6495 ( .A1(n5495), .A2(n5708), .B1(n5707), .B2(DATAI_19_), .ZN(
        n5489) );
  AOI22_X1 U6496 ( .A1(n5711), .A2(DATAI_3_), .B1(EAX_REG_19__SCAN_IN), .B2(
        n5710), .ZN(n5488) );
  NAND2_X1 U6497 ( .A1(n5489), .A2(n5488), .ZN(U2872) );
  AOI22_X1 U6498 ( .A1(n5832), .A2(REIP_REG_25__SCAN_IN), .B1(n5777), .B2(
        PHYADDRPOINTER_REG_25__SCAN_IN), .ZN(n5493) );
  AOI22_X1 U6499 ( .A1(n5491), .A2(n5768), .B1(n5774), .B2(n5490), .ZN(n5492)
         );
  OAI211_X1 U6500 ( .C1(n5773), .C2(n5494), .A(n5493), .B(n5492), .ZN(U2961)
         );
  AOI22_X1 U6501 ( .A1(n5832), .A2(REIP_REG_19__SCAN_IN), .B1(n5777), .B2(
        PHYADDRPOINTER_REG_19__SCAN_IN), .ZN(n5498) );
  AOI22_X1 U6502 ( .A1(n5496), .A2(n5774), .B1(n5768), .B2(n5495), .ZN(n5497)
         );
  OAI211_X1 U6503 ( .C1(n5773), .C2(n5499), .A(n5498), .B(n5497), .ZN(U2967)
         );
  AOI22_X1 U6504 ( .A1(n5832), .A2(REIP_REG_17__SCAN_IN), .B1(n5777), .B2(
        PHYADDRPOINTER_REG_17__SCAN_IN), .ZN(n5502) );
  AOI22_X1 U6505 ( .A1(n5500), .A2(n5774), .B1(n5768), .B2(n5709), .ZN(n5501)
         );
  OAI211_X1 U6506 ( .C1(n5773), .C2(n5575), .A(n5502), .B(n5501), .ZN(U2969)
         );
  INV_X1 U6507 ( .A(INSTADDRPOINTER_REG_18__SCAN_IN), .ZN(n5510) );
  NOR3_X1 U6508 ( .A1(INSTADDRPOINTER_REG_18__SCAN_IN), .A2(n5504), .A3(n5503), 
        .ZN(n5505) );
  AOI21_X1 U6509 ( .B1(REIP_REG_18__SCAN_IN), .B2(n5832), .A(n5505), .ZN(n5509) );
  AOI22_X1 U6510 ( .A1(n5507), .A2(n5854), .B1(n5834), .B2(n5506), .ZN(n5508)
         );
  OAI211_X1 U6511 ( .C1(n5511), .C2(n5510), .A(n5509), .B(n5508), .ZN(U3000)
         );
  OAI22_X1 U6512 ( .A1(n5513), .A2(n5824), .B1(n5848), .B2(n5512), .ZN(n5514)
         );
  INV_X1 U6513 ( .A(n5514), .ZN(n5522) );
  NAND2_X1 U6514 ( .A1(n5832), .A2(REIP_REG_16__SCAN_IN), .ZN(n5521) );
  OAI21_X1 U6515 ( .B1(n5516), .B2(n5515), .A(INSTADDRPOINTER_REG_16__SCAN_IN), 
        .ZN(n5520) );
  NOR2_X1 U6516 ( .A1(n5786), .A2(n5517), .ZN(n5518) );
  NAND3_X1 U6517 ( .A1(INSTADDRPOINTER_REG_15__SCAN_IN), .A2(n5518), .A3(n6828), .ZN(n5519) );
  NAND4_X1 U6518 ( .A1(n5522), .A2(n5521), .A3(n5520), .A4(n5519), .ZN(U3002)
         );
  AOI21_X1 U6519 ( .B1(n5524), .B2(n5834), .A(n5523), .ZN(n5538) );
  OR2_X1 U6520 ( .A1(n6661), .A2(INSTADDRPOINTER_REG_13__SCAN_IN), .ZN(n5541)
         );
  AND2_X1 U6521 ( .A1(n5526), .A2(n5525), .ZN(n5530) );
  OAI21_X1 U6522 ( .B1(n5535), .B2(n5527), .A(n5785), .ZN(n5528) );
  AOI21_X1 U6523 ( .B1(n6661), .B2(n5529), .A(n5528), .ZN(n5546) );
  OAI21_X1 U6524 ( .B1(n5541), .B2(n5530), .A(n5546), .ZN(n5531) );
  AOI22_X1 U6525 ( .A1(n5532), .A2(n5854), .B1(INSTADDRPOINTER_REG_14__SCAN_IN), .B2(n5531), .ZN(n5537) );
  NAND3_X1 U6526 ( .A1(n5535), .A2(n5534), .A3(n5533), .ZN(n5536) );
  NAND3_X1 U6527 ( .A1(n5538), .A2(n5537), .A3(n5536), .ZN(U3004) );
  AOI22_X1 U6528 ( .A1(n5539), .A2(n5834), .B1(n5832), .B2(
        REIP_REG_13__SCAN_IN), .ZN(n5540) );
  OAI21_X1 U6529 ( .B1(n5786), .B2(n5541), .A(n5540), .ZN(n5542) );
  AOI21_X1 U6530 ( .B1(n5543), .B2(n5854), .A(n5542), .ZN(n5544) );
  OAI21_X1 U6531 ( .B1(n5546), .B2(n5545), .A(n5544), .ZN(U3005) );
  NAND3_X1 U6532 ( .A1(n5655), .A2(n6606), .A3(n5547), .ZN(n5549) );
  OAI22_X1 U6533 ( .A1(n5550), .A2(n5549), .B1(n5548), .B2(n6612), .ZN(U3455)
         );
  INV_X1 U6534 ( .A(STATE_REG_2__SCAN_IN), .ZN(n6550) );
  AOI21_X1 U6535 ( .B1(STATE_REG_1__SCAN_IN), .B2(n6550), .A(n6541), .ZN(n5555) );
  INV_X1 U6536 ( .A(ADS_N_REG_SCAN_IN), .ZN(n5551) );
  AOI21_X1 U6537 ( .B1(n5555), .B2(n5551), .A(n6625), .ZN(U2789) );
  OAI21_X1 U6538 ( .B1(n5552), .B2(n6525), .A(CODEFETCH_REG_SCAN_IN), .ZN(
        n5553) );
  OAI21_X1 U6539 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6524), .A(n5553), .ZN(
        U2790) );
  INV_X2 U6540 ( .A(n6625), .ZN(n6636) );
  NOR2_X1 U6541 ( .A1(STATE_REG_2__SCAN_IN), .A2(STATE_REG_0__SCAN_IN), .ZN(
        n5556) );
  OAI21_X1 U6542 ( .B1(D_C_N_REG_SCAN_IN), .B2(n5556), .A(n6636), .ZN(n5554)
         );
  OAI21_X1 U6543 ( .B1(CODEFETCH_REG_SCAN_IN), .B2(n6636), .A(n5554), .ZN(
        U2791) );
  NOR2_X2 U6544 ( .A1(n6625), .A2(n5555), .ZN(n6594) );
  OAI21_X1 U6545 ( .B1(n5556), .B2(BS16_N), .A(n6594), .ZN(n6592) );
  OAI21_X1 U6546 ( .B1(n6594), .B2(n6286), .A(n6592), .ZN(U2792) );
  OAI21_X1 U6547 ( .B1(n5559), .B2(n5558), .A(n5557), .ZN(U2793) );
  NOR4_X1 U6548 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(
        DATAWIDTH_REG_27__SCAN_IN), .A3(DATAWIDTH_REG_28__SCAN_IN), .A4(
        DATAWIDTH_REG_29__SCAN_IN), .ZN(n5563) );
  NOR4_X1 U6549 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(DATAWIDTH_REG_9__SCAN_IN), 
        .A3(DATAWIDTH_REG_7__SCAN_IN), .A4(DATAWIDTH_REG_8__SCAN_IN), .ZN(
        n5562) );
  NOR4_X1 U6550 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(
        DATAWIDTH_REG_23__SCAN_IN), .A3(DATAWIDTH_REG_21__SCAN_IN), .A4(
        DATAWIDTH_REG_22__SCAN_IN), .ZN(n5561) );
  NOR4_X1 U6551 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(
        DATAWIDTH_REG_11__SCAN_IN), .A3(DATAWIDTH_REG_16__SCAN_IN), .A4(
        DATAWIDTH_REG_17__SCAN_IN), .ZN(n5560) );
  NAND4_X1 U6552 ( .A1(n5563), .A2(n5562), .A3(n5561), .A4(n5560), .ZN(n5568)
         );
  INV_X1 U6553 ( .A(DATAWIDTH_REG_12__SCAN_IN), .ZN(n6781) );
  INV_X1 U6554 ( .A(DATAWIDTH_REG_13__SCAN_IN), .ZN(n6772) );
  INV_X1 U6555 ( .A(DATAWIDTH_REG_14__SCAN_IN), .ZN(n6782) );
  INV_X1 U6556 ( .A(DATAWIDTH_REG_24__SCAN_IN), .ZN(n6702) );
  NAND4_X1 U6557 ( .A1(n6781), .A2(n6772), .A3(n6782), .A4(n6702), .ZN(n6662)
         );
  AOI211_X1 U6558 ( .C1(DATAWIDTH_REG_0__SCAN_IN), .C2(
        DATAWIDTH_REG_1__SCAN_IN), .A(DATAWIDTH_REG_25__SCAN_IN), .B(n6662), 
        .ZN(n5566) );
  NOR4_X1 U6559 ( .A1(DATAWIDTH_REG_19__SCAN_IN), .A2(
        DATAWIDTH_REG_20__SCAN_IN), .A3(DATAWIDTH_REG_2__SCAN_IN), .A4(
        DATAWIDTH_REG_4__SCAN_IN), .ZN(n5565) );
  NOR4_X1 U6560 ( .A1(DATAWIDTH_REG_10__SCAN_IN), .A2(DATAWIDTH_REG_3__SCAN_IN), .A3(DATAWIDTH_REG_31__SCAN_IN), .A4(DATAWIDTH_REG_5__SCAN_IN), .ZN(n5564) );
  INV_X1 U6561 ( .A(DATAWIDTH_REG_15__SCAN_IN), .ZN(n6813) );
  NAND4_X1 U6562 ( .A1(n5566), .A2(n5565), .A3(n5564), .A4(n6813), .ZN(n5567)
         );
  NOR2_X1 U6563 ( .A1(n5568), .A2(n5567), .ZN(n6620) );
  INV_X1 U6564 ( .A(BYTEENABLE_REG_1__SCAN_IN), .ZN(n5570) );
  NOR3_X1 U6565 ( .A1(DATAWIDTH_REG_0__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), 
        .A3(DATAWIDTH_REG_1__SCAN_IN), .ZN(n5571) );
  OAI21_X1 U6566 ( .B1(REIP_REG_1__SCAN_IN), .B2(n5571), .A(n6620), .ZN(n5569)
         );
  OAI21_X1 U6567 ( .B1(n6620), .B2(n5570), .A(n5569), .ZN(U2794) );
  INV_X1 U6568 ( .A(REIP_REG_1__SCAN_IN), .ZN(n6616) );
  INV_X1 U6569 ( .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6593) );
  AOI21_X1 U6570 ( .B1(n6616), .B2(n6593), .A(n5571), .ZN(n5573) );
  INV_X1 U6571 ( .A(BYTEENABLE_REG_3__SCAN_IN), .ZN(n5572) );
  INV_X1 U6572 ( .A(n6620), .ZN(n6623) );
  AOI22_X1 U6573 ( .A1(n6620), .A2(n5573), .B1(n5572), .B2(n6623), .ZN(U2795)
         );
  AOI22_X1 U6574 ( .A1(EBX_REG_17__SCAN_IN), .A2(n5693), .B1(
        PHYADDRPOINTER_REG_17__SCAN_IN), .B2(n5674), .ZN(n5574) );
  OAI211_X1 U6575 ( .C1(n5691), .C2(n5575), .A(n5640), .B(n5574), .ZN(n5576)
         );
  AOI21_X1 U6576 ( .B1(n5709), .B2(n5631), .A(n5576), .ZN(n5581) );
  INV_X1 U6577 ( .A(n5577), .ZN(n5578) );
  OAI21_X1 U6578 ( .B1(REIP_REG_17__SCAN_IN), .B2(n5579), .A(n5578), .ZN(n5580) );
  OAI211_X1 U6579 ( .C1(n5582), .C2(n5681), .A(n5581), .B(n5580), .ZN(U2810)
         );
  AOI22_X1 U6580 ( .A1(EBX_REG_15__SCAN_IN), .A2(n5693), .B1(
        REIP_REG_15__SCAN_IN), .B2(n5583), .ZN(n5584) );
  OAI21_X1 U6581 ( .B1(n5681), .B2(n5585), .A(n5584), .ZN(n5586) );
  AOI211_X1 U6582 ( .C1(n5674), .C2(PHYADDRPOINTER_REG_15__SCAN_IN), .A(n5651), 
        .B(n5586), .ZN(n5590) );
  AOI22_X1 U6583 ( .A1(n5588), .A2(n5631), .B1(n5677), .B2(n5587), .ZN(n5589)
         );
  OAI211_X1 U6584 ( .C1(REIP_REG_15__SCAN_IN), .C2(n5591), .A(n5590), .B(n5589), .ZN(U2812) );
  INV_X1 U6585 ( .A(REIP_REG_12__SCAN_IN), .ZN(n6560) );
  INV_X1 U6586 ( .A(PHYADDRPOINTER_REG_12__SCAN_IN), .ZN(n5592) );
  NOR2_X1 U6587 ( .A1(n5692), .A2(n5592), .ZN(n5593) );
  AOI211_X1 U6588 ( .C1(n5693), .C2(EBX_REG_12__SCAN_IN), .A(n5651), .B(n5593), 
        .ZN(n5596) );
  NAND2_X1 U6589 ( .A1(n5594), .A2(n5690), .ZN(n5595) );
  OAI211_X1 U6590 ( .C1(n5597), .C2(n5620), .A(n5596), .B(n5595), .ZN(n5598)
         );
  AOI21_X1 U6591 ( .B1(n5599), .B2(n5677), .A(n5598), .ZN(n5600) );
  OAI221_X1 U6592 ( .B1(REIP_REG_12__SCAN_IN), .B2(n5602), .C1(n6560), .C2(
        n5601), .A(n5600), .ZN(U2815) );
  OAI22_X1 U6593 ( .A1(n5702), .A2(n5665), .B1(n5603), .B2(n5692), .ZN(n5604)
         );
  AOI211_X1 U6594 ( .C1(REIP_REG_10__SCAN_IN), .C2(n5605), .A(n5651), .B(n5604), .ZN(n5612) );
  AOI22_X1 U6595 ( .A1(n5700), .A2(n5631), .B1(n5677), .B2(n5606), .ZN(n5611)
         );
  NAND2_X1 U6596 ( .A1(REIP_REG_9__SCAN_IN), .A2(REIP_REG_10__SCAN_IN), .ZN(
        n5607) );
  OAI211_X1 U6597 ( .C1(REIP_REG_9__SCAN_IN), .C2(REIP_REG_10__SCAN_IN), .A(
        n5608), .B(n5607), .ZN(n5610) );
  NAND2_X1 U6598 ( .A1(n5690), .A2(n5699), .ZN(n5609) );
  NAND4_X1 U6599 ( .A1(n5612), .A2(n5611), .A3(n5610), .A4(n5609), .ZN(U2817)
         );
  OAI22_X1 U6600 ( .A1(REIP_REG_7__SCAN_IN), .A2(n5614), .B1(n5681), .B2(n5613), .ZN(n5615) );
  AOI211_X1 U6601 ( .C1(n5674), .C2(PHYADDRPOINTER_REG_7__SCAN_IN), .A(n5651), 
        .B(n5615), .ZN(n5624) );
  INV_X1 U6602 ( .A(n5618), .ZN(n5616) );
  OR2_X1 U6603 ( .A1(n5653), .A2(n5616), .ZN(n5617) );
  AND2_X1 U6604 ( .A1(n5617), .A2(n5687), .ZN(n5626) );
  INV_X1 U6605 ( .A(n5626), .ZN(n5646) );
  NOR3_X1 U6606 ( .A1(n5653), .A2(REIP_REG_6__SCAN_IN), .A3(n5618), .ZN(n5628)
         );
  OAI22_X1 U6607 ( .A1(n5621), .A2(n5620), .B1(n5619), .B2(n5691), .ZN(n5622)
         );
  AOI221_X1 U6608 ( .B1(n5646), .B2(REIP_REG_7__SCAN_IN), .C1(n5628), .C2(
        REIP_REG_7__SCAN_IN), .A(n5622), .ZN(n5623) );
  OAI211_X1 U6609 ( .C1(n5625), .C2(n5665), .A(n5624), .B(n5623), .ZN(U2820)
         );
  AOI22_X1 U6610 ( .A1(PHYADDRPOINTER_REG_6__SCAN_IN), .A2(n5674), .B1(n5690), 
        .B2(n5803), .ZN(n5635) );
  NOR2_X1 U6611 ( .A1(n6557), .A2(n5626), .ZN(n5627) );
  AOI211_X1 U6612 ( .C1(n5693), .C2(EBX_REG_6__SCAN_IN), .A(n5628), .B(n5627), 
        .ZN(n5634) );
  INV_X1 U6613 ( .A(n5629), .ZN(n5632) );
  AOI22_X1 U6614 ( .A1(n5632), .A2(n5631), .B1(n5630), .B2(n5677), .ZN(n5633)
         );
  NAND4_X1 U6615 ( .A1(n5635), .A2(n5634), .A3(n5633), .A4(n5640), .ZN(U2821)
         );
  INV_X1 U6616 ( .A(n5636), .ZN(n5638) );
  INV_X1 U6617 ( .A(REIP_REG_5__SCAN_IN), .ZN(n5637) );
  OAI21_X1 U6618 ( .B1(n5653), .B2(n5638), .A(n5637), .ZN(n5647) );
  AOI22_X1 U6619 ( .A1(EBX_REG_5__SCAN_IN), .A2(n5693), .B1(
        PHYADDRPOINTER_REG_5__SCAN_IN), .B2(n5674), .ZN(n5639) );
  OAI211_X1 U6620 ( .C1(n5681), .C2(n5641), .A(n5640), .B(n5639), .ZN(n5645)
         );
  OAI22_X1 U6621 ( .A1(n5643), .A2(n5698), .B1(n5642), .B2(n5691), .ZN(n5644)
         );
  AOI211_X1 U6622 ( .C1(n5647), .C2(n5646), .A(n5645), .B(n5644), .ZN(n5648)
         );
  INV_X1 U6623 ( .A(n5648), .ZN(U2822) );
  OAI21_X1 U6624 ( .B1(n5649), .B2(n5652), .A(n5688), .ZN(n5673) );
  OAI22_X1 U6625 ( .A1(n5673), .A2(n6929), .B1(n6837), .B2(n5692), .ZN(n5650)
         );
  AOI211_X1 U6626 ( .C1(n5693), .C2(EBX_REG_4__SCAN_IN), .A(n5651), .B(n5650), 
        .ZN(n5660) );
  INV_X1 U6627 ( .A(n5698), .ZN(n5683) );
  NOR3_X1 U6628 ( .A1(n5653), .A2(REIP_REG_4__SCAN_IN), .A3(n5652), .ZN(n5654)
         );
  AOI21_X1 U6629 ( .B1(n5655), .B2(n5694), .A(n5654), .ZN(n5656) );
  OAI21_X1 U6630 ( .B1(n5681), .B2(n5812), .A(n5656), .ZN(n5657) );
  AOI21_X1 U6631 ( .B1(n5658), .B2(n5683), .A(n5657), .ZN(n5659) );
  OAI211_X1 U6632 ( .C1(n5661), .C2(n5691), .A(n5660), .B(n5659), .ZN(U2823)
         );
  INV_X1 U6633 ( .A(REIP_REG_3__SCAN_IN), .ZN(n6553) );
  INV_X1 U6634 ( .A(n5662), .ZN(n5663) );
  NAND2_X1 U6635 ( .A1(n5663), .A2(REIP_REG_2__SCAN_IN), .ZN(n5672) );
  OAI22_X1 U6636 ( .A1(n3780), .A2(n5692), .B1(n5691), .B2(n5664), .ZN(n5667)
         );
  OAI22_X1 U6637 ( .A1(n6863), .A2(n5665), .B1(n5681), .B2(n5822), .ZN(n5666)
         );
  AOI211_X1 U6638 ( .C1(n5694), .C2(n6211), .A(n5667), .B(n5666), .ZN(n5668)
         );
  OAI21_X1 U6639 ( .B1(n5669), .B2(n5698), .A(n5668), .ZN(n5670) );
  INV_X1 U6640 ( .A(n5670), .ZN(n5671) );
  OAI221_X1 U6641 ( .B1(n5673), .B2(n6553), .C1(n5673), .C2(n5672), .A(n5671), 
        .ZN(U2824) );
  AOI22_X1 U6642 ( .A1(EBX_REG_1__SCAN_IN), .A2(n5693), .B1(
        PHYADDRPOINTER_REG_1__SCAN_IN), .B2(n5674), .ZN(n5686) );
  INV_X1 U6643 ( .A(n5675), .ZN(n5680) );
  AOI22_X1 U6644 ( .A1(n5694), .A2(n4543), .B1(n5677), .B2(n5676), .ZN(n5679)
         );
  OAI211_X1 U6645 ( .C1(n5681), .C2(n5680), .A(n5679), .B(n5678), .ZN(n5682)
         );
  AOI21_X1 U6646 ( .B1(n5684), .B2(n5683), .A(n5682), .ZN(n5685) );
  OAI211_X1 U6647 ( .C1(n5687), .C2(n6616), .A(n5686), .B(n5685), .ZN(U2826)
         );
  AOI22_X1 U6648 ( .A1(n5690), .A2(n5689), .B1(REIP_REG_0__SCAN_IN), .B2(n5688), .ZN(n5697) );
  NAND2_X1 U6649 ( .A1(n5692), .A2(n5691), .ZN(n5695) );
  AOI222_X1 U6650 ( .A1(n5695), .A2(PHYADDRPOINTER_REG_0__SCAN_IN), .B1(n5694), 
        .B2(n6179), .C1(EBX_REG_0__SCAN_IN), .C2(n5693), .ZN(n5696) );
  OAI211_X1 U6651 ( .C1(n5698), .C2(n5780), .A(n5697), .B(n5696), .ZN(U2827)
         );
  AOI22_X1 U6652 ( .A1(n5700), .A2(n5703), .B1(n4502), .B2(n5699), .ZN(n5701)
         );
  OAI21_X1 U6653 ( .B1(n5706), .B2(n5702), .A(n5701), .ZN(U2849) );
  AOI22_X1 U6654 ( .A1(n5769), .A2(n5703), .B1(n4502), .B2(n5833), .ZN(n5704)
         );
  OAI21_X1 U6655 ( .B1(n5706), .B2(n5705), .A(n5704), .ZN(U2857) );
  AOI22_X1 U6656 ( .A1(n5709), .A2(n5708), .B1(n5707), .B2(DATAI_17_), .ZN(
        n5713) );
  AOI22_X1 U6657 ( .A1(n5711), .A2(DATAI_1_), .B1(EAX_REG_17__SCAN_IN), .B2(
        n5710), .ZN(n5712) );
  NAND2_X1 U6658 ( .A1(n5713), .A2(n5712), .ZN(U2874) );
  INV_X1 U6659 ( .A(DATAO_REG_30__SCAN_IN), .ZN(n6684) );
  AOI22_X1 U6660 ( .A1(n5722), .A2(EAX_REG_30__SCAN_IN), .B1(
        UWORD_REG_14__SCAN_IN), .B2(n5738), .ZN(n5715) );
  OAI21_X1 U6661 ( .B1(n6684), .B2(n5749), .A(n5715), .ZN(U2893) );
  INV_X1 U6662 ( .A(UWORD_REG_13__SCAN_IN), .ZN(n6851) );
  AOI22_X1 U6663 ( .A1(n5743), .A2(DATAO_REG_29__SCAN_IN), .B1(n5722), .B2(
        EAX_REG_29__SCAN_IN), .ZN(n5716) );
  OAI21_X1 U6664 ( .B1(n6851), .B2(n5746), .A(n5716), .ZN(U2894) );
  INV_X1 U6665 ( .A(DATAO_REG_28__SCAN_IN), .ZN(n6795) );
  AOI22_X1 U6666 ( .A1(n5722), .A2(EAX_REG_28__SCAN_IN), .B1(n5738), .B2(
        UWORD_REG_12__SCAN_IN), .ZN(n5717) );
  OAI21_X1 U6667 ( .B1(n6795), .B2(n5749), .A(n5717), .ZN(U2895) );
  AOI22_X1 U6668 ( .A1(n5743), .A2(DATAO_REG_26__SCAN_IN), .B1(n5722), .B2(
        EAX_REG_26__SCAN_IN), .ZN(n5718) );
  OAI21_X1 U6669 ( .B1(n6879), .B2(n5746), .A(n5718), .ZN(U2897) );
  INV_X1 U6670 ( .A(UWORD_REG_5__SCAN_IN), .ZN(n6914) );
  AOI22_X1 U6671 ( .A1(n5743), .A2(DATAO_REG_21__SCAN_IN), .B1(n5722), .B2(
        EAX_REG_21__SCAN_IN), .ZN(n5719) );
  OAI21_X1 U6672 ( .B1(n6914), .B2(n5746), .A(n5719), .ZN(U2902) );
  INV_X1 U6673 ( .A(UWORD_REG_3__SCAN_IN), .ZN(n6787) );
  AOI22_X1 U6674 ( .A1(n5743), .A2(DATAO_REG_19__SCAN_IN), .B1(n5722), .B2(
        EAX_REG_19__SCAN_IN), .ZN(n5720) );
  OAI21_X1 U6675 ( .B1(n6787), .B2(n5746), .A(n5720), .ZN(U2904) );
  INV_X1 U6676 ( .A(DATAO_REG_18__SCAN_IN), .ZN(n6822) );
  AOI22_X1 U6677 ( .A1(n5722), .A2(EAX_REG_18__SCAN_IN), .B1(n5738), .B2(
        UWORD_REG_2__SCAN_IN), .ZN(n5721) );
  OAI21_X1 U6678 ( .B1(n6822), .B2(n5749), .A(n5721), .ZN(U2905) );
  AOI22_X1 U6679 ( .A1(n5743), .A2(DATAO_REG_16__SCAN_IN), .B1(n5722), .B2(
        EAX_REG_16__SCAN_IN), .ZN(n5723) );
  OAI21_X1 U6680 ( .B1(n6816), .B2(n5746), .A(n5723), .ZN(U2907) );
  INV_X1 U6681 ( .A(EAX_REG_15__SCAN_IN), .ZN(n5763) );
  AOI22_X1 U6682 ( .A1(n5738), .A2(LWORD_REG_15__SCAN_IN), .B1(n5743), .B2(
        DATAO_REG_15__SCAN_IN), .ZN(n5724) );
  OAI21_X1 U6683 ( .B1(n5763), .B2(n5748), .A(n5724), .ZN(U2908) );
  AOI22_X1 U6684 ( .A1(n5738), .A2(LWORD_REG_14__SCAN_IN), .B1(n5743), .B2(
        DATAO_REG_14__SCAN_IN), .ZN(n5725) );
  OAI21_X1 U6685 ( .B1(n3935), .B2(n5748), .A(n5725), .ZN(U2909) );
  AOI22_X1 U6686 ( .A1(n5738), .A2(LWORD_REG_13__SCAN_IN), .B1(n5743), .B2(
        DATAO_REG_13__SCAN_IN), .ZN(n5726) );
  OAI21_X1 U6687 ( .B1(n5727), .B2(n5748), .A(n5726), .ZN(U2910) );
  AOI22_X1 U6688 ( .A1(n5738), .A2(LWORD_REG_12__SCAN_IN), .B1(n5743), .B2(
        DATAO_REG_12__SCAN_IN), .ZN(n5728) );
  OAI21_X1 U6689 ( .B1(n5729), .B2(n5748), .A(n5728), .ZN(U2911) );
  INV_X1 U6690 ( .A(LWORD_REG_11__SCAN_IN), .ZN(n6819) );
  INV_X1 U6691 ( .A(DATAO_REG_11__SCAN_IN), .ZN(n6770) );
  OAI222_X1 U6692 ( .A1(n5746), .A2(n6819), .B1(n5748), .B2(n6757), .C1(n6770), 
        .C2(n5749), .ZN(U2912) );
  INV_X1 U6693 ( .A(DATAO_REG_10__SCAN_IN), .ZN(n6838) );
  AOI22_X1 U6694 ( .A1(EAX_REG_10__SCAN_IN), .A2(n5739), .B1(n5738), .B2(
        LWORD_REG_10__SCAN_IN), .ZN(n5730) );
  OAI21_X1 U6695 ( .B1(n6838), .B2(n5749), .A(n5730), .ZN(U2913) );
  AOI222_X1 U6696 ( .A1(n5743), .A2(DATAO_REG_9__SCAN_IN), .B1(n5739), .B2(
        EAX_REG_9__SCAN_IN), .C1(n5738), .C2(LWORD_REG_9__SCAN_IN), .ZN(n5731)
         );
  INV_X1 U6697 ( .A(n5731), .ZN(U2914) );
  INV_X1 U6698 ( .A(DATAO_REG_8__SCAN_IN), .ZN(n6703) );
  AOI22_X1 U6699 ( .A1(EAX_REG_8__SCAN_IN), .A2(n5739), .B1(n5738), .B2(
        LWORD_REG_8__SCAN_IN), .ZN(n5732) );
  OAI21_X1 U6700 ( .B1(n6703), .B2(n5749), .A(n5732), .ZN(U2915) );
  INV_X1 U6701 ( .A(LWORD_REG_7__SCAN_IN), .ZN(n6905) );
  AOI22_X1 U6702 ( .A1(EAX_REG_7__SCAN_IN), .A2(n5739), .B1(n5743), .B2(
        DATAO_REG_7__SCAN_IN), .ZN(n5733) );
  OAI21_X1 U6703 ( .B1(n6905), .B2(n5746), .A(n5733), .ZN(U2916) );
  AOI22_X1 U6704 ( .A1(n5738), .A2(LWORD_REG_6__SCAN_IN), .B1(n5743), .B2(
        DATAO_REG_6__SCAN_IN), .ZN(n5734) );
  OAI21_X1 U6705 ( .B1(n3808), .B2(n5748), .A(n5734), .ZN(U2917) );
  AOI22_X1 U6706 ( .A1(n5738), .A2(LWORD_REG_5__SCAN_IN), .B1(n5743), .B2(
        DATAO_REG_5__SCAN_IN), .ZN(n5735) );
  OAI21_X1 U6707 ( .B1(n5736), .B2(n5748), .A(n5735), .ZN(U2918) );
  AOI222_X1 U6708 ( .A1(n5743), .A2(DATAO_REG_4__SCAN_IN), .B1(n5739), .B2(
        EAX_REG_4__SCAN_IN), .C1(n5738), .C2(LWORD_REG_4__SCAN_IN), .ZN(n5737)
         );
  INV_X1 U6709 ( .A(n5737), .ZN(U2919) );
  AOI222_X1 U6710 ( .A1(n5743), .A2(DATAO_REG_3__SCAN_IN), .B1(n5739), .B2(
        EAX_REG_3__SCAN_IN), .C1(n5738), .C2(LWORD_REG_3__SCAN_IN), .ZN(n5740)
         );
  INV_X1 U6711 ( .A(n5740), .ZN(U2920) );
  AOI22_X1 U6712 ( .A1(n5738), .A2(LWORD_REG_2__SCAN_IN), .B1(n5743), .B2(
        DATAO_REG_2__SCAN_IN), .ZN(n5741) );
  OAI21_X1 U6713 ( .B1(n5742), .B2(n5748), .A(n5741), .ZN(U2921) );
  AOI22_X1 U6714 ( .A1(n5738), .A2(LWORD_REG_1__SCAN_IN), .B1(n5743), .B2(
        DATAO_REG_1__SCAN_IN), .ZN(n5744) );
  OAI21_X1 U6715 ( .B1(n5745), .B2(n5748), .A(n5744), .ZN(U2922) );
  INV_X1 U6716 ( .A(DATAO_REG_0__SCAN_IN), .ZN(n6919) );
  INV_X1 U6717 ( .A(LWORD_REG_0__SCAN_IN), .ZN(n6848) );
  OAI222_X1 U6718 ( .A1(n5749), .A2(n6919), .B1(n5748), .B2(n5747), .C1(n5746), 
        .C2(n6848), .ZN(U2923) );
  NAND2_X1 U6719 ( .A1(n5759), .A2(DATAI_8_), .ZN(n5754) );
  INV_X1 U6720 ( .A(n5754), .ZN(n5750) );
  AOI21_X1 U6721 ( .B1(UWORD_REG_8__SCAN_IN), .B2(n5753), .A(n5750), .ZN(n5751) );
  OAI21_X1 U6722 ( .B1(n5752), .B2(n5762), .A(n5751), .ZN(U2932) );
  AOI22_X1 U6723 ( .A1(n5753), .A2(LWORD_REG_8__SCAN_IN), .B1(
        EAX_REG_8__SCAN_IN), .B2(n5756), .ZN(n5755) );
  NAND2_X1 U6724 ( .A1(n5755), .A2(n5754), .ZN(U2947) );
  AOI22_X1 U6725 ( .A1(n5760), .A2(LWORD_REG_10__SCAN_IN), .B1(
        EAX_REG_10__SCAN_IN), .B2(n5756), .ZN(n5758) );
  NAND2_X1 U6726 ( .A1(n5758), .A2(n5757), .ZN(U2949) );
  AOI22_X1 U6727 ( .A1(n5760), .A2(LWORD_REG_15__SCAN_IN), .B1(n5759), .B2(
        DATAI_15_), .ZN(n5761) );
  OAI21_X1 U6728 ( .B1(n5763), .B2(n5762), .A(n5761), .ZN(U2954) );
  AOI22_X1 U6729 ( .A1(n5832), .A2(REIP_REG_2__SCAN_IN), .B1(n5777), .B2(
        PHYADDRPOINTER_REG_2__SCAN_IN), .ZN(n5771) );
  NAND2_X1 U6730 ( .A1(n5765), .A2(n5764), .ZN(n5766) );
  XOR2_X1 U6731 ( .A(n5767), .B(n5766), .Z(n5839) );
  AOI22_X1 U6732 ( .A1(n5839), .A2(n5774), .B1(n5769), .B2(n5768), .ZN(n5770)
         );
  OAI211_X1 U6733 ( .C1(n5773), .C2(n5772), .A(n5771), .B(n5770), .ZN(U2984)
         );
  AOI22_X1 U6734 ( .A1(n5775), .A2(n5774), .B1(n5832), .B2(REIP_REG_0__SCAN_IN), .ZN(n5779) );
  OAI21_X1 U6735 ( .B1(n5777), .B2(n5776), .A(PHYADDRPOINTER_REG_0__SCAN_IN), 
        .ZN(n5778) );
  OAI211_X1 U6736 ( .C1(n5780), .C2(n5911), .A(n5779), .B(n5778), .ZN(U2986)
         );
  OAI22_X1 U6737 ( .A1(n5781), .A2(n5848), .B1(n4884), .B2(n5811), .ZN(n5782)
         );
  AOI21_X1 U6738 ( .B1(n5783), .B2(n5854), .A(n5782), .ZN(n5784) );
  OAI221_X1 U6739 ( .B1(INSTADDRPOINTER_REG_11__SCAN_IN), .B2(n5786), .C1(
        n6798), .C2(n5785), .A(n5784), .ZN(U3007) );
  AOI21_X1 U6740 ( .B1(n5788), .B2(n5834), .A(n5787), .ZN(n5792) );
  AOI22_X1 U6741 ( .A1(n5790), .A2(n5854), .B1(INSTADDRPOINTER_REG_9__SCAN_IN), 
        .B2(n5789), .ZN(n5791) );
  OAI211_X1 U6742 ( .C1(INSTADDRPOINTER_REG_9__SCAN_IN), .C2(n5793), .A(n5792), 
        .B(n5791), .ZN(U3009) );
  NOR2_X1 U6743 ( .A1(n5794), .A2(n6759), .ZN(n5797) );
  OAI22_X1 U6744 ( .A1(n5795), .A2(n5848), .B1(n6767), .B2(n5811), .ZN(n5796)
         );
  AOI211_X1 U6745 ( .C1(n5798), .C2(n5854), .A(n5797), .B(n5796), .ZN(n5802)
         );
  OAI211_X1 U6746 ( .C1(INSTADDRPOINTER_REG_7__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A(n5800), .B(n5799), .ZN(n5801) );
  NAND2_X1 U6747 ( .A1(n5802), .A2(n5801), .ZN(U3010) );
  AOI22_X1 U6748 ( .A1(n5803), .A2(n5834), .B1(n5832), .B2(REIP_REG_6__SCAN_IN), .ZN(n5804) );
  OAI21_X1 U6749 ( .B1(n5805), .B2(INSTADDRPOINTER_REG_6__SCAN_IN), .A(n5804), 
        .ZN(n5806) );
  AOI21_X1 U6750 ( .B1(n5807), .B2(n5854), .A(n5806), .ZN(n5808) );
  OAI21_X1 U6751 ( .B1(n5809), .B2(n3655), .A(n5808), .ZN(U3012) );
  OAI211_X1 U6752 ( .C1(INSTADDRPOINTER_REG_3__SCAN_IN), .C2(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A(n5819), .B(n5820), .ZN(n5817) );
  INV_X1 U6753 ( .A(n5810), .ZN(n5838) );
  AOI21_X1 U6754 ( .B1(n5835), .B2(n5837), .A(n5838), .ZN(n5831) );
  NOR2_X1 U6755 ( .A1(n5831), .A2(n3627), .ZN(n5814) );
  OAI22_X1 U6756 ( .A1(n5848), .A2(n5812), .B1(n6929), .B2(n5811), .ZN(n5813)
         );
  AOI211_X1 U6757 ( .C1(n5815), .C2(n5854), .A(n5814), .B(n5813), .ZN(n5816)
         );
  OAI21_X1 U6758 ( .B1(n5818), .B2(n5817), .A(n5816), .ZN(U3014) );
  NAND2_X1 U6759 ( .A1(n5820), .A2(n5819), .ZN(n5828) );
  OAI21_X1 U6760 ( .B1(n5848), .B2(n5822), .A(n5821), .ZN(n5823) );
  INV_X1 U6761 ( .A(n5823), .ZN(n5827) );
  OR2_X1 U6762 ( .A1(n5825), .A2(n5824), .ZN(n5826) );
  OAI211_X1 U6763 ( .C1(n5828), .C2(INSTADDRPOINTER_REG_3__SCAN_IN), .A(n5827), 
        .B(n5826), .ZN(n5829) );
  INV_X1 U6764 ( .A(n5829), .ZN(n5830) );
  OAI21_X1 U6765 ( .B1(n5831), .B2(n3615), .A(n5830), .ZN(U3015) );
  AOI22_X1 U6766 ( .A1(n5834), .A2(n5833), .B1(n5832), .B2(REIP_REG_2__SCAN_IN), .ZN(n5845) );
  OAI221_X1 U6767 ( .B1(n5837), .B2(n5836), .C1(n5837), .C2(
        INSTADDRPOINTER_REG_0__SCAN_IN), .A(n5835), .ZN(n5844) );
  AOI22_X1 U6768 ( .A1(n5839), .A2(n5854), .B1(INSTADDRPOINTER_REG_2__SCAN_IN), 
        .B2(n5838), .ZN(n5843) );
  NAND3_X1 U6769 ( .A1(INSTADDRPOINTER_REG_1__SCAN_IN), .A2(n5841), .A3(n5840), 
        .ZN(n5842) );
  NAND4_X1 U6770 ( .A1(n5845), .A2(n5844), .A3(n5843), .A4(n5842), .ZN(U3016)
         );
  OAI21_X1 U6771 ( .B1(n5848), .B2(n5847), .A(n5846), .ZN(n5849) );
  INV_X1 U6772 ( .A(n5849), .ZN(n5857) );
  INV_X1 U6773 ( .A(n5850), .ZN(n5855) );
  NOR3_X1 U6774 ( .A1(n5852), .A2(INSTADDRPOINTER_REG_1__SCAN_IN), .A3(n5851), 
        .ZN(n5853) );
  AOI21_X1 U6775 ( .B1(n5855), .B2(n5854), .A(n5853), .ZN(n5856) );
  OAI211_X1 U6776 ( .C1(n5859), .C2(n5858), .A(n5857), .B(n5856), .ZN(U3017)
         );
  NOR2_X1 U6777 ( .A1(n5861), .A2(n5860), .ZN(U3019) );
  INV_X1 U6778 ( .A(DATAI_24_), .ZN(n5862) );
  NOR2_X2 U6779 ( .A1(n4535), .A2(n6148), .ZN(n6412) );
  NOR2_X1 U6780 ( .A1(n3119), .A2(n4543), .ZN(n6181) );
  INV_X1 U6781 ( .A(n6181), .ZN(n6147) );
  OR2_X1 U6782 ( .A1(n6211), .A2(n6410), .ZN(n6152) );
  INV_X1 U6783 ( .A(n5871), .ZN(n5864) );
  NOR2_X1 U6784 ( .A1(n5864), .A2(n6511), .ZN(n6367) );
  INV_X1 U6785 ( .A(n6367), .ZN(n6146) );
  INV_X1 U6786 ( .A(n6145), .ZN(n5865) );
  OR2_X1 U6787 ( .A1(n6363), .A2(n5865), .ZN(n6018) );
  OAI22_X1 U6788 ( .A1(n6147), .A2(n6152), .B1(n6146), .B2(n6018), .ZN(n5909)
         );
  INV_X1 U6789 ( .A(n6597), .ZN(n5867) );
  NAND2_X1 U6790 ( .A1(n5907), .A2(n3407), .ZN(n6323) );
  NAND3_X1 U6791 ( .A1(n6368), .A2(n6489), .A3(n6483), .ZN(n5921) );
  NOR2_X1 U6792 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5921), .ZN(n5908)
         );
  AOI22_X1 U6793 ( .A1(n6412), .A2(n5909), .B1(n6411), .B2(n5908), .ZN(n5876)
         );
  INV_X1 U6794 ( .A(n6211), .ZN(n6288) );
  AOI21_X1 U6795 ( .B1(n5945), .B2(n6473), .A(n6286), .ZN(n5869) );
  AOI211_X1 U6796 ( .C1(n6288), .C2(n6181), .A(n6410), .B(n5869), .ZN(n5872)
         );
  INV_X1 U6797 ( .A(n6018), .ZN(n5870) );
  OAI21_X1 U6798 ( .B1(n5870), .B2(n6511), .A(n5956), .ZN(n6022) );
  NOR2_X1 U6799 ( .A1(n5871), .A2(n6511), .ZN(n6364) );
  NOR3_X1 U6800 ( .A1(n5872), .A2(n6022), .A3(n6364), .ZN(n5873) );
  INV_X1 U6801 ( .A(DATAI_16_), .ZN(n5874) );
  OR2_X1 U6802 ( .A1(n5911), .A2(n5874), .ZN(n6424) );
  INV_X1 U6803 ( .A(n6424), .ZN(n6376) );
  AOI22_X1 U6804 ( .A1(INSTQUEUE_REG_0__0__SCAN_IN), .A2(n5913), .B1(n6376), 
        .B2(n5912), .ZN(n5875) );
  OAI211_X1 U6805 ( .C1(n6379), .C2(n6473), .A(n5876), .B(n5875), .ZN(U3020)
         );
  INV_X1 U6806 ( .A(DATAI_25_), .ZN(n5877) );
  OR2_X1 U6807 ( .A1(n5911), .A2(n5877), .ZN(n6953) );
  NOR2_X2 U6808 ( .A1(n4537), .A2(n6148), .ZN(n6957) );
  NAND2_X1 U6809 ( .A1(n5907), .A2(n3397), .ZN(n6951) );
  AOI22_X1 U6810 ( .A1(n6957), .A2(n5909), .B1(n6425), .B2(n5908), .ZN(n5880)
         );
  INV_X1 U6811 ( .A(DATAI_17_), .ZN(n5878) );
  INV_X1 U6812 ( .A(n6962), .ZN(n6380) );
  AOI22_X1 U6813 ( .A1(INSTQUEUE_REG_0__1__SCAN_IN), .A2(n5913), .B1(n6380), 
        .B2(n5912), .ZN(n5879) );
  OAI211_X1 U6814 ( .C1(n6953), .C2(n6473), .A(n5880), .B(n5879), .ZN(U3021)
         );
  INV_X1 U6815 ( .A(DATAI_26_), .ZN(n5881) );
  OR2_X1 U6816 ( .A1(n5911), .A2(n5881), .ZN(n6386) );
  NOR2_X2 U6817 ( .A1(n5882), .A2(n6148), .ZN(n6430) );
  NAND2_X1 U6818 ( .A1(n5907), .A2(n4097), .ZN(n6333) );
  AOI22_X1 U6819 ( .A1(n6430), .A2(n5909), .B1(n6429), .B2(n5908), .ZN(n5885)
         );
  INV_X1 U6820 ( .A(DATAI_18_), .ZN(n5883) );
  OR2_X1 U6821 ( .A1(n5911), .A2(n5883), .ZN(n6434) );
  INV_X1 U6822 ( .A(n6434), .ZN(n6383) );
  AOI22_X1 U6823 ( .A1(INSTQUEUE_REG_0__2__SCAN_IN), .A2(n5913), .B1(n6383), 
        .B2(n5912), .ZN(n5884) );
  OAI211_X1 U6824 ( .C1(n6386), .C2(n6473), .A(n5885), .B(n5884), .ZN(U3022)
         );
  INV_X1 U6825 ( .A(DATAI_27_), .ZN(n5886) );
  OR2_X1 U6826 ( .A1(n5911), .A2(n5886), .ZN(n6437) );
  NOR2_X2 U6827 ( .A1(n5887), .A2(n6148), .ZN(n6436) );
  NAND2_X1 U6828 ( .A1(n5907), .A2(n5888), .ZN(n6339) );
  AOI22_X1 U6829 ( .A1(n6436), .A2(n5909), .B1(n6435), .B2(n5908), .ZN(n5891)
         );
  INV_X1 U6830 ( .A(DATAI_19_), .ZN(n5889) );
  OR2_X1 U6831 ( .A1(n5911), .A2(n5889), .ZN(n6441) );
  INV_X1 U6832 ( .A(n6441), .ZN(n6387) );
  AOI22_X1 U6833 ( .A1(INSTQUEUE_REG_0__3__SCAN_IN), .A2(n5913), .B1(n6387), 
        .B2(n5912), .ZN(n5890) );
  OAI211_X1 U6834 ( .C1(n6437), .C2(n6473), .A(n5891), .B(n5890), .ZN(U3023)
         );
  INV_X1 U6835 ( .A(DATAI_28_), .ZN(n5892) );
  INV_X1 U6836 ( .A(DATAI_4_), .ZN(n6708) );
  NOR2_X2 U6837 ( .A1(n6708), .A2(n6148), .ZN(n6443) );
  NAND2_X1 U6838 ( .A1(n5907), .A2(n3398), .ZN(n6343) );
  AOI22_X1 U6839 ( .A1(n6443), .A2(n5909), .B1(n6442), .B2(n5908), .ZN(n5895)
         );
  INV_X1 U6840 ( .A(DATAI_20_), .ZN(n5893) );
  OR2_X1 U6841 ( .A1(n5911), .A2(n5893), .ZN(n6448) );
  INV_X1 U6842 ( .A(n6448), .ZN(n6390) );
  AOI22_X1 U6843 ( .A1(INSTQUEUE_REG_0__4__SCAN_IN), .A2(n5913), .B1(n6390), 
        .B2(n5912), .ZN(n5894) );
  OAI211_X1 U6844 ( .C1(n6444), .C2(n6473), .A(n5895), .B(n5894), .ZN(U3024)
         );
  INV_X1 U6845 ( .A(DATAI_29_), .ZN(n5896) );
  OR2_X1 U6846 ( .A1(n5911), .A2(n5896), .ZN(n6451) );
  NOR2_X2 U6847 ( .A1(n6785), .A2(n6148), .ZN(n6450) );
  NAND2_X1 U6848 ( .A1(n5907), .A2(n3402), .ZN(n6347) );
  AOI22_X1 U6849 ( .A1(n6450), .A2(n5909), .B1(n6449), .B2(n5908), .ZN(n5899)
         );
  INV_X1 U6850 ( .A(DATAI_21_), .ZN(n5897) );
  OR2_X1 U6851 ( .A1(n5911), .A2(n5897), .ZN(n6455) );
  INV_X1 U6852 ( .A(n6455), .ZN(n6393) );
  AOI22_X1 U6853 ( .A1(INSTQUEUE_REG_0__5__SCAN_IN), .A2(n5913), .B1(n6393), 
        .B2(n5912), .ZN(n5898) );
  OAI211_X1 U6854 ( .C1(n6451), .C2(n6473), .A(n5899), .B(n5898), .ZN(U3025)
         );
  INV_X1 U6855 ( .A(DATAI_30_), .ZN(n5900) );
  OR2_X1 U6856 ( .A1(n5911), .A2(n5900), .ZN(n6458) );
  NOR2_X2 U6857 ( .A1(n5901), .A2(n6148), .ZN(n6457) );
  NAND2_X1 U6858 ( .A1(n5907), .A2(n3410), .ZN(n6351) );
  AOI22_X1 U6859 ( .A1(n6457), .A2(n5909), .B1(n6456), .B2(n5908), .ZN(n5904)
         );
  INV_X1 U6860 ( .A(DATAI_22_), .ZN(n5902) );
  OR2_X1 U6861 ( .A1(n5911), .A2(n5902), .ZN(n6462) );
  INV_X1 U6862 ( .A(n6462), .ZN(n6396) );
  AOI22_X1 U6863 ( .A1(INSTQUEUE_REG_0__6__SCAN_IN), .A2(n5913), .B1(n6396), 
        .B2(n5912), .ZN(n5903) );
  OAI211_X1 U6864 ( .C1(n6458), .C2(n6473), .A(n5904), .B(n5903), .ZN(U3026)
         );
  INV_X1 U6865 ( .A(DATAI_31_), .ZN(n5905) );
  OR2_X1 U6866 ( .A1(n5911), .A2(n5905), .ZN(n6467) );
  NOR2_X2 U6867 ( .A1(n6731), .A2(n6148), .ZN(n6466) );
  NAND2_X1 U6868 ( .A1(n5907), .A2(n5906), .ZN(n6356) );
  AOI22_X1 U6869 ( .A1(n6466), .A2(n5909), .B1(n6463), .B2(n5908), .ZN(n5915)
         );
  INV_X1 U6870 ( .A(DATAI_23_), .ZN(n5910) );
  OR2_X1 U6871 ( .A1(n5911), .A2(n5910), .ZN(n6474) );
  INV_X1 U6872 ( .A(n6474), .ZN(n6401) );
  AOI22_X1 U6873 ( .A1(INSTQUEUE_REG_0__7__SCAN_IN), .A2(n5913), .B1(n6401), 
        .B2(n5912), .ZN(n5914) );
  OAI211_X1 U6874 ( .C1(n6467), .C2(n6473), .A(n5915), .B(n5914), .ZN(U3027)
         );
  NOR2_X1 U6875 ( .A1(n6316), .A2(n5921), .ZN(n5917) );
  INV_X1 U6876 ( .A(n5917), .ZN(n5944) );
  OAI22_X1 U6877 ( .A1(n5978), .A2(n6424), .B1(n6323), .B2(n5944), .ZN(n5916)
         );
  INV_X1 U6878 ( .A(n5916), .ZN(n5925) );
  NOR2_X1 U6879 ( .A1(n6211), .A2(n6477), .ZN(n6048) );
  AOI21_X1 U6880 ( .B1(n6048), .B2(n6181), .A(n5917), .ZN(n5923) );
  NAND2_X1 U6881 ( .A1(n4688), .A2(n6419), .ZN(n5918) );
  AND2_X1 U6882 ( .A1(n6419), .A2(n6286), .ZN(n6415) );
  INV_X1 U6883 ( .A(n6415), .ZN(n5953) );
  NAND2_X1 U6884 ( .A1(n5918), .A2(n5953), .ZN(n6314) );
  AOI21_X1 U6885 ( .B1(n5982), .B2(n6419), .A(n6314), .ZN(n5922) );
  INV_X1 U6886 ( .A(n5922), .ZN(n5919) );
  AOI22_X1 U6887 ( .A1(n5923), .A2(n5919), .B1(n6410), .B2(n5921), .ZN(n5920)
         );
  NAND2_X1 U6888 ( .A1(n6418), .A2(n5920), .ZN(n5948) );
  OAI22_X1 U6889 ( .A1(n5923), .A2(n5922), .B1(n6511), .B2(n5921), .ZN(n5947)
         );
  AOI22_X1 U6890 ( .A1(INSTQUEUE_REG_1__0__SCAN_IN), .A2(n5948), .B1(n6412), 
        .B2(n5947), .ZN(n5924) );
  OAI211_X1 U6891 ( .C1(n6379), .C2(n5945), .A(n5925), .B(n5924), .ZN(U3028)
         );
  OAI22_X1 U6892 ( .A1(n5978), .A2(n6962), .B1(n6951), .B2(n5944), .ZN(n5926)
         );
  INV_X1 U6893 ( .A(n5926), .ZN(n5928) );
  AOI22_X1 U6894 ( .A1(INSTQUEUE_REG_1__1__SCAN_IN), .A2(n5948), .B1(n6957), 
        .B2(n5947), .ZN(n5927) );
  OAI211_X1 U6895 ( .C1(n6953), .C2(n5945), .A(n5928), .B(n5927), .ZN(U3029)
         );
  OAI22_X1 U6896 ( .A1(n5945), .A2(n6386), .B1(n6333), .B2(n5944), .ZN(n5929)
         );
  INV_X1 U6897 ( .A(n5929), .ZN(n5931) );
  AOI22_X1 U6898 ( .A1(INSTQUEUE_REG_1__2__SCAN_IN), .A2(n5948), .B1(n6430), 
        .B2(n5947), .ZN(n5930) );
  OAI211_X1 U6899 ( .C1(n5978), .C2(n6434), .A(n5931), .B(n5930), .ZN(U3030)
         );
  OAI22_X1 U6900 ( .A1(n5945), .A2(n6437), .B1(n6339), .B2(n5944), .ZN(n5932)
         );
  INV_X1 U6901 ( .A(n5932), .ZN(n5934) );
  AOI22_X1 U6902 ( .A1(INSTQUEUE_REG_1__3__SCAN_IN), .A2(n5948), .B1(n6436), 
        .B2(n5947), .ZN(n5933) );
  OAI211_X1 U6903 ( .C1(n5978), .C2(n6441), .A(n5934), .B(n5933), .ZN(U3031)
         );
  OAI22_X1 U6904 ( .A1(n5978), .A2(n6448), .B1(n6343), .B2(n5944), .ZN(n5935)
         );
  INV_X1 U6905 ( .A(n5935), .ZN(n5937) );
  AOI22_X1 U6906 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(n5948), .B1(n6443), 
        .B2(n5947), .ZN(n5936) );
  OAI211_X1 U6907 ( .C1(n6444), .C2(n5945), .A(n5937), .B(n5936), .ZN(U3032)
         );
  OAI22_X1 U6908 ( .A1(n5945), .A2(n6451), .B1(n6347), .B2(n5944), .ZN(n5938)
         );
  INV_X1 U6909 ( .A(n5938), .ZN(n5940) );
  AOI22_X1 U6910 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(n5948), .B1(n6450), 
        .B2(n5947), .ZN(n5939) );
  OAI211_X1 U6911 ( .C1(n5978), .C2(n6455), .A(n5940), .B(n5939), .ZN(U3033)
         );
  OAI22_X1 U6912 ( .A1(n5978), .A2(n6462), .B1(n6351), .B2(n5944), .ZN(n5941)
         );
  INV_X1 U6913 ( .A(n5941), .ZN(n5943) );
  AOI22_X1 U6914 ( .A1(INSTQUEUE_REG_1__6__SCAN_IN), .A2(n5948), .B1(n6457), 
        .B2(n5947), .ZN(n5942) );
  OAI211_X1 U6915 ( .C1(n6458), .C2(n5945), .A(n5943), .B(n5942), .ZN(U3034)
         );
  OAI22_X1 U6916 ( .A1(n5945), .A2(n6467), .B1(n6356), .B2(n5944), .ZN(n5946)
         );
  INV_X1 U6917 ( .A(n5946), .ZN(n5950) );
  AOI22_X1 U6918 ( .A1(INSTQUEUE_REG_1__7__SCAN_IN), .A2(n5948), .B1(n6466), 
        .B2(n5947), .ZN(n5949) );
  OAI211_X1 U6919 ( .C1(n5978), .C2(n6474), .A(n5950), .B(n5949), .ZN(U3035)
         );
  NOR2_X1 U6920 ( .A1(n3119), .A2(n6017), .ZN(n6212) );
  NAND2_X1 U6921 ( .A1(n6288), .A2(n6212), .ZN(n5983) );
  NAND3_X1 U6922 ( .A1(n6367), .A2(n6363), .A3(n6368), .ZN(n5951) );
  OAI21_X1 U6923 ( .B1(n5983), .B2(n6410), .A(n5951), .ZN(n5973) );
  NAND2_X1 U6924 ( .A1(n6208), .A2(n6368), .ZN(n5987) );
  NOR2_X1 U6925 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n5987), .ZN(n5972)
         );
  AOI22_X1 U6926 ( .A1(n6412), .A2(n5973), .B1(n6411), .B2(n5972), .ZN(n5959)
         );
  NAND2_X1 U6927 ( .A1(n4688), .A2(n5952), .ZN(n6207) );
  INV_X1 U6928 ( .A(n6207), .ZN(n6370) );
  INV_X1 U6929 ( .A(n5978), .ZN(n5954) );
  OAI21_X1 U6930 ( .B1(n5974), .B2(n5954), .A(n5953), .ZN(n5955) );
  AOI21_X1 U6931 ( .B1(n5955), .B2(n5983), .A(STATE2_REG_3__SCAN_IN), .ZN(
        n5957) );
  OAI21_X1 U6932 ( .B1(n6363), .B2(n6511), .A(n5956), .ZN(n6369) );
  NOR2_X1 U6933 ( .A1(n6364), .A2(n6369), .ZN(n6214) );
  AOI22_X1 U6934 ( .A1(INSTQUEUE_REG_2__0__SCAN_IN), .A2(n5975), .B1(n6376), 
        .B2(n5974), .ZN(n5958) );
  OAI211_X1 U6935 ( .C1(n6379), .C2(n5978), .A(n5959), .B(n5958), .ZN(U3036)
         );
  AOI22_X1 U6936 ( .A1(n6957), .A2(n5973), .B1(n6425), .B2(n5972), .ZN(n5961)
         );
  AOI22_X1 U6937 ( .A1(INSTQUEUE_REG_2__1__SCAN_IN), .A2(n5975), .B1(n5974), 
        .B2(n6380), .ZN(n5960) );
  OAI211_X1 U6938 ( .C1(n5978), .C2(n6953), .A(n5961), .B(n5960), .ZN(U3037)
         );
  AOI22_X1 U6939 ( .A1(n6430), .A2(n5973), .B1(n6429), .B2(n5972), .ZN(n5963)
         );
  AOI22_X1 U6940 ( .A1(INSTQUEUE_REG_2__2__SCAN_IN), .A2(n5975), .B1(n5974), 
        .B2(n6383), .ZN(n5962) );
  OAI211_X1 U6941 ( .C1(n5978), .C2(n6386), .A(n5963), .B(n5962), .ZN(U3038)
         );
  AOI22_X1 U6942 ( .A1(n6436), .A2(n5973), .B1(n6435), .B2(n5972), .ZN(n5965)
         );
  AOI22_X1 U6943 ( .A1(INSTQUEUE_REG_2__3__SCAN_IN), .A2(n5975), .B1(n5974), 
        .B2(n6387), .ZN(n5964) );
  OAI211_X1 U6944 ( .C1(n5978), .C2(n6437), .A(n5965), .B(n5964), .ZN(U3039)
         );
  AOI22_X1 U6945 ( .A1(n6443), .A2(n5973), .B1(n6442), .B2(n5972), .ZN(n5967)
         );
  AOI22_X1 U6946 ( .A1(INSTQUEUE_REG_2__4__SCAN_IN), .A2(n5975), .B1(n5974), 
        .B2(n6390), .ZN(n5966) );
  OAI211_X1 U6947 ( .C1(n5978), .C2(n6444), .A(n5967), .B(n5966), .ZN(U3040)
         );
  AOI22_X1 U6948 ( .A1(n6450), .A2(n5973), .B1(n6449), .B2(n5972), .ZN(n5969)
         );
  AOI22_X1 U6949 ( .A1(INSTQUEUE_REG_2__5__SCAN_IN), .A2(n5975), .B1(n5974), 
        .B2(n6393), .ZN(n5968) );
  OAI211_X1 U6950 ( .C1(n5978), .C2(n6451), .A(n5969), .B(n5968), .ZN(U3041)
         );
  AOI22_X1 U6951 ( .A1(n6457), .A2(n5973), .B1(n6456), .B2(n5972), .ZN(n5971)
         );
  AOI22_X1 U6952 ( .A1(INSTQUEUE_REG_2__6__SCAN_IN), .A2(n5975), .B1(n5974), 
        .B2(n6396), .ZN(n5970) );
  OAI211_X1 U6953 ( .C1(n5978), .C2(n6458), .A(n5971), .B(n5970), .ZN(U3042)
         );
  AOI22_X1 U6954 ( .A1(n6466), .A2(n5973), .B1(n6463), .B2(n5972), .ZN(n5977)
         );
  AOI22_X1 U6955 ( .A1(INSTQUEUE_REG_2__7__SCAN_IN), .A2(n5975), .B1(n5974), 
        .B2(n6401), .ZN(n5976) );
  OAI211_X1 U6956 ( .C1(n5978), .C2(n6467), .A(n5977), .B(n5976), .ZN(U3043)
         );
  INV_X1 U6957 ( .A(n5980), .ZN(n6245) );
  NAND2_X1 U6958 ( .A1(n6245), .A2(n6368), .ZN(n6010) );
  OAI22_X1 U6959 ( .A1(n6045), .A2(n6424), .B1(n6010), .B2(n6323), .ZN(n5981)
         );
  INV_X1 U6960 ( .A(n5981), .ZN(n5991) );
  OAI21_X1 U6961 ( .B1(n5982), .B2(n6247), .A(n6419), .ZN(n5989) );
  OR2_X1 U6962 ( .A1(n5983), .A2(n6477), .ZN(n5984) );
  NAND2_X1 U6963 ( .A1(n5984), .A2(n6010), .ZN(n5986) );
  NAND2_X1 U6964 ( .A1(n6410), .A2(n5987), .ZN(n5985) );
  OAI211_X1 U6965 ( .C1(n5989), .C2(n5986), .A(n6418), .B(n5985), .ZN(n6014)
         );
  INV_X1 U6966 ( .A(n5986), .ZN(n5988) );
  OAI22_X1 U6967 ( .A1(n5989), .A2(n5988), .B1(n5987), .B2(n6511), .ZN(n6013)
         );
  AOI22_X1 U6968 ( .A1(INSTQUEUE_REG_3__0__SCAN_IN), .A2(n6014), .B1(n6412), 
        .B2(n6013), .ZN(n5990) );
  OAI211_X1 U6969 ( .C1(n6379), .C2(n6011), .A(n5991), .B(n5990), .ZN(U3044)
         );
  OAI22_X1 U6970 ( .A1(n6011), .A2(n6953), .B1(n6010), .B2(n6951), .ZN(n5992)
         );
  INV_X1 U6971 ( .A(n5992), .ZN(n5994) );
  AOI22_X1 U6972 ( .A1(INSTQUEUE_REG_3__1__SCAN_IN), .A2(n6014), .B1(n6957), 
        .B2(n6013), .ZN(n5993) );
  OAI211_X1 U6973 ( .C1(n6962), .C2(n6045), .A(n5994), .B(n5993), .ZN(U3045)
         );
  OAI22_X1 U6974 ( .A1(n6011), .A2(n6386), .B1(n6010), .B2(n6333), .ZN(n5995)
         );
  INV_X1 U6975 ( .A(n5995), .ZN(n5997) );
  AOI22_X1 U6976 ( .A1(INSTQUEUE_REG_3__2__SCAN_IN), .A2(n6014), .B1(n6430), 
        .B2(n6013), .ZN(n5996) );
  OAI211_X1 U6977 ( .C1(n6434), .C2(n6045), .A(n5997), .B(n5996), .ZN(U3046)
         );
  OAI22_X1 U6978 ( .A1(n6045), .A2(n6441), .B1(n6010), .B2(n6339), .ZN(n5998)
         );
  INV_X1 U6979 ( .A(n5998), .ZN(n6000) );
  AOI22_X1 U6980 ( .A1(INSTQUEUE_REG_3__3__SCAN_IN), .A2(n6014), .B1(n6436), 
        .B2(n6013), .ZN(n5999) );
  OAI211_X1 U6981 ( .C1(n6011), .C2(n6437), .A(n6000), .B(n5999), .ZN(U3047)
         );
  OAI22_X1 U6982 ( .A1(n6011), .A2(n6444), .B1(n6010), .B2(n6343), .ZN(n6001)
         );
  INV_X1 U6983 ( .A(n6001), .ZN(n6003) );
  AOI22_X1 U6984 ( .A1(INSTQUEUE_REG_3__4__SCAN_IN), .A2(n6014), .B1(n6443), 
        .B2(n6013), .ZN(n6002) );
  OAI211_X1 U6985 ( .C1(n6448), .C2(n6045), .A(n6003), .B(n6002), .ZN(U3048)
         );
  OAI22_X1 U6986 ( .A1(n6045), .A2(n6455), .B1(n6010), .B2(n6347), .ZN(n6004)
         );
  INV_X1 U6987 ( .A(n6004), .ZN(n6006) );
  AOI22_X1 U6988 ( .A1(INSTQUEUE_REG_3__5__SCAN_IN), .A2(n6014), .B1(n6450), 
        .B2(n6013), .ZN(n6005) );
  OAI211_X1 U6989 ( .C1(n6011), .C2(n6451), .A(n6006), .B(n6005), .ZN(U3049)
         );
  OAI22_X1 U6990 ( .A1(n6045), .A2(n6462), .B1(n6010), .B2(n6351), .ZN(n6007)
         );
  INV_X1 U6991 ( .A(n6007), .ZN(n6009) );
  AOI22_X1 U6992 ( .A1(INSTQUEUE_REG_3__6__SCAN_IN), .A2(n6014), .B1(n6457), 
        .B2(n6013), .ZN(n6008) );
  OAI211_X1 U6993 ( .C1(n6011), .C2(n6458), .A(n6009), .B(n6008), .ZN(U3050)
         );
  OAI22_X1 U6994 ( .A1(n6011), .A2(n6467), .B1(n6010), .B2(n6356), .ZN(n6012)
         );
  INV_X1 U6995 ( .A(n6012), .ZN(n6016) );
  AOI22_X1 U6996 ( .A1(INSTQUEUE_REG_3__7__SCAN_IN), .A2(n6014), .B1(n6466), 
        .B2(n6013), .ZN(n6015) );
  OAI211_X1 U6997 ( .C1(n6474), .C2(n6045), .A(n6016), .B(n6015), .ZN(U3051)
         );
  NAND2_X1 U6998 ( .A1(n3119), .A2(n6017), .ZN(n6287) );
  INV_X1 U6999 ( .A(n6364), .ZN(n6284) );
  OAI22_X1 U7000 ( .A1(n6152), .A2(n6287), .B1(n6284), .B2(n6018), .ZN(n6040)
         );
  NAND3_X1 U7001 ( .A1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .A2(n6368), .A3(n6483), .ZN(n6051) );
  NOR2_X1 U7002 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6051), .ZN(n6039)
         );
  AOI22_X1 U7003 ( .A1(n6412), .A2(n6040), .B1(n6411), .B2(n6039), .ZN(n6026)
         );
  INV_X1 U7004 ( .A(n6045), .ZN(n6019) );
  NOR3_X1 U7005 ( .A1(n6019), .A2(n6041), .A3(n6410), .ZN(n6021) );
  OAI22_X1 U7006 ( .A1(n6021), .A2(n6415), .B1(n6020), .B2(n6287), .ZN(n6024)
         );
  NOR2_X1 U7007 ( .A1(n6367), .A2(n6022), .ZN(n6023) );
  AOI22_X1 U7008 ( .A1(INSTQUEUE_REG_4__0__SCAN_IN), .A2(n6042), .B1(n6376), 
        .B2(n6041), .ZN(n6025) );
  OAI211_X1 U7009 ( .C1(n6379), .C2(n6045), .A(n6026), .B(n6025), .ZN(U3052)
         );
  AOI22_X1 U7010 ( .A1(n6957), .A2(n6040), .B1(n6425), .B2(n6039), .ZN(n6028)
         );
  AOI22_X1 U7011 ( .A1(INSTQUEUE_REG_4__1__SCAN_IN), .A2(n6042), .B1(n6380), 
        .B2(n6041), .ZN(n6027) );
  OAI211_X1 U7012 ( .C1(n6953), .C2(n6045), .A(n6028), .B(n6027), .ZN(U3053)
         );
  AOI22_X1 U7013 ( .A1(n6430), .A2(n6040), .B1(n6429), .B2(n6039), .ZN(n6030)
         );
  AOI22_X1 U7014 ( .A1(INSTQUEUE_REG_4__2__SCAN_IN), .A2(n6042), .B1(n6383), 
        .B2(n6041), .ZN(n6029) );
  OAI211_X1 U7015 ( .C1(n6386), .C2(n6045), .A(n6030), .B(n6029), .ZN(U3054)
         );
  AOI22_X1 U7016 ( .A1(n6436), .A2(n6040), .B1(n6435), .B2(n6039), .ZN(n6032)
         );
  AOI22_X1 U7017 ( .A1(INSTQUEUE_REG_4__3__SCAN_IN), .A2(n6042), .B1(n6387), 
        .B2(n6041), .ZN(n6031) );
  OAI211_X1 U7018 ( .C1(n6437), .C2(n6045), .A(n6032), .B(n6031), .ZN(U3055)
         );
  AOI22_X1 U7019 ( .A1(n6443), .A2(n6040), .B1(n6442), .B2(n6039), .ZN(n6034)
         );
  AOI22_X1 U7020 ( .A1(INSTQUEUE_REG_4__4__SCAN_IN), .A2(n6042), .B1(n6390), 
        .B2(n6041), .ZN(n6033) );
  OAI211_X1 U7021 ( .C1(n6444), .C2(n6045), .A(n6034), .B(n6033), .ZN(U3056)
         );
  AOI22_X1 U7022 ( .A1(n6450), .A2(n6040), .B1(n6449), .B2(n6039), .ZN(n6036)
         );
  AOI22_X1 U7023 ( .A1(INSTQUEUE_REG_4__5__SCAN_IN), .A2(n6042), .B1(n6393), 
        .B2(n6041), .ZN(n6035) );
  OAI211_X1 U7024 ( .C1(n6451), .C2(n6045), .A(n6036), .B(n6035), .ZN(U3057)
         );
  AOI22_X1 U7025 ( .A1(n6457), .A2(n6040), .B1(n6456), .B2(n6039), .ZN(n6038)
         );
  AOI22_X1 U7026 ( .A1(INSTQUEUE_REG_4__6__SCAN_IN), .A2(n6042), .B1(n6396), 
        .B2(n6041), .ZN(n6037) );
  OAI211_X1 U7027 ( .C1(n6458), .C2(n6045), .A(n6038), .B(n6037), .ZN(U3058)
         );
  AOI22_X1 U7028 ( .A1(n6466), .A2(n6040), .B1(n6463), .B2(n6039), .ZN(n6044)
         );
  AOI22_X1 U7029 ( .A1(INSTQUEUE_REG_4__7__SCAN_IN), .A2(n6042), .B1(n6401), 
        .B2(n6041), .ZN(n6043) );
  OAI211_X1 U7030 ( .C1(n6467), .C2(n6045), .A(n6044), .B(n6043), .ZN(U3059)
         );
  NOR2_X1 U7031 ( .A1(n6316), .A2(n6051), .ZN(n6047) );
  INV_X1 U7032 ( .A(n6047), .ZN(n6074) );
  OAI22_X1 U7033 ( .A1(n6080), .A2(n6379), .B1(n6323), .B2(n6074), .ZN(n6046)
         );
  INV_X1 U7034 ( .A(n6046), .ZN(n6055) );
  INV_X1 U7035 ( .A(n6287), .ZN(n6317) );
  AOI21_X1 U7036 ( .B1(n6048), .B2(n6317), .A(n6047), .ZN(n6052) );
  AOI21_X1 U7037 ( .B1(n6110), .B2(n6419), .A(n6314), .ZN(n6053) );
  INV_X1 U7038 ( .A(n6053), .ZN(n6049) );
  AOI22_X1 U7039 ( .A1(n6052), .A2(n6049), .B1(n6410), .B2(n6051), .ZN(n6050)
         );
  NAND2_X1 U7040 ( .A1(n6418), .A2(n6050), .ZN(n6077) );
  OAI22_X1 U7041 ( .A1(n6053), .A2(n6052), .B1(n6511), .B2(n6051), .ZN(n6076)
         );
  AOI22_X1 U7042 ( .A1(INSTQUEUE_REG_5__0__SCAN_IN), .A2(n6077), .B1(n6412), 
        .B2(n6076), .ZN(n6054) );
  OAI211_X1 U7043 ( .C1(n6424), .C2(n6107), .A(n6055), .B(n6054), .ZN(U3060)
         );
  OAI22_X1 U7044 ( .A1(n6080), .A2(n6953), .B1(n6951), .B2(n6074), .ZN(n6056)
         );
  INV_X1 U7045 ( .A(n6056), .ZN(n6058) );
  AOI22_X1 U7046 ( .A1(INSTQUEUE_REG_5__1__SCAN_IN), .A2(n6077), .B1(n6957), 
        .B2(n6076), .ZN(n6057) );
  OAI211_X1 U7047 ( .C1(n6962), .C2(n6107), .A(n6058), .B(n6057), .ZN(U3061)
         );
  OAI22_X1 U7048 ( .A1(n6107), .A2(n6434), .B1(n6333), .B2(n6074), .ZN(n6059)
         );
  INV_X1 U7049 ( .A(n6059), .ZN(n6061) );
  AOI22_X1 U7050 ( .A1(INSTQUEUE_REG_5__2__SCAN_IN), .A2(n6077), .B1(n6430), 
        .B2(n6076), .ZN(n6060) );
  OAI211_X1 U7051 ( .C1(n6386), .C2(n6080), .A(n6061), .B(n6060), .ZN(U3062)
         );
  OAI22_X1 U7052 ( .A1(n6107), .A2(n6441), .B1(n6339), .B2(n6074), .ZN(n6062)
         );
  INV_X1 U7053 ( .A(n6062), .ZN(n6064) );
  AOI22_X1 U7054 ( .A1(INSTQUEUE_REG_5__3__SCAN_IN), .A2(n6077), .B1(n6436), 
        .B2(n6076), .ZN(n6063) );
  OAI211_X1 U7055 ( .C1(n6437), .C2(n6080), .A(n6064), .B(n6063), .ZN(U3063)
         );
  OAI22_X1 U7056 ( .A1(n6080), .A2(n6444), .B1(n6343), .B2(n6074), .ZN(n6065)
         );
  INV_X1 U7057 ( .A(n6065), .ZN(n6067) );
  AOI22_X1 U7058 ( .A1(INSTQUEUE_REG_5__4__SCAN_IN), .A2(n6077), .B1(n6443), 
        .B2(n6076), .ZN(n6066) );
  OAI211_X1 U7059 ( .C1(n6448), .C2(n6107), .A(n6067), .B(n6066), .ZN(U3064)
         );
  OAI22_X1 U7060 ( .A1(n6080), .A2(n6451), .B1(n6347), .B2(n6074), .ZN(n6068)
         );
  INV_X1 U7061 ( .A(n6068), .ZN(n6070) );
  AOI22_X1 U7062 ( .A1(INSTQUEUE_REG_5__5__SCAN_IN), .A2(n6077), .B1(n6450), 
        .B2(n6076), .ZN(n6069) );
  OAI211_X1 U7063 ( .C1(n6455), .C2(n6107), .A(n6070), .B(n6069), .ZN(U3065)
         );
  OAI22_X1 U7064 ( .A1(n6080), .A2(n6458), .B1(n6351), .B2(n6074), .ZN(n6071)
         );
  INV_X1 U7065 ( .A(n6071), .ZN(n6073) );
  AOI22_X1 U7066 ( .A1(INSTQUEUE_REG_5__6__SCAN_IN), .A2(n6077), .B1(n6457), 
        .B2(n6076), .ZN(n6072) );
  OAI211_X1 U7067 ( .C1(n6462), .C2(n6107), .A(n6073), .B(n6072), .ZN(U3066)
         );
  OAI22_X1 U7068 ( .A1(n6107), .A2(n6474), .B1(n6356), .B2(n6074), .ZN(n6075)
         );
  INV_X1 U7069 ( .A(n6075), .ZN(n6079) );
  AOI22_X1 U7070 ( .A1(INSTQUEUE_REG_5__7__SCAN_IN), .A2(n6077), .B1(n6466), 
        .B2(n6076), .ZN(n6078) );
  OAI211_X1 U7071 ( .C1(n6467), .C2(n6080), .A(n6079), .B(n6078), .ZN(U3067)
         );
  AND2_X1 U7072 ( .A1(n3119), .A2(n4543), .ZN(n6407) );
  INV_X1 U7073 ( .A(n6407), .ZN(n6373) );
  NAND3_X1 U7074 ( .A1(n6364), .A2(n6363), .A3(n6368), .ZN(n6081) );
  OAI21_X1 U7075 ( .B1(n6152), .B2(n6373), .A(n6081), .ZN(n6102) );
  NAND2_X1 U7076 ( .A1(n6316), .A2(n3528), .ZN(n6083) );
  INV_X1 U7077 ( .A(n6083), .ZN(n6101) );
  AOI22_X1 U7078 ( .A1(n6412), .A2(n6102), .B1(n6411), .B2(n6101), .ZN(n6088)
         );
  AOI21_X1 U7079 ( .B1(n6107), .B2(n6144), .A(n6286), .ZN(n6086) );
  NAND2_X1 U7080 ( .A1(n6407), .A2(n6082), .ZN(n6111) );
  NAND2_X1 U7081 ( .A1(n6111), .A2(n6419), .ZN(n6085) );
  AOI211_X1 U7082 ( .C1(STATE2_REG_3__SCAN_IN), .C2(n6083), .A(n6367), .B(
        n6369), .ZN(n6084) );
  OAI211_X1 U7083 ( .C1(n6086), .C2(n6085), .A(n6084), .B(n6368), .ZN(n6104)
         );
  AOI22_X1 U7084 ( .A1(INSTQUEUE_REG_6__0__SCAN_IN), .A2(n6104), .B1(n6376), 
        .B2(n6103), .ZN(n6087) );
  OAI211_X1 U7085 ( .C1(n6379), .C2(n6107), .A(n6088), .B(n6087), .ZN(U3068)
         );
  AOI22_X1 U7086 ( .A1(n6957), .A2(n6102), .B1(n6425), .B2(n6101), .ZN(n6090)
         );
  AOI22_X1 U7087 ( .A1(INSTQUEUE_REG_6__1__SCAN_IN), .A2(n6104), .B1(n6380), 
        .B2(n6103), .ZN(n6089) );
  OAI211_X1 U7088 ( .C1(n6953), .C2(n6107), .A(n6090), .B(n6089), .ZN(U3069)
         );
  AOI22_X1 U7089 ( .A1(n6430), .A2(n6102), .B1(n6429), .B2(n6101), .ZN(n6092)
         );
  AOI22_X1 U7090 ( .A1(INSTQUEUE_REG_6__2__SCAN_IN), .A2(n6104), .B1(n6383), 
        .B2(n6103), .ZN(n6091) );
  OAI211_X1 U7091 ( .C1(n6386), .C2(n6107), .A(n6092), .B(n6091), .ZN(U3070)
         );
  AOI22_X1 U7092 ( .A1(n6436), .A2(n6102), .B1(n6435), .B2(n6101), .ZN(n6094)
         );
  AOI22_X1 U7093 ( .A1(INSTQUEUE_REG_6__3__SCAN_IN), .A2(n6104), .B1(n6387), 
        .B2(n6103), .ZN(n6093) );
  OAI211_X1 U7094 ( .C1(n6437), .C2(n6107), .A(n6094), .B(n6093), .ZN(U3071)
         );
  AOI22_X1 U7095 ( .A1(n6443), .A2(n6102), .B1(n6442), .B2(n6101), .ZN(n6096)
         );
  AOI22_X1 U7096 ( .A1(INSTQUEUE_REG_6__4__SCAN_IN), .A2(n6104), .B1(n6390), 
        .B2(n6103), .ZN(n6095) );
  OAI211_X1 U7097 ( .C1(n6444), .C2(n6107), .A(n6096), .B(n6095), .ZN(U3072)
         );
  AOI22_X1 U7098 ( .A1(n6450), .A2(n6102), .B1(n6449), .B2(n6101), .ZN(n6098)
         );
  AOI22_X1 U7099 ( .A1(INSTQUEUE_REG_6__5__SCAN_IN), .A2(n6104), .B1(n6393), 
        .B2(n6103), .ZN(n6097) );
  OAI211_X1 U7100 ( .C1(n6451), .C2(n6107), .A(n6098), .B(n6097), .ZN(U3073)
         );
  AOI22_X1 U7101 ( .A1(n6457), .A2(n6102), .B1(n6456), .B2(n6101), .ZN(n6100)
         );
  AOI22_X1 U7102 ( .A1(INSTQUEUE_REG_6__6__SCAN_IN), .A2(n6104), .B1(n6396), 
        .B2(n6103), .ZN(n6099) );
  OAI211_X1 U7103 ( .C1(n6458), .C2(n6107), .A(n6100), .B(n6099), .ZN(U3074)
         );
  AOI22_X1 U7104 ( .A1(n6466), .A2(n6102), .B1(n6463), .B2(n6101), .ZN(n6106)
         );
  AOI22_X1 U7105 ( .A1(INSTQUEUE_REG_6__7__SCAN_IN), .A2(n6104), .B1(n6401), 
        .B2(n6103), .ZN(n6105) );
  OAI211_X1 U7106 ( .C1(n6467), .C2(n6107), .A(n6106), .B(n6105), .ZN(U3075)
         );
  OAI22_X1 U7107 ( .A1(n6144), .A2(n6379), .B1(n6323), .B2(n6138), .ZN(n6109)
         );
  INV_X1 U7108 ( .A(n6109), .ZN(n6119) );
  OAI21_X1 U7109 ( .B1(n6110), .B2(n6247), .A(n6419), .ZN(n6117) );
  OR2_X1 U7110 ( .A1(n6111), .A2(n6477), .ZN(n6112) );
  NAND2_X1 U7111 ( .A1(n6112), .A2(n6138), .ZN(n6114) );
  OR2_X1 U7112 ( .A1(n6117), .A2(n6114), .ZN(n6113) );
  OAI211_X1 U7113 ( .C1(n3528), .C2(n6419), .A(n6418), .B(n6113), .ZN(n6141)
         );
  INV_X1 U7114 ( .A(n6114), .ZN(n6116) );
  OAI22_X1 U7115 ( .A1(n6117), .A2(n6116), .B1(n6115), .B2(n6511), .ZN(n6140)
         );
  AOI22_X1 U7116 ( .A1(INSTQUEUE_REG_7__0__SCAN_IN), .A2(n6141), .B1(n6412), 
        .B2(n6140), .ZN(n6118) );
  OAI211_X1 U7117 ( .C1(n6424), .C2(n6176), .A(n6119), .B(n6118), .ZN(U3076)
         );
  OAI22_X1 U7118 ( .A1(n6176), .A2(n6962), .B1(n6951), .B2(n6138), .ZN(n6120)
         );
  INV_X1 U7119 ( .A(n6120), .ZN(n6122) );
  AOI22_X1 U7120 ( .A1(INSTQUEUE_REG_7__1__SCAN_IN), .A2(n6141), .B1(n6957), 
        .B2(n6140), .ZN(n6121) );
  OAI211_X1 U7121 ( .C1(n6953), .C2(n6144), .A(n6122), .B(n6121), .ZN(U3077)
         );
  OAI22_X1 U7122 ( .A1(n6144), .A2(n6386), .B1(n6333), .B2(n6138), .ZN(n6123)
         );
  INV_X1 U7123 ( .A(n6123), .ZN(n6125) );
  AOI22_X1 U7124 ( .A1(INSTQUEUE_REG_7__2__SCAN_IN), .A2(n6141), .B1(n6430), 
        .B2(n6140), .ZN(n6124) );
  OAI211_X1 U7125 ( .C1(n6434), .C2(n6176), .A(n6125), .B(n6124), .ZN(U3078)
         );
  OAI22_X1 U7126 ( .A1(n6176), .A2(n6441), .B1(n6339), .B2(n6138), .ZN(n6126)
         );
  INV_X1 U7127 ( .A(n6126), .ZN(n6128) );
  AOI22_X1 U7128 ( .A1(INSTQUEUE_REG_7__3__SCAN_IN), .A2(n6141), .B1(n6436), 
        .B2(n6140), .ZN(n6127) );
  OAI211_X1 U7129 ( .C1(n6437), .C2(n6144), .A(n6128), .B(n6127), .ZN(U3079)
         );
  OAI22_X1 U7130 ( .A1(n6144), .A2(n6444), .B1(n6343), .B2(n6138), .ZN(n6129)
         );
  INV_X1 U7131 ( .A(n6129), .ZN(n6131) );
  AOI22_X1 U7132 ( .A1(INSTQUEUE_REG_7__4__SCAN_IN), .A2(n6141), .B1(n6443), 
        .B2(n6140), .ZN(n6130) );
  OAI211_X1 U7133 ( .C1(n6448), .C2(n6176), .A(n6131), .B(n6130), .ZN(U3080)
         );
  OAI22_X1 U7134 ( .A1(n6176), .A2(n6455), .B1(n6347), .B2(n6138), .ZN(n6132)
         );
  INV_X1 U7135 ( .A(n6132), .ZN(n6134) );
  AOI22_X1 U7136 ( .A1(INSTQUEUE_REG_7__5__SCAN_IN), .A2(n6141), .B1(n6450), 
        .B2(n6140), .ZN(n6133) );
  OAI211_X1 U7137 ( .C1(n6451), .C2(n6144), .A(n6134), .B(n6133), .ZN(U3081)
         );
  OAI22_X1 U7138 ( .A1(n6176), .A2(n6462), .B1(n6351), .B2(n6138), .ZN(n6135)
         );
  INV_X1 U7139 ( .A(n6135), .ZN(n6137) );
  AOI22_X1 U7140 ( .A1(INSTQUEUE_REG_7__6__SCAN_IN), .A2(n6141), .B1(n6457), 
        .B2(n6140), .ZN(n6136) );
  OAI211_X1 U7141 ( .C1(n6458), .C2(n6144), .A(n6137), .B(n6136), .ZN(U3082)
         );
  OAI22_X1 U7142 ( .A1(n6176), .A2(n6474), .B1(n6356), .B2(n6138), .ZN(n6139)
         );
  INV_X1 U7143 ( .A(n6139), .ZN(n6143) );
  AOI22_X1 U7144 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(n6141), .B1(n6466), 
        .B2(n6140), .ZN(n6142) );
  OAI211_X1 U7145 ( .C1(n6467), .C2(n6144), .A(n6143), .B(n6142), .ZN(U3083)
         );
  NAND2_X1 U7146 ( .A1(n6211), .A2(n6419), .ZN(n6366) );
  OR2_X1 U7147 ( .A1(n6363), .A2(n6145), .ZN(n6283) );
  OAI22_X1 U7148 ( .A1(n6147), .A2(n6366), .B1(n6146), .B2(n6283), .ZN(n6171)
         );
  NAND3_X1 U7149 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6489), .A3(n6483), .ZN(n6184) );
  NOR2_X1 U7150 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6184), .ZN(n6170)
         );
  AOI22_X1 U7151 ( .A1(n6412), .A2(n6171), .B1(n6411), .B2(n6170), .ZN(n6157)
         );
  AOI21_X1 U7152 ( .B1(STATE2_REG_2__SCAN_IN), .B2(n6283), .A(n6148), .ZN(
        n6290) );
  INV_X1 U7153 ( .A(n6176), .ZN(n6151) );
  OAI21_X1 U7154 ( .B1(n6172), .B2(n6151), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6154) );
  OAI21_X1 U7155 ( .B1(n6181), .B2(n6410), .A(n6152), .ZN(n6153) );
  AOI21_X1 U7156 ( .B1(n6154), .B2(n6153), .A(n6364), .ZN(n6155) );
  AOI22_X1 U7157 ( .A1(INSTQUEUE_REG_8__0__SCAN_IN), .A2(n6173), .B1(n6376), 
        .B2(n6172), .ZN(n6156) );
  OAI211_X1 U7158 ( .C1(n6379), .C2(n6176), .A(n6157), .B(n6156), .ZN(U3084)
         );
  AOI22_X1 U7159 ( .A1(n6957), .A2(n6171), .B1(n6425), .B2(n6170), .ZN(n6159)
         );
  AOI22_X1 U7160 ( .A1(INSTQUEUE_REG_8__1__SCAN_IN), .A2(n6173), .B1(n6380), 
        .B2(n6172), .ZN(n6158) );
  OAI211_X1 U7161 ( .C1(n6953), .C2(n6176), .A(n6159), .B(n6158), .ZN(U3085)
         );
  AOI22_X1 U7162 ( .A1(n6430), .A2(n6171), .B1(n6429), .B2(n6170), .ZN(n6161)
         );
  AOI22_X1 U7163 ( .A1(INSTQUEUE_REG_8__2__SCAN_IN), .A2(n6173), .B1(n6383), 
        .B2(n6172), .ZN(n6160) );
  OAI211_X1 U7164 ( .C1(n6386), .C2(n6176), .A(n6161), .B(n6160), .ZN(U3086)
         );
  AOI22_X1 U7165 ( .A1(n6436), .A2(n6171), .B1(n6435), .B2(n6170), .ZN(n6163)
         );
  AOI22_X1 U7166 ( .A1(INSTQUEUE_REG_8__3__SCAN_IN), .A2(n6173), .B1(n6387), 
        .B2(n6172), .ZN(n6162) );
  OAI211_X1 U7167 ( .C1(n6437), .C2(n6176), .A(n6163), .B(n6162), .ZN(U3087)
         );
  AOI22_X1 U7168 ( .A1(n6443), .A2(n6171), .B1(n6442), .B2(n6170), .ZN(n6165)
         );
  AOI22_X1 U7169 ( .A1(INSTQUEUE_REG_8__4__SCAN_IN), .A2(n6173), .B1(n6390), 
        .B2(n6172), .ZN(n6164) );
  OAI211_X1 U7170 ( .C1(n6444), .C2(n6176), .A(n6165), .B(n6164), .ZN(U3088)
         );
  AOI22_X1 U7171 ( .A1(n6450), .A2(n6171), .B1(n6449), .B2(n6170), .ZN(n6167)
         );
  AOI22_X1 U7172 ( .A1(INSTQUEUE_REG_8__5__SCAN_IN), .A2(n6173), .B1(n6393), 
        .B2(n6172), .ZN(n6166) );
  OAI211_X1 U7173 ( .C1(n6451), .C2(n6176), .A(n6167), .B(n6166), .ZN(U3089)
         );
  AOI22_X1 U7174 ( .A1(n6457), .A2(n6171), .B1(n6456), .B2(n6170), .ZN(n6169)
         );
  AOI22_X1 U7175 ( .A1(INSTQUEUE_REG_8__6__SCAN_IN), .A2(n6173), .B1(n6396), 
        .B2(n6172), .ZN(n6168) );
  OAI211_X1 U7176 ( .C1(n6458), .C2(n6176), .A(n6169), .B(n6168), .ZN(U3090)
         );
  AOI22_X1 U7177 ( .A1(n6466), .A2(n6171), .B1(n6463), .B2(n6170), .ZN(n6175)
         );
  AOI22_X1 U7178 ( .A1(INSTQUEUE_REG_8__7__SCAN_IN), .A2(n6173), .B1(n6401), 
        .B2(n6172), .ZN(n6174) );
  OAI211_X1 U7179 ( .C1(n6467), .C2(n6176), .A(n6175), .B(n6174), .ZN(U3091)
         );
  NOR2_X1 U7180 ( .A1(n6316), .A2(n6184), .ZN(n6180) );
  INV_X1 U7181 ( .A(n6180), .ZN(n6952) );
  OAI22_X1 U7182 ( .A1(n6954), .A2(n6379), .B1(n6952), .B2(n6323), .ZN(n6178)
         );
  INV_X1 U7183 ( .A(n6178), .ZN(n6188) );
  AND2_X1 U7184 ( .A1(n6211), .A2(n6179), .ZN(n6408) );
  AOI21_X1 U7185 ( .B1(n6408), .B2(n6181), .A(n6180), .ZN(n6186) );
  AOI21_X1 U7186 ( .B1(n6248), .B2(n6419), .A(n6314), .ZN(n6185) );
  INV_X1 U7187 ( .A(n6185), .ZN(n6182) );
  AOI22_X1 U7188 ( .A1(n6186), .A2(n6182), .B1(n6410), .B2(n6184), .ZN(n6183)
         );
  NAND2_X1 U7189 ( .A1(n6418), .A2(n6183), .ZN(n6958) );
  OAI22_X1 U7190 ( .A1(n6186), .A2(n6185), .B1(n6511), .B2(n6184), .ZN(n6956)
         );
  AOI22_X1 U7191 ( .A1(INSTQUEUE_REG_9__0__SCAN_IN), .A2(n6958), .B1(n6412), 
        .B2(n6956), .ZN(n6187) );
  OAI211_X1 U7192 ( .C1(n6424), .C2(n6961), .A(n6188), .B(n6187), .ZN(U3092)
         );
  OAI22_X1 U7193 ( .A1(n6961), .A2(n6434), .B1(n6952), .B2(n6333), .ZN(n6189)
         );
  INV_X1 U7194 ( .A(n6189), .ZN(n6191) );
  AOI22_X1 U7195 ( .A1(INSTQUEUE_REG_9__2__SCAN_IN), .A2(n6958), .B1(n6430), 
        .B2(n6956), .ZN(n6190) );
  OAI211_X1 U7196 ( .C1(n6386), .C2(n6954), .A(n6191), .B(n6190), .ZN(U3094)
         );
  OAI22_X1 U7197 ( .A1(n6961), .A2(n6441), .B1(n6952), .B2(n6339), .ZN(n6192)
         );
  INV_X1 U7198 ( .A(n6192), .ZN(n6194) );
  AOI22_X1 U7199 ( .A1(INSTQUEUE_REG_9__3__SCAN_IN), .A2(n6958), .B1(n6436), 
        .B2(n6956), .ZN(n6193) );
  OAI211_X1 U7200 ( .C1(n6437), .C2(n6954), .A(n6194), .B(n6193), .ZN(U3095)
         );
  OAI22_X1 U7201 ( .A1(n6961), .A2(n6448), .B1(n6952), .B2(n6343), .ZN(n6195)
         );
  INV_X1 U7202 ( .A(n6195), .ZN(n6197) );
  AOI22_X1 U7203 ( .A1(INSTQUEUE_REG_9__4__SCAN_IN), .A2(n6958), .B1(n6443), 
        .B2(n6956), .ZN(n6196) );
  OAI211_X1 U7204 ( .C1(n6444), .C2(n6954), .A(n6197), .B(n6196), .ZN(U3096)
         );
  OAI22_X1 U7205 ( .A1(n6954), .A2(n6451), .B1(n6952), .B2(n6347), .ZN(n6198)
         );
  INV_X1 U7206 ( .A(n6198), .ZN(n6200) );
  AOI22_X1 U7207 ( .A1(INSTQUEUE_REG_9__5__SCAN_IN), .A2(n6958), .B1(n6450), 
        .B2(n6956), .ZN(n6199) );
  OAI211_X1 U7208 ( .C1(n6455), .C2(n6961), .A(n6200), .B(n6199), .ZN(U3097)
         );
  OAI22_X1 U7209 ( .A1(n6961), .A2(n6462), .B1(n6952), .B2(n6351), .ZN(n6201)
         );
  INV_X1 U7210 ( .A(n6201), .ZN(n6203) );
  AOI22_X1 U7211 ( .A1(INSTQUEUE_REG_9__6__SCAN_IN), .A2(n6958), .B1(n6457), 
        .B2(n6956), .ZN(n6202) );
  OAI211_X1 U7212 ( .C1(n6458), .C2(n6954), .A(n6203), .B(n6202), .ZN(U3098)
         );
  OAI22_X1 U7213 ( .A1(n6954), .A2(n6467), .B1(n6952), .B2(n6356), .ZN(n6204)
         );
  INV_X1 U7214 ( .A(n6204), .ZN(n6206) );
  AOI22_X1 U7215 ( .A1(INSTQUEUE_REG_9__7__SCAN_IN), .A2(n6958), .B1(n6466), 
        .B2(n6956), .ZN(n6205) );
  OAI211_X1 U7216 ( .C1(n6474), .C2(n6961), .A(n6206), .B(n6205), .ZN(U3099)
         );
  NAND2_X1 U7217 ( .A1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A2(n6208), .ZN(n6253) );
  OR2_X1 U7218 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6253), .ZN(n6238)
         );
  OAI22_X1 U7219 ( .A1(n6282), .A2(n6424), .B1(n6323), .B2(n6238), .ZN(n6209)
         );
  INV_X1 U7220 ( .A(n6209), .ZN(n6219) );
  AOI21_X1 U7221 ( .B1(n6282), .B2(n6961), .A(n6286), .ZN(n6210) );
  NOR2_X1 U7222 ( .A1(n6210), .A2(n6410), .ZN(n6215) );
  NAND2_X1 U7223 ( .A1(n6212), .A2(n6211), .ZN(n6249) );
  AOI22_X1 U7224 ( .A1(n6215), .A2(n6249), .B1(STATE2_REG_3__SCAN_IN), .B2(
        n6238), .ZN(n6213) );
  OAI211_X1 U7225 ( .C1(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .C2(n6511), .A(n6214), .B(n6213), .ZN(n6241) );
  INV_X1 U7226 ( .A(n6215), .ZN(n6217) );
  NAND3_X1 U7227 ( .A1(n6367), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6363), .ZN(n6216) );
  AOI22_X1 U7228 ( .A1(INSTQUEUE_REG_10__0__SCAN_IN), .A2(n6241), .B1(n6412), 
        .B2(n6240), .ZN(n6218) );
  OAI211_X1 U7229 ( .C1(n6379), .C2(n6961), .A(n6219), .B(n6218), .ZN(U3100)
         );
  OAI22_X1 U7230 ( .A1(n6961), .A2(n6953), .B1(n6238), .B2(n6951), .ZN(n6220)
         );
  INV_X1 U7231 ( .A(n6220), .ZN(n6222) );
  AOI22_X1 U7232 ( .A1(INSTQUEUE_REG_10__1__SCAN_IN), .A2(n6241), .B1(n6957), 
        .B2(n6240), .ZN(n6221) );
  OAI211_X1 U7233 ( .C1(n6962), .C2(n6282), .A(n6222), .B(n6221), .ZN(U3101)
         );
  OAI22_X1 U7234 ( .A1(n6961), .A2(n6386), .B1(n6333), .B2(n6238), .ZN(n6223)
         );
  INV_X1 U7235 ( .A(n6223), .ZN(n6225) );
  AOI22_X1 U7236 ( .A1(INSTQUEUE_REG_10__2__SCAN_IN), .A2(n6241), .B1(n6430), 
        .B2(n6240), .ZN(n6224) );
  OAI211_X1 U7237 ( .C1(n6434), .C2(n6282), .A(n6225), .B(n6224), .ZN(U3102)
         );
  OAI22_X1 U7238 ( .A1(n6961), .A2(n6437), .B1(n6339), .B2(n6238), .ZN(n6226)
         );
  INV_X1 U7239 ( .A(n6226), .ZN(n6228) );
  AOI22_X1 U7240 ( .A1(INSTQUEUE_REG_10__3__SCAN_IN), .A2(n6241), .B1(n6436), 
        .B2(n6240), .ZN(n6227) );
  OAI211_X1 U7241 ( .C1(n6441), .C2(n6282), .A(n6228), .B(n6227), .ZN(U3103)
         );
  OAI22_X1 U7242 ( .A1(n6961), .A2(n6444), .B1(n6343), .B2(n6238), .ZN(n6229)
         );
  INV_X1 U7243 ( .A(n6229), .ZN(n6231) );
  AOI22_X1 U7244 ( .A1(INSTQUEUE_REG_10__4__SCAN_IN), .A2(n6241), .B1(n6443), 
        .B2(n6240), .ZN(n6230) );
  OAI211_X1 U7245 ( .C1(n6448), .C2(n6282), .A(n6231), .B(n6230), .ZN(U3104)
         );
  OAI22_X1 U7246 ( .A1(n6282), .A2(n6455), .B1(n6238), .B2(n6347), .ZN(n6232)
         );
  INV_X1 U7247 ( .A(n6232), .ZN(n6234) );
  AOI22_X1 U7248 ( .A1(INSTQUEUE_REG_10__5__SCAN_IN), .A2(n6241), .B1(n6450), 
        .B2(n6240), .ZN(n6233) );
  OAI211_X1 U7249 ( .C1(n6451), .C2(n6961), .A(n6234), .B(n6233), .ZN(U3105)
         );
  OAI22_X1 U7250 ( .A1(n6961), .A2(n6458), .B1(n6351), .B2(n6238), .ZN(n6235)
         );
  INV_X1 U7251 ( .A(n6235), .ZN(n6237) );
  AOI22_X1 U7252 ( .A1(INSTQUEUE_REG_10__6__SCAN_IN), .A2(n6241), .B1(n6457), 
        .B2(n6240), .ZN(n6236) );
  OAI211_X1 U7253 ( .C1(n6462), .C2(n6282), .A(n6237), .B(n6236), .ZN(U3106)
         );
  OAI22_X1 U7254 ( .A1(n6282), .A2(n6474), .B1(n6238), .B2(n6356), .ZN(n6239)
         );
  INV_X1 U7255 ( .A(n6239), .ZN(n6243) );
  AOI22_X1 U7256 ( .A1(INSTQUEUE_REG_10__7__SCAN_IN), .A2(n6241), .B1(n6466), 
        .B2(n6240), .ZN(n6242) );
  OAI211_X1 U7257 ( .C1(n6467), .C2(n6961), .A(n6243), .B(n6242), .ZN(U3107)
         );
  NAND2_X1 U7258 ( .A1(n6245), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .ZN(n6276) );
  OAI22_X1 U7259 ( .A1(n6313), .A2(n6424), .B1(n6276), .B2(n6323), .ZN(n6246)
         );
  INV_X1 U7260 ( .A(n6246), .ZN(n6257) );
  OAI21_X1 U7261 ( .B1(n6248), .B2(n6247), .A(n6419), .ZN(n6255) );
  OR2_X1 U7262 ( .A1(n6249), .A2(n6477), .ZN(n6250) );
  NAND2_X1 U7263 ( .A1(n6250), .A2(n6276), .ZN(n6252) );
  NAND2_X1 U7264 ( .A1(n6410), .A2(n6253), .ZN(n6251) );
  OAI211_X1 U7265 ( .C1(n6255), .C2(n6252), .A(n6418), .B(n6251), .ZN(n6279)
         );
  INV_X1 U7266 ( .A(n6252), .ZN(n6254) );
  OAI22_X1 U7267 ( .A1(n6255), .A2(n6254), .B1(n6253), .B2(n6511), .ZN(n6278)
         );
  AOI22_X1 U7268 ( .A1(INSTQUEUE_REG_11__0__SCAN_IN), .A2(n6279), .B1(n6412), 
        .B2(n6278), .ZN(n6256) );
  OAI211_X1 U7269 ( .C1(n6379), .C2(n6282), .A(n6257), .B(n6256), .ZN(U3108)
         );
  OAI22_X1 U7270 ( .A1(n6282), .A2(n6953), .B1(n6276), .B2(n6951), .ZN(n6258)
         );
  INV_X1 U7271 ( .A(n6258), .ZN(n6260) );
  AOI22_X1 U7272 ( .A1(INSTQUEUE_REG_11__1__SCAN_IN), .A2(n6279), .B1(n6957), 
        .B2(n6278), .ZN(n6259) );
  OAI211_X1 U7273 ( .C1(n6962), .C2(n6313), .A(n6260), .B(n6259), .ZN(U3109)
         );
  OAI22_X1 U7274 ( .A1(n6282), .A2(n6386), .B1(n6276), .B2(n6333), .ZN(n6261)
         );
  INV_X1 U7275 ( .A(n6261), .ZN(n6263) );
  AOI22_X1 U7276 ( .A1(INSTQUEUE_REG_11__2__SCAN_IN), .A2(n6279), .B1(n6430), 
        .B2(n6278), .ZN(n6262) );
  OAI211_X1 U7277 ( .C1(n6434), .C2(n6313), .A(n6263), .B(n6262), .ZN(U3110)
         );
  OAI22_X1 U7278 ( .A1(n6313), .A2(n6441), .B1(n6276), .B2(n6339), .ZN(n6264)
         );
  INV_X1 U7279 ( .A(n6264), .ZN(n6266) );
  AOI22_X1 U7280 ( .A1(INSTQUEUE_REG_11__3__SCAN_IN), .A2(n6279), .B1(n6436), 
        .B2(n6278), .ZN(n6265) );
  OAI211_X1 U7281 ( .C1(n6437), .C2(n6282), .A(n6266), .B(n6265), .ZN(U3111)
         );
  OAI22_X1 U7282 ( .A1(n6313), .A2(n6448), .B1(n6276), .B2(n6343), .ZN(n6267)
         );
  INV_X1 U7283 ( .A(n6267), .ZN(n6269) );
  AOI22_X1 U7284 ( .A1(INSTQUEUE_REG_11__4__SCAN_IN), .A2(n6279), .B1(n6443), 
        .B2(n6278), .ZN(n6268) );
  OAI211_X1 U7285 ( .C1(n6444), .C2(n6282), .A(n6269), .B(n6268), .ZN(U3112)
         );
  OAI22_X1 U7286 ( .A1(n6282), .A2(n6451), .B1(n6276), .B2(n6347), .ZN(n6270)
         );
  INV_X1 U7287 ( .A(n6270), .ZN(n6272) );
  AOI22_X1 U7288 ( .A1(INSTQUEUE_REG_11__5__SCAN_IN), .A2(n6279), .B1(n6450), 
        .B2(n6278), .ZN(n6271) );
  OAI211_X1 U7289 ( .C1(n6455), .C2(n6313), .A(n6272), .B(n6271), .ZN(U3113)
         );
  OAI22_X1 U7290 ( .A1(n6282), .A2(n6458), .B1(n6276), .B2(n6351), .ZN(n6273)
         );
  INV_X1 U7291 ( .A(n6273), .ZN(n6275) );
  AOI22_X1 U7292 ( .A1(INSTQUEUE_REG_11__6__SCAN_IN), .A2(n6279), .B1(n6457), 
        .B2(n6278), .ZN(n6274) );
  OAI211_X1 U7293 ( .C1(n6462), .C2(n6313), .A(n6275), .B(n6274), .ZN(U3114)
         );
  OAI22_X1 U7294 ( .A1(n6313), .A2(n6474), .B1(n6276), .B2(n6356), .ZN(n6277)
         );
  INV_X1 U7295 ( .A(n6277), .ZN(n6281) );
  AOI22_X1 U7296 ( .A1(INSTQUEUE_REG_11__7__SCAN_IN), .A2(n6279), .B1(n6466), 
        .B2(n6278), .ZN(n6280) );
  OAI211_X1 U7297 ( .C1(n6467), .C2(n6282), .A(n6281), .B(n6280), .ZN(U3115)
         );
  OAI22_X1 U7298 ( .A1(n6366), .A2(n6287), .B1(n6284), .B2(n6283), .ZN(n6309)
         );
  NOR3_X1 U7299 ( .A1(n6489), .A2(n6368), .A3(INSTQUEUEWR_ADDR_REG_1__SCAN_IN), 
        .ZN(n6320) );
  INV_X1 U7300 ( .A(n6320), .ZN(n6325) );
  NOR2_X1 U7301 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6325), .ZN(n6308)
         );
  AOI22_X1 U7302 ( .A1(n6412), .A2(n6309), .B1(n6411), .B2(n6308), .ZN(n6295)
         );
  AOI21_X1 U7303 ( .B1(n6313), .B2(n6357), .A(n6286), .ZN(n6293) );
  OAI21_X1 U7304 ( .B1(n6288), .B2(n6287), .A(n6419), .ZN(n6292) );
  INV_X1 U7305 ( .A(n6308), .ZN(n6289) );
  AOI21_X1 U7306 ( .B1(STATE2_REG_3__SCAN_IN), .B2(n6289), .A(n6367), .ZN(
        n6291) );
  AOI22_X1 U7307 ( .A1(INSTQUEUE_REG_12__0__SCAN_IN), .A2(n6310), .B1(n6376), 
        .B2(n6335), .ZN(n6294) );
  OAI211_X1 U7308 ( .C1(n6379), .C2(n6313), .A(n6295), .B(n6294), .ZN(U3116)
         );
  AOI22_X1 U7309 ( .A1(n6957), .A2(n6309), .B1(n6425), .B2(n6308), .ZN(n6297)
         );
  AOI22_X1 U7310 ( .A1(INSTQUEUE_REG_12__1__SCAN_IN), .A2(n6310), .B1(n6380), 
        .B2(n6335), .ZN(n6296) );
  OAI211_X1 U7311 ( .C1(n6953), .C2(n6313), .A(n6297), .B(n6296), .ZN(U3117)
         );
  AOI22_X1 U7312 ( .A1(n6430), .A2(n6309), .B1(n6429), .B2(n6308), .ZN(n6299)
         );
  AOI22_X1 U7313 ( .A1(INSTQUEUE_REG_12__2__SCAN_IN), .A2(n6310), .B1(n6383), 
        .B2(n6335), .ZN(n6298) );
  OAI211_X1 U7314 ( .C1(n6386), .C2(n6313), .A(n6299), .B(n6298), .ZN(U3118)
         );
  AOI22_X1 U7315 ( .A1(n6436), .A2(n6309), .B1(n6435), .B2(n6308), .ZN(n6301)
         );
  AOI22_X1 U7316 ( .A1(INSTQUEUE_REG_12__3__SCAN_IN), .A2(n6310), .B1(n6387), 
        .B2(n6335), .ZN(n6300) );
  OAI211_X1 U7317 ( .C1(n6437), .C2(n6313), .A(n6301), .B(n6300), .ZN(U3119)
         );
  AOI22_X1 U7318 ( .A1(n6443), .A2(n6309), .B1(n6442), .B2(n6308), .ZN(n6303)
         );
  AOI22_X1 U7319 ( .A1(INSTQUEUE_REG_12__4__SCAN_IN), .A2(n6310), .B1(n6390), 
        .B2(n6335), .ZN(n6302) );
  OAI211_X1 U7320 ( .C1(n6444), .C2(n6313), .A(n6303), .B(n6302), .ZN(U3120)
         );
  AOI22_X1 U7321 ( .A1(n6450), .A2(n6309), .B1(n6449), .B2(n6308), .ZN(n6305)
         );
  AOI22_X1 U7322 ( .A1(INSTQUEUE_REG_12__5__SCAN_IN), .A2(n6310), .B1(n6393), 
        .B2(n6335), .ZN(n6304) );
  OAI211_X1 U7323 ( .C1(n6451), .C2(n6313), .A(n6305), .B(n6304), .ZN(U3121)
         );
  AOI22_X1 U7324 ( .A1(n6457), .A2(n6309), .B1(n6456), .B2(n6308), .ZN(n6307)
         );
  AOI22_X1 U7325 ( .A1(INSTQUEUE_REG_12__6__SCAN_IN), .A2(n6310), .B1(n6396), 
        .B2(n6335), .ZN(n6306) );
  OAI211_X1 U7326 ( .C1(n6458), .C2(n6313), .A(n6307), .B(n6306), .ZN(U3122)
         );
  AOI22_X1 U7327 ( .A1(n6466), .A2(n6309), .B1(n6463), .B2(n6308), .ZN(n6312)
         );
  AOI22_X1 U7328 ( .A1(INSTQUEUE_REG_12__7__SCAN_IN), .A2(n6310), .B1(n6401), 
        .B2(n6335), .ZN(n6311) );
  OAI211_X1 U7329 ( .C1(n6467), .C2(n6313), .A(n6312), .B(n6311), .ZN(U3123)
         );
  INV_X1 U7330 ( .A(n6413), .ZN(n6315) );
  NOR2_X1 U7331 ( .A1(n6315), .A2(n6314), .ZN(n6327) );
  INV_X1 U7332 ( .A(n6327), .ZN(n6318) );
  NOR2_X1 U7333 ( .A1(n6316), .A2(n6325), .ZN(n6322) );
  AOI21_X1 U7334 ( .B1(n6408), .B2(n6317), .A(n6322), .ZN(n6326) );
  NAND2_X1 U7335 ( .A1(n6318), .A2(n6326), .ZN(n6319) );
  OAI211_X1 U7336 ( .C1(n6419), .C2(n6320), .A(n6319), .B(n6418), .ZN(n6360)
         );
  INV_X1 U7337 ( .A(n6360), .ZN(n6338) );
  INV_X1 U7338 ( .A(INSTQUEUE_REG_13__0__SCAN_IN), .ZN(n6706) );
  INV_X1 U7339 ( .A(n6322), .ZN(n6355) );
  OAI22_X1 U7340 ( .A1(n6405), .A2(n6424), .B1(n6323), .B2(n6355), .ZN(n6324)
         );
  INV_X1 U7341 ( .A(n6324), .ZN(n6329) );
  INV_X1 U7342 ( .A(n6379), .ZN(n6421) );
  OAI22_X1 U7343 ( .A1(n6327), .A2(n6326), .B1(n6511), .B2(n6325), .ZN(n6359)
         );
  AOI22_X1 U7344 ( .A1(n6421), .A2(n6335), .B1(n6412), .B2(n6359), .ZN(n6328)
         );
  OAI211_X1 U7345 ( .C1(n6338), .C2(n6706), .A(n6329), .B(n6328), .ZN(U3124)
         );
  OAI22_X1 U7346 ( .A1(n6357), .A2(n6953), .B1(n6951), .B2(n6355), .ZN(n6330)
         );
  INV_X1 U7347 ( .A(n6330), .ZN(n6332) );
  AOI22_X1 U7348 ( .A1(INSTQUEUE_REG_13__1__SCAN_IN), .A2(n6360), .B1(n6957), 
        .B2(n6359), .ZN(n6331) );
  OAI211_X1 U7349 ( .C1(n6962), .C2(n6405), .A(n6332), .B(n6331), .ZN(U3125)
         );
  INV_X1 U7350 ( .A(INSTQUEUE_REG_13__2__SCAN_IN), .ZN(n6769) );
  OAI22_X1 U7351 ( .A1(n6405), .A2(n6434), .B1(n6333), .B2(n6355), .ZN(n6334)
         );
  INV_X1 U7352 ( .A(n6334), .ZN(n6337) );
  INV_X1 U7353 ( .A(n6386), .ZN(n6431) );
  AOI22_X1 U7354 ( .A1(n6431), .A2(n6335), .B1(n6430), .B2(n6359), .ZN(n6336)
         );
  OAI211_X1 U7355 ( .C1(n6338), .C2(n6769), .A(n6337), .B(n6336), .ZN(U3126)
         );
  OAI22_X1 U7356 ( .A1(n6357), .A2(n6437), .B1(n6339), .B2(n6355), .ZN(n6340)
         );
  INV_X1 U7357 ( .A(n6340), .ZN(n6342) );
  AOI22_X1 U7358 ( .A1(INSTQUEUE_REG_13__3__SCAN_IN), .A2(n6360), .B1(n6436), 
        .B2(n6359), .ZN(n6341) );
  OAI211_X1 U7359 ( .C1(n6441), .C2(n6405), .A(n6342), .B(n6341), .ZN(U3127)
         );
  OAI22_X1 U7360 ( .A1(n6357), .A2(n6444), .B1(n6343), .B2(n6355), .ZN(n6344)
         );
  INV_X1 U7361 ( .A(n6344), .ZN(n6346) );
  AOI22_X1 U7362 ( .A1(INSTQUEUE_REG_13__4__SCAN_IN), .A2(n6360), .B1(n6443), 
        .B2(n6359), .ZN(n6345) );
  OAI211_X1 U7363 ( .C1(n6448), .C2(n6405), .A(n6346), .B(n6345), .ZN(U3128)
         );
  OAI22_X1 U7364 ( .A1(n6405), .A2(n6455), .B1(n6347), .B2(n6355), .ZN(n6348)
         );
  INV_X1 U7365 ( .A(n6348), .ZN(n6350) );
  AOI22_X1 U7366 ( .A1(INSTQUEUE_REG_13__5__SCAN_IN), .A2(n6360), .B1(n6450), 
        .B2(n6359), .ZN(n6349) );
  OAI211_X1 U7367 ( .C1(n6451), .C2(n6357), .A(n6350), .B(n6349), .ZN(U3129)
         );
  OAI22_X1 U7368 ( .A1(n6405), .A2(n6462), .B1(n6351), .B2(n6355), .ZN(n6352)
         );
  INV_X1 U7369 ( .A(n6352), .ZN(n6354) );
  AOI22_X1 U7370 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(n6360), .B1(n6457), 
        .B2(n6359), .ZN(n6353) );
  OAI211_X1 U7371 ( .C1(n6458), .C2(n6357), .A(n6354), .B(n6353), .ZN(U3130)
         );
  OAI22_X1 U7372 ( .A1(n6357), .A2(n6467), .B1(n6356), .B2(n6355), .ZN(n6358)
         );
  INV_X1 U7373 ( .A(n6358), .ZN(n6362) );
  AOI22_X1 U7374 ( .A1(INSTQUEUE_REG_13__7__SCAN_IN), .A2(n6360), .B1(n6466), 
        .B2(n6359), .ZN(n6361) );
  OAI211_X1 U7375 ( .C1(n6474), .C2(n6405), .A(n6362), .B(n6361), .ZN(U3131)
         );
  NAND3_X1 U7376 ( .A1(n6364), .A2(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), .A3(n6363), .ZN(n6365) );
  OAI21_X1 U7377 ( .B1(n6366), .B2(n6373), .A(n6365), .ZN(n6400) );
  INV_X1 U7378 ( .A(n6420), .ZN(n6409) );
  NOR2_X1 U7379 ( .A1(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A2(n6409), .ZN(n6399)
         );
  AOI22_X1 U7380 ( .A1(n6412), .A2(n6400), .B1(n6411), .B2(n6399), .ZN(n6378)
         );
  NOR3_X1 U7381 ( .A1(n6369), .A2(n6368), .A3(n6367), .ZN(n6375) );
  INV_X1 U7382 ( .A(n6405), .ZN(n6371) );
  OAI21_X1 U7383 ( .B1(n6371), .B2(n6468), .A(STATEBS16_REG_SCAN_IN), .ZN(
        n6372) );
  NAND3_X1 U7384 ( .A1(n6373), .A2(n6419), .A3(n6372), .ZN(n6374) );
  AOI22_X1 U7385 ( .A1(INSTQUEUE_REG_14__0__SCAN_IN), .A2(n6402), .B1(n6376), 
        .B2(n6468), .ZN(n6377) );
  OAI211_X1 U7386 ( .C1(n6379), .C2(n6405), .A(n6378), .B(n6377), .ZN(U3132)
         );
  AOI22_X1 U7387 ( .A1(n6957), .A2(n6400), .B1(n6425), .B2(n6399), .ZN(n6382)
         );
  AOI22_X1 U7388 ( .A1(INSTQUEUE_REG_14__1__SCAN_IN), .A2(n6402), .B1(n6380), 
        .B2(n6468), .ZN(n6381) );
  OAI211_X1 U7389 ( .C1(n6953), .C2(n6405), .A(n6382), .B(n6381), .ZN(U3133)
         );
  AOI22_X1 U7390 ( .A1(n6430), .A2(n6400), .B1(n6429), .B2(n6399), .ZN(n6385)
         );
  AOI22_X1 U7391 ( .A1(INSTQUEUE_REG_14__2__SCAN_IN), .A2(n6402), .B1(n6383), 
        .B2(n6468), .ZN(n6384) );
  OAI211_X1 U7392 ( .C1(n6386), .C2(n6405), .A(n6385), .B(n6384), .ZN(U3134)
         );
  AOI22_X1 U7393 ( .A1(n6436), .A2(n6400), .B1(n6435), .B2(n6399), .ZN(n6389)
         );
  AOI22_X1 U7394 ( .A1(INSTQUEUE_REG_14__3__SCAN_IN), .A2(n6402), .B1(n6387), 
        .B2(n6468), .ZN(n6388) );
  OAI211_X1 U7395 ( .C1(n6437), .C2(n6405), .A(n6389), .B(n6388), .ZN(U3135)
         );
  AOI22_X1 U7396 ( .A1(n6443), .A2(n6400), .B1(n6442), .B2(n6399), .ZN(n6392)
         );
  AOI22_X1 U7397 ( .A1(INSTQUEUE_REG_14__4__SCAN_IN), .A2(n6402), .B1(n6390), 
        .B2(n6468), .ZN(n6391) );
  OAI211_X1 U7398 ( .C1(n6444), .C2(n6405), .A(n6392), .B(n6391), .ZN(U3136)
         );
  AOI22_X1 U7399 ( .A1(n6450), .A2(n6400), .B1(n6449), .B2(n6399), .ZN(n6395)
         );
  AOI22_X1 U7400 ( .A1(INSTQUEUE_REG_14__5__SCAN_IN), .A2(n6402), .B1(n6393), 
        .B2(n6468), .ZN(n6394) );
  OAI211_X1 U7401 ( .C1(n6451), .C2(n6405), .A(n6395), .B(n6394), .ZN(U3137)
         );
  AOI22_X1 U7402 ( .A1(n6457), .A2(n6400), .B1(n6456), .B2(n6399), .ZN(n6398)
         );
  AOI22_X1 U7403 ( .A1(INSTQUEUE_REG_14__6__SCAN_IN), .A2(n6402), .B1(n6396), 
        .B2(n6468), .ZN(n6397) );
  OAI211_X1 U7404 ( .C1(n6458), .C2(n6405), .A(n6398), .B(n6397), .ZN(U3138)
         );
  AOI22_X1 U7405 ( .A1(n6466), .A2(n6400), .B1(n6463), .B2(n6399), .ZN(n6404)
         );
  AOI22_X1 U7406 ( .A1(INSTQUEUE_REG_14__7__SCAN_IN), .A2(n6402), .B1(n6401), 
        .B2(n6468), .ZN(n6403) );
  OAI211_X1 U7407 ( .C1(n6467), .C2(n6405), .A(n6404), .B(n6403), .ZN(U3139)
         );
  INV_X1 U7408 ( .A(n6406), .ZN(n6464) );
  AOI21_X1 U7409 ( .B1(n6408), .B2(n6407), .A(n6464), .ZN(n6414) );
  OAI22_X1 U7410 ( .A1(n6414), .A2(n6410), .B1(n6409), .B2(n6511), .ZN(n6465)
         );
  AOI22_X1 U7411 ( .A1(n6412), .A2(n6465), .B1(n6464), .B2(n6411), .ZN(n6423)
         );
  AOI21_X1 U7412 ( .B1(n6413), .B2(n4688), .A(n5911), .ZN(n6416) );
  OAI21_X1 U7413 ( .B1(n6416), .B2(n6415), .A(n6414), .ZN(n6417) );
  OAI211_X1 U7414 ( .C1(n6420), .C2(n6419), .A(n6418), .B(n6417), .ZN(n6470)
         );
  AOI22_X1 U7415 ( .A1(INSTQUEUE_REG_15__0__SCAN_IN), .A2(n6470), .B1(n6421), 
        .B2(n6468), .ZN(n6422) );
  OAI211_X1 U7416 ( .C1(n6424), .C2(n6473), .A(n6423), .B(n6422), .ZN(U3140)
         );
  AOI22_X1 U7417 ( .A1(n6957), .A2(n6465), .B1(n6464), .B2(n6425), .ZN(n6428)
         );
  INV_X1 U7418 ( .A(n6953), .ZN(n6426) );
  AOI22_X1 U7419 ( .A1(INSTQUEUE_REG_15__1__SCAN_IN), .A2(n6470), .B1(n6426), 
        .B2(n6468), .ZN(n6427) );
  OAI211_X1 U7420 ( .C1(n6962), .C2(n6473), .A(n6428), .B(n6427), .ZN(U3141)
         );
  AOI22_X1 U7421 ( .A1(n6430), .A2(n6465), .B1(n6464), .B2(n6429), .ZN(n6433)
         );
  AOI22_X1 U7422 ( .A1(INSTQUEUE_REG_15__2__SCAN_IN), .A2(n6470), .B1(n6431), 
        .B2(n6468), .ZN(n6432) );
  OAI211_X1 U7423 ( .C1(n6434), .C2(n6473), .A(n6433), .B(n6432), .ZN(U3142)
         );
  AOI22_X1 U7424 ( .A1(n6436), .A2(n6465), .B1(n6464), .B2(n6435), .ZN(n6440)
         );
  INV_X1 U7425 ( .A(n6437), .ZN(n6438) );
  AOI22_X1 U7426 ( .A1(INSTQUEUE_REG_15__3__SCAN_IN), .A2(n6470), .B1(n6438), 
        .B2(n6468), .ZN(n6439) );
  OAI211_X1 U7427 ( .C1(n6441), .C2(n6473), .A(n6440), .B(n6439), .ZN(U3143)
         );
  AOI22_X1 U7428 ( .A1(n6443), .A2(n6465), .B1(n6464), .B2(n6442), .ZN(n6447)
         );
  INV_X1 U7429 ( .A(n6444), .ZN(n6445) );
  AOI22_X1 U7430 ( .A1(INSTQUEUE_REG_15__4__SCAN_IN), .A2(n6470), .B1(n6445), 
        .B2(n6468), .ZN(n6446) );
  OAI211_X1 U7431 ( .C1(n6448), .C2(n6473), .A(n6447), .B(n6446), .ZN(U3144)
         );
  AOI22_X1 U7432 ( .A1(n6450), .A2(n6465), .B1(n6464), .B2(n6449), .ZN(n6454)
         );
  INV_X1 U7433 ( .A(n6451), .ZN(n6452) );
  AOI22_X1 U7434 ( .A1(INSTQUEUE_REG_15__5__SCAN_IN), .A2(n6470), .B1(n6452), 
        .B2(n6468), .ZN(n6453) );
  OAI211_X1 U7435 ( .C1(n6455), .C2(n6473), .A(n6454), .B(n6453), .ZN(U3145)
         );
  AOI22_X1 U7436 ( .A1(n6457), .A2(n6465), .B1(n6464), .B2(n6456), .ZN(n6461)
         );
  INV_X1 U7437 ( .A(n6458), .ZN(n6459) );
  AOI22_X1 U7438 ( .A1(INSTQUEUE_REG_15__6__SCAN_IN), .A2(n6470), .B1(n6459), 
        .B2(n6468), .ZN(n6460) );
  OAI211_X1 U7439 ( .C1(n6462), .C2(n6473), .A(n6461), .B(n6460), .ZN(U3146)
         );
  AOI22_X1 U7440 ( .A1(n6466), .A2(n6465), .B1(n6464), .B2(n6463), .ZN(n6472)
         );
  INV_X1 U7441 ( .A(n6467), .ZN(n6469) );
  AOI22_X1 U7442 ( .A1(INSTQUEUE_REG_15__7__SCAN_IN), .A2(n6470), .B1(n6469), 
        .B2(n6468), .ZN(n6471) );
  OAI211_X1 U7443 ( .C1(n6474), .C2(n6473), .A(n6472), .B(n6471), .ZN(U3147)
         );
  OAI22_X1 U7444 ( .A1(n6477), .A2(n6476), .B1(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .B2(n6475), .ZN(n6607) );
  INV_X1 U7445 ( .A(n6607), .ZN(n6479) );
  OR2_X1 U7446 ( .A1(n6478), .A2(n3711), .ZN(n6615) );
  NAND3_X1 U7447 ( .A1(n6479), .A2(INSTQUEUEWR_ADDR_REG_0__SCAN_IN), .A3(n6615), .ZN(n6482) );
  OAI211_X1 U7448 ( .C1(n6483), .C2(n6482), .A(n6481), .B(n6480), .ZN(n6485)
         );
  NAND2_X1 U7449 ( .A1(n6483), .A2(n6482), .ZN(n6484) );
  NAND2_X1 U7450 ( .A1(n6485), .A2(n6484), .ZN(n6490) );
  INV_X1 U7451 ( .A(n6490), .ZN(n6487) );
  OAI21_X1 U7452 ( .B1(INSTQUEUEWR_ADDR_REG_2__SCAN_IN), .B2(n6487), .A(n6486), 
        .ZN(n6488) );
  OAI21_X1 U7453 ( .B1(n6490), .B2(n6489), .A(n6488), .ZN(n6492) );
  INV_X1 U7454 ( .A(n6492), .ZN(n6495) );
  INV_X1 U7455 ( .A(n6494), .ZN(n6491) );
  AOI21_X1 U7456 ( .B1(n6492), .B2(n6491), .A(INSTQUEUEWR_ADDR_REG_3__SCAN_IN), 
        .ZN(n6493) );
  AOI21_X1 U7457 ( .B1(n6495), .B2(n6494), .A(n6493), .ZN(n6505) );
  INV_X1 U7458 ( .A(n6496), .ZN(n6501) );
  OAI21_X1 U7459 ( .B1(FLUSH_REG_SCAN_IN), .B2(MORE_REG_SCAN_IN), .A(n6497), 
        .ZN(n6498) );
  INV_X1 U7460 ( .A(n6498), .ZN(n6500) );
  NOR4_X1 U7461 ( .A1(n6502), .A2(n6501), .A3(n6500), .A4(n6499), .ZN(n6503)
         );
  OAI211_X1 U7462 ( .C1(n6505), .C2(INSTQUEUEWR_ADDR_REG_4__SCAN_IN), .A(n6504), .B(n6503), .ZN(n6517) );
  OR2_X1 U7463 ( .A1(n6507), .A2(n6506), .ZN(n6509) );
  INV_X1 U7464 ( .A(READY_N), .ZN(n6628) );
  OAI21_X1 U7465 ( .B1(n6522), .B2(n6628), .A(n6521), .ZN(n6508) );
  AND3_X1 U7466 ( .A1(n6509), .A2(STATE2_REG_2__SCAN_IN), .A3(n6508), .ZN(
        n6512) );
  INV_X1 U7467 ( .A(n6512), .ZN(n6510) );
  AOI221_X1 U7468 ( .B1(STATE2_REG_1__SCAN_IN), .B2(STATE2_REG_0__SCAN_IN), 
        .C1(n6517), .C2(STATE2_REG_0__SCAN_IN), .A(n6510), .ZN(n6595) );
  AOI21_X1 U7469 ( .B1(READY_N), .B2(n6511), .A(n6595), .ZN(n6523) );
  NOR2_X1 U7470 ( .A1(n6598), .A2(n6529), .ZN(n6514) );
  AOI211_X1 U7471 ( .C1(n6514), .C2(n6513), .A(STATE2_REG_0__SCAN_IN), .B(
        n6512), .ZN(n6515) );
  AOI211_X1 U7472 ( .C1(n6518), .C2(n6517), .A(n6516), .B(n6515), .ZN(n6519)
         );
  OAI221_X1 U7473 ( .B1(n6521), .B2(n6523), .C1(n6521), .C2(n6520), .A(n6519), 
        .ZN(U3148) );
  NOR2_X1 U7474 ( .A1(STATE2_REG_0__SCAN_IN), .A2(STATE2_REG_2__SCAN_IN), .ZN(
        n6532) );
  NOR3_X1 U7475 ( .A1(n6532), .A2(n6523), .A3(n6522), .ZN(n6527) );
  AOI221_X1 U7476 ( .B1(READY_N), .B2(n6525), .C1(n6524), .C2(n6525), .A(n6595), .ZN(n6526) );
  OR3_X1 U7477 ( .A1(n6528), .A2(n6527), .A3(n6526), .ZN(U3149) );
  OAI211_X1 U7478 ( .C1(STATE2_REG_2__SCAN_IN), .C2(n6628), .A(n6596), .B(
        n6529), .ZN(n6531) );
  OAI21_X1 U7479 ( .B1(n6532), .B2(n6531), .A(n6530), .ZN(U3150) );
  INV_X1 U7480 ( .A(DATAWIDTH_REG_31__SCAN_IN), .ZN(n6821) );
  NOR2_X1 U7481 ( .A1(n6594), .A2(n6821), .ZN(U3151) );
  AND2_X1 U7482 ( .A1(DATAWIDTH_REG_30__SCAN_IN), .A2(n6533), .ZN(U3152) );
  AND2_X1 U7483 ( .A1(DATAWIDTH_REG_29__SCAN_IN), .A2(n6533), .ZN(U3153) );
  AND2_X1 U7484 ( .A1(DATAWIDTH_REG_28__SCAN_IN), .A2(n6533), .ZN(U3154) );
  AND2_X1 U7485 ( .A1(DATAWIDTH_REG_27__SCAN_IN), .A2(n6533), .ZN(U3155) );
  AND2_X1 U7486 ( .A1(DATAWIDTH_REG_26__SCAN_IN), .A2(n6533), .ZN(U3156) );
  INV_X1 U7487 ( .A(DATAWIDTH_REG_25__SCAN_IN), .ZN(n6888) );
  NOR2_X1 U7488 ( .A1(n6594), .A2(n6888), .ZN(U3157) );
  NOR2_X1 U7489 ( .A1(n6594), .A2(n6702), .ZN(U3158) );
  AND2_X1 U7490 ( .A1(DATAWIDTH_REG_23__SCAN_IN), .A2(n6533), .ZN(U3159) );
  AND2_X1 U7491 ( .A1(DATAWIDTH_REG_22__SCAN_IN), .A2(n6533), .ZN(U3160) );
  AND2_X1 U7492 ( .A1(DATAWIDTH_REG_21__SCAN_IN), .A2(n6533), .ZN(U3161) );
  INV_X1 U7493 ( .A(DATAWIDTH_REG_20__SCAN_IN), .ZN(n6933) );
  NOR2_X1 U7494 ( .A1(n6594), .A2(n6933), .ZN(U3162) );
  INV_X1 U7495 ( .A(DATAWIDTH_REG_19__SCAN_IN), .ZN(n6847) );
  NOR2_X1 U7496 ( .A1(n6594), .A2(n6847), .ZN(U3163) );
  AND2_X1 U7497 ( .A1(DATAWIDTH_REG_18__SCAN_IN), .A2(n6533), .ZN(U3164) );
  AND2_X1 U7498 ( .A1(DATAWIDTH_REG_17__SCAN_IN), .A2(n6533), .ZN(U3165) );
  AND2_X1 U7499 ( .A1(DATAWIDTH_REG_16__SCAN_IN), .A2(n6533), .ZN(U3166) );
  NOR2_X1 U7500 ( .A1(n6594), .A2(n6813), .ZN(U3167) );
  NOR2_X1 U7501 ( .A1(n6594), .A2(n6782), .ZN(U3168) );
  NOR2_X1 U7502 ( .A1(n6594), .A2(n6772), .ZN(U3169) );
  NOR2_X1 U7503 ( .A1(n6594), .A2(n6781), .ZN(U3170) );
  AND2_X1 U7504 ( .A1(DATAWIDTH_REG_11__SCAN_IN), .A2(n6533), .ZN(U3171) );
  INV_X1 U7505 ( .A(DATAWIDTH_REG_10__SCAN_IN), .ZN(n6718) );
  NOR2_X1 U7506 ( .A1(n6594), .A2(n6718), .ZN(U3172) );
  AND2_X1 U7507 ( .A1(DATAWIDTH_REG_9__SCAN_IN), .A2(n6533), .ZN(U3173) );
  AND2_X1 U7508 ( .A1(DATAWIDTH_REG_8__SCAN_IN), .A2(n6533), .ZN(U3174) );
  AND2_X1 U7509 ( .A1(DATAWIDTH_REG_7__SCAN_IN), .A2(n6533), .ZN(U3175) );
  AND2_X1 U7510 ( .A1(DATAWIDTH_REG_6__SCAN_IN), .A2(n6533), .ZN(U3176) );
  INV_X1 U7511 ( .A(DATAWIDTH_REG_5__SCAN_IN), .ZN(n6831) );
  NOR2_X1 U7512 ( .A1(n6594), .A2(n6831), .ZN(U3177) );
  AND2_X1 U7513 ( .A1(DATAWIDTH_REG_4__SCAN_IN), .A2(n6533), .ZN(U3178) );
  INV_X1 U7514 ( .A(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6760) );
  NOR2_X1 U7515 ( .A1(n6594), .A2(n6760), .ZN(U3179) );
  INV_X1 U7516 ( .A(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6926) );
  NOR2_X1 U7517 ( .A1(n6594), .A2(n6926), .ZN(U3180) );
  INV_X1 U7518 ( .A(STATE_REG_1__SCAN_IN), .ZN(n6540) );
  NOR2_X1 U7519 ( .A1(n6550), .A2(n6540), .ZN(n6543) );
  AOI22_X1 U7520 ( .A1(READY_N), .A2(STATE_REG_1__SCAN_IN), .B1(
        STATE_REG_2__SCAN_IN), .B2(HOLD), .ZN(n6547) );
  AND2_X1 U7521 ( .A1(STATE_REG_1__SCAN_IN), .A2(HOLD), .ZN(n6537) );
  INV_X1 U7522 ( .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6535) );
  INV_X1 U7523 ( .A(NA_N), .ZN(n6544) );
  AOI211_X1 U7524 ( .C1(STATE_REG_2__SCAN_IN), .C2(n6544), .A(
        STATE_REG_0__SCAN_IN), .B(n6543), .ZN(n6549) );
  AOI221_X1 U7525 ( .B1(n6537), .B2(n6636), .C1(n6535), .C2(n6636), .A(n6549), 
        .ZN(n6534) );
  OAI21_X1 U7526 ( .B1(n6543), .B2(n6547), .A(n6534), .ZN(U3181) );
  NOR2_X1 U7527 ( .A1(n6541), .A2(n6535), .ZN(n6545) );
  NAND2_X1 U7528 ( .A1(STATE_REG_2__SCAN_IN), .A2(HOLD), .ZN(n6536) );
  OAI21_X1 U7529 ( .B1(n6545), .B2(n6537), .A(n6536), .ZN(n6538) );
  OAI211_X1 U7530 ( .C1(n6540), .C2(n6628), .A(n6539), .B(n6538), .ZN(U3182)
         );
  AOI221_X1 U7531 ( .B1(NA_N), .B2(STATE_REG_1__SCAN_IN), .C1(n6628), .C2(
        STATE_REG_1__SCAN_IN), .A(REQUESTPENDING_REG_SCAN_IN), .ZN(n6542) );
  AOI221_X1 U7532 ( .B1(STATE_REG_2__SCAN_IN), .B2(HOLD), .C1(n6542), .C2(HOLD), .A(n6541), .ZN(n6548) );
  AOI21_X1 U7533 ( .B1(n6545), .B2(n6544), .A(n6543), .ZN(n6546) );
  OAI22_X1 U7534 ( .A1(n6549), .A2(n6548), .B1(n6547), .B2(n6546), .ZN(U3183)
         );
  NOR2_X1 U7535 ( .A1(n6550), .A2(n6636), .ZN(n6587) );
  NAND2_X1 U7536 ( .A1(n6550), .A2(n6625), .ZN(n6589) );
  AOI22_X1 U7537 ( .A1(REIP_REG_2__SCAN_IN), .A2(n6574), .B1(
        ADDRESS_REG_0__SCAN_IN), .B2(n6636), .ZN(n6551) );
  OAI21_X1 U7538 ( .B1(n6616), .B2(n6586), .A(n6551), .ZN(U3184) );
  AOI22_X1 U7539 ( .A1(REIP_REG_3__SCAN_IN), .A2(n6574), .B1(
        ADDRESS_REG_1__SCAN_IN), .B2(n6636), .ZN(n6552) );
  OAI21_X1 U7540 ( .B1(n4823), .B2(n6586), .A(n6552), .ZN(U3185) );
  INV_X1 U7541 ( .A(ADDRESS_REG_2__SCAN_IN), .ZN(n6910) );
  OAI222_X1 U7542 ( .A1(n6586), .A2(n6553), .B1(n6910), .B2(n6625), .C1(n6929), 
        .C2(n6589), .ZN(U3186) );
  AOI22_X1 U7543 ( .A1(REIP_REG_5__SCAN_IN), .A2(n6574), .B1(
        ADDRESS_REG_3__SCAN_IN), .B2(n6636), .ZN(n6554) );
  OAI21_X1 U7544 ( .B1(n6929), .B2(n6586), .A(n6554), .ZN(U3187) );
  AOI22_X1 U7545 ( .A1(REIP_REG_6__SCAN_IN), .A2(n6574), .B1(
        ADDRESS_REG_4__SCAN_IN), .B2(n6636), .ZN(n6555) );
  OAI21_X1 U7546 ( .B1(n5637), .B2(n6586), .A(n6555), .ZN(U3188) );
  AOI22_X1 U7547 ( .A1(REIP_REG_7__SCAN_IN), .A2(n6574), .B1(
        ADDRESS_REG_5__SCAN_IN), .B2(n6636), .ZN(n6556) );
  OAI21_X1 U7548 ( .B1(n6557), .B2(n6586), .A(n6556), .ZN(U3189) );
  INV_X1 U7549 ( .A(ADDRESS_REG_6__SCAN_IN), .ZN(n6719) );
  OAI222_X1 U7550 ( .A1(n6586), .A2(n6558), .B1(n6719), .B2(n6625), .C1(n6767), 
        .C2(n6589), .ZN(U3190) );
  INV_X1 U7551 ( .A(ADDRESS_REG_7__SCAN_IN), .ZN(n6936) );
  OAI222_X1 U7552 ( .A1(n6589), .A2(n4806), .B1(n6936), .B2(n6625), .C1(n6767), 
        .C2(n6586), .ZN(U3191) );
  INV_X1 U7553 ( .A(ADDRESS_REG_8__SCAN_IN), .ZN(n6861) );
  OAI222_X1 U7554 ( .A1(n6589), .A2(n4849), .B1(n6861), .B2(n6625), .C1(n4806), 
        .C2(n6586), .ZN(U3192) );
  INV_X1 U7555 ( .A(ADDRESS_REG_9__SCAN_IN), .ZN(n6700) );
  OAI222_X1 U7556 ( .A1(n6586), .A2(n4849), .B1(n6700), .B2(n6625), .C1(n4884), 
        .C2(n6589), .ZN(U3193) );
  INV_X1 U7557 ( .A(ADDRESS_REG_10__SCAN_IN), .ZN(n6853) );
  OAI222_X1 U7558 ( .A1(n6589), .A2(n6560), .B1(n6853), .B2(n6625), .C1(n4884), 
        .C2(n6586), .ZN(U3194) );
  AOI22_X1 U7559 ( .A1(REIP_REG_13__SCAN_IN), .A2(n6574), .B1(
        ADDRESS_REG_11__SCAN_IN), .B2(n6636), .ZN(n6559) );
  OAI21_X1 U7560 ( .B1(n6560), .B2(n6586), .A(n6559), .ZN(U3195) );
  AOI22_X1 U7561 ( .A1(REIP_REG_14__SCAN_IN), .A2(n6574), .B1(
        ADDRESS_REG_12__SCAN_IN), .B2(n6636), .ZN(n6561) );
  OAI21_X1 U7562 ( .B1(n6562), .B2(n6586), .A(n6561), .ZN(U3196) );
  INV_X1 U7563 ( .A(ADDRESS_REG_13__SCAN_IN), .ZN(n6927) );
  OAI222_X1 U7564 ( .A1(n6589), .A2(n6565), .B1(n6927), .B2(n6625), .C1(n6563), 
        .C2(n6586), .ZN(U3197) );
  AOI22_X1 U7565 ( .A1(REIP_REG_16__SCAN_IN), .A2(n6574), .B1(
        ADDRESS_REG_14__SCAN_IN), .B2(n6636), .ZN(n6564) );
  OAI21_X1 U7566 ( .B1(n6565), .B2(n6586), .A(n6564), .ZN(U3198) );
  AOI22_X1 U7567 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6574), .B1(
        ADDRESS_REG_15__SCAN_IN), .B2(n6636), .ZN(n6566) );
  OAI21_X1 U7568 ( .B1(n6869), .B2(n6586), .A(n6566), .ZN(U3199) );
  AOI22_X1 U7569 ( .A1(REIP_REG_17__SCAN_IN), .A2(n6587), .B1(
        ADDRESS_REG_16__SCAN_IN), .B2(n6636), .ZN(n6567) );
  OAI21_X1 U7570 ( .B1(n6569), .B2(n6589), .A(n6567), .ZN(U3200) );
  AOI22_X1 U7571 ( .A1(REIP_REG_19__SCAN_IN), .A2(n6574), .B1(
        ADDRESS_REG_17__SCAN_IN), .B2(n6636), .ZN(n6568) );
  OAI21_X1 U7572 ( .B1(n6569), .B2(n6586), .A(n6568), .ZN(U3201) );
  AOI22_X1 U7573 ( .A1(REIP_REG_20__SCAN_IN), .A2(n6574), .B1(
        ADDRESS_REG_18__SCAN_IN), .B2(n6636), .ZN(n6570) );
  OAI21_X1 U7574 ( .B1(n6738), .B2(n6586), .A(n6570), .ZN(U3202) );
  AOI22_X1 U7575 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6574), .B1(
        ADDRESS_REG_19__SCAN_IN), .B2(n6636), .ZN(n6571) );
  OAI21_X1 U7576 ( .B1(n6572), .B2(n6586), .A(n6571), .ZN(U3203) );
  AOI22_X1 U7577 ( .A1(REIP_REG_21__SCAN_IN), .A2(n6587), .B1(
        ADDRESS_REG_20__SCAN_IN), .B2(n6636), .ZN(n6573) );
  OAI21_X1 U7578 ( .B1(n6576), .B2(n6589), .A(n6573), .ZN(U3204) );
  AOI22_X1 U7579 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6574), .B1(
        ADDRESS_REG_21__SCAN_IN), .B2(n6636), .ZN(n6575) );
  OAI21_X1 U7580 ( .B1(n6576), .B2(n6586), .A(n6575), .ZN(U3205) );
  AOI22_X1 U7581 ( .A1(REIP_REG_23__SCAN_IN), .A2(n6587), .B1(
        ADDRESS_REG_22__SCAN_IN), .B2(n6636), .ZN(n6577) );
  OAI21_X1 U7582 ( .B1(n6578), .B2(n6589), .A(n6577), .ZN(U3206) );
  INV_X1 U7583 ( .A(REIP_REG_25__SCAN_IN), .ZN(n6832) );
  INV_X1 U7584 ( .A(ADDRESS_REG_23__SCAN_IN), .ZN(n6709) );
  OAI222_X1 U7585 ( .A1(n6589), .A2(n6832), .B1(n6709), .B2(n6625), .C1(n6578), 
        .C2(n6586), .ZN(U3207) );
  INV_X1 U7586 ( .A(ADDRESS_REG_24__SCAN_IN), .ZN(n6735) );
  INV_X1 U7587 ( .A(REIP_REG_26__SCAN_IN), .ZN(n6725) );
  OAI222_X1 U7588 ( .A1(n6586), .A2(n6832), .B1(n6735), .B2(n6625), .C1(n6725), 
        .C2(n6589), .ZN(U3208) );
  AOI22_X1 U7589 ( .A1(REIP_REG_26__SCAN_IN), .A2(n6587), .B1(
        ADDRESS_REG_25__SCAN_IN), .B2(n6636), .ZN(n6579) );
  OAI21_X1 U7590 ( .B1(n6580), .B2(n6589), .A(n6579), .ZN(U3209) );
  AOI22_X1 U7591 ( .A1(REIP_REG_27__SCAN_IN), .A2(n6587), .B1(
        ADDRESS_REG_26__SCAN_IN), .B2(n6636), .ZN(n6581) );
  OAI21_X1 U7592 ( .B1(n6582), .B2(n6589), .A(n6581), .ZN(U3210) );
  AOI22_X1 U7593 ( .A1(REIP_REG_28__SCAN_IN), .A2(n6587), .B1(
        ADDRESS_REG_27__SCAN_IN), .B2(n6636), .ZN(n6583) );
  OAI21_X1 U7594 ( .B1(n6585), .B2(n6589), .A(n6583), .ZN(U3211) );
  INV_X1 U7595 ( .A(ADDRESS_REG_28__SCAN_IN), .ZN(n6784) );
  OAI222_X1 U7596 ( .A1(n6586), .A2(n6585), .B1(n6784), .B2(n6625), .C1(n6584), 
        .C2(n6589), .ZN(U3212) );
  INV_X1 U7597 ( .A(REIP_REG_31__SCAN_IN), .ZN(n6590) );
  AOI22_X1 U7598 ( .A1(REIP_REG_30__SCAN_IN), .A2(n6587), .B1(
        ADDRESS_REG_29__SCAN_IN), .B2(n6636), .ZN(n6588) );
  OAI21_X1 U7599 ( .B1(n6590), .B2(n6589), .A(n6588), .ZN(U3213) );
  MUX2_X1 U7600 ( .A(BYTEENABLE_REG_3__SCAN_IN), .B(BE_N_REG_3__SCAN_IN), .S(
        n6636), .Z(U3445) );
  MUX2_X1 U7601 ( .A(BYTEENABLE_REG_2__SCAN_IN), .B(BE_N_REG_2__SCAN_IN), .S(
        n6636), .Z(U3446) );
  MUX2_X1 U7602 ( .A(BYTEENABLE_REG_1__SCAN_IN), .B(BE_N_REG_1__SCAN_IN), .S(
        n6636), .Z(U3447) );
  MUX2_X1 U7603 ( .A(BYTEENABLE_REG_0__SCAN_IN), .B(BE_N_REG_0__SCAN_IN), .S(
        n6636), .Z(U3448) );
  OAI21_X1 U7604 ( .B1(DATAWIDTH_REG_0__SCAN_IN), .B2(n6594), .A(n6592), .ZN(
        n6591) );
  INV_X1 U7605 ( .A(n6591), .ZN(U3451) );
  OAI21_X1 U7606 ( .B1(n6594), .B2(n6593), .A(n6592), .ZN(U3452) );
  INV_X1 U7607 ( .A(n6595), .ZN(n6599) );
  OAI211_X1 U7608 ( .C1(n6599), .C2(n6598), .A(n6597), .B(n6596), .ZN(U3453)
         );
  INV_X1 U7609 ( .A(n6600), .ZN(n6603) );
  OAI22_X1 U7610 ( .A1(n6603), .A2(n6614), .B1(n6602), .B2(n6601), .ZN(n6604)
         );
  MUX2_X1 U7611 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(n6604), .S(n6612), 
        .Z(U3456) );
  AOI22_X1 U7612 ( .A1(n6607), .A2(n6606), .B1(STATE2_REG_1__SCAN_IN), .B2(
        n6605), .ZN(n6610) );
  INV_X1 U7613 ( .A(n6608), .ZN(n6609) );
  NAND3_X1 U7614 ( .A1(n6612), .A2(n6610), .A3(n6609), .ZN(n6611) );
  OAI21_X1 U7615 ( .B1(n6612), .B2(INSTQUEUERD_ADDR_REG_0__SCAN_IN), .A(n6611), 
        .ZN(n6613) );
  OAI21_X1 U7616 ( .B1(n6615), .B2(n6614), .A(n6613), .ZN(U3461) );
  AOI21_X1 U7617 ( .B1(REIP_REG_0__SCAN_IN), .B2(DATAWIDTH_REG_0__SCAN_IN), 
        .A(DATAWIDTH_REG_1__SCAN_IN), .ZN(n6617) );
  AOI22_X1 U7618 ( .A1(REIP_REG_1__SCAN_IN), .A2(REIP_REG_0__SCAN_IN), .B1(
        n6617), .B2(n6616), .ZN(n6619) );
  INV_X1 U7619 ( .A(BYTEENABLE_REG_2__SCAN_IN), .ZN(n6618) );
  AOI22_X1 U7620 ( .A1(n6620), .A2(n6619), .B1(n6618), .B2(n6623), .ZN(U3468)
         );
  INV_X1 U7621 ( .A(BYTEENABLE_REG_0__SCAN_IN), .ZN(n6624) );
  NOR2_X1 U7622 ( .A1(n6623), .A2(REIP_REG_1__SCAN_IN), .ZN(n6621) );
  AOI22_X1 U7623 ( .A1(n6624), .A2(n6623), .B1(n6622), .B2(n6621), .ZN(U3469)
         );
  INV_X1 U7624 ( .A(W_R_N_REG_SCAN_IN), .ZN(n6932) );
  AOI22_X1 U7625 ( .A1(n6625), .A2(READREQUEST_REG_SCAN_IN), .B1(n6932), .B2(
        n6636), .ZN(U3470) );
  AOI211_X1 U7626 ( .C1(n5738), .C2(n6628), .A(n6627), .B(n6626), .ZN(n6635)
         );
  OAI211_X1 U7627 ( .C1(STATEBS16_REG_SCAN_IN), .C2(n6630), .A(n6629), .B(
        STATE2_REG_2__SCAN_IN), .ZN(n6632) );
  AOI21_X1 U7628 ( .B1(n6632), .B2(STATE2_REG_0__SCAN_IN), .A(n6631), .ZN(
        n6634) );
  NAND2_X1 U7629 ( .A1(n6635), .A2(REQUESTPENDING_REG_SCAN_IN), .ZN(n6633) );
  OAI21_X1 U7630 ( .B1(n6635), .B2(n6634), .A(n6633), .ZN(U3472) );
  MUX2_X1 U7631 ( .A(MEMORYFETCH_REG_SCAN_IN), .B(M_IO_N_REG_SCAN_IN), .S(
        n6636), .Z(U3473) );
  NOR4_X1 U7632 ( .A1(DATAO_REG_8__SCAN_IN), .A2(DATAO_REG_11__SCAN_IN), .A3(
        DATAO_REG_17__SCAN_IN), .A4(DATAO_REG_18__SCAN_IN), .ZN(n6640) );
  NOR4_X1 U7633 ( .A1(ADDRESS_REG_9__SCAN_IN), .A2(ADDRESS_REG_8__SCAN_IN), 
        .A3(DATAWIDTH_REG_15__SCAN_IN), .A4(DATAWIDTH_REG_25__SCAN_IN), .ZN(
        n6639) );
  NOR4_X1 U7634 ( .A1(EAX_REG_9__SCAN_IN), .A2(EAX_REG_11__SCAN_IN), .A3(
        LWORD_REG_11__SCAN_IN), .A4(LWORD_REG_0__SCAN_IN), .ZN(n6638) );
  NOR4_X1 U7635 ( .A1(PHYADDRPOINTER_REG_4__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_0__SCAN_IN), .A3(DATAO_REG_28__SCAN_IN), .A4(
        DATAWIDTH_REG_0__SCAN_IN), .ZN(n6637) );
  NAND4_X1 U7636 ( .A1(n6640), .A2(n6639), .A3(n6638), .A4(n6637), .ZN(n6681)
         );
  NOR4_X1 U7637 ( .A1(INSTQUEUE_REG_4__1__SCAN_IN), .A2(
        INSTQUEUE_REG_9__1__SCAN_IN), .A3(INSTQUEUE_REG_3__1__SCAN_IN), .A4(
        INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n6644) );
  INV_X1 U7638 ( .A(INSTQUEUE_REG_6__5__SCAN_IN), .ZN(n6865) );
  INV_X1 U7639 ( .A(INSTQUEUE_REG_15__5__SCAN_IN), .ZN(n6797) );
  NOR4_X1 U7640 ( .A1(INSTQUEUE_REG_1__5__SCAN_IN), .A2(
        INSTQUEUE_REG_12__5__SCAN_IN), .A3(n6865), .A4(n6797), .ZN(n6643) );
  NOR4_X1 U7641 ( .A1(W_R_N_REG_SCAN_IN), .A2(ADDRESS_REG_24__SCAN_IN), .A3(
        ADDRESS_REG_23__SCAN_IN), .A4(ADDRESS_REG_13__SCAN_IN), .ZN(n6642) );
  INV_X1 U7642 ( .A(INSTQUEUE_REG_7__1__SCAN_IN), .ZN(n6686) );
  NOR4_X1 U7643 ( .A1(DATAO_REG_4__SCAN_IN), .A2(ADDRESS_REG_6__SCAN_IN), .A3(
        D_C_N_REG_SCAN_IN), .A4(n6686), .ZN(n6641) );
  NAND4_X1 U7644 ( .A1(n6644), .A2(n6643), .A3(n6642), .A4(n6641), .ZN(n6680)
         );
  NAND4_X1 U7645 ( .A1(PHYADDRPOINTER_REG_18__SCAN_IN), .A2(
        DATAO_REG_30__SCAN_IN), .A3(n6708), .A4(n5897), .ZN(n6645) );
  NOR3_X1 U7646 ( .A1(EAX_REG_31__SCAN_IN), .A2(DATAI_20_), .A3(n6645), .ZN(
        n6654) );
  NAND4_X1 U7647 ( .A1(INSTADDRPOINTER_REG_9__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_13__SCAN_IN), .A3(EBX_REG_31__SCAN_IN), .A4(
        DATAI_7_), .ZN(n6652) );
  NAND4_X1 U7648 ( .A1(EBX_REG_21__SCAN_IN), .A2(PHYADDRPOINTER_REG_8__SCAN_IN), .A3(DATAWIDTH_REG_10__SCAN_IN), .A4(DATAO_REG_9__SCAN_IN), .ZN(n6651) );
  NOR4_X1 U7649 ( .A1(REIP_REG_8__SCAN_IN), .A2(REIP_REG_5__SCAN_IN), .A3(
        REIP_REG_9__SCAN_IN), .A4(REIP_REG_10__SCAN_IN), .ZN(n6649) );
  NOR4_X1 U7650 ( .A1(EAX_REG_17__SCAN_IN), .A2(REIP_REG_2__SCAN_IN), .A3(
        UWORD_REG_13__SCAN_IN), .A4(UWORD_REG_10__SCAN_IN), .ZN(n6648) );
  NOR4_X1 U7651 ( .A1(PHYADDRPOINTER_REG_20__SCAN_IN), .A2(EAX_REG_27__SCAN_IN), .A3(DATAI_12_), .A4(DATAI_5_), .ZN(n6647) );
  NOR4_X1 U7652 ( .A1(INSTADDRPOINTER_REG_27__SCAN_IN), .A2(
        EBX_REG_14__SCAN_IN), .A3(REIP_REG_16__SCAN_IN), .A4(
        CODEFETCH_REG_SCAN_IN), .ZN(n6646) );
  NAND4_X1 U7653 ( .A1(n6649), .A2(n6648), .A3(n6647), .A4(n6646), .ZN(n6650)
         );
  NOR3_X1 U7654 ( .A1(n6652), .A2(n6651), .A3(n6650), .ZN(n6653) );
  NAND4_X1 U7655 ( .A1(n6654), .A2(n6653), .A3(n6935), .A4(n6738), .ZN(n6679)
         );
  INV_X1 U7656 ( .A(INSTQUEUE_REG_15__2__SCAN_IN), .ZN(n6894) );
  NOR4_X1 U7657 ( .A1(INSTQUEUE_REG_7__7__SCAN_IN), .A2(
        INSTQUEUE_REG_5__7__SCAN_IN), .A3(INSTQUEUE_REG_1__2__SCAN_IN), .A4(
        n6894), .ZN(n6658) );
  INV_X1 U7658 ( .A(INSTQUEUE_REG_10__0__SCAN_IN), .ZN(n6895) );
  INV_X1 U7659 ( .A(INSTQUEUE_REG_2__0__SCAN_IN), .ZN(n6687) );
  INV_X1 U7660 ( .A(INSTQUEUE_REG_11__7__SCAN_IN), .ZN(n6803) );
  INV_X1 U7661 ( .A(INSTQUEUE_REG_14__7__SCAN_IN), .ZN(n6693) );
  NOR4_X1 U7662 ( .A1(n6895), .A2(n6687), .A3(n6803), .A4(n6693), .ZN(n6657)
         );
  INV_X1 U7663 ( .A(INSTQUEUE_REG_0__5__SCAN_IN), .ZN(n6699) );
  INV_X1 U7664 ( .A(INSTQUEUE_REG_4__6__SCAN_IN), .ZN(n6756) );
  NOR4_X1 U7665 ( .A1(INSTQUEUE_REG_14__5__SCAN_IN), .A2(
        INSTQUEUE_REG_7__6__SCAN_IN), .A3(n6699), .A4(n6756), .ZN(n6656) );
  NOR4_X1 U7666 ( .A1(INSTQUEUE_REG_13__6__SCAN_IN), .A2(
        INSTQUEUE_REG_5__2__SCAN_IN), .A3(n6866), .A4(n6769), .ZN(n6655) );
  NAND4_X1 U7667 ( .A1(n6658), .A2(n6657), .A3(n6656), .A4(n6655), .ZN(n6663)
         );
  INV_X1 U7668 ( .A(n6659), .ZN(n6660) );
  NOR4_X1 U7669 ( .A1(n6663), .A2(n6662), .A3(n6661), .A4(n6660), .ZN(n6677)
         );
  INV_X1 U7670 ( .A(INSTQUEUE_REG_8__0__SCAN_IN), .ZN(n6911) );
  NAND4_X1 U7671 ( .A1(INSTQUEUE_REG_1__4__SCAN_IN), .A2(
        INSTQUEUE_REG_6__0__SCAN_IN), .A3(n6911), .A4(n6706), .ZN(n6664) );
  NOR4_X1 U7672 ( .A1(REIP_REG_25__SCAN_IN), .A2(REIP_REG_26__SCAN_IN), .A3(
        n6665), .A4(n6664), .ZN(n6676) );
  NAND4_X1 U7673 ( .A1(EBX_REG_28__SCAN_IN), .A2(REIP_REG_4__SCAN_IN), .A3(
        DATAWIDTH_REG_20__SCAN_IN), .A4(ADDRESS_REG_7__SCAN_IN), .ZN(n6669) );
  NAND4_X1 U7674 ( .A1(EBX_REG_26__SCAN_IN), .A2(EBX_REG_3__SCAN_IN), .A3(
        INSTADDRPOINTER_REG_4__SCAN_IN), .A4(EAX_REG_23__SCAN_IN), .ZN(n6668)
         );
  NAND4_X1 U7675 ( .A1(UWORD_REG_5__SCAN_IN), .A2(DATAO_REG_3__SCAN_IN), .A3(
        DATAO_REG_0__SCAN_IN), .A4(DATAWIDTH_REG_2__SCAN_IN), .ZN(n6667) );
  NAND4_X1 U7676 ( .A1(PHYADDRPOINTER_REG_24__SCAN_IN), .A2(
        PHYADDRPOINTER_REG_14__SCAN_IN), .A3(LWORD_REG_7__SCAN_IN), .A4(
        ADDRESS_REG_2__SCAN_IN), .ZN(n6666) );
  NOR4_X1 U7677 ( .A1(n6669), .A2(n6668), .A3(n6667), .A4(n6666), .ZN(n6675)
         );
  NAND4_X1 U7678 ( .A1(ADDRESS_REG_28__SCAN_IN), .A2(UWORD_REG_3__SCAN_IN), 
        .A3(UWORD_REG_0__SCAN_IN), .A4(DATAWIDTH_REG_31__SCAN_IN), .ZN(n6673)
         );
  NAND4_X1 U7679 ( .A1(EBX_REG_27__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_8__SCAN_IN), .A3(PHYADDRPOINTER_REG_3__SCAN_IN), 
        .A4(DATAWIDTH_REG_3__SCAN_IN), .ZN(n6672) );
  NAND4_X1 U7680 ( .A1(EBX_REG_15__SCAN_IN), .A2(
        INSTADDRPOINTER_REG_19__SCAN_IN), .A3(DATAWIDTH_REG_19__SCAN_IN), .A4(
        ADDRESS_REG_10__SCAN_IN), .ZN(n6671) );
  NAND4_X1 U7681 ( .A1(EAX_REG_3__SCAN_IN), .A2(DATAI_14_), .A3(
        DATAWIDTH_REG_5__SCAN_IN), .A4(DATAO_REG_10__SCAN_IN), .ZN(n6670) );
  NOR4_X1 U7682 ( .A1(n6673), .A2(n6672), .A3(n6671), .A4(n6670), .ZN(n6674)
         );
  NAND4_X1 U7683 ( .A1(n6677), .A2(n6676), .A3(n6675), .A4(n6674), .ZN(n6678)
         );
  NOR4_X1 U7684 ( .A1(n6681), .A2(n6680), .A3(n6679), .A4(n6678), .ZN(n6950)
         );
  INV_X1 U7685 ( .A(INSTADDRPOINTER_REG_27__SCAN_IN), .ZN(n6683) );
  AOI22_X1 U7686 ( .A1(n6684), .A2(keyinput117), .B1(n6683), .B2(keyinput31), 
        .ZN(n6682) );
  OAI221_X1 U7687 ( .B1(n6684), .B2(keyinput117), .C1(n6683), .C2(keyinput31), 
        .A(n6682), .ZN(n6697) );
  AOI22_X1 U7688 ( .A1(n6687), .A2(keyinput29), .B1(keyinput102), .B2(n6686), 
        .ZN(n6685) );
  OAI221_X1 U7689 ( .B1(n6687), .B2(keyinput29), .C1(n6686), .C2(keyinput102), 
        .A(n6685), .ZN(n6696) );
  INV_X1 U7690 ( .A(INSTQUEUE_REG_15__1__SCAN_IN), .ZN(n6689) );
  AOI22_X1 U7691 ( .A1(n6690), .A2(keyinput77), .B1(n6689), .B2(keyinput60), 
        .ZN(n6688) );
  OAI221_X1 U7692 ( .B1(n6690), .B2(keyinput77), .C1(n6689), .C2(keyinput60), 
        .A(n6688), .ZN(n6695) );
  AOI22_X1 U7693 ( .A1(n6693), .A2(keyinput65), .B1(keyinput87), .B2(n6692), 
        .ZN(n6691) );
  OAI221_X1 U7694 ( .B1(n6693), .B2(keyinput65), .C1(n6692), .C2(keyinput87), 
        .A(n6691), .ZN(n6694) );
  NOR4_X1 U7695 ( .A1(n6697), .A2(n6696), .A3(n6695), .A4(n6694), .ZN(n6748)
         );
  AOI22_X1 U7696 ( .A1(n6700), .A2(keyinput92), .B1(n6699), .B2(keyinput51), 
        .ZN(n6698) );
  OAI221_X1 U7697 ( .B1(n6700), .B2(keyinput92), .C1(n6699), .C2(keyinput51), 
        .A(n6698), .ZN(n6713) );
  AOI22_X1 U7698 ( .A1(n6703), .A2(keyinput126), .B1(n6702), .B2(keyinput122), 
        .ZN(n6701) );
  OAI221_X1 U7699 ( .B1(n6703), .B2(keyinput126), .C1(n6702), .C2(keyinput122), 
        .A(n6701), .ZN(n6712) );
  AOI22_X1 U7700 ( .A1(n6709), .A2(keyinput121), .B1(n6708), .B2(keyinput109), 
        .ZN(n6707) );
  OAI221_X1 U7701 ( .B1(n6709), .B2(keyinput121), .C1(n6708), .C2(keyinput109), 
        .A(n6707), .ZN(n6710) );
  NOR4_X1 U7702 ( .A1(n6713), .A2(n6712), .A3(n6711), .A4(n6710), .ZN(n6747)
         );
  INV_X1 U7703 ( .A(INSTQUEUE_REG_5__7__SCAN_IN), .ZN(n6715) );
  AOI22_X1 U7704 ( .A1(n6716), .A2(keyinput127), .B1(n6715), .B2(keyinput41), 
        .ZN(n6714) );
  OAI221_X1 U7705 ( .B1(n6716), .B2(keyinput127), .C1(n6715), .C2(keyinput41), 
        .A(n6714), .ZN(n6729) );
  AOI22_X1 U7706 ( .A1(n6719), .A2(keyinput74), .B1(keyinput100), .B2(n6718), 
        .ZN(n6717) );
  OAI221_X1 U7707 ( .B1(n6719), .B2(keyinput74), .C1(n6718), .C2(keyinput100), 
        .A(n6717), .ZN(n6728) );
  INV_X1 U7708 ( .A(DATAO_REG_9__SCAN_IN), .ZN(n6721) );
  AOI22_X1 U7709 ( .A1(n6722), .A2(keyinput90), .B1(keyinput105), .B2(n6721), 
        .ZN(n6720) );
  OAI221_X1 U7710 ( .B1(n6722), .B2(keyinput90), .C1(n6721), .C2(keyinput105), 
        .A(n6720), .ZN(n6727) );
  INV_X1 U7711 ( .A(INSTQUEUE_REG_6__0__SCAN_IN), .ZN(n6724) );
  AOI22_X1 U7712 ( .A1(n6725), .A2(keyinput18), .B1(n6724), .B2(keyinput116), 
        .ZN(n6723) );
  OAI221_X1 U7713 ( .B1(n6725), .B2(keyinput18), .C1(n6724), .C2(keyinput116), 
        .A(n6723), .ZN(n6726) );
  NOR4_X1 U7714 ( .A1(n6729), .A2(n6728), .A3(n6727), .A4(n6726), .ZN(n6746)
         );
  INV_X1 U7715 ( .A(CODEFETCH_REG_SCAN_IN), .ZN(n6732) );
  AOI22_X1 U7716 ( .A1(n6732), .A2(keyinput36), .B1(n6731), .B2(keyinput3), 
        .ZN(n6730) );
  OAI221_X1 U7717 ( .B1(n6732), .B2(keyinput36), .C1(n6731), .C2(keyinput3), 
        .A(n6730), .ZN(n6744) );
  AOI22_X1 U7718 ( .A1(n6735), .A2(keyinput68), .B1(n6734), .B2(keyinput27), 
        .ZN(n6733) );
  OAI221_X1 U7719 ( .B1(n6735), .B2(keyinput68), .C1(n6734), .C2(keyinput27), 
        .A(n6733), .ZN(n6743) );
  AOI22_X1 U7720 ( .A1(n6738), .A2(keyinput123), .B1(keyinput5), .B2(n6737), 
        .ZN(n6736) );
  OAI221_X1 U7721 ( .B1(n6738), .B2(keyinput123), .C1(n6737), .C2(keyinput5), 
        .A(n6736), .ZN(n6742) );
  NOR4_X1 U7722 ( .A1(n6744), .A2(n6743), .A3(n6742), .A4(n6741), .ZN(n6745)
         );
  NAND4_X1 U7723 ( .A1(n6748), .A2(n6747), .A3(n6746), .A4(n6745), .ZN(n6948)
         );
  INV_X1 U7724 ( .A(D_C_N_REG_SCAN_IN), .ZN(n6750) );
  AOI22_X1 U7725 ( .A1(n6751), .A2(keyinput21), .B1(keyinput38), .B2(n6750), 
        .ZN(n6749) );
  OAI221_X1 U7726 ( .B1(n6751), .B2(keyinput21), .C1(n6750), .C2(keyinput38), 
        .A(n6749), .ZN(n6764) );
  INV_X1 U7727 ( .A(INSTQUEUE_REG_14__5__SCAN_IN), .ZN(n6754) );
  INV_X1 U7728 ( .A(INSTQUEUE_REG_5__2__SCAN_IN), .ZN(n6753) );
  AOI22_X1 U7729 ( .A1(n6754), .A2(keyinput26), .B1(keyinput50), .B2(n6753), 
        .ZN(n6752) );
  OAI221_X1 U7730 ( .B1(n6754), .B2(keyinput26), .C1(n6753), .C2(keyinput50), 
        .A(n6752), .ZN(n6763) );
  AOI22_X1 U7731 ( .A1(n6757), .A2(keyinput24), .B1(n6756), .B2(keyinput48), 
        .ZN(n6755) );
  OAI221_X1 U7732 ( .B1(n6757), .B2(keyinput24), .C1(n6756), .C2(keyinput48), 
        .A(n6755), .ZN(n6762) );
  AOI22_X1 U7733 ( .A1(n6760), .A2(keyinput93), .B1(n6759), .B2(keyinput34), 
        .ZN(n6758) );
  OAI221_X1 U7734 ( .B1(n6760), .B2(keyinput93), .C1(n6759), .C2(keyinput34), 
        .A(n6758), .ZN(n6761) );
  NOR4_X1 U7735 ( .A1(n6764), .A2(n6763), .A3(n6762), .A4(n6761), .ZN(n6811)
         );
  AOI22_X1 U7736 ( .A1(n6767), .A2(keyinput83), .B1(keyinput43), .B2(n6766), 
        .ZN(n6765) );
  OAI221_X1 U7737 ( .B1(n6767), .B2(keyinput83), .C1(n6766), .C2(keyinput43), 
        .A(n6765), .ZN(n6778) );
  AOI22_X1 U7738 ( .A1(n6770), .A2(keyinput13), .B1(n6769), .B2(keyinput73), 
        .ZN(n6768) );
  OAI221_X1 U7739 ( .B1(n6770), .B2(keyinput13), .C1(n6769), .C2(keyinput73), 
        .A(n6768), .ZN(n6777) );
  AOI22_X1 U7740 ( .A1(n6772), .A2(keyinput120), .B1(n5897), .B2(keyinput96), 
        .ZN(n6771) );
  OAI221_X1 U7741 ( .B1(n6772), .B2(keyinput120), .C1(n5897), .C2(keyinput96), 
        .A(n6771), .ZN(n6776) );
  XOR2_X1 U7742 ( .A(n4536), .B(keyinput86), .Z(n6774) );
  XNOR2_X1 U7743 ( .A(INSTQUEUERD_ADDR_REG_3__SCAN_IN), .B(keyinput0), .ZN(
        n6773) );
  NAND2_X1 U7744 ( .A1(n6774), .A2(n6773), .ZN(n6775) );
  NOR4_X1 U7745 ( .A1(n6778), .A2(n6777), .A3(n6776), .A4(n6775), .ZN(n6810)
         );
  AOI22_X1 U7746 ( .A1(n3780), .A2(keyinput103), .B1(keyinput69), .B2(n4806), 
        .ZN(n6779) );
  OAI221_X1 U7747 ( .B1(n3780), .B2(keyinput103), .C1(n4806), .C2(keyinput69), 
        .A(n6779), .ZN(n6792) );
  AOI22_X1 U7748 ( .A1(n6782), .A2(keyinput47), .B1(n6781), .B2(keyinput72), 
        .ZN(n6780) );
  OAI221_X1 U7749 ( .B1(n6782), .B2(keyinput47), .C1(n6781), .C2(keyinput72), 
        .A(n6780), .ZN(n6791) );
  AOI22_X1 U7750 ( .A1(n6785), .A2(keyinput119), .B1(keyinput53), .B2(n6784), 
        .ZN(n6783) );
  OAI221_X1 U7751 ( .B1(n6785), .B2(keyinput119), .C1(n6784), .C2(keyinput53), 
        .A(n6783), .ZN(n6790) );
  INV_X1 U7752 ( .A(INSTQUEUE_REG_7__6__SCAN_IN), .ZN(n6788) );
  AOI22_X1 U7753 ( .A1(n6788), .A2(keyinput78), .B1(keyinput106), .B2(n6787), 
        .ZN(n6786) );
  OAI221_X1 U7754 ( .B1(n6788), .B2(keyinput78), .C1(n6787), .C2(keyinput106), 
        .A(n6786), .ZN(n6789) );
  NOR4_X1 U7755 ( .A1(n6792), .A2(n6791), .A3(n6790), .A4(n6789), .ZN(n6809)
         );
  INV_X1 U7756 ( .A(EAX_REG_31__SCAN_IN), .ZN(n6794) );
  AOI22_X1 U7757 ( .A1(n6795), .A2(keyinput17), .B1(n6794), .B2(keyinput20), 
        .ZN(n6793) );
  OAI221_X1 U7758 ( .B1(n6795), .B2(keyinput17), .C1(n6794), .C2(keyinput20), 
        .A(n6793), .ZN(n6807) );
  AOI22_X1 U7759 ( .A1(n6798), .A2(keyinput66), .B1(n6797), .B2(keyinput80), 
        .ZN(n6796) );
  OAI221_X1 U7760 ( .B1(n6798), .B2(keyinput66), .C1(n6797), .C2(keyinput80), 
        .A(n6796), .ZN(n6806) );
  INV_X1 U7761 ( .A(INSTQUEUE_REG_7__7__SCAN_IN), .ZN(n6800) );
  AOI22_X1 U7762 ( .A1(n6801), .A2(keyinput89), .B1(keyinput101), .B2(n6800), 
        .ZN(n6799) );
  OAI221_X1 U7763 ( .B1(n6801), .B2(keyinput89), .C1(n6800), .C2(keyinput101), 
        .A(n6799), .ZN(n6805) );
  AOI22_X1 U7764 ( .A1(n6803), .A2(keyinput56), .B1(keyinput99), .B2(n5637), 
        .ZN(n6802) );
  OAI221_X1 U7765 ( .B1(n6803), .B2(keyinput56), .C1(n5637), .C2(keyinput99), 
        .A(n6802), .ZN(n6804) );
  NOR4_X1 U7766 ( .A1(n6807), .A2(n6806), .A3(n6805), .A4(n6804), .ZN(n6808)
         );
  NAND4_X1 U7767 ( .A1(n6811), .A2(n6810), .A3(n6809), .A4(n6808), .ZN(n6947)
         );
  AOI22_X1 U7768 ( .A1(n6814), .A2(keyinput37), .B1(keyinput35), .B2(n6813), 
        .ZN(n6812) );
  OAI221_X1 U7769 ( .B1(n6814), .B2(keyinput37), .C1(n6813), .C2(keyinput35), 
        .A(n6812), .ZN(n6826) );
  INV_X1 U7770 ( .A(DATAWIDTH_REG_0__SCAN_IN), .ZN(n6817) );
  AOI22_X1 U7771 ( .A1(n6817), .A2(keyinput8), .B1(keyinput110), .B2(n6816), 
        .ZN(n6815) );
  OAI221_X1 U7772 ( .B1(n6817), .B2(keyinput8), .C1(n6816), .C2(keyinput110), 
        .A(n6815), .ZN(n6825) );
  AOI22_X1 U7773 ( .A1(n4849), .A2(keyinput94), .B1(keyinput79), .B2(n6819), 
        .ZN(n6818) );
  OAI221_X1 U7774 ( .B1(n4849), .B2(keyinput94), .C1(n6819), .C2(keyinput79), 
        .A(n6818), .ZN(n6824) );
  AOI22_X1 U7775 ( .A1(n6822), .A2(keyinput115), .B1(keyinput32), .B2(n6821), 
        .ZN(n6820) );
  OAI221_X1 U7776 ( .B1(n6822), .B2(keyinput115), .C1(n6821), .C2(keyinput32), 
        .A(n6820), .ZN(n6823) );
  NOR4_X1 U7777 ( .A1(n6826), .A2(n6825), .A3(n6824), .A4(n6823), .ZN(n6877)
         );
  INV_X1 U7778 ( .A(DATAO_REG_4__SCAN_IN), .ZN(n6829) );
  AOI22_X1 U7779 ( .A1(n6829), .A2(keyinput125), .B1(n6828), .B2(keyinput76), 
        .ZN(n6827) );
  OAI221_X1 U7780 ( .B1(n6829), .B2(keyinput125), .C1(n6828), .C2(keyinput76), 
        .A(n6827), .ZN(n6842) );
  AOI22_X1 U7781 ( .A1(n6832), .A2(keyinput85), .B1(keyinput84), .B2(n6831), 
        .ZN(n6830) );
  OAI221_X1 U7782 ( .B1(n6832), .B2(keyinput85), .C1(n6831), .C2(keyinput84), 
        .A(n6830), .ZN(n6841) );
  INV_X1 U7783 ( .A(DATAI_14_), .ZN(n6834) );
  AOI22_X1 U7784 ( .A1(n6835), .A2(keyinput54), .B1(keyinput59), .B2(n6834), 
        .ZN(n6833) );
  OAI221_X1 U7785 ( .B1(n6835), .B2(keyinput54), .C1(n6834), .C2(keyinput59), 
        .A(n6833), .ZN(n6840) );
  AOI22_X1 U7786 ( .A1(n6838), .A2(keyinput104), .B1(n6837), .B2(keyinput61), 
        .ZN(n6836) );
  OAI221_X1 U7787 ( .B1(n6838), .B2(keyinput104), .C1(n6837), .C2(keyinput61), 
        .A(n6836), .ZN(n6839) );
  NOR4_X1 U7788 ( .A1(n6842), .A2(n6841), .A3(n6840), .A4(n6839), .ZN(n6876)
         );
  AOI22_X1 U7789 ( .A1(n6845), .A2(keyinput40), .B1(n6844), .B2(keyinput57), 
        .ZN(n6843) );
  OAI221_X1 U7790 ( .B1(n6845), .B2(keyinput40), .C1(n6844), .C2(keyinput57), 
        .A(n6843), .ZN(n6858) );
  AOI22_X1 U7791 ( .A1(n6848), .A2(keyinput71), .B1(keyinput88), .B2(n6847), 
        .ZN(n6846) );
  OAI221_X1 U7792 ( .B1(n6848), .B2(keyinput71), .C1(n6847), .C2(keyinput88), 
        .A(n6846), .ZN(n6857) );
  INV_X1 U7793 ( .A(INSTQUEUE_REG_1__5__SCAN_IN), .ZN(n6850) );
  AOI22_X1 U7794 ( .A1(n6851), .A2(keyinput14), .B1(n6850), .B2(keyinput12), 
        .ZN(n6849) );
  OAI221_X1 U7795 ( .B1(n6851), .B2(keyinput14), .C1(n6850), .C2(keyinput12), 
        .A(n6849), .ZN(n6856) );
  AOI22_X1 U7796 ( .A1(n6854), .A2(keyinput55), .B1(keyinput19), .B2(n6853), 
        .ZN(n6852) );
  OAI221_X1 U7797 ( .B1(n6854), .B2(keyinput55), .C1(n6853), .C2(keyinput19), 
        .A(n6852), .ZN(n6855) );
  NOR4_X1 U7798 ( .A1(n6858), .A2(n6857), .A3(n6856), .A4(n6855), .ZN(n6875)
         );
  INV_X1 U7799 ( .A(INSTQUEUE_REG_9__1__SCAN_IN), .ZN(n6860) );
  AOI22_X1 U7800 ( .A1(n6861), .A2(keyinput91), .B1(n6860), .B2(keyinput98), 
        .ZN(n6859) );
  OAI221_X1 U7801 ( .B1(n6861), .B2(keyinput91), .C1(n6860), .C2(keyinput98), 
        .A(n6859), .ZN(n6873) );
  AOI22_X1 U7802 ( .A1(n5893), .A2(keyinput107), .B1(n6863), .B2(keyinput75), 
        .ZN(n6862) );
  OAI221_X1 U7803 ( .B1(n5893), .B2(keyinput107), .C1(n6863), .C2(keyinput75), 
        .A(n6862), .ZN(n6872) );
  AOI22_X1 U7804 ( .A1(n6866), .A2(keyinput2), .B1(n6865), .B2(keyinput10), 
        .ZN(n6864) );
  OAI221_X1 U7805 ( .B1(n6866), .B2(keyinput2), .C1(n6865), .C2(keyinput10), 
        .A(n6864), .ZN(n6871) );
  AOI22_X1 U7806 ( .A1(n6869), .A2(keyinput23), .B1(n6868), .B2(keyinput22), 
        .ZN(n6867) );
  OAI221_X1 U7807 ( .B1(n6869), .B2(keyinput23), .C1(n6868), .C2(keyinput22), 
        .A(n6867), .ZN(n6870) );
  NOR4_X1 U7808 ( .A1(n6873), .A2(n6872), .A3(n6871), .A4(n6870), .ZN(n6874)
         );
  NAND4_X1 U7809 ( .A1(n6877), .A2(n6876), .A3(n6875), .A4(n6874), .ZN(n6946)
         );
  AOI22_X1 U7810 ( .A1(n6880), .A2(keyinput112), .B1(keyinput81), .B2(n6879), 
        .ZN(n6878) );
  OAI221_X1 U7811 ( .B1(n6880), .B2(keyinput112), .C1(n6879), .C2(keyinput81), 
        .A(n6878), .ZN(n6892) );
  INV_X1 U7812 ( .A(INSTQUEUE_REG_13__6__SCAN_IN), .ZN(n6882) );
  AOI22_X1 U7813 ( .A1(n6882), .A2(keyinput118), .B1(keyinput44), .B2(n3627), 
        .ZN(n6881) );
  OAI221_X1 U7814 ( .B1(n6882), .B2(keyinput118), .C1(n3627), .C2(keyinput44), 
        .A(n6881), .ZN(n6891) );
  INV_X1 U7815 ( .A(INSTQUEUE_REG_1__4__SCAN_IN), .ZN(n6884) );
  AOI22_X1 U7816 ( .A1(n6885), .A2(keyinput82), .B1(n6884), .B2(keyinput46), 
        .ZN(n6883) );
  OAI221_X1 U7817 ( .B1(n6885), .B2(keyinput82), .C1(n6884), .C2(keyinput46), 
        .A(n6883), .ZN(n6890) );
  AOI22_X1 U7818 ( .A1(n6888), .A2(keyinput33), .B1(n6887), .B2(keyinput113), 
        .ZN(n6886) );
  OAI221_X1 U7819 ( .B1(n6888), .B2(keyinput33), .C1(n6887), .C2(keyinput113), 
        .A(n6886), .ZN(n6889) );
  NOR4_X1 U7820 ( .A1(n6892), .A2(n6891), .A3(n6890), .A4(n6889), .ZN(n6944)
         );
  AOI22_X1 U7821 ( .A1(n6895), .A2(keyinput45), .B1(keyinput49), .B2(n6894), 
        .ZN(n6893) );
  OAI221_X1 U7822 ( .B1(n6895), .B2(keyinput45), .C1(n6894), .C2(keyinput49), 
        .A(n6893), .ZN(n6899) );
  XNOR2_X1 U7823 ( .A(n6896), .B(keyinput6), .ZN(n6898) );
  XNOR2_X1 U7824 ( .A(n3258), .B(keyinput9), .ZN(n6897) );
  OR3_X1 U7825 ( .A1(n6899), .A2(n6898), .A3(n6897), .ZN(n6908) );
  INV_X1 U7826 ( .A(INSTQUEUE_REG_4__1__SCAN_IN), .ZN(n6901) );
  AOI22_X1 U7827 ( .A1(n6902), .A2(keyinput25), .B1(n6901), .B2(keyinput114), 
        .ZN(n6900) );
  OAI221_X1 U7828 ( .B1(n6902), .B2(keyinput25), .C1(n6901), .C2(keyinput114), 
        .A(n6900), .ZN(n6907) );
  INV_X1 U7829 ( .A(PHYADDRPOINTER_REG_14__SCAN_IN), .ZN(n6904) );
  AOI22_X1 U7830 ( .A1(n6905), .A2(keyinput1), .B1(n6904), .B2(keyinput16), 
        .ZN(n6903) );
  OAI221_X1 U7831 ( .B1(n6905), .B2(keyinput1), .C1(n6904), .C2(keyinput16), 
        .A(n6903), .ZN(n6906) );
  NOR3_X1 U7832 ( .A1(n6908), .A2(n6907), .A3(n6906), .ZN(n6943) );
  AOI22_X1 U7833 ( .A1(n6911), .A2(keyinput30), .B1(keyinput42), .B2(n6910), 
        .ZN(n6909) );
  OAI221_X1 U7834 ( .B1(n6911), .B2(keyinput30), .C1(n6910), .C2(keyinput42), 
        .A(n6909), .ZN(n6924) );
  INV_X1 U7835 ( .A(DATAO_REG_3__SCAN_IN), .ZN(n6913) );
  AOI22_X1 U7836 ( .A1(n6914), .A2(keyinput28), .B1(keyinput124), .B2(n6913), 
        .ZN(n6912) );
  OAI221_X1 U7837 ( .B1(n6914), .B2(keyinput28), .C1(n6913), .C2(keyinput124), 
        .A(n6912), .ZN(n6923) );
  INV_X1 U7838 ( .A(PHYADDRPOINTER_REG_0__SCAN_IN), .ZN(n6917) );
  AOI22_X1 U7839 ( .A1(n6917), .A2(keyinput67), .B1(n6916), .B2(keyinput39), 
        .ZN(n6915) );
  OAI221_X1 U7840 ( .B1(n6917), .B2(keyinput67), .C1(n6916), .C2(keyinput39), 
        .A(n6915), .ZN(n6922) );
  INV_X1 U7841 ( .A(INSTQUEUE_REG_12__5__SCAN_IN), .ZN(n6920) );
  AOI22_X1 U7842 ( .A1(n6920), .A2(keyinput52), .B1(keyinput15), .B2(n6919), 
        .ZN(n6918) );
  OAI221_X1 U7843 ( .B1(n6920), .B2(keyinput52), .C1(n6919), .C2(keyinput15), 
        .A(n6918), .ZN(n6921) );
  NOR4_X1 U7844 ( .A1(n6924), .A2(n6923), .A3(n6922), .A4(n6921), .ZN(n6942)
         );
  AOI22_X1 U7845 ( .A1(n6927), .A2(keyinput111), .B1(keyinput108), .B2(n6926), 
        .ZN(n6925) );
  OAI221_X1 U7846 ( .B1(n6927), .B2(keyinput111), .C1(n6926), .C2(keyinput108), 
        .A(n6925), .ZN(n6940) );
  AOI22_X1 U7847 ( .A1(n6930), .A2(keyinput58), .B1(keyinput7), .B2(n6929), 
        .ZN(n6928) );
  OAI221_X1 U7848 ( .B1(n6930), .B2(keyinput58), .C1(n6929), .C2(keyinput7), 
        .A(n6928), .ZN(n6939) );
  AOI22_X1 U7849 ( .A1(n6933), .A2(keyinput11), .B1(n6932), .B2(keyinput4), 
        .ZN(n6931) );
  OAI221_X1 U7850 ( .B1(n6933), .B2(keyinput11), .C1(n6932), .C2(keyinput4), 
        .A(n6931), .ZN(n6938) );
  AOI22_X1 U7851 ( .A1(n6936), .A2(keyinput62), .B1(n6935), .B2(keyinput64), 
        .ZN(n6934) );
  OAI221_X1 U7852 ( .B1(n6936), .B2(keyinput62), .C1(n6935), .C2(keyinput64), 
        .A(n6934), .ZN(n6937) );
  NOR4_X1 U7853 ( .A1(n6940), .A2(n6939), .A3(n6938), .A4(n6937), .ZN(n6941)
         );
  NAND4_X1 U7854 ( .A1(n6944), .A2(n6943), .A3(n6942), .A4(n6941), .ZN(n6945)
         );
  NOR4_X1 U7855 ( .A1(n6948), .A2(n6947), .A3(n6946), .A4(n6945), .ZN(n6949)
         );
  XNOR2_X1 U7856 ( .A(n6950), .B(n6949), .ZN(n6964) );
  OAI22_X1 U7857 ( .A1(n6954), .A2(n6953), .B1(n6952), .B2(n6951), .ZN(n6955)
         );
  INV_X1 U7858 ( .A(n6955), .ZN(n6960) );
  AOI22_X1 U7859 ( .A1(INSTQUEUE_REG_9__1__SCAN_IN), .A2(n6958), .B1(n6957), 
        .B2(n6956), .ZN(n6959) );
  OAI211_X1 U7860 ( .C1(n6962), .C2(n6961), .A(n6960), .B(n6959), .ZN(n6963)
         );
  XNOR2_X1 U7861 ( .A(n6964), .B(n6963), .ZN(U3093) );
  CLKBUF_X1 U6031 ( .A(n4952), .Z(n4953) );
endmodule

